`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THTNEVnl8SALHKCB+oxzBUTqcXqI/FmN7+4IOPrbZrE0ELHJsD91ko6doh56Ha+0
I3DOeydpvpeQ2tGKb0kFxD0ozLmZ9ES3p2NaAoLA+KP+vVUYD1ox9yb4MC9pGheD
XeEBwAzWDwztzImkqJwMTiBhpn+2cP1B6DBPlXzLhIBW5RBpGwOdUD922NBS3Cxg
Zygw515u5xfaYjXsENrIBwo4+L1BboRvZPsVh062roT4NdOCto1Dv5JeqWufsemO
DV8NscCYjGzga9s6LoKTKZqNxAYZAwNyuxHWGniBrx0kPwA8xFoG7FqCFbG+0Na+
F7g2CW8ABerMve2KbcZDC7AGXWcCzAWkntR8jZ6ZhzcaExvSbcgEXW8fBBxQQJe1
7zTkXqLpKRk+fUeOilTlqbmE4KAqtNZzEttZG7EUEJQVyCi8kJyR9ooyPkeJAM7T
KvEX1Dzc5RVxjT6cY/38beg+BE6H5XzsOjkv4dG8sz0=
`protect END_PROTECTED
