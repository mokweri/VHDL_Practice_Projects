`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A/8KE9BbUncxkPuk0dzJx7OyhuptWQwX3wqpZkeIBjcRK/a4rqsT2bbzgbOXX0mf
HXxLDin/ZZdEWVQ9rVusC3OstBFAeON+eKA1Pl5wZa9Bz84ONlIXlPK/spNuvy6o
z2EU2RDJejRP+TpHTxIfqrNx2StObDEgKr/KZF4PzlW3DKTP+HlXM84gzh9LQ++6
9SVYNL9L85xgG2TX0Mi5Z4iTOzLoizfMkYJRP2UgtJ3ecCRlCfPOnd+nmyS1487S
5PwFGmTtKtEaV4x9cPX0ir3m763ZZhDI5twtjFE0BJzxI+fTM1kIIXaCjhmq1cop
tJdsyZ6G4v2OhTbnm+cZVQ4zDbCpagiSXE2A7oUsyBB1YVVbxkx1Yeu/x+D9rWwh
KPViFgskOSJn9jfWdRA1ZIiFB0T0k5RSeQv5AVQ9KQAAB1GNGWzRUPq4x0UNutBx
UQ4RLRHnJLWphebjhW7cgn68HfjKyptuPluUUdbbDQ7vyGnfbZ4iytSC+dkN35us
PRDHqyaaHkgoEJkX/A5ytqQsobkLz/PiXYr/b6Dylnaoy3aJXIkc9vYc0wfXAe8a
wXBX0tRsW04wTQ6Cs5sfT00c0mY1Lvh7ukiL3zS6pVt5EYWeH/mo+35jA0A98azx
cg20BMAtzg/P/nRtbEq5kspSTFZqexSktctqrJ4a+sP61XMRFkvG1IWmKXJSR38G
1L0cHt68SKMJWuh3i+NcNBjWkfQkfkMP7e0op8D3sE7lj4C568htYkX0d/lIZJmt
Rptb0+eernGqnEseygTa92lXk5mil+mKEUCZrlJnsANWex9NGtftkoeKl5TDhRfb
SGTEgP7du8+kldNmRCw4gguv3Sdd/8Wadj55MWg7prCpLEtchNByPrznVNisgmgX
AzqSctvhtD2YSbBhKuT8TXi4TVGFFeZBi+Tt19K8rirJTscWv13v7d/J7/hzUitv
4l0BLQ2HnbmpK+xlC0ArVc4orZ3tTdzcAfe+KXw4iY58TP5xuh/CSaTUaZOxI6ql
vbe8vvXVuwW/dQ0zr6Uy8cMdcrRqI1bMjxZb+rNPY+FOv/L1VPyY2ekYKYbaQrmj
nO4+ib33xqdfSN6TgscqeZb0BcMCw3FZ1Fqmh/to1n3zht/ooRW/HXUiLK6bsAGP
3y/SotJ4AlahkU1DczbXY6yOtX+F7fibo0580wOE7EvvBY1adM7KDDx8pmWhHdTD
qkA4VNyJoWgbFPRLD+G53rvRelgSLcOP2HyxLFCyRmh5X453q6Jd3xXme4QijYmj
sBTP/LtkgAoJyl7lyCk1U9d6TG1rLpVu2BujCH1wRL4Tf7KkHGtnWO91efnr23cv
Tf+YgjweLMVMPrCr5AIhVED4V1ry2GMubox24/7WnNQVndGlQgmFvQqXo0uLqZfU
+RyGW4q7iPQadubgOO8L+VApO3oWtnPyjW7HrlhHN38THe8y1My8xb1O1DeQnXnD
hNW+wrQlYZikw8Zw7C1OvIGpm2nij+hEjzquRF1sqThYlPXUFB/C29oLfE4u1OZa
vYrvzIiUzqdwDVRiCwON9SsV2y4C9Gww21yeAgrqIS2a6tpeYPbud9W5umUqE+hW
YCPGuyjr6v8HGHZigzm7Ij1enZoUgCHYi74eExSL7MKaiVt7uFqP9jd8ah5oR4Zf
LIw5Rv+jgU+TxPGlprbQyl4+qctNOgZiDTM1U2+y85YDagRDlbX0KAckR75csvmg
wxRUOQqPUalrREcwDHF3O4nnk0hVjo+4a0j4qj2xHhDrZj6ZvC6tIF9uQ1ntwgbv
ooJhn0TaPIbqzImA6JCL0ZYPokbXms9wovU7WwTax4wJIVfVfOqmII+D+FEKt2dB
r+w4FOY3VQlq2mYG1hNoA7YGmRL5DrwgQwbncLV1/SdKpbPI7m3SZugsXwH9Q3Wu
qsHuk5kNxGn5qs0yX9JgfJcC4Vzsbr18RiguQFB1Euq1htkOVG4r+i2nvlHgXJxQ
VJsQDRzKOh1lmWgaT3rAcjZ/0UYRNo2perp2IANbm/C7fibzvnqEOL671ocDiKv1
nT5mXN9L4bM1JFqSDX2Q0cGXJn+t9Rhx7dvOzicrvdSyTkZlkam03kkOzcQdHNAs
SM+M+hOfGcX5QL2eOOtb2OveILjxbPCZqEgDonGSb1BDi9LfPt23BtUjC9ivZCET
eSiGka4py1cY0ZtMIsEWu7ab1gefuq4WD6vYI2W2y+XxMR+rHjZFfMNnLdxWg9Lz
6l4z9zbGvA17NbL3FphHTl1GerkTdrgTuPoN5g4B0q5/8mfWdpQXyIxmG4/dbAEB
0iI9wXFKNfu1IyxWWwOWN3WrEjOIR0lViDYi3CfuH7WijkvYDzVy6bOZ7iTq0NfS
claL7k9Erz4o5dA0zumQsI7kfhgtVkd3qomkltRcu3XR9G6Eunu7qxChsvKaDKTn
JCGaMdVwI2U7tz+68MLz2eBtynG5N3hH3UaF6cgHV/FYaMP6BfNy6I8qSjwsApko
4mys/nrQ68K3YkUmDrr+4Y8iI1t2asOxgKb5Fzic/4Wc/ebcOzwtlzDgy0u9Uqzy
Zoqh8oEKqTbEuenARkHUB6wgWz1wILgBf56QaYKeUr6dfQ0tpLqvo5uzylq7tTqs
FY4wTjoEyBqpNaWA7NP7dth4of1aRdFHqGHbNQUuwZfAUbl1iiX9SaMvlKiTvHlr
hHnDJaaq/bkmh/LwGN80fHyDg03HJeOjdS3fYHyUH/+JXgL1fKrWrkKuE5eyKKaz
zSKAahcZEJEks57cZvTxThuH7YULgt9JIN4jVXzUnLtT6ikxeXlIiQGNFnFWmrZO
Pv3ku1kR99kGxYYBeUPWtikd3ELeg68fRbXstugTWfZl0gZ8MIzPBZUTIYtfHYlo
F4dTea2shJfgquX/BvEI6/sQUGHjd4yHVc/PKxVhLkE4VCNC2SIesg1Fu30H8K7k
QP1SGs/CxfqRZF2CEeZB6GI+f1OTaOMB7XzbOLu6y7zXGXOOwEv07Zir2CBdt1km
4fpvCVz7zh/sn9RR0wW0iG4ebJVEpbKpX2wLNOy2g41gJpJhSb0Z+K1nezPy9EZP
YzJWCY2+txg6tjkl3Q6fwX2EFHJc8JXchDIrDDmYTiLunMHuFwc+L6wdU3C8z5LQ
YkjL8Rq+7rUObzNM2dL0htq6yH98nI4C/B1XP11dv48G+7BNuSKcudYbXfTsqjL7
mA9ayR+Sr5IF5laM9w6b02kKyNfsbfi5FbZ8t+k3pYUh7w21U2TcOy854zSuMcM6
owDn9+AQs2dOgEwfuSktSBbjI/U7IGGOGb3rxMSt6twqxjq8CEY6EfqZrGnABnih
6oc7e557e9S3im7R9mp5CnIl9Bb8TST5Sw7uqvuS0610jBhuMnad8BNQelxXrXy1
dl8wLi6xd1ACmOs9Ign2TOXn4E3N2JsvQ7ECfB3f+tvB1WF3ArOutnZUBaENyBaY
43hDXj370xcOcIbMx9qGD08UBCAyBvH6YqvhxzWwp4+zYNwlsOWJq8MX/iWq/zZi
egZ8SVssEB2jHhveJVrALVGdRIuTHynkqhZAaBAhiJnDTsMOh6bG72586+/ruJQd
s4p3Z8OJksAt3LhXZVjGFNiW9m/UlOBOr/ZaFSn/RGqB29MwQBOL6Zeo8Hu7VbfA
W6fK6EMsh1KpcQ4QiUOaD6pzikGf06rpVVJTyVr5aNXXi0rnBdiDevUg4QTRxA5K
McTX6KvltVbBPjYQIsvA8niF8V4qPYQI5M8d3dtF1N7X+Y4dhJ3H6lKXxQbbPM+K
dT3TQc7bBE2OvvPHs9fRkH+B6OGG6mraBgx10+1jow5Xe3vNAQApERIOWeNTSpZP
dgVVelLa2fr1529xmtCGvv0/IMNAkJfSnJwrK7k5pocegLwT5cAyn202vhcJqY3h
DZNFFf9KPz5jYDN9g2tgnKhWycFWUPvxhmoCoOjW4nQbtJ1gqxTGTqKf36nILMSI
FqGLeT7m9IVbl/BmfRDdg2JPMkEyEW5E6bwVtBA79rALpAANTEpg9+pYEeDZFzPH
zg2aP22qiDUpppMNbhqL+8Np8y09f15luOSHI+MyfY2yTwzCyE3V8gMoOieQmrY4
kou9FeEaAnpzP6ao3mpsfo80ZssV4G2p5fFQS/D/bzOSEczedxs0JtlAtOuzA7Ra
2qBW9P6H7Z9aJRPIy8CzW61UsgzfK4NhoEIdtEIC7o94tp01O9GO0fWKrZoQeomV
gU7a/9KFyNyEq4Isrs+7YlBKuRG7AIszTC6h+8J1zFHvVaAhPwKyDbH2dv2q/FkQ
rVe+sQhOdZ66zYobe9u6kMKq3R7DK/RRTlurSZPGmBFM291saigPCb3yJx+9k+mf
8BtZMihnn2nKWG0w+Kj7ZY6sefg5QhTYL9fzb0bFIfzhoJymA021hMnuHO4Q0m0E
4rhvl/rQCmEKpNez9G8/gyQZfdd/ztiSxr5vUU2o+g5D5RyriZeoqTT5UHLzPKqa
+hzOJ4b2fpStjRzIqvcsh6RDgMKFMR5mGjgsjXZslPObX0zW/t34RnK84GkPOX6G
U6QIVp1HhtCtsP2d8ZUQ7v4unvTV1m9fwiE7jfo4eEUJIZZSpxl1tfa0Sbyp+30r
2/ZHtsDdCdndfGAc9hYAWfoWulgr6g0bzG+/+OadLm2GyyPnzYFXf+DdOUsXF6KO
j+zmqHXYMVzlbqFc+/kJI6v1nKuxNw+3SYp464QjEFRu6yUB6A4F8h1wKtd0zO6O
9CMKCpko3PEXhdgrJMOVPPDxQp9pcHJMIHPdZDFfYSuT1POedyh5tR5qa22Flxbl
W6frr22BxnHZh5AkElPU43sw2HM0mj+KjT7bR50ee1pl/BOsS6C4JxrKplwsuES8
d2cLzPw9TsGbXYuvPRIVei1ViPaohwcWQurnPSebsEd3gZqU/YY+PWxBmzbcJ3XF
HnLVilLx+v68cp853a6VPcP4jALdSrWWbhzKB0uICKKsfGK/UV6ip8Gavjhdch4V
3WwEU79LoLqXQai1npiF4bfwNAhuQIltMWKTqt4EVvra+FHxWce3NBU1DuLp1EjT
+QPC9oOSHnNRxexlsUuPrxiWlenKWaiMONdc6vkIPDkg5Meeg5b0li43jeKeXOIh
hCO7z1cno41gtyiCFm4sPK4sH8wAdmjNtBcMWVjHVkbNG5YT5PUTSf5CJpb/sWRV
OFBwN0P/95EDn5fqKk6T64uBqgBLmRmn7CZ5bPbsxbi9dqZbI/7DXrA8BywDOtqw
X94NE/FXvLY6YZl5v5zL9rEJw83+q5aasjjTgUUe9YFvLgFyql3YYqqxxtY3C4xn
IwYBrZdFxV85CIZQbOYk/OkRdMLBjOAbtJdGUp2ahtQOqjoZYLE0Yx6CJW6qltiD
cCRKbmDPh259M3l4vDx8ZQQXU2kTgCauOvTovGyqf8X8qj2cgBtzAa1UlGUNQrJT
dpXIVL3OX28t4h5xP36ylx5Fhq9PHeJ8KlLZB9EBjTeJuL2AY3Gqz47WI0Y4O2yg
PAJtKV6fNT+gNaFEVdsStZFMP1aY9bxw2anZTdn6pGxqKHfdbYqEMAL0BO5U90Zv
PbfI8WjcFl+xopmpCTCVXNZYzQg3QTGU6qg5WzXucJyjs3JRFcaAaZJ2r6frOmFZ
0m01vy9Oz7SZyuVbF6+4LwPKX4Xi37h7tA3+C5xLlHESUub6acCbPj1RaF5aRVB5
ydtrn8tEUYIhmXLRWxkURE7JIAueJzZI2N3Ac7anAXvgfZuE7ehU/pve9S61doBk
EvkPXdcB3s8nYBl7bQotQHy+lRnmDiagn3jw0ZfpRacpWr9OjcCKbZ938oofhXhG
ns9WSer2EPw9ayiHMrfEAFjMefhM5sX5DEM2nF9HberGVOJCR2O+teYv7ZtQxHn0
hkXplbdwErFUblzJ2KUOxlMV+MKSahPN5gXQXUmnZNSPC6dZBu5w4mC1sONM+S9P
bgqUvE/ezlrg6yrRTq8tMBFEyJUnxLimcijVfAw9yfwn02e3WkNqHzeKKWXy9HBz
5+HtB0HpUQySasry5XEG9I3t1Vk/WBeiSWh5n2mFBKOnvwOVlQhrGJ0bAJcwj+lJ
/u4Bmm/dltbw/CGBXBMxoENitdGPNE9JsPTqgdHQ+Y5UI9sW6iDaG3cvmATohIGs
+/lEWsxI/4RiwVzHXSLNkNywikeX8zkRW1qKZfe+nVZ3xU4+H9qVmJcVvdDb4HKy
lQN4sZ/ANdPX+dU8p3VSnYdzUAfSzmpIDekF8Zin4YjIRQi1SAY9kf+iy8gXUa3R
AGO1oLMDEJLxjxRmt2tDvLX7rj3aM1DSDMOilmTWhBdoOt/QreAeZAnAHNVt7SDk
kOnM8hksXOUD2i12Y5vkfKhWZ7zbEmzsuBVUd/ePgCTJ9cPn/usk2321egF/mERb
FM6qazHCYf7muRu9AjmdBo61CUgqtPDaz0073Hvi4F+3/eA2HDJ0NEAQG0amkG6w
rVBXdN2RPmW8c3yzN8j9jI5lzdmaZ3VBsZ6V2SdORvO7yxo9ucx8ISwsRQM8AmPt
kS/ziG6B+pX0sGUtulL2GpwbN5ltYfgDG751ba4ROjaO62iDC/QHx6Mh2/vXZPo9
sO8cL1Ysof4IRi2NFJgW7Nm1dqgv9s99JdH14idZCLG42FoDaY2444YHKryfk4t1
uDyLdQ6SNTdFBuorDkdqID0MhqASfTnKqq6D8P0fRlgNHs8Ep5pkc1pW9++YDc0L
OfS1NjbDrKbq1GjW1NAYJ/S5P3jGOUP/+gPeM9PFL9GcZLyeMxtBW8Jj4mJACd1f
1Bezzhe18Q1pkxY0RaGV/a/x+UPm/L40gEmNAQRJJLCBeqOJ/51E1pbR4YvYsw0j
F7bA99uZTzf4wpkRdJMXJqz0629AIbvNxtdmeFcPkNH69haLIQ+rLK24EThxZMFu
mlypocPhi5m86BOaFH7502602cFBrGq6g5X6RhD8+bkOf8sFqKMRBf8KcrClHiBX
VJpC4TsBHfR4gbOR0IH1KWO14wlIrM2w1UZS+P9XsdMM2vDspZVOaoJLXHNND7bd
d1D0EC9wXVnB1T35DobPcdS/aHiR/tklJZEGmkLT5ot7eamHWJ/ve2qT7lHB/UwC
cmiLvcYbh15CfU+fWNV0PjtLlLsxf9IiseiBg0Zlk4HH8HlfKhWuN9oQq3Kes//U
KjqBQoqmQkYLfs7VUvQXeTVucgeDWe07OgDDW33SI5MM6sWIw9qABNRz0yrYwzvW
aM7KO4jjVk89aJOL4tI8D9NzzonMUAp4lwj6ue2xvspqyCMIIYBlI7P/CSbSa40i
HW13WwqwlSv3LPcnLo2i/b9CjPapzBCelG+uzPx9UEWfvknbVB1nrNk8qCG4slWU
jsDL3VK58lT5ShRo+FRkPLTrm7fhF0p53qkB5J1yRkpUTEGSQ99HlutOPZlmH/wf
Tw9HUZDRGuku7kkMhTks0LS/jDMfkR3vkvON/YvCMK1xgdSNCNJC1vBWykHyPYGC
Q5v3fJobt2eJCJqxsVbE7vvyNQCkWPs9HWiizzosChloPQ/DfwxBZ6cK6wkmH5bL
xkbWw5g56eM8vV7iw8KAnYQr4Keyszx1bAKvt4u87rhs7y5Scb3ph3++5HYBKv5o
OhtBpJXloMb7ZZ/DhkHn85xNuJEnhoEK1UPXBTd0af/Lb46+11dkIBDTZ9Su/AJj
uo2B4ifrn3UaY7Z7XyO1XWpZWiarl6S571Nr2bCNw1hOhmCMNc6SM5teWTYDXwG5
vwLTk4jRbCx80/cwFOFZkZev+HoTmECZz7Sxb9M6vpMDC6XR1IDQEJYAwyz+qYUw
kEXrhSvuhop9QC3dvI59DEVpkgWyx+VqV8n2TGoIqlb8o+EfvEzB/oWQm+ynRLmn
z5kQhndKi0mzvXDJz9MpE9LtsS/UsLnvm5vTVfEbeo54XiUwaubkNu2tHtf/Ppld
f+u74RcFplZWdqdbXB86ViDGQfNF5AnMRBj8fJIWZ/CPm530YNuF5aLOUGW8dadD
n6MCCvqqp8oyWVP5AozrF3o97rXd38FrgcXsS0WwHBlZx3yTEREYtKv750ODQh+C
NoWtaTiNPOQ3iZy7glxru72kE3zhkuqO/PxnilxoMRhe5MNSvzWb4KYCtC3p+CQH
F2C6uE9KbDNFOcYsfdoQh7T21DQdYo/c7HwNWQIrezHRJIeeD0yMEROOBt5pgmlA
j6gbVYIx/Df8bkToDjrzZBtz9iPkudccAp6/7jChCHrPedmYP6CAFQInVxpYQ34K
d/38jya03BSdAQWrsqrTRVNyNwS3L0ys2pMfYEjqW5MGTLHx/vIJnfYuj8i1ifIP
TtIZTG3RTXo31+sZkkTUYXwHrVicg8rRFdlQ+9VBfTD5jDw69LeIrDNtzqoQRkVe
3o2ZLTHKoHb5i7QvBkXAvpHgJpQyeo9fXDvFPqGYuWTWQkuYHiX08qD4YIqpNP+d
j94fJptQbaQ2MpFhWKQ2/9IPkmxyLb+XV2XiN7DC5jZzAfulSDBVo/AQ1V1oM3Wc
YvlJ5jh1VnnmMMHH1sjscdXzztk/PQ/7Mr9ZrCIySeABCrtJoS717VELXKpyCBWR
t7VmZzzDsSpbNv5s8ErbpmSORrjIUcyfMBGY5bBF/db6Of/Y5dvWdn04Xby5z6YV
XsDmuKFziSUxUpvHtWZYnFGlqwgNPf10CC6TTzzYilHnJCzpytN8OGcZkwqi17Qo
5NlIG3bz/6fqpFLF+14H7K42RWI616UXxuGjlMIT6MH1QJ9C99Yp/ctuL8p6u+5Z
L5VzfT1GZqMxMcsQI/6X7ln1mDR45GX8ppBXqiKIowsNDylm3RKfKxCxVAmWV1+x
EzzU80fsQExQPwlCJ+1TsqdIma8Ocx9nzpGygyhRENO+FuaJRUjTbMKF28HJikk+
jjVK0BO4YdVb3LfJQ9afBxuK9uF6ksMWbKfVXUc18Iwk63Bfjl+syPrt8eSGc9lU
3+Z7ssiOCAiGH8AMG+NlCy+1wQbl5rrUwU2rM7OT6nhYthBrMW12nAX1GuSzRAHx
Uonde8X5ptLAt6KE5uhSsXBFVuz4XMmRfUzerTV0ny7TLIOEay01r8I7MhZz8vyQ
fvjeZVkXRkXtWKQ+mGCvuesnXDblxvg+SMXHlRRWIidXY9eyJbQVppcU3c5HQ4Ot
TcZYbsGDAkyZ21qvdJTnZR6vfjKh92cwC/u4PWgY1iuTjIwWKgE5vt+RATWu/tsX
vgBvst2YIKfJcxTQkBYOyy6tVD5jxMjVUCo/Rgrzz8nRRzDl19phZAApIVUpN2Gq
PhI2ym7xyWskO7y6PhFejFcQGoN59wym2dPsPHgG26iFUzNoXH3shw2GWsaDT3RV
5mirc8LybaLmkWgEfbImNbYmkNJsV1hoh80SRqTShy2AlmP87Pg5kiwTWFV2JxqI
PsFABHta8bcOnOxC9QF4wRBDPVoSDpfiM6eWZza/LgGI50uXi+6UyUNNYAbsCLHh
U8r92tsQTbBF7+scgR1QjeRlBScC/G2WqvtOk7CNaoWSrCNzZFEvV5KZS5TrkG6N
nrWKAvbm2OOpP8mRrzWg7mUsTJhjiyaKXw+woRWCWwbvu1ph+lUvYsTHqqnqATll
mkaOpEdZ5YNUbkOjianyCxGCtRA3mQC1HFn8eTfUHBga/4Gn3IoXiBF0d1iqHLVU
jlYw+JSNMut+w3yE84SXhb/k5LQrBSsVZwKEJlKrPo4QB78VpkP7cgqJiK6NZMsl
5/r/ZYaTX83g5KyxrjQKp4tcaxaWnQTDIkkzedk8QcptoLOl22zvSoxQZoduSd0U
B1MwA6ukdEsCEzc3laveDxB2iBprcJkrRIAOx5kI/wGhRKCCyj+qm9IbrWbqc+8W
tQ339XFmJKZpmCjEZ1O6Z6l9UQQOBPEj6SsoyyhZRgHoCkUBHGL2oTIsWdF01aN8
2nw+i1TaFhj9mNSW4gzPFpnk844aDH16nQOfrV+JusGhVEIH07nl6JhYn49KJhV4
jgcYJ/HagbbJR8+VJrt0MGT0HT9NQJRQ4YIYmZBWn3CgiiKKuAk5rJ4y38HqCzOg
guS9toQYFj3Hhiz0m8cHyZYHu9dm1IcUF8EoDoUTCjWx6QAWa9jDeB4nZUq5Pybr
xW9EzSY+WQ+TF26iEhkpjH4qF1dXG1LnaMcUKeZZZ6ZAJy8kNG54Ls2KH7gh9fbn
KejY0mj1EP/OgJKVw8XZ7c82iKVOFlKmt1kw5lwuPoIhIkZ8CjYpfN+4banq6/uo
BhaMy8dk4ogPNe5K8ezaQjC315UvD8uY56AxagCNH3mCqI6eTH/Zm6MH6QjIpUeL
o+81ywVAzQP5XomLzgfgiW46AwnvLiSKRMQkGG5G5KUKZ809mZQKd/d+TdCGik3o
676PpgmD+6xnHnAzKeYMKC2A11vEMBfXFuN2VKe8FwMxKidYo9oGDgsZMQRC0iJ0
iGuamS60e4/SxlGKfhRBi7/Nlel4db9rWm8rDw78iliL2OgdyDrKOIZI8gIAlV9/
k36xGxlj5g+S1mvBa4JGwhDiOJBxOhWO8+3YwP9MOs4tdhWpBApiVWIjX82HJ2oW
RQ0TU9E3uCIdqhophTpox9lTg2XstTiR/ipMKqqIv8TC76C1XccAgoZpZyWP3nni
wCFTjto3UssINre3jlfQj3S0xcbcuBYKUQaA7QjPpWCqDs7dlc/LROhphG8jzQc3
PGUt8dXaHF6x7zm9N2icZn+E/LexxfJcWX1J5Cj4lBUGXpcIyGq2O71SE3oLiktG
/aGPrdHrvoXchAv+lRhoQC2UmhaxihBOpv+V2+oC1nG2oKBE/iWt/j7522ItXSAv
LVutAD/QO02DUgui9T/uzZNb9BCX0XA9uVtjSk73wJyPn0FPe84PEWwRRXceMo2D
f40qVMaEpL+YMpCTsYrkLVOF/Lc+YnMymWkVHFESm6dNUcgYKUFwV7GuTUVk9qv8
r3uGpGX9jfWo8KXfMtKuZtwrYnE/oONe7nT5cV+hj8B9fl/XTeLwJ73WOJG4fGey
S7c4u/0f6dXZLKJkjP4AtVD5W7+Na+ixLg9Pg8VP1G2mOu/vH/m2eHJo22Cu0dSx
dbuMOHD4dwq7p/NuNkSkJ9A0qsUsssqIpxaxecUaO1bFzDjjcGMf1pvH0Up2RFfz
pAnXW/j6SHXIEQ2eKcSUnLUAbVM7PJvop63um4YD39gnGyamMu1DkSMh7rwW1fsb
g8ye+EOgdyPn4CZYONodAH3SpPCzI98HFLjuJ9cwrc/Dwou5ODkP2NZTVtP6AYwS
fWgv+0scTDHC3H/yFGaFnS6fT9EmhtTlfU25KtbO/EosAgn/H+2oNMRN7C9vYO6K
Iph/yhMT4zJ0oGbShAzlapteSLBpa4coZnjtcK9ayD5oJyRMv+7LzN2S1Lch09R1
Bg7Ag7K3hKXQdfK03Tgm8F6nEbXZs2sYT48lgLGec6i/BV1seR1IR/kRlbnR9dd0
2fSx4jzBzmyp3HM7RQpUiim8z2us/FnwcfRliOOP3Ir8dbwOYZtEBykZfmXVYdS6
+e+8t+EWhC1pFfuVhY0I+mvDSwhqdZSfi07XGvqIktZghnq4CZ8HMEwbUyTre0X6
wAcPmnCrYeUoFMfC2iFupZ6nJ3rjz66HIHmhlp34Tc+28Ctoc33lEVku5MWPnh5/
0SujoAA/EByU14Xs2REPwb8MRBNjj1hTp6JTw5UW3BB/9TDQSeHV2Zcg4ymegsOa
IHBY5fa5KPWbgQE+RGnbAZ4td3tq/dwFdEXHrWkgQ/YU+h4dyZEOpWwh9cREWUwI
3o8Sh4l/q5CL2PI7xX+liRLTfWtBGOFqaHjhRs8bBGfp6iSPBHfBQ0GHi05y3sK1
Bt+gwt58M+DWXRgz+ecj1G+xeGfQyJl9wc4iqe9REflcetyc/IKkLcjffrF04kRB
OhAAr4rZRhI0fSGPaagVC/xWIwzDTLDr1IhaK2jpaPF3CjEFKo3bTZS1fpKIL2sX
RR2uJ90K/OsuXenNbnW/qpMHDzvtt3GGImj87bP8BjDNX2m+nR6A/I96/0mYy7js
aLlun048HmbsfKIDHFrTCkXr55cMOnyQ8kzk2wV65tj4ZWPSmiKcllQj8A9/US3I
p7RmW5JgaYyTXq2yHoMyF6QlLdlsgj09TsdULu7wNUH8X9tKYZC+4gQNWjJlGxBq
26gZF+COzg8KsRSvo+4mL/qxiLNSHvy/2LJs32zE9r3Nv2PyM7kHhS3JfUgXTgSs
/o4SjiMmT+yewH7QD/2WCiRUIkjWMCRN1NuB5iY4eT0XqVrG6AF2eNU8xVFBl4mi
m1oEcHNBi1ohyxeLMRbghmwTSZlK/CkyIL6cYXYxF2yrzGF54WOaKICoBDP01TGi
MnWMzmV/4a5CVohqqCj2IOdkbIu+ZnTdBBnfwHKDFYLhuqWBstTJk5RVpQ4sWlXS
pAtiqVlYzmLprG80VkfpG/7h4xvCN9/qJVX+J4oJgOyyfTYiRrhHEOofneoxNRcA
3odRSTVmHNBOgBwoXPBV8+JkDYkPAo3nMcQHuficsNLXgTjAXLNOdqWMMvUHsLiX
QE7y064wWmVRkSAj0q1b7fKWl+34knBuR7DvjlfWY91UfBuPkuaJerIxtwFObm/S
A3uLFufhvN6VmcbYZjBx+Ev5+Y2ydepKOX0a7l+oLnrVd9P12jhDF/QDpStjCHNK
C62YNihNzHcVpnsO705BNdK7yWOvBFy/dJU6Fqe9LitdwamA1kFhbI3+mWAgLVc5
ESL6oHiHJeLcd01EaVFSbYVRpCddNTdSVVC2kDdVPd7BXAH3RlT9OZVxfgVbjzOV
CjJ+/KOrRvF5e4EgnLLo6U6kYs4gfHYRz5Z4lKQzHhWiSPCFIRRH2nxWcOd7YHpY
HGzWyo9GGn8K2OPYPiGU3jJYNA7gCZ8Zy07j2+1SKkLcLoffpTqgJxzNHq06lQ6l
Sa8f8r41lTrmpiXLggwtQJetiGdch9v4x6aezMThjd0U9i5khGQvEomnlAg66vaE
M26N0GOUOeuA1x1QfO0DnSFOi8h+F+V3shHt5jFGWDRI+Oam2XUmWsk2/w7kfHfi
UPlQgOYLySqEyd5BCk1OWiaNHccxkEORz+BGdiXlIuvk5EJf7wDXsLx4nNMdVtMP
Rnq0tHLotjt/Q3OjSGb62AdUyMsz6A1YqGbEbGWZaRnxInDZH5RULL7FUY76LjW8
Gsl7KC+nu5sMz1JTHIV2Xz9PeAzSKG7vU5pp4Q9EidplkyJ6vJZOP2vRA7kLgwww
ipBBhLnrkcg1KG9sdkJsC0eCEOYZqRRTiik7G/P6ApcUT++97SFGJiNNoCgj+3H6
/VPivPk3H0KdegFXHwSH+qKsHcNn+D8XBTBoZN6hnN2i3gJRHiPbGLfvjKG1ZkkA
EzbhHR0K57fpJIcrdpdxK5/v35MCJD/867ZoZAVlKgFl7HCz2dbtcZTqaFDVw/7+
9fnefC3reE6W1sVLggzkQpOYHJVOSipXIhWTyTH7ZnNTgunVWkYXt9dhfmagXsJ7
fF+XTKEs3OHp98lMhsiHzogMI62K+09zO4fvW1Hof0Vj88XCptpNXiL5/fav8HUL
V+xcGPx2a7QaIRlY5HMBtK8t+R+jOI1rlLoqDshrMAf+KwtUA/QB6xI+AzKvjQj4
CbQ1WDl41tqO/cf5kaCkqNn8q0VcGE52WGrTrpUYbSAQ/9TKcNOY/cOdtz7g6k0N
9+t95jqeChdWeYDCpj5yj1xApaLY542zYcDppy1pvkGVwQX3WL5oJLPCMEXs6Csu
Q6nyZYlXpzmCRI/6WWaZDtb0z29rqOU2WGyRvMmhPyqT22rGZAQe+DdJi9FxGjag
x0NDEIeUNp5u5OyLxA4nQfBZAvgnMRpktzV+joAwXB19HB4Rxa/hDPDH5eoGRaMu
+E9dgYlXG++9Q/7nSlzpgQiCXrmresrMo24ZMO9pBzD8K3SaORnMZ176u0nV8NSK
cXCVwf/VgAs0as8106iHTylfqkarFbgo+9oZDm6xUGVBX8L/181n/yA61avvDxsq
Nm4GmN8Lbw9D50rOlKxFHFunxMBKlp72K0mm5SIZT9SbgO5uVsFVtEcjevxuakzA
EX4O3dyymyO09RzlsbE+6tKltkSzSjpd7bZzizvEAQi5su/LzpObQLDcPqMKsz6/
1zFY2UWh9rhYtvOjo0jUSGfStCWtP9tk/wsbJAYYOnt1wjaNumH3UzDs7uAm+6bT
WCel//1gnE5kJr/PlUfiJbsNx/4AX7nvTNv64YW8aZKRYEH4XbutSxXwlV3vfMSz
+KfxKwELECLU3Bt7+iKq5ftTwJ0O1ctp6LcRuyCuf+IjXA+axISlUC5d3XZbOOAp
LGPRyi4r9SHEWmphuKMR0RBiIsdUoFKw1ZzL9nTHgPPI0HaT3tC5neJDPr276HRZ
CdhVFaJjGS+AshlbUBssGxo13FrS3vKgY3yMijxTIr4yn8+i3RoV1y+thwBfnYmg
QjM5sYmn+I+/K1Pzt1Wnyt7XYiJt/fNYy9UsQPKanngempnTmNxisJsx7TXA06Gd
KBSxfJV9n/G5DFgZ8T6sK/r7UuZk2xx625q+PufuKOLw8xwITTb4mZSjteuRd0mA
POUE9FeF/hAtcLZW6QW82ijxbps0iDwK+/g5DhqbpIyZFVQxOjpNmDBIMPcy4l8M
B9AWaM+Rntf9aKpurhXW8K/1koFR94JlM3MiIeGFkESd5qJgOELKNUjuCZypTJFK
baOmYR7clRE+NnO2WU/fllCPkaqltxjHZ2DXK3md/iZvXfwtfZF4N+AJDr7xaYKj
jr132MbSgsoGtQehYYe+K4VDoxfjnsw2+MVo7tIRYlH2zdS5Vm3iM0nGMy6PzoQj
KaUpi6yT9ZQvO+Wvm8ZGH/HYfwpRZSYRXjwdP2vwyZm/MA0tuauC7JwzzLvkhhKS
lgtF/j23+Gvj4THoGQx+CKKIi8GwK9KUrIM/Ltyw6Aq6s+egq/RMtD82MOjscDe+
`protect END_PROTECTED
