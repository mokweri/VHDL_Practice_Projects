`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bgA9AMLW9Kv5tWBpYo0aESQ3x+OEi7OJeqYQ4OtsmoGZJi060KOExU4IxfoDVk4
8lK7vQqEBCsuBvJ7vCr8FSn4dxm8FtW7E8QiugC5/eALQyp9PR725JRdHASVXQpi
CuhMFHnwNDTx+z0am1+khx9JVe3CSR6bbrEF2Pt/ysboCy+CdxsytF/ks0g+vD6L
rTv7Z5KgGAFltasLu8qhB8XB3dpvrDGX6ymC15x6g/RfPOEeTRtT6T8v8Yu9wWz0
xsaW8Fg3Y/K4JCTggRJDkh3iMSIm3jS/tf3UdZUJgj77mHAQ1XIrDC1neoef1vYp
5AkcA43Qnn0WyaMuavTSo1pNcAbaU2OForxoMHnj7iBnOTPz52xEfxBVtWp6BP6Q
KGAZqNia373dK6Cj+37xy7gap9oDxMiBbEGvgLJ8C0qM/mORKSEBpdZUnY5SvfFe
ycxp5OpybPUBFjgSQoMEzlwvxLRncOb2QUuZxK6KDpD/C3eEEFhgcCnAaKTH78fy
KePPdT1RuLRfqn966+kbUey1CtO72k60ivkk/IqPxd8=
`protect END_PROTECTED
