`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgPMenbKOKeCNOZmMwxtQEwtKjaNCRj9926KwZbyRBo2O5mkmZZ9QTc++nS4hzWF
OZ6ZqWZuFsNH86kCRIsikSeVuVBq3RFEBT5A3EN70Nj9F9g0TLMh9lZjx3g8OGKV
iK3loHH7RSNzAcjfIJ3UFvgr5+DIw2uauCEiWG9PhrBsVmHrX9s/GI9K3UUwdjOR
b47z6CSuK6K1r9C8P19b1KM2pv0Hdvcysc6Z9UgMUzM/gfHrldoooEIJX0yLhxfS
gOU4quxrdBC2+U2CZm6hamn7Z1YJkqWfSN7Azn4jQoILXirmWIsPOo8PWVSnzqXX
7FFBZZhK1xjtpPRZdHhr6JjPx6LoSF/IM/fQH+cB2rDaRJugHpq7i5kbnMFuoLO0
Hh8aSLwjICQdWxuOW5BQ9EVapFyN4HJNGrx3O7clmbNGNZQtZo6NZ0Sr0GEdLiYk
uIF/nGo/MHQflTVxCthCmYPaolB1s92+lZq1KdBmarbFXk758my11F9xqCbNwbJ0
8D0WzoeUUC1K9W/Mu5KSC5xuB8s5PLPJZJwVWJeuAxOlqvsmprTdL+CjEH9EklQy
71M8ffOfXDWzzRD4DsJ6mtKHgRfcbPF79lZCyhxf7ahMzztswEqTCdfIa4Efkan2
33fhCM9I1xUW0UknoHOG9ZyeFs9v/GRds3fNc3RWQo4llgtSr2rjQFm6WhsorrYK
W1GQuiVXU1JBllaILF7T3RjuX2TIKjmV1qyfkeqaVmId5TALlNa4t4shgxybXyKy
XneXZkTcfwnDRz1hjlwkr/UFOXl9IxRSaUAArsZtD6nT/SjYPT1RyVQgmtBCtBR2
Gp4z2tapZktWp7nliqh3L9W9DAt/CgIjYJrF8i5hX7xXyP/1W4W5NGD15OhipIMb
lB6dBwdg4ccC+IhbHA6lZWQgh0cw3ya/sqnt6U0NDYgJnZON5LfOzPDSVsMKh7Oi
4NYfnYIEUwHxtWpGLRVIjpZq/sPlQoGQcrM8BRro4vvCNGFlgyBy/m+9BBBkiAfV
DYyvrnO9qlm4jI1bt1pwgRR8QGJAP7jaS4G7xjVWivBAtjkkhHUa3BGf4puFI90I
bvEnUKcidFbh7TXzB584dNLlZWTmssseUpQLDG5Ulz1EkBxJtlBUH9p0g27h1/d8
dxKLJ8kInoN+lhlsmhogkjykn1nbOy0fD3fnjmnLmiyjcDVzYEtIf+G2dEr/dRoM
R3C6BVqpVGgjCxdizyRyBDf+Hbg8GFbbEbLskCZeB7vznmwplZVNohlRbSSXM7Uu
zSwOQG49YpU1EEpJmYbi3PaUnTfjJnZb7SXmwVXQfs/f+6+3xx7p+3Ksqyy5vkEi
x7wDpzx1z3x0d9A28RDzP4RzxGCKPSaOsKkGxFHMXQmrE8lA4h0+8+80+SX+xmpK
kO0z5dJL5KL2JkuZhIcETzlgn8hu5CfwROA0a+QKFiwV2n9wfZISnPKl4YQUewA8
s5WqS/XzMp0mFTjNb2VkP+w09Awco7VEcuzV+NM1tk2w7JTnNvgjBqnEF5xN3st4
H50QuFnaWmXfO8KxGKqvlliwdRAAxnzKP+8c6Rf6uIYlTLX6RwtrNRxY/0RRLRFl
RpbAHp+O45BNmYvS3tWmBR4nxUixSzbDUwhVI92XF3gX3CC01V9C82FWL1WObKTm
uMNp/0llzYxDExWqQt9lrrfzPpr5SVL2xd489+wTNFoTIQK9BsT5I5MJaiiVf3eI
08ezAq2J4HreFL0NncKm9T9XvXOv7jK8zd7kZEsQgl+b3/lEp9gQAxPHEdF5DFbz
kMmArQsnNCVEG30GujuvV6YlI2yiTX6SFIdDwo6wp5vFeZr4wgZI429CbdqnBzdy
Cr9ccBQtawas+NkS+43vDQ==
`protect END_PROTECTED
