`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KNNHxnFBCkvf/1oZVtKgPQYJx7936eI0SvkyyLbofoNAl4k4CR5tj8WqnFH2PR8Y
bB0ulaLC6n10qjBkNFymAMze2CfuwFFY3lHZjwpocRfzHkqxE6APWGHB85KAyIHu
QrF0P4qdbr7OunwuEgu0gf8NuyEkfius7URXB3IYqNk0Pu0Tu2/jOP5frmGwjJ+k
jCh7NRO/ZMbFfknh4skAs/w2PP6YmWqKKbSlw3mAdJ7+PxVZlztw6kUN3FyrMg0L
GPrCq1ISUHgiGDoE7r8EYB1vDgBVTCqKWedt9ZFesp8Imb0D2f42aYE1sf+dDtNc
0TXx5o4LPk8DACdHzXhurWDHPqb0Iigbn+hlnZrY2EDssSr8W2YIzyUB88FgY4AN
tpTWos2w3o7UiL7ZHsSS0363bq/xmQnT4HUWeg1QI/cNt0iGPzVn3gKllq8hRRKb
7AFci3QDYavD+DYj1RklBOWSY0qIpqt7JGPKTFfZkUDLcx5c7GXX6ldo5zaYO/Ox
vgCa3JGTvK5m+MVADUfukBRDKss2ePIUEY0RBs/yNq8ABRhC6CutlRKcFwHfrz8+
E7ott+WrjS1o8QldhGu8aAJWMFRDFaRgUpeDTDL8WewEyhHPImc17Jgyiw8eYsOg
jfidFYYByZXqH8zv+E75Xfy0Nn02wQjj9vM7Y/vcfDeeKlvgBJMBm38DqmYtlwzJ
fmLOeNEQ3e8yVBK5ZwJDb0U4x/c0Xi2WVSuymlguxed39PcS41WYfv4PhSzQ4mIP
VNAl+Mb2GScCRYk82H7qgazKWP5+PsLwvjfrkUO9sKgAmHCyhll9lGSJNELlzd6f
cY15f5BfQMOxcGBYWMVdPiJxyYLHfsi97Ohb3Hwhy3jIkrs3f8CpEahH/vYIRw3w
ABhEfEbFbYRgUBVcIq1+25Sr3sdjZwR29QJNx4OKuaipkKcevzoBs86DQQfjtL9T
QpHN3jX4Y1c86Q5dZ+LsBJdffqE+5t3BX5PKqt1+yFidODdaPZYGZ9PBTqTePEmA
KBhARHkpNe11Xgi11TGdLiK0wj0F15liPVrT4DTteoJ7buISfoN2YjQCCHB8JxMP
wqRgkFBX8ox9qY4rMuwuVCNvcCNPQ5PjYpmf6pAqYRsQbCpLm+9TSJjzuNT8pcsE
j4ky7HrVBYFbTmUTEmYhFLxhDKolWqQh4JNoC6CXtyBFckUMj0cokBCaUsB33crt
RsQeuRMTDluIG4SpOc5qDCPuT6gy8qeXVAdCUtOYUvbpgUlZ8KWmCcbHomu9FlqO
AcdzpO/NQRIroPkocJBsDSsKUmnQQlMRmIpFh1NP26xpkGI3frkq51Gf5ivkt/DD
dBk7cArEVd4AXnYDKLrXo3pyZO+8jJcrbTuW3yLcZ4205DPn7gVDwZTDdGI/2ndx
G/Qq6PVVUxzdaAROVFofHtJBfevy/a4/SEKekqyJ0YnF5Teo9ImF8Yp7lIEmUBX8
FAKlbE23f7eyJ/Cx0/0P35Fpo3w7oUlpPlQnWy0P/HTWLIKThdwAMYuzXjrKsRkx
NEw6xJJEoCWypGeLxc0UINQNq4W69Le+iwcVQDx7MKDje0mlULzScHR3t8FOi5j2
Mev/YVcypGEaAl+Hno6rm0el4rMGefrq6DQh0+YZjJpmQUGwBBhuUptb8X9R+2P+
avsht15UEBfqTaxzTpBg+uPZO+zc1QiPve/HhKcihQ9WPjESTp4CSqNYkk1q+K4H
ul36b3PcZG2HrxP9fxcy9aHWUaho4qtWoiYdf1SQoL5UVC1TBqbsqS9RbZcOTMwM
xsQCqkKjkDvbOvKfiEHQOg==
`protect END_PROTECTED
