`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ee37w6FJ0EbcCZyEnancugyA8KTyh4pfzikLUPv4cnHhVzucM/sGCtfhA+DEIhoV
S0VEziUml1p8H+ZX3/DhzhzHIncuW9LMlZ/LcL1HCYEFdirarHlK0rT7rHHvotyj
JzqYwdfzxOro1HKj5NJUHMyZLVC0YBv5LMKlIhB2LQpHBdzxjA+bIhWaFJEUC2Eq
eh67qhO2/mdE5lwmZojKHzUr0c9yt9yLTRlVCQwtWC81kaHDTNXt5if8RvaZ9Nfw
FNhzpCM38MLyWOjllHU9lvySQA/yV5G9bAIjD8mT4oIfB9ADkKpG+EN35f/eNZXL
m4UsNFLzPwUqqtOMxySCAaeg0rbJokTraTxNaYxoonYygfWMdLMFgJ4bzdl8oezu
n3naLKif7UenYUDmvvaZ93bfD4x/gsPQaL3h/vKgr9LXRFM+CfDe9Sc80EzczzVy
E/los4sF0hgu5KvTT+HfroFy6S7wOheRPdDq6k4UamZc2EWuhTZl3SOD2tupchos
gYgaGrBeDmWYWMKx9CG72L2mEDDz64ot8pJhO8LiP4Y88TDESQnR2wqVHnKzqpRy
5Qh/sLzeHprn6Mc7s/X25nWyWKLypSvCMoy9a3GUP0Ay3puwYPumDa6UeiTM2NyZ
VgJjhe4LINlOKsWN9uvFMp/S4H9+w1VJw7vQPev5PsBI/v+Y9gM1EE7+ko0hBIcI
19NT1tB9M3jv/RBQG2yq0XBEgR8mitE1A+dL34NCafncbXSTD9uXWBTygggRsn3L
s0q2GpeKvIfvB80B8s1kJjIh3Z5ctU5jU4iCo9CZmK2FyGv5/oTJy9v0I//SW6CN
p7wCPj+OOmOvrgbc4h1edQsVV8c76U5zDElgoctdoZwJBzQQW6P8NsU9JnqaglYN
BdN12+CyF999cL1RYLytPE/q/RQGxiPcuYkKAbYpLFlUyjvAxFh6i7K9YXnZtW4I
9zv+xFhnU+bltfZIUx1DWWNUQTqL1S+tgB3mDtNrkK0u0M66HJ1z3XEDHJW/lFgg
9D+nIVoFuXd7O9dsJ7VUXbXp4B7Nziog2ovWHXhdhTKkZPm/Irf4O7j6D5TmgZnG
QdevPJWykniSRuVkOl2k0Qj/i+AzUEP6xAP6UTBm9/A5OtdGN3vXQ4rXBaw3DSTf
jnDMZfAUWwOfBedeStgwgHLUEyJQ+HhwssAeYqtx6aM+dG1S5j4gFVTnE6IRgqtA
yMaulv+9W0eKQNOV3ijbn2fyVDtNY2ooBoGoAp98lWQCsEO3y89/b5IfPuUMOjtj
szhraVWyT0mD5pr2nrlrVNyXWCgphWlS6kcqWIlwp9Tp8iTRKCUTVcDFB/WH4KQ1
8taoCI8Gq2Le4AOSW6BxYBaMqaIuIOS61MZqKyU8ZPNC8gI2B+sNjbAmtSnIMRIN
3tvg1DGe00HZ+i1famKQUSC18fdnqUmOZcZoRstUkZcqiqlRCfb6+k1ndXH9I8Yk
sPfS+IxzBMQmXwCPmPYyhmfPxoRNAjXZr5i5LvnWsidYrHTym648oUT/lXGeFf9r
8Uv6td7vZfxffP3SUuxaVthNNcgNVA1Hn3IWrhUv9xlBjHCdpIlNgMZMx0EKky25
N7PGP5SYJgq055utpxuKU7ELiV89HAEPnw8OWZk3Q7/maKmlA2q1kIFkFGGDFRvd
melhRkmL/nJgpb5UF0UTPnrqnyh46WKBRjkPsJGZB6CnAb9JRbWopg9L5ATxbQ57
Igdj8RHOmWeZczAJ0o7TXk1pvauf8tdD5mEnf+5NHrJHa2/t7w5z+wf7gCyHuzVe
rKNR3OEWdBWA4/IDEfOzHAL9pPn5XYZBD8tcjM3xaOMo0m7qw+P5b8ylwwgIbBzH
LbUX1uTPn72dLRUrXErddwlR/SNRTNxhZRlCFG3WIY3pDjRrkS+j8h0sdiQfHn46
T5QUncxzKnc1Ms+0T8xNc6+okBAtRe/qCOLL8I5MI1I+mzLRywyRc5PNgJKwXuXR
jvGgtkZWG/SzQjPbMpjKelohw5oozz6Ci2bKm6SNfaZh0zFSuT2WyoVg9CPIndnD
ODU6BCCMOBRJWZnoqeXMytMs/v4uMBn2tObVcOA1zTVbGwb56qlQI5bzUYlSf/i8
UyVj2tJ0TARprE5+RgIloFZu/0EFdJPv4B7BbPVL7P2SEt0MqlVmWPSZkVIRe2uX
5iCn5nRTJIEhax5zVCMeqsR6jD33sWA5UQwrhudKY7MUG2uJcs011biAotFxsWYY
lhzzOyhTrf53QpAWsmub0MMQSODN6yxM5QksjdTNjfQwr63SuZ2i7mEfg7OShY6Q
qg9+OXg3moydxm7556WQO2yw7xYR6dMC7c2SbGIPUnoxlUldma9CAO64erGa6jgh
iI3JyiWTCfV2uNjEILVy1qxBWOfdKLDyRNn9NdgTG7/CQT8/fS8CdcsJpJt5TiY1
mzPk2SorDIKuPUA1UY+cXuUu7bVlMKfEU9OnVS0CU9VJNvZaFYz/AaA5wfAGrcW/
0m4ubRxcrnBKHw/PUQBn/aeF9UHkpvJT11Yd4Vf3NHRn8hnqAPqcnQdqUWqOmKeW
9lsvdvTXvpXocvnubYpmUamxWtoe5hVKhQ6GI0PCeGC0xjtg4K7K2f2TE3HT+KfT
EUksUEAOPc4TglPjHUetfBaJm4xQ78QknnuMhxn/Lj8ew9o4wFLvrTX8Zrfe0ZBT
QRDjU/IKLIYdYgV/WPiv6jw/NYLjRAr0AeKR7pyWIP2j8EPfkWiBSSN9x3IhrXNf
fkcIVy7nMrdi98aHOq4NNmmZJi+XMYIG1u/+/zeWvzpYsNwRmBAUa75plvYNKp7J
AT/+mzRBZ/iGDv/o+kz+GcAa1swnCQ37JT7PsnhYvv+xX3cyVO3xkASzOLWuoczp
JSGF3fu3ACAGJOP/GdFvp/9LqhAqPH9oaoJUnrHCwVt/lNkzJ4b/3KeFC77F9BRR
io80NPC6XPKde4ObiztpiYclmU4oEcPsGG4V78gGF+yov2STfZh7m5ZsK/BqKKBq
tdMlvpcqGdmUDpEnuZ19qtwOZ9G+WPG16zJUb9gZOJ//oUTCPnyBD/pw0Fqzcr1H
/IL6lmr0jAxPP9xISnJZoOrvkcCb8lyH6CKXIaWS1iJ+NbJLbu4SP/EuqkdnzVva
bGvIw2mk84hK1d3Up/uRhblLju+bVQwMgWaRSLMijVoNFb2Td0RKf72CX1F8SG+7
2tpAfQjJjbZis0xjVLDPWb3Rc2CyMepUgglRYUVC/YEVqAljg1R9YkmH4PU4Ye7I
yY2MHdsHAUCx4cg2N40KxrBhjO7KTIhvzB50j86XgFSGBEI02anciexFZGlRMqHq
5teWDppoUK7kljmrXX720fI1SqxrYa8m1g5t9WsScGS9xUzpVI/Mqe/Pq696rnrW
U+EdzBxADBHAfZsSZf+GBns1ExsBpdmV5+z3vqGKmZ0WRPgeB/gHRRKhjzR9pViX
c6Hg0UwSPxwLAhkxvE1QvLLMovd0rEtlpxXYJ9Nek8X5G0/y2H5MtARZCgjOgVDl
xOGg8cXV6xzKOpYtWIt4iMA995iLkMHWPNZlQzphb+35PFY1NR+kloo8k24lXeXm
U8KDgTn4DDrLSFmssmNvuGNYv65V6RJCULZRfOwdrC3+ZFMSYGoJXsPk0HwZezLE
qco3x9b77v345Rcpi7pq4yZkdH7Yuvv3n96FyqBor8Ir9+uC/y26Q2N//CS8dZlT
iSZgGTr45hLepIXpRrTuBaeSlsVLAayvUKChhlpn4qZDqy0lMs/eYjYq3KWknj96
goeMqsET9muaIWISjSqmPi6w5r87Pb0IAGY63/c87AhQmzgi7S1ScwHkkju0Zplh
GFEVl04aQNPhpGhLtKZza3ePzhTfgNiAbuhreN5UYLdaWTrvUJKjRpGugVosSE9i
GKzUuIq9f/FEbEoUftsRoarVNLcPg3aC9By8n1RpMGmBhCTmJc0rxpuxkyjTsFqx
FKNopJmvrM3hAfFBYUW6rUe9xOnzOZsN6hOSF5S2QS3oGBPiR4s3x0rawd3UisEb
bNjgfJIsi7tsVdcP7vf4aOZHJvdMWu8kWS/WqiGflvu+tk3zuYQsTxU0s8vSYWQO
O9gO15g7IfDdUxrzSFenAniVn3dKTVcQkkVv6ZpmOlLl9STMnZo1ygCP2jzvc3fa
zXHGUX9mqhGsi20KvTZbhdOqjxqg5dUCY+YlnS0fjhAnk28hAi0UIHaZivG4HHVN
NDuVWkmHsaWCw3FoEhBtB2NCpAyvkwqyVI8V7WHQuPOmXD51BlSYrewy3sHuX7Oy
/x9egjQl1X0PQKVfgOrgbVlDwfxNmO4brVflwnFJha8HkwYV0c7GSOugHUTfqbWG
iYf2zhjC/ULxi3fqVmuUF3s+cL5XDYu9sN+9Hx9EkCy0ZzbJ8FJqXeQA0U+YXutW
oxEfutVBWi3Z0Gi6SACYU4C8ZpMBtkWwhG0oGOhHD40v+Brv0Hiac1NNkZcv9u2D
kkWLMeu1C7k2GJ/mFkHCPEs9/NZnQTElSJ6W8m/lOF90Vy/lcaQDmTioxk1asJvP
9fjzDRLoXPEfe6ybgfLB+Z+ajUFyWASIAOVALtzl2kE3cghBV0t3JhzYuOQaFF1C
TnIKyqQ02u5koMXXDi7AGZ5oZfYu9/TlYbMT5xTBjA5iZJboaDSUNBj8zbrB8iQC
VfK6waUNxW621WYFygb0xIwENTmHKieotIbQlqjX60U6PRdgeQbC1CgxHQpLEH+u
hdWmFGn/57zce0vSS943tzijOa79lfFniroaM7hDELcORBVG2TgD8X5ukZkMbwFl
86CZHYs6Dyxrw802f/0jdZeBwvEcqwIKiHxAIedf83bROyRSEZLs0SHIRrDJbQ0D
hk3q/Zg82nwNDvcxT1qBvs1RkVUbhPohyMwkQddr/J/+sdc/9pcuQNCAVLqPMXuU
8T/crpa6yOuxFz9YaT7FGFjA//ZqA4JKxu1+31hguLgdunzXDA+3CJ+bYMYd3Zi6
V8yPAXN56La8jd2j/zqeQoVwE3M6iCGUO2A+ke33DxFNXVMegK6g/G3MrF+6neQE
RYshYEIhVJivcsg6cYQYAmxtI3Hvb7/Ej2vZLzthjbUWbQ1U8YqNDQn3v9Jxaady
b9I6X6OEolRizFFWlxGXlJb9b88HmPBpX+OfPNrm5l2MOzBxBHA1VhLhYklGtFht
Ylg9ZrONiiVlc2HQ2aTDk1EuM6tENzqochssqNLvQ6DcIxrdABRkY3H+XCI7fM5E
+u3T3pDzmhldxHkICSYBWcBFc+1COxbz2aqnDrWh0lARGlBsJ3ROlQihiq4hUhD+
Hi8o8yUDq6JxwfegIjXEdFbejz6mVTXMAo17NByV7Yl2NBtus9JqD3OLHrKzFQaJ
BVUA/X0Uq8Rdh4Uy9y3MpOr61RiKwxEsNxxPRvO9WOWn50sTJ4NwFhGSiFDurjEW
MwuvWToe+V04sx3kkeC8r3+rEQYpM8PBFvemz2j/jOTulWRxh5C8oBood96YtIWO
BPIhHk/Q4+Rr19WFOm3p3FKRdnp4aXMgU0+Oy9YjE8nTr+6PY8I4qdWkmYk06You
40/qFySgwLMkbIU2NZOcdHXnWcQAdzIawH5VnaLq2mePnqleOUnNiSGENsr525Rs
5IGjVMye4RVi5+XK3Ug81dm+AvgzLTcl64Q+imaRCc3tSEfLLM2rlhtvdUZRBS77
2lmawo2RqWB1MGDp/C4A0L2fuy5nIWWHTUwuIqWls3zKVRWLuRXGR7WSV3YCPtP2
f0D3hPTIx8Qc787Xm82QhiB1XNBCh5uMumvHAqcqqWKCD9fsvcKoeVlhSzrDj8yw
SdpIgUCB3EzpheKoiFSurBc54/+upj3C13cA6QaM+0CSogsB/thxlNGwyXkhLykK
wHa+mOcnKdv2qzk+5IVQ3icUklLuDStOP06ECz9QxDHNDZgN5NuI6sbGnw7GSt0W
AFVRLpWOBgI91++VJ2H0mesJRMQk9xAHI+ywgKoj9zjG1zHCZZCJ/5wqTw42cquT
Gizcy6zT6LsdPmL2OBAF/sSLg7uhK/UIiNkgNoPM2QIsaJdhn8FhZf4Sv8t1wu7a
jwyBQeKu5nkUBeFMAKJakVJn7iSF2g/bGDjQk4e0NnMmiN1yEMKF0UuMr0DR8wBo
zKJ4nkLsfWSQ5ypWErkwMP6cJoh5IvDuAc/o8FwNIbyUJBYulmLZORqBDti2F+X1
JqNGeqSQUnEVmbe8biK93BL37qRPrKQOifdOcV5vV02yOdlT/L0swtJLvA0V0qDh
r2Ytf/+jJeFA2ID9Z4dgKPHjgXnWApDM8YBgvZ9PcJfayMvcsD35f7LpRrrF9iND
ihar1E8iMYw6scb7rLCvO3vLYxalGvsImaQSnZP1L9crUbS082lxM2T0ShfeAcYe
cmzhjhQUI1F0ZdkRpYqI90c1wI0gL5oHvDA+oWJNa5WG4Dz4lyZrlWrUY7L9I5Ua
axbsMdIjxjSoXGK+BK6U4kdLhbxU0qH5bX2oAzODmFhibdUZxici4v2IK3/pv/CW
YR6rk5j4dL6elNoW4YwnUym2E+i0GBzxhrj+vZO/Z+voPlFdKdn6R808mpkFCV5B
02OhbAcaYf94XTkzpfS/KfLRb7HP5NODd4IuOj2FX9BNuLqNYY4e2SYsEAgCdTS0
Lc0yPg0xgdyNb+v6EHXGTbsUzhf/ydhR5almbooJJk2/YvQ1ngXNhmDlgQM+GCCs
qN2N8G0C/oCtDfYIUq9Zxeju8oRliCz4ECrPg7KVTaGA3vpSPg1hi1kdH5F03iVU
ho6XOxaKJGvc1QtcseQ+ktF1P5Ewnh0nZqF1mHoGrq50tlg7Foe828QlPV+cWfj2
LmVYFOwBKGfOGBsZ9+9V7I+VM4MvGJMk7+9yXC6Dv6f1+/EvfVOqqssvdPqeMAtv
6Mg43xHjR1zGGTwW7dkIpnEAaY5C2cwdkqKQ1Wyl/v1u9SNU8iQ8glPqqyAJ1vVZ
jz2wcvf6uOsCPaElsyGvs4pBEpYOMH+BY3TdwxGoxZtKMZdJjVvh5XYo96wA29VE
M5CId+HLaugz9YQRxr3bSO5FKzhTEZf4BpodqxMNpdciRjwMwXpaVexxyJCq32iz
AUfCdEK1bdX9YHoDh4P9MnAVBUgqfQws+/Yaj8CVPtBwbW9DsI88z1yrsB4gK3MH
loyGHeel/0RWBJOs/jQx+RssJZkyKJGbH21H8yMlViNw/NLkRpi+UMyIF/P2B2j1
hfQA8+44Fkpb0S3jm49Rjw/SWkd5i9S2wgMiIm4fYK0xhl8X17oT69Y16XD2mjZn
f9/cKpZrUG2CujiUMVLfsUtIvnRfvZXoTQMST1Ni3RommA8aK3d2oQY3AICoLnBh
qn87lXmcUgL8zN+o/LO8TFRtHOVqVirxObtU0xsEBIiRHG+L5bBwcTj9IvbeZvU6
zs9hH/uQ5Vn6DlEcsCKN2rDHmXfupfIvk/JHkICTkpyJ3+Sgv7iZwkw4/L3ZvCTq
B6f253qNZBVPhjy5o0fC/OKNFsAtMalKt2/hnv6+oWxZz0Zo2P8OLRGbnIkqtB/q
1V8Tt1ZFopB0grFhaXctX2gT2Oin5eGlxGwO2Gtil4+x+cKJFpvMhBzEOiPc3UdI
ozv8os7w26QSiiuhqrgbMP8lTV8XQXS8VusteG/8ghzJriWhDlR2v7lHoKpqdNZ+
VaLowRbX8oMa7/zloKZKEr4uYFMZdsxC/bgPunfOxo9W1ByU+9ijf1TH+9cNdQtP
tW6YRtilCtu+zTfBOlhrhR83RJbYYYM+uLegvNzBWYGCkotoG8tqiqV5Ql5+L+m0
4hgNwPzderIOHu0s919QemoOtiya628gh82X0dtv4969W6chUT0fDPfP0tjBkk9x
kWQO8/AEJQJ/uI8GWwYNDA6WXXBk03JJTR3uQprmNGR2XlANLW2GNc6yd+QwVQep
ie540l6b4QGGwTNvGIN8HBEAIW0xJ1aggNVbiiVefODKZjU74jjSGktYlio9Fssm
NrLKj+lvqJl5wgxybGLziE0BUCOe08KgNtQtu40BXU2rWzRN8IVOololeNdS6Jni
+tpWUIYU60SJU0IMBI8VnGQjwY8qkyVAKIuUzMqLM2dY+/nQg+avn0CbeeUNZI8S
BCY+dni8AZ5mBOu21SY5utFEEEPbVneMEuaFviMx/oVmJ9QdyCkYVpBQK9L/WJAO
cEoR8mMovhBgK14cJTid5uVLC9MQ5yh/8mndRDjtSIdgZ4P7hghOG90MFnpR6TFx
dBfIvTLFPwyi4qcBAOc3BV4jFEF8M1VePW9P24JzjRONRRdpXhIZNmM9iqF6LeF/
QFz8j88nQhq8TbeLGxxTuxSnZdn2buCiaE51DGyqkVEXCmV+web2BPq9n9KDEczM
9UrxZyhq2VYI4J30DPWWrQ+nPLlkDXKHgymtjnRnS6TsmSxJXjw3GlPCs+NIhWDH
F7/flUqAjqVcnzdYwNFCXrld9KxSwdSBD0QFr46Gnu6FDlCcYdYdyfP/7zJJi1d3
8xSmolJQzmIpRLxe68/HMi2iIFZhXOkqeVVIUxYbV7Q7EPFb/hQCsVv9GfnySDU+
FLsydLeGJv/FYlxc1llRnWzAkw1dZsmGvOpxm0ICeB3Rwh2YK+euM9pXWyM7+N6n
/s4T0PvPu67vuofH46jpn/P/9rEHI/HeJbcjLoyBCFujK0X7NCnS6adf65aVSSNd
9h+xxXlnCx5+blJq6kW0OFFfwJHDbJIz1kAMGarime7i5IhLFoOImcPeFcsLosPa
MmXgj/6al1Ug8njKnVCp6RSksOGgxTj8RkJDneUMHgCAUKrJTAYANObkvgUrDaqU
RLidmuoJ213Sv7aqxOy3irtDw5hfX9s16QGY01JW0FrBpA14XArSp732d8IMBjwG
y5tELhCEcDfXfil+8MwXRN6rb18A4GYU8Uv6kkuBT9oMIFWQiH8yWRNa3NawK202
pN5+1QpvRKuQEyPnQmHc2bqKhu6snrvWhrVafPVMB52/wgGyxWRJrst79WnoLEMA
tIR/0C24e7oQQvt8eKzcWvYpvtUjAazi+gxSxPsA9nxQM2bgTgMINGKv/vXxRWIF
W3S4lNFhv5f1PWI7WIBAPmO6wV2E8IzbtgZ30FY8eKskV/DjmUrFTh56MQUrEq/J
HzSjAa1Z1RprX7Dc4bfTu7QAL5ZKoLX3cMv/NpyAJii7YWNMLNJNGv/Rt3JKEoHy
IFLXRBSAX+wdw03kerHhcOHobMMtblk7MBqD1EZLJL0zV8/xNKwI8Q93FmFy97lW
bYm7sEU38vN4JhqNDhWRGdhSLygo9X6LtTeOCRYxRTDRGwR5G6/NRjWgeXH8RHGI
0/sMcmx3YOtBjVoITe603/7wdJ3jmnOGfGyM71i5IodatjqBz+UGoPKqXwCIL7NZ
d1Cu1CvamEZj5uMVaG9dG/T8LeuNzxZFtPp+vqn2XVaElTCiQKt0AHZBIS21s4MU
gubf3bjddjve2sMJ38vJetSFaKDcr5tUAf1gCgrAfoAj1Hvn845964FRIOclkJ4p
hLFkczL4VD+R1XYJWE5lKocLrCyfbNGi7IOdrWfiXgrf1OmPZQ9jMSvR8KXQuxRf
A9qPZ3Rb6TQnhc9TVAQotSb4gxCAiYv8+r9xFMVgzwN8Oib9Gtze8CmD0zlnVP25
UqevsbxmDVmZoznVEHpWnf/t/oagIHA07OFlhEIOF8qrTb8CE8onldJNAv1skwsO
kqVlZ320XZ+Gf5gr+FiDtzt/5XXvSPLB2VE2CmaKUCJTFBsfO5d+KLEnDoQaaGoA
er+v9CQG89xxhJ7n3WKIVNLbTmVyZspNMhjUFu8rljrtrHWXKkAbrzluG8Mfhukn
p87cmcsNjtvVpEiGPaW5WfdiMoOUTjhylP0bc0Sh0uG2KdMKa2DsQgNx0iaGKSmv
sD+AdKOrrmfb4CEAnMVLIP6iAF2EeBw2zqUdpeD7jsTnuIBlXfGtUfpFUv+33Fng
wylxpIwZ6UZD9W6WitMbh7nvj6ftsQPJL5br19Hz2wHKJA/YvGnhbHEQJARjspaZ
zRnKK+pRQVXHj8YFgt9XIZ4VciuUd1GjQQthNRik3NPZyKAHWzNhGpe5SSP5E2yb
/SKURQtr7al7G37AYZs3FS+pjVIp3wM5E1pUIJiCMP4/hiNEqMa6ZkUIU1AVwQM8
yxAGL+ritkQ7/TlK1rY6z7DnOjuZnPxbQJZZK9tmF7jAnNAW3c+2j0A8qKmkxMk2
2PbX+HmEoMZBPPar84PS4q3Rzz1qarPs2ws/Av2OPp2XaE6+hOnUpc2LZAqk5y8t
AYcy4RQ+LqSNrC0kdWo1lnoQ2dyheRjjfJdjNzlPtH8fYkZ3ulBo3WDahlQol8W6
DD8SOSxGjC7kkib0+GmU69wCzHKgLjtMzrpuih7pvEw31w7oJNmyYP8p8rYPXdkD
CGGsvLafPBXiZbsn+G6GTwCRAeSLnjfkO/1l37hs82SPLzI1Lwu4lEVHWTGvy+Q8
5pRk7AqvFJpRR8zKg3KEmuM1kDEBFEb95wNgV+qRoJ8P+SzFFYh559Vrb4K4HkDN
RAUA4GfH+Ob2LnUh7J/m5HNuL1IqZI5XsQP0LFLeCSAhjpxY8bop3+tS+G1/w08O
zZyqM9LZbFAfDvE++Ob8Bc/01x6NZyG2Q4wRWQ8AbrpP0lS/+f6C0G5xr2vGZ32q
aRDpa/6Br2+bWw2lVbUxoaWWWCSbhuqTS//vP5m15adpwj8RNS0hhKhQ6sV1xUB9
kA0xOu1g8BmkW2WC3kIdJP03WLmXmHHbrB0YASQRATcTFx6s5nDIvEY/4wMarVKx
8zEoBgEjigGwM8ilRdyQpkill8KEn7w8x1E38f+Y8ngm0XCoXp9xV/jKJuhgMYT9
Sd4bsmL4NTZY521PGhSkbQWtks1SOk14skl6gCvS8wkU/XtEk/FS3Oi8n/VKlg2e
ykvJNVjK9Em9HBkknvfESwujL+lOD33Xg0QENpdQYi070mkomfI1qHxKtw5wJSx/
FRMEmPMTRJoEPW7iaiwib7ROQByNyOkxUFiyrnzV85crnTcd5EkuR/NR7OqT7T3V
1pz6IsvE/TdCp8DkHualugCnYVq4RyFar9TQRfGYsHaH1SDqOHJEe+4IZSVtsHav
g2UH8G+aPiOwVlGhKSRh+k8/tgZpGJfR+cGSOvpOBSb9oo2/p68gxGapngEVmzgS
2Fjoe/mxpGJLW6Wn5qeoi+Fc6z6znqax7KogYYCA56Hl0s6bVO3GDcW8x44xMp2k
y+TakMeyNTgaeo2t9/BDQplLt6vPgzTyOYX2J9BTc2fIOkoU0jBp5ssNgvx/qcu0
yEj9Wenzor4UoNZQjkUKE5FMmLvVplLVyXFAtbD0r+i7ixwQGFiSwCIfSMKHSQgE
/DQq4fxjQLCx1yLDZmaQTS6UwiiilnanM45rA0ImISCU43Hs6UZNEEpL5gedA29a
YzGc6Q6R/kIBkbtfsPZRCFCkkTg6Mk3p0YVizmn6UiDp5RJeCdb3HR8g7uqeFwOC
rMriOH2qvp+laQdjRnyte91UTSuzljaWgf5rir5ysHweLD9RVXZvvjqtjWb8Iz9Y
LAiz5PrY+LWd9sdlF0n7WZCoP5Pc+gCTWTvn3BiI/s5UwT4qc+4oUJrsMN5N7em+
F3Pv3EvL3xtvZ1JrjH8VtDcDr8WWa5dWnykdCwz38qMVChrDbLEaRCWwveBTSf+j
g/fRWyDIbdmMRwLJ0fGEwtijKlp6sp+Zd62/uynwgK2dWgjPCPXwBl9e6YfCIa0L
Vns8qNoJlbhypM6XgSk4OzBe5glZjPS9A0DmXcwl8x2HYN1bcHiZWxDJ6cI0ailD
Bjn/evyuN4BUoHgEMKn5InrsZTUbS9h4DqWxFutGxf92sTI/p2lsu36ofOfmJdSS
RckDunUHrEI+rbeujzBXr8gxGA9bV39NQLtbjgtgsS/IsZr6QyNaDi6IF2DLLX/1
kFWcA2oIMTl/LG5HHb/qlCgnX5QDZklLwE16dMr6e5w6sadJ3rXe7Z6DVKrxtJzQ
rXBTWWjlilfiKG0d1e2PjwjVfTvlb5QjR3U+KTzTu4liQaPhPCbqWrpeEH+E8tKJ
WEqBBprPbeslyqOR8pnSrOEGKNmzyiIkpRr8N3lEPop0bpwtopiJKl+lcdU5/MWI
i/FlT7OndPLWFtfo4LEC2stY5E4fRhFu2Kxt2ZKJw6zKCgAKqKn3B61ihvhuZ3fa
a26HD7p2G5qGUTzkQoDy3wTAGV+nfIz/3hbH84Yr4Ek3WtXuHX5XjF/1nsdiZN7A
JNEQ1Gg1GMtCSFArUT5/V6vcSI7LXTO8NHyzttv7dplF7lqGG67ViI3704+WtODa
vgCRodnRyitCQrs4BfUg8U9+TusdiqGLF1ZwoljS3Lz64eRk8My29epeTLZ/Hl3l
QGVWsHKPq3IdaLERH/VsU3/AK7TGFku8xcAWKt0NFj3DRcFCoaMtc/XhyEbTbStq
He4kj5tc4kOl7E0JQsvAbrboXGpxREmKQRVSPElqOpSWwtBcsTpxOY0bYMBJ9Fhg
O+a4hPCryLi1yDGCwUCbjagJHZG9kABqDQtgS1FcVVmv4lIQeb3ESjkMuv3jG/0Z
wI9t8SkUIGciq5FUWxuRTv85zFfuSbylpsfFOte3GUpb4toPP46OBW+wGWVMlqcI
lK8fBfdL8fB703AqpUQU0w==
`protect END_PROTECTED
