`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+jDU0k/9ETaHBCiRyIe5Ktp9rvB/UWdyBUU5APzr7b/O56V9MDRkYJ1CA3CUOs1
xmbbJ9qcT+ZOgpkP5l063PSrQiPJGJiBeF+3H45vFxUxbXShN+D5emz9h9k8/jy8
tMnnHKGECFA9DALags2KcmZwVVGirmb4AIsK8tr/Y5kYzdPltjqRHlD7kaWcMAG0
8aU0wRdd3P5y4axHq9/I4TltLwLQXfuau+2T9LPuyHn0oifezYcHw8aSGpyvgbQx
RjfW0dXBOyenGJylrueu6cOCBpNlj56MexLzYy5B3rZIxoMlkPmxSuc0YS/WYghY
foLIr6XptQYsfcjooLsHuFkW2SGYfDZVWnCp39PMhp5LJk6anHoaacTrBS0bXsvl
rHNx/Z69GoFWRID64lDscMcLrguWVhi6EUT57DLa8Xof5dMqiN/i6zgqBvYyrJHX
pFmQ6GnAUnA94OdfVs2D/NfLWnTowrDi8lJlkawnJ/GHZ77r+/i96eYy++5/JZWf
0yhqzrU01F8XmOmxPLndw/7qqdZUnRzSoK28ll3SwLDqmmKWvmCQRY/apjAyxr67
sgLSx8wiB4GzN71y82pMDxh8lnoX6gvexaCS6FB74MzwqJkG6rgAsXAv202VEHn/
2BDq/tPiCfY4tGy8Uvuf4U9isC5KDZ6afUJOhl71fvQPwIQOU9BrCOyMx2hyfKV9
Z3gAIb1HUSyvALbwdb1+MKB1XWmOq9lVHJsQ+1MMHXulsPnv3FpxnaoI9pCx/HZK
iWUq+LmMT8FhuAXO4bvyaeP2IxZgqp1vL+Bw12otCcaNK6rc5QYD8zuGjgSPV3ta
+cv9hNE0EUHWnyWomwfkNlf/h4MgQ9QoYiVc1mILaGN7vb7Hk725WQzf2vOi5qGI
xGBHswDuTqemF4TWiHZF2ABEoVsV1cs4I7oIwODuK+yZQXCv0825XzaxRWpxxcPi
creErSTD/eq6j9enDz2pHnn40z1W7ecRFXwPNcR5Vb6PSUNEwG3A7S5w2oyI9W4j
BJNVFWjrdnSMx/+1QdmUWL++6ff+3qGmieIaAlBSLRDl9kOyxSCmknejBvBXQ6vV
GWToe2DfQIo6fgJd0qtZIUDs9ZxZflSEuv1swXuZMKwynbXsuKhJr1cqrUY7YKWB
tdgMcQhEt5L2lGPYsuI+aytEPGouQopXxUkcmzEt8Y9zzsG2mdIXBT0H1wsFFR7X
Mkt4LFwJ8IMk/7Fzun+VvT0b4gZWoamjiWGkJlb5teE0L0hqbox08b5uiU0cpCmt
7Is7gUsDgm7FKpzqwbTJN/x0dtnUo7VRTOgkI+01h5IyLK+JIYBasP/3xJpyUK7c
UqJHiaxBigHrXMe5J1wYUf5xxSKauafbl1gqOXicjRo=
`protect END_PROTECTED
