`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d5YNVr6kWXW7pv465B8idprmrB7Cs9LBoluRiPEJm0OdIj3haSh8zgwP2evpEaa2
ld15IkULSdLgBNeUiT1RUWnTgcdA4nucBKOqMtdaUuB8vsnSleQgq1adoqafypaa
nSPHzknSqJXldXXqXttvYuviWoPUU8Lmi0JbRdJOX23ecKXyXNi3aRplN2YFswPI
6YMNH6MIhBXgzlATAoxKUnkUV+zQ17jJHAF5vRRg8EAmm8js1yXG8rQE7QveDbrZ
A+kJIk8HgdJ3IkIfTlHyLu/edBUtCpOcGq7F/Rq5rJqVeSu/HvMqRjtzo+wk9sJB
lF7jMsUOsFHzNdwhDZBS+Lpx/A8h2YpnJXifzreXByfPKxLY1dx9q1GiZ1T88Yct
pAdAOCOsvTbGDEQDvgn1pEo+eznnymfZ23juLeqXl9huwcqohyBcPstwW0HYpu91
V7nKY2KAPJhPN4wjCFf/bW3oH5Eo4L9PsGJxxmsPhkRYsg5uR2eJoP8zAd2HXjTu
I9WX/1tCM8iCheYmJM+oH7EGgF1JHYJBSfL1Yxa+U3CzcsAbJgDF0WDrpkFovs0T
3KupJsUnNtDT9ASI6lf9vfCVeiRAlGZ6XybFl89ZerXPVx8kghEx/iKaF9x8sz3d
o/J+PR6c0oabGgBxhxEahnmd0vFA0x/DuceJeM5sLxDGM4mOpfUVDwD+Gr6CSbHI
Ct2lyK9EPAQaQ0ewgqOimPNsapg/1tdiZaAMeQbpIPE5jgfqLVnzTM5lGZHtJh1h
VCcaDZbCtvHR3+eoso4xwo7znoefoPdSA05Aj60RiX6lZw8esWXhBiG41QDlWjM6
WKC1F2vXEHAYRkv/yu7tBw5hQb7x/HUzmLlX7uK+pwVV0YIfZ2DLiLeA5EV3QIrJ
XqTapOIYkyDFL4ZEoUZxs3nHqQZkFqg93aP4y3qplRREWIRq9Fh4cTHgEa51+qjZ
EMeKJ3NQvhBGXva9ng/FjUihAbo5DoQ7QVzLHgu4+5uO+0p05IAhf0MluAcXDJk6
Ow5v4dEdaaEadMagDzZov0KdUKG098fLbdoKWnSIloVxT6Bq4CXp2KPCUDNxki5F
`protect END_PROTECTED
