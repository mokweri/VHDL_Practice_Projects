`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLjBCZ8vtjcVqwOEls82SPmFrrg9eU5nJRmVQM8ezPEzkYHAbbMfZFPaBxJ3T2Fh
hfy834fBE2+Hmr+avlVOkzVUrG9Af1SucLbAtxiDx0PQdtHKuW5oLY2+mL6iLBd9
7qYCIvQ7NJ12aviugwS45QjPai6hAkfQZmnvvx6lKA6npwukD3JV8xEH9SNyWrBT
W02uAPxBKDsmrhk5TQU7dnKRI4CWjlXojluxIVVjMrbw96W5OiCO7/uCBjhBUlnE
6bZf0KwTr5vjeSFhQJGdphlqRKBInlPy1MzpBaLF2jQE4ZHVCJ8gqilBBmipqp55
AJEfIdrwMhL6IzJxvvNHZRj/oGKg3ZoLeZktD1O3Xl2AgkvugLXCyY+kis8xHW9e
nxJMy0ph82JUl2kcDB+t48bSRRWgOgVrvDxwETQ+X4sOQqkxKllWYU1vJAvt2oEK
dcapHqluuoKOAdLv02j+KOTRbooM/guHXOXgkRXZ49UuAJ8hGa/N7QPTWJ4kJmKj
cpdfciy6kSgAAagtvWQ5xh23Pl4p4qpVN9lhUoU/Rw9nAb4TvjVJMHTdxh5mPv6w
UNWAShZLyYkEMZgpkKrc7RVSAd6gq0O0slG6ClmYAv/EB4yQS2Zw2mMAd4zhQ61g
Kq6RG6oe5cridOlaLpCu8BZuW+1GMMIe0sFaoLbzmTcJd0FZ7/9fQiz7DsJ/FP9Y
yaMbcXefKdnDn0zS1zrQkh2dRDftlIADc6K1548c+pgPJepjhETY+E1gKMDUrs/x
lfDwxQJihCD6uKP3RcwRFT+/rO9hiZ/xkbpNGyMdnxyFyKbl0wnh5+VMgWkOsTZY
m5My3BysT/ChhbExaEgz3CHdIj3DOivoPApNR5I5qenPi42rz06Ljd5OHEcFGKEZ
ylKSpulUriHnYNKYAjNhg9mNN2AKOHtNzlv0b3dWKLYry1ulFtMukV2AgGwSPnwj
TeqiH9bqyATTkgAX3zcibiaiFeJ6k0bX7oeoGqfw2krk7NV8fS+eKtqUjRZ568U8
R/T4N95tMxH8JDp6huy/QtYUg6Hx70fb1KG1wqn7EdBntc5OBujC+8szZyyirTfG
A3H1OM3/K3kWVGycZKufWekkiFBiuI1EU7XL56CIlIjncqfTkbwpTmZC/FgLrY3P
vehJQ6OWGbrAedT/i4p/zz2yGvHk55V35yxmWI6W33rXVy7PFcNYf/70f9ASn5y9
XnOnhYG9MfnKh3xDy+Ft6a43Qkz8Y7mi5qKIB530n0ecqXWfPi1ikIsXIYHBlONw
m7eZcDMSW2YaU2iItN/bWDiOBKypA5uysNtwW6glVpSAjx5S9LtpJ+Ayh/x7J0rS
+h+FfR1jLXS+pXTKz4FS/asnMOa1H2OBzScSJnmkq7ZHPuAOe7hWuS5l36d45W+r
JkOQdsBcsBKWeIQu36SzQVmMx7YpuQVkTdf/HBfvSvCvEM7sYYCeVmocMW1voysK
0ScUBPoINzrd8Esg8OcdjZ54ub8+gVHdMRmr3tgoWJUVmPiZWpoxmDbSiZ0plaKF
tHmeLma1w771aAKgsnCxp8pntjfmiQ+P90UF0lN3BbYmY0D4tAxN4/hCOLXT4Wj7
KCciq+GySLw88agjj7GfvXEJyzCQ74l7/3yvzrveqAnynyMKUWbu0vkW4wlwBGWw
MfaEwNwmFUFeM4WduXL7i49iDO1t625K5fHmKgF+Z0Gv8I9WHtTnxVvYbNjZmH/L
pu8sQjL6/CorsgZN4WLHV6oXYkoBXiT8V4ZbTw3uRqdCwrWypaGinM4X4mQqBeTJ
qaMkrDWRNS0gn0jjOCu6hA5Eh8AP8UciC1z8jeqjqLFl5LGNWK1cMheEScWcvVec
tHE4YeI7dR0x8p6uXZzbwDfzSgwMwADmsd4Fq4SHGV2sjeng6iMguiGr4Mfg+y49
6Yuc6ky5wNhqVi5d5WBMcHqK5U39i9P894j918z+VcFeGOVbVBPF6RhoPMSa4O/G
S3K1c2g/VX3BiRYzk93p7uB3TVSyRiZSy+UOIav8m3jtFVtQtKenQxd7eT31Yh6W
jftsdGDCUabr5KwAt6n5uOH1XLdRinICOvN4L5lK1Kep07IDtbDduqeuFlpFErfw
U6gOXKCHppZrv7IvN7/1cFq2lYw48okDwGE0WF7x3+BSzZV3hSCMvq/ruIfetYF+
Le6hIipfD9hpZY3lUTkXqHkJpqHYB1SIJR9ZmBG5JJETaBCudVrEIReYyjbCJKAd
pRirX6d2wwjc6Ls5TtdNQto0bcvTy3xB2aOgUeL2mOPk3zn+oopyUQM792muq9Lb
CYgmC2s+xec9604EOVoBF487IxwZZO7byuZecESPZWOfUfB6KB7m/bedj0h91kjg
wq69wPlw2avdnWHkboW0VDDPedcVcgpXa89UwtpgY0F9CZ3sKyK2GGUBEV9QFAX8
ThYq5OlX9yEx5dA4j6/e/iNr0GzWD/q9Ff3F5UmJsoBa56T0QMKISvTJ9UZiNInt
eCiX2gsxZj7M9dzkbFHccTRPfQiSVAsQ0fxJPem3uNm8bvGzCVZVVnkWHOkZth6A
EdkRxQL5zf7ZvCS/Q5Cv5GrmK/7fXnllSufGbVRN4gEUREu6WD0MfZL/ovYRLEx5
4YXpEiPZd3sKAcyubisrY6+zG7aLtJT40+OxJ3aXn+GQLgs4RD8ZWzOD4khoeubd
gL3zYx64bYUqr8g4WZN8CkQTmuQjTlWa/QL3Eja6yz8U81v2ioYmpIUQFiJ/bkh6
7DtczoN8Iknpwu1YKwPiO47gusr7Y+qL7mEITZ4Hr30gpH5wb1AoySWgN2cRUwSN
7LQKdYH45mHNAaCXvOkgAoLTQd/MoiQaWYwSUCE8d8sOl4EfiIAbw2wg6P427ybH
vuqKhXMSPTXppBCYkyW0FnSsVgnNIztl5umPAtRXhsXC6jQj6YbMsArevd5623YP
t4fJvi0YHlBn9JGVGZ0qfOJXA3ib1MAKz1kMVPtpHsXPQGrbJA+IRSUsWJkr/Yyr
dcMJ3w9iA1UaEAK6KVW84mP3Tx58AuDDs4wKqDCJJ/aCc7Zkh2WUWsDZl2iJBdfu
cPt4vODzfD1sPO6RNTs+i8stwoGmNcfUc1WCWp6KrAQQIpadr5SpfBwp6ZkDyhwX
1KIl1Kn9gPkWEo3m3q3xVRHbJ58hiAKRcXR2iyKMff4br33HPLcXSly0YByC2lGR
GgE5G1aKFwQWLpHtZgvvyYPkXM8PMIfuj40cIzyQlZRR0IR/pOZh2LHIfTMjKHpP
/rZzrjT4up7BBldVNaOz/oz2JWqhqd8mnrgvLSN+E9z75NB5vU1KsnzEdVC3PbJ+
RfkE97Q7RTN3pyWEuydnSROi8+kc3vZNfyuuYa+GTdjI5zGvTVUMnTAd6fTcmMD2
4x7a5Igew7ZbNn62JUh2JeZsxD1T4GGdOddiSjCg4Xd/aRpgVDwv6n0/9z9H4cQC
5LD86hBZXA/9MVjBooYhj/Gm5aI3amTgGNc4pgTxZosOuABrxaKjOnPUYyLYiZ2K
DMEADCUNMfEThrM1t/80gz55ySdCyULmxAyUaiNJXtmDlEEHy1Y5LkJqhY8uXMY7
nNtor4NeTQluqxEW1idOV17fvQk1bc1O4eNegBS1135ZtyvivSGYMCQa9bs4JhWo
M/h/teyi4DUv/3bhHf81uf9HxibjcCqU6GIg65BQMwU57ERwkCmAU17h/en1rsht
TBS1IMQ62hSLDDj02qSBJ68eaVRsyP2IOtLn5e2sv2cM6PmUaECfNED+jytYAVs/
PsBJVVZ5JNfsssPXdi5eAgEHKr0FYRlpIFDF9rI+pxwRlXoErT6FSYowEgLYLizj
+NUZgLjRoX2n6vZYyPV3RG7mc2uF077okKdOWfllrxNoMm5frmERT4LIIfaOCD8c
BmZCBayuCc2ACzdXG2F2pAcnFyHjgy8E/bL4EWUDkZYk0NzBeVNgjsB/RtiiFAlf
h5M2jKUiPuucL/e9eXg/s3IPAIIBHfOCMEy+llneOCp0hiIJ3e3bxVAe2g6Pmb2V
sgfuD9ZxJG+yqDHOMPxEzNQL2zTNmavD7NiS9UNZ4mcmtxieWz3tH+pWPjVmfdAU
WgqEqAaYIMHQouBrnGQ+B7VAESy2hIaYvmzeq5OYX/ez0dNojm/e/SttvEGz21SU
Kykert3M7ifdMbVJcZawQqEYAR2Xf3Hs0k6bgzkF/IO0nCEsilKlCFDvQogf5lBw
UrCqwVlbBjrAopV4+tjEe/NYndZlnvk9aV1ZHkcNxHQAFGJg0IEg4K2yLIYWZ8Do
gT+r3W0oUrAXefkhL70aQYQEmC8CVGkn5ZPRSDho8/og7Crz3+r6FAHk3Hm4qWwc
1BbrmcQJ4vogZzabrHM+AkkQR0Xo25nBdoBmjQZN8VOs3flqQejk4TpZfJECtlBi
yPnX/giHpAMjeOG4JZt64qhkIA+GLAtiPzENycDjMXHWXZYY6bknHRsENenFzmK8
ESv1F1DLgrGGWdxzjfyZBsEX/JPx2MIiK1IeRor8wx2MpsBmfo94sNhu1gKEhXO0
RMWeYr0GTirjfEgVcnFUXfmIy/Pmujf3MJ4+fSEARhWEXffAWrFbz3GAYh6yw/8e
FPXPBksJI/zRyM1QdJclQiCWPk4HEf7x+tJtRdUcbXAXluXEs3WluiKV2buimfIk
2VHiijGCP1mLlOlKcl9pUmer2MeWY2DhAENNe8IjJhs=
`protect END_PROTECTED
