`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sAGjVKN+8ysvjKMXPaQLW2zxbfSAw9Oz2gcL8aB8q/p2O17IKeRHtTTvpCfAQ801
3t71LbxYF8V9eM8ujoJVmsQU8cuNul5Z09Xg/QVKyuMCrMIxkPmoKW5rERAqK+8U
4jgUztPl2O3yBO4Fa8+lW9sYDrqdr1YIzcNVQMqG8mZIBWgkIUV4SIPXuu1nYTQi
1Uj3C4fA/ORhQIZKudFiQLnPMdW2jKlljQ6UnI0cZ5MnRbCdV8+tTWUWF/gritVN
sm5mNt9iZO1aE2cgS8mTNFlbWv+EMiAnEwaK/6SKRm3r6SrBubAQtslHyFzqozfv
bbf1fBew2r+c6aF99GNZAiKPUjgv0n2tg4v53BihS+E/OLDszJNYB1ZdLFaalgSN
KevL8wm77/PjPO18li+HkzNqD54yNxb/hcUdDy8y/kIs9u8q1UNOfc5xaofeRyQK
/wac0+Y12r3J9/T+yQI5KnN/dVlNtX9/3b08RqSAIHlDWQcbFWw8Rf/zMnVpiZ/W
O7MrZe4ff2pT5qRfOmpqW6s2Jij0OmBS/K8k/9HxXF8cn0zVVqG37DC4oMDOcVFC
TH0ayJU7RPr0HO3AQC+vWxJyd0zvAlC5cpx9BOHIYG5XfVNMjjZUasTqnLW0dQmU
ZPqfMAcj+sYzBjHh+URC3VmFambvfqwlob+cdVyJplRXnfaqepyCF1ADF3LMsBcJ
f1XxGI5dBcjccoOUUSNxurUOgNX34RvLSIIVLKCJsPaZTALIAjruyBewBoudkibs
8oAqOcml7nK5q8TKE6ehdajfhS9KQbEUZnBYmHRfdS6JKgfhGGuFBY4IZ6iGS6YV
R8KIMQLo7dQ5Z13Ka9oPaaUVfiYIOfYgOn+/rsyIt2pfC1UOecRBXq3kivBTsV3c
wzMkTkk6fZlbaS5ZWG1+tvlgDgtUgq7/vek7Wb8Wafmu1M0ZRb6xCx1NA/I1hpl6
YK+uWKHnnROokeK/7Uwiqcg2u0paRJTfAtYVBJ/Of0ML76FosM4JICE/ZQsO2zUa
RD9RETMpJO4zWsMOiUyMtRrx0zl32bNSQIeVjIHodsw=
`protect END_PROTECTED
