`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BmrOvaWKhIdbD4nESpLeFg+knhO+/e6wBV++V2cZJ8ZvtJWms5QZe6BsgUrHIZXf
6NBPCwCMD1GoawKBA3CwKFP5GTwvmIgc+xGWimy04iyl/abq1SToH0F8dPkrkGsl
42GZ0getQKz4mB2TETzG4X4DOLUvvK0pGwGVxFWrA338YEUMNsB1A2UNNocPoiym
bUWxaCpq/mxDyRFX50xVXsdtFZ48NXQ+K3ntwzxSojFYd4LX4AOOKo2oS46V2NNU
PxWRnxZSvPDUJFIeXJBmKqq/mB0FpAD+tWtzxjjYByvZG8+klmmx0nINH9T8zukv
fsb6yH197Fsk1gL584xvMK24/Y2ym88oD/vJCIGXZjcE+SvXMyVcXCwNpVo6nBHU
Qu0dGi7JWXCHZpcFg+0dadj1GJvg61Gio7YYVSv2EChU09mJuzLs40on1iyML1Ha
O7FGLoghCgsVRdj45mk6qkxHpm0lOntlty06b7KJsacLYDYf6J++KjYRjU2zcWeJ
w6AVsbH+uSoVzyZmiUm6Fx7a/entVgNesvW/WhWqPaqwsxzOQT0mGt8DpCQRPnIp
J41yPA5cFj9i2Dzk7V15sSkI71x4/PFtA0k0mdwaVb835x3IteIntV0s/PFUe7Lc
FLlKxDJ8x3R0hwfY0FltGb0OwFJwPtKiAd+3H9eZq849+lhigyh55TyhAFQGPQPt
hA3CUUD33rSDAtoVMKBWCxeVXFBjVe0XdyrRGFkYadPCU8V7AahsTO/IrnR3OXnX
VcKS/SPfFXMmRtyuMCeLuPRgAokqSELi9lBXACb2KJ9PANi8mllzXB9rZWIN3nv4
O1dwa3A5WxldA5SutHV6tYCPFyhsg1W6wcsda0Y/UZBmcivbljXXRev1VcnFadBm
Z9ybCQZfzxGGV9Lp8+iQTJgPKTYstZPv1vSPALlgW/kTc+XoCQD+nmEc6G1dgIM1
1uLpZhSPWQ6tW+Dc0vpBF26PyMPkEHei2yWcopAXy0Alf9LO92xg62kZ2nQriMgh
FAJM+u/tQQA1THhInU5tW6dtRNzRzNk34ro+BE3AIgrYbyPGCj/EtTYd6ew1fBdh
woqoGVLcZSshu6m/4JYNa8u7D/TzjNGxx7TdUpsospqscx7FDy5nsVygbxujMbJ3
nKBPrJJ5+0STQ7QCoKB0stKGh6m6/O5aKM27jrJi1ONbAGtFeYW7itcDYzAAeOzF
ShP38HG3vvcFqVbooCvHdT60i8hGONf9mMmOMegupFO6JvWpOg8FZ4C92p702wNA
8BoQy7hMNliUui6tscLxN7jz5+B1fEeu72WBTolvyr6Q22n3wAUAbpzuX7TjyCFB
eUzR6Uq+s4HtGI82Ld0HK8eunkQvY+luhUVJEcJo22io28MqciN7V4hzVTDQRRLR
KxdmqjPUfNHisLveef9hh3gv7Vwfyp0PwQhRQmjURMW3DaZUINCoYb7U8qUHvJs1
Hy2+vnEOHCr9shlrPaDPVVgiuJStN/LT9vS+qyuFDdmhw+dksnL/5QWUTsm8xhv9
8Ibi1rJd9UYuNZ+FfATdblwfakf5yZwFE8Z8fsVrlip5NL4iPESZCHBL/DYW1ANn
WyNnLc7PALM2YrRSYOf5dE4LhpXZ8tmZXuzmNBGWg1dQUsI669rJWvkKYT6l2DwJ
yS+GnBSTw2HtWz07NyoT6A==
`protect END_PROTECTED
