`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MSFvx6AuVF/jK9n1dkETY0I+t7OHAsTjIv+PsvAvR1/S2nJdjUw3v6/O5PxoUCKD
H2Y63zKYp6cRyPEzGmIhS01vAqjS5N/VC1CoS72HHPGPKMMr26ln7YE3Y2eeN4gx
/9bi7b4XhzOE86ziixLm7eVts4jBsfwfvhbnf226n7md779gveNwlEArYOaehCY/
6ZvOKySlsZ4e3i52rvDYre1VkeQ32dMgMrDfZnV1d5Kcu7KhwLvulm3n4JXmFWmg
nGi7Y04ys9/xYD3i+Zc47scUhzm2MNpQscyTKHwkdA5ySKeskyFFz3Zu5M9h8m0a
GjQQy3gjrg1MxgSrfzLyxR9/j5fPHa4JVi1JG49jGxg7Xwup8Ni1lGjtpS5Dsmx0
hpgrWcZpiaePLU04/BjI35WqZ4vYKhC4+9ogLBvX4k/eJNhq5OEBGiEOwRAemUtC
lsauM3evM02iBD7baQUhBvYN0/RsFddwlFc8HACJ3y9yiV/AnoWcX7EnAH7OTGyx
4e9iOt6jq5EMlo+BIaMIHcZ4p12TtVjtCTQ60TBcJ5D6Av68wDJFTh631aDx1q/d
HcCBi4ZK0tX4iVTlziry1w==
`protect END_PROTECTED
