`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Co+CjxKhyZ23hPuQ9gZa6kkM9G4WG9RqSwsfuUD45a/IMgIlgnKNsX//Qe61h/2h
BivcVzmSuyeJ5X7WEXfhIxL2mmFZYV2mFtay+DRiMNIjQAjMd4WCFE43cGXbVliR
udCjcXH4nhqYbX63vGyLCT/8ml53zcqukWZwv6Iei6CgXIzZv3u497+aWMxK32u7
NBYhpjlXyj61jF8YrFyzJOaym8NFkKT6rjpbir6odSZ2Pl0EyE+AqerVshqE24y3
uHXFjNk7cU5TTDYPCABuMpdErPRqxkFl2eWwVFHEG7pO0iurA8DSebEgRFDR5P2i
f1Fre8YJXk5tdB+PXoOz0nzmm62QVSXnDKtCOW7CzkSVvdqcKyAZUBIcmB0HSXiG
OvQIY9Trq5ikA4nxqMCuIDThyAXRmusD0s1qf4fyFUiRH8PREdLVud6oCl1q/2OV
9rGJaOuyLCFY8r+9er7bMRsIujDR1YPKFfyw15FMJBbpqnKUgNxuIodG8n0cAimU
4WXCWe0QRPniGyJd0OO0GjYpV0Ahn6Cgb9XDvE3lkP/DzU0GjEKnCcmzv7Ff+kc8
wPRiOkAyVFJbmJA5omuKtYBJ0SHZGLgcnjJ6ESRGKDHk4asEJcxnbHqgYT2D3l9v
rX1o+1WgOX6coAPxV+LdneP1lsOslylpL0vTZP3X99FOeYilf29t3Un+AGe7sgdr
WBv/uoAOw9sKUPfoSpkI2AzphCqeCEeUmok+76aMbYiyCwfzbZlB6v+esH+B+h82
Eavyk1VBkLix3+rofNA7C07j164BumI7yT6IxwQIV3esx/ut9L/cVDEFS0V+AH/h
DoqxLyfO/UBiCkVV2PuamfHluT1FKHc9vtPPGEqaSVPj14XOZHDRqqPQYEp6J7Rv
cxdqh2YV2qkji9kk66VQ3fRawKhA5m6rXVOq2BWQMOrHXle7LFpLR54h4ThL5Z6B
H6jHx2/myAphPHBeiBRbbqotTr/nBOVAE3ibOrgS2LkexaDfclTs0ujY+LrplnI9
A9uKwoAGOjywfGh74o9nV2N+JaC6ZgrJ5ncQYDAv1wLIEIjyEFz67ujUvtJoydeP
FYRC3C8bEszA1MRkqsH1mWx1Al+ln8pShbFGw6wAM5N4coHPgTTdZAARBReUb5mL
ExtJEwkaP8Amr/fBGCrwLbTiCHdBS2iht7iVVS5NlrI2/FevyhoLv1MWV5GbQAbr
8yoySdmQT4iWgzW/eSWcUO+/6beuarexaaSYCyG5oOmaHgCjAeTx7EwGw4InmP2M
JJJtjlzmwLBT/g10C0MhyGhf1PwyVcf4SQVwK3xH9qxhgFWcUzv3SodTyvp3flmT
HL1k06F2dY+afuSI9WU7iA==
`protect END_PROTECTED
