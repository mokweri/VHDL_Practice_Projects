`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9ZCteMo1Af56PM92ZPuDbu0PYNlkENcSkBy6nvQvGbmD+3P2ve3xNjxloKnUYQ/
W9sDJgyyAcyr5e6zutuve9Wf3eqaFoxiwS2BAJgWWjkGCNw7LkMk9dw28yy6Kcxg
hYJsxU9vYjedg+yNN9Ox+Q4YrsyXhiMg6noVI7T+KRkrvmsfU1aS7J1pqrQwdBCH
ny4mp81yucUFR/YwBRpo7Wc2yc0qDsdBlxB7Wp8KGJWBbuMpoBY+z9+fa2JdNoJI
BhBbrBxMXS9RVtKgDiaXqmw1CA+k/xo72dL6YIx1AJuWEwaoEKs8B8JTKtwtObPw
1mDLMZqJr71vC8t1U/vKKCZXMPS/IOXfpfHz90uayurrF4aDTy1AXrNaN1JOxa/D
dJfeY5mlNmf3Ls9Cld5BHMMBcyObMLLAMzjzC8I3BGCJcCUo7GCOsNA0kVkihL0X
wGbVWcZchZDI9t1qYpAkSSmmpqeXmbEeu+g68jXokoc6eflM+I5n2DrUxveJCiWS
nNELFcqnLbFYpIeqUusUgNNs+8DQnX2pj/nGUsi1DdT5xjJPekHvVE/XQaDn52+B
LsTiARHiqjsG0zdkmA/Cpq7kADZfKxtyhDF9RBeeZ3CCU5yfiHyvW+oak7A/y2Vj
`protect END_PROTECTED
