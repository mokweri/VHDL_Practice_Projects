`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hAazpB0HkO+x4BAkwRbCUYJpzYmOl8MMpFPphmlWBb6XDGCq2OO1Iol82dSntP8v
rTrC0cgl69tm/AsjGXXBOiK+BzJrRhb11zJWOOQZJWnRKsGUkzjykVPN3okXl+Eg
HhOhJGbI8hofhvuFvrElEGa2OTaJojes3GPgsfHIHC1LtfEjrCp17Nkyesy8W+PE
ga4BFjyFFLnufj4q1vstnzFXaAAElpcRmNN3+BhsXWw8Nj9B4ZnswRYDA0AMi7xP
diuzG4yNt6tlWE7cjs6jEEIudPkTcIeoCfK2kV5JjOU8Lw4TQIWSOBoiiuGc2VIK
cg3ChWFACg93WpfAHNVHhOM5s/voTDQF7W5uwfFO9KmO5ne32lkJik/qsrpO9LeH
+aZrEDj1WBMXsIKa3AmD3ThKtLTmIHNcfSUv+7w+jDHDMsQJFKqy9I19KaBy2SRz
J3411MBKENrw1XCHOEU5WZkJBIKmRIAfwjNrJ3DtWgW5lRtpHmWdOUiQBxGv9lhF
W5QDq3W03OwbU0Nd+OkRTdgOc3znRRWE3+rcEPygCTBUWUQC1KPV0q8M8U/Yddjc
8kbO4nWjopgoEXAfntROz+D+slGYfWrUkIIEPPY4wgGQXoRdpocsYnAToKBAkCcS
jp6L294u0nPzgiBpvZeniAkwx5Kigc3vb40te0k4FdRgIC2Fua6MLItJeY7CfX2c
vElIj/+fUjMbuWSIDahTwecPFGIe/uqAwUTMXgwxhv5yQyNEPQpmBfOxivsh6i9X
m14CQnoxgDWLPztrty2BeIMWYpVgaCEclgkSbRSxKYMKAsv/aK3L8wmkhwHo3IIc
LSlXkIp8SqOrNcTkHvdMdEEfnY5AIswHyTn/gEUSOjcmi1tNe6sl/wNxae+MC+JJ
tQEmez3njZvy56AsMlnQ3N2s5ubjCftevxqTzZ5OVF9bcWqq7ud745lu9NJ3C/vX
3UH3mJlMMmyctiRo9yI+gX0Kbxq13XZ6PvRq7sNdXN47XcwnZIsORshgG3jjaBrd
y75PAEXOxaZny56D7cKopaGTsk+hs9lOR9V4je7fC+SuTs1RzqVkDcgZ51RghL8G
ZwBB5XU59In7ofvYZBbvocJVKmJfzEzlcutIszhFG2gz4jbYhTSjxIPL1APVoy/5
xotZXWeFWOSWPxSahDMaIvDd8E7sj7PmOySFrZNLpw6EJrBNbuiVF6FZFV7f8bFF
iknA1x4uZ4QLaR/IStijWfRNkgSG1Y5759TBa42tIthalnoEbiP3EVZtxQIxMmRB
BcGCp+5nN1AuOyCh1yK0yCsJnSm4E3+MsI1CbWU8lw4+ffu8Z51p6eonIW2A3Vzl
A1V6Yqc9Jynbh820otliWX25NQ8BhKCeXK3cLmDE5FIfLqjo47hxPIiXKXPHol0H
3gOx+SA1BXbTpIpRMSBOmQDduF8XEHYRJkyEn++5BCeacK4hh4CCJeW5WPRSRrt6
yx5BOjCqOqLSl8DhBRHnmFXuVDc1HyhLDJF/4ERcZ6B37ILukKy/hTn7YBbiwy1X
PTVqBySwBB1Qcc3B59WyFUdVNYUyS21xFO90ujPuy3AXfBvwpK0Z8qPOHUQZ5JsF
LPlW7chHC6+7MyEStvU83LZJYdiycbGSBFd/NJSlWBIbKjXnDD0Ot9d9i9mQKx4w
XN3WBUNYHqaeqmg8SIEJsv1+wwhHggTXQr4oFrV3E0Zy9C1hf681x0E1UtsqKdC3
+bZeC/n/nvP0tNCSep6e7FbyBVXJEf6AOHpYc8giHGIeG/5SXJY2vpOEMJPUjFUy
ym4hixzUqbvahyoYV2gQKMOhQjgzQDOyIQUymiJCyO5Ih6tdB6HvWKB3yabiiLxs
9WcOgxA+xJNdzQdVTz2iB2CWsBI3voPpFebX9bFRf/sCPA0xGw2sVgykssu3/Ge7
8Av1obCT1dh7chermpFQJ1ONiXn9HJrx1UVYGZ53dBVGJRqcj3HyXiA0kUqfKvTO
auXI0YeEF8FSvjLw9apRurv81Pqf+ezUANK7eX4g++OWS9cO40atLtv+Cj5VFaqt
B5wFuh4tH7Rp3eQ2nDC3WXVOhanq5+3spWRegnDLR0yWvsL0J9YoPsQe1hE/9KVt
ssoemnQVYajkpgpoj4GRfaPqsta7pfk8bmuxIjPpWnu6d3/gjhDq4hJXqiV6P81H
2g3Y+RVprl+dv70jC3wpZHnccDx7Dq6Ls3URJZyzSAdisIJCkqnyFF1Qv/s+mkg6
ezyKhcia0ARu/eHsIPhPmdmqezQWU2isdJvb23FzZW29A2uJEFcn3ihhIjF2MOB/
CvFp5opOO2MYZ9wGgWZtG5do4Zu0KE12zar4fZ2SU4Ydcp35/eIpOjvoEV59Iiox
BhYzpNZ7IrAt3Rve5XRsNMi/8hkg6emV5f9pgV8Wn1/3vejp6e/T1Ie4K/PZnRRS
Y0MBt4UZyqwr+AxEoYOQ36UfPbY8xMlWB5QaqxMsux9LfCLvkakQ5seTEQNprDzE
rl/c6YM9NuA5gAGmGEA3Cc01hujobQyqN6wnjVRVT4rqDW1KmvErI+VeDrjp1uF2
wOhTwVMgVFuJ3rirujpaynVlgHgJryoQujBjymh18eFdQB8qrnkiww6iyPjB75HE
qQXocqy4AgeX7KJoB4/iGhnhvoJSUPNpom4keqBu1eydj3B9R0zy6/3RlBN0s8bY
Mjlv2xWo2hBwfHyw0FzoMveGC6Jl7nximYbTmON6x+IUBf+cT/ITDKlMCIqI3EOg
afjCnuay463wpBnFqB0+NWTMHz7cit7XURym2pFyED22s9fOgL6aUCs0xgjGBCe7
WVf3/VD10dON2HfAvrdZI1Tt5xKNGgdMgCq8qh0Jw6R72+IGsUsiEaftHhe/kTco
x2Yh4CiCUFvNJU7NleQ44B7WWec9ALfMadkh6/QgdwJjlpYA5q62kv3PdMSCDAkf
UaBO+jh5zjCtQYPqAKIli4LfvXKfI5w6Y5tUhLK9VLdeopexoKwuf8dA0ej4vvAb
R6bVLRuNqWj7WEhAzeJFF59GSv7ZwTxUL846gdPrMpDbkjTA2ZiVDcj3QJYjUPif
D+WPSvgOi2SGeShAQ6PuKl3p5JEYjAISYddUCd4TGFtkRdL0LNT1asUeJA2czd1Q
CqchoL0QTabpOgzdFEgDUXpAHIWbJqhH71OUF8KywaF5Afl8lzJ10NCahZG0Z6w+
et8+6NnrQ3Wzv5O46PoRgX6WeNQDYmTdwVdoIKpEdrFmm0gofiaffKbWoIw1yUW9
5T45q+YAbD4Ng4YzBNyR+n5/78mCO0FOW8vzZj+Cvq8PrI2SBHnyCJCIcxVG0gGJ
oD+CMIshPw4HWjyHGJUojejwG/xFds/CerGxnj+cZBMpVK8dYPRRF5AbKxZNzPxn
GIyBGJHm91J89GBMND8mRc9MDK2TkQeUdX/+vWJYP1Fi/w9EBbtwRELLAf0uJUy5
334Kkku6KDFNGQOWYtLyQn5FP60OsjmpBkRyI9uZ3PVrww4prGfhp/TS+OHs+eAi
WQyNJuCn3IHGstQiJco1rtlDqtn9lhF0mnmbVAB2aKDVnFnP4j54TtD2YaIsp9Am
WgllPP24LRPAT9bncWZGkLM7nLY4fdoMevIF+KhR88DG5pqEheu1hrUTAy/TWoHD
i1Ng6mnINHdBZxi+YIwR0BMBU0CcusQmIbtM6px2S7/u0O6ltMj5ffLf96m1b2Ev
IPboPB8VlEFmU7JgTDFdAk/ZICS7i9kbCk4b0hCT3EYCVvz7IOCDa+1Zjo+DME03
hcMmKnogH7CmhbLY5gxQQ20op7IlZ0ZRbjyD3chP+lOmyl3Lrc+Tp4Xm+CHfP2XR
hQytXvwn6CRSexpicODuEtQMP2n+XffifzmLpo9pawzIDRSNKldVqOLnlW7ZQAE0
9l6fc35eEYxcKnq2/8mzjClUogqbwAXffsBmUXyvdXRH49gGcXxFd0RcAXfdyvtW
1q6m/f1+xpU23bI3PxWABS5q9wCcXBMJomXzqpiU1VqnawOZkOJbR7mOjWgfcZIs
UmrOu8pkiwIEHStUBiliHJPA+/KgaHCHTV5YsVqRTCVsxs4F0Ieo1O0bv/J2Ybz8
QIG/gKgt562OHe+lGjBXamVw6ZgzoBxgQwsZBy+n45/+mfUDFOnSBkPybeBSxK0H
xgehnu/3W1cfzL6I2GpxCRxDD7R8AddzhKEhSaNK7XxotrRGqgoaO7Zd7CgbID8P
2TYuNl6EDMkRsbkLXRkjrGmmCYWiklklJCMUqTjtsLJHfTzR3JeEYAHQP+EDMjmt
NUJY+jbK1NmmZ2Y/dUqIY0LzbidY8cohV+YPhDrV/90dBkOCZ6Tmpym7qRQ+l7AU
VHm7uypBi4qeCFuoTmKVEQXq20FEdHuIhqATCweIX8Ksl3gaOInzbS39YtzFPsTO
dfW8aGPEXbSlDDrXb/hqM8q87eLlGzfriiahUVhua73U7xk6xzuic9jB6lvgWvt4
550u2RUqZcUxbCrMoCi8UesiM9v9NPxNMNKO+MVFv8AvRTWaCySAaUc7ZVpfyb7F
9Jt9+azxkRGA4Zb2M/dQBbNBW7k+eMIU4tHFBAASJRFwunyvaOoJN3MiyXRdU/5e
Zq4Tc6q6tTTom8Ja4n4YTfuiQUc1D1BftcLhq3vbRzk4FJvJP3jUn79PX5KhYGCw
V9wdXrgnAgZZhcfeAvKYwxEcyb9bHw3zVSY+VAt1GaTp8Y/UbxE8LC394c/3/4Va
OONSx6owzo4kAHEh747gAS9AqEX1bMV/inJuGObHrJdJdsqXESBJOnkgSe/3z6BU
3giquVjzyapJe9O8Ays2EeHjIv9XtcrBBBGuwkIxQ7A+Hb2Gc/Hn5Z6/LNr6kTeb
bAsn5dqQ4ZyLk3nW1gpxbB1yPwjM4NDSsTpBWMhvcZpUjyqthOtUcZufvyU/IudU
9KW5LCnZazwtzho76Au+utZl/y+kbtGDH+nyZwyFaZ6wrI4kVwO2+Im49nCYwppo
VSR5dCv2LRnwA6WKIG7IZ/BXmTzGrtCP5M2X+A+elzFf0I9J/6NHXvKgdMqgPGos
CdEMC255w24ppMczM7iJwmfq3Wb21PTmsk98C2gfk85vibyQYsKuRWEJgWCn7yUk
fcYM8n0wiDYd1qcck5o3pHa03mRCwJcEZuWMJvmk20V4vz9uZlBG0Hqgp3jWsUi1
huPA5y0LQydN/zWlHcrkFI6IM+5/zGlgB8Z6V7i5rpzIilBDDzU+v+nfCBR+qfsp
Bi2XgkeKrTHIsQkT6qgLDSHfzFhdHRsF9kAd7zKbIvetmKtX7amhlB17ZebK0cw2
gbOplFx5yFVDsJFRtqoauIxTZmZjEqw1RlmWoqTOx3nft6mOxmumHcpoqNCiARYB
UBj5tJIl+IbtdzdsiAFWvsm+HqZRUso2JHgqvgSV5vLSuVyus0glXSb0NkQOAL07
yCw+riFoLILC/GGJFtWybPQo3xgiB2TN5lZUujvIBNtcahTavvZzhEagBxK/0rTS
PxPlZsQq13C5Vepu3712hUCCPLXQlUXmUHT5UkaqBofrHmT1LovaL4jnv7qzxPy9
Y1PgzfRDwE/85Zw7CBGegRKP07FrXMdiS7cxqEqopqLQbXaeG4WRqXdiWFlh0FD5
c/Y4H8bUHfqDuZfGIE/+ntoG2q+L2rZwNmmLOHG9ONy/HQ3vLxdMQbfxxEcifSXg
HIMHFj0O0Uog1mDWCqSzc536UTdNJ9XXvFNvBLf/67b1M72iM/wVIEPJUMclafQr
n9aNUvmva3xitMivQpTqat/Ry8xvIdjpqO8qEAPjAlu0Z0VsKmiC+gxlE/iaJgye
zsN4w/wllPRe7U9VZWbTxbE9ax+Y1yf+0RGtI6C6ZswsM5xBHON20Oopnb9bbF0E
bloRTphVruQ1CQERTsHNzyCTxMxpQRe2RCz2rNN43SobwYN7TbzSVrgJn+4CjLRS
vvwTiqaFcWtrc1PlmT6w2GPCm3Ub1FQEX/FW45+cGpqeKU4wQtpOQTgwP0xi6t8Q
VxCU562Ccetlfhi7kjYX04l5deWl50xmqB7RjxOj/UMVlROM/Qul+QKpI0Cp+spf
RYx/la34w9KBS7WZLdcx4KZ8sjs7nexSaYs3KcgklSMB7K6Rn66/2XNG31W3oBca
281TqPmVVjOQozb7/rGjLpS78usVJ2QTni8UAnoNZAA97xuj4BTadBHMqxRoPj16
4Qns9TbjNEdEDmcu91sTwFEHCvejTS/0EC6HUI5DZFkBa9qSNr/15VglDS0bFbYr
U1cwfD49Vtk7BBmmhQ5jPIIlcEJxkBcVqmMoRH7Ixt16XzM3cktnw+C1wzWUHovS
00xu8mi3DNu8myDZpvBArFyHhGwo8MAULKv1z0GI9dPOZWt08qn2skkw34sLcVn4
r4DiynHSWmrx7oODeiIpmKPRgLJTDlI4rItiFp6gkY3yzDVGs8IytbM/q6IT+BSr
8pXcfIV0PD6oPQXFRzHjY0BugqeYnKVcDZBBPQiYV57zkOwiOR6738k8vziinnQ+
EUA29upMqygIfKMH40PY35F69nVznMpaM6jB7g3gI2XxhhuVxLWB8tHh3UkzRchr
FY8KkbgN6MrGaMuvBitzCX/Jz20rLY3bZ5wHUz2GzoSN4Iv9pYDbJJRldoMgGTLP
65U8+j/fTVO6EUh+yAKJIpOgait/sTCG8pwhiFo7M5xygfGcZtn0cNUTzpek5BxO
sn3Ar0kV+BWz3qYzF8K5dUKHek6p1WcjNSXcxtkVWrAXRRRic4xD1sIKSVL3M5S4
Pcq5yboqRZ1ERUSAcEcMBhtNRMGcrZlJGBjVPSHDSqXzxlLmrNordoqAMMRA6po4
Zwsj/dPEA7IqYF3tP4syUiwtuHWphMHkPMeRAfHPJQGsJ88glj+deI3EPnWpsYHn
BCrajgSfL74M+u+iU+yeO5TkWy8oPp26DHKAH37jAvSxKJN3Si950Nd6hTDnayT5
DgEBnf1trnoxcM5pPjmKLjZsX3nNnUwl21O6anPK9XWR9A2Yry3jkdwoaSnL6+L3
PIq/+ZxOz12UXiQTQvC/RKRTzxqtnhdjRiQts7cpNo6SW54jU6be4VlafB6hTef6
vhNOIAvFlpdSbV2PPL3E4bDpeXN+vD2OUbBkh+F5spEs+2YyMTpSbXjBC8aSDmGf
KOJnl9bd7wJZxXXSZKc1+T8QLhpMh2B0fGCqm94jja6o+pTtQZkXV0KMun1kG7vc
mgnUewnd1ObJdQlYs/AiUkFLWrAhX2KYxws7IemxiSRsQz2Wl/e0x9kkvhnVt9NI
yoTMIypbKp3CYOWOv+TEV//vXYNVZf25/We4jqASoj4DAmzNXntBRXsiH3Kx60Pv
8SfkbFok/QB+qmvY7rFhwixjq3+6IjiB9N3mLkpDpgdHh6ciUfNgdPNJ6ZtfxBKM
LsBch80E4g5jkobw+jzlGnIgZ20QEqSWOj/b0iDo0F/T+REq+sNC0ljerT9Mmpnq
GVOYpdXIvm1ktJ4P3v4W2PLV0wd+khz2Oz0gL14e5qoRDSi/t+0sY8towYoDoUkD
i3FMqNjhJq6PNlZz5nkBU8aZGqEEtmKz4rupC0TZDcdMXQU9veEjeXcxFQ63YdWq
vugtYdHuH5VDB0zjgb6nEqGw6u2hITiumYhvcrjC/5WxMmlDZ1Om7Z07N34es4u5
sIsdBrRnyVPO6stxGH1WZ+mwNbGVUjx59kU3XwAGld/7oJQBNmvFGVNVmHSkT2TK
MWuliRUrjiWpLjOHAzl/avWE3aA8RXjSGvqnOyGs2o2AdRrZ1roY9iY1nv5g7j81
DepTPkscePPROW2EPUErlDhPVRvJQqo/6irXNgwbL8N5HObGxYB++A2XNNU/KNGU
csgCGzbL//AUIsIP0nWiD1/k8MGWr/uDwn4RY+2scMw6GoQxlWrsozHWQr5M0d37
pua/JnpkBs2awcJk4PTgF48CjEfqsJ9v4/XDkomw/twCncIbKJRFxAW21Xy4E6x2
cQfru4Ct4hWmli8CvLlhnNucnQ8frP5PJRM3dKNItcdk4KITMhzcYnfZkssdr2To
OJQ4+k9X3n5KQLsPfBa/ZU/sDvM99Ov0+u+xe1dOcd8Vi3vwbQCe6b12AdjVsgwH
5oMPYu5i5TgFY7ONCSkwuiIxVHzYfqhhGOnwGDJ2O4QT6LijcxXARHdBe3F44+Eb
ShmECmmTW5sV9Us7ksCMCEpDvhEjZkwlLC/ZHUsHGWCT5RWsCRK2L1dUXBOlGoE6
cUR87vTTIl/uabtd4N//R5l2mjwtXD4J1xu9ihptt4NSeykuq8mZATK0k2ru28vH
LQW6crqd6SUIh8Q4QaV3nLTSnXPbWcOW2YRM12rqTyA/POuDWiX/BofD0TNcRd1C
b6mETh2MK5yqLDy2ocXhwwNNS75JSlrdeW32gcwUajJjBcoi9zBYVkw3Bib4fYTp
9zfuOVPArFK+YUHG/Z87KtUGwouEqofcCFwV8Y2pmgSp9YImacO58IfiAYH2Y/Ne
TTK0ooDBYFEg3M6Ac3CS1MF+AQKsXwdMZ6b0thyJpIIVGodECw1ZFRKcNZSVKg8a
VXiEss/RTC1LLMblI6o5rxaILZHCpbLYAEFkTbt8AbH1YKVFKbO5G7NzwG4JGbMC
oUmJw3KbG3rwfG+quWbfCS4Rw7Gr+DRyM0HNtulm4lQ4beDMlzi9LdvIol7hCgnc
8R9f8OXnvhLPwHhMv3oHklpyTYlwBgtIFbyiOVzPOh5cZxyxLM5+HS7JrAnti+NJ
iu7/OZ1M/MKOFXzrEDFIk5NOfV++dIusMkeacBz8GpIbcvv+IKLDuRFiZe+uci8D
rnEKN4toZmS4ZJyfnZ4MxKcsIizsVsbEknIVEIn3Sj6rBP1wGhhCRxhUZgor5nQY
iBZZHR6+WH30uwT/zqvmyZHqFuF6Jkx8b+S2uQiQ20dZ40gDBGH74VvqRfD7/C25
pfm9N35qrUt2C2x3ounTV0UynelLZr++cJKhpsnICyhp+seGx8ZzAAujC9Rtzb5A
s13SVbaIq2LtxlLEqnk9nB+VmzvR3fmM+Er5gcgolVir8GcRzN2zy/+EY11VUikP
6HPGLGFbV0bvNMhuqJQCLU5LSgvR4gk4q1u4CCQMC7fMmuuJ99WEHvt+B1yuZVV8
qotScHBC0CfNlG6IEOMMvQ9PLkq8gIOqr16NwuGTJz+t/DilUY4FGqHCHSOGYXas
AmncX/gvvdOZqLEM0E2DC6O21ayEcS7okpoI1oAIxHb+YK9dZh9ZmtJAHMQu+NLt
B52C6VUPtlSAwPTlpVtY7QlXoPCW6FfAzUO4LLrlkM+olMbWouzYcTxmkGK+auYv
Q+544vwfoDvlQy0MVz0EPoU8wofGGdVx78Q+Lwfa98/jDriGe8wr1TvsrmGhB+xM
ffMF/NcbHIDZuj25eCukHXTOt3ERSDp+YlcK42f6Vd8rRc3SNhAqRWkqrWgleptE
8uzwL/8uYvqtjCi1OpOHLU9hgHvNTG1dKa2ky3GGvMi/xGZSRdYXM5OBsYKyfeH7
j0TBB/e8RdAJpgc38WtBlY3HZ7Up0+MaPP9V7J5LbhrCCxwAFPLkJ9BPAEvw7EC3
0hlGntttbcV4LZoLZbS6QJcK89BixAYuMnav6G/uWt+nvUskjA41qeYu3I+UK/Bj
RjY+VPIyrzwlRQQE9nJXyjZywgMZYTxTgoct4AeL91JLxgIoMargdsvI4h/aPtq/
5Z9oyaDR9RWmRUUP2adqdorv7x/MFbHb+83k4NFK8kyCkBuhvVz1zTmOO6FiaOcH
pNbkH1T4oDtAk4P9sim8QTExjDfovFI1sD9KDQ/VubIVoLxeErixie+cESDTV9uR
cYU2RhtFB8tTZFo+bngJiC86xTkqKwy9RZpj03kqTffWf9ojru2UH5QBWWzF1RVg
RiSatYlf5VnlK2LVp1+GmTnlNoHI+CMVGYnR7Ka3k52kF2/5AmpUU0VS8Da4bVz/
a8H4ISG5QnjqnlbozW1kgVn+VrFbDO8N896vTv80bZHc3ouulhokROWXVAZyiVhb
g96TsQBfK3GVNWPvv7YHlPVwJpquSX5AQ2flkIkxJo8+j5Oz+cZzTo+LOIMZVQUL
UGG9QzP64hIsXWjf344yOc/QNCTdAeygGeYtxmlkmquLA15QFYEl3tAquf91ZLoE
K7YNlf5V8uTxecYmaBo+a9iV3h8mhY2Wpk8g2Hl9uqnyqgQiCCEKpR9l3ee8r0y0
UrHqcjo0K+HobpBAK2UC2jKNg+7+xTdFmJiS+zYvd8XCumLtbt4hp+zWj02knXKq
Hd8SOpYDgcPzqENCN7cFPGCRBVvkG+IZtEQJzUAqHvI/OeoIfib5s95a7672VSfH
1lk0ZSPsBZLbmWPeGqCVYYeTUVAMHkwK4EBfy5X6OjCKWKvgVjjyMNT2lpfhiI91
nAwdktyU4IKHLXwjqq6YG9kT+ql+JNoVRqoKZjgxqlUIwrO9s6raQieGMewJdMd4
Lpk0LCJDZa6otP+owsrPdAKvCAmmDSgE94E6hHfUASM02hF4mqr7UGAwsBS7KZ1C
PSI6BYkTPRcZRDgrnO4/2kFGU6gbmhC+LxPj5AqCkk8F5W1wKl6HAbKACHhLSRc9
dPTBozz9x1t8psNm4Wii0aq5TqoR3gxVXM//4fHjHDRl/pgoAZznnjWhgbcWIDAk
Z2qK3dIy5UALC3235FF6/1Jopswot6/wVdWVaAd0NG56ig6ufmDLgWFAegyXI3gj
qkf0FS9kn6tj06q/802rgoR01t7PCuMlKECJNVyDyuYjV05Z7OJKYoRzsZT9fG9B
Hscuf29YHfahZxvdos0rRNTAEkyMSywT7iMtMzZI1PXHKhKFHugqQPVHmdhXGEvy
Berb1HG32vukfLMvaGQ+0ljLYCNGsp9y5QRcIBLOX1qvjX72GNOJUxK783qadgV2
UpbnNAmVErPWTvYPKyXHOf82uNaV6e2tpb5RQE4bj5GqSmKddsXsZYsW1rvopl8R
xKh/Rxc78trKQI+tXihOOcu5d30sBu0K3sfQsI6SnrT5L6ZkmYgBI+7uTL42lL/W
bz+CEZm1FQi4+J+f4Bdj2c5yXb8FPQHOftYkVOCZN6UVzgtyqEYrkdbVbSCJOPqF
fKJG3HUL9VZEXxIxGi+u9bUAUZFdseBKE7GXc6m2RiXom18SI5EOCIAkZFF7k8Y9
ifeqPadpgQlDGDCywCDqSiDZgflLgblmXlK83/SglCX7AQs6xtyELZ/9zdlEMuPt
ula78huuAoAsLnlLsRfn5Bk2/2Fz2CcIzf30n3UVF+/BPj/cjcF/ps5WIhtCqrD+
ikmq/XX+BICRQTwbxOtH0IWpUqjcRBMj2KU7ogUr5RlLxdcALxnc5140RJf6n4DY
xWCQc+URyozFr3cQmlS/WQ90wgw1IjdDKWfjM0Pc+TEMLMPRu9YWHtTY2NF1hjM/
UBDqSGPiLtBTuMb/Pdbskjq+LgMKSjonvP7sQs6F7eoLym7RCskqvuyPuJl0TExc
dPwxsHT5dPPMFafM6ICyE5VdSBzQG/tGZwIhg6GFq5ba7n0b2covVdXKi6sEAccm
khMajfMicOmRYTTkvYjP2DkgvR/RRqysmSVybKanG510f6GGau865lufNCNtWVIQ
JJDc+T/znFXhRRQrzSCiqxDgZKNhV9iEUxu7xqFKc9sVN+zC2pctjz/AegQ+Txba
emlWgYIqlNEGi7vnygaupX1cwg1/3yAFAt5VgdzuQAxSljmJaWj6FExZQ6Yllwsx
6+Wdw319M1dpYxfnL94WGpL4Zmr1yTlTi3MpmOeOc2b1/5PtLdKzUM27xMSOKUMv
HeNa80Z55ftZb13JnGZx2yPm9i8C6fa3Lg6PrX7rwTk35rmxnnohKCH9+u6PdpAb
LRKaf07n4cbdcl4VoCnKBRkcWa2MlCPIht2GzDxWgl3leoLnBfvtLwkVGAfz/BnL
CWVm3qkQV2szaoYhHZIp75QEAmb8+mv6OiXnioO2joc1kUD6bE/mYcITUcm+foDg
ZxQnic26mTtD6+Cl19dWPsJQ87XRMgqjVvqnpO3KbCBEAwuSgtU76yGJ3U7HCRRc
r3b41zjgbGl/WZnT6WRPJAeZ+7IALydk2rQKiIX49y03kqedQzjY2Ae6HYFXTJ5a
WlL4IAYWUg8h4WYJaQsZrelssZ7pq3HwFvogcz3duzo2VhhjHRxMgGrPVcQkyKC+
AAaw0mP2jDuRnOOf2msnQgYjiCvZA7Slz+uRfdjVhSWS11VWe9MT9CTVmIajo/jA
UUfXMr4CN+1VqliUHo9AMjKuqONvry5ePqop2XoClY35hLbMSm/xzjXgmfbrfKLv
Mk/dvHZpbZ32Jz9HcZ4fWVY1ZkFMx34zJ2u0rgDAvpa8J3cGe8DmMKN4K0yUGEL2
/8ZpATzzdKAk8sHlVEJGFZE0GEBMj2df5j3x1goXLHK8b5DlDRu5Lwzzfm+3+kVN
z3EOEEkmw/hgjWxwZDV6AYwv9E8/wWXCogn9L9bl4FiY65xzkD3y00Akcuj6a/Te
/x61ScFkqJgmb4Ynes7tc5tBmbcXUARQr2//5dKXVH+KBs5gCTkhmFaqeowfb9DC
Cfvo4E4uy+PUUPesDYEIsgDj8iPcIUDPWpBPIorrqe18OqLFM/D0GJnPpKIZRShY
6R1akvMhKeT6q/h6UinnzzeK9INlobrex+HqhouRs8T8iLqDgdOXHYgrN/tBlTAT
wHoQrd//MI0CbE3oAuyDEwX8WmxdqRYHh1TLDoz1RdgiuNNIWZz8sGQR+c2dDOS1
pcNMqKv4BINBP+FVLYzH2zH/nLde2Mp3d0iMfmgB3W+nDsumvyLl2xCKepWSLXtt
5ibxHUglfRaIFpLLZKpRjhb8kwieu9M/A/Yn2VGYxXEENZNnlkK0rpwJoNY39eC8
EAGXnMBpXwAKe+EvenaZMEr7UAvu0kmHwiYkixlZSu7QT6s0jAZhg+z5vvlTzStR
nkX2oPedMU811+Z5vXbcNlQDA018uir0f7zNOJ0x8birGhfVHu/YzgNvsEmHA2/G
XBWAj8LV0ZAuDHr1dw2ykCWIsRDBoWUw63lYp17d3+IZWDfJnW5LwEHz4akpEcZk
NzaidR0UEbplbNEeBp6+yEDOLn8lbjG71A5iFy280Xfe0Tp4Q9nJaDvTqxJMWWRb
CNBxRwYGOGCCTAazXMI/nqigTe1+QaiMlozsmHEfgVqAPiJVUbgT6hoep5NvshRk
g3m2FZ5p7thB4CX9o+1esbHJhZXbU7IgdQuxSe3yoHCcA9ioTG4Cmy+VS6xwkoz3
XlgLl7WKH3ct5/ljRa7UmU3GNco8WX7I7UvAcrUfqTU+xWeJlZ6IN5vlPMijAIpf
uXtOzjRnW19J2tNFtTF7omfEWic2rMrYQiP48ML0d8reTSbqqyR3UEpkoZGJWTp7
vC8wrwnKUlfimlEic+r9QFi8hjAbVhW7doCJAGfzVczCbed0IGkxF/J6lsuYVq7G
9q3ABI/6LB/CGe+zPuNorK4GwmP5Wi3g1lMKW/Usk2FcHtKW6AxTkkLPv2JC9fXF
VcCCKnHOsKOnu895NF3fStrZIlq1f8dsVfNwjDn593HbhPS8brXWxNjYZkENROCm
EgyD6kiBX1cZZRxE2tfjCOjypbKOQEuhL9hC7niW4dgTzvsnxPXwUQKQplNxCWVe
d5pxTazGeoRPkS3MkHL2dvoKQ1ZKQbEYBdxZEEd4ORmPO65ZiaJemBHCPxdyafxE
/YCxEVT3/Mx3pnP8UI9h1KW9m6yFCFFrOtA49SyIIdDWbEtNDyRISHnljPlU52gV
Lfnhvbl3RGnyYhvrO2CNSW0WEB05gPzRgpTsNLN3NuH2UxasqDmxBykBWjKtJ1vl
ygVjnxnFKqXypvOSUml54kxnGPfenpYWRuodyKsqeLq6IPFJcIf4hzCKC5G+zM4j
BUjaK52qzGRDqQGrvSiJc7yIAkQZoeadMQSvAcMFjrX4wKmHKzdUJvswKbZaTHKc
Q7JTy37aWNZRCOM/06kRt4ulpa52ppnnJ5fjdyfqA9DDUgQxlCul0bUMZhgrLtcx
00M+fqA/K4hF7z+eYVbsx90GIGxXeaIMVyLoYUFWytnNAicFB7mTSi8fZjXZZLp4
+oEZGp+CyZN7Ky//jpjBLqEm2peRG8IaVfe3k9a1giJLKz4adoZ9Z1ZfC9m92gsf
yjrC3F7bm6yyvlXilNt7Hy3XP5oqhL8tG4HgvvNAxX5Kn2gEeN+ShvGwYSTutkDb
7BoZWA6DoroLYSEebPHwB2iEsqMJC1vxnlvdlAi41PsmTkmRFkPyDVnfBqZ3ZKPf
Fqc3u9XHgJhQYo8+d6+eCUVMz2QIEubduakU4hQyqP6L7Dm3QLW/VF1sUlj0ACVM
IagTFvRh9ZMUw+Z+7fvkTScxYgjWhJzOYJC7Un387bulh3bSLSi8VAvhc80gtnhu
PqYs46iBWoNOz0nNOosZdimVNDMvqmygr3nh73bEVAT9Q58PFPUfrEn2GZCGe1rb
WicmNlXWli+yzp8Sd/UChb/kXsvXx68gZ2HdppRY0Ln4ysZYKAswn0YLVhQ7witT
iIOzmrYO6tfZnJerT5I+0c19AoG7tqSV0gaovzIQSkNpNeABTL02YX0/tfDHhKpd
ialiQYYarKel1z1HQehq9N/xi/YBXq9CrFl8vRV5JkanZDqn24nMMkJ8xpb8pnP5
5HNhtz5OD09H7d+kx9NAtll75wRdwkMZvfEq5/Bv6m1QyfZ5gg6fDfRR+anF9yNO
Ri/mlOfy8HtZAvDJA+SY6hMNbvg3+a5xiuHg6UZ8qKz2AEnH7e22haxjsBGcuvRZ
yzo5J3bAfFZX9nRr4HhxobQAQgd/zDY95iDUzA0g+2S8+YcjPifpaowCElpZbONO
PF66h0FpemvIEFPMFkfcFiEB+s0uj1CoI8784Zphm8+tcMrpMFQgXrU08xzXT3Qu
UvmQoFQ3az9IvqIdNuHggNiHsRHcaUimNw66MSsoSaJ6Vw6GSOgMZKZ8NFhxH1ZQ
Amb9n8f4XlN4m2yjOOyx8Dqv21UW5GOvE5twjq6z0TXhYRcAkDVzD5rtEH+mZM5t
bCwqPFyPOuKFKMhh4v19iyKUDkVgG0SrW5wW1JDRnVNQt0ej7QfaWiST2sFDicwJ
7ahoi6NMgALhdty4rLgpd5lOm4AkmSNbBo58KQOup7Fgxm/k1ByzZXdFp7iJ/WYr
GPo3A63/Gr0MZHGRJwYBNpBwcL6VV7dqlbH9OGFnKf/2x8M3jdgyOjs5deXWC5jP
dSb/K9Ke5zA3Mb/AHpxUwyzi8r5kRDUMQPBNhHSvC9m8TfXyoZygM7lptM6ixU+D
3bkohrPgXZt+7V6L2NrTZNNrUUOWBpFtwcDdQ5hjhzTR0prtvIpmqr11BzNAOm6H
wpn4JNIHKVb29WeK4r+HmsPg44sEM3I2S628ZgH52dQ=
`protect END_PROTECTED
