`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yK4fDJBg4YT7So2iGSuEGpPgB/BCRd1/5ekxmbYFpLtZqnlEM7zUoKclh1P5Z5Zg
/oAbYtmWC3sFJyJta8dZ124z+AN/qPWBb3FZvcVtrDOF8DgkbIPziSejZNRv2vqv
CmciaVErwuzyiPuxQlEGkbyT/rs6GorizE+w5mKUOXGRFAJwjzbxXrK15Nh4rxA/
2A1GewAg2+MJd6SVSk97h+nlQi0z0+iev+WfQp76uONRsjt8TifqeHeDmrfLKhrx
BqNetURgOMFMQBFYY8vta+gmIrsYA4HqB9DyZSecZpQcYqbZbnAw5vUjW67d+LrM
GeAKygossc8BNNC/uwFeU+0wOLSn9qTFpofE5ktauEWYj2iGoyWdBiBIonJnqMey
dBbC5xm1skUk7p0Bw1rcsFxm0zctO/kO+zTfpyZEkIoDSOMPD7Op+UVRuUwDsvqV
qDqImY6zj1qLG2yXCARnkQ==
`protect END_PROTECTED
