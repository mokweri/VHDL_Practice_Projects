`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXbbYE79FJSD1eoNl0kkq2eOK7vmlWIsaF2m6QYZhEb3CQT4p+4jv/XUGUE1BB9N
Key+TSaabU5yMc7MKCVsObYjg08gvQZFpe1g6aRloTPFvrwSyCDd9DgMAHR2rbV1
6M4QPKiyZaKDgocNZgih7z9ALQ3pdFONqFueU78iMMVbrYPXxjgqNTrL9BQrRlFd
hyShfTzDLVCwwes56eBdhOYgdHbWrhNpe4QID9MaTY1djFLdpnu5aQZZ5MJ7lmPK
NCXw7zos4j1Girpy352OOSK3Y0YYt+GGx/EaEf2kgiabte2vdlU/zVtX4Q3EDkph
iGsyPP/El3gFntRTvQv12rIH0654T7SOF4Wql1o4OVSQJTLdEQG8g1xXJq+KIcDy
JT+Rc4RFa9nl2945EjTxpyfi07+mgTnuZCOTJ1UkDzGNi5/iMmXnYIPNP5h+Wcvq
VTQ3yfwky3Jb/vAyMoXlqSOxDHfC41//ICl8TtOQ1Q44Xmm3Uf64X0Cv8hDyPzik
8oXLlIpuSBZSPhuiLWVhcEZtl5HwsZJf/QBff/SjQsBs9zwe+wht7T5vhpoZkCcR
zYdiSmlPymsdTMX23e+uUkdM/HPbGdybuGa9jy10HHnemwUStIZqLeWGb3tH15i4
xBvlz5Hw8ouUQhR7+LnDEIZwAPaYtQo3Cvmhj16ckGHkL4pzRUHZARgHKNIVMX0q
wOwm/zmxsshdY1n2mSScUKE5IuICkDhhadMfsEfrURnD5B/lim7zl/Ok4UKZmyb0
GrcQU/e/e6FpdZ9ZBPFIMigw+1oME3wKh6JkT42bn9tbPjDvW+IdZZFxZFCgE3Ou
wf9E4xZVoDqhm6f0rsgkntegKD1XK/Tu1pB4moIQ8+soUXZsD7D79gSweysE1ChS
19kXEUvoq2+bVpDjD19QrRrlSPzpdIuUMx68ubVyJU8BHzAi29+vMG+fTEnPWtYw
dlfOV52v6A3H/JT0m8sQStUhm2US/kub5M0sr5z0EfdLMqhKDN18VWWbFI4ZuxQJ
Q4bogwTOO748DNgJZxGLCBlZF7515ZVBtDn0e2yTwmPX5LWdmfRCdSeqxhkFN4C4
ehg00Iym4+XdEDu/EfhEd8JYUGgsMaQtbFu2DaZCsCKvl7waVsCZ41BjMqxURG7h
3ejXoB7OxQRcWztplsfvpA9TtSg4ZtRpcLv8iwcISs71dvUZsFbCUSzfb9d8OcZB
qzQA3I89gatZr5jKQqGvhI74Eun+V21/JfewYpDYpjgdg0A8lNOMj7dEpTBlKF9D
xD9wg7k1WTr+iymxrv3FVJtEG9h4ejBTRUjoQ1xqk1jQPN1YvDPXBZW2AJwAFbiz
8jyqriiePA3WNCqcYZwxgQsNz/xpWjh6IUZaM8uxfc9358pLEyXVq2aD8D6iNN2s
zLfGd/XIvtdvwfnojSSAcAlFRH0CJ4frgb8UKTq+B3aY8m5pSI8bxlL20gAyEwcS
`protect END_PROTECTED
