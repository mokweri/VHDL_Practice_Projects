`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iLTO2xMThztnjpo3B0vphuERsZA6ZmXTM9wwo19H52iCWLsKUVbHu2BFCRZ2W2TC
mY05mOIpt+Q7jLKnOHZFs6ALn/lV/CrIsqfoJZ6a4hcCb4v8e4QC3CsEwW1yepM/
dR4ojDj6u9g2U6hvI8vKn4vbdB2HHrWfHJTTqYJfaALLz/KfQW4e/fa2rULhFzA4
GajFDBOToxmUL5dPaoyHnr5L5oY16FqjFHSA+ugf2EiLbFm860cGFye94lb5riRs
qurJmRzg+lkGiqX6hgTkLU3J7rd6IXwe2fcuGKtDZo8uJy7ljnBXbE3rxTozabWE
BSQkoTW5t7fsdjVcSbzQ3rolTgoZvaiNh0JAZSO939g8vI+LNVscT9+jaIOm7cG5
ten0QbxJKDY+RuxmXdbbpIdT6qp6WwsOBGIfNl/iH5mdR0RZxCwbIclT3Wn5xh6K
TLQBPu3GOeiZXiKf8ZMcym9/LaQWnUZJDJGKIaOIS2vTOJr7Au3gKd/X7MUTA8p3
EwSW52o1pSNYC/edcWlDeJjbYynJGjRVWHqReHQluSdqYZVhX2Ge//fP1yBpecsV
2hPtlTRUGvm2pl6UKGaYZ7L1HnEuJdqz4MdddeDzPBBcXfFZfMVypPy1t4jCD6PW
snQTQO18N5WkU93Kocm/dM25TUc/nb0chrH5Xm4zTNlsXF6t4CALKQagRdlk3Kto
F87eshETraDDRR0C2pb9IWj85wzJFVO+/IhIzAiYp4A2ItHtH3p2S+DrIxsgB3e4
IAWOZhEzWHdGB/N4ztojvFGWE6FxhTAd7p1OV7/iwWvJfmzAizVUIwFTIWOMyvsU
0SfHqU7nJPYN/wH0V/EoaQ9Ka5586Fuv2OWSHx/GxVZcbYX46FmGzd2AJEonLhQQ
F6jo/FBjCDNEaU7ODZ8szg7nKzlcZyUtgfpZBvdZ117A2697d74Q2ptFiB2Xu3S1
KaWRZ7ZSE7JmD+ilGYwfhxe6lNs8IOH1K0UzpaO6+Yh2fRkTQrisirDrHHKW+Ldy
n+Iqx1dOLYZLZugwR7uLbXTMh9O7kV5Uoo2QvKVlr9X/kbOtDqT1+Qwk8BkcO24x
UV1+O1VJMrCstyW0mvUIK+2gPitP10zI9CQKoSFqw0TUjuQJ/2wK4eaMLpUg93Ko
gYQzzXJ0QQjUzE9b1/wR1po8P3IcZfWIHd9A1Q2epvBveWf4J5AAmIw/KoSwwOSD
lUPxn+hA+PK0ZSMV8ObL6y7XKndAayzRrGq+ECy24qq2f/TJLzwFem3elE1kYwEz
/kP0e7yGSjZVKYzTsg7jpKR2mYKF7B39qkSVAOOKy9AGWHKFQ1tZJpk0PgRXltv9
50e8klsjd72BQWdaN72a9cIxftprpT9Y+4a0Ab2tJuqc0AW4u2SeGVg8rMG6m4YG
o6pLJN6HUFggdZs2pZNmAI/tn7cKPDSZc+Uy5teQRO1QZvuHiCTIqqpa3Q4APm65
cOSNsp7SWUpQmYEmI3OQnYrtS0FW48ISnbqrunr8LcmB0op4QM4fJq5m04vAsdQq
VxiK41ws+LXhu+fIKCWj6iyDBJP6M6JtrhPn5pzpTPnzNQx3PLysgrYuKp4x9/tg
djB+Hg08iin6mFocU42gxkoU+9LJu1J/h+SzXEOdAljI4a3aVs4uLYX7mHa+xMxG
xuZ1j7JphbXkw4vlqP1IMtgvsotxT/ijkb51KPZG9Uc7qr1YZT7Id3uTR+maPBGn
3BLQFqQteTie77K/ZhrKmdSQXpKt85xQIk+GRCg1KIe54Kuzc0ggkUhw52JB1972
XSzv4bLE+nDhkhk9DE0H/zHPdPIxbOhPIwP7TILHMGck0jvLYsXDOMrMOeVieWVl
SVHfYjCelYeVJRneE9oQnJpsg0XDLpX88DciEk7AbLGxxLShjbnH2Ln5liojeyKF
tKWwSu8hQePElssXTCNpja29FYR8ocnivvl+3SBJkLnqa4Pkb4YVkJXgORbhnhjb
fPcpKIOHjK+Gv5WYOcqK1pgxv0ljzU8f8C3Q4tBk99/RgbXmOc2scdiPg5TafD/G
H0iH0JJkmrr4NqjHiwQq4IygBij7sJHmaSgOE9FAW/w4RKVaQ65QRNG2SDAmtz6P
PYX2H4e5kLvG5DP3TLwyVwygF9pRbGguGpnuuwQrIMGwkv6jQFm7IQLxw+h+0RiR
NhDetMjyN7iFQKgBs+rqYMQwwHsoURhAh6Gh2GFMym48sZRZUFDgSniLdNev3oGa
AwSFF6Prqs1l/SYbM2Rv/OGkB7j8YVQTmvT3LtfTu/F7cxkAjk1xo8KkYuhAEoGu
B/RcOVnDdMLsyWOLkGZ0Ppm2qcx2ZkoguKgEy9zq/cnDPso7SF5L0GXxqMADz9YP
HkYWhw8g4ydDtXFFs7n39DsSSObriA8brH2zMYnf/nMFK113g3ldw1+bMvwTojrM
zmAtJX4ek0KMbCuDQw0W7TvRLfC0ABHrO8RaQC8QQMOkMsSan0qTVA6EcLosHX7L
jcrjFWg6Jyzz7GI3u9uWuGTgQbhJMJ0RjhdomvNaCHUdHQELz1bFRBbvaCAUUl/6
wrHMTeWdcx293zUnSNmDEFJgMmOWJbn7KH/L7EeVHIPtr1d4DqRI3CmkkeaKCcBe
gwdNG0CTBKgkPVShJfeWSkH+fuzFOzVIvfK7+pgSiX3QMjsEFpQkLuO2qscEKY4s
z9vJ5OYa4lLBEWLate69kChAVR3f273xvCl4Ibvjv2R/XezwCf9i1in+n36We5dn
vEeyaprC8IPhB11Cqzd4v7NKoBLKS46pF4FphRgFSdqz/ihA11i/EV9yc8ecNRSg
BW2XyGlH5aPO0QzM1YlsOoX9FRa/N+N2dJukLTY2HsxuHeqZQ2wFP4IApyLYTlYR
HfbF5RtmSmXe0TLvWHgYZKzYOGQ5eCNi+1QXBk0kK+DmgeOS000j4Lfz5bHNRhYL
zwRybEkuwcW3EYY8620cZ6saVaP5gvQGMg+W0P0ctkGhC3mJE16TjGwt9bcOUXLk
a0RI4a0/ijG8FfqukzjGAtcUaOZ195Wt5oWmgi9EkUuRmdhAyp8UdFtlETtY3k6m
JpChwTxRDmzqIUfPhA/cKmZoUTHmyDPaS+bWe/UUSsv8ixG1XcnU7vljaU58d8Az
9vczKTGtmxEh75jsPaaVGzWeQgV8FYaBhZ4rbTX6DE4vtuqN4ZNRjbgi2XkRJkt3
Jm05dXdh3A+Ux3xUD4Ax+3/v/X/lLSBBah4nmSp3vRvDa9Tz82EsmlT72hrzakDk
87p7AjEcnBlh+KH4sT6O/doLfVN0OXRJrqYTG32ik9dXLHxqTr+fi49hOvvHBFxy
E9ONcaR+vS39+i1hfuY1+Q==
`protect END_PROTECTED
