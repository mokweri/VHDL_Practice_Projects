`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXnFNjm3+e8ODQnb+AiEsaGTQGG1dFOBr6WvSTH7AlmnuWlptuTqX+kYCkSLPvhs
yWB4U5pqg/RKLM1K1AdKnR8QfOlmmSJYP7XhVFB+ooqxuiK/VTXajKy9m5vCUlp+
2bg0NcNiCOOB5d/iNyQ+2eq0q0WZCy+aZnX9ujIjE/EEbcrWoxagicNjUzQV98sx
lIFTlpVsTHdDXZLg6xuCdWjJExlCiSdfVBvkc7vlK/XU+mW/LAnhSccy8pTeSDsf
XV68KMJBys8yZVmzmX+3QlxK31XPiGPakWCX5FmlsevT9LnRdurfou3bPC3lpzy+
rZLeoBJHtVchQCJ8MRu6QRf4fvPXjlrdLcCQLdDjQjVlvZxWYoD8niv9FQ+0qQJV
yMQN/vCP0HUbm6sTPY2VsilNHly1Qey+BFZE+F33sAeHiYphNTC2JuQfdsSYV6qT
hC2twc9Ad8p7FQnjRTxgMDS7SSbxEERUF3HM+lvCeMTfO+cE0keTa3mXDXwghERB
JSjx8v4bfJRhZMaUVWJcEPcdqE2ywBN6N3uiUnzXQ/xmNcxh8sBP+ivt407Oh9yC
lin82gei2syIubNBG2DSJTsgkASn/kqhtEmexyD+AGcNrLdrhJTbGDMcyzphxSFe
jThkoneAjueQZsMHkszM84Y7FC+lgHx4tRxD0eY0wO516gZo103VIhNeTgiyAQeq
BxmVhWk4NmXfZas7Z0IojDqWPWPmE1JxRltZ8hs87jXc1WeZkk8t31VsaUlqVEbO
vCCxaSClqThmQlBjJuC4lz6gV/OKeanty3eme3g31YGRMQ4ffcOu2+QhK7XSu7Rj
GWE/JOMu1oCft3UZE5GBRshxQ96qiE1vrIzkY4S0tyLsL4t3GWJ6jh18H897hAji
srVcXf6V3KYyLdiKvt6A1ynf2T1keMecsBEfwZLasduf5N0OxPzuZk4Oy7Q0la5S
MwhxyIauEuZCpMD8KkyyHggy96ymYfm2H6Y5uELb5TpUnDLLH2gtS0wBftr5H/EN
d/TUW8nwy91YdeU+yT6quuJ0CLumHLosMdf7+zg20l5+lIa014HMZNolqzL/Xcqf
N2m0rbyznzQ0PcauymanOoEwCebrhLxvPQnwUHODhepBJROKh41W6WuyzXOWWhTF
VXbh06exMPMdUJym6tZGZfk4XJeDWIH9V4bOhpDraNGY1+6Qhu9Hcc+XRdNZAq6m
kkb4gSVsf6MZCQVpfdVfMQz3rGo7chOgunZZwuPkFZpzayxAdFvMdy20Wu1C7uWb
vJIXtVP8WpQH5vAVFNsV1uwBYmS3qy8KW2rHgTPIzth69XPFR3kWSHYQA+hsGF94
6jNUnFu/V5AF3P5sE/4BuyqYN1IIwH03M0YHJldd7K35XVi0PLJBcz1YnxMY1qiz
1CsQwneReNHG9yie1DxZ0vtWHg0HlECUhN8j/rAozOhBJsczyTjbYTDFzfLuJ11t
kYcwquod6Nh8rmkD/H8Mk3+ZEKJkGCTtOD0woICdbxNwhR7fTZWuWEMBwDt0tqA/
+ADzCGsUsugmppTtvMZ0PkTJpQxIIvq7rwy9eq+ez4Z5m/6CAU5h9O8xoAqKCzZh
m5BWZNtxzWKbUb1DtWJvkCdIg+8j7XhFxCXImNrVeh7lnOscN7jwQ+PwWkzjeiZU
05lDGc7eymu6aUoHuMAT2aEqt1bvY+tK/eiKY0w4z6tOqIK07vPpInxliLo+95CW
anSVRA7F4u4b0JiHGfHWL2/AMSLTkVA+7L3E3nAXM8sCYzirhX7Bz5yWD1cJOVVl
g3AxqCkHaR1Gb8lblZM9Y0gZ1i7L1cN2a2CCD9vnZbieusec6dzY++wzQSm8DKaG
fi9bDY+Ha4GO/96rMOf/i09XIVET9ugtiQnd4NhKFY4M0heTrSEPRRWF6LfT1UCt
DnN1ONoIQJucF6VEnKemMtdjkKb4j24xkfXMhcXdNJ5XNiRYAbdH//HObmTRKl+F
atuaeYeSaG9YqBhJZ6N62jsOjT6iMoUwcESKjCwO8fnDDwHIaTbGSm5zC+L9JBu5
5bC4S4+9TYJqYsEzVWjwM6a3Vo1EqY4GhlBPZ02LPOreQI1FGqg8p0geUTsRiTwU
WNRekxe9vUP3ZAE/9dgt29cZKlI0UUQf44TpwlJLK/Q5SBL0kzOQEGlh92Dr6bib
Q7vo1x2qQ9B8H/cYCwXhM2GsgCZxg5erBG8xXJjsRv6atrrpi7BswyLgTLHIGokc
yy/lDTakeHBmOBWudHsxiekSQsC4uffmIFGcKCCm8rw5qBvmMCp0rqEb7w+v+N5Y
GJZ/8GrppnYewRI6GZdJ0WfmofrtewQkSqZo4JoV59Oms4WlgP43F58hqNv88IIQ
TKQD5SvbRo9khvvZWDXt5WjjLVnunrD/k1tlUMaCxPAfTzGL45ErMIz4nRfPmb8V
AqEjDmHE1yyKbQeRJIVlqGlqdqO3+vG7ESv/ygPW/pn6yfUjOXp4nPlXsReoX+c9
9juKiiRcLVng4/Pz1E976A2bXiefqJ+D6RAJFjqsZEpJtDeXywp9gzxnFDj59ceQ
CoTJFrj08WSw990ozgaNjx1fBGC2aNrA1S9NGEvrbTJtQPN/bsZHztW93maaLn9p
Oc/E2xvsverC46Z38O5j0L4E2KFmnCrSv7Gv1I30aW7zNrtO8PQHHXjfQdsU1bws
szre9bC3r+BHBq9re5zSqikGTxlNmPSVt76OL6Gier2JvP+DFkkAnxVmMxitwjtJ
jYgI4cSv+nY+bVr7lJPS7ity3dT9TCIAhpVIc3KXijFy+L4IfXQEfxDI7mkjuAet
OElXrpOgBhadBVLK7KeDJA/7u4AdpDgmTr7UlDZpPdn+y9c/WtiLPF+kv2QDYhL5
sF04Ko4/xUqvc4AUOaF5qhZqlDWlSUjMvxitMwmZq1r93XYeAbTnK6WHAoE3imuC
+HpsJD0vZtDJyZScqM4b8XlU1q0VAD2LbXKUm9InZAIjnAFNdgTvYrTarSE1p3vP
h4cIU4lxtM1Ve0rCKPROwwSM5qNQLQpmLW4EfC1QoiYlUAyezeKd2B12hQqFbEk1
Eol4Id0VtHAS8BP4rWJm2Dvb+bUR/e4S3+kzIZLPNlLA6kCAuQAB4do7DfPhKOv4
mV6V0/8nF5ddv0hF+fQ9ew8+FBZxoMGHlOvlmAZMHU4r/kLRArMcbsHVyXQHzjsJ
ZixGW0JayJ8n3rXJZgrzQ2c956c1VdKuIk8l3TiNIfRYXgfEuC3+II2/mxh40Qw6
IDGrYGY3CYPXYMO53/j9tfTuWEIwDbk6Pa49Fb7FMP3pfHWq2OMVysHMdmsXb1lf
ao+TQzHwumD7hTC/vb1W5Y1HDH9zj8MkVSeomlvPZj4xKcD3EiyCilVIa8TDB13a
Dp2vH65aL8lpuT1/IhqbwV3puGsgQ/AWLTDPuHfO3wHXlgGOTYHm0GkfWtAEqL9n
t5iPbFOTTeQUo3E5hO9K5n8wtcOBd2WFSo83YAqJHBk3sTaDnJuhQuNAeZK8aQiJ
+wcpE1STZCL7hyM3ASoVrLrpL4I7FAmGh6ECzPOilMPbVn/tgftTyduyGoK8bDmk
wHoqfwLvKpOyRH2aI8bnPanfS0dGZNpvl5LIpFlkEkp9EXX/wFrgUAj5CsqZXVP/
aUxwrsw6A1En8SHkVHpzkxXPlQerHASyisnOCv5c2ZMlo2/dhclzv1y8chQCtErx
xn/8XfmHok6abC8t4P2tZkVT+eJlxDEVIw5+IbRb4leAGw2ZQ62CN/eUvSIX77ui
HbUXpN3L8OTzkJjI360mF5n4Wbryz8j/X6qpMx0tIDWXWF2W5bHP64izIo6wIhoN
YfEfR+o8MRdxKtIJB8fJz9CJfGXRomWeiB5cdslu4wi8wAxSTyhuMwzUsZjY5WZn
U3dnAXslrW6WxyS2aM9znoHWPEBaactGSJ2jEWECEmg///mGrtIg/GblvJ++d1IX
RB4ZaKjglDVHWM5kPdDym+9aIz3ajUq1L2c95o3auP/a/bLmtdRKAZI+LaP7QEJP
ONNgNVx3LZhttaXGJQmQ/lO3NluMwUKCAALcRIURPfWeLuFoRjLqcBwZXp6ZL6IF
7KzdBJH413ZVpfbYHXFi56siNF6AbiAT1jEcbqm6bKX1JyxwY2GsDcTTXRaO9lz5
S+VlznPbXsvhukkYe8iEeCUB9DP/ECBG5qP/dHgm3p/hjjdJ9BNKo4mLuwp/aeK4
hlIMOnBqFZG2727Zu7QxfiQbv50YX69kywmTDj/UCw7GH46P2fjHUHQzfRcPPGQ2
dFrxVOTILv1luNqPsXKWPPPA278IALxOjtczTLfymMZs5U3XD/WobfRrDOOiVxBl
/DvfoB2tp1pq5TzrLJlZtbo8XqbGXFeXB7p8Xphmq8LqrJmINfBMUXqXm6z4HnGl
2CWSbc7OS8jSZSNH3rWNKy8Iizrwhjl+BSV2hMhjiCym0UgrRvTj3SNe84/A7mmo
+d34jaaBYeimqSpZ5oDAp09ACVUAWxjjVnNt8ApOSRKcLZgLdmqmYP3YmCxJDIpe
nxuR3aGi2Mu1+awg9mgCZi4P+GhRMaA5qwvgj9lV1noYovYwZnWJIygoWspLNWgd
u3ZlVFu/h4vqz8EM94YNj3L24VHA7IKJ1ezYt4N0mYqAPAP6lJiogBfSEkDTHpMu
vAA5ji7EJ2uv20NuFBHFLKdT7ObMhVAsZu9DEPCNOvM4qCCe0D3OAzSczP30Avnx
wPfll8EA9HUD/vg0JGyVjkVnPHrrd6SNWdK3S7Jt0RTWz2nz18/28Aot9GNVbRkB
OCO2z6TXGJ7HJD0O/tqSjWEaAj29iJhUaHR9pEXN34fMUgQLCX9bVuULP9da3qWu
9xQv1PcnpH8ffzjpbTwX0os04xg+7bNQiIadr8bua6wjcy2YdRghzfzYlyvf/6aM
RAQgI8SW3jdEDtYMc/yXkJhHStzwpOEoRG6xpDTH+4tTomQlSc3mswhLnO3IuykB
C11q6RdAw4cocLubNJIkYWhyB7pEpOmGDF/N91NsmprO+E8f2yzf+DlUyELC4ZiA
myBHbKV7pXWlAnhcRYiXnQ8PXErF4dT0/MrQDoQX2IvlowrDLRCjvRkYM8cnLOqa
1dccX3OeW72nx45cqP/r6X5VQslZCT5g5aN6xbPTJhQfHCZmbgdOvCtsqaYB8bac
ByDL+Zl0cHU27N3XQmNlVZStKFtDEcuLEYkVd3kIM5jNUCtbcpN2JR/2tEeQgMwa
kG3W51CR8UTEalbvZUQWMpGlslvY8Uoq+NeIt0kErJ042Av00gZRmJGkTZcd8pts
W7e+OoeLJVJ9jYUL8KEgT4b6UocnUwgOMxRv0Iw8w0sHd4yicyWPCPWeCIdb++jy
7j356LuBNuYw546ClOeXEeE917rkEX+q/LVlwDENwEUdDWOPMSRycGSrKyDbBUsg
yOYNs/K0EALnJZEAIDOSLVC3Uk1h7x2mre5UJ81FHMXyVXcl6r9RHLOyJQ14Pdgy
VI2sq6quKFYPQZbnLTkvINdmUK9fysrBeSbGxXkKER2emSe1G6gPG3usRfcXIswi
1MCSdCS/c7dpwy4fwBNwF5gOETMe7D0apMuKV/ZN0Uyknlin3wg7uqu/VzXhpUNg
1REhNQ4EPxDosc66kjt4hWm0maMKGC2fh1KKRqXyioNZUK0GK3FrKlO7cgvfDOyw
jNGXGOpkOpbhfNSHjWqufHBzV2eOVMM+fji9ZJouLByL/Mcus5OUrtIX+CXgpkO5
WgSihqBUYYwmefJaJmxKbdvnGgaduLyhiqCy4aTpdaSz900Xcc7ZT0pIbONwaKMq
x7PQUqIjOHYmLfGc00xJShWz5f8mNZue7u7X0pxdWCGYbn7/sGV1SVaVcd0C7K9q
eLnwq/teikcmlmpiTNR92AaPWN8JKxW1bEvFWF+fLlYwOhBtih3DNFjLmNNJK1hD
YkKVcCSb3QGeDoG4czvM10If4vZyfarp8Q+j7fNdA+6CEJ2WeToPO79HTwPlFn2N
iqq8qknQuLUgFZ5HK5qsiXySxR3nmNnHYkQJgdLaaoLW/YO8CegeuuvaH8toRskU
aXv+Ne9Qzh9H/wuCO4nT7Qczk6etRMkl4QLetSJcO41CYC+9dLDAorawg2DlwYZ+
a69bQ0FsoGZs2kIr/5SSD/NSOGgf7hLBabgHr45TG3pWxBoZwh2y4yC6OgPRcaLV
n3A/Te8eQ5icbjp2GgjKTo8Fe4dETjMYd8E+d6vg+rgOCoArOmIau0a52seQ9dXH
QXAbvqek9oxCLrqSXKUyoAD+10JnXWyaqmZaF6WryaJifNwsXue8eIXkhuy4TzA0
PyZXMEa3ME2Tbf4xWdFsREPGBpWsdxx66fKwyQJMQbQmCKLEeuyryr+TbykMMVHQ
akadqe2wYRbO7n5kMNdrGkdaLovqBz9ue1cOVonZ2+gpBD/QbdpNoFIBerv70pWK
gt+rFSVAm1oARK0q9zAKUvXFyiESAJzQwZ8v06szyP5VfbfYZso7lTr6Yb836EUe
ftnKiKv6ZRYnvQyyNrmT9EuFS8rYNT+AGw1/KS1UOp+9/ZzDd7uiq+rhRRFf7Ai3
FCDuXwaonLWXSyZ0T9OxGgoQbk+y+YTJ4nBrYfQXVgAwH+WqwpZDGFSyrIuioDgA
asN1CtkWxE7JV8z2obYscLIZy6gp1z/zy1IWLYBR2iZ3XREkxUN76cy42zI8wgJE
A4RFTrELK4PY1fvwtI8Qa5zSZfShU8w1WwkBq26RzTyVv/OwjUp/7TOJvIFmJ4Wz
RAveJ1oDpukvx3ASw/bR0HqC5lyl255WkKdQrd6s4Yl8ssxvylnwThNGtu8tGWA3
SEFRIu/g6x1arfR4MA9s17OAZMGWN6EC55cAEN2IRGJ1jV/PR0CoAYR8LTM3rgH3
yf/JLy5SSgYgZYTQJQ5eAuc2Hp0KBSvX2GqgG7W18+OVm0TlcPEvodvYL8eaqhUU
9FRLu3FY5D9KYMK/N+TI7VpHoQjLw/S96eIyhev6Hwlbriedpu7hs1icoY5/zpcZ
YKI3TRZ4KchKOsEn8X1OeNQfpt9jIgliLAlmknjVTqZ7lE6tn9nZH3gKBxHFVyHV
3Mp/MVyaB4/D9NPoTvAfdfb+as3ZU6K3J3J6ijZgtPLCH7MAVD1WemkINkvilZr4
BbHE4SufdsJa8MkLha1I1gVlxV2cS8r6PDoCYPrVckgM5zRu/LQcgAPmIp574244
IEeIVnCv5uYXgCR6PpWkjuSXbsQ1oriMwebd/RAQWxrB8tuN3+vCloJxqx0q30B/
tGC6KUw1/UsOUHZuI9ZQEV4tLlB0w3AZt5m1dVsNbBk5tcflFr5vasJv/SqTI2uU
Fr82hcRdmkZVUQSoz+/hFjvMJLMWgWCD3d4Ghr5dMaHmU6/8mySgPmk0+APvb818
Xa/eGX9tFHusfZkUUlUS6+9Mww6Kwe7FZIpNgQOdEdUEslV3ISstJAQjxviPysk3
6B2TlTGbE3RTyQyCm881Uhu9nJ+S1mUprHZLZoDnx2WWWLMjU7K7nDyD5TL1dGEP
WnSMGLwu28Pq68ALu3socC/G/+epfIMEPixr57I7IzGv8zOHmwPNeirrwJNyVzsh
eSSjjO+npDuL8WCj1yv37lnV7RfAEogzl3CMDjZBcwETmi5el+wCYtr0baI8hcDd
gDeKwNcU7nkBNrXFpo2gxKJllB2Zl7j8EWmRQg9ZloU5oqeefehFU50a+oeQXXgW
dbwECQYOekh2eyTE8UdZcKglR53o1bejvxv5K86aYTEueSWxmvvXP4QU99vow5Yi
f4C0y/KH3mJMx4nv4Q23/py6KLjtu4np6c8q3g5n9nbd9+yPeToc8nSw00uKQdc9
/HFv6rJ+FVFDiLQ+US3X+foBkdcswUq5Wf82BD1rwWBnPxw4IRHIfUev0cwLabpk
j7pYZQM+p/dwm02yS7AkPMuHPiwQXxY3j4JlFuEJakLR6OIt8diOYrMGzemEY1ps
ajNSZCUFvo2zBvL4uPbQcDMvc3kHcS4wlWIG36Omu+emLZBZt4dGAKpgBauYVGwZ
ljQpsbp+LngGPvCA93PAQ4Ksef4ij+jnOBH42P1ul3cV9V2LPNOaPr3u1bBbBDJY
66dS22xKqCKJhph7+/8jyRxh0IRegdFp2Osq4PUrcA8RVcEF/mDBXmTVCvTOduxb
rZvUTnxj5ujekRsC2IvFM2LELXfWwaIAwnnw3r+KY0wI71hCPYz9l1R36RyE1MZB
wJeHQtW1Q/ltxppngkzMskCMq1+q0ujOS0zTXqDjT1gRcEjMQO3ROwN9Gz+xleQH
k70fZAfJfLJqS20lVFE7P7hp6QZSWLBi3iObgQskCd3Aa9g86NI3CSJzqW6FC9Vi
SM5EQl7d9n57J/lWLqSFxlm3cVw3E69wA4HPndm63xHzEGzJxBEYmSJYs75oxJ8T
tULSIKAk2jklU6i0Pr07RrbmbCXur+SuLr8SgRBLfU2Q4b3usNFkCVDdO1rKIXzs
Ot552ckVgWsZ9Sq1QJoHoUxLH5IYu42bLIUJS8T6U69/PqrXQpP+diMVyj0Jt/uO
NFRt7ln1GgqMAYk5oCbWYxgip4/EDl4anbtc//iSCH5w1t4PQ75zZAp92i0Syas2
W89gQlcdgvwtK5HR4DZPT69NTtPv964OBczAXVBLhYHJ2UfSpdHzHF5TKxfUJsgY
nbtglOKVbIvHMuHNw/XXPiSsmHCKWdwm6yfhkWLfWA2elCguDwEQHjBCe6JOzBnJ
SV33i8Edmg02xcIP0END0jDWbDKYaD/ypINN6RS9s5w85GShLAhevIDSVCsGyPtt
Sgd3M2vugH1xP+3rVaAtfo1RwYITOKhKg3xWs8pPaBtFHxu3mmSiKYU4V9+7DHZb
wFgruPACittGyhO90Rk9ks4DdaYHqgnDG5lWBMmkcnpkpdHh/071fuGShhXwgU+P
vYTtnNXNl4hrpOhqGfhSupZquBTVOkz50LY6b0NWDQFUddqKWAzUVcn/tdA/oKnJ
b4Lv5Ot//SXFp3npWlyuBwqi7PbIKfAmOgij/24A5TQ1GaApQ6Qi+1Me93SIABYe
BHq4IqgI+yvsnsciWeo1CyGsLZ/8WycwTguOfd1dZo5c8Q4x2BZoiyVoWawbki+W
rabDEdc3xsIMDSeTYtDdD5aKCjUl31GpfbX8zoR8wNtWMSUQibcDQ1r54hX7eIu9
XYi7vRiawhoG5xxPHHUIXt3PTZabBKdvRK7L8/v/LV+j5PQ6UJVUWPwJ36uF3HHp
bjfjeQ7N5AoSLzukRpADV1ytbl5u2q2jmqDoFvblu9UDbQQvxJ7bcCwvKrQT7H/c
X7L0/VweUWJV0iAQA+xHLzC6eLGFrLjAG1bs6K8af3Rka+BX2M3wd7UJP7Z5XScI
1AFbZY5b606ika97bh4dj//xI/otwINkhdPXvRiSguzyYeboP+kqh1iOqTSULZVo
MK7nkW8Yvdv+ItYaaknGLDN3d2+Y/fmGH8UYXdxXt8ZkbtM7Tztsj984Uk15MEPl
7sK/QvA8/a8nSGSm/9ALsDXsb2DgoqW07TAl+PQRoXiy8KCqiGSR+lghy9yH7DPj
QdV3dQ6CHVPd32B0Dhhiz0WlZtkLHGg8Sz1HKs21fQ91OlFg5bvZCCz8RkuMotyU
gFEdmarBoTPqQFx81tATtVFk8Rd/9fL/kL67jG2+6MR4Ku0J0Pg24PS1g/8Uf9PS
mEXMKzsFE76KKDxps8H+cH/VXOkOM81NwfdYFkPLOnDV2+Iy1XikkcZarqzD6uQD
oZ72u9GnnjQyyjUkYKZU8hM2RiETVPWmrYAbjLc4r7+cjDb4uWlDdNl8F8oxiWBc
BMX0byq6xUAEHyc9JuaL6DIxSQb6d/Jv1mGtStTP7INtxnUZXioteXAV/ELTCSAA
xuW2mUowk1I/hPHrLvA7cyKNvFcHyarZ9InquNe4B/mCXRTF7Qvmvs0/wG08o2jF
oZ7n9nqcZ8D9/j8cCfjJo/Gm/tAqExHNciIm9s1MVvUWGjpvOawNHH/FArA246s/
T/NT6+V2dxRyEM+U17pLOPi0fdl94DLn3L6MvOEmq9RZJV+Kx2Xxi5H7U+EdinJh
nmJN67FZTRtUuN7KNsxaMQuq2gFov81lbkO7oV4AcyzYI8fCN7ON7KyzYCRMmtIZ
q9kq3azIbDZgEFjB3Ge5QP4R3SNPbDi8jZp2Wl8pbWyG96koP+E3fTBhekBGJxP4
N0IdL9t6NMcZ8jvDG8GIJutEZ4J5x5QylkXR4YryJ4PlfuecyZQoMbxLH7xMFQvk
bIzhmvYkQktF8Nao19MURvTTFpyUGg2zZbn9nDPrveffkJey9cXw/L5lONA0Q+sa
mbCs6BkFd79MGnJnYYsKVtn/FK6kTe442+QgIxsrc2V4wFz3vHP5OJBbLO/P/0rK
d5RUYiLcodf9ciSrApG6Z0pigEZMARu8DBzfmfS3a2j4jBE16ec74V1SWy+WFyXV
HEYVZQZBcY1PFwNmF4siSgPNWzYxVc/XH35UEiMV6LMYQTdNOmTexEWbJI+UtXeq
K0qR9FJNaI+akW4rpwRL9lALt1fV3YAJhHKjV9yoNtpeVXbg4m9mHXETcmjdvAjo
3i1wpgz8nvkzbsVuDTPFSkrg7EsRXm3FnXi9ZIryFgFGkwEeqlSk6JdCVnQ4Rxd5
v7btEc2Vif3ml/9ZG7rFgNo2IvN9hS08Ig4r2nlj5n1iZV2WCUNHvlFKYen0uNO9
4AsnTwlebLmAM+9Banrfkw7S1/SafQJu02Bek+zY7HYyuMsczehA7fbbdeYHh3ZJ
mGTVpzUsQb9x9+viPzHjmU2jlVyPEojMZQ1xRK1lMj3vmsltw903CJQX9nSYb6J6
c25ZcwM4NwbFuQktynq0WcHCsu4tkRqj6QRUHD+H7I2N3slLoOy8UCJuKEFea7ys
6KkNsM5MPu9Cl1yXTv3e5SMoTmoc6uKFMcB+onmSu2d6oVrMLAvrRYj+WTfytfL0
jxroDMNHh0xRM8fDH2k3pwjrE0U3eOYoX2HQAfuKLwL4eLvVxrK+qGFPmYY+u75i
YmJ93i2O5HitLJq19f3TiPPDLiKTuivok77fY7ydamHWcUBvnZLJ0PEMUZTfdaei
NzWIpRaLjJLOC8BCPlLCe2QJ7DaSEn/1B6fFSye20LVkdBTP+Z31QHxDp5v7P+xQ
kBY66p4i2VwUclHjpWO3kfjLvD5cOPbhLLlKd1Rf+lZz7thBzx+D367fYrg5gv6B
k4SyzZIyz6uA1Z+Sh12OFugxNpC7MmQhESrxBHeUj43rBhZJC6lviTlybWF4J5Dz
a2Dw5/CkvBrtEHHMTsZnpXW9BoWnBFupx3gNg5Yvpe9GuCxIywaaP+VWW88Y0yKI
Rc63zTXKAFkWiPuU+9uaaSq0yRc4cba+fk8G8MgdQaN5TYdKGiis197Y7kp9e6kc
cqNMoZZNo3DLHvD6Fwdd3wsPwp1Fbto8GxZyL/xM5xdsB7Ttcc0bHWtoLOkJfFtd
OwvF7uQxzQ/OZIl+KXRX7Ux2QiKSNBTrPIqf2I6c4jRjy+QnUryJpfQHgXVmD5ko
DwuFPfZQzOj2ZofsHkcAeTsh/pzTkJzVo2AcBQLV+WhmtElIQow4F5vUNopbvy/c
WRpUJIVlo8KMvkKmZQvp2Q4XYmThgQgXRs7N6+Ko0h3nSM03txNp4fPbBDPisjzt
qEH0hW8jsWucnyDlyjnOtVacnSM63e+6g2/dsCzXAPE0MrzvkVHmjV98e1PToG7r
IXJqWwTx11Xh/G9YFuOvh/3if9ygDmriwVINa3poTJ06UmbVLVlkXES02tA3NUg+
KS6giSoUhtJOEaCoSs0UKMM991e9zmVSifY1pLtq9pQYHl84XergQp7IYD6pBoBW
hx2MFkPnHHE0J217KYMMAqrcJk7X6wG7bhBP674NrlfXpuIOti4wQZAFa2Qg1M4V
N1QUwuxwmEZu5/XhKYFhXApMQ5hUpkYXVoYr4UauD4a94Ijgg4lPm5DJBUDpPsvZ
SSxHabR2SROqNiJq+/xV80KSVeNDlunUScRFQCdQYjUXAbM29H/Wqp5EiRlffOuW
27fuxRlwb7PQkkgqzf28+km1Y6tivL6Mz+ty3gBlVRRdqXN2hpyUClyDKoxvZPBK
FT1I/4YN2wd9N2SGvm38AiYXNO6BFi1MxpsEsjMaxZoqQAPnj04REk9LLfNIa6On
2RSHoc8EUwKpjH69Rs8u3CVdNtfw6l1Op2w3gSKxu+OM07lzgIR/3ojl67qstlte
o5Zz9PJY0ufFGW/hYNHH7FZw8glt3oFBox+BhI9jj3zzI9SBlEsfr1Oz5PEDma8a
b+pZlEiGjKgGG1CqDmRki8sg0Ev8iM/rmyxpOoIeNCnmZF37xcITLKM1dzA/UwmY
e0nv5+eg9jHR90pOLobMQTzope8fkD/8uNBfU0QVV6WPcIZK/UAswpY5dh7ZILh9
wSbBk0b3g9g0pwnecoxdEHvNepc4T8ftnR2+haRGCIRxVeDnToMMif2HWmQNqyFk
0YEsHTZ71x3vO4pz35HMSnoXUeJsyRbXI5eNcX+722FhX0t8h7+mHBrOKEh9FH/E
uKOSGxVzukHQx0hdLEN6IHj0mLR9dViTnZwDOdQI//ky7jEoUtz4kcK0zgGM4vEk
2Xj/dVpz5CHmCMmR9uV3/Bd36lHJ5QoEPBNztAwpmsirkxO2Vkf3kWXOcTLfoIbZ
sVpjmzixaWoUax3sQGbj/dYy3bXUdTs/Slzr4/knERa33RYbL2MPgiE+CqOU1NOc
txJNjfkl4Qcke81DzDSgebMjnvnoVxX5QR2mNCbQOFhxL2uKFYzCwidadd8CV4cK
HUcfNuTEO5/c6mVxRSTCXjYmnHlMBlFSUBHnusF9X5qVAO7R+F/pTlSbTHLjjqDX
gtHowE/H2KlEU6LC0NiVjwjM3+pPoVFfpWgwmJ4lFxmG9n8mn3YlbpZiCkCzogKU
uF3UXCkguk5gAOL0X4EKMudRDLaIAt/dsHDZ6IOQdPnf5WGbX/QUlWjJ7q70luUC
Sm6/LJGFtONsD6rhgq9stldDNhcjLrEoHwnPOnZTxz7ShuDOTIkk4PP7pSFK3Z+t
aDnZRFjfRiUZEX1UOtJWbylWFjDS1GvsSUpkGzQ6cXoRMsZr3NbuquQBA6fAMs+C
T3pNAwwifm0C7woN32xXT5IyQKYZTL+KvWVNyQeNrwy4j983jrQd/DED5LRcDrLW
fqFAW+7AzXbMrpgkK7AMpe4B2IGe0vTwfZs9IGJLqjxZwHyuefHzmD2pwTopHwGT
kvg0Cl87dx/2C9X5osLMGKvV24Y15U9bGQQORDbRfxekRqH/PpSewULFUqmi6cMs
sJqvmIzStgkSzK1zLYG3OtjQlkhIZMfKQoBXbPtqOLCS89OkqfaadSsvowGKgVbj
FA1VfScZa0nKMwErI614STEBxGkc7SynqL9rkBTpBJlLO8SJ7T5f+QaZNLq0HUDe
Ir+zkwoYk717bo0AAkR/yiSqzm0XFJiwCtXB6LSQRRW+wSm4/aA13U5czCVBdoyr
78OjbYW1ecZMV/oIFblcE8+5Q+FFaTrf72QjSUgUz8+ckvoGgXhnHGad5e4sKJi7
A8d/H4PwHryIQetIj9qxuwOwKSKRwjqPgs6Sq4GAxMDmdpmiImmP/pEUeg/q2XHo
ijgDMEcmm8mLiEDpNTHO3MTCxahut+k7TBpAF67KDv6jarl4z7ifGfAiRsOzrd3D
TcriZSDp7gSoC2PuON4U54rL3Gg+F8vuLy8NNciyctBPqJQeguEjg49OBflisWeD
Xk4kbG1pQ1Itlsyef7xCRe3+jIqYUZ2CpseDOw/zYbLbLKO+o1aHxQFDVSZzfgBy
HCXwDzklGndHeh+qoS/scSHe2rWpXgi7K6TUQyo1eTc4UYsAmVQ1SXUFd2zAAZed
sh3HBtZiiUpgPvSPuoJHTEH4lGIPUmNqVDUB3z5b2d+8Sefl4z43M1WhNCJq4e96
NqCvbiaculuMF7wLqg6AHOsxMZ8Fb6ba7I29fOzWxJJ0+GDl+3Zzqmv7jxfD8Ju+
WYL6/7BaY/7HK9lAMIacGvUWMz2ZdRJJOkaBiTQT4/1CX798yqD+zAcEqPbeZKn/
kyq3au0qpwh7dvOO6rgOHMGByHzKmYJOfaXnS7auuiM2ycttjdRNkzujC/WgCEbu
+1N4x2IhzHRx9CFUv6dYn+zczMmDNZ1ChnDVdNFEcKJ7Fw9Q7ZWuc+5VsEua9xSv
yR40NVip9n4260HplTSs58iXHhNdCIOzwlZOMtKRBklpIFHxF7XlnbC+gfMYkP8T
u1D9kZhlsuFWUqJYYh+kWZbBo18iYOIS8K2/qKKJhDVNZZffAIx+ynuupT4KDlq4
E06A9jDtBLkIgIF2xi0Tpd6JO+k4Ujj8uNY9xbhzLp17suk4jceTdQcMDWdR53qJ
WwDZi83LnqnXUrIdMcIuqRxFQx4uVRTIdziluuNs60a95LGyylA1PzWn13ghtQfr
txKZ0tgnGTrRe1scgEiq3sbaHeIM/ZcPFx6pgtT0cSl7WlZ8YFvsBQ5H8geoGUlC
Ux1Yw81d3W/74tcDu+Qy3795JjfrigMCTwqXEfsEba85maVTAGsFlTnwmPIwChRP
B5Ur1SH6+LmcpE7AXSV4wRFyvhn6uailDasj+/3+CGv/i0L6ojPUfR6+pO3Lif0x
BJKb3BZmCzUeOGLpulWErJji1iJPUwedjNZcIT36LAo9zJQqJFSQttBb2qfKRh7F
2lidkjUqWixyz1WiVWSAzAX9w3n3gaKciamGRff6UgIjFc9RAKUOBMoX+aL7P5eC
g7ZxGavmV/ljfLIOOG3cKBnLhc2wx7N03xjsdz14YfJfU8YU8pAJ8yA/BoWY02BR
o5NxCU48BIEqNkCr3GYId69esqK8iHEqDl164Cq903vQjShhZjfHh7pxFABJE+k7
f7kuZdVXyXSkzQ6JHO0BJZXGAHixdOu6rpmlOwydlth/aLcjVYk9ftalgRyB8Uwo
n16FZehS7Qz33hrKXPXtVca1tczm+/4qbt4mTX3LgrK4DYtSn+wPtKT4hXsbgG+L
rfcD4hVHZQJn2OISl96WyVvP/NQ6R5ffc1KPm0b6yju3wRxv3KxjRVcBxmASOWwI
MeVi0L6V2cenF0TVfhtcnyqMaFxRgwbRDv7KhTvP+gCmOkRatNoxX3b3BcykF+0V
PvYGsrmEi8V+Rx9n1ev9vp50sOQ9UpplhdayIUQ3t8jp5H2HvhIG5iB3rd1QjQn2
XLvxaSLM8ZB/3yraHCsb05cWXQxzsWwfJCeVeb6VfF3Q0L0FNdyejx2njDPD9laY
pGJUmq1P0HHpVipdNktVN7X5Nsqzthx9EKSJ8YoQv01R6T0m1oRthGw7aSymUcED
D1lndRiHyn4vEvg7Wi7L2n8HgnR+g3pbDYLXcHONHFvivCxfvNXm05n6/n2EYI5o
lvlPJFPZm6iF+2mnME+Z2SreWI+ulx+vp13ZPIw6povDLYoB8+nrd2hvSzR617PM
Mx39q6RaEyxK7GSZ9q1cssZg3iWcEPwd5LhajbD06LddoWBGF/iiglyIYgPTYSM7
HKlyj2LPaWb1E3yA7/cZrgrRsmxzC4UG1gD7Pts/LPH/Ss4EuLSvaZhjPmuMp0PR
x5YssJoWPyC1/FxHCX3f8M4GJ4XFm01BjghPeId1KlQTGtv3VXQPchaCuaR0AL7w
7zRGgFhYNguDRRFQe6uwEPUl/Suco4QDveTlWoYkKiO6+Hb0ajgIMLocUrLNKO0c
9YJeX3sROy66uJaN1fOtkkMzAYzn1ot4OmcDINOzubA92wBLKI54srD6fxZGh3tv
wA7ReO+E6H6lIpf+gYmNiuJS1VIwnQxuy9+F8OkP5SfoS38JmFhT0bbMgYlJQ2yN
EfXXeuu01Dk63vWSZi7fnqlKOkj0675dt0RzExreEYpEx9/qTgzRejiLFmqsi3n5
5WVankE6Sl9UbCKQqiW2F70vIlMK+DR+QhrolBqblxlWqhBoY7pdhPOgMg4hI7Un
B92vUX+2KeAXSFkpi/BqChEfbrNj1+2Ydf3zc8d/yVDgoaWr0mOr4Dkujt4T6wrv
O78O20CY1YR3MCfTKev3u23d2GZBTWGiuenqe5cz3pnF6CCfgN73ysA9tzOCqtbv
LcVSM4umhX5H3Gas/TPl5jq9D7B+/zH+oYKCwrVSsNk6ipO8Bsx/MzWRP1kCAU+p
Ct8R2uwoRi56PRXkUcMQSE2MkrFv1CcFlncoJkZ0WAAygPvIZmgr7ZBFXhATseye
BeQHwAvTaxudgGkOExjulpMakY6PRQqEcBFzt/pB3yR7Rab6iqHDgNqo2aOqi8BT
BTE6Hl1Ns3nwuZ+CcQYTX0mkSA+ez/p9bd1Cox0yDkw0B/3DRp0dNgjjeQcUcANS
KlFIc0VXmRX5Sn+kkNBKttEvMD+fQZU7kb+f74bCDf8pBgbLfjp2bcSPbOF7KZeI
wvOSji2YpiY78MiwndZlNBu/BWTj6JzRIzsgXLbyKEULxHr8JxSKXWIeMuMLKmbG
Wp5RsHYtIa74nCcCqLts4FQuXfP9xT5FzPg8YRSMEYX+ig3snbsDjh+DmU732PDO
RdiN2w7QZgBCI7273ycMlLlSaGTcJg7LAb6qnWCHesFaPFkEGdDR9XivVDdZV4EJ
saQfegvav4lzmLrWdtpvik91NgUk9teyBaK+aOqSv8AlABYpWXpSTCziYDYKRuyS
qnHHi1yDBp6e9II/C3tHmtxf6QrRoAJhwRiTqEjUc1whOuPyj4L/7mjunLypJtcq
Ufcf5fLil0zWbEgg2NnwIpW4e5sYzzlZHlhTv6+D6V5d9hwOfFBYFtnb4G1OVlgG
2wSDS8SIt8rdZYZziDc0vikHkTWhXNyGHva+9qE5t4CwYhuVmEWMMNTsK3zvxI4z
hCkXkDRv6mUSP+8dSHx0HFgK9iGFJwevO8PYD03lByzSaVMLjNsOGR2MEFpJTaIk
aZlr9xcA6bps9ykikTF0zzzyuhozrPfzIyjBj8adIxzW4wCf0oWp09VZfTDImPcV
Z3yEi+DK8B0tqBgvq3X/iv82Hd3c/4va4k/YUrOceQh7nLhwerXTRG/oveCwEz2L
bvg0/olQ7t24vEW17kcOKNZvqL4/RSNXpBYv2Z7/csZPcgHDXl4p1jU1Uu2YBZ9Z
YH0ioerar1TcVQI8VhsdVvC8QLKECw944ZsIkPay+WrwOp0ypKxip76kEuh2oj3M
ELrMj2PdHdM4PxcOxBmbarg+4u5isqE2et50ahV79to6GERZBOIMZaFWLmPkB4+y
68vLpTav/bgK9iU2/qe4fxcHCGk0d7DtWar2/gnXu9lkii1tYEtuRVY6xAL5o7RX
+0ZfDPxH7Mmtsng3CdK5MhmWNYk056ICKfJ9CRxp931rpHzaqVexD4vS9iLtyrvu
iYE/MColnsVPvxaV+SWbaIOSS9bYBSI7mQmROi/HhZg+Na/+CqdidblOveMYhlmS
0z9GOed0oXf21KNsNsNdmMYmOk+u3aZ3Ihzm/RHO1wQNpKrvbGQk4gfb/fr9wbIs
tXu9ttuuYsxN8b9nHQCBHGlY0TxbU5GaMwAeDpHBXojryLp+QLuWbN5BkgXQjoYo
pS0RB0NlgiOlwoKiAvEBsQB3K60JBVJE27B9dTcc3iwrMjmRkjytvhYg/0wFU/Ow
jdR28e1bbfe7OqnoCu3g7DeueGUEn2D2G1tQw+FvXSldwvmyQk+3HdXYD5YI1GTQ
KtirUdrYS3WoEo+6/PaUrOmqhOVI0cft0DnJJJoV1Mf2CcFjffXd68LZEaCXHwTq
XrGSXyk3rZRzRUcuZ+fmgpFMax/d+AoQ/I6wi/dyHEkV/YJ+abwA4U4E7kSuWgr9
1gu1W8vNwnw9vn8pNYjHrqO+iojLWyp/PNSYdcRwEsok+sV2p1ircRzl+fk0+aR0
9PnKitLNCPfM3L9yMQNXvSy96RC5aE7y6f194MCMTScGT4ohrykrtVyUN/xbdIak
aRuFjSQRmtN58msXNiak15+9mLVfSqjKbWlL8ifD33+eOPb4h1KRWc/4YM9uwPyp
/IB4blNP1yhVb7fQbKBjhVk7XxQ1K7sObrIqHtBfARErRylByGvUtZi3eMkuUgOo
gFU1eXmQ36EjPvkcX/bcJKHv7W5JubBk3YpRRUvwQjbN6AOVHqsxSEdRVN+tb0YF
lvFVhOhKYg7pFSXfc0xJq0/tGD3Y0YoOjGXYhPihqUXgkuUxzhQAAkCEtnvmxkCx
Erk0BDX2l+Zw5ii6MTT4vlodARgU8n6fmUyfPpsife8IZ4ReL1lGRCBS+AvIlEY7
aiRjj9pFju3jtnn2peO1B9bcfhYDkM99dHLCB5wFyx2XZE435Bqjl/3AN1G5vip5
7+uMbg/jQxuLBNzS79iU5g0pykFtymKh9eRsWFA30Q21FuV4YkD9e0ffnS9PRMWZ
eG0P6uaymLt7LL9D8kfGOvhZWI+uS5XYmA/fl6O6NG8ymKT45ejmkrwdBvZJAMzd
VcMAyDnSTC4FqkdlpUjraHIH+sBnAJFv6+X9nQFTx97Dx4/s0MklYVRODFIAVkry
xMIOC1hN4DX4NRnA3HnfW5ipk6I/oE3JIp251zDJv5lpGllf96+9eYn2J5PLFkrg
yLSj8jU+2WlYGCeUuDprlj3U7ASjl5YqdE+9dXOsonXCjBdSBtK5504XqJ/ARX8N
hgb1FXNdjwUhOrsR+eYn6xI2s9knhX2pyA5+7yez/WEhasw/jc0/sDLsr/D9SqSi
z7KQHrn6zy2D/sOl4/NYOJ+Zwen8hb1GBPugevkRpBllOyFkCfmcQkp9DQG8hy6Z
4/F73gkU+MBylegg3gp6MvUe3M4Bi+wXVXoIKvn7uWhFM2Jn4VO1waGKXDlrehqo
PM8VAWnB6WN+YKdkLpJ2cxLYNH+JimShZNnXgRBlR5/GiiLOrSJh9xhpEtzMCcAF
4EHmkurI8lqGVGyGSoomNLoj944/pa4SGyn8fyQyursTdTdzrUjzZQK8L2KKC3+k
IrQmUx6kxpJvcIuzEzw7aFG7y3d2yznSOmae6LrF6BLHAdiB5hI5LfyS7Q6kx0Hw
T2BtoS9wETsmK8FmorZJ5UmFgiWg7aHU2UX6zsM0B8xd9nTW0qrkOZtZJ4aWcIfn
x969taRyTavoBf9S9UQS4I0hcG1WC/76absPHLzNtF98qndhvphhub6nKmyRqAkB
UtNeHPGms1M/sNCVDRmIkdygj265JCmLS7k8iNjleRfwNWWJ6nDoZ7f1G9SJLDrc
aSdDcPeSDE2WXDXfzG1o9JSQLUqZi661aECdi7ff/GuSw72a0p8Mm2+EnzPSGRpp
wtR+Tyza2lZzdvJdfA8ZvKQ244JjtRaDU8nay5oimGIM3OPoFbJLy+IMtEt77LPD
CZlzPdqua500lcviXcZM+9yOdppxnzTYkwlUHYD+aBPt8pn9hsGod+HhxoBoJSs+
hWAnB982oGFGUmzSRSusr97Lx2Au+A3PuDic2wdPWmjzXZpRiiAvAPztngN7G4Mw
k6BVXthYHPTIqPLpfp4/Z/iBWtFJHgIQ+26K484B8cGejBx5bb5X6UP/kNvKPY4z
NlrjP4b1Pzy4TY9ySw03icQ101yA5lLkduiyoPvvty4+wOMnRK0H7wMM+wS6zQJR
XO7zUYhB9eK9e5XFwn2MzoAngiSatGFndhN/uc4yViVMJb0MaxYm0NCikFK/+4hZ
b74ytinUcYku9v+Hjlvi4yVtyWXOGF8v+gJpu9Blf8vDqAQJUEJTbyk66BzB1cLh
gQ4EKTKNNc+y5v60yWdi1T5Ivl2bUTdyj18EsROmva4qdwPfReetBLyo+9QqYSPO
s29PA3ZEH5nmnax0oq9cZzMXUT4OclFvixpq16zhwapCvFrDgVrOXm6/KNpW2+s6
EoXY05o4p9ZMjd/EJ/KAEDs+Re+f8CcimeXPr5Tww89N1w+89z+ENgdEJ6rH/iIn
1O9BpWQ2fqlGGDe2MC6GHQ0SiqT6sWJvXO3uc4azXag+h1zfEnxyN5gHegi/+vJJ
u+x/z1mBd4Xy1SombbVeElQBi5l29s9L1PJTCFdzTyaNbvhcdV9ZiHQDBVhG+Q5B
V9+MZ85g+1UCB7tJdvIKkEF52WYl1FSgGO9Tl4IpHwrYheCp5AWhvfdzV2+toDJc
IG/T4cJOsnmYH59KpjNTwjLVgzvkeccokg+8/TlZLAYq7hT+6rTXZ2s4EIoaZMTw
hHsZdi/p92cHwvIxTnKsaKjQVUEny/SJaa8752XQj8ktshBH3Zk/QL/NiKAi70s+
3Hi9RYEbNdrIvnwtgVlzYZjBwxh233zdX2MOJZVU9xP0Ln/ofuXy1geJbI11lZYi
Q3JKRshhc8sjN9+Z2QljWcXp4XJvwuSeGtYRx3tnvB80910X/n3dCu+PNQR2b46x
HgVGr4tp69S0jAWpVU+SQgh1FDiUZ9Aax07H6Q7jUIVUoR5KY6i7tQRos7Hvko4I
xkAB4isMQCaQ7lCAtl8AjYspxtZxIQpJRIX67/ezvziNOxzvioYyaJQh+th8qxoP
/nagoBJiNmttwCv6DxoVaCcS/LYAvyqWp/pOyjVl6pn+7nYCq8csr2+5dnFwqqrb
74iO2JlwcrTj81dYLH5Y8xXO8/8QsDCy7vo0kDi2Ots/vM31wedMMYWteKLv9bL6
yx5jET/ED8xewasZvkyB+YsfpKbni23TTeWUmXZD2DqI0ztqJQ6qShazaGfgZZS7
NNo5/XgMjnW88+apf5u5NZbpD5nV3eoCk7o4oqep6wh7b+04IDI9+xDWOfBYhTDl
wwnNvAxv7eZer46NO+PjAfAMZnpKCiXrOh8wVjFljIdB5jvL9eYBYAHSGswxagDW
2dGQQbXxbYlKEo1y1GW88hBHs2F/qZhPjo6nRHi497XFj3NLJ5SK9IB6DdBowqiY
Wa3MKane3Bvq1JI5Zz0cfPSL3sQqzv3/7K9GJNQeNxQZXz8oBOkCHQJuTnp89fM2
HrDuiQ6/LJKtqvdGYI31KgBeNNXYuhEGRwP//euHQiELnLatVinzdYxXmOQ2gqmv
Tnz7J7mYtLdR7tFI7LnLEXgZX9YduB6/X+kiz+m2ej2MD2I1yxIAEtAjmf+k39uM
SGTjfdRWMnQhVVK01AYk8n0JDjJGovf9/4gWiCZsvyIBZSV6ik5BAnKdzwAbscBK
kQlf0tLcwZ9P/LvY9Fmx07bFHJT1zR0qOpdoVQK/lWfjxF7XwAHbht+wEb9xlVFq
sjg0yo7y3XINcOSii2MwlkO4e5okTPJrCqkG1YD3QKuu53ZBUme5YvwN9GWbbPz9
wbWm1fHmSbfrecK5JH5PJ+p8vVs70xl1jaNq23j0XtM1UhvNEKYzQSsm8XGKJ740
0NOPPZ2wRQCrbc/2n6Vk5LLWpkvzxVs/ZQx8ZeM01HO4EdM+T+3XrUPIOODeXtif
eVZND6bCZDFUTx6Bj+OtopYyTiSbZOGixX88dqtLu3Q63ix7dnfbEnC9NkRnANKs
pbAILGDwvnpqrmw5D8QxMk1vXnwUSSzWFqge1McWeYAXcFr45LBFzNa8rFwiZlfm
seQ2chwKWsdyNZ/wFp4+Kw6kwQUS1eNN7IDNLq7/gVk0PW0FBpkY4wRbNYOFJLTz
bj2XYEmRHpd7jrOg9WYewHRwxx0jFVx9yiLPf1OmcFulzo++5xxtzG8EkpPZOg8L
5h7PMy7KyDSrAWFUO2bw1AGIBDYq1Beb64LqA7/rkC6RrEFybqicGdHxZmDgV8Vr
21Y7WQZli/A/yF2hI4NiPnvHgJxbHobOmdp8TRnBJ+t2Z/V9EmeEY2WZuCPNXHg9
LWv+BnqMmiHZKxZTVSNawBApEpjq9AxhV1Pwqy+NvvYpQrUUvkLsGAL1D202iPE3
Y2uiJMVpTDkMSzWWJXI04EkQFzsd8HXnCsCz6iIrjvIvZusY3xlMKhQWP3zUPplX
OLzb+byuKUC3QuWGBT+TlAZ+Hy/AodLEHSpC7sYkDsd7PKjNCdde0Ez17VSMBKu5
HNW45qShp/rbT472hQGLZR0s21W5ylbYsbfPffO+Ccy3eKbxjft1Yi2feVNcWGBM
vZvead05uTSsqY0jk1l6lnQdE5+eDxbI5rSoMVRfCVdF9tPKEICAxhW97YC/TUjF
TMH7ZKJiuO3oYeU2k+Bq24epy4ASy8I1DcoqY6G8JMaHY6QZa+Nk5KiO6BI9ej1L
LtbKpEKZFXjhBTyyyEbqrtc6i2O/f6JKubpVXsQJMQkOsZVKsNHr6dXrY0MsDcta
Nx3i5xH6p0XCBUwcSMmAlpjizuCP+cKxrgmbLcJcpD0NjXy4YolNeKKvh0Zg8E74
Dn8DQkqNJAHwN8YSG8l84WJOsKxRcSubrzbPrbbWFMHmUBAacJM5UM3LE/ze0BEe
UNMhzOtm5jVtfgVHH/chjGLBixSRzNaUQH7rGDyHcFD/H3p5kF0TgK+X/K9z3/Q0
Z4yigpj0B3DGv0bb9HxH4iYFwl1f6Nsedns6WceNTmnSYhfrEOt44utpBiIl3e5T
k91QJ280Mqpp82PD549hOJChKqellbwr3Q4iBgqn35rseNjkEEXMykimMdZuxxJ/
/si+6A/Qn/tQqchiH8gHvCKAdfVVXJUV1wp3lYNrZ3LVpRip5IEiUV0LYCtGJrMC
j7N1OLMIv38KCkubkMgepoeYwRhSzEaMrFEY8PvmuNs9kJnOflBZFubFutMAhu1n
X1Mx8AE5zXY95I984mHhBuOgR19WQWpBYMb+ewAu/soI0NwgMObmtwvf3RM5OoJx
Lth/ERHIyhhT3l0Z15PwoBuOoyytuxrjWKqsBF5NDgCY2A2R1hI5sNo91j7X786p
nwI2iKH5aAewQajoMCvNZ+aWV+9HxHlF+d3IyzqpsX5OpEfWZT39WiDWYCpP4PwE
GiQOGRrSsN6KlpsBEwRA4s3ANw0WBr+B9drkIbNiV4WbXWZVPccfNH8aMm6F8Ofm
S9nma5xCYfUSOM9JEIsrtxOQzY7P+sIqfhf2lT9qUg5rtXxyxRcQozbHfH8JXJg0
jpw/zIP6cnsU/km8W69vE5sEQra+y3ip9XhGkwoFPj3C99pugefDg6gFuppnFuOx
bVNScJN3ezWn8VNwG5KJtEiIw4yTAKmt9XGWEurgWIj74ogyNE/b40tdcuqQsW9k
XFKA7YQCW2aRuO6pkjWoJN7Dpe9ELNmzPMA7BA+BEvA36x1qwd4pIi35cc/2+toQ
K7oEwY0hr8c8EFdA3DRrPpyByHFu//Cdz3zsvy1EtipxStvBQGCu+t4f0Asl0VVI
SzCu9OuhIiCsSybojbM13znK/f7giN3jTXfRgj/2CrPHXn8IqWy1o8ui+BRd0+vU
zx39bETTMud7UU7ZkizCulOJMBryU+0OiFXvgV119ZGm52Dc8LvPjb0aItaZq1yb
+7Y6nkNDWK5PBs2/P6tfXJYK1cM1siUAietHhkAaqLj+jFbanJlNV7R/bd6DWCDk
YYasRe/JcohilXJnzJ++VJPpNQYhhewD0rf2lO88LawS2YrAJeCQLnzmpqXDsMJF
sKFGpTglZOGIVivIZbL2JFLUHZLTLTFYCpuISsZpH7pjZFmmJxgJEFkXCQpZjc8c
xJQ1Q5MVbOHwmPK2NLWr/2Q5y4ta+ULfxrifCDOkTydhV7iJnTQy8k5J+YTa5hsE
2jILVQQ5a8MFPeulhY8352k8loUQ0Up9VmnQKi9Os5giw5PP/ZYx7mLESdDtXi7k
axXs/+cbzYfp7PjrexnA/vncx4Oc0VOgxz2XcFkcqYG6YEWuK40xEaJg6cbhuPdd
OvDioX/zXsvceUrJR2AtY5FC4NMLH964lQ3ftvNBZtbFowyVjwr1YXPFo1e+0tu+
oPt/VMEDd1dKf47pCVUQECfrp2x4a3kk6jaYhJjCACVLwV/TjSho8+BUR9t76lIt
wdjVO1CJkEFDbnZ/XFMaXMF0de7XvhwYXHaV+UdzxSHqa9vzuoVPuxLXmU7b+i6O
yvHRmB/P2E2pZwgQgSFfVe8Q/sDV+w3Ms1ky1sNXANBiXLO4NZZSmukcWfJJDDOB
+XyB/ycn0pvF8QjfBHUJQePfSnxsrGE+1Eo2jNgqBo+BW+7y7SONMTODohqSaUWk
7R3VxXLPbtuIMOwdA5aW9PDzdNCO+KmpgSL6m7orN36UFJzWr+zz9f2UzAg70NDQ
l3vKDmZ1pO1jLmD1JO0ax8OVT28S4+iMOdTwXdxKQKObvnFIYOvYhNk0H0ZyLO8z
sS5ysQ2mHEb5h7j+3cwZdWwSbDpla8vI24XadPt2kpf0HOYqSUJgzpZbsz+Emv7N
RZJ032iCnBZbbZqQrnemr+RelUWf4Ig4oPprDdm7KBYhbnLlUiWNoiuZpZEGXhmj
9FbyjMjNEyUyWMXPdQ4wAxmOtD5Re1wezHN4WUs+zLtvOxiSVTatEU4dpOPTDVZi
jPTDWIZ7o7/4Ux5bHLjq3ajpHdfQ5fF9j2NgBYGI9BL1WqeoJKpEV5H7fNIjUeDN
Up+6YE3nbDjB2u82fwjmdtn0EDTGlshETtxWXVshQxqkHRq84rRXP5WGCFfx1IIk
QiZTQkKjYMExU3GQifH9zpo3C0Y6RcIB313vHWObGbUf+lnz0Yk+v556b3Nbhtjk
VyJmTS6As9ycGr0cJbJCm56xAxnkkECSHf4GuY7gdp2MbiYHHOHWTQcqTesB2r6+
2kKaQU9ws84DUNHXax17zUD/DU/E1A/Ymj6727R4RxsCGGbvtYI/tJf4krPhAfCK
JP/LZNkTLrv4d04Ovjs5NfEygvjR+CrvJjd8dMaw81dMUv6RMld1UGlZ7GIMlVO8
v69s75YAesdxi0GKk8zXD/8NJUk9+g4bccuIuwjPXKEO9rQ7Id7ngNjTMhaXyi/2
WHiBTecmApSWKDWTy5uWL7BYy9cckAMY+jVhsWgc9uReZACDIlkBZfJX+l2BsxNl
LdDifcL7WCnQAI1kvzCYD7ISqSHgR8+khbPvnO2nNK2rLH1SD1889raKXDHUmRUb
j1N+P3BaWiEZF1ptzY7Mmv1am5O5CI8MY6SAIQG91sEHPLZrc3L8p4vNuZFyj8XS
l6nGZxf02++/qzTj/PcQlhbl/zo/fa0ajUwnWDE4e2xBybxvBqqfnKndcyD3sKdS
pp5Ua7TFFbx5+iA7BDVnnJ+BWrU9xSH+XGFBhkUnz+WXaCjvgX3bAIrg9I0J3lCs
8g1NeuQHD7P4QR1cQbYAOvHm9kIDBQ+jfjADqK81+N+cf/7kj7zatFnbiVwRJ3Me
xcFg/B+DcrloMmTuPhfrzH/kyN2+5x5Xl7Uf/xlanazI+c8JmxSdQBGStHE2QlfR
NnZ3704QJmNLbkHzSrwyx2qSR714ePs0Q8147d9nl5N0g4C5eL5p7hDnT9l7TLyI
O92nwDZDqXBVU5Rax3UEDs3J4RSplhh6ypRH6gwYwna4opn0twzGgESK9vZIpc5O
5/xiBXUE5y73c+qBHNchK/KxgffaQXAbiAHUwNP9HRvho1lX8sL5PTecmRadrOpY
b06rWR7hnYBam7T9tTMH+yp4BXYx+uyYnqNfMsoMx6mvZ0cWS7LlpBBd9zbTmU6w
vohn0bljksw2i9eNnah9ZY1sQjao0GLU93Wq/4CnuwEm8pt1Q6iE7lNtlyW2a5au
m45Nx62YAtPk0Ux+GCtl19BlI10r2Jk0gIxLNulbMGOu+sWsXH13SjFB+2VQV8sz
G3Kmf9ijInSa2argrDaw8z4ahVgnk9W+vTnjG/syeJjkx5JaPwwJPM3D/3JCt3gQ
kLtXqiUtLc6I/IkKHMKkA7jijAbDTdDkry/1uTsM5VLXkm7c3WEBZ1AOYbDnoFoS
UpOENxFgp0jyCYEVJkdIl9B1wLrb+ksK7gInNxVSkqQFwcfooJmzTuDK2SBFUhGP
fTdMMGaXwYpP/dHGhBJyyTfcrd6nm97tRjJW/44xvv8H0nvc562S7C6LFfgcMyJm
qg0hxmcV3sU/RRDmcpomeQMxbBMKITPLXAlvdEAEdy0yL++CHyZBlvsBR3KXOpi0
72IQosDN18L3Byl8JMf8up6kUjXrcWtd/WNlUI9irb90Wmdtb0kG4rz2igYXflkK
mXPy0RhTFSny6ibW3HD8BQ+uuPe+O4f3YymyoBhjrpbb8xfk5OpiOMWa1EGq1EVp
o51HktQ3MRDFMAbLz8oUl60GPbDSYX+SnQu03kcFY1QE7bi3vZ0AHue4umWvYy6d
6hEW9OSTSFPFDzsJlaMakvp9eUFMST2UEQCVgYP6HWr05uae9tl3gOKG46T/iQyq
xpkp1r5AMGQ6dRo/WgmSYSV10ioi/osdxTEPEZb8rOl3445afcbJxA/EMQ8J+mva
tNaeR/lRsuNSItttnCqFoYhhRwhd2HNASUsK+m8mDyGiSaa0qlUiuubtmO5KX+vX
JIoE9sW1XrCoYc7teubXTspB/nerkbSQ8GpRB7mdPsEBx2uJfmERLDJfx0def0xq
FnbcwLETv+5o6pnTfKqoMQWHmNcVnlK1asMIeMFRMQ3xbHTcLsmX2ZVuPm6LYBSH
g+PXhtHI58Cr5btRvrRmWMuedTmZAbTSPnuQIyqQlaqOpc7kwNuElRZX5YXd8Wdd
LudcQganKeyt0STG6UmoaWxtYTfIBS8/py1pjWu2pxV4qwiNaHiZEATfLNWxZta6
hYWKl8fFavex3jIuKOPeS9aCkeSgg/R/dqS4BUkricWUSQ3cpVYH05JW25+WhxCF
AvcbXzUPn/ngqPwr3QXWw3/gO3R4G85wlhw0r8H/f6xmEOJASIm1+bphyXVz3qEK
prT/sX1eUe1ltoiIWgYrh0fssBQPzmmrA0e+t7+zrszyhaQoCI4rRsSYj4N+jtnY
Ij7z1zDgG/g70yzpi71jx+mSvaWMmXfmoeE1KYGtP0dzt5iN0Jl9wB/7Tgxvzypf
DIyXQAw2c/+kSVN7/51Eev0ImQN+o7y6pwN8juXdzip4T2x8vIyAPTZ5H0HYbQ84
QGSMsQjKJSmSeQY7bObN9pmaDKM7edFBFPKB4dYIRBovoiJRzxRjWb77VJHQi+t4
ZUmaNxp9mNGM5gv6bdomYduZWQufOLs+Vvwd6ozPZT+F8fublZSPU4RSL/2/eGCt
NrW0yQOdnzHrQe6SlMQo2WL7jNW/Kl3Aj3UDGEzqCqZElG4kZIJp8LCev9459u2c
gH8nPA0Jf0I4Hv6OpYP11xS6mU0ZsP78iqagXRgzz1gM8yi16CfhhCdqHhq6INDf
lbu7jFeu7xRznAUFxHMMCWmGF3h3h/DmQgq4As3EmmqVSMcCtQ+VRNaAgvVz1bEd
IuUUP7TWYJyeUBJQyE7GaFs/joKaIZDmrltWX1CoqK1Q5XiPHupO9/XN/n/DNL+H
RYaTjOe3NQqRYAmP1KXXdnCQY0dupkH2UuY5oiJR6R/R09QHFoqtlaD9zT3cKl9w
7VW25sc0OlsGPkl48Q533d7z20dbH+m8ZSpatNwRK3LiIf7M/Wd7RZcSwZJvZkvh
d7vmQDowfxgwAuCD4HMful3T2dHr7WpUmLxMRobqltj9YNqtkymOhfSIDcPoUTlI
B0CXW0FzAlWoqJiBF5HEDjyvfn6dAmWkkWr3NWV/BpNb6VzutOwJ/yEuAj/U5QOa
Xq+OEsJU8NzlqJpxiMjDJDlUNaSvNZtjgdg31EEObKEJ2trI0qgpt4dcYEptLWNU
9K+AoWDQRSHChhBiUWYGebLxZJV+1qhGistmRpzn8UDa4uIX/GXNjCKz3+u1e1vv
fEcdW3kktAx5ovEsZ+ViL/tOeVMgljelR8i2GNzVD5MN/qKtTrTMPy0g3NIrbxCb
6EZYWuFmNFAexvdUhE/BKRzhx/3O3yW8R/vzEjFrlaG0EBQEXludPRbI9wAAgPzv
nddMa/9S+vH8G7JTVe2NWEEZVAwi1PE8MMuPUfPXUM44PDKwQsQET5imuu7UrUea
LKGtIVVqbEir9qsZeKAPNYTUVbxLRZ9ohuxxW5GLG2c+vNx1L5WrWbGPgtHa1IEh
egYrrblMbm0CL4FO0wF7/KsbIomOo7W+1sCdko49giS+5kiSJUmzV7hfG4xxg51b
AQqAw4IytBL5+BpuqANZK4TJ/DNTZXdBsFg+0WM17oAhhu+ca4wqv6g4PrKpBSYK
qJbwGPR+szO6K+pOB29vwwub6eqSvZl3Cl1oYLxW68UNODm0o/07RbvMSQxpsYaf
sRpoKIo33WUBaV6sf83b5fiwWg31luV+d8K02F+4kTXlJbUfb/l/0JDCBPBTCD95
ZHgoFacjFmOgBPlDrPtpCyyQA7vTOgy8UezSTi8cbhqev7Nz+3ZV68Spbi5mAQa6
aoz8aTYId3H7HgJ8FoYA30+OXtNG4f48g/rW8EDvsl83pY59oKKk6EJyB3kxweE4
5EKl06hTtfa8Au2vhA+uhlGvhonvQ848kj34bcQKBeGYz2qVrg0YRNUyRUaSjLCo
hKDs628n3kagXMGf0KqaD+QZcFvZAvFNluqE59hMse51xEL8qr94r8w1hB1JBqqd
bewtAiDXxbeZzwqbc/nXvZDif9sCLFD7eKjG3rPg47bG3N2JQ8GdQ6CFAhd7Twr+
9zL8ORtABCfPY3SlyQoniaA3Rtp50v3GFQIWOa19SydBjLeQvbJt3bh/jtEWLKfa
jgfSfzDd5dWoT6FHKHdq9hZ+/kNxcCPUBUpdfkJSB9ZI2HoTryJOmyLAUD9xM4wI
8P65TWRY3ScqXqYl4MenE4J7B2XNbEnpwaqWlvA2ubKnb2md+jmDKEyq5phM3aVu
t7XIsEMe+24gkLwg2EcmOorxSiLDXtOJlZHUWk87MgCnIP+KCiYpynfFVuEL0XNZ
wzwSPdKl/KnbQU3xv285UUizFJ9U778VtPP+8TQd9zO9FMg6phar7y4oF18LJl2t
bnihsLVVwSBbiAC7JbosQaVwpG+N/KBANYU91pSdQPBjPjFhAlPbnGHC/0ttPGGP
qmbtgfnAN0qrv+5fTT1VaQhzMUSrtSzyR392G2BEYZL5QEYq8GniEAwudnvELvHV
/aBl/sORbKvSAUJw/6I86RSkZZYTuZKOvqcTD8Q/Qyhd3SF6AK44Jgo/pmpFpVab
9ezAUjq9m2FGvKUnhgUWaAmrC6bSFs552VXgz9QIMqYh/cye0E1VNH5B+xm8oT/j
WRnYrophlSjUiJwIkhlIegEAiC8iODxBKES63HxNPgw6H5gmlEdeuLYpdPlu4JYP
wrG0QAyuIU6r+cAlQf6YQu8I5xRc1re6oNs9o0PYgeho7pzGqCcHToU6mLzwTNB3
RbaqtVXR+ofEwvnxLjPxA/h+b4HepQicoPecqEkbzXmEKdylWCIm+B47n1GpYwXD
NfIvM6VWAwuVJhUpIA2tUzEsbr4M+VSRXZp/yYQgQCn3GFoTnIzegWXI+DHFDCrh
5G2eD9+A1tYZjgmqjcYWE5VtTb3jwxWqudt0BJWnOIk2xhzyjz6xYAOr0ZH/+s+q
O70TZZwwh7ky9GWw9kHA8kYemmfrRB5b3H5Z8YJI1TqQF3etndErKwtf0PPP0VAM
VMl1pkPFKm5fdeQtSeO8bOT5oruolm9wMTvcpcUwg5R90xjLelmMvbZMiLvCa/up
sOz4CMwbLNftJbaAvEwkhD3trdVxjzEt/ZbuM3WRbALb95EWmz9lsbAGJDBD3aE4
gpb7nARwCCZiT0xe1LdNjxZGocEnNbvTSPGrHaI/fULhmoj7xZco/QIohbwA1Shs
rlluAg1hV5aCgqatMu7l6gJTvdTQ9ViuCTRm+1pohEO84we2Ix5iVMI3aA0J7I/5
MlQyZtLqM7cUtS8xpox70J+CXiADH7tZ3RrL7nqg+hMmewH62xI6ICgnOSitggI3
+hfVXaSxH9RdK7CSDKebLPyq7zEqlrp5XiItWaYrfceeXG7Nef4k0ULjklkA7nGP
LZwBM6hXeCdR+QitfbOmZj92Ts+sM5/YmooPRDAQqxc37S36sHB/yHd0gyvCnbzl
+UKrH4tXUk/RcGnOp4m4DdlT/tQHaZBUpfFa3qGwKCe6h+d0bP7ixa+ipP78Xphx
mBtxhldAuVdeH8J5zq2zjjPEVujK4PEzLuRMVDK8YgAXJ+hgMZq3YVw2cghOyxY2
/qlLVrsaHZvXKew9XBwNwbzGz2feUu4FOMZ7cDiN6AOX0Ih0codonR/zuMKeegvt
++xm4cZ+HwiVcR+E7/32LlzopbPA7NpXaQ/94wk9GJPeA4EGe1kWTmm3e61u5ZRE
3J0aAwccgXovbeQz3AKubG9q0JSFg69oI2DdYzzl34EcUhkyo12rlC0m/e/oEHgE
qhWWwOwGF3cwzP8linO0ULhFw6sCUUR7S6V2nYsr2W3xzVi2SQ6yP+d6EkXnK+na
VUBR99a0lpAJVsDepZIsI9iev6cHQp98DwwTBXvyPqxCfIFaHBYJz22NE+VsZ6xA
8YpJeMnRxYTOoZHRLaFOs+9ikU4GChorf6IB0f+kXyWkl98I0I/Y0O2dqhW7PVWC
MUb7GlYnpuo1Z7gNSof4zal0p+vf7VMAoJLrt52fWiHpcfYxH61WBaSsNIr1VOvr
fG3K7vhWdvxRQYm+b4frufwyKMntxNcSNcPhJ5eIQn7tlYi8Df2bSrmdFL+/oGbD
FQ/7ORDcvsqkZaBlVYxmr0HZBPkLMKuM6VYpfqzk8HnidK5+qu+Kl9In8vVfH3es
K9NWHDHoMLr+YrNXHZMguLNfp4UzGHByJ3DMzauX/mtihX07MgB76KF0lIXtvT8a
TM0nBrsXeBbU50gCONddZpHW2VnaYOmPqxXGYccA+OOhWFX50lKivnJkXxh3vYYt
H6sB5RD2TT3s2tA7OHGHfb9zx63K5eCg2sXUZFV0J/rzil6Tbwa4ALu4IYkX/17L
3jb/ecATPGyefJUs8s8d0wd00BaoiFu/E7p9W8HYmFhhYaWA0SaTisyOd0Q8qMqb
Iazg47v3vC4yhtrY0m+CLVkxUGYCovuKPqVvWdt4NsrPqezYPc4VKxHG+yfJqN4t
qr1iHeAhzZvUpo4wbWgHg8ZKpuFfeUNjdrvamDKn3K0BDHX6wj//lw64qtnBu2xK
av22f2UAJFwRFIsx4oOT1YHWFsaFPikQkSHT85GuNoebVOAOn7QFgUQjyoEGZYsy
7ZEceAmszvfEhnTTRtK6zhVk/s0X6tDuKSnMEeT8dZeVY9m+q4m4GfajwCJl7Lce
Wfa+7wKileOLAkXuCFhxHr2GnY1WU87vc84fF33LkqgxaHMyfUF9Jbzr2686GJOV
6ZMfLj/7pVLax7a47Y/pk3DsQkYXTmgTAuOmULwsFVrzpqGB+7+CCo+WfLTcV+DZ
SUJ6Tn+a2kaFpykPWLAqcICg82camQI0IHnREYCtxTWv3QhCpEwg8GSgnMKuwcjH
N9dj+Qp8Zok33FNo/8KEhUf9nLVkwG1mKeScazOhkdXXGUEkK4IOZKXa59dZagWA
LNLwZccKHfQh5/DPZDL4jKgmJpZaIvalUI9nYqnSqeOlFZ+UKtqbGA6ZRMenIusn
Db3iQmZNw5t6Pr/QSgr6pXL1FS8SgLYnVIUuX9Sgn0fcoIo+u2Q49VI+Gv+arO4Y
6rX8Hw9/xbHMts4cFpnzLe/SjZKBOQslYuz0nHh3kMAVIeqpHplqjkaKBerssxkU
zJrZxXN/k1VyjY4dt+td6IbYIWUgu4TWGRHmuIhGUGCpM+gKcs658GVVDvoICcPD
ozOAgCekHLLLf5Q2lJn/v9MH21UAhkeGLWqCxEUgK2TvH6FG6v8xJdNcbb7F+iHp
wu3JnnT5zQJR3ZvyJXNeWxXjBLmDV9x6wEb8iOWEhHcqA6npbJiwpqfcQCtzKe76
HJb7s+qhduIhyvoRXVAOo6J9Q1dZqLLQdb7gL52CaYvQjxYTlKpiWL4M1b41pX8X
EIRjkGwcUUbU9WmSW2pMjCpdSfBZfsYpYZZXIUL2MIGURB1hu6o7z5Mi3/agLS+o
wAH4DiKEsv/H2A15OnntdcixHRbehWMT14tKa1S+8l0v9uGWdXY1hUltAdeCaJAL
JbvQvbo9bvbUtcvyqIHBvxHKfh9Exyii5SwOYC0qwd4vlWn4fNupZHT6z0e2Qm8d
uzaksnzxciuzo6kZ1W6SBf4vQhJdGOFf+H7V6pQThZs/By8CCQShDRC5HUxpKTrQ
G7nb4oqVKheojSySFWQfZQrd15V55GEZQGKOUdiwPa1UH4o2bkVw13WNuRa8nqXb
pPU4DJPGFMs7EhQ7in6vu/bRE+Hj2dn6VRhj0DPsruptqqOJS4IAgZPpnd7UOZ0r
HKYFdMGbJgpyL0hr1hZ0L4AQCmymq/LZoJcSgEce3lvk+XvLL6Ir1w/UGSTWiSti
3IimXs0lbKbUB0536/cB8wux418K9NiWANJM9BDXucNeAsxT8CwFxwW45yy3b30a
G0WWomh9qA31JcMhdn2FM4nWKcq/J5+l9v7KhR5FWQYf+qkZDJthhybLW8dpa+PA
C4tDNxzL1nO+VmaRGM9u+ffFCbBCWJZ4WboPzSixRtCA1x0azyeI9SKCHFOPYSMV
IunonlsijGI9XkgL7b56vHMy+MuDimbKV42MeQYAwKN3YdDvL/sG4gPkXS+jisg8
D9u6MfFn48wTyfBVAN8fEQcjpNV9YuwiJ+TNIwsAMeP1uany1t3+MTa9rqQ8YH0d
vKy8AEWAVxxf++eoLUnwgum+TTuiOAwufVtmrTAgm9dla6Bj3xuKiNEu9fYsvCWr
pBAJX5LDzwLgJeYZbNEaA0hndyEdji9ryJYl32VAALOgFn34Dz6hbNHRzI8Nhla0
6Xxi1vTgZp9sNbmRVJe2G0RfkJBvwy62Fg0+0Dq3iwZJMIOaacAkm0RuO1lRuBOR
b+tTyz+FFcWM+bQjx1NSyW6CTFJISNufLFo9v3yMGXADbMW5GJz32eRATXOfLB6w
He91DDx/LJ5/XrftZ74w1X4SaAnLWP3nPaVdjTnADOrcMsHnuFeUzc2/NhsscKp7
pMx45b0gdrcJknY8DJzoUY0j5qLSErP9/YcD6Ph6/A4+Zu5lFQAIOhMErlgjdnm7
zceX1MBoPlPiAIB4Djt/IYpIqcF8ZE3ceLrTgaIvn/89nUa/F75tKfOnNyIstmNa
BeLlR3yfAO1B7LOD+q9Cva/2n+1PMxbT1VJauBh1PMkQrg2/6K5sn6O6T9xlI7Zv
M6eliYDdP6wEgEq2lklu6cZd/XFJyF9HTLo7oGqMUf7CNRdRzOqamKBwmafWBPDm
Vo/XE2tdIHyWhglnBSPe/8pwbMiVNbbczlN8MIbNbrzPvFlChhIMDaci+dvnFplx
TVluqRXZr8umJr/SxzE/O1e6NEVdMIzqEj9sv5Eta/GgDxGlUW8G7ynaOpNPfTA+
kCNlISO+51zzLSSWVog2MHdvwJO/Enr9Xr8Ss1kqQBqV7hqIrhcVes3boIIy7t1q
da2QC+xtWNJ6KeGwtf3oLti1WyFb3zWzlv+McHF4IETyOzvJr5rBlJJj5I3fg/o6
xe8CGU2jm8zoqiJBWESkpwKlH78X7ke6drl0Mzns4yFqVyXW8kIWYK3fQZhDDRUa
GQ2M8jR8S1r3lpz3XwEytYrjd5EL8pXXnFLTTmiluduck8Lvq9nxzxI5Krz/xgbq
MGqtzt2DGNP2LJp17pXFh4mOzK1iJhp7VWayF+MAtmXkFzFAu7cQgCGz+tP0gBTr
V1imLdx3BAZJMqf+l8083qXVO0GRhRSd0se5x5Lm6FN9+69nQLA7p8xaQhzGf+J9
2VS9ydlIy8DW8CnXryxCgTnFcb72F/sJp6Gw8nPqoWAmkR7/4kCm0OJMnmvh91MT
h6z6Jcsqr3nLTvSR+DiQE0eyFXXTx7+pZXbph+8ZbnOdeLdY2wV4pAKPe/MQhX5j
khNKuD7TYVkXAFZhF+R7Msr9R1dsOmxY0qXstkQwmP7zUv3T9rsdkGPbueW08ia/
0+Q1abO50/npWpbMtcOXtLGdu4gKnad7IhOKzm9X76Jvcha+ju+3astQybybsDCe
4eKjbjYmlMqroWvvRPhzaPHf35fqkZ/GSX/Gmjr0mIh7fpUGEWoYQJTdvpHgD0Ac
rWw/Ayd2L2rXEimZS7HWmK87J6If5P63oG8ggOwhjH5HTSoN/vof1GzduFpwUviE
i5FlgfJr3tBP6BPeCb1+utAVNfMJAPVY+iVTBNiAkK0L4XbvGMdY1p6UtkT/vq09
nCxQ9N4VXXq5BgNW8KbPmDQ9FaKcm9u6zKkXs+tEpTeGDf70stZ++/a0rOxmK1Z8
Zw1svC1xXLXs8uQWxAlqO4qsXZ4+ENE3vrf1GMUYZ/vFKsFffY7AnJVtqHTHFKjb
ujDI/xfjnRcFqlzvAv/AKlZXhosCOuRGa+2XMiq7N9H2IvI8q8Q5zt7v0akN6Kca
wbHApLWsFP5/gq5AhWUzlOC48IurYs3f79upO9GfQ1upf15Im+W5t6/QLG6A70rD
Arky9xhGQR+xhfgULgTkEV5f7O62ASqICDqd/STAGLdf8OmFoEQYrOqpf8nz9PXY
gfaVtghr6w2uKYJGORzGY/9xFXmORiuE6nNSxzl9rmFcttbZ8Hjx7ka+THfXe5mF
1/lYgXQNDaH5qERb+Um4BD3oJA6DyCaVhaLs+4zsCejycl0e569RYENggmK96onc
vJS9b/mMTtcdM/+1JENWwPTQAOtyubECczOHpejHn9MSuZAnicUy9GV+pejAs9tK
xP+l3Zn3rQ0j1fPM8WIkR6XiDyPzupo1VQHZsWSqs5eVetpfnPYzvR0jUxiuCVKy
q6wqU6LEUCfWrKw94bY42QlsWBAT7y8bjMdOTERAuz8RqlZ+3hd0cH4iNqmnhUsi
sX+bvPPEJ3oxMdVeW63jXV3TCUFlfoYdkKCSWflte8bkgLPke6uSNYpKy89OVWsb
JKoU+LB9k0xU67U+5Kf0mVyXVJ1+s5/4GEAjITIAGT5pfbQ7LUpa8HkvX/T73El7
o/dF6LDKaZeC/z8EGaM0KOWW6BCFUOlJ+sh4tqSThxJIA96Ter7tVFPPU/9Uiy3Q
hJQTLLVpGiFka5xJ+2+HEUhTPxM1bSjs9qpp7hSBk92T5Ei8mrFkPZqdSKNF9tFN
uljcY2E3JoF9BRuXgS69ztAZeNn/2p1uYWmUs9zFKo5heMqNpDZYLsQuOOpHg43X
MPSrTwkiNEo6V8kufoKlFUlLzIfLsU3CrnNxqpk4TYbJoUXNXFLP/a31bdBWi3nQ
uYvdFTGdJV25qGuSgWTreZoFmYAjH/Z5g4ZIxbdczQB8KZK1a3w3JAZoEx807Feq
rcPsgkjlnyIaK2deqaFzr/NgcTAQN8KTjrTP4qhnfdmQQyUZRjRoJxJilv0EKs+3
QvfzegvRfUhynVbyCsvQnSdzucq7v7iQz3b1CJXPOpO0FDcYzi4c0xHoExc+vtAq
3IfkVAda0sOOZ2bRedPnGQUdjXUkuU3cOirGA99QdOUU6+vl5ekEChz9bYaGSpEd
i0KKZha3GoYuh+2aHnuv6+kKhN0Ts6H3A/+iHefxY5PlmlsbA9oNosTj7y33jxMc
OKW2Vo1Oc5vmaxdbW38rxlAXHMqo9sd3kTxOvjJ1JNviL9/k+rKK6Ux+Q/Zwg6Bw
00jmBaLiAouhlwegB16f30UEJASRdvN8R97s4yOo1+KjvPzl46eDm76MUW0CFxKa
kLBUkAz+W0HF8doZhbPPTdmn/5qZ5N0Fg6Fg6BxFtNu61I3jrGX5ovHCKp27Ofzt
ygJW4WhXYJmHVfZh/xhnaA3C2AkM4Z9RF8LGTLsz+5qTn0PQP4+ZDRYx+9E4VQDz
wypWGZDeqhnxS/MLKIRlHpEh7U1qVaiQ4j9eGNGmg0G/a74u9M8JPsSA8Zpnw56q
/WW0KHxjhETqOvYtSRbPFk0vIp4/F3GWsQlC4gE6DGuCopyMpeb1oDo4GTvgvKCL
7KxOXGRUUP774upb27qGbEe3NhWMI5CjiwhWRDTu/+IHbt5t07gxoqZFRFDHBaJB
ucbh6D4Ly2FUpij/IgyT05cYrUckO3039L2Ug2A3rXU5qroKQiVvPm/b5TeT6ZsT
6yRMTpQ3eNS+bz1/xO3P3/1YC9FArSkfYEvZXEEXGwBIDa3h/mi8l2OouLNJBipM
4H70OVIaL5obzaGjiyM16vMsa8bFMTTrL3738CN++FE2iHixM9Y9nBfpCHw0oH0h
zGqfLsGjHMKu+xNNko5Ogv2IT37t+Pj8BCSZ+v0ywD2aybJsnawnfJ8na8Q+Q8JM
5Jx47ilGkqgGYc0GJnovx0fklInokvke7cFH4AITIiV1cshweaDKRixv3l19Oyk8
fi99kyx7+bAETSDN5+4WSff6KEJoeL7O7pPuTXdAyeTqFvdoZmTeYPJk5Zpnn9Op
mV24K7zTkBFCT1GVXCX50lxRB9A8WIvERODw/rIICmhWibeTQluNeZrqFAwspJf1
h2Dx8ly/kV1X7hVlYFqbsu+C1pGNi95lhCJ4ngQvgkDBu6idhejktCjap+iN8qgO
wS3b+2eabmW+RhGoxMh/dV3GpPvsHVlWB4dreAX16x1i97azaf5fOemdOfFAk0R1
mym6VYxgK9jCuN9NjsGEZEw+RSL6FVoUppqsinvPljCv3Nu+jTjHWvwBeHtKX+z0
hF4Oybk90YZYa2rRF1uvdFRp2bGhWUV4kGM7yaLjqOSmo6T7xU+QaC1F4w2ahr0j
8sMewr9Zfv+Ps2eMnwugFLcVLjXUjmbGdip8dLioGQoENtggoFLVDnPwC3rkygwf
SiANboV3ccH82mOtFG4oSlKNNww8sT9zaNhL3/6rxhXvL+GQhOklA69LzuyUw7Ow
R6LCoOecZyIN6uSsZZyBaeJHvZGghfULleQt40gdF70SsLIW1V+HzCKZhzoFANbc
EWZr/qVpqI+mFbqSJjgVXpxUsJbPBc8HlUCunoYNEYAyYaJbgkEgxUSo6wJyb+3J
pftcEMCQUdKCogBitiU0JoCK80z78csYJ9OOKvMgJ5QX2PiQDjGb44Xd9Xyn0aQl
635xIJmWxjZ7Lx2CtdSqZHtrs7ecgQfFXs1dh48OtrL+YJ93LFEoKrLm818RD77k
EozHKO+UA2RnQeDkh2dPGPKpgCYjOAypXDtdaTQxuxIW5+3lc0FUCpRZv9KwCPs0
H/DY/2MWjuBMl7A2pNEU+krbokojsHNZQZKVvyqKPg/tcLpG4UUZP0GYXYi5iRfj
tCmBE5eI26NMnNnYBkjpIVkCQDX1FeQ1lOycRTL8qwRBUVAmOdV1JO6M8H2mzTcI
TezjJg39XeZYJmb4SCJqpB7c3b5oqIM3NNRto+lZDx1vdUxKcB2j1rK2dpiLPpK9
IBvQxt1cw4U13I++qSJMcq85VesdbbHVsIu3/NEEvJhC8T86qka8U1pPTl2yX2uQ
4GvhGaBuH21+RE+fJnZNjvq61NFS6Q2pGhwJeCzvwGS7bBtGnXmypkcUL5A0Owkf
QgDqhFqL85tnLLb5rOmFZ8NusdSSpGN59422OleHBivjdP6IMlnArIl5SnFogBhA
xbWHGkEqPWDN6pyOkVaTq4rGOTjQo4gcM41NjYHEpkFeRFHUA+b82klrVCrwnaZN
Wqkp4pAwkQbky+KH+SggMJYhXB85ggiNjNkD+Ly1zoJkRFDDNOxkB7/notRFpatn
LNl0XKYiHKdP6Z4SHtQM1cUUlKAHyGAUEmGM8CZ1vvBdswT3Dsgr4PNLrmMJlXQR
Xfv7QSm+nDLYwYBvolDFvsHTJzJO+iwkqcijLIPQ8sgxRq+yloJ3SNLKTZHU+M2N
YXBVrPUEE/ld6ohAqHQoUoRmubOJF90cLoz0A0o+8frBFenT+KfptbxaS5+/iKwT
ZwQcxfg7ajoRdeIZkgOTNMAHO+EdvbLlfp97yszmL+50xg6waOLn0iwzRDG2eiYV
DfRgi+sdOb4m7uT7pS1vgKcgKhJ0tK7Ep2BrZsp+R1ame5eztqO9Woswb8mHJusw
XWNopDns3QqpxipbCRPf5QNQ6niC3Imffa563nSZN2cVUavl1VYgD2FFp+bhSmVH
0Km5ptToSCxA7SabraGWpBGL522rhOsXO06Djq66OJHC2EDP+WMjgvna7lfIrT5h
qT9ojhNkSbNYeZelXEqu9LBCcOyRUwLFOWyPp3EiCyUC9CYNanrkM/QUIeMESjbP
Mbq8wEsZXqlYUtZ5n2IdCnMRLvSeHLwijRqT1Sx8eYYuEcn6XXHMjhcsxF6XQmPu
822QSM9+x/mBxGiDIkD2uUAez3cA0WXVHIN3BL970JaslApU6aMDRoCh8nY/PNam
qUMkJsN7s8Ay16yhF/ClOWWkNtKTRkqdjI8w9esU6y+I+K4//mzpf2jAKyFlss/d
a2EdDxNoEDYwXMvrOK9X/kqSjZGaeidiVOnGxVgGkvnXllnJSts5nI4FG5zAaLEM
Lk7kSKNlm8UGewKdw/p06kzQCBhB1NuYVGS+veTdinF1dsPGo6o2EeHfBEn5/DXa
zSvcH4jQqyUnuRVKG49fCXr5AoazGiL7/O9ryFzd3qNSHIy0iW9DExGQ019Ol4gN
M6hpA5RV54AZq/m45ZOj/EMLyoWBRsfSIHpDiGV2mdP70sdoYB/7X3x17gDxJ26O
HafIcXfEX6bBAZ9/jZA1jW9ESwKOyDL7x53AgegAGgKiYI1O13A3kRFrOP1PXYFb
JH5HmWIQCFOAAGUwDhehDW1BONGHi0hQKHr44J7TrzjcgKIS3woYNjM1HEyjHxij
rbvbGHYXV3Jy9jiGU+wH/D2pzOr05X895yCjI247S15atO9wSNjU5X8EdSoQQ/qv
ukGQ9kSFo6n/4I6ta2WRkQrdLUbGhhzAyWEXNZ3BdNPDdq7/TLcFMFmj/GUNF07s
74fBU2hHHKYSunb+NeceCIhl6KJUeC2OzOOKv8bgI8zMBoBmSdclw0Y98BpVogzq
VlB+LpRQZaTnuW1sgcND+MVU7DcMIQs3JZLcBO7YWbAolRvgpjaJAgB/qqOIRQ/7
2LcUvPLL+D5ZHbkGzrYVuAPcETf1Kh3Lgf6QqZ7Q3I49jq4Q5xsohpNIMpNJNYus
XTfALRpLhCNTJIqoks05PNCZozcemAZ+dFP3KyodALb6dJKQgjHH51fteqqD6Mxt
aP6B0TPzzrTMIFDmpCKTNzmlb9mXw9Xwy0KoSniHarkHBkwmIR6euyQfZNAQUZ4K
QRdvYqMs8w6MbjdxtI4fLnuScb3rcIC5Zvx7ZgegiI5WERP1zY6OQrjfE5MTB125
FPBpvkjwytt7aIyIhRmvhof0zBDD3CXQ+nlWzWcrF1lHW/OdMsWPMYcq0OJwZN6a
p9nZXgEvUyChVjylZ5yoKVHs8Ompo26/586j/n05gMfXdnYpRXIOr0hJSaZgfJQT
FEsmS4IE330Ufi59VTZP2nCxgMpcMcnoafiWRJ6ddWYHGuyyAvXaafAT734gbk6j
ezZHitunV0j1ceVKyFXsvVL1AXpbQcrYFtCY6eKudzResDTDu9KUALVz6I+MpVpU
s7RTQowaicfXdUPlL1Xr7Z9XtGzgEticStT7z9a74Sxiqq3Bz/m0RQWDMSn/44vk
4JVJOoXTODyA4yo9TOwSw91uAqn4nyhlXb05NWgXVOtXJb+DcyTlEPboywSWAUtM
nTMEXQV7imhZn7ocXZy+9Si3R0wnXUMhTB6hjz4Z4lp0fM3lQdItK/A58yJEf7V5
gpOrvhc1cNU0OlU3ZPOKJkWEHqgYZZuki26DvvvpugH0ElOcvzSHY3jbTAhmySMe
fe3ugY9mMpBQral0OWEdfNLSQ/dibV2MAu0ieKlYzRVlw76tJMd/P6HwJhdQyjwm
vtrJK1s+YGUR2XhonJ3qmOfJbZi+4cg4z0A/rE+mrjaGvajRjCqGYMN+K+Izz4ha
1uFAtpc7l29CGwbwKToFvbAspNaV+9A8Rg1yT5LCj1kLuI3q1gDPVFCHWBfHhyU0
4F11/9faJaOSmIgTm7POXtEPeAtWL/F9y9HeyTfVJwW4xSjS625jgSDmFbEtK/Tt
YyWHm4qYAbilWwx5jqywwVKBuLxMWEzP+sqnDDNwfQcQ/PjOWKK0Khnd4yfJWFDo
ViWouXT+9l9Ccpp2X5wuzNsxSCJXIZIP6h/fooyPaeC0/hE9yMLzcQS2F0CThxJs
EpWjCRJLxIdUYl5/VfMFkPWb63dNSCNqELdStMEAYKo+b7WKvgd4zpAXMEAsdcjV
94yVYTB58eCHuierbV5d5Moqq3J/3Y5Ew2jldTGuCmR+Ilzc8vLcGI0kI69M7Y54
igd7HR4lyZLNnbHyDjH2I7LpD3D50ni9ViubYmBsGRv6Y6vOYChr9q/3SGPaqMQP
guv+ctdAgtWjU0fG9ze9gxmzQHZycgYkPjBi6P3TCsXwNTLn3T7F6CwYA8kUbxUx
SD4I/6ITJY84pJIAPLiRFRxBF6AZ9p0ay3AlJMCz84+SlkpeAnIXfu3u1he6i7lj
jwNyzj9mthMn4N694lTe4HDx8fw56RJSp8qgv89Wpijvh5ePw57UUVYHqfppL75Z
ASH8dTsDF1ffmNYAMNgZD5SLqgm1AONzT0jtrD+lk2I+GXiX5zvoI27UShzsvPTw
fe51V2k6CSsCJWj4/oX324uvbQwzjY3RClZbwnFHEvIfgcpolNWIUbM9o5LN6xFN
yB59nwR38chCM+YVxCto8NOHZf6uVwb6woGzKxR0Y5PZEJIySMLFPhbJkY/9ofAk
ZV9fkEYHOKhdHvB9e4ux0GJ8eTHGb5Sr/v7qHFH0lFhk4WMCM1feAeUQy4GP/9c5
r7xbtrY+cVrv3ptgkgdjEFBm08IfSHRi5AHmZ2yQ6nY4LY9iiSxqzZCFczlO+f/e
yEBz3ZN5vHPxYQhgu4XOJprKY33rcCTN6c+JD3Q4CDKSzrHFXC3myIJNbseSjSM1
EgERTaiWLcBv4eC+qKKjKw2K3gce7sjrDOkt3seRBfKJu7KYLOV0L1HlfTeQfo/K
PQMmGS3yOqj6Aj8noTnyQqgGUsfTUhpYu1nCwvqvqLGPhakazet68rs+QBiKNQD1
akPh5gMg4y4bLUV57oqF0OvtT69ea8a+KOhtQHrBzSappBgNsS0c4MAmvMAvXzYE
Qazi+VXg3sW/EkLCsqdvQQvKGOMcxg2RZWgcflJsLHlUCE/oZuoxNjsIwKOgi21r
VEVIcD72ebDfr66PpgjVAjzI/H38A02zPg/TuglsXQ01GyetLNhA+MSHspEgkA6x
JiYZO2v20YMn61IONDcvJmVBkxjm3GCKfMnzyj1sLsNfwVZVmU9FXFeKJtugXxah
Bm9oF+XAJImtGvIYRPVTH1sH7LpLd7SHSvqWK+z7gDBXWyMHDnKGI/SlMqY63zs4
PJxiY0KF/fThXeQXFODqj0Z507sZt5QU5el7HpyJfIlwykjDNFrB29Lolw0dsJEt
OvIGLbKrAOSWMrMpsRPnlqhEdr+EfBd3CZe+nIVCGxTiVxRtbbemAlK1k///mWXo
fzaCe221qfeyDRCR9+xXJQfFBqou0fC/ch+lJMZieLtgU4aREbhvrcjy3D7YipQp
rRoUaSkBu/etSkp37yDFRH+D3byeEpK97Pftxryt/NcWcQ+7pYhY7koCqcEWw93b
vvmAuODfi9fojauy2TfbQ9T1VLdKcNDELuuipwSLr78m/vPbOVV0zJp3PUxg0DJU
kkMs+XUoCrZ+F7dtbz0XNbDGxWCTMR60j+U8fipkeOsWRYLqV5acaw1f5EyqzUJp
WTrT6/hk6jppcXoT1ExW5lx4w+HABpMOU6UV2iqR4FGUF1fHFrSq55k/nNK//9X/
hFW7XD8APV0iMCl0JPEph+FOStOHQLqJ96MIhGmAb/e2FcvNbidcnIrR6owP/75b
do6omiG5apGhcYz9JfY+eEK/dznKdyogBlxjJBwLeGMj13RuQNisE8oqxQeuOKhs
hG8aBNKVo8ipYDpFnaH6XylXoLzMSrzFUafIiuXUbtM+S/dJMKfubLNYPspAQGtn
zmLv7V2bYEte61BzrWc4zw+/+DKhyuluSs+iyWcgCjxG7KbG9bgiPW003T8zux86
ug8+SD0KvfGYfEUUCrgeAG4ZV1r3g0jiALg0koJ9soAtHuKhcj5bqbq36aE9Z7AP
cKO51q1nIxpDTVQDg5nBwnmutZUVpGNIS6eHMaVpeMDat6BT85GX/W7ggnW2jx5d
G852MfvR972f4D93azaokf5q2XGsUqFm7SDVJ4EM4CaCw2qFBLcuyXrnIX9TzpxW
yDOvwUDU2qNnHtpaYNvVTAyxkvcq9kJRNw3bfyWogqbTq/hAts+IfubHBsqxxSut
buP96UHAKncbuJOEs5Zrd5bYvhWoSpxqRIcNVQy6tQR4pR17GJW9Np/FHkwRQzTS
yUec+sd8/K+uvBQurG116d52VJeDG8slJH1iiUFvWgVpxVDeas60aYs+hp5Qm+xi
kuZNx+3OxalpCCXLRcXhYWvw4nYsiYe455H/u3rXDF+XtEe6o3URatoLa+7Yvq8Z
/tkTR8aDw8NUvsBP3gV0+aagbKKA6KPE+60UynByop1kguTM5h8HWuQi6YrmHQyj
S5COLZQxIDXIZSMLD85koct0E5Z2fNfAG+P/jEc8ba7SBolUFC7DsyGuLc3PY4wE
LN08aIlNwW3BHjS2houZpQlARk8F1BaqLyoelrO4aygZOANYngpH7D4NhjmWc5SN
w6YDQjwBIjqLhZtQAYl1k7NnupPgXfL0kF5Iz3vUVHBqE7ei3tgAse8XdOe+Q3Il
iCwNeGz/xSeV5fWaHZNJWAgLrP//7Eyd1HvKtwbIxYM7oNrh9yKLzVm6Jhvk5u6Q
XWwtQH4OqZKgKXo4chyhYbPnhkKTQn20BkaiQ1PKdCKw6yQY2alEMwHs1Yj+EFsS
/kqmQaV/8G89jnxv6RoMp7NRip5/tb2Ov7RF46Zee8Q4JvDR/5uOwko8B11z4AGp
+GTghNEkoYlpFFa7pV+ztyW4BBENVxEuvI9GKjXV0SRIR/hFWcRuvfDdahLPib37
dP1XD9cVawbWDv9NM4cvlJJ0lqOKu1D8o3ZlvN86vXlrw4FJPq4TeGgNdVf+awnF
e+gcgOoKasbKezlhltW9tq4AT+E0wuq3fWWBu9TuzC7mxUKBgJIe9BxkUvEqJJ2U
v7TKvOQj6VROVaUnVKY2+ToMvN1f+LXMzMPG9oaMvY2LtBTAhaVoRXVNYXCxmXaT
G3teUUn97h7K9+SyRG9tjfGCJdtCkjjxOV4UGiiMa59i9R56mDRX01lT1A9/aKDK
3XIvekBcgc3R3qvI5Dp7GkVq5mzjNtcFush96lGjX7O83lwWgZImUiDNUdw4r39o
w9V5oAuKOk8pCHp2PguHwqL3CAWbQ4irKhPWsHdL5j7DsMNM5EPnhR8CFTZiGPYt
FbzEK2lC2cvFnBWe+VLYN57PYTWoyUAGbRkJ5ecRlHRVG62ySjITLfqWQdWtDAmp
A8AvoBWerTuUh7xI099mp/MYgb1c9lX9FbMgdn4CcCXzMtCn3TIhoOBdZFQwj+7y
IgC1urKN/jQ/0nS/nFXhNVgD3/DY6Fla+AebpPqO5e2SDxjxXOLJq/AKDOD/TrIE
1V70w/QbJf1ARr8WAkv3Ckvs15Q5pg/T4VABozB81OmrlpDMRqqOygRsYi7IWG2t
UbgdG8OTknSF5+Ao35M3NwrVlu6PXkiHxlhY/YT5q2X1BgOQP/IaZrr5RhfNNKMP
K7jdNQIVsUasM8MH46I4H8QQWurQZwWaT2bov8JkFY2kvLT2Gv9Br4eznnY+zob0
WxZqs0bKX1rsip6z3/Ba+TzGImE5dAToe+gMklDGEhqCyfrRjFYkWldNGAY42nA1
529lApJ5w2EIlEs87FBZW0Xp0lB6xRER3XbngxIeULu4sXKPLjrPU7uxXvl3bN4T
PTW215nKIlA8m9rF518bKpgP/VK4Khq0prtQu1LIm/RVFO1T6+OryYHSCH+OtRtB
TO7TfSmi8Ufpm/FferthX/4BwATyrkkJdt/pc9A7aSu5RSPf3aU40q1anAQRvwTw
6xiBmkIRCxK4LdtezYr4srht7xGVHKb+bEYEgIaJ7WbDhFH757+Fz3/kr03M9wbP
xF2GvVsQ9WdQaUhsjg2dDEnBuyElgOaNndVngozTnMv9yf5pR4Y3Zt+jOZff4aZB
iwiRygZotqCD9VuZLOWMcEzXhpfBVdgUaCil0kYESNQUibwwJw1r6hUSc80UTiRW
sy1zdEq2Cy4qQHzm8BaCSgH2Dk4vzJbbut96GWz1VkuPsPBUt/X2VgDbTMNQZMGb
s3CiO30FvMYDcEFMRbOYmNz+eUUdTvqlBwrLEc4RALmc9ozNCHzGTEHvfgwxe+h0
c4qYFfPj+hZYNBOIXMVfv0WGz4QBQyimhZ+w+wgR3I2EJGUi7ntnyQ0fkXJdh8+R
KTh7fib6E5SqKzSFQ4BWnA/w3xyW9YtKJDIVCsP/d6dyZXVx+gHedPqnPFBbUZZT
skr6c8bALCQ//apMCKYVIfBn9lWqvOB+YlpUltbqXBKYPDYn7Ahgi352ytNipnDH
iGpACJdOo8t9JoGhmbPj5BOnsa3a80vExCV3cNNWaOX7Yy3uYdavSp400Ap35i5r
Y+FmDWmmr8wlTXghp2qLioLZoup+4l6wanu+PvWI+tFdVwogDd+yx7tLuA71xXwZ
e3pfQbmI4m68pO4HpN1pLNVFMzsvivNywytbdKH/JmXW0sRpsbwZZ8rm/dVojVg1
AjU3vptTQ2cway01RyII8FAGND3Yps+O8CVUJvzBWW2DQ/oSFuLC8XiyGgbzK5U5
l5g1ogcUUv3VtM8mg4chNs1uebLKicCkkB41WO9+imwzj0JFqOlarLbExsEJ4nG3
mo4X+YbVtVEcLRfOIQGVKeWJ9LjWQjquGrxLIBjPikSyiwxC2KBsS5aVnyzisLNs
qchvS7yV/I20bFyj0IgYSNCfYdr41X46zEmeiuTyWYmcnfxogN1RAbmQdE6zbwjP
iHo9cXQJd2AXyqrNyvHifVoz3ZwfTTh8+Cj2rtgDkj19Q77VuG1+yRaQuwL/0Ifh
ZWy+a4rBkmdqseBL3RtW1+dk2U+e2/HFqACi+urwDRPd/6eZVOx0ANnMCcTelMn8
tB/q7i0lqk2Vc1T5aILpQA5ZxJuAMdHmMMLgiU6ZEH5a4TNWt8AB9OIIW5MvwMGj
awlQwyFUUZswIrGlEZVMtHw8HHK1hLU/sikmgi9qLJwhgbS3jtuaIFJ/YMHCCTFa
sq/Q07A/Ota7Y+DuhMAYunq0lYkJ/Lny3lr+uxFUx7Z/cacoT8TyDmqwFDbB2jhf
PT05jR9w46uFhByAN5HFJLugCZMHVKMKBY7jDXSIhm4N4/+gGGbqvkuV5jIAUbua
U3jVpA5/EqnckYkLPkEaP+U2PiKH0vzRNeiaSrG7ckVXLVC6LB+4o2xTBCiP37L8
ekSsqPMiKPf9psy0IzQUJUbcCDdNfjnBn9tqbAmynXlEsSoUUMF6JHDCmiOCw/2w
RK6UFbma+tUcOF1VVkmGXufJZ2h1Oj2BtVtAb5cKqDjvyXQcehxe/RkRp3akbsoe
7LHTueq2ifGZcnoHosqkjuQZEiXzP309FWFHP5YWuJ8z24rlRhZfb0ad5KaI99AL
fQZ5RpolvW9ILgae2K2ym2kw+aVUGfAxvQh9ELmqa0FfwuK5D8f3XL9jnuOC+Xtv
LPc91hfw2izzkfSVvTjVWfuMwQVanseDNNE7EXAUQkFOwudAcUK9U4e4NrXPCwKJ
jKIfRJRgPsO7Ajh1JJxl6Fk9mQiZ8XJl9SsCaic1bUMroolLSZW0wsnhpy/w4pAx
36bchc1aOerCD/rdQJXiORAObuC8vptKaifOl5bG8TJV7nl4yBSxNKdVwu13Ooqv
6r93sZqvGo4wq5e5AL2TdjQM9WEzPp7D0EdQyFuwQkI/Z1pnF0csuw21uk2vieLT
cBuCjerOrzlsWLHVfDIN2SiQZo8FFq3IIuVYXOX8j2CRd+kPKzSDrVjavINYzr2M
RHfKwk9oPLUt2lwzy9faweyg5egZ4j6IXm18ruJebg64tpAfuPmvj46j9EO7bQav
1aYxgPQ5PgTBqRk+q2pAYW3aCqJoOaVaLcaa7TkQwDhBQ0qMxgjCmE0t9C6DrDaW
auq9NVlBzv7pHDSYHoDl5WS9uikvNUEszEZe/D3/kG29N8SEvAp/dYyEvW6NDHcB
eSbz3o/Oy0dakv2FYP5rfU3kE3I95zqVoPdqSIWNIYjbWJnsZDygewvKdf+FIbLL
k6SacEUu6iezlyktbzoT2sopGS/OUHlHpBYSmtOm7bOTj0fs2fW4bE9ht2bGEy2R
Lp83eMl4d6MCbceySIl6RKv8wsBjxJRYclyQcGmbSSAyqfqVxF7aJ5qXxrjPjYXj
CTqs58iSRkI6hihlQsvHJUutfQ9JujyacBHTH2w8uERoQ50mxGVA8032NIBSvfyG
WV5xVWoKkip5TyUfBPLZGEtKsavItd41DOW+G4zyfmYWKIGAfeiO6D8rb7MU2Vcd
PAAg4nRS8n1YpL/LeQHUQcFvUPCrkMtE4dOMYM9E24e3d5CytU6ZHd1RCGztO1pN
2a0AtCr4WALj5IGYztZJ3zsmX9U/aL6diZ3iBDk9ySOGoBERF9h+jMxKX9xP1w4O
OnTUctiik+92oNE9p1WUo7MwJ0h5bSWKas0DTLtbUfx+NNzNuOH7vFCfpn0Xvr22
14K2FuorgYAhYhbsTo9mldVg20sbYBuD0PNrFmySzdW5eopoN0AXlpqT9zgugnl0
CzrHXE0hDnXkwQsvlKyGt+Jx6PpBOg0e+uAc8aY0xZDPF/vfc1YbvhFTRX2ixX3r
6GIVsrv59LRWgHTwD4TaKbyyjCxiPU4iOTpr90ry6WlYr1IMa0XqUgoEv1pY9gGI
OPOwX6DRylgB8kETBX+E0SavZdycRK3jg9vtTDfosEjQxr6ruJn30iwUB6AfNue7
wOj7N4kD5esjiN37MiQ3ZqXtYajbWp4K4rnTMhJtikwuOWaou7Mb9cjggSdDZrXk
FhVjMDFtYUneRt7iCy0SuIWtmIqwegSvHx5ngd+wyN4QyxO+jT3vm4HRBkc5ZeeG
PmFJbIIzlNhcoDvI4D8GLAvADCR2v5pC5ESkQ6Tm0vwr9mQoRTJETuAHWFr8Z7Wy
rY0PFjjz1JE2DYF4PukDMUJduDvdu/MY+VxpMfMhqeTxBzjeiTwxi8NvtDoT+7mS
3SrcCowXp7o1+N6IJLWgHdcZdJsq13pzs89dWOtkmCoOlfEXQVDzbyhaL49IFUqk
wwzWfTwha3Fea9+UZk9UV5NQJG+rKgAu4TMqMWt8V9ZjAPi+Bn52ubRtrvPk+e+T
wOLeBUcVn8jZNavFO4StuuyheHZzkdUa3B9d7FsmwCko4M4u06JlIc9CCeUxBgDA
vtKy7NpWj7W68KDgfLjpYq6q0Fr41THrLHp6C7pMq1wM01J/2wk53a6xX848wDsX
Q+scsJ5P+jK8G82brmCyxRZJeb1n4E/4gq9QZ7e4OVVQOgCtAb7bTPL/T2s14vO7
sSVfY95G21Pu/fngufnTOjxblLI6fch95eHfRSSi0kE/Nd19QEHHjARQcpjqHL28
4+XJ15bADyHRDHq/n4dOX4u5oxKE4Ui/TDF3NVAlSP4tgBDn4e6ill/hANVqnGtu
jO5absVCIN+hlht0DpZr1d4dI1++Sqdzmg1GT3T38bl1sf10JAzR38e8aM2FuRb9
di+9FnQvN3DTL5HCVoj1Ac8g374LVnw006nFtnLRBVgP+xszl3ijccbZX9l3v+Di
GWEbEZ1BSqZCe9cv3QWPq1gpjIEmVGXg9nY+zpb2uR6ckNjHTkl33dJV5B9oyMMr
2RlNw4pzkSLpQZHACcQWfASsvuIB6sy6bV8H3lEOk7bc+vxW05axtziDBCKQPDL1
yBFMXRZMOgG55OM2ZDnWckBvS0fJL36KtVyWrT6px3C/E4iAN+q2xOarBxnUdKKI
CNtHjEh+fZMsidfQq3nmBR9/JxmF/pebKw1FUVUFG7BiuioK5bGm/txsw0KmNqdh
GJckWmpbtqP5/hD77nKs/rpJO/RGwAgCynMeuPUFwOabd9NkwG/Mx7ocXoXaOenI
7l+/nxMV78xLsocHg4hMcwwKlzG3O/a2pM3K0UFxXZ/PfHa8jHa1tLSl8hC0NVyg
CLyW3hKtv7gfs+0M4DjQgcVjPQSyEBQm1NkpcKbJX/tJxGg2W2cQwTK+e/g2+Xu5
y1GAaMZ8xn9mt0gGLWeoQvMJSZhh0XRuUFoN7TpxSa+kWXn0QCKC9vW69aK/eJai
ioYkQMkNQMeNEZP4WTZTVMMHy5EcQhbaLAj2CjgVE14B9jyPl5WJBL6z79GQ+HB1
xp/+Cgx07gCw5tWkgiHP4QPtIOE6EPMkf+ynZZ5sVwEKkx9eForrB61PTHW60jwp
tZxVo5FW88iOUWJ2t1BWbRJVV0DQntLmZ5wWDmuggZi7x9gEWXMpLKwBumu01gmr
uphRQMG7Djp0UcUSyOiyWUT2LqkprtKReVw+GeWutcGlHMIIfrN60cIDidt99yCX
1G+d/LHI3ouBfGGZZ/GFls+eFB4GPoXEAt7+pLiiuW91jx1oUCl7KK35TuNSlZNs
AMmIPBjeI0A5EOrFabYvAfZd8EAarmgFLjUickz+gioYjwiDm3xMIFKPvieMDTOn
N8NHK9ilQbdBLzjPXUv/9fsiPvyDjq93FN3ycfhaKlNoBY2FPKZ+EAAM8FD7g4oe
4hgFX24d9PywKDrBpqyyjyq8ZYNLMIxq1ve0ZLcxum/ohaUjCZhS1rn2TLUQynKN
5My7/A1L14te1JT6pr1QQnONNcYXPXtSbWxPybMspvefEYIWFzwQONfEvt/IIHQn
3c+0wdD6x0ELBXHXzAp0FIF7wV72RQc11rIkC4t/Gho/Hn7o0/awvrifTyuv9ilP
WQSrZIyYhcyJ2GY8z9eUfNUJ5fJel/x19yylydR6ydIHQrkEjatRFIBtv95Kd56J
aEr8qsbzZeqbqzlj9AuNNnwAaXNW18CPCK7HPW/WcGd9JZHgevIJfuicZCXZVh7q
zrflSbe1Mmjo3wbzEik8xXSV+nOvSkl2JjdsEb37PP2QVMAevXDVhbeV3nPbMpEM
mqznluSkvAmCtHGe+kUiZAD3avOI2RsAE1fbbVPdrpVqIPkFSpP5ous0uRJlikBc
+BWX29F+46TcGdyTrj/4Ow61LLvPVClGPOUDx7aLFHSmZHJk5c7ygj14bAVczw/n
vRyIF8ZrvlIiY6H2HUYVos7lpBV3cbXsQm9tT/MWlnx8PNQ5HbqmGqr2K6ocSm2c
sWVIwIcJdaBHK+ZnJAHhCb6ZhS66ZKLdNQ90vrtdKWs/j+ldMpW7wjhRUf4Lg29H
dQwPDZ2ZpR6XaY82CJ7FA0eDIi3zQpdS1irPQqPFp2tM1kvO9T5P9plpQyUCYdJ1
dLhVo7eehFrBUO3W1yoKyENE6Ep8C8LNwSVKnxpmTWpnrjKYOba9pj7BALLWynLT
chU7qvr5o8RQJk/UsTTSqINMDP8EeuiqO8ReeSkZeSQ6xL5SiqTri12eeA/CxG7K
xDmRueaVVHF64zOcdUlO4PhDoRDd7Y6i0sfKLyo3UIfYo1Za9QcfguE3XTC05sBi
8hKlAlxts1NokQW9fvb1w+qK2W925L8q5EBiIpSdmlg2JcEv209PD9UL8/7b5UGg
PSeH3ytwZT8663qQR2/Q7ZwTxasrHYa6vaULjBQgvGD7o/tYnpWe6qo35dBFWlS0
pWZZPAI097WJZa8UaPIhWnfmcvJ9jhlo4zHniaovylS+eiPxkbsrdiLtOXtHdLf6
M16Zf1TxEVlsQbUSm+/IDvq6c5bNu7CY0ck5RmX62dP3ZO8AR8AD8FliYm2rty+6
iMJDDxp19FaIEkBvsL33HEFkxUBMmqL11QewPGrq/kAobeIVh+EuzaQsozHcA8v3
03LCoQCiMe5m30Da3UrcCrHdn4/zbcgbfYc/CReEVjmSVZEh5Tj2W7xIwFL+vil+
N+mfrO69hwxSFyIWP1HdXqgp0rr1SNj3oNM7b8z25RatAU940LCY5AqaXuylep3U
jPgeu+lP4Wrwbkz5rKC7Yc3zSDcUk91CJMuDEa6k/FkxY7NxPYisXIAgifuQ2mj0
OyvIs6287yaIpYkg08TH7y8DIGcUaPbR51PT/NtF2A28+dCyCEHqGqkRb1mOqW1B
GJ0SjqUpw/0w8W0a0Xbf/93GKRrFpWf9yAcUF3rmVxQ4fjbX9lP8UDt+v59zoUcB
FDFK1D1m4R4+hZvALpRdEKZ5PlYnf3vT95wqV0C3Lfm3pGayFESHJCrB2kHmVrUL
iyseR9yUqN64p1Tlg2FnICPTv3M89Hq28KFWi5raU0H5uDvJjX5H2nQHdFFl7mDW
P48JNZACbFTyVOdHfbqObiQlRKWOA4i/36DozZKT5/sxzTuCvZ1SVnxIJGCPJ66Y
yiKmzV46UIs3Bpew2Y5KaO23BcfZl998bp5JnOjmW+/4cCPQVu6T5w9FPtuZBPeM
bKeNfBu+UInOEsrNb2hA6ZuvpDSvAUAS2L+ZH5NZmp3ckiBq78y/wvAaFHbjdtjO
IFDJa9bfWR1JupzpllfqStA3ndfEfFp7qfuDeG05UxqV4Kt/VVBATw3skn5HlVRG
S39goNA8oGl27I9FNs0rjHSJYi7xuuESpCzQ14B5VvLs1CDRKcxoNazSBAiRtg2r
L6rzaU7l1QnAakCVwPPIE69yvqMCYS7BUiKv2t2nLpLdbc4dYaPvyi7fNdSlmuEd
il0r/1A+7YaoRNEkLwA5krZG23ch5fNEvBoU4GA2sWZYJobTUd5SJRtywT8x6e8F
X5DpK6ZeQKKDsVEUdzPCdtv6/hhsR9KFiItpdmRFwvI8vvgTCIazOUugDuOJRjla
HBolZUsivpqZlaHJpA0ESec3GKZT4KVdbbJNNOi9+eDyMkHnnDf0BBICjdQimgI5
sT2P7XMBirZelWsCdXlGFCpHPwWjGDykA/vXbrWbKIOOY3m/HU3ub+Q6ZCNrGRGp
xCb89OoEthYCmq1x9/xI9/GWRzYH77YaPls3Qfr4KrZvYZCKEK3SyQyisLvy7YSF
gjDO67rJ0kJ4cvoZ829CdWVs8g05IEWLx62ZZtzYhmsh1gJDrS8FKaIH70GGNDlS
oRPpMKNEEeXUSKUc5nDswTVleeOFFTlwYdAX91K1YXVLFViCSX/xBmt7DI8WpPJW
kv9pu4zf1gmewef7Gx6MFzILL/opc/bltfc57RuH5ClhyWTZJbx0jzCPGrdBRchn
4ev5KQ+YnuhAN2LWHYvZiIoq8EMHzhTktrCa8usFgKRla+JIcbjvasbqvmTP3ITq
Vd2yISWMX0XToV3VDWF3k+yhOjEymvm5oDy8jJe1k+Wk2bGLIInffMuziYZFtjU1
7Sdoy/243sJ9ZPFun0Bf/gwtM0pEtJDW9vEJMCHwQLC1qGQpi91c8/PCxb89dKXb
MBI+1wkIRTL/n+X+OPXomx6vWj9s/6KWsz2MvqH9ABaj/Rp11YCaWDUc4bJLd2t2
uEgj82V0eeNGouOk15rjCEEbc2xEbON5//sMNTC98i3ULryR4vPiJ9Dg1gVjEOld
qWOKK85x2faj4BEaEssZKQ890oeB49LNUyix4Dha89QdIDcHF6J2NXZHRbCvl9rm
8/wqRI1qSk8/UsW+sr5OjbFfoGzQ0jlWao1JktMZNwQuqOza72iEmQ3w5dfnl3n3
FCdBmN7iJCx7OzGspeeYPvPfMHF0w1ajWD5gLklVFd8A+9ZV+EIIlSUbNri/CwpR
Q1F62cGhRUw0sm9lDwtaxj2C13fEF5yKs8ITNl82uUjEdC+eQ0hQc/mxmY3LEkAl
Vx/4d+1kr42BpshR9ASzUmS2l3N9hB+quYb5YqvvD+M80dZhEETEc/6ycBwb/wFr
wr3oiEXp3ElVPxts6IBhpRKwiu2Vy2atkm1l91iZLvx1pY3LIFO3mJE29/3/05r8
NKYiwpZ4/M+dWa5ZSEmhL6r+g7jRTYA1V9FCSkJyiX+oIYLHVYEsY6TGHZxBO4rr
+po2lsXiqCSbl0PsC/tuo4d/B6QXavbo1ptK6x9CwZRpoWoeXLqXosgL3x2bLgxc
XGaEgkfqyWW+dplz6S7376pwp9F656H+M34X9+ZVZ8ixlojovkosMrSVbb1wP/BO
fQ8DkUZeBTKpybvRegfoq1lTJLW91RSqIQm3DzaUOXOsBdAUhlngA4TWODEyAq5d
iyv/uTDoDpN+Udmhmak4d5k3jOu7W+u9nz6paw4iGA3GJ8ksXAT4r2VRKdAbZszB
nRhSVbVHo+ZqrOQjMMMr35hfScyVqnJU2tpAv3HlrEKleYeQ+b8ptkfYHV9N4/7D
Kw6RhtTHWxpyJzIKU8R6mm1357Ej/LlDpirIKH5Iey2ZPvog7V9X3B2/8UVPXWH9
PY7e6zNroLjQkFnDdqiMH0rCga/BX/6OdJ+97ZjDjY5XeNPC71ddy5Fp7K9HEtLc
m3RzYzi4N7gPctR0aBYIRlpJTlwSAps4+OUf1n3odr7Kp0qxTwBk0iA3Nqr3W8o/
oLuGxaJeBSgQW5bwuhlYSO07yewGTk6UUti5vOCe08lttSrG8J0Wf5xEjugeRjML
hNr0phwpa0OwrFUil+zb7NU1iGByxzhhLj5nTgnoXEe61v6KP6nPEXVZ9lmjCjvh
7pUYPbgJUnkNvuuXX2/xN59EQ9SLcGKdMrEEmbpVkoIWoSeFMVrf8kWraBz6TRbk
l5zKC7ktko5H7AbJzeitS+q/LJt3gNTtwYWfBdz1Rw1RLJ7JIOcJHz+TmS8jfyzN
WfQIFowIP0/BNw4jrS8cnYeiUho37dMVr8R8PZWKY9n39lD70fZZcU84tfX7/Zjd
twro7KRQZrTBewUY2hbjy6GNUmLWcUxPJDhX4N6nfmHsi4aSLjT+SpIK/Axf3nL7
Rt07ccBLZ4n9JUAZiQb7VNmRThuMxCshaz6+yCEpHvBl7Ka1Y3IiOEYd7MuWKRgn
Vj+ZMTJOX/8IzoIepI1S/BTdtmOr9Q4VBDXZvAZ6RNupKWfOY0xNHYwKXXAjHCR+
+LLiJOGmlVRmtcBVpTci/5gmvbbSTYn/iifW57rbrbUcJKc4UUOYQEK7y3GZEPSo
+PIP4GJmcKBwhiRgORkpHz62Sy0vBAfFqQgplpc7VJjNmW112YAXE4Wo27vngfFx
2Hd915sjPsFlp16VnMnExEHgx7lwF7fWzIJXnrcooxER7Vo8mNRjwzODahfZnHHQ
n2j5HQa+9tePM65OkqtCOHYMh2W29JxoizdHUzAeC0eA8OnzEXhgYKPNNFuiqJ9p
uGT9yTvTiDPX/BoNThAgf24Wc688fP5WpfBFNB4OEzKLX4/gi7zUX99grO7tf0Rk
JVKGNb6W8RCb+1A/BAptykaWOfz/udcwM6vX5iiJbt20YJGCFoklqzDMTfSEJ3oc
nP3I+gaZVgi8pOInSSPsgvds8GrKrUtEQJHG0vRfKxCXYBUiqHrWqnovBdSwv12+
Rvx4/EYwsoZxIqxhF6Am8sCXWiXUcbjuYeW1+heWMjSQXqJxGox7rZuvdSJc6PgJ
b6ooFYapJx1vmTTolJkaXZJR/uV2sIFEUQf/tlXesSZxT0Ymoc9uQz+rTx2S1RYz
LNLUxd89EDF6/o5cpdKw/o5vWDg9orF37sTjDsxbAPlKl32nwDYnAXTqHA813jUD
r37nnDokm6Rt0wgNqQ9TaWY5raftp0Wje0uDh59twUIoItnLsUGirvkYXKNezDSm
gB6n6Y4TJfXXZu8forwPDfwQHQ/EtR+8n78Vg5mSElkEg8wh183WmKcBEy/36eIM
1rokv6ETNRx7regxYdCig+KMXDyqrD7D/PwV0NNYlKmo4FvafvCQpAHGHqM30GyG
op9KEWpa/FekLq+2WxJx2vZ2Zp2nFM42o0hpVtjI+VqPyT1s6yDEs+iR+9uISDvm
qgJyc/+31dQOikj3twPpYN2W1W1TzYk/UAuJZhV4Jh9Zl/CBMOB9+NQX/kk7W6Zs
cFll+G14kpfimi0XxfTyXUsM9wKPZ5Veu/UWMVnxK2njN2LBui6Eua3AyvMhzxKw
4sCKTaeamEKGV+b2+q5nilXXd9IrVR9ssupYIiNZt0B/CWB3ofHSrbf/SnGFC9oW
7/0z0mUlOG3nv3fOJakmhjjM52W9rAdn2auhowk+dw+SW09hxtmLQckbBccCmGfh
Cmm6e8+1izHhqypQudjYbBnKqpcSa48zO1JY1MQkuVzq8mZfe1CU4aH5SLeQwrX7
KJ5PnC4QJ/RIfPRegkgJm+dVfN1KZwT/s1xXaGinUQsTzkWf39A0msUC6VAQNXC7
ljm16yjClhQerxy7zFzqiJFxJ6bMlhyGQKPgTtkj0orpv4zbBWYnCoMOSFSoN2a/
GxtELKpEBOwK9DsohQSwUQllWH+SKR4z+6U84IE7Wv7xCpF79uxsypBTtYkmtc2o
DWCaY0Qbl6OWM5M55GdsxfU3h0Gpc4oZuD1R/yF/yRjM6A44DKUZ2vU3GMsdsQ6v
tJfZo8BZhjqfn6ZA4Fjg80C7pl1wVK0Ke+7jb7RCcbiCzOBkyVVrVBvQYwpjo4+M
4cdqKHiKmM79qI7idb/V1ifk/qHNraiGV4KVdImupPe/EhMMDHiXo+pjiwS2rbzN
/VvT7vwPxNLteFKn7DOVm6IzkgtZIJldXl7MPH9sezi1wqulY5k2AeUsdYgQe/bN
0vf57zr70Z5MZ22HJVOZ2h+vYVHGkSaelQPdK4s4KMSk4bMLnn5eUXPnysG4haFL
i5WOhZKEvQiLP3etvFERhR09riAgfdAs8JW9DVthcbVr9HuWMwg5OXUS3HIu5VKl
IPNGSweJKKQLkojZ/zujF6h+z9BZs9y9gJSaOSc7O+6a31p3Zgu+b6sfUd6REjHi
mo+m6AfFA7m12eFq9GbBFk4qrkM/s7KgRNg5C0DOWsWA3urNnlstM9eTjPQCFHTE
62Q4jJNbHcCzqhfo1nsGKk75q4J2enH7QIYmw8ADds8BBzNKjlcOhl4sPG7TfcPP
Wqx+Le/8KMLXfPYWKDrrf24bbvirG79VX2j4BGuliJeMNjYx8d+5IXScE5fl1NU9
O0KyMRn5kamxo0t52ZwXu5p1wUMMtH80FnAwhrPNI3OV8SKgeMjh0yqr5WhgwmCW
BgMPu/GP8opuyxwkC1xkFaOIRe+569L2bzz/hIslM2EmqmHFjC/iKE56/KNHGCKr
0oQ0J8oK6iEXSW74chxvcDbiVw40E0l5XHP5Yt4oX0zee2Mwp6iSLgyPTgpf3YYx
DoF/DM4XTQEkyuAS1X/zGIkaPvB903CfPI0HXgpyzDScayFmNMcd3MszMwAinleh
6j9cW26exylIn1DipXLbAd6c/YUbRfmROPRAiTUiJaar1Kf7Kef0iQ4dCBpId//x
E0uPA3+7fFKH+qXJ1vzNA0WOSl8zVOfORj9wlvFTDnkYAsQJ2VYC8sC97sIgl/lq
YlZhstUFM+tEIOIAN8XvE6Xdp6dNPU+UCPlhNSXw0UNRpdMJ18TXXv4yDJ2z3KRc
9BVfZgnXTweXV+86xVzEGp97M0/ZpLGcCIW1G9cBdIik09qYuK2eo6uGVEanZmI4
euDJrVd2SCbL5svX61cMLjbFqoIVMZWupgjG6IQlG4ofB4EJZ48544G5f2wrxUwu
C6NcAF5CVSMQaG3oquKBVStFLLEu/NVvUhqyl0ZBb2a9A4JUrDtEyDsBQQ4Em//6
qZkPaFbLUGRI1xn5ZVbPjru3fTF0m8/u8XM4p7DhDqvJCAy8ABmZrXhugpouQvPy
oqDmq6tV42vF6ayltAYIfE8zu/claDkMPHs0pNQasBc7nHeQ4I/UvisPLBNjyn+n
5tMGLgHy6+b9Kd87Ct1ru46ZE3UEmQb3Ro9sw1JV3ZLaUb8Ku/UhPAxFmU1K46z8
u/4k06sQsQp9tbW8GFHQ9GNtRidPFXQneg2pO5ZcAJL0IGYt4d5E3a3fyq4x5koy
vegsKfNPx6TqNykxoAV7wo+RQStjK2BbQINFkcGgboLayK4ZuhJ+ufqbKgp/s06r
e1/FfdbfFbwztBDkYUATw1KfffNlbYeCpZpa4E3xkY7D28PW/VrSX7x9hqCQKyQC
znylKfNu9P31HyQPxXXHrCYrq01P6hU41UyXnf/3JTPfTC4Id8hLCuD6YTwkomyE
koaECtU5YDSZoLnPS3QHmXe54OjJH95Opg4GaMmZV1/tnu+OW3qat8zFJp6f1jv7
t8xbPL/wloopa2+jNuxXfqqKpgIn882X4SBcGWbHCM4k5Y11BY0FISyJyVQ1ovKx
7GlvU5w2+tWUU97DghoBGmb9AqPRn/x7lyf4JersTNtVhn1AoWhdXt6ye3HKgOTK
I6Vh+y7jeHRkF9GMtC6OqUoPdFuXUUjiLW7/8O9X+jA6IujMbUeuq0B21SE7OpKD
GuZrIkE446mJF/vgZgRpZ9yNkPXq7STaR0brAK0w4vx2660SQszP0XtyXELt133Y
vJ29XVCcCObAav/2r/J/SW3KBbBPzyixQ3kPWsUeckuUQxJBxvQVY2XCnhCB+52W
dvKs8Z2bvLZ8kvIKMzX8+O+bAkdSvwyhIYO6awmBnkhkKftHlTSdImZjBSTRNaBk
iN6uCAqZDOFUzRYn7b+yJoFcKo2VTptD/iPyyptGFuANHQ8hzRZLKtPew1UHF32j
5VbsksZXzF4Cf6HVwGbcN3q96J4KOc0dskQImy6dLXF1lLjnVwlwcP4/riYGE58/
mSbpMoMwVhIULPBBGDLziXvmubTV4IBHuPbGcSPo+bfmC6OKfSYuz6CEUIWpsQMl
rZUdkwZ0yMku8DQpiGvFRulrn9Gs8vBxjjDVR26otaHy/XCgfdBIFQB5r5VqDmEI
EGUd4uflQEMmq/rWRtSQMMQ30AZLdL4FQYUzGd0kMiwX2kwkDH1uaiUqbFg7K0c+
eHCT753p8+7M1yNR6c6Z8Ul/paYArmGUmUQfzcNXb4eeW6QVgsirEp7l/biO7D8b
caT+Y4MZHfmnMjgfR2cREEDwr245qT4fiSnqp2+GUtQph9kM08Pikg3nNgRU7OdR
rFNb6be1IBSofL83Zet2VcX/N9yYZzqeEUL/kxmMqOCTbDtf8QaYpo4+Yt9Ro/XR
7H+iGUh7qBV9oX55cnbx6KBnEoMcpxwY0j8UkvWz690PPRVkAJEqO9xtFvBqgv7+
dG+h9Rpzya0+qTnCD8+gHKXdIps15B+kzN58xyBnrfSF+wrvrUBPAK9h17C5/7ih
q4Gk0V9Nq6Z4X7w3vVMjh00rqHnUzpVwku3XDgK82MEoBdpVoGzoRja1ZmpIuUuN
LWFkDj3WoTIHEmETqbbomM9VmJYw4X2nfSt8arSupYYGpnzLzZYHl2hrJInuv6SV
gicYAWW3GeEnWyFkhGH+vuzcbhxWsfNtIE8/wjv2B+Nc2LBoENgfEPT/zvMJEhgD
5yEC90qnr0OzOjQcBQj/4QABwyAA+xwHqzDLamoU4fNV6KsqiHYveELgoa70kX2S
nI6zn7kbycf6BorITzCOALOFQjbuPfIAouMI8k9Tvd1RKZ6aZ+UpG6Yy8dkaFUbv
xjNDke5VocnD2SIF428aKGixaSeIhwuE5dDP486udHzjv4giQdR3GhBfQvHXl/Zf
DCR59rRRH0pvA8uOEWtjZgyw2FiKY11FbJLOf40wEfeMba4qGUeut66oO5a77JxD
6o/CIzD1L6qSXtvcQ8r2UB0AxEObY1PeE+Dff+z/HEOfnT16+x3J6RM6+vjFg4HG
bPh6UBBFkE1DGMBOzCKJJPi5XTzeVqim809v2EppBnOJympeZSlacArbyEAeT6el
46Bu+g8ceZkR6MepALWiaQkqmBrVU4spBqZnFFYUzwCZk05LrWZmUrJtfy3wWcOq
u7tg1etf5JVAIJTQB4Luu2u/UHJACCzcpw7nw9vUQDsLgEkjrGzOvm2ig0+O3JQ6
knFfP3POFgakXgLPIqMuNuQLx9qJOZd5sDjP4pvdu9B/uvQ5Rv6dYY/+Ztp1SBcJ
kyd0cdEP9W7BaSLPNAZtZFqZNaTQZjhKJNbauNEWBrUdCHbL7unh7ukKcLma+sQA
qJs/m2sBXwmLDt0tggpvha7O94vrb2oEafK5ANph2sivx0dVwDnASh6zMykYRWGz
SFy0EJE416i5EDNVeV+Bcqcs5vbqANcU3fuj24YJxgwp9rHD2xrgqR+m2XZfd8L/
Ztx3jPAb2E6PXkmi1J1lXnvqr4ybi6BPM2ra6n6EYUi5e6x6b/B/qHzZ5qcfQmjb
eT1vsJozLsFuACiJXbZoP3tfQisocgn3d1pmNhD+7rmVswXrEmKokhtd5scCWHlV
U/YZ5vWQ0LOA6fSV3gbUUcPGf4pbptuH1RVZRKnFP8/E/AdCuQeeUXMCGQTQkD9v
qMP+py4nzzlISymiZkyrhBTYpU+Y2SCfm1PkOyGO3UWeaWXTkwR8QSqrep/PuhPq
N62MbOqIsnW7RMoKvJZ40X7AcieHsAynA821hV0pP8CaHeL27Y+hXJjx8CMCthCe
TMy4CPorfwv8yZxNCvSii0B99lJooZP8FxkBRiDqDtTcFNsrtfPTYBcGLQrd9cfj
iDFLInUuH9tiZY6XWZfuML/NjuzohqPe3+eSWZlt0j5U9gtQkA8GKf9NFa8tG1ww
cijmvXL+TcVpIA+OQvQqfI14cbBXjZHa+ILmCq/D9VmPUGtqp5KjUedRcsBgHGWe
q/RbkmZy3zWWGQbWUom047HAsukGwLY03eeLGLz+ApK+AP+8gqEX/BZLQlD44zlz
21QD8XZ8sDj0gzP1Rx2SZyVKL5CfcP6+h3i0jBLJyVIxM7muoKiXG0LnKLBhNanF
2AF9k5vAfk9CvLTSffX6QzJHs1J6k5ofQUXXj3PjO1aLcD09aB5McUt6nQfSAxNI
l/mzfDESF1HiYmdYmgJbxTaPIq60TncHMo4rqUQlsIfRx9lOlbVOk++10sjACGkb
WAks5MEoNRixEbl2ef3YvO52dITdnPbBRhcRXM1oJ+KpvKjXpPjbaX2iLZLJZ4OG
2iD+cyuRhIRp854sfrqfgUPDOr0oWZygk/ifhGTLm83SWV1M2UH37LuxXJFtpZmg
5fs9nhjD0kuW2NiSahwb+1oUNrJlirNCwv+TmkLq1hyLdLXLR2RP4z6sOE02AgP/
MBvUf8KAe/KWQcy5X9pldKLp/4uEDGeFVbIl/upca8dQZ97e+7RbCrzkRZcjcCy5
c2zYCKLLKUgfJYg65v2H8sddGclEr2iC0LgbDBYh6dVJcY5qvfz7Xmn0nffmOT1y
xf6UzrirjORovCBsUhL0Ys+fZsPyANorIdyBeJWp5xRamioaAXlPhwU2MsX5Qeap
FnKx8TT8ZN196wI+hLj2hPMx1GK2jT+bL1VyoSnpJMURyN32GtXJHLqJZUy5k5nn
G/505vKIp2DrlWgx4s3hIlFe3H5NO7J4wig3SN5N3uj8BTG7EFbuIlxsFda0PgnC
I/nGjUORM3sh1qvyeYn1WwoFPI+C6giNixvWM+vkACip98sspRwq4P6McVOZYMON
QQsvU6XMYJypKg+1G420dslEqXe02/rQ/8rEqKUlwfZQHW3sj3CDLR3PGcR08f92
Eeb5xd5Hw2f/TNd6vzLmXEqQhLcVpFRrw2GJCRbjgcDnIfwBsK2Z5tBQlnb1tSUA
h5eQmgWkMQ3bPYUxcS3CcICy95kqnJeXpUgA1uI662OO4opT/367VoyFJoZTA8oW
xZmWKg5K1YoweJBA5pIgvaXrhLwDiHQX5mbOzcp5NZPhFxU1+g0KiuTKkQ1ewobd
OvQalhXt4gSR1tN2SOqtJGvZp8nZgclot0tSficlMGgXz+g0v3VBc+fC9f0wlPMC
m+MxVi/NLvPryo7ZI2lVsAZdc6FtBi5X/hRKlOW5taPDdJf0mLwEyGcsP1XrcCtr
B8yvQzc4k/4AYHlyVYVUngmqhxAzeUT4HTox5yzZwXKMqq0IDMvO5MXbVsUvmg7b
kC824es4ZcBARRQ8OYR9R5DmKXyysxsaxkXFI0SQQfHJ7CPJLgMbpv4R5ZVZKvOg
8kINj3o4X9u548QE9M6lieL4T5HqJmm6YyBu+oAcGwU/Y/+aKcCzRk1ZTTu3LcU3
fIjV6udGDfMYET8RBMjr7oSlPF+MbYrIFL5jlBvQstxvcLuN1gYLIsoXoCj9qfFz
ncUuySs8JJjvqeWBW3j/4QvRJYGXoIZzKhi+Gwq4FM/yphKh+gfAo+SBMgHZAo4x
leQ8t37RWNfHSyNuPwQ35fYM2ZA+hABHToW2nvJEy0G4a/HOrZvfLaECtE+fR+9j
dFX3c1cSKtOPTYhPidEUDIjHquBDLM69bpPssuIwO17GDgD5zmPIlSwxlLcba++o
hEEDCSYMzR8Tzwfize7ESxsG8LzqutU+A7KznwEbB9DQa0+NfnhBRCfqJ6STOJOs
Au3RgecOKCWBzkmZ3XFk5j8gkflNFEx/z51FFA0OT5lUwKO3eH8JkQ3Gznsx8fDS
+AAmeA7ET2vSFp97zOYUoe5cTTLtaxZSN492ag34jt1dwxbDG+UNXsOfubHMNkUl
Bs22vIxR6qmzCtGH6oKhlviL7VytkPTjh79BTqxjIYDKdMY9/y2BLhVBiEbKIJMe
hn99TMGcrtjqXEgmSZWv8yqExBizFD76u+UJqMw9t9MLbd4XhpxIp5woFBpBWFr+
QmK41NKZQZDB6m4BJiGZQ9t0VX2W7hccdxMdywcDIteG0Xpv8VlpaWG/uEVQDxh6
upqOauvsxpdnbITVX8tSuRRQPqkTbDAaThqb3+Oto7u9Ic/WeuFXKR5U/TWQgV+K
RqLIDgREg+AHjFXkWKLSvX6ndftgTQTaYi2JMM3LmQpo8CCmDxzM19J8FKoEDvH/
RarD9F4Y1mSTP0huPrxkHusamFWEaoujmxR8ibSPHda9sUbPiYqo6jwJ9UnjDTBL
3jHZ9HmpRY/Buh9IUIZuvAPBG3Nz+GsHZBnsogMHFbQaWYqP2BHVACq67KgYjBQc
Eu3B9QW2oVnPyZhrHzmw3CF6LRSTS/HD1vmMJe62JXon0O815v7yvVagL92z4DfA
BVMCJTn/N9H8FPSHS/KapFk/hqOAqIwfG8xfPs9gnG+fVh0+6Ii6b6KbS9ZCMbhU
nKjvZwAUifFuRetvb2jH9pWhqax9NdqMV/Y+eWff1LboLIpGNkxGVa4OxJeZv8vh
jz/PHDMLVLMZD1P5XgzPPzSQNSBwzsdZwAi36genSLgb0LT556JJ/OFstpPaWTAN
llqSMs6mGmHFuYysCQe+T8GHht9haf06/9fPIDUMsJ8zzJl343S8/DC8ZDGNBMgz
BGgSX5zsKxWH45HnHXwlAkGy+8PNEI8Q2UitzmcI3fTwzv0hpIacFmSSqbMI2u5l
8yU7MH1b5wCAyWNFy4B/OIIeBEUQZIvMWwEZBuJIZNZc4zh1JhtVB/QhZq5O15AK
82rBaZ24zqJMXnpBDBjpj0rTZ2sjq9dyT4IMIsEnYc5qnXdmZ7FLAnLYypJ5SEVu
PZrtxQP29HQKrv1YLFPAmZuUpRQAlGh2TrgcsrzocYe8tboytQWB2iqalJBHNey/
VqOuFRK0IiG/oT4ohWaKfIUaU5don5kM9q8LU8g+pMT29wd1ksotDXYW1bO99Iwq
IfF52Ouhl8RusoyEOZ5DSAWxO6UuG7XyqZQ0oG81DRDqYbglIln8FKfzE40Evby8
NudcmQKXxrJf2QogAuoMVjskUfuhHfcPpXx9M+NExKW8ZlFpgCut7VSMCdZEYRB1
jid2YXZ8tOFHYrcdNUtcvCOLl52seBpVJxwCUJoQ5LbLgtlvK12FvLNjKS0S4K6n
i/euzOY7QwTR4+lKfn7MwW1awfydTv91gp9ARhWixI1ZMmDoMS76p2z9Twk/js8w
ixgMRvUwiKL8NZqm76PXDy7modO7D+Ckf1nFTk//h7FERGdCy80BB6K3PVLKWxvP
fBzrw+cXlLVT5LDBDCEHCt86MhSVb/+/9BULQZ8Hthi5ArOXl1HWkizKezvVyZWX
AUa+ex7RYA5Ptt7s8208Pv8RoCqfxzw3u6Sin0AYkcYSKUbyicYZrP6jJ8N7tyvr
eiduoxUd3g65QvhoRZb56sjZ997JK53I1qCrJihBkwxVG6w16GNS7RiVYiuUzdqN
U14JQuYXkKvOIkwdd+Nq9CFDBkAhjiX1J2Had+huLn3MImC8fMFgg296mrixrtbj
y2xNs0d3xF0EiB6PMbkduacMKwp/sAmOxyGmXdrGCc4NWxrFhKUHJTJ+jnau6iZg
Ob+1zueQ0n24s+RziV5H5Z4HIof2hPSfNxwEEliWDM4B48kBVCd4GcTUgAQBWTzC
9aOKmfkgt4IL/a/9ARkqcxIrYKkfcwm4TKaab4V801VUSfAiAzxG84i6K1HAzzYe
MSumpr2aB6MODXUykHp+G+r1b9OHCC0TeSUixL7fGbzDKtibZeJs6ZU7zoXimynV
OFSxvxN5a7pYCEpmlmejtS0aDI4u75tWW/XMWp80VhsREpkbdhRrsiotnLppRxtJ
KTSgJjyYsmwxSTLM9GbYzqpduIthaIQnR6MOsgOaTjh5lQ+tJRD9gTFV3pSFFJcZ
c2S0EIIJRBc9Ks4lq7b3eGAn06tpVPtdD+053niiEkWy7/281KFw4YapIiLXpHcf
Xmjc8bYcCSJkMylCZyc3XZEhNSVpkbWJIxREBzX9TYPqLRDfNSCnIv5oQG/CaUNm
7L4auKCOWEo6gbXSv2MwGkb/S27PUtCkqarVV0+DDgNToZ7GztFHvrAxvLu+/1T+
EgWYYIpY2vYGr0sRRthhrXTp1uPlPXlqeR//Sd/512J5H6gzJZrhr8zxtUjDQGHt
e7OwAo/lnjLDigZcEoMP6bYhN/Q0woM305EDBkXxbXpOFhyNrKC6fdN8BeV8eqY9
Npr+km5hwWmjbiJlRjOdYkcbucIWKRGhaKwh1r7V5rv5J4EUcuEXwEZENcGPLV1Q
5dnn3D/V6zkZs/J2B0rAtE6j7o4OWsHeQpYS3sbzBK+EUqmWlZtMNYXZW0xn6kM3
/kroveWnFFg6NeSs10/DPbwfQG6oxLCcynk5putS1rEUW+JTabCJIyuL/rjtOPjN
RvFV5+7Qr/pR8thMMMMAmkC+2+QtCiZMPTIViFmrJfuZXZhIFFXJq9KF8AeYiAL/
LMpPFOO/W525hhM9UoVSQUTGuNBuF6kI2RebSflY1+1SA3TtzoQPX0DVbE0TvcOu
UTw3WcaI1duEgnRF/9Fxk8EFE9+HkHjybNuBgz4xD7OmfP+KLmfz8nbPqX+KAvub
xUL2+zHhvW9oixPgncW7hOIjztZkrDbV9pk9OYlj03lsBShbYKqaPn6FFfp7u9F+
U8dI6JoxfHdw3o/C5cPO4Zr5Q88e2VIxvfW/9r6OSN30fqSDo0nX5DoPDYGJZ/z/
7aB7fS6W0AdeUsxI6hal1o0OXUBRcLBIKwMhG2BGbRf69KRlLaezy/j07RpiO39g
Ac4YXhOrIvKiX8LfKZ0enXV6/UpvcTJVSW8V1TIV4mjDw3lNs51zNsuAFX2je7K1
GVLJM0Uq3s+VVpzrhNIATsU7tdxqnkZT34dydMD9z6+x3Z482K7OLnRTNZgwHJHo
uD2+oc5pi+gLEPchk4kPye7vWtRKEP57M3wIscYcy+Xiv5oEBDs7qhZ06BahyZi0
Y2xZkd35Dt28G+yc74yx3dVk7Oy0EOcZIPDcckhVB9ne2rNxTrJXgMT0xqkFHLne
ZNfW4I7h/U/NTrzzuzSn8bnAX4sOLR2QcSgx/EM+3lRUYZ+kFLb+60ERfKs5/zrT
zVZottNXpcqG84KkdjyrROA5EEpqq2Byd0Ry7/t1u0Ds5myiZI/JROdGtOBnPJEU
Tne3tsm2Ttt8mEswzqlp2ngfRFiBPiSIJRxAzGnD3FUyZmGpy3+lawK7lLxL1Xh3
QqO8HRBEHRv5cgIkodaJ8QNWMEZZOGWwtUTFUuWEoVWqQFKOewy5wvbDTec69Uu9
tfkmCf5BotNGG/n1eXpPsblYoe+AeQe2toX7w1D/ieaX4L98az2jLXWnBVxSagBu
0Vp68Ekfzv8/lGs08lYaGsDUKieAaGBgBUFV76xnyLEXZS3c8yAcEntlb31n/kkc
KHz3Dmdh7REdu1cwqb8nj6vyPo9wTCyHz94UO6IZS68w9TxaoIcVmpH4SZXuu2kw
ANAecyIVPt1FfZtRCYduq2/5klmWH4aWGM8h5y2rDAGAS+wdV+hOA+pL/1kNJbW6
4KCwoQ4XnBBx1XyP7n05QxRgJ4bwe7uCtR58tkk8aonO+XtGuvrJTcm8BTFulRz8
cw83gSHr43sLLmPrNp0OUea5OETgwbpW7prl2/NcxkdNk63qgvhBl09jfDS135a+
7FPLooyGiJ+kS2nT8annssy1UIzhVjwqbocn2I0v6xn2EGawbqZCpNQoIg42NxlS
CNnVvq2waYqFbtje8ANYygJcdiXyXgAq44a8VLuOsuBC0yZKQzemAmQh9S1k8Lzm
PpgeZ3X1lKImf34m1L/z4kq1I88dtzzuROB69Vp+3XM8SOGCGVGzhgmKo/FiACWm
VVsZ/vn3CU0wh8ISF3U/ohraK1U1fqyc8CiActZ+iN6vXUSLMMY8QcFPcDpgCz4V
I0UAZjxj/WXXXmuwj4ZF5yvKb7DwmdFnVsRY/67oy37I1vfRKzB+GfC1MVNGgtWu
Ay0pKf7fIwOZlw0qJYzsROizw/AGDIR5RgukqkAvW3j8isfDlX+y6weY8VnkELha
E8gFn6nJQ56FlWCz7C6YAqunViX0rXHsv0wsGsQbuleSF3N8nqYxGDJ2EV+kev6m
b+i7lnzKU/nUq3vxfZPXOxH/eBNF2vSBqIHFFzeEf4yaA5Ap5m3loZ0bICMvzDmt
Gu5TaOQG/Zb/gsKAtTDUMhTzESz+6TIwQkvVZxztgmSL7PP/mjAcXbXaiuK7GPML
aeYUE8wsxKDvRLM3usSdyx6c3t16kVzlp54PzZ3fqUwz6FzGOam7j4Z3t4gRHfJk
jA4lGVmyVUemHmVPCAhBV47iErhjkOS47Su33c6qTrIlC/foyLcjEzOpQN6yKRHm
Had1KnCaroL1pLfdPadOtVHL5wI5u0E6yNHvDMHH1AiFifv3/yOpqO7qEOdQHsZd
mLke8s1DW2kcUmYh7v2N3BByJ9zJrjMROzO8YOseatjPp84xF/BStNCPqXvZQEHU
AZBqHdmlkQlN+LjLzUrY6awQD706u2tkNmbECwrWFNN7bPQVVZTJ7H7Aaimuhw36
oaxXKy+vjP97YXMbfzsKMsCzdBDkMoRRJvUfKZcpYYSplMAT4NjmPgW1E25P/9iC
ddN2rkBVjE9t466bPftMeFVeH0uzlDV+GYcnzqoJnv9QQ/zmSJDp44HEdrwJxu2U
cn1VUbfe1sJeQrzqFXuhmdg3b6S4EhgGS8bQr4euDwoiTAVXFPKvvEv9JC39szgu
NhLpmIXeVKcqM/1Ewz8bGvnuUCW4dxpg9MBH0pmXQt+E+gN15hk0SrZB4sfwHgy3
b3tSYzF9TzpPnM8EDiJZXxgkQFzmUfrll7rJhj5oV23tNWN9hhiRaoQ0SP+1xTPm
ZYPcjNcrFTFsBG/ZCtMMpbwzYleTWyW8Bt79tuIzcd9t5RKtEyJZ4ms9lv3xogbr
uN5zcF/iMWHa/5Z5mHQIkimdACGkm99Q9aNWidMg9HnFepUaUQS1eFSDwWi+vpq0
+4X4WSB/oWCBb4fVizNTV1I85/DAXb0CwwTsXqH9BXfMTfj1xACQgu7mcgW3/JTv
a1zkvYNIVtKkADPHUvqwsL+5dk8NoVERXk89Mnz5tLQVwPxtTWHTHSd1nhkPqxb4
bdw0SzRZjOKDG0+JzEQi+BnEAW8BaNW+CW9MyJylVcYmOQ6vps12xTOWiPqPJI8g
tIzjvDNLeiyW7FZ6Fky+85Gija5BcTXoZH5iXI32V5sOvFv1IrhkahK/AflEerx4
UwYsvkNEKzzi3UAKqOLvqLqmDDknj2DVWGlhvZQpOOv8rpJ+XEy2Ln+cdLBxpVeR
etk7fJby2pPHvZhBbdtVlj930PqU6MRRlUlCrsLgLSv0+HoL6BNL2Pxn14K5HwFb
d4fGs0L2V5dPwN1NbS7JPw9OX2OnLQB2nwKQst5KAh5aOE3t4g2+XoqB2cCSVxqC
CqxmecYRbMUQT+bSGLhj0OvRrQ9eMvh+Fg1WUyPvIT/dTKGnUdfmwPaQFq1Xix4B
uxTcF4v0y2/m2xjikkQM17P/fvO11gtUfy9Ck272qtxyAsF4BQEiRUClGpBioctI
1quwjB5CaxbNjUi3SmaI20javvEY7qS2Q0xHt73PQC5SjHlS8efRBnUboRM3vJja
Vu/ZiWDuNDWbQa2w/Aj400BTdfeDwlDHVmmqnoI/88ETWTNhPQ5LwIi3NYK3x9Sj
qmD67X2Be6NwDnguRfEk8DyvccggrGjV7sQlrfzzfiCM3QTvfaVooHSxNxasD8h8
25YAHlMbLQq05crz+sDy2qexNZAvTcwzpfKHfScZNesvnUymWHQ5uayQkRoDbypi
UyekR60jNxuizN262/W2heK3hWbRUyqfrmKEmOGw6D+UhjWLL6Fp/8yTQVDoXGSO
bWCuGI3TgEE+vyq83B+nvmxDrAvu5Ca52X6r+G2FN//8EM7NgzPUpJoYdqbIH74D
KSWfES+/30/96doiubjlpV/BpwpZdGDj42Ipz62PJzOZ7FaKkkjkGtJpo/On8Zh5
Si/5z0O8lFoTxRFeLYCImxcvbvcOvUSqSyzZ8MFPVfRh4qmPNCo0eK+2e2nDOrUY
/neI36iQYY25/kHUqbLC0hHsLze0VjTP54qWEM6nU3qWIsFs0D4sCNq2sxioMcVy
PMKcpjAzOm1Uehmby5Orda3G8ZkZOabIvpDlzveSbrNrnJOKDbXy8cYSLVovFqp/
+Wkk4DbKfND6q5emnPjJtctivxEnIobSO068HPd0nUUuqzpkMgmPMhlEfFmZ1vRK
YsxA4r4vogJ/E1n+mmgQkt116S7dSkPktfqPPRiIclZJ79BYkHOiVMv51sc3iyFY
krQTiKPxRr34Ivb4IvBL93rRbv02ns2H1BzgQc/qmn/GlQyyB8FJhXz6vZRZ8SjK
BXh6a5CcFoNqvpO7tSNpC2qm1xF/1HEwgH8vfWzOJYDtfxWfBtDgD7kysAlzpc2k
2jqU4DYO2hsfdJqd84WmCqgXfsuhk28sHvGTcsfvuOwFx0ph4gnnn2mkFeZvxnMB
1ZDN60TT/Kp8AQdWhZvL1h8prWfp+L+G0XNbVXYuSci6Lw/X/KOW32b/TRO/I0Eo
sHX5RDmCerFFF8v3tSNJbS4lr9P6z5sStkFyQ4T1uXWhwihPsx5vEL1efPyNBR/K
xEdZG8pnwShzQU3HnJSqy1399iIKMZvVIQP/izKg5pNwxK+SmbLE9t7siL1FoTDg
cdIzFAlUdaXLCODi4JKwtbqI1EgCFO/bEjIFaZdZGJniSOuLOLuwbuQMGGC2YTPZ
AgvgH3e4q7Fb1tkeiTBAeHhCOC09ErvMrFly0QyaWgGIApe1mHVeADXorHkj2IlJ
yf4jspCwpydbZ1tIxLjPIH5kgRuGU0sF1nkgeZ4BHuEyApSjB2NathmWrwVW72Eb
qeXnpFS6h79P8o+1RD+uV4XzW3PR36gnH6x5psTTCZ+KEg6Lboh01y5k8zFH6YsE
qNiBtZAbGtqwkWcBIrxwP34gjY/nhuh6J4K0zO6YFWP1BmA63QF13M09dR/EX2zf
EStqfD8VUqdMnfnK1XvP2XHjw6Cj5xovKUxP7xnqxmuowHJF0+mC6YMj4/QzO7Ii
EJNhT2iin4uVmNauH41QgT09xe1LN8rgdxRfpVc3dYNCRslSJdrObaXEdmO9T6Qe
bL1CE/aGYjpZAjeCohkxZXZLYNK3ZbhM80lSOX4Klnf1q4hiw+DQgYTZ/zY4Rhm4
rkuzUyHZYM4d/AUk11va0rwRPl2Gec3Ip9E0hicfTsh7O+kBgCCky9rsLfa1Jtpo
Mq7Zs108X4422NAPpDlhMnjM3g5M98ZL/Wa7YjbF51iE7PRArk4c1giwBTxd8sJZ
uyY6XOYOtZzVYsQpGaGv05fjTAh9/pzb7EATTai2XQ6jgp22QWIus8pPOAZTLZbw
aFKAsnBMCWGEiGdVBazBKY1NR3wj0AWmjLiy1iuV1gWPeNX2mf/rvSLdbTxqvjja
NyUc894K3mfjMn90sQhHpRYP154DKF9RbuD9E8agN1+Z8HQFfAbBbJ4scj1aHPm7
YVHaRaXIBGcAQsm6BxHizv93BEKX4pe6euYsfnasmm504HOG+WwbkGbZtbobyONk
AKsBKUDkKKRzHP6A5F9k/5jiGsKMvC2iMkwG5mWyS5KcRid5ZDXN3Iejmr1LkeJH
CWfpm2amPFmobA5t4tuaz1TDmtVdni/DykUnRqaDHhWEIeO3GD2Y6Y6eF/1Plosx
LmvULdWZYOUcKN46Ik8ztkHkfnu0aPgF8J+6aWoEW0cjxiqBK5gUvIkuFQBV1YwZ
855FzcDipQRYkKR7oX/P37uDPgqGx7Jjp41ljWX4ILzle573y7nhltfw4fBDuHKt
38K2wpnRtmGUMPQloBd3N+JvpSLVjcDlK98VOa4F+v/2ojGIfvs5bv5ygu39UXYa
fOo1q0fNe1UCuI2dBrjRKfmgqH5JFAJrXRLf7FzJFdcJVm8a6FEwyZwkoji4FimA
gqNWjZMBI0yDep+h2g79lfeaHo2Cfwge2EZ6402Do0H6MGjmQJIgRJEP6AGXyj84
quriCT4C5B2QPLzHmS8eftc0MUbrbmwFn6KzzMA9iULdvZeeHWj9P2tOWTiGbx7c
FcI2fOrtiV2KXr2J4fkry6d+2jzfDHLj5lZfzHOKBlRx5woaUi4wsApwEWSrDkf9
8JdV8XTbKV0pASr1LiuMLEJnTSczBgT5nzv0hIXryE1MiNzURdfezK5cNj+koQ2I
rCdsdesUgX2dPaXWwHyreFPya3bsmrLsGl7dWJn3eKU0oSMnCr9cAgbBFVd27/rq
tGd0msil93TsjwAOR3ciqBloSJjo37U6xnDBDB2OptGe4uYP2HpagjxJai3Um3zx
CdpvrUINzWsTZmVT1wm3SbkxvlZsm9aa+kcIRJSPtKsjYhaRYQhy+hYisu3EKEAV
MdDFQ5LrN79dN9bx69gaeGAljlpY7KSktrlsRRusq+Ln8ZMHLg4vS4JGXcrFNLMc
sR1+EInC50nvYi/W9e8ZHnJpg5W5gzcGOG6roaAW1pGbJDv374N2RzvKlcgr54eo
3LOjHMdL/6xuVPwpeEVROnFnTKnZ2z+sz/EBwtzqVw45uFzjqO9e7qN2f4SFZJGd
jhZce1zmUT30BaH154V3j9cpGEadi6lWmwOePeWbQAQLn8tn+Pg3o3ov40YOy+B+
+a5e18lhA2TvLTDXmi9dZNb2TM6WNIjs1PLIe3Z/lNSORYPoWZOfTncnQvhfJxqO
m3b2uZf3opvIqhn4mEq2G/KtJQTetIFycF/Z7ZVhU245+8FJ8hbK1OpHBAN0cF4E
soqcYmia3M6rFihy1Qdr6ToNQmyn07Xip8vrc7yZ/CDSv33D4yEd8HyfmAgn8VXN
jbKBGVj2UYZyUlMqHH12oapH/xZXL072EfpjnEG5ZXCQvNr1699zbJlaZXuSbRLP
t9UQOaarLQj2QgwldSQSQ4dpzg2HNpHVgBnkgaT+1JNjkdqSU4LqPYDkfM45tq6g
ULCrjtEAvW+tU4ZfYcFDYZmrKVU6UN8H1ft/ftZ+FSU+ILlphPr8zCGnlxn7Hioi
KMGqkVWX28s/pOvilbV5QA2B9t2MZUVWvYkC98neGfDeC3tZg/mFP3sjIzhFCy/t
fWRekrcxWBSrBIyg7E5y1CSjfp/fHafrjXU4wi1xlh/CBirMWnqEPrmYjZncZeTD
3VWBtLPAGRfsWoEmEnDXcliZwsTq34+H1SZy+L3cVGC8NiXLpPlzJSfzDWJjEwTG
h40n5iH3nRjYw1C9n2n0UvKf18zWnwCST1tMQEu+kGomd28658S7rzJHnwyrA5PF
g06NqirF+LWbsmsyCCckMYPhKh8wm2//caKFb/LHX7agPGtp0f0mfUJhJ+exBZid
jGO903Lmgnu/yuVi3UfaHENxilZcx/7NWMdpbk8nmu5wBTeN96S8blfrD+oE755A
Bq/V8Opb4ZmTeMimKnsLE65SL2WpxLVjmzMregpQyNNgIsqRND0y6i5zQGwyz59i
L6l0hMKeReJS8GwudBYl2RgH1B7t/Dv8+GzqGC1DM65LCHEoq8wyaa7GXmBLCEf4
agv6sSWf6LpPiYrbVMAWRetAQIC7vDwMfwmJ1RDXWKpDCiFOXWD881XlYaV12L6N
FFRaX1CaZNQbtz2hIKjZ/vfPLoqLeSWlLz78/E9IKmKZbtnWfFYKeJ7v/bD/cIyW
QCuVz6syCZb7fBpn+eHL4iW9y3ZG6IuKfn+c1GQlt5IvDzHyk3ChV3ByUpJBTwjq
JzesIQYjsnX+rS4xPGBpbXE3qrLkSGY9BNmPD+wNLAxGKvmqvk5WuGVuiFOW2KkU
Dm0T1NkgAS0e3dGbTJvSzktrfW64oZ8qJNxjIiMbhQ9SCePuBRM1NaI76kB5GXiy
jyxq5McQ7vyvkYO+i1uzmYSzt6Wl04lMVJUCC5SyvsehdvfkKuUUw3OAbU1ONc5I
fV+JcJwFXcxxEpQomRVF08KUnc5hqhgz4Le5j55ePJA9bn19Myk3ieMJ41LI9WJR
ekQa6aL6/ZPmlmXX7wUH3R6qseBp4BRyiEfO29vjExucMl+eQKzrb5qWisrFTO6Y
cX91MiAydw4jBNlWtK36Ozl9+ZuZEwnhzlc4AKcMiy66k8CRRf70qkIGmi9zNRKI
3G3aAYpzvRqm4NQGRaF2La844sxs3IlSViAc30i+s+LhBWVnSGA4W7eQaf51IV9X
j5zi20MBRJ207P5WzSPv2XyrzsN2JKWPS3Ujxq2E6MLBJFkFovzYYIpjt7k8fTPL
s1z3NuUS+sev4KyO996tD6CozLwtfWRsNP+HVi5oYs6C9fnYnaf90Oje761uI5ei
QNqPRzVbTQABywrYH2LKsn1HAiWk49vkpFhCL5q9kWq7rIaYA8SsOjfcd4d6lJ0Z
gGZwuo569zZgQuR31xa86axZEyDLNTNCsbAos0PMN1BqaYXzB1DjCvuJ+HibK869
1NBqbKHHeCJj/8fToq2tP2A2s51hOv0i1AKZZiRl/j2gP9yOIrmNp4q5JcEzqI0c
QE1OI3cXeMqtTQgvE8QhlY7ifUdu7QqsSMgJGmi1YjnkzlF4XJp6YXOUBZyM9xJ9
uabubiGIgUS9RfZywhZrz+LhMFrDY1sUagcT2xDgCN2N7Td9P61YdjmtZFAxsGqd
8TcJ7jYSYRaz7hBm8f5XHOQRbWK9vmAlMb+SMT+qVkSf5WnbeGrHThxZWXFjh2sJ
XmB7tK8frGeOGN1vQtVGquWM1bS11nefb7VAJX+xxBmblhKiiZMYQ98+jj7AN/1F
6QnWIkq27IxagbUPcq3qO+FE0wF6aKz0Ca9Xbrq9NDQjY9WSFa9kK7ZTpsesOjAv
ITomGN4QpvUqYvA3PUtnmrQCjGtCTVvJeRU7pnJCDpA8LcYsPYugj5iq/W3j0pth
ZISL+SOHmTx/kNm1CMYPt3iSdER97A0px5ZzXySXPpvRaPiz3EnMz3O5hfx1jqfM
H+q07AvABz23/W+TNcdS8iPf0Y00hfY7wM2CyS2yHeAsrRFYe+Il4tslA6Inygbn
cSEdqmh8k6qz4pChUcnvGVPVkznN57e+m+pQkb/OjGmpJ6OtYyX5267N0tUGBTKL
S3Z1ei027GEZJxjIs/Dn2/b8Nde1Ei9PAA0Qo01K+dnr1ZBvdFzSwsb7icHE8RTq
dYRJaOvFEpLjZuNks1V8MVezjz2o8g871u+ef39YcFXAUPtib/Pp2zsKnwK0ADwP
JpR8G0Q1nKQLAkL3hBKCS1JXC5130T+/CPlaHWl/8CUlY5Z8LiWCwRk4/QHr82dQ
MVTH1xEwjEmv/YZsp6EHoQmYMhthEWLQeEa+j6WH6oIPf1YnQmZjCzfdFpdjBTPU
55fD8b9rZoL75LZvpLSjwiG3UXePQAlY9AatcPf/T3c44VKW8k+/Pxx8n6TnZaVn
eQ8nvGFkO/jxsa7441mLrxTF+//egYvbPm0CnP3bR2UiZ8Xgap44txq2R9KJr330
lKWLy+3x01NhtOFhaH3sgRQ9wXCvLNaZm1qAMSaSwIWd7e2pVOFMqnQMCZJkLA9Q
1q4xMO69X6+tLDD7cUlTXwj80x91sd/LrMQz8+63LwCgFRI6cH0eK/OjEJID2z6S
wNpxuyFXijL97OTN9XdGGCAT7Sdn9VbdB0MZBn9jJBRoDWORQGIwjvi2tA+KgTtn
oj3lKiKjIB5LMuI7cwTLFr9QhkSbQrXs6puSHrmpQ46fAW4SZ8CVQUm3JzG7CMSz
m5Si+qnrmmyU657bQd2vTdNPjl7R4kd57RZ9yq9pYXy9mIXocZXqpjaXWMGdIBQf
LoArqLRstKpDTCNTbv5/dRBdLSOEsHcvZ7i548ulmyVKe0MHKz68Md1AU+CModNo
cOwwMOtZyMS0ToeTkitXgNCXtQVJxKM5XVapgq/qjbtKoWMPWbR18LB5YNL7zIzb
U4b+DNxjsul+cafaNW+ClbQRiXVAtHNOVn1vn/briDb0k3noe/feLf1icP095ndj
1Ddn4JPCDm8UENVGAiIM+nNOfQo7S+4ylcIjeSmvp66EDvoQQCqPBfrqXixfxdXE
otQ6vHwl1mUxGX91Qr5L7JCv9e4BTUmoCFaQZ5JskhjgmPV0/7FwSpKwPfkI5j08
TOU3q3UZRJQi8CSlc3QFShwe05VNG7CXlIx7XWJc5dPoJenIP/ec3wLyHS9I6qjq
Yfpzzc6LcJyAJIP4rKFo3TNE4x48sNb/F7KCxA+pV1MFnk+PckO03bJ3GDJHCzUd
dZhu/XU7tSdO+8WOL8yzWYgxcWwMUbkF6nv/2GxZqae9TZnH6PJ62l0ThDeURGTs
mMrfpP63lkXAIVckv5x0PouWyL9TOntuXiXXGGJql9pPc9s6UiQ59/PohYUQIdzN
ZtldQZxp1EMs0uLm2KyE9vOq2fXHB43U8NsNWxlRQbNAGLA1euqkYmWGcH9ijtsg
3l3sx3LfWUgNvexSoCDkE+lz6vANMJb5Ius3ptn4uyI=
`protect END_PROTECTED
