`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n2HDDTK9VIDOnGuxhfhJvAtWqkjTzhjW2BYzh8k/NeZpCqNuvHqvFDxaILg8M7Za
JxH55lyMqSeyiZVkGR+FfVjOVOZ7aU289KuremSLwCtU92v0cbxJAlwUrcxfn73S
GesxLmYgowbLYHUshTFzJO/qx228pwmFkWbMo+EM6+izb2+bAetbJCNcvDorkGfx
TKKjcdT59QLBtl2fpYanXtvbJoXD+llF4d4PkmAWhAGIo3xZWrsASt3MmhAMkaKK
9twFCqRUadl3XB2yZhrhT69XTiWy7UDxopawTAyVBySJi9EAQCknica8T6Hpo3LX
BTL07EBQege3eRFaRz7ZssDqW33h2tc28UboTctBcsQUC8yL53OcJrfXQFXO+0IW
I45I7sloXCjIWKPCvPhl2+4Fjx0C0fj5slhukuaP3s0gO90HajNK0wgdbOYDgoZO
7+u3fOAoBXV2iueVz4bqzfpNxR3DGLOeSjmOm7k94Fh5WgmXgYGg1FiVaw/AXWJZ
zAJ/fZzyBJphmMyseDo12tBKS/el+jrUUMC9oIqGg30ClMKJpEuY6Hx5wv2LHt76
E6eYVLsv7I8/9wTn10/MAfyB2o5vsutt1M+3YsJpPMrYx4sRullEDz8MR8KqUx8Y
PyUO744m6QORVydWNADz+WzPfmLBbRfnJvGv3VdnpUs6yRWbPk01j1sMuEUVSSgJ
qJmu1WukCNOj71gmgiQdUYaOrcD6rTMpBQupQZKoibxiWttHS5D0Z+1xrmzeJF8I
jurpqTCXISRcMoqtn+cY6dIINuKEVaElE88otdwP1fkrWceGPqdDs3EKGWbJCLir
aGxj2VHkx973Y6bT5jai0qR8YN1wQ3kVMaHxwJJcg/mJsZX0y5m/8uBI4gr+NssL
t620tfPYKlb7h3AEaK8i0F9coPWnRUT9IEoZmoMpVkFIVipMJFiroklbEcaqcGQF
D6Xwp4fI+8PPJahfBuNYGxaq4yy65Ofaqh14QExuG1LFpawvDKR0bNrd8TNVJ3nw
vhWe50vVWW6eWO1nhGcguwCoXhXXQ6kZONqZ3OtlGdb1g65lkiK+ebKc79mHoCGa
CfMqKtdG4o9bicnIraKubu3K4yJ4iApTsvvD8/PdjAHRc+mx3QjrMhaiSzh6cr6d
O4vMrUeY1vmthSXBfbIq0EVLW9MUoyTvQFDx82mbC8XznDesKLiEGfZ4nWzMlccq
l0vRyBPkrE5ZTG80oIl6VlRWzds+FrssbE+t0N/zdYtDeKNFoELgh/fcDg5ds3bz
OE+7gxft2GZKzjVl3sxZRreKeXRZ4KFrOQU7KB8h2S8=
`protect END_PROTECTED
