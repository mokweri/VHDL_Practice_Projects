`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XztZBEffZsklXVSr876yAc110t6VqKH/9BuS0Y4RXNI/RKe9mnVNaAOrl7/Oa7BZ
y21hkAIb66kFknFiIbYZgxIaWZBPHEpgJ8t9FPGNfD28XJjhtojWgIc9s2YzXgWe
yLgu65DiJJk1S5Dvks5ZZnDoXRRaMm7fToITXt9eQCcNo8G+AvBkZA0TcpC4C3sH
f6+2/JuC+5G7/QbQnp7X15sDTFkR9PwtKM+arRnDYIB5NCuepLTiVbUWoaVB/k7D
CIDAgN9nrJYhe1QnRqoZjH74If/mlIfpW5NKpXY4acQiJn97hEPiM3pYn1a9MmFZ
fNayUgnwrZ/l7uSzsuqlc3tNfGBuSqqUH01xbmnO2snSGOTdB/1aURYjx9HJ4KSv
oUqLGS9XfbpDO0fYdWocy8HHq2Sjn0m8yrrhQVJSUJ/Ux6YRTGZ5UEqmcqeYVVww
TDRWKo4kgwpfQuGJhTB72sQCbBZSKu8PUgEOK5SpbxhN1aWx8KMxJya9JPMAFMU7
JK0inpxZ2lUxhaAcLTFn6VLtzBUDPDFnz+s4Tq1vu0MV6t7UCR75DW6OdM4t59aZ
gOikpZSbXFvpj2ZsoihdFDmANygKxOlJy0VoxcJmfL5B7Nj4igoC8CQptVZsSg5m
UofcEgOwmOWdRvt19Ex/T0lYkJyLirKHLQPvgfsqc3R++jok4eVTwC5xkd0qhd+1
sfU/G5n0gHk8QWQ8xGaM2Z1URgCIxcVu8GTlOnWHymKKnXSTbtVBNBkjeKBz1O4n
oioZ3oUD2GRgNHm+JtXhsB7urfm65mNLlNl+JFGkqr41oQY2khfsBWLK8jbB5dHL
2MAbjm/pbzKu5Jf/JgRB8yFUAW//oQcQpW4I1lWNpp1gWfLgePUIHIvA48yLuI4R
e6NtdgGYT2njaIDA1IMQHH/O/nozttnASz1K9Rye393vZL3oTO7ZJa005n+/OKrC
h3BVlyU3JNAArLAqoav3fQtiLlRiSrpp2UfdcRZvC6o6pH5HGlG35RJGtYeBcMaZ
V32m3riM0WWHHUyZkdVIaVKUCWGYmQSkHeWGlmO5O7xjkrU8HbQSdliZjrUxkPiT
X1Fnkr52ZYFnlMIWLqflThfuFFAPvc7VdH5hZqZrYK5/RM6/pOK9vcF4wBXkWMjQ
Q471W9gsLn+xdrbD4GAvsGyB5tdKzEm3TLs7tjFm3Bra/SFIBaMa+Eo6evHVwu2k
XNxdvtRlcABK7sjoXRKVw08DPcR4JTXeJLG0Xm7XfEse9UCiVihjXgBJY8SYYGUV
`protect END_PROTECTED
