`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FaiUvHLxsWJVHgNlj7JVySnsgDvcdxxxZxxJkMDZDS6rpOt4uOvUaiPInm21oIzg
z6Vumqyc1/dLcEBle7/TFEsSYd8nbqWZW8Pna8UxKd4rp8QJT+mPr6GuAkFUDHr0
gSSCJ/Ww484vDl81WdnQU6LMSqZifcG1btj9+BDEbxporFtT98Y8GMOveKhBgFXb
feD7R9rx9S8uKsqMdsPaUZ0XlcyVBAJeTx2rFjewkX48aOraxerRmmebMhZ/Vpil
aUvLfCVNc2K5PO5L0ywsCDytKFPFdi0RUmdxZn1ljwQYyQTUci0zM+tBdlZeWIvr
v+fLZXj/gB6os3rx2fzp3MS3HvUIg5GBWw2HSC9GiPpsI8QcotPJE864mpqP9FAg
l17vhBreoWNCaKoJsDPkDKbfx89oyNeiOrp7F42nXJOLUpro8Z6b6c/Uw+D6mlYW
kL7DED4mFRjujvCKHhxqHHJacfJeVQd3XiW/H0ytNWcuSw8QFfB/5OBfhe/w4zFJ
fD2ZHuLeYqoe68fMMZqsm/VgaOU+BQ24Wosy5/9Jte4sif16KzAyG3enmG0qt4UC
Xu9U4xZuqmblgjVRFlCqnhBto0ouWROkf0z8P7F2VYssOpSvy7zf3R8qI7b//d4y
PGG2rl5dV4JQI/MmUskiSdwZCkM4ARNIiE3q8DUymjbdQwZcsq6tq4jJl74JAn4/
vznzxBjG/IYQ7wXbBRw8AA+/N1TWWxxTZyrORh4Kw8hu3XTjDW7keP6ZG71LzhW2
Sx/O2gYdl+xoy7x+aAFjK8EPuXlrges3MsA+DeYcPxbckdsrYs7w1PVuUjsANIRm
i57ebBZezkJP1Zuy0+rtd11teI+5WZsqzF+1JReqUlJ4ArLHu51Tgv7QNpkFrB+o
+29B51O2yg8qskCefI6TvkofeFO//yr18t8z52ZeMuEPAmqFsQejZ9IxO3qk9wRx
wAmaCcCl+IDUb+M8a1KoAgJIadQ3hS/uML5x+x8DCk4sv+g2arCW4ennJ3B8V/td
NhjUWfl0fTzl0l6ReBV9c2xI/iUzxX8j6MYg+Tu9uOoy04J3SQM2/J26LSy2Hteg
wAIof2DwehKc+/FyMDT2+BP6lssl6KAihJ52+DKDqhcKRAp93TQOqjhDrbrjqMMa
lupnPivcsoiY6Merw5aMJPh+DP6fJtosdS8Jv3lAE2EeUh0vOr1Dfi9mzzqcIfC5
SJE0AWbhZH/XOwp/H2tOG67t7BUA4lB7fAB56nKjE7S/eDph58QkI2pyvraV7oUU
qFtH8SLyf6gqWO/xV1kNgqCute1psoEjlQOKXVOiV/Tt7FXBt25VVJ/n/LMgJMaF
l6WQgQjgn35+bdnH+rlW7jseoOyoeFMhyFyoXQAfzG0lxQj48gAGlHLBxuHOe/E4
m6fpyCRmLxwFemTBWFZXkfyCcgeEN+de9Y1MGMDnSFZqLWbGEA94GJ5V23wk/kW7
q5jy/jcmKkfVO8yPTOapOER+pLX3bsmUiBvBEuw5OD6ng5K+GDwyR13zchZLgvEn
c8/yOKaEhNtaiTkZxpY6TLp02/1s6f884WnDKuw7LYrPyhuNO/pBjdsz8nwEo4FJ
MnFdO8c91yB3gMkTBsR568/XcF3XIBYXT5JGoyIQgFA8LNGsK4ehvRy5cu3uWOQD
h45PJrKCkkgiOo5zFHiihp9Xb1kB9QMAlevYjlFpRlISx6g66djSLYZM/Cau35k8
jSdz+xA28sLz2LgRPBaYLMKz1U4iDkI8ZhJQrEPd+lfXBKewCSgCmy8DO4E/Bh2b
R/2TGFlcAi2QTdAbCY5IhUEEAHoKRnh0UPiMKQWYS+uH8tjmENO2k3BFphA8Yoyy
3IOUMFFHojT+LdjoDhYqYIBy+AhXC5edh0uBN1y4p63X/cPq68wzBYm1w/yLEBUZ
MQ/lmRKRRdvtUurIC7oiu8iGC3qPdYyiYLMA9zsneGEsAWDWIHQ1fKvTl69RE8sX
fx4X4nCBGLnYEZDcS2fy9bWUu7wfBy84fC/1MQHOJJCq3EP3GEqS7rxC+RAG9f7P
qHVJRr4ZM/hXOU/cmgogVU2SpR4DNTxSa4CdfJyXD2Wbr4sPuIQz7UG4zzj7JfY0
7hPQxZ782vQ2C4Xw8/vTXvbRhlPaWUlWgowV8nWYPnBp1+MeGoX1Jfg0f5QrB9u0
S9fqmdQstVfOChNkXd5dDP9CgL5wySn8uLmQKBWooNqUIDxHBUNUGjnyDGJJQRtj
95JePQWef/PYr594+Gf5GkbbuvZREmQK0xAPAZAhGl6meVK3qqbdMlGI9b75J92g
uj+jwLqUtANWyW84LUael55vlgxw6ay+IOEaHy9IP/yxvUvAoazIJQmZ9ChD82/L
ZC6loV//SprXBQ3qRRVpfo1cNk4XscWFSy08YSnoz2D5/E/pyy7lYXF0+saSbwqI
PRgPZhCBN6BYmg9Y6Sybdf5ssFSBWvB5D0DuG7by0hfpzom7cUD07rfneETpxSEq
gSjpzXNwQH4j5guaQhZdiN0d3ytmoN77tkWIYVpLn/wvrKFm8DzzSLUhKK/Y3D4c
4Kxmg6DRn2INCGzTGJ1zjvFv2sC2+lwzmT6PkpY7q0xqWUGwb5Lmg/O53xUc10HA
1DN/WSn+MdI0jURXhadFsPSg8OYXhdgI+oKugJlO25H56EMkJE5vlJcmuM6Iicjt
MOA41GUuy2dy8hBBNoJhnMbznIDpNTMaAFlGoZilhjmlIrOmow5jaoPOOCwe9/G8
WGrCeewMG8XESQtZLKgwP1CZBy8bNtLyAtqlZzQn7S+JXgZRxiHLvrWBgDi93DyS
Z+F9gxsFCuv38orvd7uKInITnf4Cc8SS2GGGaRZuB2ZKFiWUU4ZDqqZsJWm0KSNC
j8SQBFfTRMWdm4SPQvBYhtssdAuSha6EGJ7FUlpncfZCB67SoucNExacvftGcZgM
vHJwEn4GBHEns1ZHQFL3bNBRy4ioxFVKfs2PfBPlDgHV73cSNlS4HO1PqfB8VvDT
U+7oQLwpKpBelKHd/4UMn6Ljkf4rk9r7SqFujHscAwkPxb+QvKrpK1EK6navWNkz
TyYWB49Hkz6JvOz0TIPaRJSKB7LO9Ge6aL8Wc2dlHG3qjD6y+jj8a72fiWDLpPCE
yo7naRy1rak/77bF7KzzubLOBQR9WzK0rHhpVSHsK1fhO2Otm3ChkvexOroTvv2b
xGcfUkp/p3f/xK0Nx2z0thCg+Y7pgy0+CrmkddlloiwFCNnpKyqYf6HG/fQxQyFD
LunhQ6TSgl7McfSTePrbHw==
`protect END_PROTECTED
