`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1uqz2iFIc0tvhQfUhhTkwFiDUep5cEjQniGKw9dJqbwlj+dRTJDRwq0EXJMmot3p
o8h3LOidviREfsC8pAwY3EofVd5Nb4gERRxe2LzH/L0O1eOYQq+U8Eru6beBu8Pw
9d8wvI29Q/biirSWrN9c9keDiYKnijNcuh1XV8xH80B36M3ld3AeeHJylWjMXBb3
MPi8gHowmgNY/8qJcltrIAWmt9HKFtOJLBapdH2/5v8twQueqRHyYfnwK4f0dxLU
BaTjSsUy1vjBU4XfosvBk2/r47UdTa7ByUYKJ6x2EG/aBVaUAhuMilEfsKNetYSO
3iHNlrJJC/XeqSmQD1NGbrI9ap+ulqqYy3K/5Y92TxjV5MqnXirV25VaFzfpQWrX
0tWH3dMHfiyegvArK6Bz0OwHB2HSp4N6ezo8xaO049KvFA6SACswsmS/rW3HOAow
VwSGxyUktsOK95jjwQRKTb6m7mWv9xpW5Br0CbWUg5m0/JuZPT4H8VazeR8iUHsZ
HcuTGVEdEaWc+i6ghq5thqWQZ7GtiYIfohhgR0lpJwMeRXyGLTAJabY5dHTFWOlo
+JCvqzwZ+NAc+LlwYYZFqX0dNUBEA5ZZbdAae0GiA4owGp4uEP0OJx8yhYXHeY++
1qfSwlJ4qAOsQwvwNKlPuQv2ybbBJ13/0lpqlW/1UOlH65bFgrjfCsfCnJScyRux
1fAHi5jEhvNJ5djfttLqCtpvGfWov1cIIVc8FENM8TpLtCGSm/UqKHkfWsgqO/Of
g6XnRWriTVQ35UhUUg3E8GeMpYAD0Q6Cpor8H3S4HYavi08JvDAvxqwl8q0moldK
n49Qn0xV8SCBDvgUfAND1X67NM0a5uxCmYDIwYOLul8H2/0odSj1+BP8NZ8u1ez1
KxD/FhSYS1h0R9XvT2tpMDjKUPYRAfb0mxocx9tcfV3d3dWZGmWWw2lJrgY5GIFn
n6qIgZzBOsFbEMTP9qGNu+2ZkyQnIE9Wzm1bbVXebzWW1KiwtgtLsKmPf6bWaUFs
0VXoEFcDhTvvUiWbfE0nA5du/JK/+PY5dDq1DbAVUyTJEgKihHd64nqtcw99cQuv
eO6xYvjALar4Ey6S/Jihf13RipbHj6oQrctoKli6PikhI2w6UYIQ4GmUQuEbDHiN
sCGQGffJdzxMhtwm9gfz9K6BvZOyzUX9Ekr2v0pwChsz7ntH0vcToVHeE2Sa4f8G
mom3tvtIKjLMMUpM8xx4NiNa376VUg/azhLa+0bhqUw=
`protect END_PROTECTED
