`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaqoqVSOdBo0Hqb5Re1vxuRvF9lJUCxdYJsfaPEAllT/PM+2/EZW0BvVajfNoWCV
14OpuyKC8OrXhAc8iLy01B3hA+QCXBkegyO6lFJDW6JifuRpioHElQdexcej65D+
wyGoqwh9dAgmVX/+9ZU5PCiIQqQ34+r4bNAUjXM9saQH7f33Ckf0RY9DRcH9H2Dm
5n2EI7Wvrc9JokGdtkBzvXaBXDjVqhSFJGkFLG/KRlqIJUIQzIUoAk5oFy2e7w5e
Rvwqx96HV8gTB0qiJctbqOncm5OZh8gO2RqLWkPXCiTURwfkkpEZBj5sogkEcI7s
vZ0K54EKZNmjkE0+6MbEQwFqnwjllLJeedk00dMa12rfo72pEnipbScvm7xghc8n
3Jh4ISwByloUk5utVeXjExL8l/6HVgM8/X1ZZ1GwocGBZyGWzHWqrgWBEXj/jyS6
Bf4U4zUpndAXl/WPcEZZ9QMVBpna0VALVpx3neGSfvDISgilXxiRcKqtTXDw+B77
glJikkhNhOaAXRKHl4QHTULuYwhL6eeDLhGQ/bp0KEu3C0KvyLy+/tyXqZkWJ1qH
Z2Djqhr6UpH/4N1h53YQAUI0GSs0AnQmQDcW7p9fnsoNU8j/ZcyZw1ukKyc0dPiY
PZ+bSZllhykbbn4lFYfwFVAbsyHYONJUwN+zvKqHnu9wMmiGArzVCGLNk5lJ//Uf
e9b7TYRTc8+eKmIJ9/88L8O4Yg1zMujSxCzlXAcJDqDmR7I0M4rKspUpCR9eFhSU
ShYzaMHH/+7oFjKGTG8afY0t9jAoFWwCqIMtM93UjUZgdUHJRU8fBWjG69h+xwyn
ti5MZ2QttKEzk09G3pcAmccUgVVU6iMT/cBvrEkac2UWnxWNgTD2CNIPj4LRqADB
afpDQT0uEntUw9qwblc4AnWJMuYeIOu1S1uzyRr6ioSedJMUrV0Ov60F/+BGznk0
LcQKXhIO0kNStMx3ZFOpmNnqg+PwmVaHcbN5UepKRURswknaiTePIXaryy1hPnll
xAH4dif5ok3/k4oB0XGmGbDInlJ/r98iqXckK67+AFbNtdMteQAWogYVAm+n2ROQ
KdivIMwlZhl5APumGNy1dSy+6siykft7WcR9dF2t+IQDGf/dcXO1ZIB0c2FB25zt
jxsMbLujzvlElaXxfydYPuvotuNGGA++X/6S5GZAmcDzl05jVBMIFY8u3I3OfKMX
D45E/HV0ls+lUzZl8G9YFSbuFuSoXeuCfQenvWFvHiUVVkvqstm/KrElhDQaUGcX
dwcq1ef4+FikFAIAnHmjEg3Lhep66iKLYe7HZ0qgyoytbYYpO2wH0HtN7VznMNsx
1CkQzUbUE3F4MNLulXJ/53gKz4lABwrbE7xfb/kvkhSmhKuliNOOQKas6JxA8jZ+
BMoT2HqJcDvwp3U7IlvKgc5odq0xj6njrdtR7YCtTM0ssRjDjPBm3OVUq2TI4WQD
gepkzs087PJCZwxLHddrYGAYe6vm7x4KJXPdq91C3HlqvCPT7ZgKsFrjbVH1QJ0e
9gmUS9oAea6yX+uwr7ST59LhpDf/Rct/fxGbIX7ytABD4CmXgVdSIWPMUfmkrmC2
610N0uxnuWShdNAGPLcMgZHBrCIyAUO9DzU153LPZydJ2RShh9Q9XqdJyDQ447tA
Uit5P0saTkVuzcf/Gu5u1azLZlu2JgKs5MjidfZ84d9YG8diqZY9oDC+K48NV32t
ry5LTvyeXE/+csojUebdUpl/5yJwyHCbAt/q5ypTM2gw+qDL8HT5LoMdtRh7wMQD
J4C9GbblJk6RtOET+R/LezbvwGCwKz2SuPy+8Lv7DDxnxhrCVEspDTVHdoZPA5xx
XnUFxMBJV8Tc9zHupAZJAowT+2ikejehrSA8WHxFYAfMejP2P8W4rqPZ2lVa6mQb
eumBX0KZ5XfHh727gMNynFKImxxuNr4TBBGtgp6e5L6oor5KpVSo8dQ/2naQpQ96
zKFCMGL2a2DNFMoxgvwIKw/6RyXa/mVFOX/SlzKheRAMM/IVJqpqWzfsmATXmQ71
HjxfJ6s5UwPHQgf5nspSEeTmI91FGVDS6/0OhLmd8NsgriFwdFmpa5QRKoLN+8J6
lmiBLLWyrdftQZG984Lhvrhm8WuOLKMtqcoASP7465Tc4eKr47eUU9sJzcjvmUbR
Ly3asQYxQpaz9XZQu5XVpquBv/NEvun5nyFs4cF0zKDg7uviU+fyJ9IXjoaPZt5d
LJsUAGYNoWnnMJPHazu3HmoftSFv+XupZLWd28+yxGKj12SzLW6FfHzAFD+9C9fI
sB4mTqhx68KOCBAZw3P+WqUFZP48iArU2Raog4seU0VyJMhxha1CUpPAbkcTtDt1
wJ2XtTYguTzpG0DQ1oYN773xNzK66xeJyxkRP2tFA3plbOHMmzMHMIbuwAiW7tkB
dZhqWF2AVO4iV1B3/g8bw7Hza+gwVpqdub/2xjCSePJTNFiSVUuMRRVLyn3pBqcG
bVCApAzb4ZSzWA1VioghGVAvpcJvcWrj27edTektpGM90OJUe8QYDBNb4iNd28kM
IycDTKsrLt9asEMx/96yIUw7WXcAW4Q1U1bX4T/9rtThitSFSZ6I/vjBQYSkTd8l
QC4P4LWZRkvRDMZv0nUTFDpwXs8GJzY4NJbWc47tFZ7Hf/pSOZdiMrwNwl9VsFtO
CZ1ESKLpIDrLxXn1+Fmo10ntvKhd9/QOxwld6JKcQ6+LokJVXPEeO/Jo1sYaUuC+
a1rZTF3PR0EqTXg/IL89yhSG5h4zDRW80LAiZLLAIYl1VK1V0DjsYFokSLlk6qmM
v/bHm1d9+OTs0jIUwMyQGHXAF1+bHdrdziTqwUD7e/33RIZzcKw0PME8KfAWMQLw
6dYI2UdcvcnXYUT0qgniGtGbRUZ7B+5QQOmlcdBZ2/TYPE+g4362Hmp8t1oHT4T7
DXzlPcSh5fUFQAdBL7aG81yxLvpSqFFlvK+IL9kJ6dWYDV4rSZPu4uy0OhWbRPc7
uuhelPYaucxoxN+LTiYu3dIjMgC6WSTC/v/Kvv9NsPqkZRVnXNlg4prDwVfVqFkV
9vdi2V8iKYKOKky9fEPFh10DF5/8dryU4d7SnYrHDtoW7sJObmCqfhziSDoHJulH
n4V757lfaf5Zgm3se2BIrvTWqIZlPfRUxnjIWqa5QEqTjSecrjrmMJESWPpCpQjN
ZYynpx6+2reMvQAvjglvi+wL3XU6/68KI/fUMfb/+ArsuDg7pAs3eEQPmLs0/tDP
N4r+MkxAROktPdA0YQNkkWG6rCGlME02pM4MtcYLDdCjuhV+4DdNufssyKlmi352
LaM7DSM1c2WS6Hx6N2eg/YV7pLfWS6XnijMgoIt+Ak4rcSGmZ+i5Tdaf+ERHePgS
/GLlgcqIOSutCdrG3OVDmIXmM0NAHpudOIry9+4CqDjJ/DwdOnRmqGYGq0QQxNdr
Bo4LMa3xJcypeP1PgIr//mqkXSeEaQToC/yoEWCz6jYmExqMI0aHLR/WbMtGnQ8T
vCbfmgTDm/2+uj/B7/eNQA2u6VsA/4+eZZkcgGguT9lmjlGejhHkkO+4l8XMYV6+
wOuWeuVRbTDh4fVWo/VKSA41tw3j0SJYQHVdf5p7kvIsWUaWtMzva+efF+sFeGaw
wE8/+b/GXAQvT8l08IqJ9HUF4YeU3PHkPpgKVDMuJzHJlt3W0wAUat1BajPQ7nP/
aDE+oNJk8pO94g9596rRcHQcI0BpW9GqXygf91WPVZ6rZSqejD01FlEIFvubEQpC
1fHPHJrzST/W0m3jIPfL4cUCdibCZq9goVB4wnxFNoSx8SMVfBtmU5BeWY6m1Q9J
c8WnR7S6UwYHOY1RoZF3F9IhZD8L51SOZldOkuf71hRtXK+OATBwib+oWRYlamC4
MJ7uPFrRXb9E5SPKlsR5d9bPAbMBruDaDagwtowooOISOdzgPQETnslWNSrdXECe
xoKPaWxW8cIwdOyWXpK5s8IWQ7wl3FwG5BuvUDCs5Ik/pcmmqmMnIccG0p3fHPg6
XJC5J0ggQJw16GhBt04mI3N+rmWIKhK0CECedNj7QqN7lQoGp/IMlsuAegIQE3Xd
a6MBPFGItNQ+dozOQ9T+V7XTJD4jxWlOoywE9XwABY17u5IdnQGrW4i6RTTzhFAM
RP5nd65v7sx45LZ0D3UmRZV8hDo4zS3T436nC8IiMYwqbE/vzov/giEjzWq7hPrB
i3mi//wTmfZvo5h6sytd6MH/wLtTEpnsVK7egtsLUWw4KZ9RQUDgsC408DMmzpOm
atKbMunu+B2m9WXfXtzDu8mapbD9Cj1u3+n6ELO/DNSJeTWk0KxdTOUs/FP/EXBl
mfFSGVXf7tdmrasomEaGpRRT35ac4BK1D/uSsgiFVd6yZZ7Pe8JnXleyIFsG6f53
hHExKMi34Kz1Sk46u2ZbilyTQr4VdVPq3PNvVKjkdU7JF87rwVsGlNqw68PhvNhg
8M98VoJQz9b15dD2JyH3DRNlkWTFtzw7PN7EeVhsFJiMHIITClxRKTL7+E013iaa
Rk4v/50dLQtkttKrbZf7Ef1d+F/Hjttkkd6dsCmKsFHRKpCKGaOKSeIEp/o7m/2a
f1iW++wrUbdSC+g/1eDxzLDdVviB/vvMYWTpYaEoaEvB1qj/oNP5WzDOel5chHp3
BmTw4yvgcgw5CQnIjLOGL9psJNRQ/+wmvcVOrmE7JOLrC4dIWDrMPMNTGbqs/CpU
5gEgdFGQOaogjZjyOg24Ud1zXhB0h71MM0PNiWCIdcudDDkEk/TcUOOpJa4a0IWx
W6wjMKIaqwcryQTgyQes90KFwlgc2gPFYYQ4sIbfvP27fsgpm+QKS/o3Yy0XGBHQ
O20rKpJZlRzBPmuPsagnqDNm9UEmz/eTJvBgJbiFLt5H5QH/G8kWhVCOA6PtQSzC
dVewTM9zb2iHFgdje7Ce/NSpHL0NV/t4r1nxt4EFswqh8E6M5i09FIEmlJs3waTc
HUvVy5m7IVSuv8eoOuQvPiN59Xbwbrm/J8pRGWsWsy+n3mEID3G3t2MIDlXg5NSw
gMcuWHybfXtw7WFK/2xjQm8xUxhMCQ75ZPfhi/WfB7qWbqBjqpEMGXbP6ssOYiv2
UGWg5xDNDlYZWb4IVf0x7AWxmnHPRtdVqBJwCTNTcca/noR9sdOTmSDFncniighA
wZG6tvHnPGlMF4kS3OVilDbExFGjM42PIxnJsVynQqSpZ8XXl8Y8qpCmaPTUH1Mm
flMq08jWUkJskU4gHT3q8/wRXW3VrpJZyNtldeCidGTocpuESc/UJyktyVCfzp2t
VymcfH8Sz7nghpzXazXDjxIMRgMok3u8dIfpYnfH0sW6oLxf3ohzYB4JGgEguuTZ
KDxjp3Zd+NAd3VQK9EaFkyY+uc1/m07eJYthmo8MbT+E/OND3yvDqd5LO6cdI6hA
+F5IKJPT4OahcDdbVQ3NZQVFywWKmyCYEf1SsYytt8aZr3XKjvwkFo6RHxEukWYY
ia43cog1z+uYhQqAtUT3qIHmdSKJkP0lXGLsj0kl9lsy55b9pKFGLf4M+Gk610z6
nwoB/vw3FRZBftBOKyUYgzyp5C4zAwTn/ui8pL5VkiacizVs6fXBx9TpJD3h6bP3
mmKch3n/tEhJ4++p+RRM/erMZzBWnVqb5D+pYxPZQx/MDV9m2YuvM4v6nfHc2rwv
yyNSTzb369qiuhnXsUSmnIPQ5a8Do7ugkXaKERjqSxYJUZ+7LV04CXuNlOW2YxtF
K44rSSASNiXPFIjNxqr9Pl5GXJ5Z0wF9itDvabiw2yxeg+hlimLUGL8uGVkM5Bf6
UcVYLngWbDT+0I35nANG6kyVz5cvFKuLzLc7VIU+c2iFrTrjkRF3tSqYS2LOMMLF
tjlNuUPJ175DJfwn6f1pHNpIo56J/MI9w/7ZtnOgU5V6xkLo/FYlGClZRmQrqCYk
QJZO3FaTiYwER3YbkNxnBiISAtB+brzgG5K1e9eVbHxsBQXgP1g3dSC/9MaugyEw
+ARRVe7DrWWDBufmSZriFyyfhNFD6imaKgvqQ4CB9z9lLUqXdRjt2TWcwpn+UYTv
6rblFuQRbrbG/mwh49gku13xL9dbbx/bE6SUcJzuB9QpujM6rMbIjQTeVZHAhpEE
C53JFR5wBUsOeJHosEDwf9hK7LYfkeSJ5wr1l6wwMwPT36JapGSxyX1Asl/S3L08
8pc3bCvZQQB4qkU+oDuRJ6Xv+Kbjk0tx5TMsuzmjk+AnsVV1LP2JwzVqwLi6Yt+s
Iu0aAGZlul7CCWnFoGLOaKnJZUs80Zn38Ohi7ihypZFA4z8ARZJKwuxANQxT0wIP
iX2COVNn9fAlCRBZ8SbtKPGnCTFLNawRtkQ3i191W9sqTnrpHlacWRhvhj2Jfpbu
WF+AyM9CCCCseC3BDZeb68Y9+MrK+oqex/xJjh06PJKCZFnY8A+aqd01yXbTHmoN
iIamSBJTzy2yi2fFKEOZH70hKOTU8WSy0ay+alnE6KoyX+DzUvAsfO70WXT69B+v
2/xgPGLgR1/zOWw3xNgLj+IugHydBajg7bMsdBSqnp9Y7S23lSDoK/rJbz23nZzL
3rARMkMm/fDQfHQgcZ3wkqS9ed7T8tzQzCiWo4bfwn6+lO8JF8V9jCQ9ikBWiV+v
N0CbWNDSKx3UkNcbnXQfOnSGjp6+WZcfc2jrD5Iov1sWAwdOC4YBvEXPqCxBpYtp
oGZsmuQjdd10unAVFFR6yXUcCL4YSeGax7X+4sSUX0lEF4LI5ycvBdwrv7HiGSTW
ByaI6rLD0EOJ9MXzN46jmyiKn4SwEHZz+pJgLPNOCpbgqX9hpCeraGue0wclIIZZ
VFB8afKOgfvaslyFFCjG4WArz6oPoxKJl12TzoaSwOQrKVgxtOx6glhv3JkX8leT
z8zZN+BzCqPZmHsvfw9Cybv5qdNl7Ubd4bCEpQF1ChVVneSe/i2v4T81XP4vWYOb
Z7aQJOrw+uAofCfRcxyEuXWMI9iZNEUxFQEPnxRmLY2rJBAkrxZhJulTspap5r4P
fIoYVAn88aF2ZTo5kgqq4A25+tYOW6/YoaZxcXZNMgBHeYMPux2R6n0Zni+i0Jvj
vLdKG20JmcEyw5hAFiqTVqFnlIgmquTb0W+Y+SI4E4QV7AReEe4GfSa4YbI1kc9u
BJ8tAOf+u2xmSjlHRYJ32UzvZgQ7mxwYa/ztrd9+uVP0xV3cTX22GOZC0D231T/P
aAHZkWd7An9jIbdgZplgTk3fg6RsC79ZAFfgiWQRn+lNMcn3FJsgnC1iADBlRBEg
ezQJGuj4oxVMnY195liKj3Fe3+yN7FlIQadz5OLpF7C89Bd1SnOudFwM9ZTDZFic
t8rEjSwiAqY3z1WuhAbRDt+v8NEifR2csPuYAWwCbvUm3vO7ZDcH9SvpGENl7Gn7
NdMOgKTzVxkZLawG3LHtdlTgY84fwlMPJLuoudvub+32Y1lzfm8FvQsVr1OhtkNh
gKdkWlcw2XFXvLoq0WtIFmFc0Xm3QsLeB5+OyU8iy0yGgtQy2FylxWvxIzvDBw/J
LNLx47eYtd2IKPCBgp9RqkYd/gOXfBVde+X4M/tpr/EjVotckkEFhifaTAv9zh3Y
4MUr6s63p7EgQb2zj/ZmePvOCTuNJLp0QA1GRoMvJt0pVDZvj9SsscfRd/+TkPVV
TfvjTZNGtuGKE4WNk5xaVwICDX+0hBm2y0bcj8BaNW797LPV4Dmr73U5n+vN1aB0
1n8dg1ZLrQHhtCGnzZpaA1BE+RuWUbw79CcIFOuGdWHW/5+ZxEmXGpy6gUDfEQcM
UNegLZyEndvX+83q0DZrVCadPpBffEMP3JGgYuLMup8sTyyKNsLGxnVny1RUTSNK
gsB1L5MY1xhe78mSwwDTyqexlp9h+NcmZ15vP7LkyHL7r2rVYEZQQ9Uapi437glY
UiyEluGEKx7Ea4Ast+qZ0mSg8Nagg23gpzgFXcgVI9JMotWx7kqVXh9awFPIfOek
3fppYrEJpmwvsh4OZI0InleN0ZLxIP9CJ7eSK+uaHy0x2mGp/7ppJ/UhxSORZ8Rw
16f0wkxDta05vG8DE0Sdk6K6TN8dODgRNNGCAlup00gh2BIe+etkDVvW8AOCCWbs
VW2sX7MDK5KiuQR4yxnj2tg4J+OWZfXLjtd+WPI5Kv47O9vCrTn2qe/X8wZ8qaJJ
6kKw6YyMijUu+UiicHd/5vlFXu97P5Skl5dzrosgKm6f+fXw3DhOg0x9r76cErdF
lKX2jUKXBfOCmyaVS+i2ek2iMPlubTBIromb3A+o4k9DbuW6XtXU01creYUfVsfD
Cp0Xpp84vbvrB42esh5ygIj2NU6hDU7d04KZRUVEwgxqpDhvOaVF/Nt047rWWHVa
Su0v7wF3nVfD6sWKLmtFRZ0+luTYSIpe7ANmBrn0lFE/Iyd6l3Q5ISrWhZOAgeqp
h6kH0MMBsrSVmZYWZW+zwGQBAIl3jZaPFMtdMBPKcQX7FmGSRY33AyGyCmRoT1im
l9Fab7vSGAMoflhjbG/DueVM2pu50ITo9PQdG9sArO1zGAfW2igROQw/ee8h0nxJ
iASJb4jBMwz5tnhCgOCSl9um0Qgo+OVGXCaN23hKF9Up8/IChN1iPPTdsAfqoD7n
qNHRgCQW9b3pRySD+f1skdNS5yIyOdHs0KS3GLygzFGQHi+OEeacWNfJfuIPsrCc
AvmFN724wNgyGmKpSSfY0bjVHC/9eL+sgOHYZcX5PbfrRw3JVddCFLxmjTkM/kdq
L/gJJ+6wzWlIHTanVUPNAXFqK5HqNZr7ZNCGS06CcFIzV0Ao/amkWW6MAk3XlxP6
BgbOFsbWidLhyz7ugpQO/tS81/DnMSQbkrVXTDh0Vj6vLhr7wBWw/7GBQ/agCbCB
4vudbF4z9qMBngvkoNDHbcdfE3mtU2xa4fNCJ6NIZzEtHkZNd5h9y54w1VWanbTB
5K+sqL2lWxXH/QiDOicPm4Z/Ul7iMFK5lCNzVF4rbpQLAZc0iYjXknFLav22J/rh
0o2JPThSL8lX+7tvXJVh6C7cVPS837cBVTCzUWcNRyOiXXN632jJr0MNRZpDnSt8
twDBrdl3AkH2W0MamGQfHKegp1TG388Zb/QRF0LT2LD//jHuHX76Er52qCbBNW6u
iNznuVy2O16SzqALozGYgAGJl+IwXtdg/GYEscLeTbEZ5Sle1gcKmMuFTWZ00zaD
L1wkzf8cRVWHU3LHG9KRsqtPsdovEN/90iwAUJ+9YZ81nK5ZPqs/AtFSEVscq0w4
TtBRTvfWN1LTisBdQTOwwTkQVfnKxoqAtSbWj2hdPjvYkNpZMh6LSESroCUINMVn
5JjP20JEZbjHJsYOTDUUPED+abT5EbJwCuAaulI5sM2+A4UsERcnuXnDFivoCTnZ
SDP0CVOYsyo513WI6sz/k4ZC1tWUr0duVlrQH/znA6NBjj043jerZ9UxIb5i7Zb1
VDmeGpq8lbLwHkfk93WGWbgx6Y40uWojQAFBde66FfM8PbYlxYWoxQSKtmx5vOx3
7hq6m4b7flEBZ32cCXsPGmedrw/euJVVopA8bH5Tu4LHsnrID7O4y8jZFuC24Am+
h05hq05OuvPGV7h5KZxx18zFBLQfmEyVH4rQ9l+vbwfIGGGINVlYFKHeubBrXyXg
IuDRUzG4ohhjID/UbsqRaVrRzlSYsZtz77frQ/kft7sQ0eKLFZN5B9mzoPniKrcb
YBGcATZOYvO1qsOXG0W7dEDUfVYKJicBiNLT8CHrpR7ECXwxQ4S8xId71Lk59yqA
oEFMDDVZCtfB8DxhvmG9Skmuu/xNQB1nW1wYyXwEGFkUIIPuK3ZibeMAyQbTlW+b
oIbNNBTbT2ZkCujs5hwQnBfCjOwP/q+SMcjht6AW0kNoIKlHQaU5cms6nM10SkqD
1yJPCkiUH9olK4AQ+Y7My9rr63M2LNDy61bY8yqa1OM+ScV+O3JUFmz8YWcg88gb
UEGt/oOMhwfHpoXPpnrxZa79NM7cjkdQPK8PXzavjO98g64pEh5kLOsnU2n7QZVw
LZFmShppv60tqEBznZtHoZiRhczxVBLjtERHNda6i8BebjcX2kCwHUObyJNXQTxF
LZU732rYrmMiUqpDnvAQiNEwv413Jd4FSLiK/LSrnRDug2h59ByGHuWcjdJeEzZG
/QBYgZGK/UewWQfMpoFc62CPc4rxpV6Y+IheegcPknWkBc7FzRASW6jmid2ciBFK
XsmY1cq8kOSPwvGvjVnxBiDScc2Bp+OMA+hBZ3pWMAlcg9Q6YML1p/q7ZB7PyDji
zpAPHK/v5l91qUdOTzsTaAzEaYy7e3izeP6V2+7Ov4sn16aO7jlcxX6VKvX3kXDk
2wF/3+rkfy79U6I/FPuYFBokF3fCX4SifJRF2G75t8DvmCBVth9KvT4i5Un3qCe/
R82TDopLPkKmyPgsoHBZPyulC405tGu67Ru5vx0WQ0jg7nyeLYzxvRTYPia+BXgW
g8bMO6du0Vfh8gjbEMog4OYKSTaqeyIq5OFpzUMmPeyObP9k/72pdyOUxww+hc8H
Ugo9zy/8M5RDu4/QgYELoFhODF+L6y7XCoKy324DvVwlYptk8vJROfP1ahrGyBDC
xuj+4tdHk25WN4gZ2Ifa3/TpvCbaGpQKTDPV/FVtXOWFIwxoOhSkdLa2ZAO9pCRx
zu5k06riK0hVcxRGlROWHw==
`protect END_PROTECTED
