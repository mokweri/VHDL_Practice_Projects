`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6haTnsxHk5A77MnboDHYtZCZi042uOe0VoWTIPI++FskcJowrwbpZnp9EVEYSsBX
+v6Qa4YA3D20aYC9Gf3JN0uujR5khQgiUAiOLwiQ5BOK6ZhQ6aHNrgvzLuJzwdOY
VOYqsL08iEmA/jGlOzBi3z2dtl1giOqNrF/snAnS4HPt45Ia8z8TyBtahhS3Ls36
CjXk/qbxYWqao/eSONVoRGYK3goWG+Lv4tgR03KPA8/ZMS4newYCiwv+LVmFPQsy
LjFBhQZY4fWRIxVxbKHAhF4wBku28+XwBp7rgUhW+VY++8FeziDKihWvLktIIwb+
aFEoFMxOXZHFQfVpH4OU35/+BEB4mm0m3g6CdHf5Tzc=
`protect END_PROTECTED
