`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ajxZIa+1aVQQWoRW4/YpcAU9kSQK5TkKV7j6tUvRx27ldQUrV1MAQrX3YjsrEaG9
fE+8oWm/h8JF294ThWrdjGj4BGSGF5H6+eHNq9LhOFnMUF3m/bxwxQo9vyG0BKNP
B3zoE0pHIVEPHReRwAGkTyV9ZyKibC1xbRVEWtfRaCs7gjmzHk+oDYhh6QKdVVaj
BsTW0r4tDcH6OoIVdL4H4lEV8G28DVdYl+9xGCx+5dQoOalqE2aSNtLq9xy7IF4x
vxXtygJHWgWl4fqK6sseMFYeVPbCzPPCrl7CiXdWnuZceWW+dD6kQsRowOGiK4IV
xSTDYFLKHje0qZZj1xB38i2n9MH1xRsKD+uUZ/YBS5ctiQsCnPMU7Utm2vZ/hU3b
+LyaRmfrpPuoLNWhqyBX7FOIAnYqGVwleBvg2him3kJpxpKH0j2TGhvNb0kHPno9
q95PX0YwJXMzbc2PMAsy2F1ejSJEDc/E4gSwNCtSxLc2/GyjoB5uIXJJSws3LbE7
iC+EgQYUaJhvSHPt1OnzC8/jN2qRxBF6SHYpyIdMO9j8ZPJI5pZFVxsaGK4nH6nE
+Nv6OPqeVVydj3nldv4kyFJ+dj6hUQNXJv0M8CEUHCnb0HYgmDLkctrFJdCqIX14
QvTZjiy/7Wl+ZwA4DknHMl13eJ28kXxxEX+n5oRMs27cpmi5dTwPkeW8ZFB0TGQW
gwARQQNE1GxrAVhF8Y7ebYfY0z9ZpwrSxA66Y2WIg4tFsJZ+mjL4m/PJqHASb4Ri
yPL2WPKx37H86j+1dSH0qdGDV15JwRwCQv08rhXzaGGDQL1QL4m5ZTo0MCnedvOs
6RlygqA8VCNHez453hyaHxFuUsv/H6pxcOim4nh+kwPL4hYVOgkCfPOMd0cIWy2v
I6Ft0CFBtU4gpV5B/8EG+vGtiBKeIRQg9Jl0tmTMKgFKg9Uod7ICBjGGoBRAsSby
O2oITgMj8G9vBqNFZzd4nPyTPgr05nMe97hXucQX5/Zu/WGaaxb5zx4n8gyXFOgq
OBsZtc3TMHGEfSg63F1szchyTV59alQasT2axkkkWgwUT/M3PIerj6MUKiHjw17n
vQw5UZpiKsQRZY8cPmWUcTZadYsMCrWnNuMDr4jxDq+a2AV8bLL95ybP1Xm6s7pE
fFrMHXUP6Hz6Wf8iId9wXQmTwOmSDDccp2yTQ2nqesGVg1MZywhc6hT0gtY0NO3y
12UpiMm+fxbr59++msh7iMhF+v39bmilKkD/UGF+LPJZJ5Wlb8tYmUIVZQfUv9xS
qm7C/EeHjSu8v8C+Qc42AS1LFofcLQKl3K9l7DGIFNSW1QGxJrgNB8sbSUqi6r3k
FT9txY8Y+eYBEkzv6rBtpeDTqlM+uUVvMzXyoCg1byqc7G1Im7Z1hgC5v1ebMtnC
r7OOtGdQ+Rvt2we1VtXS1WskAAWAFJK/vvkD6kQ9j5oXtjDGDuuDv2xCVJOjrgO5
8v6iHHTwpcO24lHkQl6Nvhe9IU3Fcmc2rF9+yUw3EGH4Yxi1yvOmI5NVHuKepG43
MXrCgRsuJ4s1c5rWrhJNVQ4fJlx1NRAqVxfSp0CGkGK+6NI5l891rqmptot9AJ0b
ryUraxaNrk1IiOXBEm1IIuGKx259FOPmKtlqE+IggfTKx7Ti+Kqs8NTkMy7bVCrx
M9Q9SYHIF2dUK+Zd4miVXo6zvSLeR24DffRH+17KWfNKSIEqTvp0pay929K1IcBE
izJHGZxWdoyUCSONaCouvsgOwB+hbS62eB7qyydl1D8fTeUB+I/zds24w4E3Hj58
6jaWywl6AveOWJjda7aqXqkqid17sZA1B9ZWoxdB60nMn1yArg+HbaI95ZuNod7u
oEsPUASveLD9GFCcZQbzRMMLBNjQdtFi8PMXAoz2nItHskr+4aZNCUMABvwvJc/I
UsRltUQklyZ5zV7vn7k77H2FgXLkgS4APhLVJuhag2pWsG/uUevkDkOgWgmqauQQ
AxTcNwJDgCWjBdzN1DMfjr/Cp5acJyr9jZ7OVQ7LU7V+MJDwtiS3nwjgwnWL/MKQ
t9xw8nAqJLLW6H8PCgaTMLAsjohAzjyIMhYjLsuv5i2xhijW8U3CUs78nhmmMPbd
HFNuMulmcqLQ07ZDqI7p9bQOnKcAU5H8G0aRy2Nv/pC604kk6M/xUVwpJiNPoJ8B
r+TZvF12U+ehqp86X/kB9NhjFtYBIXvvkRvlrNgvI5E2CSgNXbH747yGQnA8u9Pi
CI+LmXPe7SdqolCEMqX2E3uQxNKSrpv2QyGLGzPLDc3L+YPbboHwz5ZcppWBRBd6
oNLK2HgY1zB8BzHAQZnryQ9YgfH0JWPuW4CeVuUMiHsQaEtQiEZCck8CzJ+Hh9y1
GYZL0U2FaZRpjRSGPWRdktHOwyzZxQXOunUF6D+W35NeG9Zv9uFo/XSi0bH5vmkK
rRhMEWrSn27NtwCvmRwaepINCu+LI7uFqfTs0zYgC9HIr3beC0HFPqlLsU82P1HI
wKoD8wxOjJe5oej+30wIbjCGUnLkmmKJdKEira1M22RQy5/0jSxK9omA53K96xDh
cwIHGplFY7VulIMdHkV6XSynFzxeVmIsudetGOjvDm0V+eb6WgNBldkvw4I5iOeZ
KD0Bxhha+sZXw4Oe4NWF5Hq7Ifjq8uBPAHyei7SJwtO52+odT/qVowA2qZahUk76
1RLAfCod3VWq2419iITG66ojJcM5YG/S7eqX7ssNTrKu8NS1yuwisVeyrnX/LklZ
z1IIYj2SmPBlL5K6ULOap8GRAxPZHtSI34ojmPqogYHmPVO/WME2hQJORcF456Fs
qMQXyXYQ/bZCUZ1p8JiQYnYeP1z3S87pgDUkWlaAK1sfSpLjeAja2hY8ciw75i5c
7wrVNq6Q4NeyVLzQCi11hxF5AOxRKRjtY83ACq8+1dhpYmpISSIvtmsWbOzJL1eA
/jdSGpNxVo6W4fx2XL2rXQQuRDPjqbIhAXMpqGXHwSzPPuYZR65nukj7ovz+pvss
UXIfrcH6JwcMdmEJkMI6vKroMeyMXugjmXDFLGd1wSH9pJH9RDTlfvrvi7UFVzct
a1M2rlcXTyRKj5Lg1J8wCWagelDEGu3so21RvSNjYeh8O3W9YwhDAKikJbq1Tz6C
ueghWKriFpm7OcmxuhJLx/9SSj1Zv8RRb+/aH66mWsjxzMCC7Xfj1eou5gEOWNuj
vexLruN9RTMJkNjdjElWz8Sxkb0v14cx5OTn0OxpxERHvPlDDHxbKpZXil49jBhZ
YpJFmV7TmEneVVU69FjGxWANkzmu+CjuTBA1oFSF/e/1TvXjZXl3zUUbKTVeY/Nl
Mv3Lodcmv3YQ1RngvQi5E9d344HulXvWy0CDTOUG5PHYN6hDZ0xiz3ehkSNKQkZE
264k9gsrxFkw71jLeNsHzRSwxhDYjLmPlx/Q6dQtp9Q3yUyOvIP0vKcqJ+nxI40s
cTzh1yFDCH6SjJL7+FRlMvDCEZBgl41TJ2sp9d2GynQusY2x+K/1GwymT8uQ11KH
oz4GpqyNwjGVd9MZ8m7xxNfR91al8lUEjM65L/hYwRPvQzTeMxz/vTTMKviT0/Et
AFctTtEdVCHJK8TWuNePIByeFLh8Zk/COfvO+ITnKu7OKRSGua4WvUKJMQSwSOVs
RqM0sT2uVUiXedauHVCvVClvQ5FmVLr9mUrHT2RNl+pK/cgh8jX7tKX0VmvJS5bC
lIL6A5OxufT74y8QonGJViijVHVZurB2SaBHIYQXQJuwa4JWAkufn8xdk9EVlOzo
TGND4KnIZbgQj9+ZVkEOjvh+EtKnZAnhkWB4Ols2ACmeAZGRyzZM6Onz6dQ3/6Yt
RWhAwJU66miO1Fuegue4m43ebdb88NgEcW/Yj+M9Bhi03e291dezrtYVsIEb2eyb
fGZh423SwEbhDwvVJTPipZJTsB0wNH2mqtvVV40adpw0cjt8yt2DbmW1StyffSO7
TWmu15dUc8USKfTVoC1F2yc01rSIozTpJ89XVQkJi2KGOa6Q7Nsyau9QTpoQSugq
yPN++YyWgEhF6CLkYYN5WXodDYdCS5I2OQtYcwfERUzyZcF7yRP6gWaiDVk+0HZu
sNWT46WQ8ZeGptdUNC1Y0n8RI+30qAVaqyGhwkjMJtGxHVXKEvW9m8SQDjxeFyay
zM2gkUPsdk1eJI0wCzTjWGvKU86PyekIEAl1JRVmQ24WgWmno0NAL/vV8d5v5Pcj
wvbDMmrscXN4vzvGXWoD8a4CPcFqopsMMu6fd7jFbf3E/V5/UlyA77U3zK7q4O5D
dHT4JrxJsQMw6Cr1NTdcCip6xLObkoFBwQvD/OvJqIzg+xr4EAC+YzJmtDAd8Cv6
LJpo3hoGvw54Azz+1IdxZgPUVdHntr6n/6QmSemjUjhpFK++VnWBvnkvyLFZTrzj
xrVypk22u168xcOtZdRFlWz5RyJ/BrhcEog68C5DTO90ISuG7Mewbdu5lQcDhX34
t3fSKcoiaTlV1kbXJa8NPcFpRf6UlRqOsuAoSC3FeknYipu8iYa1rHw88Z7ICglY
sM8uVcRtnI9b8qeeKs1a+rq207BKkv9+KcRl7aiWK1AuTFzcDTAnmEsHfG/HddO7
y5ooPuxGq45ytlkXuNUKvgz/RqhdqIdvpCIHSoJ2hMKrGGTlVYynd3yaU8kKo9UW
gBVn4hard46I68wU8bYql1+j6eWOEmpHr/8hhjKU+xJcxMq7iwBUiZcfQwosRc9B
Q1n1sTgU/IROy/wWyfmnKB8hBNYz8xTjEi2p5K2+HEg2b0d5kXBk7DvTPkht5JQo
ou2crgycuDqgH906lrQUpA7j+PWwhf2jYXBGUr9H10cv9wiF2j3inyl3gbSrlwI6
Z/fIQh3D8QYPLC3BnpPmQhNHbVMyYmeDd7tioNfLPYEczSzp8J3MZe02nesEE+GS
I7dqGc1t/CdN2HXKd6kPSPZXgbsap3cnrDu1hYziaqBxz59jlXljSlD8uKkdReDr
RsH0N1rFKTkJpaeD0bGzJDRMzGPQRg8qgIfDRaxGU87cGvZn8kdsb4g4OUQtBhrv
teAa3gPuaHqlsx7VWiCFPmMw95MNeLgk4Oh4XTDQUjP2SUeHxIR88t/jnV1EnDIh
MdkXHwdYT9Yj2JZdYA2/Pvp4RZDeAxeGBBVQZVjxKi8oQ5lD0LQZ/2V6okx/ENe6
aYQSnm3fbrgaITrHI44T8FkzPP67obiMFxhcJUnEkk3jGe1IWy+oeuWEs7WNCeF5
038ipmEmiSfF+luT3gwc17uKp5WgAfcRuC3eY7btU8S7Dtkez1pNqPG4HgFZKa0R
6JFd7J06azWvpTd4lhEIRtNvvtCy/j/mzE3wRPLux5qRy4vDBs+4mB8E04a1mNzr
HrgX4UKcCi6+LOEzjB/wNiAfIA/TcZay3xD7MAl5H5ysik1lzHR2/HY+RATmqy7Y
ERzUA51ZSkhA2KalkFfv2rH9KuO3+Wph5El8/lVgMbyx9s4I51XQW6dEvRlR1pKc
4GE2osRvDPMZ15erk8hC6r0AiomE+k9UI/b+irIvP32n/mKdL/33tsTtsFUh8orv
nmTWh5tefxFBfD5FC/EGLoXtXAp/4mSupccjMgew437PGe1ERtZUJF1bgSH6mLhU
Dtunw9srTQg6d/Po/xSKvVFz9SSCj4MRJuqxBoUG+nbS+e68r/nambxR1Sz7QHx5
ul3g8yCSnq4e+A8dPTiewIFHpg0fNd8zDuoK1gPvYcPfKb5jwu9mx9/RSCHOetiO
dpZ885/6S+5FdcvsKRyZQnqvbEdojGfpXNqDQh9/Y386HQzMCvzmVUUNaeaSXJli
LPtbZwDz7qCERI7BWtLk0KuN82bKGBVvoF1R0CyGrwT15rCPqhfuJL4xrDq8iDUk
nbV7NPZZcUuGfjSC2ckSTTi2bhu3IMhYuWty5VrU2aYum1xHn6agRqmi+hr84O5h
pVW6GAk4+QcpZO4X6FqwIvz4IV9V4njL6QlpCbY21m/hzeK8jewOnoXo205a6Wsr
`protect END_PROTECTED
