`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGnTf9Q7cdA8zOO8gPywFW9WA06T12befFmE+Va1WZvGmwwZWKYL9S5+n/i5jfJL
frqkhW0CDxj6FmHqOUOl/XxMbW5QFbQh+fi6/pgUlVPWSOYResx1RaJQOgfeed/q
kX/63bN4RykrOK3y7I+V2rYRNbWnOc/GKoxXMcR/1z5YG4+duqiCd79qZSmGogL0
WBang/dJ6xKAWB9kCFu9GU0TmI2BrKkLvzeDwohRKQoT4pIEh6+x/W1YuAsU6c47
vnuL8Rqp4DuPDxxxZ7n7LxEwxggbhhl4NeG7r/vv3Rbz1In9aG7KeKZCww1JOcju
GaT597qrG30braDq9IyWKxFJ72xcqcjYLkBcW0jmpew/KG0i5oqP6TCVTvwCb8mD
5+qi/8JmR6ycaBwqR80qM+6Vpx2yC+445QsAzEkC1Mi9o5yVN8StMoAWfKUXHkMN
TseZLp+/7GC8tmEsQ9KsDb1ceJL5DedDvcpSW0/u/pP8RdWEDY4N+ZyysnQJo3Aq
AognhO9T5mtLudJPDaXBEZdOMA9ODPuuYZTavjN2gPhzyYfK1T3L/aPLs09oApXn
/FYdR9ebtRpxRB3KzxWtZT33BeM8VlVSstvU+X8QafSxPC7Obig6JFOnBtRok/m6
L+sQSYSsKk6tT+cCNrRfh6KGNVSeyOrIky7YHGnnbjAlau3isJwQG3tCPCQi8yYN
vu4dCXgtn5Kj0IyKbMDe6QtVYbNZ8M1b7N4RHL0yw95/lkROxk88Md9wcbJRMk72
ntiOWpuNFYBObNqsHht/PLFiiXg3rlniL4xMs9tqioh6Zqh2zYaJaL6X2yuMsyEQ
/2l6yp6FCo9zyZCW8sM6iccMiLq8vUq3FC8cKUmQPN9Z44c8jwlCaSCecHtvIwny
vVBcX07Pc/chNlDXtbhSLaWmoKvst5H2iD3eHRT0g0qugRGpS7aihrSYP71JdLHO
dt8tXJj9uejPsrsUUJa6mSB9DCEHMkhuDZUdgMzaWxlLFjIIpoWkgTAKHu2oMG0F
REcJxA9KLXDP7qHC+r8i+ZTodpMcY8Ljh1wSMpoU2qGXYd2zICxVar8K/GXSd5oJ
/Xix8B2MqHVsBNOW83TLeuuLr88tp6fTqA5tV6sf39poT8XkMAeO9a7RqE5oUHTq
yaw4yZXjaDcJTtTmIppTtqEs0LKns4c9dC0V1i2HRUltdEkLyTU+A8HTgfavkDfM
KFSXkJtt+aQo5bumbQfZynXUcS7mp7Dh2JxkmzkTdEK6pCOaj6nEu59kY68+R9Dv
haKnf1RcboiY5BohUXlmBH9Fm+qjdpPK+yyAb0poR9RjaP1A2hei+E7wB5Y8LSRg
UZWt41awdKNAUJC18EOEPv6KiMhD+GFiqdMb6yuXOwumMM9cJyGOOVG7rkCvVtQ1
aGg3GANCrt8wdPBsfrvx6Uf0CGrzUKK+5qGy08ORnNreLVgG4NlA41wqZMrbMz/1
XxhVeWRfOfSKcUS0Aw6RrL+Nms1ocOHu8VO/fhdsmjGwmysPogqG6rAy7tJjvxpa
CbwFHcV92TzymzPMNN24VfAb/6fijvShYTxkwF0m9XZDB0nt6+W9ERp0NBc9Rppt
I2B5jdCyf14SDCf3WFdxlyJDwMnWhfICYnufQ7oNPKtBa6Zl65GgY7zT2Wm2dgT2
l0KuJVhmxz6be3Cag/ZMBVqytZSCnb+yr2hYGEkaz1Ubsllwdc2jVOnUB5YpdJBS
MtF/d08z97ukNriXVb7OLiES/6s5dmpHQhxUkNEeDfPRlPrv4wqiSlcQ327zuHKT
0UROWhI4X6/9Vjt4EURkQ+HTp/ssWRqSIYWd8ELG+amI3LGKduLMjIcZcRccg2G6
nAJ8lL6Vx7sph4NPWHU0u5/kAIcjRUGV9gV7M7VVjFrYUSyFA78q2HNBb5V4+4vM
1ZfDAy1tjc8a+995jMVKOaDZVQ63MKBBysa9DPr9aWLWwpuQvVAhhqqeXw6fnMri
8OTS+d0YWIFdr65+/12jEBSycKOgM/r2BlreDwYZjMd8eY4Y6h0VWT50BIvSjQXk
ZHVdVmD3L9wQ04xXRVjITyF8vLqAniOGW2QsvmQ5EXe9NrmYRWq4lFVTuw9b0aX0
nm90bxgLA0R+/XCephhA3VKC7XttdTFIjS1CbmN2n/CMNGPFXEjb7YqxJcGrtvRM
o9v61UJqM4NXPVa4zkV34p6hZ4uAiW+4Plb7/7Av69aExO8Tc1MxFeYRteJHDsck
A3NTtpTaBG8jK7yIO4xl2aZwpG+x11RNaVA5aUPVgGYGfP95oS1n5Q4DCQ5gVCjU
5ySUgpFboNpKFIl4VM9mJ61oj8CR1uet3AxWNC7tllGIM7aaQ+TqtvG1jazjJSXn
WvkPybCtKn2Ue2PxV7BvWk/yvw2j+Jf0fQavLqTg/rymJRo6QrtoMIkq/fM3QTC+
plvRWUMb3JjNhDbqHiMV51+iJbHcatEyvj+EqOkbOjCOirViqgUo0pxygp32uBNZ
Q8ybp8ZDfgtooOQgRtuDEoaFIaT5WSU6DdmEJMgzTevOlvF4C2oIn6YGfZ35NKxb
re7c0OZycjG9My0vS1tsoag9FW/J6MfNCVC8bOTdt9HWkqhX6j3IuTnGh1cLQa4j
oses6+yNX0VCCu72f61GYsIolFww2/uuOoDP4DE6HMAo5LDSauyl6l4gp+8p5hLw
`protect END_PROTECTED
