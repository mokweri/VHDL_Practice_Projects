`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6A3ZGEqXlqmVNGT1xSYvB85CcnnuaG7ka7BMYHvudMQmnaslISKdJ3V1CJBPqEW
bLwiROQ3zOUXwGNtBL4qo4qanM/+d/kt7Kc9ZH1Y/xUHARpYjTYzSSW1HAGOX0gr
MoM21BQLb2B/bbQRar1Oq2xRxcQ18IyCvtI27ul/BRWcQVOO8MlGKup+lJzmMzkt
E+Of2+AWY4eb5bFyVQoXl3V12T33eEcjke2l+oIYGhbMk3FUpZ9YnZE6VkWMpZwL
65+nLAVH0rk/uBaGYUWYQx42xArj8x3uFVPfjGEEWqYDuIe3o/n0CJhB0cMpXelo
1sQWNwJalsReAtAahL6NLnMh1fQxeBSf72X/a74ESLFOt7E/cJEfFNm26LSaOLO9
q57r+G1fMd/5IWFkP3NXRqQDEDGiSTkzRgeTitclUARXQcduhmY34eXW3oBaj1lp
66nc2/R8C/lGAkaxRyAzXhEzps+6rgJl1X07UdISNKIjiw9fcIm32RkBCmmHjcxv
Aj0CCkzEcG2fG9n0atgaOm6PdUBUcqBJODtHfQh5ON5dFcs9kPYvZW2zWi1w41l3
P5qERtOsp7UPCEf2byaWbEE36qboOXleEjvGR9uFvCo0ERbS1Slfi9t3iT8hvVM2
dlyirhoV06Jq7YG0pBDowBm8W/n0csU9mWBrLRJXwtqugnjy895Xlr0PLKvXg4ZM
xWHoWA+T91reMJwRFwDVR9h/Lu1G/azqcsqCnEnLKZ61gmqQuXvZF8vsIk0NbeEp
7vzZEaEWbNhdDlrzCBrhqXYu0DB9P1KQKF3b2QtR2TK/hCx0WXxx+uKmcfeRmEte
8e+6k6rXKnN2wqmnPjNCc85L8GnMGnMmdP3ZNBr6bbBrYWG5eNPTwEbgmC+SxKL5
eYhK1994U8Fa6p+xAJ0NBs5fK2nhpDjJNQZjXRq10Fnh/2TmvNUlggeXc59x5J2G
4g8LLvh4U1Py1oADV42Mf+I6N+MccR9nbUI6d18/Hl6+yJyNQvjlNLhiceTyB8KI
HdEiQsjO9+oW95ROkoBBNDaC6iE5Oq8TsANQHmPgmCtgaTliwPT08oqdhaIpZMZL
70kxFAz6+cV2Rqn1WRhDmWaQUpre02QTS7nwbqrHI8O0xj6bgZWqg28GgkvcRSR3
v1fP3w5MIWmLZLFPud+8iIzDsD4iZ48oXP1LfaNCanUiGdnzx6fsNnM3m+giim73
76IfX24W+Q6FcFyStWvvHL4AMzuI/7hoUoS2EuTu1db0RNzP+ZzsIFoyQNZJa+m8
4pzgFavyHKaNWTTaQ/ghtUwHZW1QDId/oOGzQCJ33uvPgDR5fA9rhrckz65cw9Iv
ZVG+6AwSRjGV3On2j75Qc4K60tF00V3VOp27O2xSk3VQCCJ4RpcuX8wVBQFQmAW2
ft00gn+S2ZaOr7dXbyPqTbLbniqbR9p+X0gMowJeHgAOnjOpKP6XeUu7JrzK7QzI
PPcURrRLlO2g0nNwNLxOZsMGqkkgmHo1ns2pb6tjX2brkwDHueTduTJmBZQ88oZl
31x86V3JFqzbjRucn6U6ZeG5H2LXn6sK5y0t2y5hAOD0YxRQYDyo68ptKjCMG7cD
J6VbaXenh5/S4Ndufy0tPQ8SOtooT7Fy2o76yZmcx7F3bk/jszT6OP50NJSXncNj
mRpZud8ttHIvHlLvNLkx5zEAlDTAIkr2kKSNMz0sK5HDEiTyZ8ZTID/t+Wu0cq4r
jE4HqrVlJmoIRghylQArvGpIMRYR94HjHPksYtZMRWqUTnEeHymKFzi0RNmpxJaY
GkQZQFKHs9LAdZxUPrWxLMzCxmCTFEVuRefZ0ubNWtHEdN9GOoHlVwIjxK3Otb9m
jzT9yEeiUBNY8nCUMZ7tnawa5QksTjWXBEUMhT/vWYErxWMbMr2FzuQ8dNpWdvDo
q3M4qUd3ZqC4nwJs0KpTx93raN7GDy5k7UfJKSuJsK4nER4SU0IpXL7K/08qZ88g
fM9Q3ZCAB+wR7NdSLUoxz4J7+fc0pRGq21MLo5cjwOED9Hus0OIyJc8T1kpqKbYg
L8DfBvJAsDpXS/MmvjhoV7pIBd5jxoZTbW8qulvgLIhYxziSvgEIZ351Rq9UHG+n
mSF4db0ecJwxT1pxm9+xIi9XlHARfYGfgTFdfe6IUF6h52BzX3alzmQB6KCA/jbY
zVmkOXQ9tZx98AbUWTPOKru8qAtkT87e2utdA3sm4Zt5PVVvaXWjiK0VISiKS9H4
5iSeJBEZ9scwNOPb4aU6Crq2OUkwY0IuCKwn4tN7sTn9LbpOZEJNN5RIzT8P+r7V
exR2pPIPNzP2gYN0Y2BtSMpSyHsKeByeCkEAnVa+ryOpsc2dLJhfASQ6bc0H95c6
PtBDIzZMhy42vC/8JxBWm86pyIBVJqnbtq+R520NIwlod7PRRxTGxZLoEytsho1X
Ak9Vt/gQ1Gra3vf2TOfAy2QiUqYrucN1MAxY3u9XZGATP5rnFuhHi2e2GWUbNqRk
d5VrjX2Ba87y3nIcMAI7mJa6+8ZYjcSoNWCdm+fD9Eb1mfKCbGUs2dcVhHvG0qRL
VJYZbFiLNwOkADUa4YFwMIJ+jrHCQ3u55Iqrn3N65rU7FAGtoSfbnDq72qfHzTMb
o6XAimGsv22FPlOrvjrGF7yJ4+Iu5Zf3582JzC6D7aK8Q+TjEHTmiTbqYq3UeIRh
XFfR9dv14Hx79mUKzAlzpn4163gSdU58M4lALYTEYBT/m7gv1rukv5hlCAqoDpq+
Hs/SxyxQf6TLTPKsV2vBLCePtWLdpLHHuvBOzAeIsBIKugwy+I88jp/MAvl4a4L9
4TlKaDpTGihFZ6WfbdN5YQ5VOhlS8KC3skgJm/vovY5vMciHvgcNBI0/OeINZ/rx
wbFAQkJP/vebh66EYE3W7D2oqcJaIgO4yx9278QymR+Cno94sNGYhaKZaJI1wibL
ggh4lDzdK5Vol4ACtccLvlzFtJy1957Y/2Fimab85WcjrdDPDh6nFxeg5v14T2az
dUoQuHyxRzzkSa1atPUc99hDifLiSqupc2D+qKb5SpaHnerjt3B2q/0zAbeD/OlX
1TCtMLzy7FtzZH+ORczrYjkyjJsk+rjCMpJOi2fSr2zEbSvY9/G6sYyImYzrOihK
SbwqBEf+Z3uzZIug8ngg3Wx09XpAuoCVE2wrPMdv8pemIpm+Df2Oed/lGQrfXD54
hm0U+xZokz6HuBfoM84v8v5O6Z58Yn1EQRru1JsX/kf4LHksPBF3ZgHXBZODGEoT
jgS1JKLS1CLQrO4DOxX+XcbxQxR5qstbpZPZ+ar6uSlkyQuV5chxQQXdQJ/g8FFu
pMcQEWXY8FhZUo1TV11FvYaAzkZz5pV8letuIEBk2ObUXeW/QVfoQdGJ6lg/SAqV
+3o4ej2EVveYzBTcGL4oDE8rDDzz7MmPCYptwI0rWRiJjASP5coHHJ+GSQ6Jhjl7
UmfWy81n5LQ+3NTuAFc3PkO6nTC9GVl/3+ahnoyIA4f/swNdPctK92QwsLXJIcVu
AHc+43QFgGziRh8Mt86pIhtmLCn1vDYzohN5IMWTqWMNfiaQOVpHp2PlFvJTSy+t
cQSilO9Z5BCIkhoeHL6Y8Mf95GU4p7qho2izL1RQ3+emUy8tOV0mkJA4fWvzkmZe
TSlRbOEoesA/cty6/7Sahg==
`protect END_PROTECTED
