`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzhJmDuWC1hdRAimeth341UL2rIpLECkrOYvpcXBKfsVdvbvlQssVAB/jk3by/2x
p34O21ULbXGUz+Kg74AzTdCcNYstVmTv9jxc/P0o1Dz51e6C/k3/HEAKprooRhFf
ZhpO5aHQbG6L8j618KFP/KMZ4fb75Dvv5b5bxbFB6DKJyII/r2Z+SdLLB4byMXww
Uz+nipiFu4iWfu5Cu4NeofyCbJ2InnUdXu2GU2+SfS/ayeCs+dM3unVmSBEw6W1X
NJegORkJTheS//V1D16RdhUJ5udhhgJOm1OFP5Ev1uHmdGr4Ab8ULGfyvyFe3wQu
ZqR8OJ0M/jJKFVP0ijARY+/hRzFq0CDP2jdJVxXqgdolN6mJXZmWyLQqle0vJxrt
eZQ6k7SqiXw7uHQ0kBzg/ZxIeGjGRixcI/9QS4sj8bBtqNvibIF1Oxgc9jQ0vNIK
Ah4Qn8WLb3HhsOAiPej7YtLTzu207Zvw1yuJipTH2wXVU+T0bhv1pqwZALWReuG6
0Y5f5ktDIn5dz+W6cW9XStp6nlPzFoAOsRVoa7Y+w4i+mb5piSUHN7Rdt1iJBwsG
OguPP6EdrUvpk9Wa/YGSlEpOHJ7OuwWSZ2mwjBEXP/zryloDrVv3gIG1uSldP9JC
dNgKI2S1FjyRGybbaxv1NeUJsbYe5ltksEKtWFUZ0rOruA07V8jeDWLn7PN/x3Mm
CpGRDV0gaa0syywQVc5bNdPSxkRh1vS3NP36WcLy6A9h6WfQvG7krom8cIdK3SNG
FrKMXH3/tiFq0HBt5Hnvb9PJmpTTQiBX6OEbRMcUwivbuMIWoMT7TQxxFS0eU28m
COKtC1DO1x0zBA88++fKP8HzclV9/PGW6WBvKfbAQie/E7qfX48y1Svor/MsRgkd
Aj9J1TuD+ryoNT0UGlVcmuCgu5/B2XO6wDf9C4VLEyHg/CDAtFOt/88/SmZXzuoX
Zc80QrP4+EguxkAv90vNRBIYk+uefEb9DWqCXswn89iV0/jCfjweNseiEqw9gORK
0uNTi1RMi+yHgULw/gXykMWVmbQig1Dea40VeqKvE7aFdE1+mKS0NRaAfRq5eD/b
CWUwZr/piJEj3zRZyzh1C25kHSDpvCkDnITJNnp4RMBzdWkgotUIfoqR/6Ap7t4t
ZDQ7wP74FzK0VTZqYk37GmTgK2/juFHnS8zH2AkMYubFnJBy/47Qy61oMFYJTkNb
VamC0HQLg7UmbsIaAsqqQn9aVAIQmr/1riJYcxa1fMs=
`protect END_PROTECTED
