`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
deJ6wsaD4oWBcHjNAa71uawlFO/qntNnPH8XRaPYeioLQj5j5vvrbB9shPdPZSz8
ySG9XuS/n5sKse+IFCyI2oLNRhEvARmv8SChPriHzkLBdA83RBVs6nJoj0oE/khP
uH3MS6aGHmylsP50c0085APBRyg8N5WrkN6g0GMeYH1b3+Awtznux8Pw9bzwqJhB
8w7T/uZdvArWPBo3ngp3edUL9bbh2z9lp5a/WLEqNiusxDHWEicBFESCF/M4V7+a
DCXwkiCUfwv/SShh+ZGFXwkQ63QWStgbN9D+HrBh5uWoYksC3BvmL5drNZorNd/N
esZOJarez5AAVROLZczR9EMkpWSTW9Cg5KY6IDwxCmCUXObCBEZtj8bkNCKm0r7Y
ZN+LprVTHJ8+YBBNi1aEFOxAVy2w9e6lZ4ktThRWVBnRTp6FEU0UCyCQ2Nc9vXIq
OTcuGUlqM51/vokyrLnK6+pnoXVKMEgvnBpzFXG9pGwm9q2sXrXIiZwbFniZhtTZ
phdkRrmuwNexr7sM3zTeNEfnpv72YIjfJxp8RmhPXQDx3n8sc+ndJrjqpFPx10Yf
XGwYaPFDFiucgqhlD7Pvty492/4xX340za+QQ9bITuMTMvZd6fSjolteJzQzyJOs
us1J3t7tjlkWshdHJTGI3BToVQ7xW78xMwPAlLZP9vB8qcjHaH+zcWOaq3Y7DNqG
0QUdH4nhEH2UXREGmCu/ryMrguyotMpCYv7OtAoZM6A/73D5jc92VWxSBThqDZN8
sxTnlrZ3osOr4m02Db8urwfKM4edykBMbAPiRYyoHazi3Xr2f5cyLOFnqBhLR5tV
EQq5BfDd8IgN58Mbdro+dUTf8ZomrA0nOP5y2eqBy6QPROWOrjvRoFUOgWA8DiMB
vp6lHNpz2oiJS2NocVdd4gL4E2grU6UlOHmoufoocRvNPkargatQM/cd8i1Yxt4Q
XodYsI1zzpkR/JQbKTPkiGB1UJ1dkbBFikiUbH8272D18ZbDuhPjZBfmZsFka/iH
FUOTzUB9vETgMMu1gOkEIK7d0+JYDUNaqC7a2sRIjl1E3BlktfrgQplVfmiLP4hI
`protect END_PROTECTED
