`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESV6xsaxBgsh5PQdd8+Z+Q/0ZsaB24/KFHaWVHMUmoc5yyOTC25hJcYvWVEjvwTG
bkIZA+phTwLB35iTaVsG5XfDTYFmG8/FasDTyrVx/G4o63iMsU8Sc6ktPnn7DLSW
3T/AiYH7bgPABWvmYgMG5d49tTagw/dgJYNl7DE9nrXfV2iP2ZgCoOHi7gZKrYFR
jE2ioJ4/eVmFJhNB3Lu4WY9HwEWYbsbtnqzn5Y6wAe/Nenf+/3mmVU8mPJWxbAzE
aoOjEJzQUdok/AiabPAO65xzSGR5clxgzHYzyWs42CMXlMFais5I2rF/9rPz74T6
Xz3xj+F0452mo5WgilNmc2NjQCCmROn6LZZ3UvYpOjql+r3Rla9SwTslC7IN3YR7
cP1kyMVuZIP6dVQdpQrPmikhQI6uwQ13WeGp5n4r675Az4oaz59zZeWV0MX6OA12
jjMbsbLjCJsRgqbzoGeg07/HnggmwjLnWcvQyBGleXurOi4vi+mZo0w6kaLk9Qk8
j4n3Xf5Q1ApBSOrHp4W5GjfG6zsho/roklup530AzpyKucp4ppzOEaRYOQjoAU2H
+fascdTXM3IInkTCmINWLgT7zwuF8rULFhCcTCactTGe2gjo10Ot5sfMSceCLymA
MwSu7YsrAEfKiZWXrVGkGgUzT03Kbc0ESpm0gD5aXlRLcnK3iPS48b/XLyj6J8+x
hosmu1UpzDhCYZFxIuSJOCvQOPne8xMKHBNVtj6FfwueQ/9W5LKZd97LbkSbJ9gX
EG43TLtecT0/k/ZZRi9QbJ2Aj/ABY5urQI2VtAYxVVGRueN4I+/zxLeYM9hWHhft
BK6I/nDnXDujiiUUbkdn9dgMqCV2N66NA/yt62W3TpItZgCKbXMscJ0wjSQV+Mbo
A5eYcaOMT4kFhe6SfydT14RWYgs5hAGPOkiaK6q2Zwin45VYyJsk24sWneS7WF/A
MHU42WTVvUa5J51b33XrPs/RydNuGvtC93mm3av+8OYi9N2Ix7eJovxWtlY1sJu4
5FbxCMfM40mWaGTnyjO0wnEVQ/yj3UkbUtqUNrZbSpKT+nyadfz6WXz5ygcGg1Ml
6cnCcAJXILJl799uM5PypfGGnaJB1xFIIlGTQ5P8jPjnGot+LkiF4KiB5KhI8C4h
ILPEqnF016BmFhbiP1WYGugj/afD2zmzB2mkN6L2llalnXVJ7kuCaYJkMd7799d0
BfvVfAHHCFndmG6RMKLnoOhn7TPaCBXfwfy8BLXvd+rkYBhK/l+gSzOzaMZ8Zklr
rVABr7Ym/PNUKwfIS1zeNDPOrrcOW1cj/yMGmifEQyECpSldCX/Aleuslh4Od32A
5M5fgTOFtsmK1jzQ2FbWKRbRWLOWAw9RCRiISDlvUpCfbchHv9VOqhEuoC8IhwZ1
riwyiH/OGxgneInQy0bDPuHz/v+SBYlQdNnD+2C2DIhonL6khe15gzc7/7+yxRVb
Or/Hxv8Q0ePqJW+4DBIRy4SDkiCs4EaUquWL9tcAYbOLkdPjRW6GGo+CUyMhUqj3
iTZSD3HcaxEjbdKkBa9p4Z0+5uBFxpef77get8Rk2XmumEqJLVf+ikxxm8Xnj8jY
odm/QRzRaWQB2LJhZxtp6xDHPukjFMrm5gX/j5GIByXar9GiF5NhndUxgptLy0fr
jYNVqkvT45lpKJy9Grfg78nk0YDUmJJsyd4sTD2VWHYdduw0ItTdTi/JSXs411iT
SQ6J3BhjCFiTqp011TGi+lwTJY44COfaWZ7wCh1KjolZyLdCn9kChpMSZfP63S4r
ByrWpHqC8Exo1GEaavLJ1q1M1ffv7h1LqNN7rjPGonT9y0WdENeupaUqIKL8QGTi
yvv1QNwNjjtPLFRmq9mf6yPez4kBXCK+9il+q644ubWDOBKIB+kq6hOyom8OXOcL
eHR6BeTHiJUKEJMEGPUIqjR98xjo+IptXqtabZcUXuorWv9Zor1nB2GmTIfLpxZM
rNWUGkbMsxUrJXLE2HaWlPiJP6NiXOoZf8ovJcE+vw4D6Q2ddp3RvSA1i6GqFm/9
6SGDvlMfcnspO3HC1lcFa/0PCBqJEjALzMrlp5OVU9aBlW6fj+JFSoyZsfh/vCKW
mZmTzTK7KZXmr+GxQhVVMuXZ0G2W8wM8UtWxg6V9MKSLhA85u4ZCxyea8hdT1ZRf
EDcg2CzZeU8pt7l+6IV+1W/KuuZ5J5doIQu+bMaiIl80b1j9qd22lWFfTe0InwCX
o2R51vWkT3opp9Z//IhrCol2IncJ3+CdV+3ZOTh1zRljCs1dOUr3xIfnpibJGbn2
exTzOhvW6Ch/Gy1Cj+Ist6AFPdw4/Jp+dA4yAB3gOEpy+5jKaK+N/Is4f1qGOaDd
wU1yb+OPFKC8+E7uTNiTYVVYwEuFNn8LUtBL5dysbiLiYoVYUl1huhyq4NzIF1LH
9eDM5uhsdJ6M6v8g/1c9PoFmaBhbXKKkRU6HKQORlO87n9XdSVznOAOw16J5XG73
8h5pCjjI/7BTwjDz/mY9X3+YBj3+kh1I/oW/ba5TjIm2+A5z0CywSlLMjrtMcwZC
7Tyge3k8bW2/NLOpABOb1r1dqUGR17WBcOEsKBnQsaqoT4tW4UeODhi6jEqG86iH
Avo4+bUQLGW+KdoCw/xd8iQH1cPmf6Om1K7F9PQ2PnnJKjH5M3052DHh0rIkzrg6
/B8wVB8GYqJBG0FeIRBcwakha6Bcq8RqLkFdFaEjRScNg1g1EjYa+qcwvdzwdMQh
+hH/X7X/dL7GiIPm/0ea1zNoPKETG0o9IUhCTrdmQuF1wosZ40uymWy8YAFdI9/6
zqMFIfg8EtMm15EkimsZZ31Mm8ProFY81WwXLpaXN1rTLiHFjHN8wT+A9v7vJB86
sHBhsCuam57wWj/awmwXYbAaIO6Ah9GTKGpwQSyy2XsAjMHoAtPQCvWo5RQATUZP
QIiT3EOx4Q7f8QLmMmdHcuM1lZc6Y/PLlRDNaMqbtJKE1VAY4Hthsjmgxp89lDm4
zRNuY4o2zyRLo1EoGS2oLyZ89IWcjpQA4Pu1IUZL7elIJnEvsO8e92qbsrve6Ggb
ZVouFuew7ZT7+TAHIny4AORl/grogeRx0YhVo8BkA68jHJCmkSkwhD/UYFeh1W7s
LF68QJIsvNEC4ZsJsxt1Aft8e5zjfrbiVxNPpyZO6NM+YrWaY/LG7ZBSWN/QXjNX
fceSha38BalUU7Jt4zHuzOltrFKOicO6yEwLBHQPaZCdi/1lo0QJ6A7Gxbwd/yjf
weWiQTH/bHv9kIAcJikgCroRnB5M6qKrrCycB/YDdYCO49fbETLkazeUcNXpwEHR
bNk3+4hZGIqft/FWmqzCH9qrEFQMg2VcDpMCuZ7wa61wXPysds0nxhwlWZcNv9Jy
GQi2DLKHOuzrQ7YTccZuMU50fX2Q36E+NR7iM0sPAuhm4v+iKngfoM0QIkrQWnkq
KCvPlwcG5b6OUiC8TAh948s7Oyhp99pQC0ymJdJk6Qbq23J2uj5Ww9kYb0EvB92T
P2x/Pfll/QOPUc/fYDtSxXP+8oquPlhDk0CQAdQuYBwdVEJLbAIGTHkn6Z3q8Jiu
jzkj68Bse1/iywD3XnSjRGY8t0NM7GRR2dTCelHwBamNsuZJ9Pcf1sS7IkB0uFFj
x/TjjgAHZGTtgDL2NxjuMfZKLktqlZcGK47jZ1UAKkQCsr8NdVG5Q8w7zixTEMh0
/VURPFe5S7qPHLcnwyWry/jwCWuN7RVi7Y/lg1X72znW8SSzQW+Vsc3yUiPoxj5Q
cgNlZ4EMjBOE0sd2BXvm+gOb+hG8I4KPeAXZNrEYRHsBtKhKBgdOv1fO642a01YS
9+LlsCd8XTQi/K7TLfw5vzR7AJSFdFAbDMICwxCDWh2W75IVTL22ORQV7GOGf+Q1
CF42WMjX8fbKyPlpfP53vZVayVAkgo/wSt9wOORCxY54Ywl5vrq0DAuQFUNv90+B
lXZUpHP3tpKLWVPXrvNGpGDQtxLZ3YHdovbSVT+QI8SUgtWZ/owI6p4OCwqHQNcW
qj0RCoTwy6j1saD/83zvIU+K8VJ/jVxCq3aNCVqq+jRrLOWrt6kACNinwvPpCFXc
MRmxMlX/t6CanktiPtKjx/rAPoGu6o7gDiISvk2EPrVA/J1YtVwrbBPFrIW9OOcx
OZlkvALs+bazV5WhWESWbgXZqgrdsmmyZ6hQayHZIywZyvEP+DNzYIRd5DFRJN8f
GMW2tjMiMa+8ivyDRvYz3sDGH7WUuiSecipMFlpGafUoSD5id7F1f/8n8HwM2qzd
cbjPWkjDBZyvjd8a+LpyLVCukCLs8dRerfLN5bI9rE3iqlR0I9wJChDs9rhoPbEn
ZXWlCu1LBkKmWxzt7Aa1F+1EO/7Mt3IVJ2YfufBc+fRZhlIjtyn8SNDdXv1FpK+/
irlh2HXVjeMDK79N5MgLbn4gRKdTJrQb9uV8AQ2ZQ3h/gSA2ejxLsRlYL48/KG73
GqmzpIL0n9772tCtJ1vUMsp5upBZlxTJCFpJZvcTY+k5/FuA6lH1XxIlN//E7FQh
MmpgZfgKP5ub+wJwf/3bJ7JirzeDof+mDhz1IpV+lqILNlJhavqD9BLtoOIC5iIk
ud9K9cvZURAuhOfGdyhucb/SUGRXdLxvw0p2YVaIKWrfIhU6O5VTHRAw/lxs70W6
tQNDuDUgYy3Im4mz1I5cnRX/rz8tOqV3gonIeHHAypA2jnum8378XkN+6vcEzX/0
awugKx+xl/LcDOVxUkfp8CwY3n1tRWex292Y4neDmwI2eq+bN/Iln874QCwYvPLR
L33U+GSQr4OgpI3qEzhpHgMK3YE4GMa1R1l4S06Xm+JIE3gpxfO8RshhNW8FEtdU
NLawdc/nxM24ZY9k8yB5GI1Xail6VLl2mAsNyxN2thuXTXxeniVijQTzYiF5iYyE
mCi5Sf+JYJw45+00VA18IMQEcCKb23GzkHtG0czfkU6+hUrgQ235O1wn7VJbKbPv
JsjteukJ4ipPIUeoJIQuaGgWEtdaUC6PR6wGVEj+L0RZlBXAB9n75K2mQ2RGI+Eg
lFuL7bQND1yhvwutCM8xziHh+FiQNlGsIfuf0xOxoUCBdLw5qCaB0jj60WsTMWeC
41UcTlqfOHtU084cFSBNVXtZ6kQ66dfChnE7odaHOBiVehjMrZ9FPLUPhLH4oh3H
bMeqA9v9xDORLJhP/D0UJnB8rOhZvNUeMtJIP73Pi3Y1CBV3DjoE/IqJzwlVc+TW
6x94d/XvMdCv9hCVLkuGTMVeGhoViJYIdxDYEfreKGQ9PyxgjmhxBKvzh3p6lKUB
gHnt2w1B4WBm2uwO+NSwaZbpem0NGyF/Ygo4r9NvC1tgbdR9LRB7io5/tFRjy1sI
/yFttAU54DGPavABUeHNTojR0H38ZknkTvJ1UZTN9DBQKnXGCh2hDs9SQwSFO7Zf
z4pOUJFVTl2QPnCxGQ7xjW6K2E50QMWTPJAg49xXMQqdg1mdozHQvCQ1TLUnjvWo
MP8/VQP9l5JXhO4XjrY6gXJjcLoyXgrQH8eUhMPvcHcWx9x+pT95g9rff11MOCBv
cGpqH1+f1uTHbls7/LMyxwD1jnYxr4GLcf42ntdtUrSRAZuNYV/awZIJWLanYFaB
FHJUSdHhlG+fPa5GQCVZSC/V5YZdxKH27xr8wIIzyY67yIujpo13/InwB3ttDK9u
hGssZ8iwK+SvUqJeCAXOGpqR7eDza6ToOw4/jf4Bd6CeFDjqNnIAi2yV/j6k8+3J
7/c6RJxpgIZaU3cOiE30SUxazn9LuCQ2cIQCBpM6ZPIn6k62/FeQLTxs+RO0kWUY
1RGtxow77U3KZnliWg78EzGmEZYTBoLnS0GETW/R0I8socuSvHvaruysI2TrOLAT
B2dp6OOUv+QMDPkmiRZuemUwYowIf0uVcEFNrU/Q8NQ1MftnUo54y+kdvJdyJEti
G00t4kTVIURMwl9yYna1CyWBVoD9OA6fhQa+TQhec68ICsjz41u230sSBKElG6Xu
M2Ep+PWQQ6r2Ma+nWt7czVqHIafGMNGhAO99HTbqdx5bKzJfkJIE1AFPUYZKFC0x
5+lZlfogZzvfpaYp7ZG+URXS0n7ZgRPnlYMQktw4DxISGJRUXdDWyYUc8satilYu
I38ZomsfdvV2GGEOSO50OwnVQBE1/P3amiRBl/Hs8JhtCZIAnnYvrYsLITBQtC/x
/UpNesF+q+E9hivxyhiLl04W+m1rIQOGNiaZJySt1Q68HA5gBCGo4xdu9VwxFQY3
LEezrszqaJ1N1TBks3ElHbMDLnGCbMqXVCm/URLTsVdb+De9JmcCHNhxdH9s7aMP
xlXHXwxpm7+9SLeJ0CgcYvvcrZYaed0Qkyt7uTuNmfEUydm8EHv55WhoqyKkDlB4
C/1u2508NTGuA83yelGjOHH98qLPV1UjJaIEcHh9ooQ6UzDSqNPxRTHG+BVhMR/1
JJCG9U4R0gnwvoleSqE40fPfuG5m0kEOkTYT5TabhuFX57BDiyt0E54Goem1bYKV
7TSCdyc4/2L+87vRe6ti9eHJWRVhEfkJirBqA1Du/1sdc5Kj79e8OBmkyq0ZBW/v
yN7m7IdhQcGkE3Rn+27ZmSAN+vJNXlxs+dnVtqeqmpP26dsqcHCiMCRLSczw8hZ+
qN65hXUIDCy8YLra9gNqOZ55BnMyM2utoCgF1/GSIUQi6EV9rZv3Qt/TDF+238eh
ErPzrN8zxfKuOZ5KLghySfz7Mn2hkN125M2nMjAlKNStGf9xhFnrTlP7cxw1DxAG
bOjSHfQoKnh0ZWfTcvvaGMSTosw2G887i78VAY7BCEh7N7wBbkZ8QeIkO3jPMosn
NkIW0vKTpw5E836S28bwJxFO8c6MennVaRjBmLde7WkyUx3WnJ4XLJdFgY2OsEgH
cvf/xCunb5TNOJj+6nT1HZk9QyPVuNtQYY6zsC2yDT5BSwMMwskN+KrgDb9rmVvG
TlwcoRsjrskTBbhBLRCbBHxOfFbcVH9KcnK6V7aUQjsdhzA2L9/BdsqkXXG6wlde
DEkbktlFuMpNVRNr2V8PXFsSFKSnr6t58A5xSuCcKpTVEkLzivpCc50PlB8U8Prt
QUekj7nsc6M8DFYSwbjFcEW7gmJrX2UYj7bqNG8ry66w7FjHGV9wF/A7CatLHO1w
rOranQkEizSEVrQ25Up1qgUCcnsd956q/JPMSj/SS45a/1cNbdlBn4z5dqu9akbR
5UkXoN8JthE+gODCu+j7DzqnfCefBFQwIoVyVHwAsazt8d4WPwPN8MDJe3TkpKW9
tyqboRieHjrvCEVQU4hMjkwucvIubMJ4DnsfIXEOLVtF8hIMIv0H86ZXTpk5PiZa
POGhY61L2lx6rFBxkYtCeURBEmqMIVAZ1i28hYCPLJcS5/TS7uPyVG5eRzphog78
Ejya0Hv5bIFQ1u68e4V1RRfFVKvU6++ZL5oAXqW+DU3BaqtYfwaDok3MhgwUg08F
Mc64R5EHh9njrSOAdQUHPfhSXusMc/Ymhf1QvHelGruO7YBEfsdc3uhXTy59kL6q
JpCuNhpfC8W3xp0k2MJdjaKzyDTDigSbzLbH6S48JX2ZNUJVEsJlnF9M8m/RlEDV
o/a5vSIn0/pVZ5SBp+O5L8/6i2V10VSdpZVnFiBwsIhTAo79Qp2WWOGZRHvOcffW
3WYZXl8MWO0Z2EN9doSPRokmYquIz/pIpiVCDSGP5DIYuHYoVxZIxM8OVZ3ePSTb
kBcQQmRf0y20hVHw4+TMMJkWhLBmRT6jUFBfMDdjWsrJ8DE19yXKr/iixieG1PZZ
9M58Nk3hFrV89ZZfZoR40bsLoAOKEzI3bDm0FArUF4AJXc3ZT3TP9jmGP/Khi29Y
VTZbsBHLUyoZjMOXe2aXk8SSOyUEB2V/MepzTn9VRquASreVszOyrFpamu1FE+M2
GnQBU6FHtAZ2FDAtWAAggnZaucRmWDaTcNvKtXi1iBUCr12NMFioZ2L6m7R/FsSf
jXjr446m2gt4yKsrmEaKIIQJeTGpvOEL5cr5RScy+cg5yYjhn6k0im02Thmr5fpB
NjY2wD04yBSkFZCkbiQ/cNtnRLYZkglFv4LRWIrLykDTwkeBir0+yD+O6BVkD+3R
tgkVCf5QwtcbhWiwJJljun4gcf5c8K4Ud3bjTfbxX9oFQnQTlamcYEC51uBWfJqE
hZvQyldNdiaXnlZJQYMAbr7v7OBIMcRebFx4Z54mXAa8XLC9l2DO5wCyVJl8AsLj
Grdmnbvf2WRqm7qFc7rfqNxnlDSIY5YOGkfNJ5B2ldvkLpP5EEqKG8etFmUkWLpt
cMOXAzTw+Wewipk/kF2a/Y1/NKlBH1alUluDnAZuFFgbF7h9q0djhf3P6WjJsxr3
X9gvL6Linne1STcdFDoOY86ID9U6oL1ZOsQHE5jR9AVVDPiP2W3OdWELXn+M24YX
WqKzNucrQmRBMZ/b80HBs4bFyzBUVPS8A580GbBrBo7zUmMxBnBz8a2RsqRBapuZ
10Hg4bFApxL53JwSWn2wapjL/5LMkEbHmENmB9jowmZXk5S9w9hZAcOHM+laKrur
o1RdxKFQzgA3MlWHs0v19R9Ccnm3pBQpLfEcp1tWrPeOVusdEZzF1JY50pYi+8G5
GNQR+xQfb4OVuATDaXcZ5KZCeVzrQix+YW8g9ZZd9cHk5W7oz4380cvMC0EL0Axf
FwnqOhA40JKI7OoDYhYCtZrx4dgFx3Zi4EUbYmyggrDu5xxfyB1ChmrgpDuYxd9K
vtsbg8OrV0xE3KT8Dx3R7yySLa345lWlM1pmxE1lBA8OdSXkMXIDGU0Jhu7YvDum
VfN34RAQfgqJsIUtq3momZfA/IVySV7hTQdgu6nv36LVs8qHI5j2GcXyaL0ZA2Sm
EmPTRb0RDXuaEb3Wmchj/0Jfd5LeCqx8nEQL6qLX/9UCyrQr983Ybslrj6HiUXvQ
/vC5ozk/9TB7w+Th/+jfq0zGcO7g8WGcZxI1Het/s4CqSOwU3zIIiZicxd8CwiyO
CIlWwa89QTDNT/blrMOB4pry+FGev9bbttopxa5/qCcce+5jmdsg5OOoGHSMASLg
I6uOQNWN3MI9O4FYkvVFbNDOFPbdyHRi2t23JyHuwjtGxJLersjgMg3rEohoBoVT
AVb7LK2DoFXK0JQ0bs29I2GAnIr0zHYkHWlWGIvI/mQwduo5bRFujERw9PxEYkQg
chD48UoauYrYdG87mZN3OD2zSGs2IbiSt/upC6qUTM/Al+xJLOVcdq1XlGfzs3pj
5nUZ9j8UZieArMYMfeTO1SIooVQ3CWuoNwSWTyAq9a2pct3XyTMn6ms3DZY71apW
EXUSnZefbdkXUzJlBEiaY1PUiVWIrFDkN3iZfbAT7GBvKwpeXcSLbb64fL3hp6FB
fN4KEDOoKo14u+UAGZ8g2H8F3pXNcyqm7JhMSV8njgPuL+tczvtteZle7/mElNos
y1chcGNWMTC1qvIzRdPLBPvMIssV+CnnvUlp0pw3ZOvi2/Sakrk+aUJJclSnIT+/
X5sStV/lJlyTM5ait1WE+swQuLRsboqrLHniTKP1nP+Etc12vXL+2MQqrWKXKv7b
eySoaFWYIUL0L35+N4oxV4rxjnovghGA1NWx6gksZ4nySIrxevH3Np9+Ugnyy/mg
G6w5/fYMrXjQXatfYgPh2HDuOUoW5PY5IpAbOc4/lNoDIeX4VqDXOzsvK2TlBMJS
kJTuMBcCKCNtrqqRLdNsWZN9HwkpTe0ve40Wd7mN7MBTxPDcnAf5hasghf04S2Hf
hH5ebTuSliwOwwnuQv9tkKonRvZal16EnK2Cme6NMM7zy+yy9HKL/k7GwQ1QIGJx
BZGUlb2ELTJakmuTiN1JWmsutiaoyR+YuJ2W4O3NNZjzpHcapJmSY/Ru/oP3tjdg
Vb8BGI5Lfwr/5mbIhGqSZP/u7/RGbhVUxL72luiI29gggbXydQl1myujinQ/tj1+
FtbT4VkCP9+Aexyb6PShwKAU78tl2dKs/lRc1vFRfBAWjWPIEkjhkXR/IAYVfK7B
ZbmUmzLjXns1z6ipUAgiVnWfKsv0JqSkom0xYrsoNzsDJ3si7fu3lSZAGNaiHk2F
9KB+AbZyD7U5T+dgR7gLOoY/Nn4ykHiIpqsLSlg5b53f+aWFe9TbqFj2NyA+G3Nk
0VfaSebP47R/rX0QzQXY8WnvdvCrmeP8K9nnch9MAIiKjQoDb4Sms2uTVunBM9Ms
Qhnm+/79S+drbOTgiy5K9w5E1Wgpv/n+0dpFqQ5JcThEqQkrhcLilj7PKbHWt6N/
7uhKqJ2x6qI/pDLHjQoejmamgGMrWdoKOMqfVQbe086EHPnz+5ENK4xoZK8CcYOf
6DxFFiD8VTFQv+IMS71gIef+EpM7iLDu3o48Z2IhxtlfRJA0+SeOV7Lr1pz00NIH
46p91L3ZG/I8a+yRKDv4gsPuH+xdgVA3zAFkdPOR88y8/KtzzDlgy62f9/RQ0fDT
Hbb3/x28vec4dHybLSV8R3h7Yqla71WRxIlxsmxzxtiCZZki8lwYVzmUrED5X/Ve
TpSbf4eB0kDntqhG7R0vRzIWxLsynkrNB/AEHYqSK8LTyvHWGXKPMvb99rlWjZso
MK8ip6MppziuPPnEcVjVF2/A/yekHNvnNOnyuUlXi1Xsre7dWfE9XhU06xClE22u
BfHJPeYi1ZFc6RH95vzxV9RqXdEXVYPR9l3bp7zYv8SyhrI+uEU4yV0odKCln9Tz
ikGXyHkVjwSw02wUlCCSL1FFomStCikbCaPfldkUOYu8UMz2JMIeeAlcPDucVV0e
nE//H2oKIMwOUMULsPNQRiThANKm/PrKeN2UfboCbevSS7omYbPB20jma0M+1aye
K54RJSKu2tgkI5QKN4B/inxDogRAljWEM1Xyng5CCHlXO7hR2swzMxgs7PvKLfeK
4Vlb/Ap7hx0WVXAwKDWZCa3pVZ2tETeE0GUlEv/vAyZeGHF26xDSOoUFU6OMge5f
wuqpwfh4KgQwVbpqY/Y/KorsqcEsETXF8wOo2fY6gzPkEHR5XZGUTBChoscUbgCM
tZS2pyQGit64zOxXaMQDnsTrsx+IvrLii0Q4IQdHHGBM9sBXd/CfBpP+fuCmK+NQ
GUHRH3b/9SxeqbOQFNd7qPVG8l5ST0UGvXKJWAM5X18DoQeltc4WrXd/RbDrbe3E
IlL1HOUAD+OhaIeKl7zDgccJTiw6KV+kIMQhYoHAGr17wgUZIfKfA6NiwJ7gNeQH
urNDOarutrok74ao68ps/PYzVxkqplS0UvOXiWXFCbiEviQmbv1Z91M67GbTUL1P
1aP//hSjORoMDW+c2xox3rI+2k9prkEU9HTitfTATK+i3++DYShl5bh89TvMEBeT
Ro8b1Bncp4AbtFsj3ceJ17mPv4ChWEQjdRWuwNwZ0hcd/ydw7PaSCPxWKgz7qPXL
2xYInZhqxgw1DmkJSxxVZypQK+yw0WRfWqWmma0KxjRr04tfpUDleBJQcQ068ucO
xrOZ4L4rVQXkKlOgOyxgZ9TBzHZPWCJe3mGGxC0YdM9WKIkT0pF9WMrkRbs65T2D
AuLiwsqJslzMuzJGx4ZAvAByojzTCEnm2sw6BgqmYywhTBMrcgTkz41PTHtD9moJ
U7Tvo0XAabD06L4Swz2QE2reGY6jlfNGTFx9NdI/hGuffRimPUY6BYEtUCSTwA4Q
/wOMZk7hOGTRS0fRNemtQZaaj3grtLmL71vuWsIDkmahdAZgp7xY/kUD2PN/v4Y6
4YeEKPvjoCHr4Iy0FawsvDWBE/IfpSwkZr46KZIb72KOENqnn5NxWsbR+CqDXqZt
KvS5Buj92JecO1xA/ir/ccdfKozLcV80dXHQIbt5b4rzWLwJF6zRqI9G0ZYn4hgq
WRx+ER8ejpXpXgX3lQkq4NCXFiFX988p1MgRBZpilF564GmBhthF2qbsEjHhL/VK
z0fBSu+er1y1WdLAUqeV81LYsWFprfuVF4ANHxnHEy4Asjc0TgxOUbwqunKaFRyt
42ox+WHFiZ6Gjz8Pt/kW7ooYFW2rwuNukhrMFouS6JF0xL3nxWB0d/2vzA+i/cWP
2vrjgEFpwQkLuWNsDceEr4SDL1rAuWjHsCicUHPb5DQjZGSUV6yiXoYDxExenVOz
zuJ4YJXl+JLTJ9mdWOYRrpvDh9LkrL+658jpUsu6cAP/evKpHLp2opIWS/DuOHf7
hwT+ZszoBoDxzF9Z6n8QZ+CT+C3JHUW78LWy2Lway1dR66X0JneillnSs7v0NDwG
RFgqTCXl2+ejNFbVg4/x24SZvon0ZZlFqtoW5FKkwgHLSOGWr1AD/6hg7bhnaZkv
enz4KAWfrfQWocP4Xhn0Q9NQkCVoGDmHnCja4IPdmaQpVoRzQJ5C2iPde0g16gWa
fNO63AklD+Jk7qJuv1esAmR0XzAdGuQA1gd1DXp9UuFkIAD8+kHWILEnljbVpXdL
BKNNdnyAw3f0jW+D/uG71MbOZJEqvhYru6TSL++eSik+x1bu0RRbIPvBb0TYiYpC
ad+qzzwADvjC4aV6wbdri1NfG5kVCOMSRbuzgpgwiOGMyesZlEpKEgvxnE8INC4U
dS7r1s8RMbdFpo0qSxzXg/X8P7pRw6t85yOJych1B7Hn9c3XHuZRzX3OEoX9D1CI
jYnvJp6Arts7cmu/57PMnRmrfLDfGgJkkjYfRxUEVRsogo7qND8gmb4BX9Ea1xRj
Kuv843oSywt4OqNSvt7HwXMTlEBIDxT8S/cpgvos45kzXblUNgAwGdEN12aS/t2p
9Zs4+ihiZQ73+yiqltyThEGBHujY2HqzAZ7Rrptgmsvo1dCfH7TtVqRHeDSpw8ae
SdWeqRLT4s/Ma+zGdoxmgaz6d2D8W+trRDcXApHZnK7V1eUy50GHXVkJPBwS+kC/
tueFaZUNm/KfEh/9lwX7p3qxs4VL3lkBZtADX9H0lZpsyLciKdPtwasBp8ZyEzNx
V/p3L3L2SJQc4xEqlohwQulU1I3j+fHVoZn4lfIqBjb29KAm8D1WTkRhfh5++IdK
0S+/9+3SVHXKAcVzgLjp8ZRa7tPMjhTPhQ+pVl+5cKHKPtkSbCuA5CfwcAjTVvv4
bp7/2TKG/DJg7CIonE/+5hLgRUvHh6xXOMSReY9d4grUG+roP5outu6aUsjyPjvL
PN/bIVbFXhXHXvbHDVSNhNZ/Vuibg8AgYOPXVwJZZRHQ81RYybjcgv1aB7Ca/BeL
QjTiEFmOApoIafgw7i6bHgGUgfaOLcyU+RAB4gTLVqgMCL1HWJQPB6+uSaGZWol7
dFbEWMApkiuIrZiASPPF2xDy/AxVZCx1RO8omu1qWd04TC47N36R9Qi+SLZw9kqf
f4CXubunzkgW14NCy8vzeVfQzp2fuR+DZkRlk4pHrwrbiE+r3lRrN6eIByHepWJ6
5G99bv4dBxO8b+cFlQ4YxtgcdfkshIkg/eynufAkPUlvUArv8ctBP8A2Z2uPjJef
4fWzsMYLDFjwsB9VemnuLb+OdTwvZArelIX7osjhq2gG2rRF7kqFaEKvjoeqke6T
rA2kT+o26Itkb0As9Zl31NQNcF5eSvEZtOBqwJ9vWRixlNzFnNqxJRhON5EuXrRQ
/JuYj/flf4ZXueE9KKfUsR+HoUlF6NnvK05/PN2hKdhuTd2zagK1JMgxPAAAPHvB
1RSdumzeACTbwWrE1kmHJXUuiPu1z1X3onGsb7jtzVyIq39OiQI2ZOlV7Ar6tt0J
5et81R43barbsw9Ag7Q4S0f/h6ID1LtRVNDnt3xUqSRYt/ooT24ujR52tenYLb/D
UeKOcX6m7WhCMHUEnIfpFTVv6YDi69Od6hClb85akpi5j9iifAie5pBkx4GbwtIV
qGMn0MbfGHKq7sqXJaXjp5LDbuKfhMNPm0CYEV6muq0M/S0kFKZVF4H/GDSYBq79
u1NN7vmqx6v9C8P72SxGafqh6np3tsj8G0ua0w88Tfat7p/LHsGk9nich3l3IOss
oeR9u9hBEmiaWzzxtTOpbfGXUsGDZ1S7rnLU+dOUFq7TBje1k5/XJC+J9VttyyNK
F3QlQnHSO9vKil/I2ZJEMWcdD62E6X7z/pwuW84uuxsPHvawtRqyaOMXzd1i5wYL
Xu2FlsgE03AZIRjbbjLGqcEWuvrirKeiHPjdArn0loOeJjXY7nkXyhn98FBOs8Qz
EY2K0+ylKHBVw4IlKwg2JtOejZ55B/FCaU0JxW2ygNPSFBueGSrc4JQhHciSZ/jz
3blBSUpQVt/fTfC/1KmUSDvHaPt+GuqV85rHY89wwWf/v7zDGvvvG+De2n6MqZwM
XdA0t6zFy/qgbC6V35znQ5y4XmhC7z5x4dtHDNN+caFvOweAWgV39rd8ZK0D7d5P
Gtj+zj2ty0uVlWSkfnoUl28hopQjELAjHiQK8mnq0LcAeBeILRlkk1SfiBVdjzRA
XN9u4mUctdy9Q+vjIEFHKifFe25Ah2cbnTm8HJbdVchenLS2zg25jVbmFc01X0ge
jYxm8vDxVfkbs/KmzBLdPTHTYnIaT/cM6C+43PF1IzTEQVHkDsH5D/A/0qNyEG4f
T53yhMepdznN6LYwcWvuha4c4mTJiTGkCtjb824ChDrd2Cl7tdsXWYhU7C2ISAVc
JbypqQo4YTyUeviNxODFMM0CGH/4wqw4ER6xjJzj8Zf5oxvaJ34x5rTEU+EgtLRz
IVImOr2SYPVtjFl0O1rqco8uXzVbctkCAsIEHV+DQ4JvMrY/6ta3TWLVCVr8iw7I
ktRNyYdPc1w0dR4QonFtsA==
`protect END_PROTECTED
