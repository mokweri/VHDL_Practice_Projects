`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8T1yvt8JyotxuGnk83uJoGyHL8GKzOFr9g0wZ3fAY2tiYxmZi54R4ldLDkVmSuAa
31U2uJ5OsUFFZI3lyHXLLTxj4TF8NxCFKxdnAOf3K4701f/qwwJ/+2t/RigmBs1f
dr/T2sEzrkrccmhasqJaNV5t8/9KyqNVWNMl4l6lFx8iwKkmHplSiCacsteZZBDU
eA/lzuG1pGs3nzBjalnp2hx9T33fAy3e+Nb/eF1vORlvmqIE05kPh5D1buH5CMze
xUahCk2j0P6gGmQAirkXB4cE0KCO2BQmaeTeEiSpWQFQiP1X5V9O1t4imAIhVx55
8uNRdtgU0Tw9RTPErlOFF3x+1wkq2m4m0olyyEL0pvWmsQ3ryyszFXwL8Qss6WSL
gHeeNdFJC9JuTsK/JM4PV/Uo7BGcLcW0oLXbvrjliiodVEtbhXmSiLOIGfjw6FK0
I9rqCP2txBQCKTkaWppboQnDwsmfLCiwo19f3vT/6lIox765+7YhVSAyJmNAIGHz
QNKcK+v42+PGewe1cfCSfLTSvqqemId+YQVDsNk2V4ksDrbUYGk3p29tjJELYGjm
HRxt66bALV1XS+glBkt+MdSli+L6Xr8OsT7jLJsyawVQMP3KBUJ1Cfa6guH6LOs5
S3J5Slrdb8H+AZ5rQ6Nyxw5iz7d6GcGxAPB6r0Ddf3+OT9pJK4DbnRiMrRWJPPcF
gxNqO6sjElqDHG2BlaO/HG+QJoeVRSU73PNtgC38liAF7qHKHk3godgoPZxV9b3l
jh4fRSO72LLDGs9E9WpA+Ttyw0h6rJa7urjkEzPek4mMV8jS24sRCNdY5dv1KlID
5o6Rb58XZUhfDG71TxgHU2WUDgI7BPRJSmMbrOS2+PMtEPvKLXXiOPraUwSrVRPb
xK4D4dmmcYWEVjOJefJ+wVvm5naoRyB1GQ2tnSZgK4IvmfdZMrLiVTkO+De8bUSP
DjDoWDINELaga5HZpstDQbbNIBrtsDe2hLX18w61NzayA5Y3NqL2mc4g8K5/oFAg
Y40PLW45uGpyin8l+xWGV9sbJzMW8QX6fUqwUf0HOxzLhUefjNKp7yM6NQcxi7DJ
Y1lpceI2untVH1wz6qhybxZWrw2i7aMj109dVSYDNZyIu8Aw35fbh67bJIa23KVV
e6Pk4o6AA83hEaeq+oXZkeaIySBhJl6BBnPq6+1iFXoFCSBTuN+CF33ZblG/9Sa1
Ha/IxTLqh9T2dJkvnA9dhgg1rupx4sl/cfKigSB3w9qYnQFFXzXOcH/wll9706oR
zzYgFjKcX0/Qm7a2wxYQRg/tOIW2lwnJ1xl5EdTNzVTNHOtZ8Z0fkYbJSB2gKKoG
ilUREWainvg2dsKzae2AAzxbL+8MWokbUi6vcjh7o/WEZRCIY5O2LL2M9o6XpnyC
5c8g2rJ+GIsNTjDAEBC5HNkkwk2U+J1AYFtaQqn1T7DGDTGvTrlhw5psYMzLWRRJ
2FI+TazNr0TcG2DKwiFiVMedVdm503PB40S2vDnMtOR2BveHAGwxgZnnYrm3vn/6
C57BlTMYX/jetmGjmbXOJA==
`protect END_PROTECTED
