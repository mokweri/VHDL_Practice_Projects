`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xMsIDtmd0F/q3TmHfMikhR+6u4LE48geJMVS+LFCu3cyj2QcPisF3iLBjm/+NapF
qOH0h0BSyzdw+23zVIhG5pyWB4JAQXjnTpx/rpSUVr4s1wiVhTLsBhGVXMrLznoK
gUyY2gkm7q8JHbAfE8aLIPCVIvga3UPFs4ntHu5JxTjrs+jKrKI3ZImaCODQqu/4
LnNJ3ARskr5pJAK7Z4Wo+g==
`protect END_PROTECTED
