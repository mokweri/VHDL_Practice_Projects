`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBNMw3wxPzXKffdcV7T2i23GpRKmg4Uh4ooiX2kJE4xy2GIuASYh2a50BU8UUJSt
dLcr0E8rBQIPRfQZoEZ65jU0mV6hKPMQq2+RcH9nibZkTkqQLYW2wTheqWUC2Ojd
j1vBG18ETtwVdZN8CZ/8j8vi4K3JrNOTtQxZq1Za1luP1E1npyz+Vvu4WaYwK+Dm
oIAL8ZACP+mnQeHU27gAuN0lookRwDFHe6+1nHlTdAptxuAdQaw9k+G47cg9lDks
wBIwyr8CVS9aTvgBCcXowUKioxQirorbqueLvj1D0Fg5XjpwCHb0Fo2n92JtBoSB
ichHczi6R/giNxsD4rkWsGrovEOJCccTigUm546QBowVRLQjLODfQLOTmZAmgaB9
MeA9jyFWEr5jWwDBrtrZeWB3uAoXdxoUp/9kjDkQRNnObDWlUnf7t1CKziztQ+ZW
5ZSb3GVbQp0s0JnKos4n7sWdMVbVZxLhg2gvUipa20lrOry4lXyhtADWJ0ivKuRD
g2/Acv8xJQJvOHtNDvF3894LdKmA7qux3hJrA/8FD8WrJQj15GtcbzxuTEQ5HNMb
AxX5nXZLLbugtzQL5HqF9oElyNBknOLF9KEqggDGjCtkC6T58DiF1a+VHPvyafWv
mpZ1maCg3t3myj+jEgWSlBBvoQ8Rd3nFLQkclXdNj9wPNr8PkVz//P8eQj0QxGXp
dhhMgyOx/dXyVHvxFMxSNB6YN1bGfXDkRJqTgHlCAyqQMWbQqfBro62Dq0oulbF2
GxMbWtqFW//fztWUz7H29GrPzBRzmUG6DULtDY9qBBKF0CNL4D1oGKSBaCO6z6IA
OSbzLk3a6ltYc7QuYnYsfY7/yhvL975Gt6FkXD9mClTNJOKbVQ14izeVQKZub44X
UaulNgBUveilhN7YD1jnXWX10VjigV6EDoKUCib/n0uRz4I1Te3Clbk0IEMyBh+Q
aMXydPdo6h7ezdsOznZQAFY63j5HLgkpocW7NHRVZcf7bUqxs0XBUM9RIzYeTlFU
ogQH4aQg73iDmXgyvGpptDhPfF95X2z3s+5NQjffhAAXM7dnZDChJFM7lR1aptu/
CMTIhz1NG5Q4c2yqAk0WX1UGZ2aOqFCWgVaIDkry45D6NNGiUNQ94WJAD5cxjbmy
icXfAm7d6uJndCaLnV0qJtMPrbn9BB+Q15zD+4Acn8hXAYVA9a4/4AAedifcyS04
dPMMljXqy3GypZyTvMQoBbA24vcm4PIuTqEofxoFIfNJ9OCfx6o/kX6+FdwnqZqX
Nl+jsmU3nvy+HlCcwH2WZuVrkv+EWRHIIhLZu+pLF1suA6PtJ8So3F0Wem7O2k2Z
juzDYn09SO3oYB6971OlL21pSyr1zdiVV2ON2bdYlv8xooVJsQur9/ZnEeKPv27r
18valyvJT4h9yLJX1nSIL5j0yOuCaH0eBFNRkn+zTQGVegg+41P+ZlD9JO1B+nD3
temm3q29VbqTNNtYG86TUwduWP3PW02CRPkVwvy4BbohxWqFoXItAMIl9Vd4lY2I
Hwn9hADUAPn/X28mCE+1fli3eMOAk69WAKXiyVDmWLNVSyjm8mdUL3VcFavFHKLU
a6+dtIBk8iOYWVFca63nkLzuFSHgAONvlqb9rMQZYCBBioWEiWYEDOZHVa2KD6/o
nolk2HVjZ+PESeTi7q2xryDW4oZURxrYL+uypOC/k78ppas4s63Iv0nLUg3NmBhH
Ddq8HaTVmBTg+Uey8VtGsh3gIV83AckI3iH0WRBSgm2gud/abXs2fhZ2GRQbXSGD
NbPx+VdugStUwe1t1Sma0FCBbldXWYpBwi1A5LZbefgB0MQ32TApv3JdjrvhZG2p
+o0eD4nJpezR1tVIBm0ar+//wkEadXFeW/gPLCYIcQytRwb85L9QgR5W1AgQ9iDf
xg6qf5qdheb6yOADSgidUwDqVspx2ERY/eXXxADZfwWKNMo1pk3P8KshSOqRnGc1
yEIpxBa7aJcvcSNmhtIGnQ7RlnbAetzGhHvJg5f4DWDPaq+F5rLHNJ71Cc/BNSEq
5h21a9W5BRhBi+u5xdGSZqE7eEFgHc9e3IKzqINxsDV6D824IVBpRDv/k5Lq4N81
jtHKpCPbc9Cg/2/GsI6kwrG6V37w7ws+vzMEjAFDrBs6W6klRhTrS5H3WEQ21kQp
+XsJ0SxfCLYPMIsMCJM+UxCC7xyl1lsi9oFy9roNt8qUUr3+nySypHIJdr+n9kv1
RQujd8tUtc6Y7p3Od2/iBpiO8Ufk1waKPxZOWnCE9lzf8iPMZKxZ6Sw1Py/T1dZ0
gQjktgQvHGaA77zYkCff6aictT7Z6vWlrJJZ7AJ7dBQxLfvoUEUKaXuDsswAA/rL
PKTr4GgD2nlZpgbVseyt7OhErWd7PJCDs1R9EF62YEUOb0JJa+6VGX4SUnY898tD
91wAtSqXHQONrrcYKje3ImPzBqrbm0befcZHtnfuiksuE/I4nHMDM/Mbz79o2uyB
GU67ADqhVONb1PQOKzjH1Cfhc5dD5IT71ECNorp9B6Jm8nt0s1LygGSjt/i1Nxun
irUdwVg+UADGzeElPXYMLeZMiWLMBJ/lm0q/Y5E4VKtOMrv3X2ORPSbVt5/5FWCb
K/lg+U58Ou8INiFmtcHPXYqxNa3BDCBsF/2WxvwDPz2gxy0LpT6CTCT7TeluDnvv
cQ4FueEgFBPnISVVl5zSikNXtV5BBd00b6Tiavwt9Gdq/a0gF98EiuY84345j05p
ZUpSOon4px4RI25BARitIVOrXu5sCJTcpkIgQfS3peTFpCb5Q9RjAiYJo1ZPA/V4
8lg4Ve/uTdkIYGS/QrRLAOLFkUxyzprZSw6Mi8/XA+R9ju/HRtlm+W3mMqxjzP8Z
pvyD/fCFQhXRL6aErGOC4dZ1mxN286MlHPbvsZlpQCyoWkPPwQHYg4GmOJ+EK3w7
osnpZ4+aQ+1SLPod1elG607B6Wy/KVvOVEW56xeoUHGgp4DOgFU+TNL7lC2/a0eC
1mFqcHcbz5F2umm7suh2Y2UskA34wLtUx/JR3B01Ov7ZFkz1oPfligXhh99YZRC9
tcMKisbO9CWk5qnqsooklYWAstWFwl1gagoievYaZWtkuT/ePOUf5ZSpfle7AnCC
Pd3PKxxkiCTReMuvgXnZinGeKkluyrBDQpqQwLUBu1l25lLaetxeHGf6HTSvG2MQ
sMlQi3sd0ufibOYTgIU81IhSOAeNilX1mJMEQoUOlI0ycpdHIO4omAr3Q1J5hGn+
XlSPLieR/qai7vZaj2LJFZ+hi8ZWQg++t1tyRaL5pXJiuwifTp7XrB4tDBezfyWL
Hu3kHDV1K0afTb/ww4f3DeMYXu7SgQAyaEHnLncdHZdNfNkt3SLqORUW7dvVxWZw
cecfNpnZu8zNiHLJICpoZp6WDgxTI9pjxVNGf5yhKlC/noU9enE+8Blhqz8v3Crc
ApOaKQoiom8CSAJfq/xasfkkmI+hNYgOb0FGk+8Wv5c=
`protect END_PROTECTED
