`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGqIs+/cUvHLXMvJHzi6462DIjHfYsKwIahJ9/XBcirq+bm8Ku96qx3HPkA/++3P
7STFI3tTZOA/iS7o+nXshJ+PVp4s0NsfwocyBUSXN0PCMkpOvRWtf9o+d8ZugGTC
e3vgXRmWhbLmWS54p5gIKVRc8vbLrL/uCIOoXOJHk5bMR/qZ2Er12iDmerQDVcoE
HgRAaf5UM15y70mlc2XXX7WO+fxbqzjctKvhURZVuwjQrs7WTaCbOU9WlaGeJ6gd
MdGQ5v9iKGC3XUDuE0r8WHiPfQ1O1BsjDFo1REvQoLDHLNS2z4p+u8r9HeS+xAg0
73R0wNmbAGy/x010Nv0TtJzbbh5RXmpCTOfIbJgdTLTgdSrSLD0FIVzE2qtzs/qO
RWXhj2CFONI39+NPSd2W7uRswn0Bhk2RN0f9yks85SzE7r4ROhsGEolhqsW80vnY
YFz10kfX7z3HHir8LyT3ZSX7El5bTtKNQx4v4E/gUJsUxfHYFtCC550C5966TmMC
7lIEvbR3wgdm0tDunCg9uA==
`protect END_PROTECTED
