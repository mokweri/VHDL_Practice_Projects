`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dIF0QNcDLHdzUcNufPxu0tTDhnI12ia0wSa8lVeJzoc6SS4/vDa+i5355Xm1K9rx
IAlTi+SUUhWKEpRNKNoiZJaX0s11uEO+LFghQQVPeK+w87G44z36IDHsfDNiTATd
eB7EU5zMS9Es2Ac0KHp0xR4liVlJuXPqK4KjthUf0feme4ykkWqKmA+a1haKM2Kw
qNBEIKTgfdfN/4LpknHpBILY+zO8OYGlvn6hh1TyHRTVW0p9UxVmmvsi95BCtlue
UigsMZn9eG8PHXl+BBffCS3q2gXA48+NSlKpB7Akjp+gN0Ip3hOKOGFA5gUg4dil
OQvqC9XwrBNMhiIx+gD+TTXS2W939MiTYbrczM7VgUPn75c1fPDyYrqbJdkf98Op
vYsLw0Z4XieSRn916P4KqoSzZQz9YljhXf9NT2KDdrZgO7jtw5dHgLZubS+gCcCt
GSw8QDf4G9g3Zz4FryCwX08Oj7Tgip0j6dvLTCVsvfxIz5S890cPsa+p7Z0o+oaG
DcgCy8h6CoizfNwfKPpButaYOe0T5bu0VFsxyPXMgmxmS43j/TRxR/I8NTF3zvk8
I+zY2OpzCQj09I96BWOpCIw3ou08mU7tTjSmM8+kpiH36F1MFIXSRe3/Zgn6qLW8
vJ5cb36tjICW1fORTIBlVnXj6qAJh+X4/hgrSZX71ou2xsYC5qUnB3lLFPKdjJ94
UPB4Be4630RJrYUv/PmTKlQO2QQoloG2dIrPYcAJqeuxIiHr5cMIOCmOqfYXgjvX
sq4B+gBYJsaVgBw48ZGM7xt1KEZUmGX8JWeofeJfwAWEWYi3W6t9NKYVQsSzX/LX
JyU5OHY4KEPsDqleQ4p7KtTkxvTNHJLVJDu6iqxC83wPL3pvR5oa4+I3KEVUjm/X
ISMjoNzLlz1IHzHofUBeTtWjfPyCTN7DFduUhBtdOGx9bSQHNdlm7O2npNr60Uvx
M0+UubN9mG45Hn8NiRc10i9yjwSS7iWHBmz568ft2KY=
`protect END_PROTECTED
