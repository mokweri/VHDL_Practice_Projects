`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MxA0MhDN2s3+eNrVxE6r/g0RiJ0Y7mM+WJoQXy/544ivBbmhORML6vatQQFx22JE
e94YNfZgcMMZthRMJiX63CyMODaIKcM4mWR0xQGK2B3IHnUG6XISmZaNUK9nNfos
fg91sAl15TAzstO0Ln3Df1MbYIbXi2PNaaROBtnRPqRd+Gw5+DBd+tpv8q3nMRmT
cbqsV+CHojjhllYiBpUPJSe9U4Tusmko4Qtdv9U2a6Ipsx6zpgOBZeEgI5N5ip8u
1Vjj/DICVSIicuFFDcnaDOt0cDO9VElKNY0qtHz+gwBwcxiAABca9e5Ch2wRSdJS
fqXw4JcILMZ3+7hk4XKrlvTQ2MadXmTczFoivWDqugu9gd727H0s8zk8nzIs4rOh
0lGRWMJ4RSJDktIqggBAivAidMwnBwQBMS0rqAWEC3Rn8Cd+P2jKdcbpKMBmR5sS
kvPFh29fwxOQzRMxjW/rFBiNEZLsbTWF2dooUZKQO61WTSvuuqC8SAV9daPHtiU7
LEBoRG8TUABgv/YmpCKdBaGiCQ3GnLazg3ygwVPkJ1d0BMSZSlP73x22GxRVUST6
`protect END_PROTECTED
