`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AVZmjcvIa5iJ07sYTdYT5gfVLjCCeoA2A2E6NCL7PmJpS3jwv+2Ki94g5DyH623N
gXkQlhymLhyywG371rDLVG6q5GHI1mXdj4JnJzk9wt27/nAJ4B354I7zOBG1fT0P
tps3VPqMnttXJKS1l7MFURmlly5HkXWkeDH8hdnQnVi+1taZV7a03q2+oJ/e1x/v
8qwY5KUznbeLsSvrFNlyzLVCPxprqxoN5O+vLiiI75bfPGBWlZDxo33q7qpxPWm3
0Hmf4tbolJ9S620DLwfeqe1MHDA7yv6hoT4wvYMxMcCekmuNygKpxCQKodq+HA+P
UG0Qq5gisbrQcJWz2NMpM6J65dyjb2ekdX1LaA1gmMysMd84sKadLsHrpR1uu91E
npCKnWwSPDg8qwVMu9loW7HMiDMAdzORx9K/4EWZ08ysd4GjhSY0TjaqXIG2KSsj
3cgTP48qQWHxZ2uz+C6UEvQJrH0H2Go2zPzPlrAevHCVNNtko4lHS8E4i25BYA7m
9puWaqKgrvxKs/j2oQTMPx/1ij/aJlxDNrzjEeTCD1QK6ZmoK+ylmFH7KwcHSxuP
qS534sWFPLcwoOitYdgMZGL6zykZXgtjdTCTkGIhkRSdbAL2X4aBWoH7+OEpYEBr
98zogu/Of+dUvbtAEymMAiFuXjuN60MiiAvPpJ+4Ed7HiX+s3w+vQW4F2DoJhJ+N
thEJfGqq/6dMFLgQguQt3bPlJz3T72udJZnOOm+MsX6+eI34SRZeKcRrQVHnH7iZ
57Z5Bn8veI5XMQ/xu0FnkL9QXS7Cw9yuRYcgt9vkOzU3nmM3vngiQtt7TfjYG+wn
r4/XfZo53SdywrMBsjN8LFrxLuIrtI2egxW1ZwpMdwoCTFUpD3CuyhPJ0PUG/CKW
8zXF1W5tLf9vCtqRhb3Dcpgd+hpBXhFsr1+IVHtKJASROS+G6dX8d+bB4tIOssAT
bZX12E/PPezwycgdmXDKE2GFrZod+3dJQAxk1uPKE56Z6Rv87UfVW9JrA6UB/DkF
a9hAEqrumrmFuEGMXjVLLQ/ChuYLRAeZB1ps7UeO9rbMQJIjq/fxwLuYgiWlv1ov
7DW/JJTqJcDr6oWeGRvon1+4wWlfXT0DSbLE+UHgWMXL0032Z20qob21uorj6pjC
cDTVkXJRc/nRQ/wPmPwRt/Hfb5cDFbTZ+jihbjdzkitM2XVaq0DmrP4sZIbR3qUU
YYPpYHRFefr/QbwPvyJLMtZ+5Vfd8xHcSKDP9IjL/uedoAVG2wsohn5QlCxbfqjr
TRjINOwsGzEf43n8EU+aN6sFrgU1zMg4AYZ4PCOAJAwAAW2zjc3Yoursm9YOdLjn
wMhjjdLhTPr6xQvHpkRrZEJ0vglHsiBa36Gp+17nxVIgIkzfOl3u2AAn+Sz6mZz2
9yKixGt7eQ6Yp/jeoIZw8mqf4W8XiKqPUvIUMA4uO4my1W4/Vh6JJ/SbaQbrUlUO
L3JvniOUq0YTa0xWHEuko8dtfp1YdAnhPPqhZsKY+AGf6pc0Ta29fwqagvphHNHs
l1eXjNgaY87q9vAGgvYIK2CAl5UOFx1jg3KeIUIeIKBmEYCCP1fPPeQhP5IoLRAL
1P4aZeB6SiX1swzDxGW6pNfS7VFx+Lw9mTdFK/Ra/3vLXcoxYZbXFfzdwBdTb8dp
WTzTYJf5Lv4oI5sI+RM/2/oqdQEfDxw9ZELhXjk3rMYlaQcDgA+dhk1sBnNBQPXH
q9c/AL8IBYNWTY5+//tGyQsA4jgJIOjn8tHq4Q+S/2rk5mSd8WAa9Hz3j+mJ3xtE
WjHCuy9sPWoZ4W/tr0EGwZjhv2bHSyAI46jKDx+0slr1TsB9UYNDAM4N+Mvq8L/S
fBRCLez/+yJj3rk/G4JtSHBy1xo/sXVt/L7jYhK5C2dWCtRi4PtBXs41hTE5zsSA
vswP13uAwbphKFehF/subUS4BiwKvIWSU+nH0Kwbxs26i+d74LrtTOgWEgudhOBw
3iIc+ipsVf6hG53NHgKmphRoVo8HmkfdJvXGLrtS7J0QyQXdpbv/VnSDZgHHvOpe
kdlG9avRQZPrQrtIIFkKUUOOqVdDSPjikrVA+t6ZHkrQLz/Nbauh58etU3nBlG6U
BI1a+bp2VuTaZG90uOplKpRlmoBzqsKgnKExtnN7TypsLQyyqScgCY74wQLKwBs1
puQqZchRaN7MJgNw0EXx7qjTrBfFD8UucV2z1MoFWyLzrTkilIwZKIjFbOubvq1d
7tl+cQrguVekycYfKNm3WadhrlMGCnUMj8N1EPJZtPr+lNAKfSmNOpKwaq5587Sz
RslioASKTo1Nr6FokMWmF0ChGgOPfLP0BA+W/6d2lfFRp5qzUskoR128JPnj66+f
pkyjJcnYP61I4QeRG+c7BK/R7g9O9P3L1VALCNNHCy2lkrCfHAF6BBNj8LYQrK76
pc+voQbB9jWlL77nlBdGrbnImAjoMhcKkLiUhfzi9c2n8iZUY27f/NIsKK0sAQXC
spgYkMwGr+TLNgTNgwIb0F5/wL31CK7+QHici/DwpX5uHYV+0Tj4s6Myy5YbtGNS
LBjhtU2sa/hVtkNqZmYB0KuuaUCQbaWiRRhQ8/4p1DYOmittImGHh/glSz4COVkV
W2n9asZ/GNS790StMI2nFr3xKF0F55ccEw7sMfbMygdrvgHFU0BoRxt4jxioMxxD
tkAvqj+gE2uULZAFuuAheu7hC+CuBZgCHw4NrLJb3ZeTuSdHoS2ApjtN0Fod0/cM
BjibLMQpUspJIWFM1udsVHsZheGL4SO4EfFFRloqCm25m/jtvIe45+1qWqRN8E4l
IYUOs6od5iGDgxcq0NqvIKxjT6PJdaslVZHGzaYpGXoyixVicgQqRZb0CRGADUXX
VayPNMFqwYu+V6YxjC2VLTqI8559si45qeowIXMtxZpGBzPh0rSY9/AW9P5K/XmF
yeHs9zQcwsuwNm79Ts2vHiV2oxV6U04Xo13/6Tt5TZ2KxmsNzRYev2E5WoFNfpus
Itk3dz0srOypULZMa0EQAFTP0rAgMH6BOpAiaqYP9GAEsxO3bHwm65bGPJ3nWOIX
0jv7i8Q5zUuYC6hNDrKHCK06sleB5LU3y/UX7TMyE0t+b9D7F7UbzL3S7R20X6VX
tqin0wc/LKiVXdoa2gnUnHgCckBYwQMiA+LBYug1QdkpiECVKukc5QUKzwTBazS0
9MQ2N9hGfqUZLY4l1H3cfYvSkJiAjDI6a0E7rFn2/3N9yCtjjFh4SYy3OWJ14ztn
cbb0SqwqbPOlYoV/N4mzoNJgxccMhoHGhz2U74tCwYntIeURuw0w7Vo/kv51yIMb
g1AYiGldHFWO9s69vurUKD5MJrVzCblIBl2w49VzDrTy5pSEEN2H0+hqe2ePVh4s
KrR/h5D30HuRc/l3sKszAHUpcLIL00bpKfn/dZBbYqlZqWr4SpElnhxYEY8X/siJ
vexryTCIsmFOIufckyfIir34od1wFQCi053lfTAdTwGwNl1ra6A/q/syI46oO6Db
d4Zvt5a6pXHOiSuodoc3weWHtg6VB5hx4btJM7LZy96VHMN8MqreQoWn7esfFVsZ
d6d5iA/zeSKA6xLE9rKbkFxQ8kShY5cVm9959P8f91ynmiwOIBk6fV+Idoy6FAZX
O2IKyEvsKmm8sdAZHLSGpkf1jkz3lzaEM9k1PAdGsUoZqH291prVTFu6eSvnT0q5
w+6nWy0TlWzTC/LdVU3jzRtE2eXGpqkLCM6fUAQwmXusJr31fUu0oISLrC9jlNkR
H5Idx5Kh7nOPBvebNw0/jv9dbxdDH9u696wmuboPXkWAcZVA8xkH8kkpUgHoPO+a
QBlFR6E6Vt3HosjBpAcqCyjx8Db1MWSgdJuO548BVUWX9j/GIni4mjvLBemHQc4j
eDpCVz74BVC2J8zMq3dgn6WkJEfjY4+LkH+bMLzEXHzAkHX6vxF+022/XnVECgd3
6CGTu7T1EUCV51oeNb9umofhpeNCU3zgD+iY+vNH6zaMe0Ao/3pKZhgMz+03gVXY
DqBzobQPbwpVfg1TtH3vzjlgmX/yYtn7K/5wBdHbVvokBHdtydhCq6/l3ZjBXOrk
+f20nq7oQ24c/assokTrHhWLsf3Y5jFTAWsp4ZtbOhQSdrx5a193FheRDFBMrHFn
khSP5D68iVa6CRmsZoJF5Bnir+RuqoOGFTxLkTEvKCx02CvTViVXp0cCIl2Z2eG5
NhAvIwfXMVNHHCjiV4trnJ5hEoibVaRA4wSWs1P0XEy8hlZizHZRrN/lffQVbnnV
ph+PYfTVwhrP+uGtSRxAyn1yDwXmRFg7bMh+Y5LQUhHaItO5Ut9jIhwSlGe8WLeF
O9FszCvRD24X6FcH3o5DH/vYJsztNxUu/94VnsVPOxjFEgYU+lOiNNnThjh0x6IJ
iTPW7hYlqW8VCzlQqQ0CzMFyVAhrboH0Yhe7ski7Ha4nl1WknQD/mhyzRdgpBEe7
S12JSVGxz555pWAoVd+ri9FIKydnIvp0NPNniCj60YrDTxKm1Fb8LDydMtiMp5hI
HxEtheZnifO0xOd3c044pGeL0HWE84VcxTUtE1fD115YUpC277EjchEbe8+xulOq
6icIJGe4O+zVQeeBvGz8U0E6DrUivUMgfRJmbdbuOiyiMAUzwmnIDc85BOYfhF/w
ruD8GAnKq0uoG3UZwZG7wLf+57mzlV1t7igTS767PZ7Mb76DtlcbRU7fUKktyZ9X
0XR91ZTmH94RIZBIe3RAqf4lU+givbtUDoXaN28ZCndmDtV+Cl/Zy8sLBFBFYcSP
5tmE886/Kf+XNIj1lk7hdMU4FTI7LY6LikRzfJeCX+YiYHboMfBSBBBRBcB3gwVy
J03r/x21FswcJ09F7g+SzfEzYp5FujuzOq0whnto9zSPQvK0r6tkBQC5nPPtKj9B
PLGT6N2anYWLXN0abvFpAVFdGPJZXeU4dNOc4jzy7cjhSW2OQOb6kTn2GnxX7yEZ
UFnfFf/jDOr+AxFJ+rrOh13A/kAUkuR+A4xXVizrr1qSjmXzr19PNFeX9ecLB5eR
tC1zH9tdmeT5uPqoDYjaNVDH7pqRsVtEleeLdCO4CxbJ5arPBdUnbnd99EhAPXZJ
GfvbekZg47Hv/MU1VffPT1z1ituIV9v79V87cdFzb8FawlWT303DrwNHMxRqv48f
xmLge7+Qaws3yuEaVnByx8dt79mnDNwsOg7luhbmDcWjeYmghmQ8ZG19J7ZJ55F6
uGdT6+WJmtnqkx+Z6hSF42LtiB5zim/OoRj5AiefvucqR9AVgODcv7PiWpbW9fK9
7apugNA6EpbMZ/PyVZd9YqRLAhr8nrepXk4mUQwmRB9FRozwZV2Zl7bepH+xDHow
7E5jilRgtgNmG1Xtps/p0OSl8Y3DUKAgyPi5Rz5ta2ts9p5xgo2CqqXtqAcN35uJ
RtpE3++yHAx9IFiaXc89QwGPN9egiA2oao5t6Q4UpsHGozWMt5KjumO77UQDYKqY
WRWdEENZ7wpnw3Uuqvy3fRg7t+hZ/i+PfhUDeJbKa0Yk0KeJZZh9I7Ff528MqDR6
GBctPXgzFn4PyaFDDQFj89bo1bL60wGLdafOF9Hy1F2L5U0cD9hS0m3+JDCBbAzP
OscUStIcO0YOhhtfGgiXw5gezMQIVTVTJBI1SkRbIvaPQoZnf7yPYZpQCgGjT6VX
FVb/RBw25meOTw0KZnkSFohKJynnEMd9xeTLdAQBJap18ITcb9VHbQxATReQoiSC
f4fsBhltp2l0GUaMRUKxDAOpFqRgKXoU8n89xt/Lsv7SSoEYZumAzZgT/DVLnC35
Uv6EVf63gFvjMUOMRBSGvC3lqVd7+artyaS8Ow2EIMjyLvkEE2fgUtQETcNNIJze
Yoce8wORBCxXcXR+9p9+87hMwyPir2OqOgN92SiWm+XY6u4qLVrgRhOhjEYgBH9N
ThtrpDZK545EQwO7OIVXohMYAashx9ye3eTsYkYE6T3q594eE5XYq3Pmpv7F7/KP
muO7ofsHhgawC+fl/M4bK0DX8Je9XSEtBdUiVRg/BVNv8a+Uxar2cFaN0VLkg8Ex
+znj6gMzOk97nZCRvzPMJW8i7Zo/tZ3IfzBnp8SNg+bBN5ov+UPgRQSlPSPr1BDw
grK1e60bmchsEQCZm4KHppGUtpMkY4Xu3Bv3aoapzjU8Nrt0JG2ZYr4xx30ze/5h
COITCtaB1neLMIhnlV50zMqrlcvU9dtaSO69chUWXdwugdnnGM8d6boGySA1xS7f
RwwsVP/yk56TbH7Ek1KqPJuhLM/KI8q9lxVZIhZT7BucOu0OLJ3N6v9kShJxkmEh
/PGCDhn766h7KjoteIQdd8HbUDYArvRjI+8nVziWJro1LPuZhk5H1BG3rmDJVFZ6
+Q4bGnhu6A/tdQnGvvvt70yWoWyDVIWlImmgoh92Nk3+xFnDbY0JYZF1qDsKQoaB
raamLN+rApFoFmHiSoTIh3Bs5N2c4KWEt078tv9eAN9r7zyyrnYEWccfnh1098lX
b/gphMZfpq1QHh6/TIRY8Q8PfayQvI0G9UNf2wTannrlvPaizI4gL3FRhh7y3TrD
+/9Ydfi8kNrGf3L6kNWAX2B9+fRw35ceDdSUDwHuqxUNoJtaSnoadpQ52O7xe1KI
iJ9IrLc914fI3xraOaF3KajOWoLQRzlCQbrk1mR8xebi6FVe4QVNq1muPuWJdlOA
g3mWLxOXIbyQYSqLToFqLWVreG8pdjQE7j7usrnzu8BHpgUOJhDxELTYUXqXVwMR
4w0/Z82DjjRf/HE51+KdgCPJkgaWZx3pxE2sgyj1tx0fH2euyu4cI7kKDZsDGu0X
u6jOQi2TlRxf8+lIsj0Vv0GnVgrT1/q6+O6cS43KAF1TvFhi35xLBbDC1dlA92U6
3yGnWb/PJ7fBPiuAyC4EL1rcefKv19l7ktLWk3cvQjlLpcx+Tl5LUHyP0Oc+V05n
qE7nonjLzh4Au8e7zYhzBZga7uJdwORwKuDFbHuaxcfAq/yq8urPP3oHQrL9QvKh
GBevQqaEUYHTIFs14lEHfWv7PvqUKECI8OFbIvVj0xx8xpCDFMMqk2f2gVvJA9rl
k0GmKbGJYEpAz8a4YiOd1Zwa0tVnVu8Rf2ZPg2WKnv1BJ4h6WGsLGHR5qxj5qDwe
dn4NMSOKHVzHJl3+t1UmiwqR+/5dzj+UJ8UT5y8Fq11K2GgtGZtEAdta81SgDhWu
4kplakfsUqxbKtuqyxGmPNbtzASFbZQh065tkdzxmm+OYCLvgIf5ZeB1xOy5VKwX
Qv2oZ73qvZKqTsWP6xgsi00S3Ph2ogYQ4JsejNyjrkhbo+Fq6PhUXGeB1mzLRJBj
vckS8qxd3V5v3Io/xPX3m2JUG81ZIqunFwAVlz+lQ7kVc0eSmExl7Al0ImuOZAUF
2DhnDCgi5SugpWR2eq6l3X6r9dlzcckaurXN4A376NKD7WPxAEWfRfmOEL7AuPQD
AKmvsnpEVQZQqwBsSSXp+/NUWZzmOYqHNkzpfIvc41I73cYP+NUNUnb0XY00ApUB
jkQqQYe7EccvCxHAzNqrGF37/oNnRbHouf4ICweVcf45cQsE/nuRSgSEZfQv/iRP
aTG8Z+KMFHavh6NxqncWl0L+6YQg/zSMXroEUPdMydOhRqqNYVBK+LbS/lLRU5s+
b4reEdH9KAW/bHVXthU6Ezx0tjftDn5is7gcdMn2ThQTlllcg/qt58ynfxmp+wFY
jJFchJ7S9fk3FyCMBzs4wNSNjQ1mNi/VpXwtltv+b4d7un9kOlsoVxRAOIDyXjWg
uB6ivUlbk6xVITkVJcwdzv/Fi+FZRQutYyViS877oBcFVwmjpQESA/6GK4s0s9YE
W9d2uVFY/Q6Olc6rhvBeQznCgisutIwP3PkGCnlQgBhUDKNp9fya6+3DPBgh5/5o
EeET6lqBoyYvv49qOkpShMUH+K+IJwV0dCDJj56AIp7BL01WJECCnh+SD5DDeRLv
EUf2mq4oGi4yGdLPoDzmZ1+XlhF4wtVLgKHOOVXaRz/nJEt4zHE0+WpJjaGPBCfo
B5L3Rev2uQfACKcHgQ3YVp7jj79IQuzTDTXv03nD+QDh/UXlBVQ3dWRKzEj+oMdq
wTS1/SQNSm82nmF9ssm+Y2VV8DWMNsx/mb5aUX7b9BdechdcoOY+oKsdfO5y+a6D
y7iIHPDeU1d5K0fEu9ZFzKm4CsZfmqV8Q90l8GO/ZyZDrrSIU0iueu5Go3w2IEMz
L6v1B4pQyAIToJpV5cH3gZb/UdOuywDyAfi+IakABdSfZt7hbutXU/d6TzzZ5FNM
F8xQkR5fppre+8xgDHD/+gH5CqDWNG2CzDdke8kVl9/v2RNd3E+jsMitoh920FIO
FQJhMynjd39vhIF4wviOEZIH5S9uKHuOJVvx9Zx36R0CD+8Gv5PER05BXc2Hgmox
sxPyfzoBXTNEdN/TMA1Lp2Xv1QSeyxZyXsewVfJxj6fXVqeQA3smcjrMq8otX26u
/ixhxHhqqBr4rzTjrToLyTZ3O5emq0iONFyybtj9A2FrSeLUbNH/XJXM8h78Yd0s
HU7jSEhT1tupLU+AvezqB0Uy7bA7Lbr089JjydnFon0ITkfnnz7IOW8iRm7R/UM2
xJVTSSQmaCkPiX/XBvA1TjXoQM5UQpgC4JpjR8aoOdS3D1/5CBz/m00iyY1nIQCo
lNAMaVR6O2HyhMOth8UfJHqMLjParrAhvoY6Sik9Ppp8SQRANutLdF0AMt8msApC
EX6L+lNL9oMXy0fc3xtnTSrJHq/J9E1s4ZddM1HGJjBns3SZHNeGH5ruG3mW9Q9w
mMC3k+MrUalswwR4n70D1dESBLiG3sF2fJTfxkArAXo94Ojrf+8wKH7o86gAGBoJ
aBwLFacq44XMSLUQr9wUsUwfyXysSBM+Gms8qdlM4bVwaJjYcYLXDPUDRZwspnUq
jGgsMAU2LC6W0Z2abFcnKt8YKnST2dCOSRK1Ou9ASp32cTFz5PbBdw+HJApxGztW
3JS8BZtCz65usU6RCPEdxC+O3QSW8gScsbzT9v5hDhSr6Z2Op25OsGdLD+0oApTt
yKrhsZ0WsebhqeIdbmBJEO8b460tMJyJWw1QdsHpPy50lNVWNuWVUP/+O2KNTwcT
tA+FqjIKO1f7DF42OTr5rvZ6LuYa2xH/gtu7534oio+Hj8ZHowB8LPifUmHdCMc6
leaIPhVcOM8UAi4evK8HEdzpJ4fM+eT4NZIHsPum7H7hsEMgNCSp8XF6qJ8z/nBQ
4FpIJ2KtQdM8b15mp9s5N2ZP8RmArqTwj0u0eui1m3HKYLwkTAw0Whd7CDbIXqLi
zs5JPADWqDYRf/5cFJc5pkpIDs1Bd2AZoNb0Ly7hL4ZuaogAkkGX3H+Z7RFFolyi
xvdALkGgqVSP1eiHhxVf0w/4Phi+TVHDkyRmUEG30rEQljc3hlgtUKfmPfuqAdEW
2DrPx7fNkFawtQGhIznbOd5mZV4PS2Wsg9syx6R/lyBAv5VoX7sJL2vPnUp2av9h
JbICzEQxV461fPbMGf/btPTuI9AOoRNk6MQGaIE+xZpCfd4gMWZCM9qKviPtkp8h
l7UUhiDOoPP9c8zbdTJ4ngeFpJPBRg88De2velM7/mgvGUWitnc74+uklrsAP8z7
JKq9IG2vVHzyS1DgWsTwkGDulR93xOteEt/nRfZ9z5InJnIWbSzjElkeJhdQOMtF
jGB1FpzxBXGcefEh9zS5dB37jmuvMK8eTsYzuHHLjjMnj2Q6IQQj1x+juHTB+zwS
/txybAv+Yx865wHX73e/8b1MJxdRhHFAjz7MI1r1Gfisuv7fGjTlRFNi22WlZ2D/
KUTXKah3gCTE36vt+FaiokW6zXgOfQZ9vqu7M44scH5odK8Ddy2c4yAM9Wg56GiW
3gzS4udf2sghMfyZP/FCPillpFGoPmuQ2Y1Wo54U9xaQ+I4PeK2iopU/splfYFdz
4tByeijQcaV0PrVfofh8xpt0B/R+N+c2M7wBYpeGahUJF99nBpLOgk5q9XGHBsQt
vzJqTtGWFFcLxCINMJ00dtfaGiRGrckw8XFfYAvOR6j/M4JvbPg4GBLGuNJ4zydh
1CC51n1tatAbvbjeWhaMA6rPwD0e647yK2zfMzWg+Uu6KCLvfyz0FbmSvQiEKTiu
Dsage23N8RTtEV/EqY7jag4sgc+AHQutU7YX/sP4Mf8ENAVTkXNgRA9dlCgspYlq
tW7QzyCA1KmGjRIPni/Z80/GyU06U9Q9g2/FEMopMMuKSef7UrrePmHZDXiLoJyE
AlykYpSMqhBT8jODj6YkA0KcNlBe5wwnwzczxCOVxLbzrm3TksAjPQeOgGRn36ml
WYVYenxYydYi4tUEs4I/WvRjd/8TgqCV1vhxaISuzdl9Yf3XB2EBwZXHI07Br9GO
Jf7pQLGTmto9YOTkAFglyaoaK+IBNGL63ijESeCqGGK2vB5M1eKHPnd0A0FGeJSX
nPek1hbXkjWKNxcWbYw7vZSzsUvt1mjoy64P4KUFAzb1u9eqPMm9RnIzDtO62uvZ
Im0aNK3zgOJq3+7BYLr47QOICECnu+gWQaU64M8Nd27MRRofvCMDPIMREXZFSJok
Ro/UzS16tBRnUPx92tkQryF3c4o0mWCvYeROEcX4kLU2ALywc9snL80QV0ADw4O/
X7jhYef1o/XWh0p+JMqehuzfB1Al/6bDrqwXXvvvQpGZOSCYHfmYk5tnUDTQkMnS
hghuKfklH1bTgSfs/LqtVuWCermaiw++Cnd4bNhVL+QIU1SWZUPJ9QE4gR4AeVIx
zPRjIxdHl83PZlZLJ4FLBFJXdgHXHTfJIHd/bFukMH9Upw6P56ghCgeKkoN2bF9/
+qpbuZN6i9iZ/ECFco277tiI4KAK8iFsMU0fr8ZyziQaSun3ZX97mOnrUBFIHZwS
Xxx9x/iuObf6sph41givvGukgiW5raBFgQulbCTjdnBRaNsdRbDreuA8m7ZtIyYe
185117L1Pc6vr7T8mz1homrdJxp6yEk+SX/4XHnJYWbDyHOlEUk8wp8rEYDHwjfV
BDhKVGkiMmxEmP7jf2CHDmL0GQSbRFcuqzZhbfwCWimzdQwb9UD22R1mmJNqkX7D
1Gk6P4JH2AsaUN+enq6u5wzAcuQ+fkgy/W1qc3p9NA39uSSn3NgconSXm7bxfFMH
47dpLjrAg4kGx0eNuYbd9EbLLzBoArNaOUjDCsDwk822YFNxVBslIfCKF/KqrXXT
b3Rl+tJRjOjDYlMcTfhD0yMQ63YzFCla/UzKFG1HkCmgPMa7RFd634NUQFnK5zCw
pxgtkdraxMNFR/2KBWFA7+1LJnDMg/BiFmXNwfD56IAlAjsYAmHpLtvgqdG2c9DI
ESb25S1OGSg0mItT7fR83RLXVmQ34Ajl4DVmXG3zyztfWyeqgIclDGkczg2Ae+b7
TiXVnrxRdioxfLC9gZddSybKcCQK419ZdGADRg2YUzZVL4I3ANUZ9u8xiY3YTFmN
ZnijeGOawekB7x1YfdaUSfMhR0hQjI2Frtr5BapUr3FtL2LXgunh/APWwL5XanSM
RPrs6e0VA9GpjAsVvqp6rNtyEvpNOJG1/0OBq20hnEew+mWi9mz0yQ8IeoASoExH
kZPDpDyCG1I91CTPnvKp5fnnzF2034pXB1qBignrKYgx2hXmwCFbvdn9EL0m9Okz
tUYEHdAD9sd6rGamdOVClZYvmiil9w1d77x5/UPTQTbaNAzQCA2KEpfHCIzE0pKV
2K1oONPqH0T+WWt07Xarks3jfC698cPWrX3xPjj6RmSPSRt8gT99QV7PZU4xYwmj
SFJQvPFte7+qwI4HRwGHFdzIkPZHUFy9UCfFhWGaX1BoVKmtuUKeJ8Gebj4DOfKs
Wil4g9R4WjiEaRsWGMLISf2EOfPWIngp2gzExNG9Y6eQOGiUoDJDTRuaxqZSbFSp
G5kw9GHEwrt63Vzx1AJE3jpFuOtcIDYGXh0pgMVwmHPUTy7bEwqjrsarNBC+QQlA
725cPJPyLBHXkENiYt3EhBl45ywZVPQWmWTHvxciFFt9JrqAr3lgszROqI3eXhdF
hF8reY6ai66a+JDXLnRXoZfx7HpASWhTl8Eag5Vcy6iOF6EdHoCKjZTHjblKpAY9
ZMtnELzdi32uctbD01SBlH6GcZ2CHlBuTpHHaXunPihX/qlfTh5BHOBAdqu44/lN
1Au5HYiYeUEsalHKWM84P4jWKyKeiSmNQtrSHe1cPCBHVJdNxDWD4p7wI3I2eOxY
RspOImcd0v1ANHwEmJTU9NRkNOdUxtvcbHvL5OWSLtLk8ULzt5M6yR2nZCwK8zSD
BQZj4F+NvS5NnPDkvfmKU4x2PxSXcMYypArulk2rkChPD+jT6Tt6KY0SM1JLJXii
wKxiKtZlFB0HTYIx0doD/sWRnyOroo+gsRQb7O1B9l9QkQXAJTyu5xozHlvb246+
DlzUeyE9PVaOpH99SIhGmg==
`protect END_PROTECTED
