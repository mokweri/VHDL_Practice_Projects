`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPepK3iUv97KQ5nxVDYh6wygYO4TN2I+2rWX4Ekpdntg8QJ2+zePrrvZg5lwo6yy
78hcc7fLAqEat07GYLpB6xt7P6ZUYck7uh7xJpAWgUpkcndl8He3XnSSerfdwLU6
lv7fsn4XluLFUawNu59oWz7n/HExX22WOtG9TYCwEFV8Z4j/uqzELOa6DXlKo8Wz
+2WF5FdSQUf0un/eID+O/TQ4Mgz7bVVozuMaF+PaKDHyzUKHs9ICvRjhGK4bL5Kk
HbHbPlJ+wlGdFxfYFV5pC78FVdzHuuEmqGwn/Juflgi5OKHki+bMsAY4h5qYTMsv
Id8VdwK+E1zAJdWzdO/5NmtUjkzXrRVJEAjASENIPCm+s2fJEGUwcfIV06GodGLC
oa4oKxWOZf4ykmeOawOJHvYUEfUelVZ6ajyWBRAGewD3DmHXbhQtRBb9aVF8np1V
S0IVDR3HVyykTvq6+53c2HKH1ZVUvx0yn1hOrvAAqpkZljFYYdJh8xeDAYsVSpYn
3coWt1IF0Qp/R0nFmGdCMHtf24G8WVzN4DkdRWdcfu7/RjOIKq//ezrJnQQYKbBc
sm3TkoYrzYkV00Abs/64MstC8+ash/77uhrEq4ve7ik5bu7ICRzMgk6z1LN8EnU6
y80/V9wq3x+hPIZFXiUKoc6h5TuVccnZgJNTUtGtaagTK5XtY4pk/yTieeMcNfd0
x9VM1UrwlrD0J13G01YnxDIXzcddwG/XWuizITl+IQHptbX5ZVIjc3Dcc6wjcL5z
TeLWHAsHwZQ5OOik1rJ9pp2eOJE+PTpB5NF+Csz3jkhjVP0hMCSUzTH91aGGzhGv
/iNiOI/cYYMDq2n6IyWpvXzZrjvrtxpSTrTx4hmQAWfAN51iIrvqcE6NZoOzze9a
Sjf6OfbDwv5aLAs1i7wnj5XAA2QTMCMBFMbO/1cSvZdUHi2Rz0zdFmIfEX3s7k+Q
z52BYezkkO1eWHDKyvr4dhcs2nBGptqRQQ+yYbK/kB2mj1Icw6ugl/DcmR9IoOw3
0jkwbKQnU1NI7tab4baOEPwcQCEKXv3hdbWgA41HIPQe3um9U8gUHHy+1BzRHKHe
t+JqHu1o6SiAZoZumzsUm07thTKHjD2v0C9Vx1N+Qbq3y1FY5nTZt5eA4KQhu8m8
RudHB0Yzt7EgvicKaXpCQkaM9mUvb1QVL95GH2PvjgoVXQT9ng9ZMEMFRb/p0l/s
EEbEX6aswJQloCCq6F4I4YU9AHrW+bR1pcFb+fpO4pR+ORO2+mRplOrDXtClQ7oj
lTKZ6yX+BHJVbI1HitiNJvp9ABeOkRv6AWky6GVUe0Y1TzyhlBS/m7sbvpAvClpt
Hh91cohYszKsVjuagzYM4McL7RonUBQCQVhGiCi+nW3eyBA+8lltT3EYt4CHLpMQ
`protect END_PROTECTED
