`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lA5K87YxF/3F7R/zbDt6rjUC3o5t/QU33/GiLJmHX7wI2rQVVr5bjn6mWtbaGW8X
tIsoHeKPicKz/hbj3m7HRSSW6hiEN/GKlYmXfZu9XFfZ2xCVogfSo1p1L33KTxG3
0miDc7QkpVi6dWQEohEJiixXabjfrmgIXU/SgKJBekKJorYupGdTL77w6EVGta7m
7VoOrK3K/JGlK9dPlNB0lw1LhfFpCt9PDVRxflzU676bPz75DFRCOYv41HgM7LsY
i3YQSs2a7iioT1B43zNQDqPjBa67dOlB04346xYcRkZMCptJMmG5iyyLP9fkn1+f
Xnxvyd0EH74Z7bwn0jfMmhXQ8xqZXZf3yhAsFhA1LyHAkOG3GYBLR+EVYUQ5cYzz
AIdlxNZO4wYYlipbhV5LWNmssTBFHDp+r+tDgYYJ64okFw5bK+En6yP5EVvn3wdX
ZqfbQH7JdRDhkRLsCMgdoUmi3J5ZKVw15gcHz7UTzyL7iP0ThnfJ58hge9+V2N8N
JW0E7o0xmIyvNBQYnE4lGbggeDLGE5Ig/inxGvBvEzZwHV6akvstVIH+/d0Qoc7W
Cs5Mj5KdAq+7ejJc+VIG7mJhyiInKtVVi0o6gbtVxUqB4DpFvgOxMVxJLl2NUhB0
pBe1oul2vWCKyQX3vLlrBAz5Cw3FoTl/d3QP3VSffnmjsyT9PM1yqN3dXe+cVNYF
SpZcFWTKHA9J/YDzli5uz2z/A3lTQnQ7gHttrhOf6xtQHfqg2nIudZCkNOAH+VbV
2g6HxtO3t92mkZorOSg/iz/IsBTi6Qt84A7eNZWYQ6GS224S+oA8KT5GfFEESckZ
r0qQDmOVinTpoPiFlphGllww6fPvYVcdQbDVP9kz+dYNhl97S7JysJ2lqc/UH4uc
gYeybRTitOmIwQ3+1JyhMbpC4C/p3C67GGMjwlmlNSzXOT0xydOcWQ2E4HOs/+xW
fqUOv6dqEJhUU8aPkq3EaicgLjXw2nQ6VBfCBzMKgnpUJ+VZ8Xg2H+LPTSac48JI
PHDEUubrlF2zcqv67G9jmGdaYanqJBK5G2x3hBNhPT/SHMyA37ogVTcx/pB05wn7
nepKYi5/7TyHRsJdndIg39jBCwjNATUSEFrJD3pJ6QEIbk9ddkiZ7zqIvmrl/R4g
7CfaxRoEzYuAcWdNDvlOscOUOtYM4oqQ4L6MxsBthEfzFiCk5/r4Cr8lRzXnlvrI
yk8ovSh6Mel49zOZvvL1k4mC8KZ9xcRQYFk6wuKIBAFMCvYkssSFm+VmXohFr/sY
hIbOcZsJ64UvHF7kJ1345kwB2xrb5WG3pADqLIiZkD3a1ukWNCjcOKhDQrbINnaw
W/AA848Z8YB7gZY8qa+j/j/o1k026KLCLMnUXrGf2edXcGKXk9awaB7/AwZUUb2b
KM7Qbnmaw/mi8QVuqWIBaiAjUn5MNbiVld8RbuSFIY40RdgvCgnjubEoMYa7IlDh
AMrzsQ4B0fYXvSLyxHQJOD+vKyR/HZin2N4ZURTUcXpZjKCXDcNV6RsKx9cusWYt
3/f3fJnRhwYEhh5Cxq+XmrGNHdD6H1qRViSUIddGjDH4qmP3re0wIa/KhCMQVD3Q
tEK3Ie7yvTF9LikFkQTBO5OwPlRkqsemPCgbIQmYojhJYRebcep6OBQWuWnd8uxG
eF/pzbctRdt8N7P5grVfQDnzTYEvzyaajwEoGLL6dSERKclCOVrU3J4a26rBe/SW
EUjRV58ckKbqJcHhaa7JHSuUpPgWm0v6Z/xpO8ZQoRv/aFCYb1oO/now7zP5kmRR
Ujw8eLN27wed/mcbR6+xQ67QH/hUpUe94TKsu0Dp0mtguD0dSPf97h34IuFGOW0R
vFkgaaO3q+yZeWsfl4h1kQy7ocl8HbuzIdiBaoRpSstwKr969uXp8TppEofxJaMY
ep0uzfWXiF6729vOZ7R+zA==
`protect END_PROTECTED
