`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/bVgG4DmCcmAnZU78rJoGRFtqvrBbdLZTroXwvISi7G55rdyLy5KwvWuMPvmXK9
JryRzU3MuymKtwDtXqT/0FUXgpDEvdcEzbC9CZBgbiiU/6PHYX9makHyUV83o3Ds
S5Yt3asUZAJ+MrQrGQqhQwSc52zi4duP8HwdVuBGIw8bXtC2KZJvD/qqYOnTVMD1
WNgzi8ZR3ybMoB/CP6YkmRtZaneCknygWsdv2FgOB9dmEoi3Q1vSESEKM8J2z2Af
eq2qgvCoplguWpGVGcDbrw7Wm71X/Zvwa9/WWnmC/BAYF09pGcGQDZekYY5Cm2JI
FgBi7qQjvAunWqClOi7yn/Gs7r3EDt80xrZ3JDamdehLbdJrxuz3kvKcJBMR5d6t
aTCDj7WNJUID1uEiBWlGE4Z4wTz+8wPF0Rq1We489b+gXkx2axNAxHKRuUlGQpk6
OD72fVDPzhjGojnkxXzlueXB769fLbc0F/YijjYwTcp98NCL/DeUvcVHziIBt+QS
g7Gr1cs1U+oybA77pGG4cUGBhSNOtsYLgb1PXKCRJ0m2yFtIrmaavtyv7vM/Nhtb
l7IBarIwfyHqpYbFT99KoKuRw2qhJyA2izbq5MMtYLqs8yJLrRCBq5Id6gViZ13b
mdRLdItLHETfn8XF/l05ssE2DdYwQkMo0fU86CiCjFok5Gox4IUzO2fQfFAB0vmE
ABprbRbGKxyvu9sYhEzGZHC+l+51Yy9IXIlSNVa3Ng4UQ+d503GzAzoeQIkndH7U
aiIaP+yrZ/Np45XsxG5TPsuvdFtGn9LzyJISX3ogX9iBC5livkijtnd6hhda/SNW
6jRZtK54rbn/uykNqidftjNyLpgjKwlCsow+KYTbZVABI0/eA6OgImBUUamEldly
ML27CyzzlgKVwbWMlT+KZg4CEeALqIglPOagi16Oinf8pdgPkoWqG/L8TYlfT6YY
2bgrt2mkCk4RbiaJ7Xi47nj+CM6CiAPUPw5Wbr/tI2k7myMJt9J5X3K2YRr+odVO
036DIsKYyv4wAWfPSuVEbzwL3g7tbi1fTA9mbkwSQcjwqiXAum+IMYhGeH6z5mgX
/RxGgWefAKowWF040qg2E0XfVrO7Bq3/iyIaCr0wTj3YZNbdwr9BYfk7MNJu33AM
D2Cdjm+lRjFsbXNMX9YBiRtlXHO4cAChRnCYQXnbKS2DDZ0v1+ZHbxWIyReSfjJI
Cu0CnbQhck0NYzBHdGsUbSbXLJ48jHdw0fAG90BR9TGbgs4BgTLuWHXZNeUKlmDs
DFJtp1qtTgoj98gjrKfVP2uvAe+SG7BqPsHp1nmFMoC8B7k6uYkSG+k0CjHaP+1k
dzOuSTf2zrWHB8iT1CbY/EQhhnuMe4C9tm7W6JbVE3ynYvnVDXdW65jQf2tvKnqK
TowVABUfKLohi8m18N9TAnkRU76IpEqqB+bKbNzX+mHdFOLACAicJITsegTlBOgJ
U2KBHNNMBljFnsWup3ydBxM9AkElzXQzKFAZipHuUiNMatCmG54hIAn3UUS5Ltpa
FH4vr6c44/un/nJF0wxfITWieOKtCZ3R1SYNI4c+PSrLMEVVtQ0DNzI1IUZfg8rT
FCtyQCydSAhj9vJf8n2h35K8CAFq5nO1W/YZt4sxySAUm2BxuWadkYW0dGJX2Pf5
zyfjXXMkZZtmeZM2jqsA0x+cKQDMNBE06aOicpr8FmsAbZDodaNCNzZk+EDbbTu2
XfVRG7ITgX5VN4nZQ2LwMhjqmZgQAqU5UqObGQxC0sFDEYwQChRoCzrlh5Og4KB+
IaVGgjUXqiY7d9kidwpbXKn62gsFnF/u2VOjHCUosQ1OtlAe8uy2O1pgqzgrUXtu
X9QFtewpjrjd+w1Cwys+/JL7QAV3efjbqfsBcExzXEXU3y1otdqmohQkzWBhKZhe
jLNEWhnn5/BxiC/n9c2oSqlxNtLENopLQ6nMsvp3WPAJ/rDKbLAKF7aOZZeukkzo
VDV8EQ1a4ndV/hBgGBu6U/UdzFJ0rlPG6y+TWr4QXpDChGbKMF6iN1vAbgH4xsXj
w9gbXPMyYaD4/zu0I9J3wpwxlqgVDr+kxE1Td1kL5tUXKXHMF30h5Ud/AK39JnGi
WmtfkeVEnxUM/Wfhb8opGkHfqckBK9oxjg5lD8iJgHNoMz8xP1p6NVKxoMxntWAZ
bHR3G3c+z+HGXJ/TMpXwXafywh2OOnV10FxyGun62c1IpgCKX6/pjiNuEKHzC8R7
RNCAqb+QvqN/zfSpFpt1rrXfJNWodA2Xmg+vEV8j3XhZaUDoiA4H+hRUDZBvefET
8S3iKinYeT1I70gZ8w6BFZw0VQJU4yadA0Ym4Fvtfl7otVK66hSUpbeNfl80WLei
Jjqu1qbTnmjh7xKTIWeTj9geVt4nAaQ6dhv0m3wZ2BovsW6U03lXxAfek+J2Ow0R
3eCz9RufsEIFrxyb98Qeo1ok5Pmbd7chP5zWWTeSz9j9TThSBUkEXc7rp4ZH5glA
6aNWXJKkjQnEmZrqAKGg52KqKVJ1vlBg9CTYBgIkdpG6j94g15Otr6R6tSbseima
jQMjdDU/atbCrSriVI/rcyCtKEXr8IsWtiu6vBqiknFl/j9C+i003Jrkd7t0tOa3
64P+nfbd10wcqLHm78ba9i3scKmhEO8/QbrtD2Ra0Fh/ECYU+G0Sq36HVHz/MqHC
4KHOkNGF8jkYx96Mc9NaDDhnXf+FW9+1pNDLjImkaY5/gtTiTHfgsOhjOG9GdP6Y
Okjset0wDjLxFzrJ15JTPp2Umoqc0E6HVxCTtW9ziJQFDDjygrilY/KpmzeCkkHP
rszlIXbK278MPSld4DEMjGFYmkW5BDd7lfPNSq6W38Ld05klnWZn+FgKVRF07jEX
n4Bu5W4wYL+0QCu+uSI97gcUse1FLoPdJ85MS55e+uJl6KnuCEuAFDH/yHOa4J5j
bzvEAxEEP8q49bE0yMjCV3TivntaACXaTr7i2lyUZd/wd8PLeeJqUwhH37rqXAvZ
Pvseo4ryBInjdOML4UQrpCSc1P+AnPXsfyPwPfgSLFpEeiYDcvoQ/jrMm0GIu4Pj
jA3KWJyzcBBdn8iwuZgUx0k04Pp9XQkXjIq5qitHQxLKcxvKsfpikEyVCSgPwD5T
IP5Q2w+aVVxlej+8JzC0kz19ZFmDTgYzxg5BWxIlJ3GtY1J147RTE4qTW0HFi9eu
inogxNqjDHbPcW7HzrGOMxmXuyLf0BSj0LzPVIZsIUinBHLMA5yfqFsEB0UOr3B8
1uIetJ4iB2M1VB2nZO/VuXD3ltVzxPuSkGRDjIPxCKsQUsX9YoYdV4VpAJ6ObveD
yEYwzgsFoHEJnDJh1c3rKTpFk41i5zF85wfcOeXMPKbERsn4s4/MVsGuDtlkNVbt
L9PWeBe/sLh4ZH/881oU5glvG9B4VQi9UyC/Bhye6F78tFZWd26JXhjRmW3eA2oE
0cbraFi0zcl5LCoQZK6vbYZ/kicHLV69uRs+DIRyW/yRlw+0Q3QB4lbP8xUb8Vib
RJr93dKi7KUAZUVxbjBnnxaEF/luEVHQxaXG7HDH+Te3++7GkGIYky2l0EaCAmR7
hq8d8Qup86n+I+Yc0rF67HTOzNx99RnFe4ZEFhA6NoL0U4IqS+oGIo4Mn5lohkwj
PsgxBLyqQ8C8biGrdF47a3r4unFvzcsT5aVlIXpZZD+Ypu2VJqSUDd7oHg2A5OXD
DMioqPZLukqx5DMEuZKoW/LCtkH6iUqoIknW8IcGAmAvvCc8IVKg20Qh4Xybl2uk
sYYTQa4m0OPlvxadmFlvu52ssWdwhbH3C8zW6e64jTYK2xTy7HD9+doM9rNyuyuo
Rkv34RNFj/G458xQNSkF2SEpOIrcjVQ7+j8KZYYQDhVktQjyBVyhhAw4nEHeY5di
vABxdKX3zpewOj+TQFilGO4yZrbwW6ReXmw7+BKv8AHFQtN8w50rVeIAH7cFpWRm
PwN3Oi6CC6odaYGHNVs3cvvMU9eGvTFCiurZwwmXO2SYipqzhkyP1PWn0eFHxJIU
TbAj0USgtfy6jWagyafmc8piCXbUClBmyzM4tc1PiCKNhx15d7kNqT3Bj2EPird8
AVvzgUtwDs20MHnCK5a1emaxQ3Xh9CCOY83auXrx7ZuviyrW3qYKbVwfvOWOQNip
XOSQRAK55UlRfhNqf/F6sv7enDAOi4Qngk4xEMu9segnsKP1Ck5PGE5ogLVEr8VO
/dQBRnDELxK4ZbOsLYIcQNtmSRmd3cs5+MIbOdbJ+9GMxfzN2xem1sOR1px6vNeW
FZydNY+b9cwXwfvxPiQO33guGRk9uBF68OUKKc5HUiMWoITqwVlk9GiMfUkEcJTj
kguGk+ulw0QFoILloxpbKmlOl2LLGsftUImiIWTDI66ibzerferL6oSTmbMWT5Xb
oFFFpYShgOX/K4PWV9h+fDoLJ8NVvcX2gA0xoBGt/hP+Mh2WKddMA/lW+DQdG5W4
1+hYQiNNx5TI/Nz8GGOSNTmX2YHOVDoZ82ewFp4C8HyE14vTTsNnB1jzTJr5WFIc
nhUfNClv8z6zYe/q6vC1QQPuWXsDrsZNULkCvhJnLW60lZseLTA6vQak4IhQMUL/
5wH8JZguqWMXtPQAaKV0iCawkFRKMmoJkmdIBjQh0H8kS28qMnfQgcNihGjQYVVh
sk2dFQojbm8BgXRHFjPraU5jh5N54pu3o9hv8jnNPbfx6pz9/uceepEG3JRDOZaD
QLicaBlUBmu4FznDj52chMjvKOMPygVdKRAJQnOFr4RR3TGjEboA8JUEntiRljE4
pFIQxawk4T62atsZeUlbrdL/GkkDGRVM4CFi3o1/4uIyZo0KL1YnmBVyAKCN7+hE
MeH2z8bcsobTGkbZYLMEnECDu/fUw2dWCCfZ6tvq67c+TPiL+uMxotzlt8FOEjWG
1f0Q0XvIIbI3Mr7GXqYcEBn6bWGEaqaRpD8Um6jFNo+lzUorJqGiiSh2XeKutH/O
lqRXMtyllfTHDBD1zKrX763FAfjueWBKka5ozXGgf7+A9nYrMVfg2/aea4VXlQAk
MXF0v3BUFNeOdvbaswTNvdeFc6dY/WGjMjtNGI0VM0OiflQw4bu/PbgKnP03hiqi
tAxeo0qS/eQU4pf32dN16KuW9PzdGJGggxeDQHcmqMiLhrZQ7Z4Ji37JMzHwrA4W
eYkERp0db8hU7b9y+bGoBM9WC2TsaO437ZAWwGyznknvC9kV0eEtdlcDLtwnt1J1
rfy7lnkyw06vJC+xftPZv26TCdJ0KbEeuSztCAyzBfoF5I6WNDA4Vk77qLiL4x5O
nA6FI0NtizmAxn6XWmGfsE1iJR2P9DcTYc+WV+W6K2UgP0/VNnPGGept16GLaKol
vGaWvF+X3e4MaMa+E0T3w4bVX5AHKChAQEdFa4Zgn6tlIWHBYAWPY6VZIHXk0iIv
3Y1+5KHjMulSazv5I1MbMN0ujnjaWc/dSCFUyh9nId1ka/6zHBFAa0kZGpM9oBv5
HgUZlIE84JJwn8bv4LOsC6BhGv6Lral8vd5XzUrj3ywxZacP7U5cXXxiaj719Yi/
/XJIYpmaxZQh+xPItb4aEPPePogNWmcw/Lfp/vjlDoKrqEP3m4ubPuS3TuQC8/+x
nr0Eqxivs4wc6u+C8K7SuWth4+Pq3JTRcXKbZkuxkXLsRy4RmrAptLLgc6VG8h+N
0prnwAqjIB6CJlv8LWnKOgUQWluvnKgMdUHpiL73bssUslTR69YTvLvAmF35nK84
ZDtiVdR1kodjXPnfFTHHNmg1VXZvoZ7HusxyxUyoPCmEXTKu8V3/6vo0FWdtsn/C
MGkiaCdcdOgpTqj7Q9S3bBRFszq5YfdaHJz3cSr4elEUdScs5LuNjSdbP2naUyfN
WEMh5Ee/1Dxc7DuRKHcOYFvjQ1+W28SlLOTRhq6KCYZmHvV4pz7+oIvsDwDeLq1s
SoqA6rW7ncEHMdzMKFOL5RSczglINlkIALkojCK/g+hh79X7R1rz432z2NIT3SV5
+KxjwN3p0Jt9nffsDC3mOiIwbU7AQNo3IIhwFTk3mCQ7uE+iwROwYCP01CSK9ow/
ykPnchTULZjtNB/g6s6MLXoZ4c5UKA64Vgm+BvN3J3s4+IKY9UVqYF6qAgWcAgIR
aFZEUJRh6dASbSOIOFDfFJRZNmi/3k8PAqaoBMYCZ8/gBMvWXtTQqKRZYidT35vr
rLdnC/Ip/Oks7pJ4lh/QJdbl3pU+iAS0h9cyd6UA5WXI53xcCsyNNt9DOOgmRbbp
d2eqlyX2WAOXkVnD0Zjon9L/ACZBuzK29a7QRdieChTAOhcq8KEtbc56BKFV/cY6
Q0pBPcSgijqGTbqdzRQ7ivNOw0uIMBRHDdNrRfkUQaRdQdTEXNAmGOGJ1HjfpYxl
3Tti3nol+YWT9JviYdDyNAmFPPOPiLO6lB4uHJOL2ksxIJpWX2p02BQDvzGXXBc0
6C7z0HEq1iovQbXNh9d6WW2cpyu7Vn5r6Qvo3AXhZF39nEjqeRIl2P+o6gvZ5GPJ
vMlEvmAeRbEtC1596clmTB3SruGTquPGjMNNe5cwBfaA0qyWvxjc3vxww9gzfoY/
vhhNjd76wQcDRi4A/mPLbr0OIeqdU6c1kR6rVZoaXUFKD2UPV25qokeVaVb2MmVo
75BCfRB/3L2LtwrYOzsFwsDbBgK3SGjhOTCY4w4LJOKQjcmaYz4UHzOPvi/Y/12W
3BrwJox5SuD9weLNaOU0WZKQo+so+HE264NavhLSD5VNfYSg6LIk+C6eUbKetAOx
r8ArtP+sUBfTD6teujoTl+fNNvwuNJLTZDjHowY6W7sIEmqi3ogho+6bAkyWL+Qf
jIQx9zgW3Biwc3Z+P354BkQexoiqlqmv79VsGZjoVTBOxusEUMn6HDmI1TPQMU0x
qXxtzAOg64cfhtdHFz8x6yVfn49gmKd1yAKiv8YMLl8O5f2E4CZbRcvmmIzVY+dO
8HbRqNO5pYKS9qmgvNyEf5k+Axhwxkpso95V0REeG/PZ/Y+Cr5KZaEFH4ihj+WWj
cTYUkvqH0xWUu6YwgTABl/T8/ZuDtPWsHO/eHx8YwYUSeeaz1ZRP8t8FSwN3abvZ
RruqGt53Cq/QKLSI+EogtU9AcWqCVvbr66rzf8Bav2xdDVnaN7mQmgaEFnRwyjJQ
ACRrDBz5V+eMflcmp4oqXJOL0AlwbgOKC2thShLZFXUMjh1zoN0mOfhQLah+c7NX
4GW+irLKUkWq4hNbj792hLfZjUC9DZ5Xo4xWRligZ1CHDYisZRoSyCig62VXG9rW
Zp3qCZY0oBQGf0VOZrpjdhXdEvsSjQIIOp9FPKU6Ql4JNDrnbS3eKS7kdvL7rKYk
jvxb4MsirGSN7vdmwAgs91t0YAs+Y+3e9nNBWMyvZn5t4TEVyMLGKthq/MmcCEsc
+vDwvcJ29G7FKGHJdLxNdFw1pUyFsaYJGWBZsyrxJcIQWASzrs5SeOQ6CT/BZ+zN
mx5iPpYdUx2wWH0BcA51XApYM6i5zA5x3movVWPb4cLQ6cyPiFYGB9pFuaArkuV6
aOQ75AcvvSRFmaF0V/BtH8JYOEK9LgC9L6+yHGdLmclA2Q8H1kUR6D8bkLdaAeMu
80dE3KwWYmrHYo0QKOG626w4uiofojwoHL2jgWsSnWpq7jMS5DZgCDm7IrDNpsFA
S+rs8pUKXQUI/JkKUjy4MTcASfTYdMwQveOM5knas0zpjA+6ACGTTerq018BbepM
+D2/R2zmPT9T8XqUPbDJMDbhMjp0okzQDAHn6EhrLu1w/hoAijF3n4WanlzpqN1Y
tZFi/A1AkPMT74QFZI6CJiRrM3+25WiS67EIuDda4UiWRiUK6QKNNDKpsI76JB4X
eghwb8FjXwzfV3eXGq28evAWR6W6tQamWDeBWuejN7MG1Djy7x+uU/HlZmfK7HZm
RT1XBD8cDjWuZV5pUDxeQ1If7s6XEwSkUQ36pFkAAsHpfitOb/nsk/j6SecMbA87
J7iXsb1FNQCL9V2t5v0/shmlGM1Pvp9sh/sSn8HKmufAdcIewp1rvB2iNFjB/dzU
EEehj4w0pRBe58QDFSWRNAIsX6l7ROOW1kdvHugaHjxoUev++Hs5/A/pFsvhCO4Z
Hm8Q5y8NKEEFVzX6Mnv1NbGFhf7r46cHCR2BDrsvsCr34NIFlYD7ugRgjKyngddb
o/cY2zgonvSTGeK3KvynQClLnON2mS7geqPtf0aElwC3cOB4HRiFF3fZmK3nh2BT
b5frTff/4/AX16WvE+6Q1XSR7nV2FC49D0Qj6ORCzH9FI0uk3mUciJgyJM3yp0oj
YBXTQITVqDVbm7W/+wjq2JuVsTONhA5z3vVJN474BA9mw89BI6zzCWE50lrAKrZy
8Or/iXH8SZMTmqinuJDhW+HaUGab9eAuoGWzhWhgCqGYd3KIS4G0fSLvF6Ep5+7J
1HZclpwcF0Mu0lAkzuUF9z6rlg2Ee4or9rY7AKIxozBKhKFQNbtYcXJbAurgyA/y
SIrIUukQ2OQFg0UZYUx+ufH7LA9Q5hxdUD46WXY695YWFYmpOJ5EXkRgpPl4mG78
wDlt7Ik4KJYQnwvMsguuANu6Tsg+Jqad/QgaEhJ/i/4KhTsZkKgiTeA/uz78V4Qr
sHLkoLlMOMlAF7QSrMZOJJIMsutvJ1izA3pIg7Ne1GTp8i5vVSznphvdvDw3JcEg
iqUu9uJJs+M8DYKl0SQQGuFKM1i3xtK0IcvrngF0tVY67Iu42CUpXaszaw/TfArc
ui3EXb7BPrXq7b5roWT1xdQUr8aZXSH7biXk4S+5q6Qm5sDtsxA34XAUSRgHJAQd
rXz6HO5lbTJY0zt89z9NiRzLxG/0VYYkSZyydj/JggmJjqC2xHQFNBsO8iXO1CtR
d1uSxTmERP1hpmiME8H9vWraG0re9wk4Jv5gCxVRVYvnunsLCuvY51DzQ2DeUGwA
cOB4jp2XstlYqopqFYAeP7LiVHeNIcu+kRj9lWYdsMjypZ7gz1p4Ol8I7oKKJFcJ
Kh33pcGj8aqta7QOIBQNh/81b3kWL0qZC0B8d7d/+Owe2tD+PiStvW1UsQuE4InD
cB4+qC3EX4nNPFmdIdQz940AS+wXfQDLp9v259K2at0Yu0BM6FYzbVLb9/wu0pS+
zubsO6ELjJn+iAmI7tuj1BP9WVg/CTJB23lTKW8tioLOhLm7RoO1zudXkxO+f1X8
WoOYWeojHAhwHhyxusHuG6Sf2hKSC53iUXvuw1vmGQEO7MRJuVTmaEDyNwf6/U5F
6+aL5ohb+/61WX9JW8PHYoJOyhhgkT/YjYHNSJbXn0L86zspnw7++Y26Q95D2uJ9
D8on+WmFO09vOHWoyAA9aYnnD7rOqPByBRA5cdotyp3TrXoV1Eq0LCF5kO7tX3Nw
ZB+YaD265Dbf7ah1sIvsIy8J5CemiAkmyMnm9b0s6qsnw62iEqiwQYk5ZMwrT7EZ
lbbZGW4weVV6m8AO4mdw4nWOJzsv08XP6Vg3BA7hNNPKRN8PNBupFzxCZqaOH5mp
Lq9RfQiIjU+DVSB+M4TGdf79j3btE50xGPEdXR9GIRo3cmHu6HlSRyrWhIbldHRH
bOQ12F68iLfCCx4IKZbrejEXnZunYdwZ+LhLEV7mmvG0s+1mEjA1lKrLlP5CI/SN
6kM1Mdr225gxmUyhSPNHUoz/wYFpUKva3Z32juOsTBVqbwMg++kc01TLFYeAXTBJ
5xKDvV9HSv/F3b7QD+6eC9XUz640KWHZaTv7u+8MvK2MZ/+Lt7ib1DRlXy7V2G8j
/7x3qK3luvPFtm0vuJxNFQFXTILhZg5T98aiSKNQmjV9hMqWjjDGNhPlsDDwx5KW
gViOU8F1oPuZjMf+wNZXQkcNhIBGKC8MwX/cReWzKApnI04nc40xoGC/lZ/39j/s
UM1tElte36GefAaeaxwmFtISns0ZcXRymP+q9+tHCiUshF7qK0BOwIVVmTQkeWP0
OPS97Jj2mLwDbVkgQNcCEsztGYItAO22XeN/786yblG7dQ3AhJEXzuWM3tJf1++W
Uld9QNGcFZs9XifEQHvwlnzGJSHGuJre/w+VBV9LwUpNoWdcxYZ1RBztj5l+grmA
DgWTKoVfFe+MoaKNW87h64BhgEi5dZ6B9wymvoZsoHQ7wY8yYdzrI7FoBZMlNZG0
WnhyfbhPs6kSAM9KR50GyX+QS4G/UuRDOJIzmuDF01g7ODiiCAbC7MarnNxZNjZs
1yxl0HrDJJfy/hELSbC64fVruF5H+pVecaiHxuVien4=
`protect END_PROTECTED
