`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nXCvmuNfwNnMr1d4vkbWeIeX1sp/HHle45ZJ3byv2mmG7kMehTuf6XoeqzJOSQn1
QR0+I1Vo2TSxtJ6Gbbcb6ool9r2y9/6lQkDfPUJZsiyCXXTrW9JZmxBt6YdVi7UU
21qSH7Ein9V3re9zFEJZR7sP5zDCK0Gw36IMrZajTN9rSbk4LC+rp5nGbjtm0g08
F9rf9wFVCtLkZFRVJrG2W+qxQDQ28ZremiJmnw/gs/iAqaWpdnNyaQPhhgcEwdDs
/UdDs8J34V61m4MaQRIsiFiLXvpW9vDMNFtSeNek5PTG5rG/nNhdP0s3WgBpcO+M
t2EHKgi6EnXGybBHvJM0ldP0zj2RsEMnBg2Xl0WT28eqg0vTeTcESKUv39i8gMLd
CkSLk8sqvV7tN1LIQfDhcVOTtEoHQAtALZE8+oFp/fstVPOy9LEXDDDsleuK6W/O
OOYXK/mpJrsl14kU9jIN9ubyG6D1dF6rA0le2p5g1bReMkMM+e3KubtDtRIZiRGH
qnodBopV2y1OUi/YUE9RFCmaMTXBv1W/wSFnx6upM5IpHF25XKlmg2Aiib2FtEnK
+fWH1/a6QzKgqJyYgZrORA0s1jsBOamFzIIeP32SqmgpY+/Xouoh1+DDBHnKdA7h
/Ky7TUdBYCO8oJgmPBgd1PEna1P0CrzfMk2FfL8oZFhveU7WHOBRGQUJMJ5quAO2
CqDnqXCvRT/0qJdYjvFQE8C7ECWTdCPHbomKWrEZcbzhdYVaZ6Epnt19/+RGUcxA
o6dZdkCeWyjP127R61d8JW6wfxYYLJet13Fil72fRVnzqNxB0g34RsqHr/S7vlVe
8N2igV/xM6yfM5NoSa3S7NEfevz2l1x7CnoAFW3BJ9hbt9dz6tPdErgxggRRkowQ
E5Z7zXbDRQb6V/hNvgisP3k6aclv5HybxVXTnoG+/8ZGQkcMAORRh5HovhkP4avI
IeQ7mq4yYvgsDvG5BO25crmfo60IQM6bdaZKcZX3mYdTLhbz/OYxqM+3VMLLIszI
+y9jm+FVbo1ZKWrzfHR6OzaKLRPT6SbzP9v3uMI3G+mVyv1jrL7AY5/cAV0UyO5P
8P+ci5o/twwtFfY64TwEKgMVH6h1rNyIpYFn7L2oNGReMWBwNhhEcAckTiHNtgzZ
tTeDO64h07XiUfglPiGUViq45U8rCx5MaKJjkmP3LnTpGxAdGuEel5s61MGIm+7t
BfjCBsQonrg12d+3ulQpuY0eUgOtKYCR+v8y3gnAGPd9v5CxcAL8hkWYJw2+gGcj
ajyH+wLReTlkTduikCTOwqYlHNLBUNFYn6kYLhbgtfp0ucgtZTPwEfLCkrVEPfmw
xbNPx/m54du1BqlQYEoV4Tk6VeHpRJXl1iQ3hlUQEx0u+lLAa4PyRyRbQRcpdus+
8K1O0ClEKadzimxM/90byBUMooXLlBMNjZCPgli9HSa5emIDAZKe+5ub5Jx7zuBI
dUKw18Xz7wDa30wlaERcYi671O7d/W4C4UX3Rqjk5p9GNeR26CsAZmIcxWRL8xXw
W/CVu+PMX+9tmHidhI8pu9PCuEoB/tXGII3F7V3t9/eLUGjQVEtyQYTFiZBd9Hp6
falBTfcvYhWWx3/ZpfYz1hU5fw0UvOd3YavVnSs28S1iDfB1jqV0Z3z5hR/XI7Uy
qYLe2RBL3e0PDFYJOKLzryZ+XlHIsyBtK60Lb6T6uy9Z+6T+Au1b5r+XOXoEqw34
kC4MpIyU9Z5HuTzFHFsOigtqY9IcVqlygeM0HFRtv6+IlUHTcoA7LvgBwal/jbLr
dks1L3MQtlciNM3QyrZIlA91bPdMGJJoyEa16h5cj9U8mgIDQLZuRih1T7GR7CAL
7EfcWkgYQ29p7fQr4roKyTwCq1rixUQRDAv8wKz54POjB4v4MN5hh1OwH5bQTz90
G8IchSfS2Fhz3+VGO4wfQtimpIFJzgG3G+whYb168XrGXz9r0IrqtMeP4jwcFuf/
EVr7eYqMR0uN/AQIluwlF8UHYmR3XBFAfizcJtd60affcWquZLQ6n+2VaaG/dflc
n69imZ0QP3loDCAZYBXdgCh0s7HCxF5zHPUVfsS7SEVL+YQuZLLBPohvC7Dv82fq
q4UebKaSL1YXVTkXOHzgzhtSw1FcB5QTuAA3h/T3x+MXdPETfB+18E+oHmb9NY24
OfziVtX3Lmn4eJEeFVbmiNl0cfwfKpOapKfSFDp7zaTHp4AaCFDBq9bnjp/0KNY4
PqXK9Yao4Xcr2jD5TGE2/uD0bXcG1TTjHfXwv04Lz0frbPHLwYXLXAchM4IHRPRF
9EbKqtUTBKFT8OJEf7Aj4inprSF6QbycCdctDBBko3NafQy5N72KkWDlw6emvlXM
JLZUgHU+z3CY6uiIpF0t4kIxZgVVEm180AT73eLyGisIPxDDUgpZyjHmgmhaI/W+
Cop3u/6jtUbOgAlA08fJtXRDqNEnFHPhMSHELetKkav/TJiNbkARxgi4E/uwuHio
JEcp2y96q4mYh4AQydqe/Bp1uyyOBACaK34E7cZ5w2hB7hlswZsThsfzYbcYefQy
eI5HZgSdLftX0WrvdeyaFqcvwLXdOQHK0ELwHNMvR7VSjvxItqrgw808wyPhz9Zs
5AH/A20ZiP/85ruv756AgVd9Ln/JLpB1g370RcNbrh+rrdtVrKk/8f2tHzWHMyTc
Ck2rk9wzTd5QJru+2F6P3LTI+CguJWxTQUJfN2K8vRT5lCilkMk9T5Y9r9f14IW9
a3Y+qbst23SO3yBQlK1nUm9aXQ1z3r3y3mtmzA3gENkqxX864K0VtIhGWFGd1CpN
qFuU6ToS5zFoWPJuyCZwSH6vDlMKKHwp4PgB7mBAyQblG2qAm6oIPIrrgObTN6pj
pgIBxQa4c61pefjZiQt16hCzcd+XCRaouK92c4X6aKXgjLEboXJ5QWDHZ0i3KxrS
6iewO4r8fRqr4t7WJhegcWCXoTspFIZW8+rjXY8qx9Bd4DPcZ6OhehChcg7to4KD
YxRS5rhSe0P17ZfICvqvUP9pGZnSnszyObvqNk6ai8KQsH7cSTg7Xjls2LNsXxd9
UagIrbd4nTgi/TZ6X6AjLSLsywT2xIb1O6GhcPa7CxNVW5BiBWDQbbfoiJ6TWRO6
zyBFzaHgMCtY8TadU2rqdoff7hjPgjZPBvSvqg/TcG7BViTOqWfDN4ouqiQWi+cy
15et8IyIGjzBiq59TeoFppXtRqMtaDAFjppvRH2V7A2LkLWQpNvecH1PJG7lEJHR
jgJB5ia8H8Wv1UP0XxiGa3IYBQ+B+NWRaMPmwWaUJ/R64LIeX5trV9kCfCxTf6Nt
RvRe32F+8/pUPJWoc42d1So5B+5WNZ81zeKr6zGy/33chdEFab/ENioWdCqwgqev
aENlw33JFd7U2VFqMenAFV9yJskbFON+NvtQxTDQnwGwLIFVmI0a1dCO+RNhN01I
IforQQjntyIojL3gxoBIby8c5Jy5U/XrhB63/dwxMqR8dC9Fn5rMk+T88/K8SWzb
XxsuZi6hQYUs6OaWXsy32PZZxfdXbjOKgJLx6caNJ4lHGh27oYbM5OZMJhxzxhLf
DBwyYz+dXDsAZ1d5du1xzwhxTO+FvGlFo9jXLKAJVfKTF1zWYeCXE3lYRb9qLVe6
p/WPAKwrmrtaj2bdk6LA5XKhbOwb8F1TWFTEfuL/yR4PgZHTih3fJvrM7gi1nfrc
D5imXrtO/5jYc6zjx6LTLiZKitcTsJ4WMiaGeXb4yMeHFpvwzz7hd8+b3BxdD30J
Lc3iRWVoBVf03DJ0ypC3gCmWG9U58VNs3bDZZlmoMcQLH60r0/urmf26tklTSw30
DlyrelHrScpCsk42ACvYIZ/4xaDpz/xtPyaAtsQETQ4eYALV5RdfqqyVR5IwXeYz
IPHtGEdwWjS4vp8ougUOY+YNyxpUKZ66KiuH3JiorcdDANLL/RHEznCC4FZYBeFX
/k7B+/RP5BN0ipWGNbTaMT9BQtZYy6LFIwxhzWHvR/MV/i8UB0OVhrbDhpcyrzhG
tfq9waVAS2ALfK1Sx6iMOwvnLKWOEJtGoyIKWYigz9zMq2wfba+D4QKd5Hka/iZv
nkqyCK77QWXwL1Nrf0WuD0I4vF4PEmXWmLe6CxfBVhtASCEAxITnkXy9JGfrWkKp
zH9VkRKG8EZDaTzscH6767R5y3a/VFxrv0Vp7wq6YXVLudnC3BdEx8bNEA4Vb6NZ
gh5vuqNiPqXQNK65U/6BtiHoqk/GvgxndhvB8M9uWmagECV4rb/iUco9lhRV5dpr
OBZg8JX8jVicXQWiY4DFCD1SmTd4nOQl2herurFrFNj346qUbguW6p9+n15h1dZc
QrgYYC9+QaDTuwxjVNfE5T+3J9ElCbeObHfZ9r9pQ++tefXxmlii3Gn/zOsdUjzr
si8U42vrKrCZbQwjcDBQZJ4sS/6oKgcQZ7zbag72T6aY26r/DgYMPDnvH56ys+wd
qTLg5suSUd3QMqeB+anjf9ybTZXKlsPNJXMrZ0BWIgNMjZFzKoOHpfDSt0LiKfnW
qh8+7HwVOQydXABmPrExv3NjDtPvwEN8uyvsu+81b0MApU6u8QugMF5uSiLjflm7
EBWRLbjA2LLCZqk8TnsHvNo4OLu7NznxoCnQJCz0m8/65a3Bq2q4XzgQHJ8S5q0L
GxPtHCc3Zwl4UbBY7HKCs9Uyf3B3ek6kMdTKNkPvdrim6Ewbwq5hNf42Hjk7c0Xq
zpnAp1zLMYbtD0iLtwbpD5rrmg22Yqst/G65ewt1ekB0zTRynRcW7kql2tee/rG3
er1qUnx/etCBCJQkjJj92XQ21uln/YCAR8Q0ZDlsYoJSOeZD0dJAvwV8AY8TJvpL
S2KBDoUDFMpNFqtmXyLe+6A2CLDU7aGSCymZI16K8O9u/pDYH0OA0oGtQuzT7rrB
HnmuntoxcuS9il7885rDywbE0hb/5xh2LWJzKIBUDTtpSQM0s9IyTT3QXPNcTXJX
snMzavmT42/ExtTyMU6xMOJEYGtIKkSH/dBq9z3feoClcbE5s96njcsowv++cYcS
cWqvkR2p3ptJVT31ayaHtkuh2u8IRzM5ldOEJyB0wlxqrCQElvCJ20mhXY/2x45u
8Rsn5aCkJpohOsMMYbxti9lkzjDD53ac8bAoD2Kv/ybfNl1y2UyQJ9qc15KetE+i
FU9v2unAsJQYTj13sirz7qPEm9JdXsXzEobW38kb+nGI2sToGKVc+/V87rfft9b9
a7pDf1oUIqOVCkgRpd9RNZB1T1wyHpwA3C8d37+8y/siskQP45Jm4qb1b6EEEHLw
NL7TzhgVySIcAXwPHdxWKEhLVWZqISkzYHPmitd9UAkZPEnaxOzy8nVX7sqPO5Wh
OCoaocFw8y1Jji8OybaKxORoQAFOrDYC9KqJ4QQ47HcRAdPEuM8YuRMFnytxKv3I
HtFmUfvgiPN9mWBqrV5Ph3aJXzmZDcwSzWnh+RpJNY+yHNVH2hybVooe50OiMefB
AWgP671/EneyUjJompwV3788OUS08VdBS4ezQWgPgdW59+KUwvaA+9a2JcLG4cbz
cpgXa7jJHZ8234P+Jk6zZkBsanYRhP6igze5LoJ4jnqaJg0Et9QAxTvxsQVlRTbs
CnJlfG881tsau7Se/VS+nfd53suoKeMGHqkB07InLDvjpRgM1X+++MS+Sxj+/qns
E7hEddxk2e2D6J0ic4MrYgJ6NlOtM6mJzUwLb00Q5jnaV9apsekLp+aUarIqFRvG
8BfITZQwSSV+o+WSW53hlSA+KgYZgiwqWFXQF2hAABius8ulXlvRhwxfsDwjqI+9
V2deRRAbJHluyGffjwzJVb/Vxtr5r70EpWTGe+HWK0KQptwoUM8U6qE0tQMTMB9o
gBPBmCGyV2a1HUqj3+V2L5uUUAA9Bi+yxjQVefGHtOBCFUkCEV16TQ+/9Noe7c/b
pz9c0jWgdWeSSQW/prF9RwyYf6Sl0xhTpDUaZI4ILaO7MLpbonyAbEmgnfZEr2Tg
Cyw9ZxGVnZByfjEHA9WbD7826Ses+Ofz77GFdGC2M8fUVIRE9X7cv8wgKQHieiSd
O5LthkqTYCbZt6B5PzvtqGnerg4bflo0ris9D9k9lwaYftvwDF1wydFv9xmoAyRr
OmuyeuVF4dlHTdEDrwaW2HWbQDcKt3WtoDrjFU7RUwodnwVJ8eko6s6RD9XJdUCA
88u1BA5GGCa4oI18CH3qoW8pHROuJv5twVUMpTZ1WEQKvCx6qzZ+3jPiolXp4Qgy
OEGSoTh1E6oDNvuYoE0Qj25cfGF/8eNIOMemDgVE71WccLmweuyrqB3hVtbfrkLC
bRTW7lqIed9FAvQ3Peu3AaIzvDTvSyjvf+tH38S/W9ek8I9zFVx3IY0DksTaQ897
g0GR8yg+av4WRA1hyyrCBQiZeCppc/YJtqTysn99xi1N1o+K8qsCUTUTW6XYkW0q
dyVSXsLCCD7cPYaFG59TpnGxcHmwbtkDfeiFxP81MsVG3OhDdBxWfT+rOwHOivm4
JMFfqwqaDUkjv4ezFNOSogtSRbnUqN0COPEqRFlRa9Fq8khCDNXq5KLZAGfrlxkD
N7c8bT1OIQ32KUeLZbPBzYKXVvo1yz8MncUBS0u5C2Tqi9KBGPDKvUMcDHqhIF+V
WTIdOGnn5JFkDzvASMbpnmtKFat3s/dMGoiFK/mzwVrpUrVnPnDTVNpsbh8KGCiK
Z9xQHkdjeUSaMWolS03RUYQA43iGuhEom3wRuJbnyFU/uQzc83o/xGuw21Y7wJHJ
hi9zrLF/AaVYhoWUiUuNZbFBmDkYuvr5qDOyNk4RsXvoE0PCJrlCb4gWDRO8C7s1
PRsl5rgzmcdRrRe1wNFuFXve4A9RWDJA6roZyE9bBVCJkjZw71c3xbEgX4d+vWSw
pLDI0x+NfR7Slffs7bGSJ+kEnB8bjC1fmNNzZdCq49xWlRUTMxDEvgQV5fDTvflm
sYqB+jDNfod1CXqMAQYxWChqfIRkyBJmsvYuXQZZ7Ngyoony9OF54cPkezAITblR
jJ2dRFXdyMQs7TSSSkEvBOvaRosdKvUku5DXenA3XIzwCwYX+285pPVvpmttYyrC
sO6ky41biCn7NsZdOsRra1ujQu4icUIM8Wb8BLnIpeXOZo78j0+uLWDEEvRw7WPz
t9wVnqGAHdp21+glE9g34o1CQDILmmhY7vOij6s5iFsAZNSfa6QkWbitTjTH9P8Z
NOrbqB3tWfeNaUtrfgg3w8RcdsXFAlb/fgqZxLgL+JHr/mzsLlWje73SptObTqxX
DBFJpVsFTg6AC+MHLRnw6uYkV1AYdxcuIiwjsFgMvZO053qAf73StPgbyrdB3LH2
Fa7zu0Cs28kOx9aZjYEHlH35aT2z5N1mFwKNXS1bESX9FN3yxR+xsNFBt3FShxqn
c7898nc6fiPwOzHBqhKZA6/T4XtZ87+vMhF4qyejwqWaN0hjBLKWEj4NMQjseEtU
KEUZh8ebPAYnQVnhf/NBqqncX80SA/G0xfzM3yGpjNO0ynvYPMXa29wFHQ0PjisK
HgY2pEDg0ylLmHvcb+2NquodTCCLHTz+ko4w+L1MA2cT4VyhOzB7OTftVYfF7vGf
DhTIytpWoNBFNj41TI9uanEsuwr6ayOfFacnlz+ILQluEFOfVKC6QXhTBAFaesGI
NSaCsJP8d3KO2Ltl977jo+zyzL+cUGwUuw0aFAxxnAVum/KoKsQI4gQaye/G8Hvp
Gh0a2moPrDgALN4aowmLqUTXEvnFNicgpG2zb3K86BnJ67Iw5lEzidH+mmMSnyQk
g/QaoTka9MIGxaPxhNP52tNTMdOhdkoAWbERXw+dgZOU6qRIBSBCQrKo+MWRZPjG
Nk9STJOLHY2lrLY68RXXsALfYjEPAhR8ABBSMfe4wFoldg3tlJGSqjold0wDFZZL
zilvh+7N0kdH/rN1cr5UN5HXWqoyWyaFwPW7rpNB8LHlbi2o6qUsR8qkhXDHffOo
PPamN+p0XvJhI/bD4cu0WeBy5bKUCmQLc5r53RDerakBpIqyDIllimQExiVM2X/I
UaCFy6ca0UU235uDh1P9R+sEc4SJYYYHN8Arcwb0DIEvCb/97HLteFDLizkPy7sr
xT60BRW6ksj+V5kH+fIJPkJ7Uy6r/+KF0nQZbG/1CNYwwCQrnfJXDxdAYcsEeOz2
9vSj4rC4LJTiWuN/GrtemZ5tETjU2ZkPv++1ejNmjJA2LG/74pcxy+u73RxBnngy
aS6HTxKFlEpJHS1JHZq2CHT4VkqoGQ5AQjfdSeENCYNP4T/TWCJx2eqn6dfbyN19
nlNxd3eHPl3eoOKqu1fGS5g2L82W6PxmrY2lfl0E/Ieuv5IKxSMT9htbh3S9Cpuj
M/ybSUBMHJx0OdqY0zsTdHHJR0+xVQeXffa2XQ9hCtY5EAC1OrJzho/QkHone1zt
AVPbkLb6uFRQEQhpZC3hJWmYLkaPwBPpcxXhjN07fm5SyGzjrGGGBA06R3DvwvGX
NepJv2OSSIxLluz5bWr6ez3H0xzM+BSY9VYRL+XCiTVqrdvZ3WXibg/fcrp8Vib+
5lQ/HkTjOgdxwMmbSVpwXZkG4aNiewVGmkOqTXPgahFTrE1Y1oHpuDMFcFluVQTX
yO3vAi333Rxozhdp/O2ctexViyv2KFjdvhBDxp4qJ+I6BjLPJ5+udozWDNihrtLX
qOp4K0G/JWncE8Y/RnRBW+pSoxDWm0iNyCgjfOEO/dwOe/yfbx6YqTnN7LV1MdCC
7HsR2HBkQAXwBeuYy4SyOM2LWlOuJbz3xuytMz7l+03p1FZUJXs44rjOyjlWRMDi
GVhMFNOISJ0Giah/ZrO6sy/VXbWANYawKWMhOA8fqcUy5kjD9URsBGi/x+zgeoVF
gpZKuFzoAabPqCXEazFY77skE2FlqkN244Wc0BSxWUzjRHNz5LJj/WirNCW7ujM0
LtWEGg7pdL96y2meQOazLlzKzwLz6dTpJCW1y/jgAGM9HHyk12XA5J9u5zPcUZA/
0UqipcpO6xVhgCEr7RxnIRQyGzvv+QwvHWMJBncWLhPV7UTZFBT+A0q0BYTHydY6
DCJQtVqm7c4YHm7Jo0JwhJR6HUHMniUPDXOkZkX7Rbyff+V62x6U5hQyN6iN/MIZ
m4iIhRWrKSFeg1X7sqtETAIoZgTL7QkGw7AqegNymIBbEtzig0qPayt3ePaRhOZf
+51CipFGT0En+4mO1ORqex9/Tz8/9UG/u/lroxhbMr/UAeH5ZEs0GXTuULdMAt9Z
QklZL8JUcPiRTaSWMqhIfr5h+a/gD6XfeKWsuhY/jIPQ+yDuAasjumRndNKzMrxH
LdnRRu4qPhzzcneMqMc9TpvazoQS4urFBK8DAH+Zjz/Uaxv94wcpDf9vYUY1cmMZ
RzoH7/khQJRKAJd2F/lGBE4A9pFm7JZl2n61e3TcCZnLviY0f8Hs+JOz2f7iJts8
Ej0K7tfcJG2yCFZO8y6bELNiMX3V4BdOckwV0XKmL6BXLuY0PE++mAZoo1Sr5ayE
OHjVRxX592NmoyFBSxK4a/K+uNfkG0uiYsrIrKNgHFhVJP7/JZ4AEZF593tWYrd7
0CfNl6giZLu2sF7lMGeqawCBLAVNqCtLsMG0b5YwmBo+pq5rgnV7StxNWKB1/Hih
KAbwMoWGlmyKwQMbAXMHOAWRisyADV6iM9X2iYIQxfGVfAI0X8NR31HDlL7xFB4W
fA+hZSWv5FZlfNDvF7ZEyy1ejy/YblFD+WueISSJTcWwi741ZkAECBUHJnF/enaE
sJFeIAwj/TZgOBDeTrMUWBSEBK+QXqUe5vJSz2ECx7xhjT2KR2CWLYLqJUxOyzou
JTi7U+Xg8FNSVo/E6zRtHcyAJW7Bbc8/P1DcUJQ7Akcwkqzev19aC6RuvydEaubP
cg4gdbxhMUveZTqj8baRZMaO6MQOFcC6JmKxEgugO78ueo8FdVNAhnqpbZjssYjn
Rhh+Ry2oa9/eeRo3uc1OtDO2aL3gbx15cYpgixXbqUFXx1uZ2zl9PZdsr8jMGpCu
SPPjXazJ7JOPeamz8cAwnqEcbhjHadOPKm3PcvqGLXl4waJ0d77ayZfD9G5Ufr7V
z4BUdT7HUxVJs/fyd+LnUEQwpCBcRy1siiv2W98XaBBAXvZNUz/Fwx2MxrC+rcsF
EsleWwwDa19OzzDrf3kVmz9Om3+aU97Co4Ou8Mqyt6QzX2gF/seXkq6Sfct07J34
svS4a1hSORrLisc8XQvZZzR+GHiXCMdjenooqkgc8ZCK6MGNlWN5yux1gZFcVzt2
Ubv48fpViifRbsDVCRZ1ReKtDEZ+ioDBG9YA2EWE9gzF0lF+3Nj4XhtrBlraFL+5
62WHamwtKTStxVGj4WdEKsHqAfny6lkBVSYXpPwlIXdmZVJCgVl4qAdbksELI71R
CqvsKHZX9MhvdS0tOKdZ8XkFdBmDl2voW3yJBa1MC54FpnHEt03aHGepmqoIKdHM
LHrql0OD+moc3pJtNLXWny6EERkc4WYRpO6jCd5XfQ6e62NCm11wp4DDS+XyvvMw
GAdsxlzNCEjIv7PLT/gxFkTwUd7ORznC05YNiaEQWh0Q1/3k5sHs/j1XpilV/Z6R
0Jyvp3CMkG8xwN37HGuZYIdtPpzBiVisKUn1NrHY+6TkCis1bnRwtij9TMSc4Hm2
QkwqmvO//qjmblwdwRhnELNGeDGCPnVr3NOQjtc1MDZxzr1vrnF4LVux3J8ycKGL
4CMMIXFxj3d5vN/ld3zgcQhxjh7gR64D61naRCFRjEdLzhPhv9Q7t4KWTMl7B3F6
tvykiF7fpAeSC/3S79My0h9vdOik1p1cgSxkfnt4dA72+qJUvx6l0YCGluXIYYjV
AnSuRq7NHfvnIv5lhj3V5OTEKtqD0CbEsofu++nw2EHsUxhc40OMwjrBK7ylEMtf
XDTU2FvkMyMQ+GvSaT1Kv+VZTY8xABNL+C2qpum1bGl6tC6VjIWKCCV/l1PNhKuu
lU4IfZDoqBmSYWgzEQDIA3HIns5khqKN47wDgkbNAzJThERcEbZc++tmxKfVieN+
q57ykaQJvZcn56mcJx8JjwxhFsmElu4R70c+8hoMV5V5orYiSXHQtLlip7BvQhoh
SRXkS4cwoHjKc5sZx+PDR/zNyLxOH0UPT3TB05UlKqc9zXRxep3uosksEjcwnPPY
hCn/QfCYbGCHMqN8X8/Ww75d8O6b9X6+4SdiyRCM+IPN1LX6RCkqt69SoUVuHXr4
p5HiiC6zzS0Qe6xFuldzrFAK4NyNwQLlrl/xe6E8fLX+wlkgXIiw11ZvSGR9i+fE
Yuikk7xKhtPXBEENj+gsZm+IzCivus/KRd/B8X9i1nT3Myp+XuELTnd/v6xjQ4gw
Mv19p2Nsbls1hcZx0G0iCGoQWyxHrGNtsaBmxemvx7W6Uf81ejAPvK+CLiWkqRR2
6iUm7FJgdXs3owD8zZ1NY3XE23CmQKT5Xor1vDi9H5Gm9C9qKpnCscdwUBbLQej8
LnTL1FSh5zNQyzbZ9aPt4PpcQ/EubFOvXQMoaghwR7akgmeZSsvZKzl3E27JcQ7+
uHkAn2sVqYUI/mY9GlaQHosOTeE39t+cvpJjgw8fxfKJy8bAt3+o2mFbXDLOgXju
4ndcDFtqsS4TTgHLKRV/HWJR2Sp2qIzOdMjDS4eEFSKPdHPuinPK7Y1BPFoqy8hD
evr64p0JpCS/v/7qz3No+YKQPGBsEpLX9DEyQGOwLCh3ABPkV+3u9ZBLDOe6xWI7
P8jm+0VyIWt5TZRe3GZntk8EBLl/hV1TKOMRbzR8lZc3X8zOLA7XOu7pnXdfDoZG
EhIfNskPQ242yTyH+bj5SGb2qddBReC26RKWct0dxhc9cATeEqxn2i9gmkQRePgJ
krQJjFAfNGCiyWU+gyAicWfRn6YIyHfxwCLoTL97uETZC4CNY+s/WT9BcyIIG4gb
bzfc7I5MSfrRDdr4NMU9KeiFyoeS4krFvIelCtz1HabGqxyHk2ga19JJmWHTRbmn
YvY1lusGFdyOVEwjGNacMpPKKNVe994MAl2kc+RWrxe39ZMoy25WNQJIN/CJkLmP
Gwpoo53SZ16jGu/uYokfyo3UTsgdIZLOiuWATVYffJhMfrTexewUDQ31N2VZaPxB
8p1d/cuJUyyK5WtFPDzf1EKHVgvnBWl/coRm9c8CrzwfjKPNdB4kCXzD+jx8DkiT
M503vabL9eyZC9jvRCDhdcS24oo0nYLzS0YLYCMnhpKSyZ9ZV9K+qP9suCCGEP3W
cC72WWPO5YOT/Hwf0qGZV6PfwFYOUe3k+SnACHQz8Ir3PdCjU4rJCRWn5Q1hocMK
UwWFG5saI2wZtUvXkRLK8ZgkGbupMzavs9xP/Z1xWrV5CM+zeAzIe/fHY3yq1YjH
dDIlt7skqjvS4HvQCBxKT1hYW0HA2p81/h8dxHq4i5hDaZKkE+b8LRCcVFq64ap3
MB3pRU04HPOaHk8wYfYhR4v9+1xSDPqtO0o2lj1ad4OOH3cwsqG+CIjv0Gegn71/
EdFHwcj+CDvQCORJJc9XOp0WhQ6dPsPgGPnNfcH7jU/g2AjmzAS3YLyJtd3iB0p8
k0dN2BqPXYaxQBf+k31PFBHUaIfFtRunp7jawWwvE8EM8MrkxrEQgqa+/5q4hRGs
WchcS1BP7iFS87Ppfj9BUe0KxPhNiQ8Fk4FJbC5DraIDLmv6U1wpBatyGpu0aTqH
Gjzo2pZYH3o4CFmK01qxB81jMEEjjyw8BkqZ36YwUmoFnEjdqqdLTo8s7Szrg9oo
LLQqChs8tT50ucvZXp4MgsJKfkZNFLexAZO7MMZRdjljY4eT4AX6Q5fISG3AdLT0
tQx7kBczqnoWP1mnheFQ4yamf2aqcjFkUtbSCXLpQvpQIB6iGLqLp4HqFyJUjfT4
dCVvFThlpsp+kNnSk5HQvwZyEfsBqWwRHWGSjpnhcSPF88LQUchwy1ROZS5vx0KR
cCvHRtD7jFfcgIRubgvgj3RnDbL/GwMPOrRhhAOWOt2McsXz7nr55xE7GCrGFozV
BF7AP1+QQWYz2MS/RM7cGaYFcUPRD2O/PG5MJnQkO2caRiJg+Bx41LtRhbKBCidN
jUl/y3Sbjtih2YGzRiEnwc4u8mcNFWN1SYPJBqqxAjRReIzA+NeI3PWf9qId0x43
ieiGTX9CBU70mxi7viTOmuv8xfncEi1ughSflFySFFPVhB5tQSvv4Ua2lELgWSY8
I2b+kF/svAryGuLyl1ow7aTbWDYGKbk3hsGgsRID/dWK44Qvyz0CGgaHOx5Mq+oH
7H/tBGA/9P6vC48xszr64UAXZc0tBH1zj6W2RY83t0B8hQfzO/Jx4zN7D65bEuyM
15gMKSET8l5FS/+0JSmw+2Mf2z7Cv/ObUrRbdOpstP6qg/bH8IvI6/2fGC4o4F0U
W3mSLiIphuP8GCxMNjg3BFmS13lXyJ9jrIoGEQEj1NoKr0O9womh/tvHBzMNutqM
AmI1pbwvGAKNdy1RPA3czXKS5Fwi+lT8S9ul1kO5b2Vw2OW5yR60CCNETlS/I6Lg
ym7hwsWBe9R0TlgrdJNbvPAqBwfVmQdz+WlZAY8BBQRbtRokoZCbL5ScauCMVmf3
HBtjnWd+wiaznFefCnHZIDM49r6WjR9pMzie1V/azEYSWNMkS2H3Dv5JOSo2B3hp
XPDY5LGcd+IhA4uyrvADD7ZVRpfcl6rHSA/ZBDXbH92MCAfCqIHUXLV0UNOHVswz
p8Z1fZp4wcYM5e5qGk1DtT8BZJiU9lARJ920YjLd7fKO2kI11ZDM2pDeBJ2Skyjq
UR/dZ+dbB0WIx6RtvUBl7aO8f6JrFNvIOHqPc/Vz4BtM98P6O6xjg0IlgTIp0tts
TyVEdysqM6CyG4uz69Q31ii763fiu7uA9NhDaZzGRBfr+FZ785r++3DbX9wQl9XB
LCHef4Qr3cr7vMaCyEDqLsr+LF4rvs9GrAceyzAhrpV2i2V1fieJVlgBIVAVkXFX
V1QT3E1dP4q9+GNeUYzaZkC7diyrJi/Ru9FJBSYljz36oqzCfnKxwQ+y12FaaFs8
Sohl6Qbe+jGkCXJK+cRuWYwdHNBiwRAXDopn9jl5TSPQxR7p+gtm90olWM2l4cVk
Du/22ABExMtKbY+lYh0V2ZCKhdiRu4eq+lxbsFpWkcenmebzR7e+dQ93pxt30s2Q
wdbPYSMZGnC9SF3+mkqe67WahyLk1l0mtYdfh3NbonThomFjQhgHUOnQ+DbXL1YV
BrxO0cqRpDuudUr1d6jBGdmOC9kDhfKYPHTzGIAIrYHf1+trDydJRQ8J4/WJoaDa
+nGNeAMlTcDSFpsDJ6etbaiUfiZc8Y5jPBuJKkbbpcR1SvQeF89rekpiGO2AObSH
/OsrxlyGE1aXTLPzDhHtVtMBuXbEoDI+PZ93Z1zeD/iFfr5Xv6Etd4IsAeryUK7z
fcpuZZXfCBjHln+eyRh700G058puQBXKI9zDixmrw9i5A7YUeoBeApEGAjLYnE10
gVUGqsA+wvqgIUSJIi/Kga2eipjM0OGZANquVfZ3w8tj/T7ExdZgYHnDw7mTJRGw
AgcSHRkYDlMKSOHEDSkBH8smFiE0hlTUDrvVMg9Li3HBBo8AuhzGWHIaQZQOi8Pj
MsAogG2/EJvCusn3+0JBrSjPnx3RFgaiU7BmCa0uowCoJHKEPCaYIiY5kHUtz2Rq
AmS8Fhwq5HxUrvwjbVse65REtxLImEwLk+xYcSP8oo+Lt+I2pf81Gze9obo+Uzhz
7m9JOo6vsiBtoZVCnFrqcamZMsAT+wfVHd8G9t5vWuLmwpup4Ptz8UbPU/uILikT
XVxnItk/mEBqUQLWGIbnxD5eFoDZCll918sMAVmmyLMK7RxRh0eJ2W3g3rl5IZuu
gM93wGs+63OciUkFKZKYWzuKOl7OLGcqLjypQk4PIh3BRm7UUdKRjO/A1TU9swAl
evpLTXO1xrX9GVHsmmu3E4o2SqTKckHgrGDE1VGoZyhsgUGBIgN/TQIIJJ65HGQX
aWnseFVmChOPK6A+/OuM/gs6uXjfzKa+kBfAgrkKAld9b1kLZbPlbyWg7DN0JIVW
BNvYQ2/6MzZVZzyg89V7Sh38f3wZN5H4bbu5TNgyJ5kgniukrUOhB7PwnwNqCkuT
mCyRy1gei/jAnRSvViS+XCcMG9WgcB63pqdQmokI++ermUd3F1iTi5Vweg0JtpPF
ggak2lmTgBNJppfk6YVPjzA0egdv2i69s7Ws8tSUoNwR5p3G7VN+6dJaeL3uZc+H
NJUpLhlC9kKEhBRzQh8PpJLuSzeInnuIaVwtGOIP0L5Wv5VVi5olBB3lbF1hWnMK
uSPQ3NBm0k5GdaXKcgxKrhGWwT56a2gLtSGF8KJd9C8GyqfB/ES5TdKOeaedvsBx
29c1pYkp9fYZYcsl/8Zsom43W9qz3uJu3QjMEt9EfjawLyX5Uf0A6T9cURFZkkg8
a3Dw+r4ST8RIwh0r2h7AGQDArlcGWNX3o3tKDTyaDK8=
`protect END_PROTECTED
