`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
icIkGuoD9vXUgEcx1viUtKMLCCqB5rshaYJxo9ZPIRCy7sJBB2HuEndJklXel4q1
qWesEx9p8h6wFnQhYCT/3q8eAzxXW4E7sZ7w/ifzdFiFYyFT96gu5S8eY66XKFRE
ZbN7UtuP+RjsLy2wiz5YCTt4kzjZV76IWZqZ7w4yvoAZCj1fBB+aa3cGhEH/NJZe
8S4BrqA0lI2maAvGTR0UdqU92lqDKM+NM3N7WrzaMLKN0uTioGEzsgHbIzIFalb0
xfbRF9SCUoTnTwzG8x5NJcR6A550InO6B69sS2ZoFdBw0gH98bvkvCBi6MGZkoIj
8MhDOwpu4Naoxh+AkM7G0kMV9Qoicdcj8jd7libQUQ7PTl6vFVa8tyoPtax1LDoX
4E7qFKECr42h8N1KvGXQdDvtVxLjU+NClt5wWFe0CD8PEVJTX7qGFeGKWqjdHvSP
DY/s/BUFlbcy0Kx6sXSJkq9BLuUikyYt0jvCR6qZckz8F+o79cG98Z5uREgYylE4
mjSF+ty9CrWtpg0JSb85yyrUcH1go3BToJhaVJqqUZwSp3MF8PNkBOZ7bgdAzdoM
wI4ssgv4v1mMDCqx5hhLDDTZMMYwiPJPV0N9OcEruv0mhR+PCNodfNXT0M0CCqBc
qt2V0i/QoX2E0CI3byYl5sx2iVwvYOki0t75+srW8EJhK/SGjjG9kn5OQCNbQc3V
qWR70gmtNgxMyr9gNEFrdy8M35JOCLaYOsOP4XXP6mzgJugzRdJ72+MTMI+A47JA
FRenvjnNwFOMTy8xlc8wpPMU/4cKnja66FcgRjf8Dn9dk83jOrGUoDIV6c6KWn/N
kk/pvAYgBec+5G5z/26Xx8lLm1+uAOPIKTFvlBWp92r4Kf+5Cu/cS4Y9VOAtpxl0
BN2Xwt+ITnDOGyRVGfkp/EDS9OIXB6zQlpQfbL2frb5NHHhQKPHLvxBWlwKYXn+M
fr1AXgbOqDtjk8LVWswt7uQXYxcT2Jvb4Mk1vnm7jx1Js0OFgyn6B1aboF+RD8Fj
7GvfBt8oDJ+Wbel/JSnqFSci7zDXFBhSkMnEOphFLK9vislqF1VrH4EPY+F2S3hH
sQZ5qG8clRjtDu+ig/XVxpsxTXxYE+KxPHUYJk5iyYyL6zU1EfeTMUi/9DXHLzVL
gUNwJs8qHqIxoA9tdCxkhuBaKghL6vhFxxk4suEkc/leU0F6DGnvOVUiyakkzobU
HFGJeGY8g3qkOmaOiZ4i6F9miPGdxz96EAzXhRHtZm6FqaWRxCNt+EQIaY25d9Zn
CXrG6mCgenna9ePLAxv4ebcHXr/qafgSRKRHfw65xVVk1OEfWxckuDSZg70bUCpG
lBXV6fbbwrLcJF4R2iphK1mwT9C6w4Ucnojl/HATei9zhJitHjWBiwYr8SwPIWQj
cpK7uYGUWsNGHpzaP+K/zpJBepO8jPd0E81sdueToR3gZJ8n8BaUn2jsEfNJzlMf
zhs/5jbCHWvsJjvNrpGQEcbJLQiuBbK22s7Ycu0foPJv+nCqzylIx2b9AM1Ks6hf
VavzekyaHNowfvBKgy7Hs6lrTHRTYMgFXmVUa/0BqFSfcCMh2i+LiO/G8GgKSQ20
qwZW7r7Uhndlaz7nJ0iJbas7u19TqZ32NEE3N4OS/zMbbHjXeuvped9C63qNiW3T
4dbGRk2W9jBk5yTnVkw96E02tgwNMJF5GXAcNaChTdL5RiVYwdpNRr8gYj7RxGX0
AzxKJuhSDUOqPhqmRKr6WNhyQtWDz7oEuBQ4PnxPlKeRup9Bn8/yJOIkvbDRYiJY
2VagbQimIpFad08NO0YkMbQkja60qp08ln80HmjjYmcG/5UbIdn9zSrsaNHtUiai
jyQEXCLkfa7+YzdonE8eXo67pXyRlRdyIEZDT+i9Oh828bSdmkgYWz/jRHNCrBof
b2cxlfC73hNb2djEQhwyy62BgfEu7Zi3clW7AkvNgR8vJC6isvgH/+jH76uLXTuN
thF0oqz1cKWw+g1IXCrAPXeXR2oKXJ2/p83MFeGH2atB5a9TU5ZPGnvcoPNpNb3F
BwUFyMDQZWoQisZmOsJqY67IJD7KQvEn4abdR6113l/g040m2F4UDDLqf9JctWIo
IKu/yKHLvo4EEGOJYgPYGck8L6mjY4ktTqSSw1T7QlW+gTzL8NbBLwogY+34NEkO
TN7qcJIh/zzOUBx2x4Bn+Cw7oGroomqKCFkToUMEQ4oCK12SH551bT2eSXJeZ9vH
2PpUJA5/H8Bp6OSNxQ6CvDMUCO2GblP//sjjzJJrRXOFUJ7TOJlvjE0vXJVTTrPE
L2uLqroWllN/FavDV0KACvmV31IYsWx/eYMswDSZ4OKvYh8SDt3xPtII0eQ8SKWx
zc5jgWItVN08WRc+SKu5rUyrMsQwq+mQocKfn+nT5r3Z/llfI+chefSEPxKzFSp7
lcqUymiXo2D03x73YZpeSS6+YFMJOtiHw+jZ7DJxO2/Nrispoe9rOOWegQ+/tLQA
grajOn9xQovUxQ1gVjTV2Q==
`protect END_PROTECTED
