`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCtMp9SQbPrfimhM7FfuBC34BPJGkFjelhR9KskRQpE3YTLl9Bm7o4SGv3/naju6
r46to9z3Px+GUUmHI/oqWv9CWKJTbTT1JbGkipgRmLk8gYWuO3DRYG32qLLwfTa8
uDJ7RiP1A0NK10edidggwD4GL6g0HevZWu7NE9vG1q69fGmD94D85HFxvmVPJlTD
PBplRZ43h2HW0DY2p7CxnuZZc48Xfkhg+XqULLvICW1PaFq9jvPceLcqCjdaLrpq
Qf7zCardAtGuKnLbMBZigpoGYJAfzp5updluw8EkzjVYc3EPQy5cagXFEMQ9KyJc
DheFuWqTSlkjzmKa0zUoxtxvIym4Y+g81lsIQAbCeTtfDJWQMNH3eG+7+jl59GMX
WJytPVOjvGsKIKuht4IzFUq6Jc60eX8y/Yu3Jn0gQSDOYJsL/rGdpGmtKy/SLevt
EKrPabz3am4CUfGiJMbdOfeCInvY4AXklftZRQB+xtLP3dWVmoWGbiVsJ0/1hlCK
A+s9epb6aCqGdOGuG+7h8m/PL8rGazb2mDm52TTt1Ed2nfKwsDr8IbakQzHLBzDa
p9E07+zfHFHlYiYZR7dyUFQPp/oFwjkpBOIdVsAZ5wFUCnErmrMLEpg07Ozh/hVP
z8zC0ofjx96OYHuHKW1eW6na9+tscCguhBkqs+iGW1gGiEH8pGwT1HS9XruNh2MG
/rVFJFWACzQ8a4yAkR8jAPYjSDpmUVaW5o2YT7THNiVlwq5irqW+FSHR567PTMUl
FjC5Nn8rZAa5t83vySOvPfs6QQcEKnF5oChfDiNWlWpQQ5wq0el21pifeChOq7nr
RGCMuvDo41k6mMX0dqkugsUQvxNJxoD4iPyMHBZrTC+g5Z57WxZ86kB71BxhECV/
m4Wg5miEfugrDndwOLo3jJCo++UwDr10sLOF3v/9/HQgE9fbGVjqLJ07Y313Zie8
Hk/GodeI+Hrf5fVRJyf4IviCptTVEkN6a22ea+AKYkNHKTCLoDoocjUZsSPXYHU3
TOvvtApUxMdueH/4QLRN0upcydsroZGXUkxJYNdscIIJOXMFMch5IV1yM+wX1a3u
lBwIdonAFxmyfdK/MNPBQ6J1/qwuh5LgU9OOy+u0q5Gf23QJWi/Us1LzOdQodl7j
XmL+AKLGxkRZERMguRw/dFDaDd7VnZLTTs7QmMKwig2ux32zOC5skVs03+HNxEz7
x3gNEBZOxKWKF5M/rd+e319zlfd2JVsXjT1eSUMeowCbP5jpD/08S0OLa2QbxsTV
NUJ/VXqn9rxREHiHVpxbqiYnBIPAUflnFiHwOwPy6GD/qD66e0TAkGT/w5vqwWx3
NfDC/QdYYchP12rBb1BDalI15FKzW2CGRXjwk/2Akf3GIT3YPMoaNVOGACJlk6Wr
k+S7HhQEvcjNAZxOerDre8ePOuTg+vxMZJROFQAgv78=
`protect END_PROTECTED
