`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AtT2gRXzGwNfv17AHfVdv7oQ4R5e4XYKY+zA9m+afUZigW1j52GP/tehMyFEg0/Z
bVyfSjwVC2hF1kSJZszJr16SMJdGJWkLCfRqc4sp/hLoh1r59Wh1C5THblKCux3d
JrR+A3ZPAX/IqtdAfLQHlBSNBZSlxTzvrw5uQZ3wmFEIe6+g1esavZru1Yu+x6hc
UcEew83sBqRrYOPDefNVPCwB4teRbsc+bZl4MP6w7cJ3ldqufs2FRmGx7cqDfbfK
BlNN0EYxSPRdD5q/KaPEZYd460HdEhkxcbXE0gt1us7F6Jld/+0rMcCwybwCCyKH
IRHS0k2E/6mScJIM/LsYtbziq8o+7rgprpD+MHivaPY/1qYQf+rurvyGhf+ul1lA
/GF2aP5ARSxUYk6oEvFFgW9ZQf8piIgS61EoB7/sfctvdcNYfkoJD+9utml+5lsS
dvFykKo0/X9Rr3JYhu74G66LA2CkfZnD9LrGMJfp651Sa8yQrq0jdBbNRAuINmB4
jLddsbwaB61+RbwsWVL9jzFZ5OLiAMVY+4lX4Iv1PTmxqAe3YlkkF2HaIyhRAi4t
ObnVQK5e4y5PVnbhLa2yjkvckyu6VPfWOK4JNgtVVQdaTl/9UsqJpXATGnNHTVE1
+zkHhUZkSA8jbmg+hQhpgG60R442b4GPwzjk4LuZ0oF/Hsrik4mB4JreYoqwdwlc
71ViIDjbG4udrcuj1c1mT1cCC/lsqsGiv2LPNtb9FTStTuZZEwURYpZO+LnfjMNv
qgU5c/XYQXgF2b6+HIBsRQHcynGeAcK2KVnxShvOY1aRpfEt9hHnkkECCNwTHLn3
1Fet5Cn8QZzjGnaI62VUgak5PsIOB+d9AtcWQh+1aNQ=
`protect END_PROTECTED
