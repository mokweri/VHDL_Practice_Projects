`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qn9L6TORFqVUkDJ1xvelLvBDVEJddVzqyDNO1/ZupQh+Vwg0J2XR6T4hkhGo70ba
33poN3NZv4TpesShTq+oqXt/JHebhCXWhUmdDR1dCBEoodLpuqkeOhgmcD7HoGqo
MAh25R4VQ6YrjvgyQxGvbRrUHwVzU+0bGOHipkFNfAb2mAJmuJEn7e5pvVeE4bft
ojhE0sWqQ4pEmweNoX6J0E8epXNjWEWwStHzlJ65vPTNz7jLTh22+BcPUABTRUiH
E4SMHxJQzc1/2/ifz0DBrFK2XsmeZHavyihWbsrcuDByYTKOhKzErVnMxhsU+qDq
0pkt0fpzwnjAXEWoCPTCv0UJkwOp1P6SZaJBslh5ccI7raX4JPXRVdYB9pyUWp2l
7PHs3mnxzY+1CVf0VEBk8efWMAwWt0eMMFvC92k7LTixF2plHvVlWg1MngqmQ1JN
GTopV6L8cseTNHZ3v+U6i3vHFdrQRgpn7ls6KvKmu1iuLgCpqFTMI19Ne8OhUueV
djSebwsWy2FGlqPnW8UcDQjG0hYZEQg2fs9UtD6UtZmqNjMgi7hR8mLXf8n++BLP
H1iEhihUdwFSoEWQrbg+jzRP2CVF2F8Ws/ykHBl2rza5d40oTT+EdRttN4B6DFxb
syWL7Q7h17C6TVn8rEcilz7xfOYEqy+h9WcRX/qC3LJwBQwIlsxJNcp7OoRUGM4e
YlBKkL7azxO5vCUbF2dijitR0ia01bq50n9UATso4GJLEE5vPV5htX5zf8g+RXsy
qnQ5jqaSEmlSVuYxq4ITRXnvt99WhzYnH9v92I4Ga1mPdK/y004jP/BgiY1BqYYV
wGbynBQq7UL8YzOap+n4rtvb6fvDdyy0j5UNmrD1TeRqeVQCnug4CRLhpDiLG0Js
4hCQvZCBU0XUSB34Gyiu5S/QQdly37+LWreAQdT4wcNrLBkp/b+Bb7Q5NNoR5ZKD
nwgoF+P989Xpibw3rd0G5mVNsSOFlGoHqzu1zt3UP/zHfDklzZdtYlNTkSLIDCIP
xpKnvEtWG5mFyeTnoqPY5kLCn4AfpbanQNxkZdrJogYThSFLyfqkWsRRGV4xYZ+a
eXwQvtGUquFrnuQxb749PRJyOXdm1DtHfcUhnWD0KKK7zwWRIbqMps3JylQq5Pkc
jWNAAqWxGBDaRXvtHtDDff+kQpiGWHMNVnagWK/dgSCA6gEO118ts7gquOQ9E0Mm
XxV4KCOnQuKhMFz1gxrMPWp5YG97W1Ff6BViU5E+59wr0kK0ZiTGACdUabvbAcgh
2E4rVG/KBB93W0+OCNatrNSI5FANxqFD8siiMgxUyK5hM6z3tru90AuQY9fHYQlz
cG/fgHGdo6TemqZ0BC/U6xIeQCW9wDmGGuBgGjCzPZ/6km+bctS6Z68kB27pH8tV
GuMvZxg580gX6DXC9Z6o2jSERkHlWJYQpiebbXI0m0A/id3WGSpMFxkOu84AoBdu
cVBmYT3dJngZt5i/kJDEocnY7uKopBhTRggTaL41SFnKWdyMLMtcCxn8qRqOlVLb
onS53RfrFbdLqV3K4GGQfl/QY6K3pJq/HQUJN5YB2NIR9BKseNeGMcJHq2tATCyF
4Q48aM595pPl6AcXkihaINd9qh3fgHMOZTJiIa7V05V6ZR+vIOnsU08xNsGyhKSJ
SsJZEabMmAU/m1D4EKlj/ZXIP+vBN3m3HbKDpnzSGjjRRvTKVI3TyH8GoEiSDwZC
8D1BqkNNzPkuqIZVoPr5+53tdriylBjZXr14AK5uT6YIZPo1DBnDVNPXZbVf1wFg
JWz2VNxb8iz2hh72Ty7+2+5tvA7ouhIce34bZF4liBFSK6GRFRmUU2ZeGb4QRqd8
A//EgC9ep9EliwnLzu3TvPE796Tno8Z2CjmKxeilVP7Pnx+WyNXp233Apx11ET78
TfjjIdfgvUMxUMzGXv2IJ6fGPfdq+GKgAcRSXO/M+Daoi6NFbxJZ1LG/uqJeo9WG
`protect END_PROTECTED
