`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TowLSWL0of8X78WXTnf366pV2lhjEiMVEtqJLGD83mgR9zdioxRvth4KrLIH8e8q
1wcweGxY74ltXulNiuaJCe2Wb9bznnZuDjN6jKvHmlJ6NTIREJ/C7lE9japmH3S+
apvVC82H3BJy03vMjrgihu73hbwmjzUdZJsjXX2b1xCMJybGSCogQmiqmx+xdC9q
+n8aFYZzx9hd98iRJGZVflCDOEjUekdXrTyN+hlrkYtCeZld6W03J6dV76HNYKDY
o7Dlq5TqLAIuh5D/n7RyWKqpOrHzDOYyY6Va6YdUgr+G+cFsk0FSk5qtOZIvr2UO
nIef3rvGxnHeDlewG+ANVQsu5N3H5OsTRFtlWW9e3V31PqNPmIN+1Mhf97Cy9yqT
086vUnc/OllLCka/7fob13NoyEnUcmh+HJBUtsBGiMOez4CEdNfHIQXQA4my8fcn
XlXt+J9e//LJUqGMGORuaub36KAba3mJc8YJs8yKVUuspkw4bSC6K0Zkoe4fwe93
OD6TazACffUeZxxiAYXToh0AGJL78JLSDaauluR47sOIKniYwIKZDaHYLCt45/8n
IA0KzH3gd8v9SEIqiqhZhj3epWjS6tdifLtDNxYD2UZRpoHUsSYNX4TKL+mPWzlj
2rmnFLzu16ItxtmXwrgdqAtz3ztzfZaWFxqi3mlHpaFFcN6Dfv7q2CCZUip7kBYF
41Vm3LV3SZPWqF6kYXgndaFXOudSEj/TDUvN4VKB0Jr7Lw731juFzc1Ngfjj+jPw
3W833aQFVUBK/Px4uLBQorjavcpgTZkwKsaURGBDiSOYIbxQCwNHXGfgMnIxm8gj
x/M8sM2YswE/DJCQm4xNzkqiwYfiV1eAqLEWG/INy5Nlz9KW6euwHzA+0U0SaIJc
Fc9ziUT1g6tLzj3DMmuzCWiQtrZf820M0Xzr030uDKy2L978GKxd6MQ+NjQdT05b
+9uvvSpfJfSe3x8We7kmdfgjdmjpUtzEiIBSivVXVpTIUb+bjRdFulHEtUdorEGz
YMvvN3e4tMZk3yIBj+J25QtyUzjFYuQSr+KSsSE/p8c8DO0YLr6x22b6WkNpF5W+
WgD+fUiXVQZCuT/oBZMHl0prW/SxhAVRgLepeen/2d9hQsI3B9uIAgORaydLjdAt
qjE4rhSkWrBjZ4RlMBAE1buXzgNaKYNIlEtaJU6mn/j9qujD+isLUzzjGtto6pik
nUc/aU9+b8Q8Pw8c9dFp1ZAaJ9zqBDw/WBQtoL5pa4ok+h9tJ61bbAhZrDPRdZVM
eXX9mEaIHuCqZY6rNm6U3KO3O/IYJI7g1i+3ZohpC/2JI4quWNE4jVxgDKyouo+9
JOKs954N3VPfNttAYW1+lsLo0bWwAp1jRKgOB6Ii3zG8/KPEvT99sBPEq3ootNvv
0h5G5SJRn49NmQDpZq9aLhWoauzwH4wSLkKnu+fiddOoFbU0Dsuo6kWD3g+jGy5n
IMDnvOEsDJQaTIcyZB9Z4nXnMO2k0k7yjk/Wnr03Nn0Qy8AzhM29QTytqeNLaEha
lF7wq/lCMtE6FHk2Y37McbrTtRcdcCJd3LvBYNUbv7fjD0TIvNZK3WpE+lY+lUBG
EIkbUJZVdEhG19PtAIEaKz+IPs817NPtDkDS2xseJmSK9wjTDhUpphptGLWaSDJg
8Un2wp4oJqeznAohpSmaFLbDe6RKkASL/BFL0V0KNQFwIEd8SjajFRfPTIocPUjN
7zSXg2pCKN9bFgLUWzjh3b5atgGrLlunqIWsEu/x36OK2lnihVO9V3O4npVHPm1t
9oIwLjLIY/lZS6pa9JtqSj2RAg6fIxL9ZMm+TptakglsK2RHmc5gezUPqKRj50we
cxu9WJW7FFkiI5dr6nDtRvxQpASQIaptDcCjF7OhmM0wamv/UeWrTtEMY/RZRZH0
Eug/j7SJFAzW1UboR5mdjPt0DFiNmzIpDqFuSnGJXcXt1bW59XMwenNbZ7yFlzNa
lslebZi1M9/CsI4wve9V1mEVP5XwyiPteRP+MfPGVFQze5qDHs2EhNmyXIH1MFGg
qRxWQZeOxhWTBJInU++WLuHfdadJsdqOUBj9CCcXKpX5LyKmc9nvqGHDNm03KS6x
+erzuMcX7YLC+/buQdI8Ru11OrCZFZiRLOo4VC2qa/4PFgxPNsJcCVa8c618a73W
T+yeZaaWRzzHUVelmtvMZMNY9CnRtLfhT6GecN22yGlmuwWFAe19+uP4cXTThK/6
4Up1D3iTBLrhkLHkc44N9ZzG7A0guWofJzUv59DfTAT2neDGujKGoKoyMuShuh3i
Qi4zmiNe8MMRHcC9azkr3rU3JkP8ah+zQjLxigKtTeZ7F6TGRXAKtc1DiZMQ3sHK
FvmGpRfQZTdw7AtsocI5qzVHIbIhb6oQKJyesHNjnHr6AFS5GKHnXe/4HmVa2Gz4
kQKY+8DKJTqrlKSMCqUcGLSnTNv5wOw5Ert4njgqbZO83cSwnljUC9+JW+W1rqM0
R2In9oCXpOS8nHtkN8Ifv7hfIYIP/xDJl4fkld8v/s8EK5FOICdFIUs+ZX82AB8a
cLFqglqHLaCulPu8i8MFvzv4c/zSgT9mfCBPsV/nrIZkz5jRXsEFyNK24v1DIBKK
MQAJEuLKKlNa3Is+BvT5QaHdsdvdtaoGZtTQXt9L2sjy/9xZTMaJPi5DGvC7w9P3
Ve4Tpfl3e4P2lBhyHMYairAHXis2EsSxNIPYVHZ7b8lhXBI/TatOZGeAnucig306
`protect END_PROTECTED
