`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o34p3bmLUb6iT0jhsbpti7+EZQxWF07uocEQnFbcfV8q58ED4zmlO3aOAHVlINmI
NzMR9gwIsQphqeffLovoM+Rf9RBmIjHwFpmHrq3ldCpn9HJY+CD/vF+rKAmMuEn1
5peS2SX1ZCS8mf8WETwRJy7X4fyVFujQ6Tsy6XqwB/Q4rmJa8+XjsIskEAyZ2Pm6
YW2yAMTA+xtVsEd/pf88/qq+KJujMw9KqHn3+6OBHNTo6cN3Yvo4Tsl0hEgwOvHC
ybdGIiGDJ/MRfgjp2ISHYycHjmJNG9qDcRe/GrXhcz6jDFpA7ywFOfnwK1Zys1by
8TRk2+Rf1vZwS60g8a5sZp51C18c6gFxg+5Ad2/DCvKmPZ7RboauBOr9es/Idlc+
bC1ZfUYW/lyEcFQg1LNkvoihEvL5FN+flZ3TffpY4BAMj5d4B+oWo4Ui6/MZCl+F
L7CPXpDmkOy6yM8sdDxW4+0I0uJgFkYD4vvFBvew179PhtVRsEtmsDRPygU9J9Q/
9EC9wB/j4ZVAObY/m6BmuLiWhf0aBNcNe95VJC+20NANsTCiZLOkYn1uBEtnr32M
9b7OGtU+UGtzFR6H3rRP8vJZTyrgAvBFDvu6thr+Mxs/aeHOq/WCblngwp7kBDab
xrfVeNu0NwMnwNA9/cxtBFnJxiCk8y3ylzQ+CgenrKrmNmYcKo9HyQ0yvtBY/Rw2
63LsKtOLapslmIb0AksoF1GetNAiNBTkvsSJJzjuf0H/E3TwysVPxkH/I9X3sW1F
vt1MVZV8cuzfQJOjeCZPF3NgAwOs5I0y4dPxud5WiQm3vwsle+EuJ1NQr8KZ/+ar
yPkkEBtQ7vZ5s+GEEVbRrZX/w0hcnltRPn4Jfxd25obEZURdKYueECWPutokG7fN
v+/L/fsKzkMlNNwmMh/VftMT07BOEb77+tayetgfTFoQKsrMOEU3yIPeXhAfcNBy
ktyI9SWTeUN3yqPd3hg1nW0keV3aLKazug1HvOEDr1VvyyrTRh+UQn/fp/CKlgXh
XIo25pW0q4JmZ5mXLscDo4MpZY+7xSOH94uetFgU46c6fvrsJlbYv+CsduSfpKCl
7tnPo8xis1+bRJzYSYtBZ1w6JUm+9F8qTHQOiCzyhzCLiJbx7iq2g4CT6ElQdBrJ
BRlolfwu5YybIp26GjWIAoh9qUrDvJIw32g7+mrg4VQjMko2Xo89nttYmHynnQai
lEKVBznlyMluwYUlRd6SB7XbtMwQtvIhizkGKFGuTdgq+RAuvW6OR+z9B3wtD6me
Xs3llK20wjlXJkx2sAGPLV5gG58dtDcQcnZW8Rd8+keIQjzbSQWrUg/MmWXq7cr6
nk3h/fGS8wnRtXWTNEDWywN6r8u655iCqUAzLbhEpkHa90kcU+EvRm6/v40auQ3l
bwBSYiXBA7tSgJVcdFhSXRQfMn2LL5V9OtbX8AY34UMUBkeD55O+nWzoO9HixNSb
ASAOs+dNPOv2+/n7DAWdwgMEuMiQenDn941/ud8N6jRz8K3mOLj3G/YWGQnvKAXp
VAQTrkx0Iw0jzO4kFPlIkpfYIvVTFvRzp8p+iF8sMXIDzw9TcyZqSrNFvr0Ms1MS
Jp8JEZB1ggQ1TXf5Vkdo34ssRz21iD0s8Gx1WkPxym3HVqgpcN3AhgzClG/BTBCt
pb3kHKUbLCzGvf/s0ep9eTC7MKssyx4f0IAUdv4M+u9OLClFx2ro4lXHvtGr8+JG
IU1fz7hiPHQOMYe2sOyUQF2I8jp5Ue1tze3kI5Wvk8R1t8WceQek/mD6QT2bIdOO
yhEENzADSbySjVu5jMw8H3NfVfokthLcJWT3WXRYVOhj/9P0U3iL9ILbsSQ53RV+
FiOmV/mKgEo2qH1v/XG47g==
`protect END_PROTECTED
