`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/BXQdtf3RkIxyiLgOPBj1quc8LJrb5qLyo4Ui19bMwb2PNxRfL23KCsJtkztXv8
+zj90Omu9TO8e6xW6MQjMViCpmp55yiEnUtUOujQnwwkXUAvr4L6s+CwMM6EKsTQ
d6DfICExF+CwbTgOFTLuyIABdsDYaJh5GDKPyakk9vL5lbCJw8WXBFjG2+r5IpqR
zTXmcOMGk5/QIloL20qI7AQCxQUk4H7/3j9h2Tiv50Ry96VOAmAJ0D1g5N58OkUp
NrhxxLzhMnz9cEkD2cnEb2rXqTcjqSo6ME+q5PCGbOM5HuXcF1b7c6t0dfCO8qJr
VmLmYPQ6PBpWuiHsx+10hry81e/SaV8V9leHf0PL2mSnVi92WFqNC3GQ+vVNc5wj
6Mvk9aeKTxAP5SxpvoXOcjawE9ZgqyopIgpcAUAnuh9DlXs1JX728iJ8sBFV3RUr
VWX/Z2kyuWLt0SF2al2JHB9eJOY5CN8atoFz4OhfxC50oZp796Ghoyt53cEkdYwC
iYT/DXBdtN6eC1ogLOsZRltLCyv/tBvD9M573VlGlq2Lm+jBM8SA0sXV5ZXytOGt
5LVUi3d91PYkeeFhL9n77OdDnDkqOvDeJHcNSVsBhdwZB+4BjMhfUOaS9kXx6NBd
WGALavvEZDkHIIOcFS+r4lupZYJ3eIXnAr+ulpPfWxTj3Ij6Jo7Jn27XaNsGC30N
dyXY4dmdWkQcSeLpnceSaedGJau1EXpMfB/627n1jHwWaQQvnckcMzkWCOOQhXSR
Sho3vBEYoNjpJPwoVOkQ0RVEpn6gkjFxuoLQWdNnRn0E4G1OluYmohaAZrtya1Sn
`protect END_PROTECTED
