`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mOCxuvbj+Wk3m2uGQgEjPDV9wr1tbBIWH6IbKBrpFV3DDhgnesR0IKUQzHr9ePhb
gDCHiqx4bEBd0pZ8gEH9lCqrfrmJmGumK4h/wdRoKm8ZE5cUVkobeAMCRDoozGq5
g9EVVbcKHfH/PUsY8RhgeV1aJDfxCJwcPCK7hOjTZwNNZ4PuV+c66Dtq8893eMls
lOI2AMsYANJReUuQZIWYkP3bUlppTTGIZ1w68UZTV/dFTWa77BXWNgJVyh6BWC+F
fZgCNiX0SxkRuajETYB/zvgC7eUgu36IDVeNu85ddYh1zEsKekFx43j+wu854iiV
lrQGsNB7o/OjNRSbjvp6E4FyAsfwciWS1HSbQmqbHhH5cAz0LIvFCYd+yCxMJdrw
0nXN/uiPZFJBcTJNcLT0/01TwohW+05WbbxHKORInvvce3FvF9ARoNGlRetgTJ8q
S0z45iTJOEvRGcHg/7YYhfQ4qpOdlVFCS6LrkF8w4GCb2qksYyjqRCXTaAVZ7Q0Y
lfNteN8HpRaYIE+vbIWvV7wlVG6ALg0gwQzYy808YHOU8rAVgeEbMzewbXgN1jmW
Rtrg1NjMV5QZXfgIHrMje/H9ovO2mTIwd72kVzMvqI0b5py/8F3ZkAEcJy3xIibl
nvfnwV0J4j+fI9wH8o/o6V/y2SZofHmFwsi7MrA29r1wIfjxetOXgRiqee6Zsdfl
+l1Jia2O3OaFDUERRglsVRro8cl1ye/iMKLO7G4qwg4SPte5c1zMk4gxiyrtGXHp
DMAluTU/9uwv3ENmBcZTUOe7Lr4EDyFXXpJ2wOFf3YU=
`protect END_PROTECTED
