`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RPrEyL05qq3Qsyh9EIyk2aMcCyMpFMFEeoC8ITJBCb3Md3wV5OY0+e88x//5mDn
3Uj19eGat9E5ICc9IJqyO4dMVOLdsdpEK1KEZGy9IUX2Xk0eP80q2XR9LMelMZD2
1iL+PRVME2qtp8n76sles/qlmDlWGeZFK653YfQ90fuP+nackB9OVc4An6zEW3Av
tlNnrRYq4v6XuSb5ux9j0RMHFL+r6E9gUx1hHADTUqFy90HTXQ/wWMAvmtCgHIo9
nAFoZPhpcG6TW1+mzsKfvksB8b/N9YZEGAiJgOlMTS+4Y1m4C/jgkEt1T03rtMoU
+B/6Aa/zWAlRSbVx5tWMms4vcPqH2fRkgiZlXDPTxDXnOryIqcr98XMEnd79Ip5w
qj8uPhDy7LpSFUw04EZojN837+ocLB7Y8eYYkATPZOXQuDr54IcxQtjJtitFsmUz
HqPVimCIo7nzNDuaot6iqrWHsexbUZWBZg8MHfVeNscbxdrlIupJ1He4Y28m/B70
EuYTHdotsYd76NwEkN+11Ck2TahwLVbBLacyZIBVgLEivzMZkwj7AT5CD2r8wx/t
3bbEVLhm15o0fDmVcnpJwDPBvJVfLbFpKjRU9uWs7ybW23A7PYvDTLm4d9qv7JKN
SNEEnIiyhTtmwxZYch3CXaBUIrVebm7kDCdABr0YFenDJKYL+UUfTa4eo5UIBGr8
ApZn85Dj8mZ3SUCNNOnrqI322KhnV1I6NYMcZ5gUVCSJDoeQF0+U3AcH8Z+EiVfW
+/VwPLMdZk3qV1QWVIwim07LvXuQuVuY26pp8/m18fiiPZdzvXfparGbY4TxIWEB
XwwX+srcj7o9QGIl40Qn9+eMDblLWwUMDe2VzUov3K7UQglS8oPOT1JnsIY0Bs/l
nJSypoS+qWGxRSNgbtYgRipneTAiMeGx4tvLKl5DjEtO9OmagLAD82jDIvznqnsX
oB0NnPgBf0ct9tMEf56LYLQjbBAB8frxJkMFt2A4DAXw5H52/KpKS5mDw2eHlhFA
bkKKqdFDZ7YKiDDNKSxnRAhn0Vhxt0olOhIyPb1HuU/JsxIBCAcUaOMss/4dRTpL
J/xNMfWdUsvRcF/JTcAyIdQrnuAyUtqvRlda7Jr7qLERAnVnhi3nkwEsDyv+tToF
lR3L7779OzsuBh4e5CuHvjd61/PQpTGZSNa5apmcIPuOaTiFfxySL/SkHzMwJDrm
d99c9vH30nVfVKHVBWFTy93zTpUjjyE9sj1IoFCbPuZ1fxni8UFV3J9spP6bGr7M
FTP9tczmilwRphAv+pnv734ApzQFEHMK/9YQ6uMD+Rtav9xiKSbejvJmdMB294IL
t2HXMiGndDfksnslvQiiadrSBUGwAjXIpfllh0vFzQc2V92S2+PWvOh1kTshcgBk
0/jNyH33MswasFpXjjETt4SU5Bfd02wC/ZIlqgOYXoJMH9WtBwaJyrDl2Eu3C7tL
PIaIWZn/OpsCjMJtXCGxpRjhNSNIX7AzfLTEAXuVdQemcLK45L2OhDuxKc/JwJK6
xcRN0LEjkEbY1RXExlsW7h3co1qgx4tQlrpQGYAGS8E1Z8cKIDaiDE8UGwnNuuZ/
w10A3f9MdZtnEE4nKFg0h5ya5JZ10aDm7KEsXFoy1nea3L6WUM7wZWeARODscpKk
alWXyV2Hr7+X5dCCQMiqNZqmTnAyUnMctwM/V6Zdj81UNUURELb3Sr4kd65Bt4O/
xGxu10gi00/zy9QRSkhJyCsSJPnDOIrginH4rjZvbo5dsWeUXgYPYI6scf3efnLS
c/bJx6VXuxd2QkXd+MddqY9VoMg0Azw0hpba4388crymNb5EQohSpTYJWtjMAfe+
8q701TjdKZRHeGlsPIfx1T1uPSmBsPm1XY8CaTORy7Gpt2A2Kz2+Bo8jRepgUgmm
jFrlYRECWWL8vjGO0phJibihD4/oTqGHIWky8U0tZdDfEI2MAdHi0rHwpFjpCQVX
bL1B6p8acb5dfephSCQ3XGJCt0HlSEgtbNZJlcKhRJSD9wmekFj80W8CFtzrZHPg
NUVI32ihC60j2FgjV7tYKyNO7k9H6Gt6dPECpF4B9JtwUolG90vjc6jTSJ3xX8fK
dbl1HnRrtZp3u88XGs4+wVbtiwIMC8Sy8b7ujMOPEsLs+u+b55XFZZFZmOvZv8Bc
3cuV1LndEqwzR79g55JefmkICTBUItUJInb9uYwjqXe7LfX7a7K463Re8tflNnmn
0FHpKq07vZF2G3tWGojeCItTcPNqz8N0+1xoFugVYleRaleDher4D2FM7rxU1Pq3
XH2Fr9fP8C5mr9KOkyilPE8J4GomglAprQ31Z3jfamkU7XYBfjL6/KEpy+/kxRM/
5RhU6uu6n6srKDXIhEI5AcsZ+jangtdqp0ZvfvW2r1Dse2DZaN4qCo/1NBbSvHnG
rFWK+ArjpIKvKzGNj5Zke44X2GksSQf7ymVMX1CaxmwjlEvZoY3pon2U+mKzD/bf
n2JDqEyd7jI1Iyun5gH1brAqAILSi696jY3+t7fsRH1DzQ1ryQ40qH8WbFrp/1uM
W7NM+N32M6/1DtdWChW40iA3hRG1045CTfVvD9x90abk2bXA51MeBtIaxc2TFi6e
XOFtw5N+svncUE9mXnlitZ7qSm8aZW4K/htwbgB5k3+tgLwjCD4mKpQtxyXXrDQL
kJSuEWeFvlKXA2h0ev2At0uOGmiEbHY/FwZDGmWtVgisIS36qiLOcbcIFeWF8dOu
ml0h0NK9UNJASm2yhJBwxZEy3cVQdZoN2GniBs6QJMCjpghyh3wpo8JdLjBsulTq
4sX0ZBzGd5AFaosd5icO3/17w1CowU2WpAF87DRZ0fr6LgwXLN9QK1YU3WGxR+c8
t9zeacY6ftOgKPwfNnpt8yuSv5BcU/3+YZT1978b1M0os/XXndDSCj+OenGIBXc/
iMKVn+fhM7ODvQqnUkIVX9OGxY0p/WX3YAb4SXZ2ouT5SKkV7gdW17fOPGttkHgG
EFClFvnAommSHPma0MV4Xvzm1vlOUziG1J/Tj2O3oaWhbwCgdmTiBqqG9c9IILpF
c7cKlVSGf4PurZnlztwYNWc8ZfIPyJ3wTt1xxNahNwZV9g0t0ZxWerUsJNxreSSp
DPWaDVo9KfG7B3bO7yi5UswIiPf6L/5BVbFu68HmLNdywMMxAIcijfIDdaPN5bX3
TP+igTZ2y3QKw9NCVVoF5u36gZTt87VA0qsUKLdSlKinzca6LxjdYWRtk47jsm/J
a1vSYvQqBKr8pfaYpcPF/l4W1Qf+W99nEYaDIMQFJBQRE7a64LOF/2/bH/BA7rwQ
ZTtvHK5ZA74d5/Mgn8ajyJedrgITeecJzFXTUml4dEDM/938XFeuCqjJ9Wy1UARB
OY2fRfKfbO2XN2JOB6DLTy2zWYf/UfTJjqrmqWWqGwTSHFsxKOErn5u5TWpwNDFf
piM55AlaRG/aVHnzVLDHrDN8iqM6O4Cjj5E9HTZ8MHsM4K1MaIhPQmvAfYfwpbtR
kF2rPbwATRpW46OKpQ0KIB9NbIjqmC+MNesNfUpxmcklgfRjM92l5zp3xlCDpf/V
/wxfy3BSxZhxOOWq/Yizg0k3IjSXsSjH38SP122Fm04xEPa/3J2wlF/HX5mtPfqP
PYbzbvCwiBwk3YpOx8mk1pnye+CXM+aNJ5GhQQDcM8gQeuObLiSqI5XD0Y5LqyHp
g7EauX1ysR75Ryk6t45R/nZVkEBZDDHjt2Tr5gqh8UKPiUSB5ZYJO0X85ehSYcI5
V7jDEE43NW1N8MTwI8LQxmRsAtw1PMXRdZt0a8WRZPzHTv7joGFIQYfxPRPSRHNO
Mhy6Zl6A9dWKDsete+bewSlYTNxvdFdNj2pL9M7gGmylZ5sXnOrROVKAHSV/Dl+N
nAgXDSBy9RrPW0kbGfVVpi4J/3hMRxJrE9TcSLWCCDM51VIxDQEx+T97rLe/Lcdx
lfOhAl77YRRdnWjWgS098jFkXZtFyRjOnINLIGJ+L5J98gKOaz8I50I5b4tbpy9G
iCZlVWSzXzbmM1j/dVNURs8dVdCK8dopT9bLcwnSykBXSjuwbMgWLCECPr0CVmgi
hLlAN/xAZP4F7bTZQ1eqyEZWSGPEB1bZ8fyxjr7JyBn4W9Ob3xz5ghHNdFtZgYLZ
3RQZuZcQDv2YkPTeka2Z2+05bhDHrIJW+CzU2+HfObZAbZrw0qH9pLGLaVO1uAjP
4Y2qB91Li0QHXoDtjYA6xMQ8dvJgLxkASM/gXkzHBX650UjukLm6chvqwWd8Ave4
7F9cMVVb0djRoVlD8uCyCsU/TRo0TNCe1HWKN3hc8AnIJgg7bLAckE5g9pK4gOU3
3/YpmduoxQYnBYWG6+/RTZeiB9adNGDUcu0JX2G5n9kyOu8uwlHtM0VriMlPYt/X
5951p520VjhMYRHCEH4V0OUVBK1s1lMsubqJIsDGdQCIOj7SsJvisW8GFUmjKlxK
Iq8UVs9UYp5VE8iGkx+HpwN+FSgDI3kz0XfLUedXgPWKP62pJqY4yuE6HDxUsLOL
PEJe1h7s1V1uilu0WS2p+Ma6n/rVxV2m2xWL8yOTkVuYnTUtaSMtYcebcpwBv0Uy
Q1OxHzAXKTqn67KLbJEzoKKpbL/SZSOo6G7ruwIfJreGW7WLhABUZmTvKSC3Kcdd
iu416CmielJEIxOXa+fj5hV4Qvh3zGrJJgxP2SykM6VKgnOiO6FsqeRlDcGoYyrI
nlLdEwEb698G5gUwxBNpkV8+PGVLI5duk9+xRKQ3hQHsSc9wHOaavuTJp+m6aD1k
TF3Z8908OLm/WBs1Om+e/HNT9aph6tkJKvxov8AVUTmMN0wOHJxA80g6Ujp/JPx3
XRqESlYJ5u7SpfYh3X/S5r7U1/qiW2yWgp8Mpk3Wk8iSAj9bwVmuv+nu36q0K/Gz
1W3SVzwoo6Xw1KHaZi4YYsovFX6RLOEdi8LbJqI9OSZ+I7fG6wwiCYHRUZ2Iln3B
EF6VnaMCt4HI6uEMqA0yJl5WhrumiPpb86qip2Hqr+yvLpxxjRcG/4MVwc8DIVV9
eDqMUfygJ5djKL0WRbMbM6JRdV1NYHWHN2AieFhSK0qNl9ChtNnv9RXmsFZq/9I5
SAeFoV+Vry9dd4a7+tVbsJTzzbyeR6wb2oDy1eNWnljGyJ2QhE4ehIIOghZ2PWeB
89dVbub5Oxq4UtBaUi7H3+WlpKz6GV1Mbez4YZ1yWIyO0ZTbEgcq6IGbhiw2Kqpw
w5+m+jIuNT0SvSYGCJ2vFANIQFfojtjgBE3h9tlyXNSKqPLRbkXlpFX9TVMadx3i
7bDl8oHRZq8tcErEmI4bNtpjmEEh1U+UPsRCqmJt46uA1LHJu4db58BzusZIH5bb
pw4yag+P5zwJNAnIF9lrtkJimkNkZ1zKA8UMby/zrsT6h+R1ojr8zxxd6pVeURPZ
zRdGy+73ZLNIH2xNoIaUXdwhtWRE9IyXgBhbN23u8wOcg1ThT/GU6q7UJBe9gjik
bmm42CASWUmOsTfiI48G4Nm4GeiXVx4X2DUjrT7Ws6C1E8juqb1mFdz6lRlQhkU4
HYUKghDzCoslJkOfS6KUjxtcphvRHRRK30x4GTT+7+edlVfIsQgtf78wEbImk60t
HL0Unt/IBPz2Qgds14vv+8PmjxaoeocpcJ7gE+j6QkmpxFV5zxNao+Q56QyoJ4Tb
ZOYlSxvTAROXmG8PYn2NSX/4PdrR8DfoKot3cwJKS8W/xXC2elr2OyS1pQy48DoD
23/tXGf+Ke0hdhfnqm3LbwpfcQjYKXGNYwIfSnse9St1R3hwRIsIRxWtx3ZdOLkI
6RUI6EgzxVekO7xkffZJSO4P3nKTEgnhbNiFlJzt0XOdWgadzWdScgyFIXK+H2f1
rfT+9HVPl8RBfikl6VKHYlpFY5KOEE+EhSL4FM0nhChtRNEC5Rznnyv3nYIIDj77
Bfc6DMBuJXbqh9pdkX3SAW6lCylCySmeDZiuFjwQYMV/cBJ7ANQcFo+nf2oX2U9w
5SEyIVqKYzSmWntWYO/U9BbYbTi8wgVb/KZrtd/94gXMWaLt0Vt0gvNRkLQdl/se
Q3R2yATzWtlxy2SdWNUbr1x2J4QhXJhdxciueijbsEBOLR4nlMHHY8A43UcAHm4d
z7KWmnvAkMuF53vyj4DGDT5Dc3MfoFnfaSwExa+NEb4r/0EZVOzR7hDlibPHN9Yk
BI96TeE0c9y8UklV4ki0vVr6MpBv+IOSbTazD6MqbRU+BN4xgpp58k4AGH7x0MlL
majgILYObCsDVGFx24RmvlQksFgV7ldp1PMaS6sHKG1/QJo6GMvzP1VKKoxx0xfk
+dA69OpRPwTD+74aejrhJGjZnanubLN7Q3WbcvrBHhBIVpDi5aIM4ylb8Rudg9xf
NhC2Q8Hr76fgrBU9Jeb7/ytbcrttUELO1goR20Iu6kwNbuQdh6y24hya6RNe2CfN
9ulLbV/eT+3n2MqeWp28i0JL0B+ZCpUsN6CspNu9jOksH4mgjjher3p45wH+uxjg
OHf3y+A+dlUAuQ3Me0Nrlv2XrI5+cL2OzcghS6oy6qCilijtKpFFhwzrhWAMPlNn
OOzVS3vC1xK5+Zocly3THou/ILbi1LHIAMVtGeIcEoxWNFQt05TW5qtm0AWvkNrs
tsQYXdTa/iEx1uVI+GlI60pyp65q+zdGxRfeGCVBT0hc24HR1cGlJNLqlqOEB6jJ
h+Sahw37w4pS/I1A/D57kd9Bzn2m+oLPzsU9hPNZsouge67wpzU7A46dEkmCRE2U
HFnOQ18KVABjoBhyjIcKwlQnKMS2M/0O87SqVrPV6vZiIBCGYmh9JStD+ZHGuNv1
5C5fHjeHNUL+HB2lhYzdGP/XB+U7YvBH3d3HbwhOVLoswMI6LOSJwTnuYVR4a2vO
7lR38I4UhBpNP1cLsLuqf5QHu8nhzUpONpL3+ieVVPmSbezYh0EpHAuCk7YdyK0P
0QSTfWyJZWVAIFdpGFmXE/qDy15CN+2gVzHDcAnyB3fixpiZ3xEO7nKnrZ2Kqeyj
2c0hB8Xd7YegdUiSf4pItSB26c7ekOCybZdfceDQeYjpViQ/v6L+UD8DEFHDSJsF
oPIL8L7pMdNTfBJ9W94I+BN0U4J7+b5tIv6i+7JEZIz0/RqDmEzxscfKTbFYxKgi
LD2OTJ8GfoI25I1ZVeFyCE2vC3CGME5iPtP8hFOlOTAKa+W1aRKMJjUSzoCv/pXm
z5mXIf5NH93nzcxspu5Fz/hIPf0ejerCgvrbDl1iM+g=
`protect END_PROTECTED
