`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRMD2Nj1VTBVu/v1gDI3LIFjb+dteSSyOOfD2v2L2n8y2YpTZ2ieyuLQFkq+pmqE
aEjBlTi4Mbw8FEr8zl7yiyfkE+3Q4Fl2v2cEsdADhCzYK7zZE13YRZg4N2anase5
vftiwVHa39CwR27E6JE3CPoXmgUswZjxyOOhTUi+j/AGniNPLr097/q9FJ2y/ELm
hD03EGp54s9YcuU9qz4WnK2MJLduV3s1Ma0GozTxqVsJ18V7K/fj4ZSz5ZfwEFu3
qmeE4OBaQ6sj1yX2/ZggyiNZy04soKlvNaDSGd0sfpzMOvY/co8ySv7kGvToHF9s
exmjbqyTV7fkM9AJ02syrMB2jl8s3eca2GEXKiO3a8P/P1b4gM2Gjj50J5Offn6+
sDIOnV9xaSGuPKyWiWuiDXSjshfeAFgJW58dohkzFR2o4kglnL3SpgInllfYccPj
sk0I8ma8YqOYtu6KZntydDu9VRFgGCq3uKhw47oz7iK3kk+A7bI/jrCME91ir2+H
XdrL++hmjyJjCAR2nGOqd1EnxzNwbKtcMwjuWZ1L3pwTldK2Uoww/TSoxgoI4oUj
OLXHbLEYnL6KVrcN5jxDpnBIW2R8JbuK1KIkr3457bk2Ix1LJbSsid2IeyDeTCQ4
q7wn8QM0SBymo/lIVPDYv4jPuk4X9F3Khb3ncZBWhM1yhwenkJGxohcYlqq7qw3z
39N7DA0udnQ+GpwPzluuvjiVrypgaE3JsG0HP/3vvn5dN8jxu2pSOQn/R4lwVmnd
1zs/98/wP0Pg/UVO5l/Ve5Rf/tMu/O7m/IX1DiOsxoce67iUeFKJmrpkuxJpLJkw
9p4j4Rqp93i3Bn5x9TcdyISzTRDP+/HU4SmdJkGgSfWmbK+WjJIVoFSnowQnwFVM
k5FZRtUS5Km0VfedSiChUkvqdBZEnGCULToC8/ZKRoOHsM6gN45fN3HwCtvnhnNh
xNNyWZXJjZ3vhtTXOyVvt6EOb+Ewk7BNsSsaOYflS2Wlul7nYwo6731t22MsQra4
pDb/3LqOHQuMB8/VgA4v9jONA3xk6ZTybCm1XhmGMJBhBj+e9ggF4XTeprklE4Bd
jzj6qxbNA3xSFFR3Cm4zuLafhWSbe9doImCp5D8bpuZxHn4spW/E3KroAa9ltkow
8Ugy5VE4aGJga6yUMjmStzkmVMC1My0QPWVyRWn4cOkMtGVQVNwXDySd/BRQ8g5g
679eko3po0Y8Hp/+krocR06Txe+/O90TA8wO1B6UH9A6LqTBoO7Yu/Z41aSMLqNc
G2BS4rXi6nPcwT5V0f7NNAiL7mOeQvEIcOfC6mOfu4JRUXztsSc6z2i/EMfqBYBx
Xlv9RG/SP41ONGhrchMrgEgxYXhUI/Cpyt/evLtYvZJwoiD0sJ0VMluunADHJxBI
tbxnFpHeTd77vfVmajOykIV4ov3cWuQObFan34n9bRO52Fl3+FU/dMWvGh8/t6LK
09IqHU/UMtmSX6TeQ8ip1SG2Izwqxo+wbJjjamJXdVRaZhKrVqqwFfzVANA8WVRk
FaozGv9tbjSwxU2OiW2nonbJUAcPNMttn/48j1hp5jZZ1ZS+/VNedIhSz9thFma5
NORsAcwpLOY+TG/p2WMYQXn3tzZRuNN7e5m+5jalPu3jHh9BJCvBW4NGihHwO66c
LZ1cwUMP+/T9PO1XD2eWFEogPRgkJAxF+c4k6MtHuwoGlvH5vO4aKf3QKB26Ike0
MKPVi/Ar5HfcxNFA1nzfGnmOSgk0BG8ROdfM+pS2aDpgqQamdW0xPhCpPtTYq7jO
4rp+jlftxrDB7glesxdTZMo9W5boWX7It0pffAj1nnrdF7gSVLUeLlSA7kBGQJq0
tIbKYlujwxGGeKXg8LQVg48m069l7zNVj2FHyTVhu1saTJ/z9PCfPefxSTe4dhQw
XIMY8TFvJeCmWSekH11fuUD0i+T9bXHiZw9V0ywT2EkgyNJBnZGnk0uf6w90Duwm
B+525nTRcIyWUC1LRlFQaJk775w4mgF4TX9CY80E12k6JKSXgAVnI1IVxniVBaAr
U8e0Li4OPjrr/NfBJfGwrTb/+1ID3mptgSZ7yFNGt6S/niyuBk7U3Mkmu2iAVQWP
U1e8ZlKZSVXtPWUhAHdDdcEc7U94BeBnpfzboBSOJ7LQRY1YIuhejeBJQhE0iuIU
NJZdpKFtLNVaC3VdeCnKSgNt8HvcZXgNxYZfsWHXmonfyE7xKbJPziTD3TO+aASV
xwigmAJUYzTKOcc9qxjMVmOkdmxZBVZs2Wn6UGtpXCVa5xk2YjminGPWg4gFX1rZ
A4az5cbAfB5rGCMZaEm6soUu6s0mv04unsLmuDcYeVnUqUL5qAXHmapAN5ZeB7P1
pmM8eTLqpBvW7RTR0h7Zi+werbF6ztz/6M09L/9BRWYgNpPj/c1o6W5mtDsbvF8z
pH0Hv2vgyzeLMu7IeYYENpxtYyRUvRqUqZZ+rPcTFVdfkV1yCWNXZgCs7O5ABzzX
J+Q8fYv+AVKjjpWrDqgVhbGMI/zN1l1wr9SWys2LM5XKvYONxPuV4q3b+aX7vNq+
ormW1Qvol3nPlnFQfp424sC1qP7bnVOq714NyuZ6SOthbxg7tE/lwoTDsCRyKw/W
q91XFinbYDs+X+DDYwrSkyPoRpgwcfSQAE/f1i16N/+AJVyADqJUotq0e9bPSiaC
upv7kcpP0tR2WAXzQ4p4xi/M/4ImW6/MbyrZNFBJmsEnX7++EZP5f3fXSaNOOtdX
VsKxQXJp/yzIlg8suSUaIPWUoqELHaDgbwELJOgSsEuiBs1gAMBQIh2TTFlBN2HH
LoliXUep8GTA3osnUg8OUNK7ph8TCa6fFd21VOMQqqCbzH7Abk7nhr+q6ms9FrWp
BxRN0tJeZnN+XQubzCVzeUe+yAOglQp3lJmqbRK8ciSgkOgJbyT/Ck3dmI5aCHe3
Wi52K3nh805y3Yv4RF0KjLZd4quD4IhoQK4tEZgT2GSfCEqt3DJ+t4NOsgu+NK8j
vvCw+EEnaLQXS8zTeZQQOHZugOD+nBz/DECtUDUXYqMBxE8Ft5Esok5Ix8tOoY3Z
cQA18HYgYe2VeAkMrLDQOWRd9Tv2qPqtRrjtSjhE2v9CFJOstMr/CgJEr6w+2aLd
G8eMvOCKBqqJ8hDQRJaakuWVqCpvjVwxIDJX8c4iuqT/bDEqPmPuh/llTZn/iQdf
coswPRDTN67T3DE7ik+gD0l21ETZPI0O6onhC73Z+InxUAaRouLk4twVK7DcDpuS
xBcHgpm2o0uRRgqF/8fdR+SL8fruVWBS2U5+7xKvvKLbmPjib6IqPvrtnBoOpKGN
6HEpc/rkekzBXX12IAVv99T9Jo1yGT4CA+2peDk+BoFN2n1emCzs9rrocM50lwEn
2gyGcQR6I8rf/TKxF7AtrOO7dDmAy6VSvjEgg4rDBczAlCdS8bCY3b9eEe0IOVIE
c3snsb9elQqpLTuNt7FHP5N2J4cn67PDK9AaAk7AXQx3T+ujPPBsEfS+hTE5GlkF
cAn/vCvnr88bfhkghu1niI01/RM6Cxedr0lzsE1E3bS7s9FvYWwkCE0ub43JE8+D
RS0iNI8rb0AumSvx8PwS573gl8HbaqWhzXvQ34wQI9AJVwEoMqs4v0/tvowq0va6
cSCJ3/IkTob4/kYIoMPlCeITRkI535LyrVrj2jffH+g=
`protect END_PROTECTED
