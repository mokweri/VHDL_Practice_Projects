`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ipjc6Y7g0AmlG3z52yOvN5wyiwk23VPCYW923wbkufLxnaKMCTAskyWx1tvQesXR
D+gmmkw9w894P8U63FMobva3V/rAYfCBqGBR/pTNwC/PPff3Vg74KeK1lDNVDEso
jaEr1zNJiw6atCTxqqpURJrLalNMl9MU99ZFt99O+n8ZOI0bSQqmgJr3UYnz57k4
lYfb8T23ROUjGSoQ6jBKRGC5COoL3bSQvcD7et7E3JD5iPPam/KPCMQKhLSaL9p1
zrcGPkkdWs0LEYwzVresiYSCzcgrQ3+XiJtE59tlYzoOwGCf48NNHa/Aaw8qtR58
osNvsoN6kyHoLTZmHdZDupgofJ1f73M0tCd3/bRi0+WKFnUUsOmEWn1iBg5v7fv0
OmpP91cc2tROKmr3K8Muawohzpl7PuiMbcrvgh2IrVS+UQwIpbYogqyeE4x8CMzD
fRl6WAPGXlRCW31XMl624QcOeGFRsfYsk+j4nd2waa4+YuFPejKnYr4gZqO3P6AS
/A/KnjPTkEGjhRvq1PDagtpradTnk5DN0c4uWceQZaDygZefUXaVGc3zV4CF4tcp
2NP1hjvoqh1X73lg3POLU2jAJ2zNeYcEhN5HIcFYmPlP8SD+WNPv+SogXThzz7oa
XlgmpFMTDu5S/rz3pG35vxqHwm2jab9GeACrBLqivUr19rYuj50VAKyuQGwymUUC
O5cSUBOsLo+qDTKNl+a0mNxhJIxnbGnWq9qmqbY+4Itr3/YLfvwNmvp89GFd+W+e
Nc/XFDqC8TERfXZ42kbzVQhf2M9jdSt7VACL+oA9scfACJ7atsKYR+4dX0i2u8JM
F+XVqa8DK5sXIF4dNiUiSPOBuYZFYpbsD+H060UEWSWX14y955sa5ViwDGvO0Poh
ybbQSBT0utFG+6C6DrZWO7qxVAEw2+Ey+d+43qz7RWiHJ7Oj1ppUYz0x1TVqZ9Al
fcv385o4Kk9KeD99mGpyS/u6Fr9PTAsJ3MpJRDeC03KyBB2oNxfh11Y0VHCvOH1R
pIabr5cSqYdGYB5OtMOk8LwNxAsJzo68ScZHO2J6me/sv744uZwT9OXMqNE3Cioj
+j/zzkHoNSImFWw/x5izJxkHC6udTAy34nNbsONLyYWxzm6SlpljtBaur2WZzFGf
nEDQ7W+OIrOySxnVCYXMgGz0svd0WpljngokhMJQmMQ38IlesSQXvevzL6rPTI8I
AKghZaEGInE7u7zpiuxsMBNSwVYgL616EuPZTyA/3zuo6JXntZDvFpSsN1f17v4p
Kq4oQ3ivpqGS9Cb5AbYaNA0EZ7RiFWqF6/4NFnz/M91aq08j3LnWZm9DzIL3I9Uw
X2Jm4/JLxFlYYUOkLaULzmnSEzOcZga0wEBF0HbGxbraOCQ52r58WcJWlMgS8+9H
jJNMOOqMJ7tSIN0/oyVF5ePSLIZM6QV/Swo6xpCtlrVH4Ocy0ktH4ARmQt7+bbW7
4148q4GdBACeJ0JguSQRmiCgcQUlY23+168lEB3Z+BbJXQfT/ISuysKsN1gHgNk/
6cKj5VuVB9zoeMFIWg98ZtL/LbaZpadKpt6Xoi1lvMfzkv5RyrWirSe35/01AyEa
QJOMfKL+pEOt3+bUthNDXaueP5QlCIeJa5ZJ3Ao3+ILWkG/geDl7b8dMrqYigmHt
KwNZHRFX6mbmUU4rO/YO989HaYVH++uONjB18C4FoiksbEwOXBu4pDUEUnWTyaPG
qkOpUDCa+wgaAnTYtL9ZsSukFMcMY8XEBV0/UGX2rB+9tUzHgwOROgWF6vdfqlQ4
f+1xKrvwZ46ZFdd1eTTJJzpP3kQeFSWwZD4f29TgnxYOJkaxwioVYSqcijE0XdGE
aBkZCezrj+7LxmAbz0S5haQA6dAyjhZF6jCG0Uv/NCWlOlRJbsjjQ20Bg17tc1n3
HfK4NJ+SxnuCGVH05y400FrBQSBdsvaaOva9dBOxL4KWdI469vtIH/z9ZW3t6JtH
w/NMK+z9553d+OaYADgVH1KjlsNL6VBSXmoG21cTbztvmhKC+nHOi4ZN9mz3PFkJ
NcqJbkPHipU9U03/aBIBfpAknxMSqDbh4gbtvkHNrrOSLRVffRL1TPA3h3c6X/fL
07licCVv0ZECTg/lXql6rtr7BmYWY9BI2fW2f0/K/BZY4VtvRMBw0bepqNxhsvZQ
4B5K+9U239xiS0pCGf0BgpQwU7Trvw9aJaObVLFYYYsXxF+vCSzFRNBQdFDp5Igk
lGQUcxSh3SucUC7dfYcmSz/M7UsNIbu5SkHiLVZhrBEIu4Q2k6nHZM3VZWs2ZI0W
sQcm6MhbVwLmrtCYVwTGYghqLhIukszOHgWwwfoxxg91QJUwAcVWuCvEPcD2Yk7z
ro1zlOEZLUDaS/rFyVlWHWsT+btmiSMRa6USy14MoAEjEaOy3eyEScjGM/1JtARJ
/nym/4VRKaCy6C63hF/soUIFxQjLAJwS0pU5t6n9ltEBxuqqasgXIQXSiHRUE0wC
7kYx8XSD22GFgLBaL3HY8ORq2Y6rPZLBAGQr5OK4CWfIKwH5X16YqKLeuZq1JNa7
ml5yFjEJ3GZpQ6+Gk9EPdafwtUTjq3tJx+nvBlUZmtd3jAIe1OjWJ/OQLVfyo+G1
Z0BGrPu9BRJ36DQZJLB5KIdlohnppCjBWfpwN3tM/QsWgKX/NOuf2ZaAvrNO2VTp
BAN/7EJ4q6mVOQJ57cvjwH1UEqMKK1Sx0c+atnKRzgbooVvbjporSfE+31AfqhIm
m85k6tJ+NqFzUM9opxxR/4gRn0Pfpxemp4VxHU7xBRu4DTU4pCrPE95VolKjVXQ0
2P3iNjbvjZNR6qKl4sYAdT226eAl4gwTWmwWlbN/C7L8aONfwLZHF9CdSett6r+b
SH0fgjhPQ/U9r3VaOBfx0yf10KrHRkoUFJoPkaCYKX8UuqGpU/RIyHrwzF2dzzy1
HSBJp6L/CqcUj674HliP+CPkW2QnRWIyu/xtjhmfOLWBdAD1iT14axihtEk4S2hO
Ars/FZ+0o0LlU9uh8ywhbYKDc9ttjhY5vNCyL4VsiHUGPDm2fVONWVP2cwo8f+0B
eK01xxsOF/BvKJJDm2igiopx9famcW8C+8R4slX63ZZi/sBUt91gInSM9BC2xelW
KUNZ6yo/fg/Y8UhP6Ni3sC4wZdI2o+iPE+awmOsFW+779uZus8fEDPp2N4LHJj4Y
xRuZucUp90hrBS2YqHwTMwAn7qBoQbnE+Uem7tBDVkdYQa8X9XUo7FAFW0balPjr
bw2fjVqqCLYybK2FTrhElpCy4tpBPorEtX0P8Zzzp4YI6xxWFJPEt0C3wKS/Do04
`protect END_PROTECTED
