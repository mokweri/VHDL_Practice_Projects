`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8RZEn5MmxHGNTXrT7CZOmsk55dsUfxgJu64iQHOFyy5lMnKq49jQ7nr+4Gy7asx
2qqFV2jjtM3T7lofzHYAJcAAUR+IppX0iBkKoBaJB6f3Rm3Vi0yaO/I35gfAGBFm
+MJoB1jQ5QS+UK6JkNdJSHBeqPbUb3qgY9T8J3vsN/b5XE51OVsuc7LQsC3DBH6/
AkfOQpGS4EyA4MeaxfrxK47zvSmOnqTyu43hRXarEwnMXHJH0/FGqmJccOdy6tOT
4d0pqYFpBjPAWNdoB4jow6PDbSDHZAlJ3Z+dVYgXKP7wNJFZ+hmcPa36J/ZdASj2
JD2DwKCRoFa/Hufl2IRPqWyO9SDywhZD1Qm+qtuNWm6w1lQ0pDdL+cRBd08QY+qJ
7vmxl+/L6v/QeRN90kbl5QfUqK5RHsnBXmlFaDR+huQFpybIfcmBe36mSg6a0eGl
OW5zj9JnKWChBKZLaFabtKyqETrY5UhPd+Gh/juQPfLgwav7Fbr5nJv7awipq55u
7kKx1cG/Jc3bRdVo2qVLzEbvqktoTQ4jopPhZGujMySLDSH1BtUdUZ3BN79Y4Vm8
5RsCoVWoSejg++U7oAtQ0x9MKlPAcmC5ixS4OOAKYnW0dK8vdYONY1EBRyowLAUG
fujaDz+1V4xxBJntv/MQX4mZgVDaQHwzToM5g3hbIXpVxfZZsksAERGo1c83pkQb
`protect END_PROTECTED
