`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaeJ7FMMngjG4ctoSzfji0AhTuqvte+YnfNAiyXieJYQf978eyXYxmPUimFX8DDR
AkPpAspQXYpaWTEhcBroR2rqk34HJYqvbKhZNLNgJs4NQjFvQNNFGRfBEYAp8jyT
jIGa3EFxjyKufna4JXAS7dO4yU3G+gKMshMTEKMb3i4FeqLVDx8PsP+Qm+U0J/id
aPqN4uQFM6/In2MmjkQSNyFaOQdAWD2UkGbm0zAASaIrJ40PgbZT0efuwTGu9f0G
a56BVUtbwCoQOz1AdLikxD/Uvy8+M7OLg4rASJg0zayRGx7D7LxS3X146VoFlwhr
r4XrlteORlXx8XzmceNECHBqzAHetT/NP68zQYqct42XRrI3CrdAClNUm2uQ1t9m
TtobFmHYf4HSjF0nhMp5lHY4ryt5ONdFf/52ncpxXukk+FxvyrgpimmX/FvYkJXf
aJlQIvWjo8Qt8Q4jW+4+1/FQvt28bTpLBcH3IltIh7WFWYW/6afHqwDqxrGlvHnC
LUWCkS7TbkDhLW5CxBTsfkopbsPNqxezOkfIh56BfTXYrPIqd8L2QFL0R32g7z+5
PGm/StMNZtAxCEhNRinLRFKOXDV8LGdid7GA1pzk6Xn80OCV6BQhBTbGyMgg6EKn
rt4WGhGeKuYpLQ4mvdPpmp+oH0Pj//OpvXBKaSmFnzIyGp0FNIVEDyV0imw9/b8u
j+bqQFqdwk9dFYjf9uxv9j0BfXNB5HXnrVYi6Vna1WnyUF+cEduHfISe2Mf0tdqo
E2rYQ4k39stvxP9xB6XUagF9pHmWA2zTRhU044o1muWZ6grwVCpmIHqFLtTYUPfh
kmksRPsjQjWceul3rXtvJfGGcq10T0q/mgULZorb+qMNiLD9DvhcZwcUekjiVxvm
ySKbSz5yJjwxj+ItXTqgK1zSGGjqP6xltFqp8A9Aj3gJxIg196/SJIPmVZKhEqIe
fAtx3qtH2S5mY6d1J9zpVpmYDtDDzvF/U3YMXNGuIq6T+d7Zw7MmJpkvylarqnn/
Bs5qtXxB8F8mjhsb7GQLRpXrvznoKdfPNPhTZmp6CF/bUGbKZhU5U7epNQz0KGaY
1SOmc1i+wTh6plGvUU/qikhjDcOl5NQXFse/pCWVrS/xhOHXRI0z8H3z3gSUTZp6
q9ABUpkk4cnXnL6MYKpbVQNFPh6/kCPGH38l+qL37op1nWBEcacKy1T+KAO4SIXS
9OeFG5AsiPiHWpooTSvEguQC/4tsNwN4osFI6EpJ4MgSX07TPyMM+0py5rEo8hxm
scbBEi3T9kv2JF//N5gi1MylnJPsfLLRWHjHc7KyeHqdo5nxMalfrCZFCE4G7lJd
uSaJgUmOn8YDt4eKJXys4VC5/li2GLke8VdxuIkG5Wz5Gxp8QLhZweZtPeTXVgRw
x+u86oJ8kJ5F0dTeIa/NZffEK5Jr6BleX72y7dLXiB/kijhhwp5xCkulC1M2ErLg
XYhHUWifdxl/1uQO8d5yaA==
`protect END_PROTECTED
