`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfioyI00DwmZLtngNkNIucUM4rpcCYGJZRaMiUFPcSJSz9MTRA1Qu1+e/LsJhhrA
CfSska/2iUCG+ZBCoWPTMnUqkAW+L2rq90M4kvI1VsEVrWzo2vuhyoULRo3fSEBM
Phmi4DbQYrsLv/+MJBswRorXXyvDMp2/Cm/15hnzB9HjJVsSNV1e5j7ojREKjKuh
u2bw56rhJmeYR8CJRyec5sVnp8TF/yNPQKWxM3W7CobnouRqBYG9sdSh/uicu4UC
wX6cmHSVFdB1z1+1QYUaoJ+ZUYN64C65uGf51orVtsePxgbt+Aead//4tkUMT1Wl
hDoVElQHoN/gJcUmxcOgyDCQuvXrIkHUwRa9h3RVH2XkhoR+k/B6C+xk6RdYM5Zx
1GNqpjgOpi5xIdNxQ5jIbHUAIY/BT8pB0T63ITfSXP7B4d2X8Jz5rDOcP2jvnfvQ
niMI0m2UrmsClmm/3S+Vj+7QNfgJM9cs1bWfuTUucNJB7JpXh2pw4sMzH1sQtbfN
5PASweGrB2Wd2BFB5ycJ3K5c2NrPiQqxUXossPRHn7Vcztxnb87BFxUr8bdUHvhk
rkSb5lwFU418iMVAFzOjHblEIqVK8iUZsZXsufSlOy48qCKf++OyLlbAHwmpwv3Y
I2P5OfaldiLfmlkTGXRCdn06aY54n2zJMWsdIFP2GnZrIDXUVAdEPS3J3R6xuBWD
rVXGCR6R7xoGGaYnWBs4W+8G7PyX3J/c3yAmS0ExJzijIzAIgaZiNQmSKJFOPep6
NmjtKn2cJAH6JqxAIOxj4w5FRFao9pJo3tD9oCvC8kuwmP+C0opnjj1345eUnhS7
osX5dkb2XKGDd2xqNIiP6dJMv6n9R8snD3tnYm+zYzFtbG/a7Z5x2VTRJkVzY6Ay
morvHdy4zjPAxMflTBaUiWtSz0ecdcFWvO7TKjP2pGvd4Qw5ICgyJ6FHJr2ZFd8+
3mNJ95zKZoOAKzXWd2Kf0DGZtFJcmjbg0uPWBNt01/YXxnR6ZbAAU7Q7i6NMgImb
u3E+fzn2OkhI2Rk0MUYsqH48YSbGqYY/jxhk/gYBngnwYev+/mco9md7Trojna3G
PzXd5ym2Fv/pHGvho70AeKVdu8IMGpxmktABHc1S/rpL3C6Fvjn7z8VFHVniZqBx
Tk4E5oSB93Rc2MAJAOesIL4SVYX6PROVeT8pNxgPQ+F7+IpUdy38rwYhvJSjB+s3
nYPxFwxaoE5YcAGLnr5kVE5ntYGUE2YiHgpj8GXWVaVyEvQlD7Whs3GRd4pF3bE5
/USA03lt4YQt8ltrgagsLE2jgjr4P8tVqalF0rILdCa1ujZVyNaWgQHSHw0omE7E
76AM/VbU1fMNwsDrqn43lCmZMwWZI7ZrNW68YwqkiPvzocjGj2ZFxhRH0raC4Qze
GT6MNzpAFcw7bEqYOahklwW2UwFcxvpyahjMD/RVJcgGhcbcndbI/PWT2qG4YWkR
XPaB35NcCdZBE9XtmzEtqC5N9d6hYiozpq+CfBXcZjovtV2VnNhxVyjjr7EgfCsm
GiC3cqxjpp/mKpPeA8Y3NU9oBmYq2b37o/pNRqUSBubBlkQp/n12ixMSv1uVVqyp
9Z/YroJomE+91/rBt0PQW5TTx8WwdLC01H6xooK4o0o+2hHw3XKAWnpY60Ic5pI0
mtAXI6jvDqcf28QZx0oCx4b0yFZRLpNk56FWcScKeb+LCSaMiCt1yWUYkyfonqu0
miK6ndFnaCeOMiTZJX8mBkFOjVHa2/7xNGIYuZLBmqZfzkUbX2Is4EHgW3Jp7r/Z
d//IsCnwjF1Ip9fVIurFdYegZXLetjEys/C5A7d+Xlt6zljvBRl+3y0EONFTDewZ
lgSuKkrEIK6oBK+Af/4g2qXKo6pyMy5gUQEERlQMHolvjl2Jkf2VNwD/OJ42lU+i
+NhsoVndl/1NOJDPR9Dgprf2/DdWdGdN2jz7xbwV1HMSsp72OaAc8k39HWLw/K2x
k1HAAkUk9Q5zGYj0n3U7PbEw8e18W4yfyagKGkqWEzD/Im5Ib4VUzHsxVIb877ms
BhQ8/vmTtn7w8p7PDGJiAEKJ6Blf5u0m81LIXLLMSsQCTV+BmzFAPEMSOvnzrrmA
pGCkKufBPNbk/zbZdiajdAi8YDI3eKKMReO8C29ZdKiQPBMPf3q19fvJ8BdXAFgG
bFbT3lHUZj7meD8CJSzjiPSDjKSVf/lDAv1F25zVVUtUN9ROxyIBSKRYPz/A2Kyj
wrvzRXqmm8PX5GjrIKRIlCetk8kTSen0fDUIyPCJqJ5TPDSQ3iZGM5Vfr1o1Rbax
w1kU+zm5LiyPxhRTvPosh+PsnJepiwop2ABg5M/nAq9w9pQWg6iDVxAzHNiBD2mr
P5R4L8A4F1doX+VfNiG9g/PCdAjUTXTS1+Kl8CyO84Z6gLVHaVXeY+YmZn4oDkun
wQ1uQOHiWqZ9DlDR9Xtyu/KLrvxY/fRcbgB8/le3TxhJE8aR5p/Ing/wX8eVucvp
ruf+MjTVeofcZF7JwVl0vRK8ZDF7bZaK5X4WHhRbkWjK5yD+6RpZTunBwteFR2Z4
UAphcggeOohWIYFEeCXkBfl0XNyi3nIoHUB8Arxmx44DXkmh3Xx2eqTBX3mwvX+/
A7I9jCBQImG8bMtP99kUQ49GyzAaTvFO0uXInV2VHaaFhLR9/hZxIZhZbkyL5lne
PkRpRrB1X80hPPDRImz0zIQ/DjD0sLdqVNkBzzWmqc7RkQ7YVdAxH6IALbg19UH6
JgYMyFce7z2OF+n38C8hPUHeT8z/7af4omTCNKQWr4+dDEJrZrmcRjAtXo2ZukBw
2wp8bLnFBWC5eF9r1obl4LdwbRp1hyIWtoAD+fvbDbZhtuv11sQIbF62fSOsDEFj
cwgJJBeS3h9GPaLniSS4ayL0ltQHHpLwmkr0odmKQx1a9J/O8sVP3QtJ/S6YMXU1
PVNhO3pg9aEcUEj/NiXgYaf0+pNFks19Irlgjwyv3aIUtNLLVLtosOiYN3ekW4j2
UIJzitEtotnBA/W9n0p7nLvJKsuba4bliNMQLs71xSpsjubAX7eBdZ5IxLbRyQBp
o9LAlyWZQpFkzIzxgvuYi6XHCsD/kjss6Y5SevuX8n7tZL8Vn+KPCdw7Kihfaw5I
iKnx7jKK3O+zTHVE2YpRRZetjW4xVoITO7o0/wBjxCHXrLKwlaJ2o2NjSYdgB9T3
0vxhzQFVuAleB7xmFz2koRvWMxoMBuBlaIOkF6cJeeRs1N4TZGGllGkDf4j2Pv5i
mTYcMuGf6djbTuH3J5WKAyt7kdaifexaJn62Hlax+u53gUTSA1v2wz9LBuOEWXgd
Rdu7tJolCQ6+oZHgduyCo1fNhfG8SieqIrJd5oefqpbcQGR59wbG+ndmS5q1cN0d
XG4orN9jcyPrxwaYzZEfoP/mUHXvZaNJKeamJn0ANyV5bxJ1PZoBh02HHRk8V0zX
5K4DW+P2aST6OKqtl3XnBvjSS02Ej774z/2CUDOFwHQ5uCnv3nx/ajbILJvpi7nN
FvkmquaYn+e/1G6wYiEfVLePXvUACFvA+9GogRplE5Cj/rH0mMy+xNM8kkTaiXFp
I45WOLEhII9amxRGInvCVB0fCRyWkTLx+pEe+oBgK5MyGEjpXZtN+WmMgqA1cuUA
HSboNXgCrPy3+pQ00w2nqdQkMx2LbOWaBMQHFdkom1S/XF/5z5HgdvS/EsyX19+a
VpSppclDw729fLzuVKH3rR7ZCLOunosXedgBbENdrq3FCDONIyVaJnG0xfkO5V09
hKK9sNSHAkAwlR36vOWDIjxsrtaLE/UVlTtZqEQsgA/SywA8hgNh+CbbRZW37nR6
dqGDniC6XVYEo/Nou3cVpWHBJsOlRJ8cmCGWcY0oyt2zAxItsE95gjeOq6WU+k5M
ZwXrKAhI45yXoxjXsmf3aHS3DhNIKQ5tmFifABBXqBFs0uFWbaET1LjxYjRr/3uG
vockXqLTw8oqMhtJRLbWylHuu/G+/UASsINi+zCiiS8=
`protect END_PROTECTED
