`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWaOnt8PhPAlOO+rpXI3AWYs65L5CCNE4xk288YjbF4AMrZxoSMYUIeGj1/gcnRv
FjHbhZG5ZsWAyqqfnRtbnxJ5JETVcXQopVDGtNPUPBOQL83TJ4KCIJLHarLsae0c
HbvL3sTLhiXMxgLIefcQqRM1HNakzgenAfarFzYqIOxXBCf9+EaTazIed8PsZ51c
ZhD5FIWxOdLGwClpJAKads4u7hpipBgcuYjrx0x9azsEMXbXeTmfsoJr6Dh4G/JU
JixQ8Mqu04jvLCyjQuQC3/ivp2Xq0DdWecZfcafCWGg5yPou8BgshZ/R98Jcas+K
HEWyQKMc8dnwMRJna/BCf2DwWXAx2WOgsBbJ0qVkLmPCi+nNBzfVGwL/a8jj/nCv
LHs1vRiv3vVziV+y2ziKgr7uhON3t1Utjsjw9w3yebkFBKz2qYsSoW2EwtVhi9BO
yjyBkPnLTK43LgDepOpNjt0TjV8vNkoz1UdyjdBaxMbcSaVyCQsW0D/6501rtYjE
Gk2p+VyeEAJjNtAmMFpqB1R5ALH7PNn/Z/QPYFu7xr1MH4MXwGsEw3h6FVKR6k/g
dVeuq/ujCqJa2zN1V2SInR5pxgW/YJeMiZFxgFZ0FBy+4JvANeq45zkNDNwdOYVj
08aOvWRmPlaVtCIzop+7UAil7EilCkGp243Prz5KgH9iVCkwQxzdktqJltY1k2g/
m4ymTxIDL5FJSZ9McvXKA37X5Ey8HQXEO6C7sDXezkVhlFMnTwve3rZqtEysyuBq
wO4s238CGzn3NQKRPQMpU4YvXKx+DXMPK+y6Eb0q8lEIijsFfptgsYyV6sFs1XZZ
6fLZrzleOnejGYXIgHXokbeugbAJHtr3ntF8OyNP23Lx9Bpfxb9FZQ+GIkz4/EkJ
fEvTxNv4vi2lkZdFzLKHjSfA8JpsuVPZdIy/HdKHP/VK/qCDpjo7rJexGmsLlRAk
zMqx3fAZe2F8HDaCpM9k912EPIs5v3QBpL4be95rpN1Qt1yM5Umg5ySPQZKXRids
jmBMSotT5Dy5/v6rlEjOt6Joy06V5AdbLW/4COiEPdZC6BVxmfnr/iUP5pAHpGSX
bBjpCOTFEYAFwaTLSd1gMG5UBmUuC4P6lv4ACFpQvtxUOdUpt+IrfVMjXR8flpVd
NG0scQpYD8/d9TeNKAuKwSXH+Qcgnpm4aRXH8WZMPKyGRz5ScS5IQ+Cn/+GOXt8f
TqFEd5vNRoivTr7Vjg9aytXrEhHKe/PfTsrKRv7PTYb5DXdyAOoa+V6XGaev2fUD
meo9eJrBNZIKQszJmhBtgznOWZnjiNDGuYR9iK32II4mFOi31fAIJdLDHNymcmay
p9gkgC4fFi+AYBOSCQG2ow/HF2ylI7p+e1c5bKwx0+/cLtv+sKbO8LXa47mNmzgi
UGH0Ej2b58s+DL+NdTpk+y1yelRdSBK6xxAGpa933tzHrH0x1+84nFM2BU5EHVji
vrVsmUZ5ByD/MMGvWG5W/3yB0ivjMrD/5NqY9ogjLESxb3tAqPRk+pfcv26U3GN+
G0zNqwAdCFeuFpywx4sgqZ16S4LFt0FbOoc2G61up8kgpdFFsl8/rUtu2MqFd7s+
JAZyCd6pont5IzfDRdxQpgcDgH57YbohKLzR8b5wG1bQTl7hllaFHO7t/sG8AcUf
52WEa00xxBrUa8MAxdmlyZpbNIM6V0kNyI3a0lJswDSGEZ0vLxW2BqDwlMF5scXY
HJv42rE9Sq17rG3cltv+7Cum+jk5n7EhnPi1GCSbGWsV7llRIMJY7WtBUNVG4KqE
rVVLDvMCMxl9Epw+6NxTilO43gVE+f35xzI4BK/wzBY1xnhZPPI5poEn2DodQayW
JYxunz/GKRwh+BHbEZrgIFbYbONcLwCn2zG2qpbIpBs3QWgUY9KWK4snvuXT5au5
K0apvBrCOZV1hVdPLndVI3dtKvfw2lPGmtgJzl1cjSakKO7Pd5OaQ799tjFryEty
uPuUMWPujEF3vYURuKRetUMDeIicCkvP7dMiheXbeYOoKfXKLa2misfUQPsUAioc
mErewhYFvC9cx9PQ/V4hfonus2DVpCWfHpy2Ds7y/9LVLFA5Nz2kxgbAeT9bAG11
+NZ+Cgu7uLjn6WkCG/gjfgvzI+2D6UIYCks30YuflPSaGQ3JbGGcf6a7fpJij6Re
+hLhTzNrW0/iWyOzbRU59zygMbeZpKVi90bRgPb6UQ4mA8jkCIFuvW2QTijUlEHb
iq3qf3ip6EogTDVJMNXw82hZqf8eUjVQ6GAhZkGCFlDnBqQQ+aoKxWkLjSto0fO7
q1JdJp/aSQFy0OTzFoj0OaetYzZ3FLe+vZkOtfAaoqwEVh5aN6+BaEXKnFBaNzZM
dWhTyYKSIFxfYRo5RK6JOe2ATlYP4QM4OZObpfvAxTe2J1RGFq3EIxA9q4A4WNkM
tJ0Z97mgC+8/QxzMrknueqN42UPUofIF3k/B538iP7OZR9PNaMOn7WNTw8hEcBRt
cbcas/Uw6K3Sxi8KooNjJBsmh4KZGMj0rTdtRqrNShTo4ve/yAozkGcIHfsbLj+h
q+imniV9KKL+3iV9dd1IgFJStl7an/aPVxJFT1Sjo3BiDbDK51KURCE6Hk0BftIG
funrk9r/rbtdPY/SW/46LIq+tdHVXWgCGmSeRd444umTmHvleJ+BuD1NEYW27Dxy
9B+DwnAb3GoxiVrhkfWmPiYfv+stZhTBKbP2Ur1XZFOazB3JEx95KVuv8NwjIiYh
x86B/zu52hr1sKtQhxBg4i+Pi+Va9r4Uhf0bHnqejRz46ETYHMOp+8ejlYk9AGSL
by/B7OSvT/4XbmJJB3Wq4Srvgm2c3NkjddvfFMuJ0lKWdMBorUJRjaGSch9ZwvZO
r8m/5srANSQPmV9gw4vWnIm8ES19JDeUf4YZRXHJhqp5F2UFPNVYu/I8f3JlnoTE
JbEZEb3AEk9pxjmcksJLhenrlvCaWp3NAtSPHfjrRsTHPfp3i9d/aFurz81PsFPs
RKkTa+8+FkvVIl6mrh+eY3pirajcAp76g5ESX1fCeFxNrK4Yv3/sBx6oxrMV4QU9
S7jm+9JQCpp1QqSHD8P+HC4kKO+i9ttYvVaFIkbcN6ZVKpTmIEQps7OLpAU7TUw2
mGKsf2bZ10RdRVB3X2ZQM1z8Prom85zioP6rXNDCsfbUA4TUUmiK9mWqq8wcROIX
GYzQe2dOEkToDM/22n9cgro6b/ns40WHx/QTZnlsjjKR4tF4WLxSpS95WW9PK0Uw
6x5vG6TzVEsqprYIGw1XXs6amzB3uZmJH7q1BOlqbIePxNPFUB041CxtVUhYCvPq
JMNHkoortd51bzxbOt3vKrePhcgd42XISRKnBDv8bv7xnT0Obd/vBVqcq9MqQIac
TDRmhAdRUgFJ/G4W+ZYr1gKdJNBAGztAQKn6aHzpJkq6pVJvpWh8VWlMrZHzCO8I
fhvzGr8ZFq9ttidpbHh5pmvyIJHtepb+fLAI1s42nvBhKxWGfhrHzFR4GxT6SJ9L
eq/QOaxXXb2Mn4ymSa1PIRhUkNKcP8ZgfxE4981CkJdSX/WecDatRg/ysP/nbOV2
Vy6z3gAtjW3cWaySD5heTbetfYSJa7KLuns3is9f+Re22LMU/2ikgj826iggtegY
wdMHF+Wy1CCqe2Ez7idtwteNEW+gPPjrMQWT+FhOPfOtQey8vI6y22F5ZGzYvRHf
8g0VZi9KNXHYKDebBt1hbFu3/+kGb2rFX/Yfa7Ab+vyDMcrJDmfHhm4tU/5iH/0C
CBNX3qMIRBgCff3/IML6EoeFc92dyII8TEV87g1qysuI8ie5qSxPUfwIqybSbALo
3BZMhpBTzU4aXE4M29d5v99FMOkySZa6FUYUx/yx5P1BH24BsfRY8FS0wx33UGIQ
kipu2wmFiEI4pYnQLem2ayqW0DJv1026g+oD6jTEVcFS3Aaz6jXvX9rf/zKa/XQl
vOTHl7twmHqFUg+wwiplvhTpk9P1LAPahAa5Eh/8TwX3TVQGPzKhSfMqKiwohQ3Z
oTiKFUupFbwlxc3TsNQEpuyFRib6pqvd66e+aDIfT9conVTAmI6+kY7RmrcZ0yms
hZTjLvJDMHVArM7GAZ4dEe/rTOaC4vCmKm3cFAhTPb/Z5Z6idPgysTtizXBP6AVP
hqlqFcd4QsfW2+7ymAMPT/ePPWiqq4k/lrPNgH9DXNb8K7rpzjblSBrp2qlLd09u
wt05f6qp7zt7gJgi5OvmhgHsmiJkaYQbB46yUd8PiwK/sujLUgq7NDvqpSli5BIG
RYfFgaCXn6A6UaKp5vfO7Yzb9Oa0eeY1Zf/e5qhQ25NnbbFrFbn2+3nJHPkKHeAj
yEgCBgxZzeYMCFdtdejAahGRBEawM2Rowjylbe35ZD5ZWC9f3hNPTCHN2Iw91Z14
wbRYjCRWuVcqkWTpZ4hqDcj3/KhAlDiuCjnuQp0ZHlYAgSxEBauBgDK6HmQ/3cVF
pucO/BoEIargXfgS9SNt4KM5f0GYXbp+cZ7TZZGp5WcGCZCOptFgR/pVVhT6mS/y
/krV8f7VEAOAJVk/i2y2a6HrXlqEGMtAe8RxwP+3Y5zz62gNIwqfQ+tX0l8OeLbV
hrWoWDQ/3uFGV7nOxacZRRBDkH6JMX3zjZxxVbjo5/NYMAJM7X9hQx8gJ/8GxL+6
B3aNKORHP8oPPRgTyrvD0XWmiactq5tyTWpfA3kDKNv7zZnwagykFIsZyb1dE4lZ
NlS3RNEAVo0z8/+wPBHhry6GdNmD9C3HdupQal26n3xtvtGpenO6bbz4IwgAUnz1
FpxKbOtvbviQxbl/3TuRe/Ki9O1lV1Rue/sL3AxFc47/1wgUV6g33X0bGuE/pj/F
03aB+wsGTAammq15JVNyVGqPmXQq9lKPV/fwSYOu0YuUCIW1iHCOoojQ0I1YQOZl
Cy/OmCAb0xxWbwvfaSGP/y54SdheWuNxzd2Q6hpvrF6D6Zr8lIszs5QGUIXSSIEi
bTl6vVg6Y30Udl9pYyRYo0lQfIWBKVUwtTzxQz+Bal3t+lXxaMVzEahAEuu9M6oP
97FjEq/xS1EELCqjfZanbCju8TnolBSamklGMJZI3JIohi9gBdfgb3dzb0O0mzbX
7AzhqumOwmHrOTgYGrr7UW1SUdx6ob6/X7E7hIZuIwPhalFSAjeS/8cykefeP8kU
s0MGE+8nCqbcstcpdVTfEOQdqfmnxcrm67Eem4MFfcmQIhnBtE9cx1MVog9XtjhU
Log4hJtQYZgrPNQtMFweXqStFlyCbHRvZYZIuVFC0bONYcpbLLQxpBUYnOLb9ezt
obk9ZmUZNKL+q6RrGSShAxHVZ3VP+MTlBOEnDgs3f5W4VQpUA0EtUuVi1tctKjRj
3crSPOYDyvsokZhl/UkRRRYqL5KSn66CdLrn66RNFlZB7LcZrWK/Maim3Xztc1xl
Q77L97l9cIV+8NMVQeP1mo6hwItT6ijoUM4p81AVxwzWBWjngzLZbwNFBb4kKMY2
S2ERTmImBkuqDRpJrzBtoLS1zlJSZeUAUFHZme0+4l7Jhvlmy8hG8p+8xPs9nmtt
7TYme82iCUVbNDYTv6eUGXiaDiIPv8ZUqZRJJjT+jUslHEOkD8eHr2XTLlyZqpVT
H38pmvTB+sKod9Zl834I+SB2SMF/7jE8PfPcs4ze1/srcYGoWpTghbpwYLHBC/p6
wQo9wG0VHa2Xi5ouxzapfon8RAWd4wlpqmopXkuChkbRaNQRrD3TJocvCMI/XWT7
V3MUxXca2RyI6U85XcdGatIjxy6Pq+m5ZOS/u7840KHI6a3L1Eb0GmGi6xP8efIL
QID7uPpXanlCavRGTwxjUpLXNniIrJg2Qzj+A35Cs3Hs9WhsJ3AwTVyXAdr0ZqqA
uJ9JDq7ksW6xqTQRG63QjZ69mxnjhlCCMa+ShWCipVCRnojzRDy67eW69Z5rR1Yd
uK85pV0KyjP7Vo8O2iOYf4W9F+Su2/wqeQ7pCg2ks1aWaqyR5M7jdA1di0+jLIO2
YyYno5OytPFzFEtWfLHQa2FF0I6avORev9MiK36/kCfqJS2neyxk4w49TJ43orh0
6PguZoF7xbkfNyG8eLjzfRUzB07S/hyXDR8/EZV0h13Cl/8j63dXSZ2GDBCIdDMj
VefottOPh3ZR/ZPyCthfgUPyUI27K7kyRf0zog2jifttYE6H4TPuYWUU7QuWQdtz
2w/935szgwlY+FVrBDmeCgMVshVQ3DZaEcIJelF40sNk9YOqHxyFUWd41wqWfmCa
bX1SgxnuxYicyCLuCuiJPCU+x0QJrBRyRJqPjigZkf9CS2WpI1o9YHCe9Negnlcx
XhGU3n5QbZvCnPviMySn0yPajy94IXm/byZ7mkPRlbi2FUE3qq5l6QahvOh2bFDQ
uXP5dw/Ik1uCfOTuFaq5ftcVVPLTdjS9Jq+ZtAsrJFLfATDmbB06ctbcHEPye40U
pd6nPLtbO05tR/BYEXOVjq9x62XI0aCppKp8ocvdTugItRhhZP2VsVClEGi9g55L
bEL6YYUfpITAVuV+WpSQ0Em0R8sFdW2mfQtRWP0u62XnFFztdk+FMd4kE3cOeOR8
nsn40Bb3ihTmYVdL6xLmlJZikJbwBQLwHTfCCvGQmDe69sOyHHQlZLglRg2rofEE
ulqKEFMGeY+fqQ0uxhKB/wkiq/r3GupDVg+ng1hSDNxxw6f4CoP2m19wioTW/RFY
cuM2JncMBdANycUCS8kaMoa21XjOozgn958iOMmF96dola++LtRGJZ3WkKe44+up
1oROMel1cpA3xcmttQXCzkzJHQ7ghhR1MHA9iMJc+Dmciq/Si2bCRjvhG46WPGal
KFdRo8qZoPvQHEdYWWgaEe6WGk/LuihbjEcYwPGB1mEC5z8n0ooOBNpEx8AObl2g
E63XCmbVaAd9vgo6KnE4FO1KQ7ZIrjmy6etOo5ErOrn00fbW/DkbQDWnFsFaVI3s
Y2TH7Yzdv9a9fMX4z06sknCM2xzdOjflnqddNo4Y569k6H1gPixFdKwfLYT76rZk
y7JYWpwdLWZY6rxK8xNqRXo3l0/JLOH1AYDFDnAi5j3LgVXjhE/DEw75GCN74C2q
wyjzRbKwCf/0LfGOQlW7DxQ20cTGP5W8EFBRlHGirMWChH6IP2qOVoTZGQ4hmVkG
Os4C23WFedwppkLspcyzf/tJamImXIfbrMasA7ICCQtoPvz6td3oov2So9wENB0F
phg+O6xWaivk17TJt2c2v25/3uGupjsc3gU08P/pXNrs0pBZXNHqVY28C1M6pYRo
8fIFJWLtgqRgDF6v4HBifcCVhaMf8bITybiT3TWYzrajI1Vvy1y13ksjMbTjkuAz
mbP+VxxgfPx1v0WvKNuv9aCFzXHUClaYQ1k0AqpII1YxmIlxpaPSMpekDCsXNSIY
Q11GaF2/8soKQrA13dNJ2TiPrtJic6+whfs9K3Be5Y3uvdMg1SZs3Gnv4EnSNYnt
gIZ5Fbd2sUCG4ZMUqOZ1ZGVBrcRMOQm2B3+GCK+mVfaqSUFkmOCOGuSB5pb7k+lo
QEGEWhLwjlqYOgzZnG+0mnAqw9ivGQn5zHY1Tx+qKZcP2e/+nLImUeNLeGf/N6qE
+jOn1/kTYiVDIqwZjNYhNJFruRaB67d37rxDA+r3pW65irBuiKTmhMPN9R7DD7+Y
k5wlgCfYnVsStzcBFqxDIOpmaHFjmFQRhmTPiIQ+OuUmd0YvyM/gm4rSndblWixl
d46+WfftIP/gpHZxEx0ff7JjHNrykHYXlL95ScP4Sj1O1hxMrvDLd/fPl8zyGIka
9rIoc3POFK6b4t8ajQeB2jShzix/zCNU9iAcVPu3OYDmDIr675c9kgCP+RWqlvbm
OEH6+LI0A7WDBa2QAV4hlSCArZGDzicaBen4PPTR9Cj0saQJPdOizhXe+YsrU0YZ
SY+hkzXKnZtFeR/sjWDXhZhoI0n3KekHW4uX/MmZF1SOiFwYAdMDNLZMITjzl0U8
9UFSlSiRhSTqI9ngqEDAorYGPxbgHh8esMOfcOmnsdqh6rKz1ssruTjiVzyHnYmo
EYw0hE1k+JPWA1awzJBdgYaLrmtV0T6GeaYhUdR85RefzRshq7mT4Dp+QtEk+uN/
cH6UZ2nRVeCCIy1snm6SOlv/muF4nHUbKtZ3EgQNfQFabqoLev+qzffyRHKPGroJ
ydRDoXdWDJgcUY5KvM14AVAZSCQhkcs/595XZpyrJSx4aH75xR0PZFlAiVi+KPrJ
Txo87VOCXaeBMlMVH5Ozy8dznhO90hYSyYiCB+61DutG2eQsbj0xRZ7BC/mMuKW/
5G199A0E1blmfFc+TSeWpjsdXl8RwqxtNW04kvvAY1jCgo/8QEO5Y0z1Lyt2JNHR
/u/gJlLXgMbNGCayzIAt47kf+CyGe91JQW7Q6EbS8i7NwPF3Ha+l8DX3muR/HxfZ
FJwOIrNBcyYHe7ShxzIReWDIWWM1YPWqDDjcSFHgjr57y8RNAkOQosUvlPKbENjC
v/9AhReaZccqh3FYBgWrb3c3T25n3TAK1TrB5KvPrYcS10H4J8Qa5TiLCZO/Ae9r
oDRSh4fdfgcj7N8c0ZuehMz0Z0SANtdSSu9L115iCGgAWetji+AEM63mFExf8pKm
4dxy/1Ng31ZOlbulrg9GfEk5hJmMYw6l4w0jVmGilKlDXS1XjkmCTCqLNPGQpTFj
37TVV8ge0Vl+d+lGHpF/zhB+R0FOtLDFvp9K8aI/VNMIaQzb/8fyynk0DV4BPF0K
oeW9O6jg3y43FUzdH1iU40qLohi2du+P4b/4qfTeI6lQZOmOBQx5e4Q8g9V5GoC9
3bm+UL/8awHTH/GZX6SjTdQDU+pCM8R44IomGpnU5N3eKNuMWpm86IHW8OpI/6KY
T6GDUyCmxYV8E9/A5A9dIzY11YlCje2WM03yyWOtXUu/p6OL2QqIPGq161kFS7nE
UsfqTa2QgnyV7RQZElKRNkNHsY1GPJ6hWzu/pfa78vGp81HZWdAPHrcL9uGNT+3O
JpXaYmCz1JoLFXygsH8LNUQemn7mWFpprhF0IJbT/MC4AGoOuiNOEF8u9uuhbkit
S3tztfoQcl7HEsobUo9K48/h8Eu7Ah4UDmNpMLDpnuQvJUg9rO9EBLEQyLWbUT20
qM8IMM7OXv7hzVhUm0HKYQ75MhKoLO51e4b3KZqDV5Dbj7YhRZY2gP9WzCEAovLm
IWvvwQ1juGtRx2+C99dxLt2YtzmS9v/6yBV6lc6CEAOlqAhvolvB4ow+CjCWBy93
Rv+F78jy3QzSFqtvXNphKvSOPwOmksMdUduBl6DtIEyMEGrXdo9qirlcfsP4BAQM
B45Zyq24FlHsqYA7FPBy/5N1+J1upr4bdDSQXsAOfMoV5OdnvBaXhi+SEHv7KaBs
GsGY/pZYhvEZi4Rg10J/LKjDQXDPe9jrDda0gA2hHjuo7Xy8RXCdcc2mcFHsSFge
dn33QwjXp2ap6qmnm2CGOPxhyMbYCG5563rhb3lPM1skuf7eGB6asnAlvHCZQzx6
C07f1AWIjp0YTFEuwvkJ2OQf2hNcoBhIgCE0LzBT/ONQf/Fbns2eCrHQddkZWDDJ
1/4vVZ9b6PNkxwXD4ObeczbLsrzM94gYjOW3C7kgKtKt5PF7ZkMbXcDnEBALoAzS
gjBUwom64arrsnvINJVDS5DKTq2pA4e/MAgw5NFuqSSiS+YNZoDqRZgt8Mfx8QkG
mSzH6/kn5/L56RUw/wcYrqzeqQwHT6PJsckMvNxLgX4YvEcsPexRERMvon0Waf2h
GmdkteYHhjL6rH1GaWvj1xktBEWx2AJBixwqv3WBrksntmAbkJvbKXrVjqU9QrwJ
ohpquA9G7KfS6JgQgHa+qAKY4HFu1nuZ33NE49+194ZUOTZSZOlXtxZgp3WtmiFm
Yx8f7CLVh0t53grcdfKd1IDhVEUCtfFTmhzMrDD+4t5BtniVnOEptr5+MVVX08Ng
IfSQKQmXDCMi09E9PPGGYsBL6pDjdphzifAHKnikooTKrz/F4IINc5ysQJmYlkVU
juLwFToDW7vd5o1Mt7zOL5pskJ6WUiryxItUW6xHat1Hne9iGPDRPVpKU9NLaxN9
qIvvugjFgU+9w8rSkd14n1wzUVnNQHmBAoDpaQBmeBeeZ1/w34VHXemQa/VPs4pp
ZHmpg9VYXVdOIKvFMpqpIGS6WlL5tqhfU5YaVyc0LnmNvxgvHWqjoWJ/517+LvCx
ChYeo5rbbkbXWp3CFMPHWh+/uBQRRMEe31KYb90ZV/Fpk+YhmiOsQiryUmNVIR5k
H+j3Hn+XGxYLmmWm3p6wEd24zF70LoT+HQc74ogYuE+fiHpbCvcXz1/QaKLx2Z2n
CMB5xzmjcUPKzcfbsngAt99ol2ocMCig+t/2vw8bU94p4B88PU8x79kGPl7o0Zju
ywllqS+ydK7Ht6OkN8A97qmeztAffDSxFFlHDQNws0yS841gkDYglbN3HhXm4Tef
ohfK5KVrLZQtylFtbrV8gxoKd98XEU38TggB5llZR7L6fVoACvaxVWW8PjoAZZrL
Qng4YMzgaSmP7lAC5cJrOEZwxUPiybydnNq7NltXeJx6PGf++WU+Iuj/MfYGopwW
GE0+p3Wdq+/pNnYNkssnyDHisrZeDCneK1iLM/VVL6gMtx7doAFYNj9CRMyV+50M
IZd+tdJ92xPxbTI6bv7WgmLokjxj/yjdhFhkNvDcybSee1PYq1lNJTL91fWgkv1a
GEBf8GaXyKj47zQ24PQHrD7TaeiIWxon7Ti0561O0kg//u0i0waT89H1JmSrcDu1
hdYJEKYHvd4nRUGiUcWqGDfNKcdC6jxgJMNhVBnDifbzfbNFNaggngVyJvnv8QKl
E0aYIOV12L0tjqkrA7OWvDaazfEeI6qn14VJnd1/0jIlcc/bNf0zI3yhCZtNu9p1
7D3FqSaMjheA+Y+8Im8UH58TN4fYNfn2Aj5TJxbsZI+16AC5AOocAtR8oj0z9FCi
TUnolnpCo1O33SMO04rofLmJtVrY7L01c4JZpYDPHOisOSyvZaao9jbiluv8uYJ4
BPhV5QX/Li4oltHc77uZaLAALAUQbXDxIYqg6BDoJGYhiFJRkfvc4pi3PQFrYYFc
pANFT7lMPhZihdtY2JOeCJjXYTnLcM4iNKBv7KNPgItdvt1O4HnaeeqAI92Mf+AH
uR9HIMqH4tQgCIXCpBaDu4Ig59FA11sP9yf+UaNmvf6ouYdPtSBz9dajeEICLn54
NVBIcGyEOtNPekbw1Ay5NxzdFBG9oclRDa4drcXBJofrpLf+M59grRSlfr9ZS9o7
pzOwRexFCmpgxF2/B1AZPYCkEOqgyc1rIE/UCfJWaVyvD3wR3tfmWTV0J4lP1aY5
1ewfuuS1EIPG5d9yDaOmgNdddd653Tkxsw+d8rSgcF8Al1vDpNVqhcj5EXdnOnII
IYOwWSjYkwj7/+AZ74lw9UAFA7qaknC2wiFPsE9xqnmnViraSQUh+ZOS1XgUXvcT
lYqzBpWiQQ08h7PZCfjZBFOK+q+Ab/c4HbfAsottm06pwp4AuHVFuwWsSiIbE+nB
BgBCG/TDIoSdXebmejywwp5/y0t94UfqCwKs3T68Ge1wAKcn2JhyxJhWy5lFTcNJ
0RaGCNeFv8ZCOYaofhwQHEgMkGae48FoheYErKb0MhYSvMRTkP80kv/iKjQAjs+s
NsUwJdCKJtd2jaZNojRmmV7sC0LyjJliOs1fI6Aezu3ptSObBzmSAZRMCXTKJI6Q
NehytwFzkdSiM8DFaDU5Sh03qQpYPVyXzTmX/Cskn3749rLcKIMAhGelxTaRDbPf
1FXSs1f6YfUmdwdCQVJNOqrCn7n5ZNuFn+k26bKmVp7I71Ua6CQqrnYeQJ+n09Hh
f0Tv1HsdFhCEDKBl7Mup4ufCswgilJNzRXTSnhuwvV6QwYD3vsCb+J/gP3eER80K
p07x+s0nD4rNygE0d/PBSvVgWicA0thHzHhp3sJ33m76sw6/RwkYc9AJ/dUFqRRc
rBW9BJt0yjG+kH2RU28YaxTaopt95lqF53FO2XR85wShZuLARpS80zsHberHpnbC
ihvVKS9afqc9SRbfH4wqe2it7LH1M74aVkb1QP0Ok22Tr/vZNoUVe0AbDTXwYDYg
q4+T9VqMT3MXvCLR6VQZvl3+BpRUw0p8pIXbUvMyssHYf3WUqRbRrDEB0UihOTfV
Eg04QFwPuTTyHFIQY8zD9X7YDi6kV6uo7fK0ZeuOYIhGoN2OxMZD5dG0PxMHsAbu
fADsV6mxHfOTaorAqQ3uddb9pj+9DHK3+5pK8Bs1+E1ht9oUU3wnEXXRNjoqQvzY
3y7N/XJUEHQrrMckcUI4ngUGHiF/fee3Zf+VdfdWzncOM5cV0STbyXZKhrqlyoQ1
U+MfubJ41Vgh0t7bvmfqQwplwO7K6yTljhEtIMEfw393yN2R/8Pc0VYvhBV8u5uK
NAWxlftbc0hbrLoZJt+kSQzHt8rF+1Zlv0bFWVejWornq9B8EkTQ4iheDltRBfom
lMJP46gVfXQaKMAcaYSVgzHMllculzn9PoiPOQ8jDy6dpwMRaL9XRCm7/KpsbzYp
1vuj8mjR8FyfNnfZ+B+ArDdRuqKBK637gKHjEXZs5KVV5o9CVGJWrEwpJ4juzOY3
CLbVyz9msvjhDGBE+mz/5bddTyCkNB1/ABb0tyn4V1dV8MVu8yfCtz/a5OieS/Uv
U1rJLhIgTADiOL7Z8qaVQRzz5A2EIh0EUsAO7VmlKJn8qSIICB20QlMkErU5vleg
KA/Q7oMN6rHSsHKy0XVIyUSp5Ph67Y1BYQwdXcnVb5cfrN0eIrt3Zu0nurYHe7I9
XIBAjRDr5Yv3xK4yRWHaZxfvps6VnaCyGZJyT1EeNyXMJ1BVkw8cGvFNfiHYpHhB
Cn7XaWdhgFWcvqdf+reklwKY+CpVYqvRoQsZ/kzQzRX8akZo0LlutkSCru11A5cR
yQ8z5DNMNxQvwLPYGGds4eDaLM+GDTehv7cqxAORM5Cgd4kKCj36w9EKHj3ev/xW
INae5oQ91F1vYtiunsYsTQgA5R8ZWHKFdChF8dVVeb4YQmce5jNceY0AHHBPmU2a
WIWzYPOf14OIOctA74Js3Sijdr+wRwYwebrMMDjt64SmIF8FhWuA+KpAgBRtR0b+
HI51CronP9aPQW8lc9dlh+ENTVFEqUJTzjKwxVbqrVaev4pnrxvgnKvoIgNW7lIa
+sGXfLkMwyhVd6x0wl3+9mA9Dw2bB4qra2yAoMO6pzoAZDupacGb8F57qQM4KY8h
YKiVXNmQKiOJgx8vktewEnt0eAJlVra1Mg3OfKv1ZLPzTB3W2sfiOaSZJWSNTHgd
+hxhP6+eZhPYWmjkU56MTwgoAEg0/ApCGbMEK2QFg9/AcxlikyfOk7f8i0zMzwmQ
Evs1/jGHuCd0bQhO/JOmRoXGnniwv9WGHMG2Q9UmBmcDzh3ms2trDGLQFRWijwS1
CYQN8buGM6mu/IwxMunrqMunRUzrhbgmcHA7UrqAIxNAvqetqTGYJYiCbnNd/ufq
HY9vo8y90m/DchSV0bnNWzorcFpunaxicnFpI9/rOPNnUvPhpmIAATnw+509DdbD
o8HCubBXuRAa6ZMmMqz00w0aXHATT+Zp7FtQg5sVcxzMtvXTYeMH5941mOmefJOk
kmmLaOLLjdiBaSThxHl28WGg5JTIpqJYMebDfKd4Id1VpfRzPZIjq+62PMeiX1Y5
tQMO1x1nUCEs4etPncLHgoXYWqbgmgMcRwmjFU3r5/Nm2uAZz3dR6rYoXojy+Cx1
FbMUy6bwj5TCLKg+70k0Pf1/kpuCuh/wuR8R3SnpCjab6ECYu+1igLKeZEORyeFt
Fnaeqepi6C8mqOvuP6rJXNW62sQ5JD5mE1bxSFQ/brCXefjA/Y8WW7X6mC7RJcUs
jLhsOClAIbbQXzIFod35HHU1O6LBChkron/KYTIR7veyO7JqlK+wwgqnmsMUf6KJ
WtiH5FDpcK7GmbO18gEisnB9TB7V4TdGcOyguz16St9rnUr7W8Ktt1mQ7AX89rjx
oyY0/I+8JYtL1CbXgPkkqNfIkryPvaaT1htMscy0Am75u4p9N/eGDiuoWXh1FXKM
LrLaKhjjeHWqzGo9OWrBEdUOG+0rrA4or4eOqykrA2P5LdDPnfC9N+QoPmObAJcz
5W1iyqsOerk/jAIQVY+5tJkyXsKkBScGPbtmx7zP9Ng28BFfaGb8u1LXINmX+YTr
Wby9QymW3HnzL+a91sruZGdDmRk5MyuRscvW77i+LSQt6m84gwmMMq+fcQgTFbOo
nQ+/WthUWAcSlpkbFcmF4bixN3sR5ugADGM1G6mKJL/EmQjy5PNByDijHF70aV5V
65gTPW3F3xuDXWQ+1m32wD5Xqj4NAChzdLOV+SnDEX5yN+C3JP9/RLJgUFv15rY3
Cunt7xABJD3rDyaQYOjcAEwsKBh+UqP+cBv+sDeEzVB4GcCrCbr4QN49R31P8/+d
E98B8LyroGll+/jSu1ulvzlGi9D4Nnyv4VNUa9UiZm1gi4xAaTBd8YvwXYf41rft
PM9qRUULMI/N9t8axhUatgRtzChnYmKfKHPuJYxYPwRw4DpzYl18U0y2rSoupDAr
ePMA83iLARldMfgKqkbxtBjK4QEwgcIaiU4+Oh3jhFpUtThzQI6nMcpliJAIlL3h
0Fr7SjhoaB+WD2yz7d06f+hYRD4A1B7Zr8gSAqVO655y3L8pGAmkN/vyNaGO1W1q
rFZMOvidtnx2fGKMlCY0YlwzxJkUqhq9eJQ1I6hsc6EHcrylBra0C+OME1CO2LLX
Ep3bCfgKagtsuV7xFrKt20ZkgXxdp54vkkGndNsuuEJRRTHhTqab7GodIL2j2abR
hiZ2lxITL/Pp0RXnzqPyVWT63Sw6AeJZYboO8Wo86Fp3jxJd/HDdvnIfUxhg/rex
ab8u3L3Bif4Z/PnCAw4Yu2qV7qd080UEeNWvzXbsK3Fk07UQOt1Pt7WnCGPZTW80
wXQSMfCQJiezNDg7PtxYLG1LbwOKw/+Cqtz+bpDwpShmgX+ImKc2sj9WUmTvd4Xt
a4bIdTaIVN0BiVkhrEdQMZpsMmCA9zKP4ERENuC7HM0hDOs4fDs3FSPXfGoZBZWl
o/IAH5ylE70ZftYjK7L8EU2Dg14bw+FQM+dkh0vLrnsMhh9/STAAmFTxqI+GC8S2
04gwgt36ALwECxIJEjPcooVfMLxhhIcLkczmNNObYfqhnU9t+EiW2vqRc9sNjAW2
4Y6Cf7mgtPqVeHIz0FBrxsrjBbexnvODzedE5nMxMYyc3H7dfpgMWPCoBpIH5Z8E
QXqchJkICgZSY8qbT7M5h8u+bge2N34VnhjfvYzgWIC9M6twC5cgXjk1MtHakF8z
etS2JUR2XV6A21+TwMkNinngsPwk7w+VYzrGhpS++qylbidVGzDmyr0htxXQkuTS
pP2/q79bJLA4i8hbBIIpH00+mzjBq3IZ2TMA//n/0WPu0f0rRPmy6mUYDYSc7EVT
rT5YcaO9KYI7HhdW5UymrCAkhhpd/cIg4A3l9DmR2ZVKuDm85Wdv5KUrXKA/CxWA
h/2qfSGcCjCa9xPbAd4JQiuAH/RiJVNAE2ggH8eMuc1Uel/Q+wwxSfzhlMwZhgr+
jyjPjY7m05Es9YSTXSKBC/DiGjCtsIV068/e6hc+SYzKcWYpm56GMYfLoCt/jpQe
144cje10XAHyBy+ziXlxhEta9MrOnaA4DaI6xsUDwkkKsPsBa1QDdeX7LX7CnApg
Cneu20q7Jkg9heCP2sAJkP1uWCWknmAPY3JvSoTsPhMxpS8zvRAsj9vCQpT3Rizt
/o7kjXrSvCtDnFhSlJ7Vbusutvist2r5Nomf9x8aV+oRs+zUNkG/8NxqX06rqVyK
mo2dx8ddHPAPI5EMO7szf6x9cy/VnEFUbr5t0MsAMOc4B62nfx51P+6dgOnTtGpF
8DCY9cMOdQY8vvO+pdAKUf+ZX8AnPBehqlFUu9MP8lSEU8UVN9wYvjfLcaKXuNY/
aty54t5I4sKzYFq2zsSyBU0F9v0GkbIC0k/2Z+eRDOeGUTX5dBJGT8xjUre4pP2w
d57KlYq4ryuE4XmhbyzGZ/qOw1+/B6t3kUKL1F8Xnn3ezsKaQCQEbyGyd7IKN7O8
qeWSFnvVeJfBI+92aOJCQZW2OmYlW/MMMxYDBNhUVtwHttYGhecigR3lROgsdmgc
jAu11C+DlsMxRZR1sypvhFzLNFO+Ifah2uoNi/zW9dByWEbexN8xcQikLRuwv+Aj
nRPjgg9OoJC0ppwUafgvHi0LCYGr3RB6pVj6kB4Jo+ucPbdU3ZwV8O/pFawycL7j
GkF2jHyYsE9QqWZ6vj/ipetJa+Vih/7eSvOio4xqzHvSyvZUCEnXSnC+BcPcF5WX
WHvw9n23nNnPa9saggxUwzoEbeVWjofIsWY5jSOVgW0driSkEoU9s/LRSmbp50Pl
6YJoAiXxJfb5PMTtp6sN2NIukwW9HEGPSgg0PyHgmO5jz9hAy+n2n7YiICgSEbsJ
bbInuBXotBIg8x7VOZJpicsk/QyCDME8D1SoaRuOgyusJmktSNpHft3DM757sa0r
mdQgTC/IBaseOGx2V9ifJ0GrT1zD56IvwXanMJZb2u7+6h5uxO98Me/QRUhO+Nsq
cKJnt9Cj0917oXst/hRD6ZYW0P1kAckVbiy/gY/VugSh4CF4uyu9eQ9fgB47wk5t
1HRTQmPIWzTUMaX0czffrh0Azcgs7U2np/vNusQbyUTHhdc3zGtSJHbl/hC9iEK3
Ss4AlqcxAfz4au/R7jRh0G2dkkO4FxPwntVikx12eTJyIDQP9xMkRQR0CyyQeja+
HsHE7JcLQCuKt9TU0PoncT6hG5gDZs0b56KqhdT7cfSJTdjWdeJ+vUqvA037Q/6t
+c/lPrQqZpVKvUuEwzx6NoksefyW0rvyXvor69735iOLnmIriqxtDtB/X5z8OF+Z
RUmueIfy+P30MUwZsMATqdLTL7QU+HPebwR5sGexl/UHeS4RRs2U//W9Td8uFmPz
+ED1b6TSz4HSvJtn+1fH1s7xbgHAcFz16Ary8nV5h9ciueX1O/LCKRYky2a8YW2N
4diTY9P5gH/0ia8UoFgydOOoV5fNAGvjIMPscCUo5K7TCpPk680v1ZnIkEWREQVV
TSMatnXetcObglzU7mMS1RpB61yWwcx3ZF9ueAuh8hJA1LwevlFEIZhZv1WA3Tip
avA2YPhiAE4s0TtO742jz/t02ibc7pJ8yo5/LsyY0IdDHF8ac5mjE0ag/gu3riXD
2GLTjH5hgQJ2IIxvYx+GGggkIwtWutolPv4IUPB7NKap7kXK1TijYAeP43ZQkELr
y3LT5/cPKPgcFrWGM2ExuNyOfeQ99uhejkExJdiAlwC8mgq2oyxCrkVfTLnlNNCB
Xp6cOzw8P0hggOrpdB47qtBNjvaYCQzc41Zxy8rtaS/nLuhCZ3ENWE1C8qvlgQJg
2qa+6oPURaGdaDw0YaiiyAzBMFaOWU2K341wLtwQ5oajGF2aZNValo5k5Kd0jmpz
QS9CWsA7Dzgud7j5KV3YnSlihiPa+vdAUoY0dwF0Hc/SCrI3P/134L9EL7RMW8Nj
yVU2QGeoNgfay7ULh0ccc8nOJw08kCBlgvnpjzKB4/65p3LmW0GJ4aEtc8DWgjd+
b6txEvIkCG9qlrtPv4LBV06cRY/xsv0Olyrr3v51ZZ2Cz4TLWjo7GHV8OaRDUvie
FMXBCJOy+pMnpb38NVKGXkiw4/PahOUJJQzov/sp3Nk7+8lmoSrlGyeUe4CAN0nz
2Pe51qLrdkmx6xN9qosi9s223CMlY8XYhNjRFYxf7LA8KB94uaAKdTm4n2i1aDkG
BPgDbEVmD8HU3Os/SzBpUXaV6u32bBHgJq5i3iVePk4XQsgOjX8OAgERWia4AnAA
2ftjekg/YYhKEan/a+2ExGjOXD5p29nvGr8EMsWOTGWgeIMFWSCzBnhFDUBFvXk+
xzy298kUkDIF1P+DY3AMFcuqWX72B2htZJLQTAKSjUa5KOxPmJGVOW/YshLPmyLZ
DETl7cMyDR0wLwsttUVBhr6ywmn+zGJhrJITQltSq57NqSyCS58TG9SEp+uJo+Lp
+2njeUVlaHiBwNRyjE2a+7cOCaOAskeXOQ+XUwRC0beSF6eLrYwKmNVk11tffv54
gR/lePQf11NJlt0EhjoO5GU6dR3mMUJGoqhMLKhuSLvbGL2s3CV7OVzJfaIlcXCE
7jDtTqMT0aTuUYDMOrPm7eh0xF+3XceaMbyldoZdbOAx5fDmLr0p+91RUCHDD8kR
QkVuVBOAe23pkSoeXxwWG6xnf5W6VyMyK4eMVhGKUdOWv+vfmePd4hyJXGuZto8R
HayZwty2q4EsPXSwOAnaHIoI7/QHidYFLmL+V62RFregV0zA3bZssctEYks6rdrT
QP8nj+hIM150dmpPRlxdIJTEhvo18H+2cIkM9hfC9LL2R3CFyAGKCTytPSQW9H67
SYwfBp3tgMbryTVEt55sk5W/0gHR97idUPs73sANtDczIg1Cj4upJaY9IEJKjdzF
X6Um44ZAcaJxjLnrnKUHYdA3SUAcqxP4v0CIdFxxlgrNme5KOb/ZeAl3s2y7wieI
QR5jSac3JXdnGc4iTX80y/swKgnNpQABjdX87/xMh2aAY82zMTLW2LQd8WQEDlqv
gjSOURm5b0czx+JthkLeTPz8Q/xChrOyAyAgysaXUWjanwE7+Qu+bl0SIzYjWyCa
FO8kzSIGCJc1FBsg/WzE/JdedLRPWNr01FRnV7PzCtyHxWDKfprSEm490AHG5PIW
xCd+cAk2cTwUZ7Tff7j8N1HIL4Bl6SQMr4h9EzbSZlWxN8mPf3Rgl8UmkKr4GwQt
fCIPIQDCSBD8VcJbFcGQjH+sbGCmUVGv53Wq1vzAoqZi+CyOJ4R4LN9KJb1DPW60
ErlQ3V+H7Rcu0EWJWfi5RH7XZfvR+WtiPzsV90A8HxyINAX9jtK1B8IVdZbg1jg4
gGSLrbX8jYkH4BshdRzK6rHr9Ihzlv4KdgevkOUukzLPjwbx7xC4IQGP1OikOKjf
zP3R1Euk2lUkug9D9OxqplBhVIUen5fH7ZYC3edoSMK9CD0wlNr6wgNrzUTVfCpl
ymtDUMsWpU/i4HfdfgswK7khzNkuWsEOq+KRCs59wZvNZQmxWbk6DTrDQdjbdau9
IIAT5VoRoyhYqvsutxAB2QKqLaKCkj/P6MUKTDkO2DXZ75x7bk6IIKvPUAWnGaVv
/VE+m6eurvFz2qK0WTRUxx8E3C/YIwllDXcAD3dP4BtKktiQEV4g9tTIUNu7D9PP
UIFZEPPVogvAO4gM30j/ep+R+PDz8/6pYgZJ8dlt4RfqVcfpCIu/XrAIRtdLsRix
7cYipqyNENmKmtX1UoyXOL0tfeTvXQXb3Vvp0sdQp+AigRb8loDZ8AJ5TRxlRoOk
zotG03TN3lpVlNyn+4JsmIZaMkfdCshSI48n+74PMLa/fafNFQk3au+iI9Me3N4X
AlAVazxOmZywgbaXwYRNKZmxFzej1TnVgFQ+2yuAIqXGIzjObGQeo3xAv78BkWTp
S8yJzpnZw5ZJxpl4OUltxUjHZtmXeNHN0LMOgD+PLE0+GUgd8YMCqriJDCE0FINz
/PnxHgGyjiwqopMVfR6vCO+lPasmhJUDCOEJ8C33UBJTZcB7GAzB0O6D7RQyecWq
M4mZMaCEzS0SfRQs0v+WtwYSNmdpwN332qD2uqF7H8yvjKzl0Njt/kvYSbgK1B/8
flfO5e4fGNuvnQ9cut7yo5aOSnK9KBQVWzSm7qfhgTemu0FNYVBdyMn9+2X5UgiB
g8ZbW+/q+UgnFkUUtPu0dVXE4azeR8Q4SsDcJR0C6CKc4SgcinUyjPOh9Ebe31Fq
yRy/6H8nmFoor5G/BEgYmrN0e5qzMK5MibrKNbN3N7TLpJ6ERGANcIbFmiUpc0kQ
GXIF5HorsCzfZYICp3hi9R9KtYyxivGN/g2rw2R+elM5H1fpNsuuRBvPW9tgatsK
hNguwpVVygLY1ep3p0d7L9KtB/3ysK0oHPcUH6NQO029CRs2OUwmE2biww0Z7h1h
j1eoKsZsiuu8TvY5SnZ6rOG+BvkJGu/xv6z/lw1yync6Mz0lN3p7stfqhy43KKuR
u7a/K8AuB23Yx94wwkPNpLBXeazzZ65K2IU7JtNtF2aRgMdqJM4AGYsTS6OJmpJM
vGY2tunGU+6OdmKKCnLPRyGUnl8A6FLCijI3kEyCuuzrqb1SOm9XCxO9FJsPrKNq
a3OrMxZ7Ej3wPMJAP84xIStW05AR7ubki0kompgInENmV3BhDlitFkN9oPEC63bj
d1Sb44hAsXEJSFI3Wsu42KfBgmwLRBbMnIXh7imPfH0bWIAKp9kSds/4z5r1Prku
iEXTptzKPo4fDVgJ7tmEHHwKttjUpBszw4407ETdeUEgp8ef8Pcm/PCMSrg6B/MK
+teUz04Nw+Ql90f2NG9yCkJ0Uqg+LIiPJRBCRCMMucWo5ABpH47ZYLzCB6vzHaOg
ML+cd6YhuQM5Y11hncWRA/bLQ6V7cpQ9nZod5pifE3WXARG+xubSZoRb8wxjXRo1
YpUXzcmDDKnys64PDB1xUbQAZjTsHQPQX2R2OrJq4Tfzlr7muU32c315mvDpTSb+
wNBEXTwovQeoCPE1vl7gaj0RofMxG9ZsHBjUqPFYHUzA0IIlCp/5xgtWnEWAEkWm
ofrYHU8jh47BsDwvMVuJUOGvJpk/5kkIduL7iJoroT6m2z95Ipe5V9dK2V/1SfCa
bfRXSR1xB0OqLTozi+rmAnRgVtqCU93LXo2Imk7G04dNcnuvoL5zIrc8o7fCbWEl
05YRTty1jJ4f7xyJ73Zs7j87RqdVeb7EytFGa/g1mm283CCEiS6D6nZCmXQ80epl
Y8i3gvC8mTSj7zz0pIW+biCjvSAiUk3pk+i7Sot/nBcSmBo7eLSj6FzL4VbI3xBK
ACGfNV2xvAa3fNhi7CR5JQp5aya14yBcCOkVE55uEwNmuMvz/JVWf1UQkDK4AXLD
wVlzmw0bnkqoVtLn5Tzl8yMFvXS1VlMIIBcqKMjPqS+yO5d0iX43254cJ8eDV+Vu
h1cN+4PMeJovULlOfDFjL/7q2P+KTfOhGAWyDbm+yQN4nEcyB12jZVSqLDPVJhDN
FvOWznUlgIjq12gsQsnOf5YP0+hJZX1JnoZuo1yj+IhNDl9dJPUVqQ3dC1pL7xox
zhFE+9y+8P2IdCFLP/ypbfK+l05xkQXfyspj73RfaYLOW+yY7OWIoovhLEWBabcH
Q8Ecke6IjATDKQG/btjcINLrGFvvTuMTD0sUgXEGLg+kvwjOIuQ+WDxEG9zDYzJb
CoKSa6n9WmmrkL9avu8ZPNo1wDG8pHp/371vOIsX81sVLqGJHALrcvoly6LIIPII
QT4fOSPqjKFDJ7NFE8n4SE8lLAElAa/z7H6rpjUhzgWpjS/3zaHU+XLO5jfycL6T
4+4l/fsqi23RVXhIKNkN7D0gYlLt2bI0t9r/CbdnHFenMXQ1RsQYMvTfxGjyRfyQ
bQNTs3BlBftp/TLIcpG/4G9YJO9Nb3/eu6W2MB4V8dNdS5RDhQjJlB5BRrI4jUSS
cGYxzDBGl2q7RmkTbOQ8uuEB0pNTvzQgmjBlYNI/SVj5IVN/Eet2eAU3B+5uIUUq
t6rNsKBgtfht/4ae9Llm5QaF+4Wvqgy/v1pG8eZiMGJtL4bfF7x2Ka0CRjVFs6OI
PK/ojupoqkjfc8US+L3SxsbXVpG1s0Eroc9uRGQpI9Sd5mZfDAtL3wcxyd/ofA4b
wSBy5ZABuaZq+GsLJSoFf8eINw2wAMjP6mnQG6MOwDuSHiBZjqBSWjgubFV+GC03
PywCzWz8wJCADkXPXDXvhbbUOZvGnBOKMdHzG2vnmTj3gqhEoAK/me1zH7BJB12/
jfSwL/55DbS3cbppAg5jYmBYoJahOtp+5USYFcYBi6dKGMrGjyMX6eYUQiFKn1W3
yoS6bT5Js0QIuIVSV2mM0zWLw80/Oogjffv16Ejq5cR5oZnqJZ69wvYC2GxS+M5A
9l8DJ5IuQ7+eCnQPLwFIU1jedpqMb46K5zZvlsnb2hT+SUGUDYylN5JYZe/bOAYh
JrrUPyCgOK/WhGAErdboKqGz3+3zDP+5jqjABd+GySo3i3dPVYHx+OA8w+44As6V
TadeM2XMToxGts7xTidc1Rs+IL/82AT0AliglUrUaOYvUvrJ0cfe85d6TSt9zYSK
D9Nvq0QoAeHnKsjyWBZxduK4ZIe199lnTS1dPxT0h2N1hnlIhVDgxqajUOXA/J3e
0bAu64mTsMI+J2891S5UT8xyjOux/uQo7GDspNa+WBpRsEYpwEl1ThL8qjl2P3Ex
y83R4edAr2TmVxigwgAB7UFCl4x3mXrgUljbsSTIPXbxRb57ZeygvpkhuULxNfRN
Inqlfzizie7/sWYWYAbvjGXbcsHoW9EpEaH6CnQCCTnglrC8Oy0VFsL7GA/QZXky
UMDT4r1siLo7GOXwjSiPS19bydprqnR09fVkESLm8ZSG/PGLWzkTiN9/R9sZVX5W
IS2djLFODMGOh2vPR83nAqq2PBEcJIQxzlOFrF+QpNOyMPtsftMy9c4u85d6xza5
4Xs1cm7B+DF7rJh6XqeUIB/tHwrQxGk2JUYrpPRTrMZp8NF3mVJJxLdzbagxKv5m
PvRdqoGlC1zWHybFueDbhv/J++ft3CnKMI0Lmoi4pqeyNnZcdN9HXfoP46TEHCr4
dgTPago2j6V45glF9AlHy3fcfd12oqCgFGpnLqcp3zG2+N6svhyVdFK7uBWuTQYo
G/lJRVGzrbjcd47ZSsHNzVK/F4lr8HpuYxOg/P0YCU+TeZmTnCgZeNC/1vX2HkTN
0Os5XjfNkUqU7WFp36/S4r1mi9vULM95tnddnA70/PosbhvDpaqzQb/x1/ogk1QT
i/nUjJO93m/T2vrPc5gg5v8skRpGrEbntxVuq43eNXiMzlHE3VhM5QTz0KgNIuHX
CenW9Z1ARzHnaXkH/adGwHOQmLgGaJGpoJGrBHETEaA06sGF+ymytVYAS+QTfBaD
tC43s6boyLv+ALoS2HXMH+MlLw3fjsGMPvpPL4X535QVMFeKWJZC9VIqkT1ui1ul
Yk1ScDwrTcp7/w8joj1IzHf1EpPv0gBpu9pnKMqQ4ruD39m8uay+Vl4Z4pO/yfdE
TrHIMPnC+M6q+SqmRjpZh1MZdaBw0QpydQA8OvhOFlSBBVZIikSMIcqf0gwqd4IV
OtBqJXlzMYHm0RHmspEVmImoGGuhQJBqzBYfQkFHFLtgh7F/hv3vuB5JBQO3WkOC
I7GfWRr11pSpJoFEniBAfjuPdJEvCMPusOZgzcsmhf3pD2CLhT83QkxaYRNhaPQh
8M7+0MX1bIB7xMMnPrks0sRfE6FZUJsYsY9J3AHPLhjqWs60+4RgIzf4a5pgujtu
eB7Cn1ybt7g/Lf5NkoNvMyUbEw4zaqawBfqMRHcgtHQwB8Ybn08ukMXVFEeUpIp/
8lmECuM+YCOIKdsEy87xnQiaQT0QH6GxMxtVKOfZnimkzFV9XjOrKNmkNvsdybS0
iyEdK4ga4VzFOAbQszp++GYD2UIPwXJhQhje/hdJ5zDY7b3JMlOzKnuvYqZ7A47i
Dvk6T5xBbAyoohakmoyxglpi+pOwPlRxFp1ADTLm+9GPOyVmXTJX6sE7QYRbCJvu
b1J9rwbMPD7bQTViTRx/yhUncGV46pnrY4qhRU1kqDqxDwdn039V2f2k8rBn7T7S
hVh1gY7QVGUk85MvoZ1W+90kaWaxrBppRMBIPJTjgpKntzHdlXqph3pzFELJMQ8h
XakY0ZwPANfx1IVk7OJ8audxHAJsfNLMsNLwEfvFrRbHnV5Y8Cra31hOo9v3NYyP
AqzhSJICCR3QIS/fDUr/9/GFXRvJKP4hkMWw1dMM615xGUKD6kCKvu9E1rBJNrmn
exszEAQOwqXhUYeGx9mOpiTykMFPufjWbhNuyXzOCF+fMOSmJLXDEsHMtpFNZD55
02cfYwmPQ72l0GKp3yOw2IAK/OCn5seEKfoMFyHoBTKAauq1iDp24Fgc1QaIfYAU
YN0VebXEOxt9bBKizAUk/FTi4wE1NmadA43TtlMl3mVfQMLZGE3cSTzcV0G8TuVd
MZT/HBti/TW7QA+ZNBoSlvYPRIDLsut8oVknvac8WfpvV7cCB16x8Rn1Vz9qASuP
ljJyJVgbrsMdNzvE4nWL2qgP95/EvSthYe1wgpf3Uom8/0E1tzoqt88OyEmonTeq
DOVMAN5AOONSPkwCmHKDdLC1/scbJF5M1wcBMtI3fFneooBQsRkwQD1dyARRpQvh
qqNfHi4oeNCpFtbz3G0wppeWAhEOx7Q7M5fYX+CSDOWExPBYZGcup/CMzfgvgVmC
2Gq9zh1QOF+/gdoqYgbpshADj9ZEDWQZy05OvJiYsIGczBaCPvxKc769ryfTKap7
nBDtqTE6Fl4Rritt/m5J/pbbIJvAGflfEIdNtVANMd6CAJEAf9KUu9QXDpNJ8ScE
YltOqyeOEdl7YspjK54hT263giKu5GOHIKlMHkLW7ePHIiRfsteYOkgtM7hdZ/3N
T3eLynv2VQo1giCe+rLEygrSnsXIvGK+OL7HKl/wCLBZGTM0howqbxN+6fzHaH1i
wpm5vpS5zE+DCFZ6ACXmgh/f36TZFxv/4t73kwcgPchl1HNL3ahtFaOAbKEGswj+
OKfRscPcdEBJtu60QV3QUW6grelzJK0LJqBU7Lw4caMQJvW1pGLiR7yz5oHQu+KF
nuKBQOdepcNFmS17eeEmqD4tjBiEIiKANkSK1XUOFzNTdCbrSrVHaMuisrtoDcUG
MlvwwncZvKHfALXsF5/d/TkRqA28Z7xgH4xTJpNlMtb+FOUKZAMqPCPPB6qTfI/Q
y64vFZ9yAD/UuaVTCnWJJAXI7142zr0TomfREl7toDRYayGiRfHUM2av7TIsexsp
K+zV0lgoUsq7WgDUWaAdPNbk5/AE0OVMY+cVbqTOTPw4CWTPbhtwge3sGq7XMh9x
B7nL3sTDCmpgH4L1pXm2ikUupAfz8lVJPqiO2r8uXyFW1KcMU4neZ8Iv7g9Cwms0
fW4frnKYZgDl5ePSNHd3uwuFEC8BmC0ers/R5PVilA9XlXKN0/f3GanKxq2k60X9
23p/a5jf9RNR3f6YtZO1FjSVmOrD8072Aj4aJQO8hePlmrrk0PCCB8PCFejgSKd/
Bp4JbPyyY3bTV0eOc+t7dCqLuN0h5sFbitQ+nFIGnQUQu+PXMqezktTiaYv8TE9P
7KIBMdxlOLb05CNX2AonuyHnYHR+zxTi8+Yo4EZxRehwM+zYlnR9OC/3/b0ovFLT
e/fsCa3nHjIfnrgxDma27MVvULEGI6ILWjr5bO082lYdpV7Fdw7JwYKwV0qFWIGg
oSuOTXezmFoAo3MaY229ZlpOQKMaDI7Eaezht5RXJgxH7sszssXRTnM97nCAQ3zz
8iA0FtEV9zizCblyCJ0b8Jxp8iRkUPRpASIKVP5VOUcLqNw5DRWUs8DSZSlpfb1u
YvEjZ40GgFgshPe5gnySyu1MNPTfekwsKLIYrQ1EAdZZJ0FIQ5PatTNDYOCeJn4B
5VMKX/nhJk1AULecL2oZHirVBNnDRHxnXcFoOk7f4sxEav+1MQlUUuu+HP66Vbt+
OCvU7pqJ8gutr+PpDYY9ydSvfR50DzIwR5vfGxNzRdjZ2CH6iTVafp45UFGTNWNq
KhB0ls5ChpIK47PBYeU4PuJd1ugFPm7OVgq/F5iscduViZ1177MOXtnqaF3HKJFR
LdJVLNdga7jpuQQl8unaeQiB53tV0oRg4FgELldiuyU1vXH269y+kvystAMKWBB2
okmwbgqlVxjI/uG/PleIgrnMGkRxE2kmLNNlXsdIYy5he64kO6fLhXqiZbCD/E7Q
vxOPE3l0lsFGsNErOGytExJxqpZTSVURZGAn5dRov4z9DrVl0GpG43HAarlBwmNZ
vkGbmbe4MJSKYubhvqgbKgkkBKvqsD8VbSg9P7+MVQry249Ob4p5zDICBvq/3epj
pj175GVr8aUpdFxINBZikc+UmBuLhGhB3J43XOJqFiWHRv3PU4l9ik0uhKxYhP2L
iSPBdUXtnkEmvoknvzooYDgZB7JgcE/I3bvQaMa4UD4squ0THa6XftR6OUKogSol
T29tTkvIOykamhqI1FjFJB6RJ/dKwtZhiI1vR0UyNZbWH5+aXWrGNZodG4sW9Rpl
I+Q8U2yD7y6KIDBootfIfgIlRc3ucNeuDA2xg2VvpjN5LEOpj0KgUkO6SngOj5rN
QEB+kE8TmbnZPFXcmcwhU66VqdOoD5DJh9Vaa4HmuqpIEt591JAbOo+rIOILBcYh
al2Hgmr+wV3TDDZTchJW94u+Je9bvsLDesJ5A7SUQeVPGmkGH/7Ja92jI3mLT6wt
JVpKePJIEski9qKh1fjg0LORcE/Fz8W874two//iHeuRkdGOlMzTZBbf4NiImc9I
x/LJg9rWAz2EJEaSQEAjgMt9cj+RuRH79qR14rjwsRZDhj2Dzso6+OsgjacZISPd
qZ/R94s6sJMZnHvqpFdwRSdFj+J8YILjPCrZNqzk3yfkWRG2sbMUkO8XqGqrrecl
UvBcAGeLWNEaGwys9NHcyLmZfl9/gj+3GfAfJlG7PvssUZ4FHUq+dKpKGkVoLIN9
f3JaM4FTifzsECwEYbP18ZlsqkfTebaAZdJ4r/1k4YCy+y0UQ/NJY+0lfnWnWart
0hp89exMb65g7oZOH720AJfrjGXxRRZuNDvapqgPrd5qcF73eUbflC7FIFE2UOqL
7V+v9CUe+Ggssys0ioKCeg2Uqv592GZ6Sn/nQRlmUZV9fnR3ItOx7uXNzl5SlZuC
+ib74BOpvYrMhFMZsYWEgZGRHJp6hChArH9RtBzaMk7sE7p6H3eel6sigDubjCnX
QDPRqYOCbxlR/b9ZXCe4CZ8IFYsBSj7YP88HI0E7eq3tok2evDU7t6RjOwPQxNqN
+5Yoagq0Dwn6xNHWENIepIVBrxEq/k8QMegbMYGR8MMm6HsmOhOqrYV1uRNvGE39
kVlNd4AvEqRuJqs6vkRf32dpwNaswrQmFkeQpOM8qtqua6uZyhb5v75mjzSH/NVH
LI2qmp1tMo0mzTG8O6PFM+p+uqEGgCoxA/MBlT5MXKnJoS66oAeBHAC+BES7Gpfl
0HauiuRykWNIC30hvY4VFWNvQSTD/DpHut6aY+umEfW76r3xG3eZJvZV51bsiRbm
545cKuufZqOABckTYrSGRHidONOqeahY8kAzoW1RVkOGEhR1mkQOlZ9HmzJVX6wI
PUHD89p7H7yLzWWUE2mm2PxN/G9FIpiteLB82jJJjmKHfucahGgb7NziNAB1FWPz
YyjFUtc7FXDiXWRqglQxtcH2u85l0kRYuSQfjxxOlBA2mYWFPlGPb3RRAKptCoTE
dRk4iO6/FZ0FGZrJBFHy0FFZPW9Xrcv/6fthV/cPkw81qR+whB8kzTVuyv6jWon/
hPeqbMhdGP+2DcSACETXQ7pO97cLyTphs2pYDQMO29QUkZpx8+LOX6cH7Lh5HtbL
ZixZ6hd1oa71KIwhb83ch4lwZ/TctaNR0dU9qNosCD15g6mrAzJ+XSqDvUWxKctQ
AB3b9+fc2zy53BJMHqA18l0j/cI48+xleAjA+JxrTP3ln/P7xwxjA8Phu5wBc1YR
pn8xQVH4kx6ydAIOOJNPRSWpn1ItEa04WmgVCsS4sGb9c+QDzZAJPky0MN+jOYMD
pQwbWfZ2eU0mDr1pGtD0uuPj9GdvTrnienTpQTvjDCnTDH6z1jvErjn34MwUowRS
lzRcQAe8M9TJyz0BKcuv69CPbnQ5Z3iDpIEPsQIwSHBpZpcy9wQ1afIDgvYtGesf
rSYfffYDw3kZk94r+oU/Hr7Vj17UCGarVNKIqKqu0rMz0NqE4Ae4eEadiLVmxF8r
D+hEZI0Jx4gaSn/puI0Y8rCuLj8HWr3tVfTQ8efgNc7TIMp5KQiIbJwsoRvsgH7r
hgMDZ2s7x1P2nvutEDexbJYDtVe4gJKJo2KtV/YdBQkr1Xyoysv0DC1twBq1lYFr
TdC6uSCgTUtFRmWicwvksad6UBQ4MTSAuJzJ6YuKaQZq8uqFIQjcr+P1tFPKVV+B
mMXfFiHVspUiwGO3X4XBaEHlrtaiqegrn6w4tX0UArxCE4eJqQqk1hptMW/+lsFw
WlbWxazmHQcPCh4/OAnZ+R2N1o62jCWuWoIpw3Frc8hh339aREj2q+nDJDGg9zVc
n+lGa6EzIWSQ1cj9tqXrHMYOigEEwRiv6ljjFN9CFuKE970UXPvQhBZ3Vj83BcJw
P4tb1hNsskr3N10JZ9EshaZbU1arRGgDuDs3tdVSUNk9z2U2mkJzvQ4HuMNFmVz8
TwLhHEd04d+Rs4vqpw9aZcTBgfP+jZx5LXBA0bhHucXE/tAAJUEUp90ARk5mXWqZ
dKu2Bof8EK+xTubnqTg2JEv+1+CCna6bA49siJ7ZPb1ugpJXGh6eVqWAKvlqiYrq
G37G5J2XXLZ7AtlKcQWIiPvIiQ/SVgeb9KQYaqNaKPXGnkI/8rkCKt73+8j5uKJc
koHSwWAQF7xHd/IIHH5LeTeyGLknIo6vsh4bUJyECCeURDZJh7UFxaAvOe9/zEKy
AJBC+jAvymxlSLtwehu9qZEiKfdAYhMg1Xerg10vy0Z+odcjWOuvCUcSFCCpb17b
C2S7S8ddwaPRwqLppR9HUUbgQpLPmTY9gvv56d723q49euZZkacu8nm9ffD89hPl
RoSuPI24ZxE70l5tl07lSmDKksufjSYy85OGEpSbZKAFSD69U53w2OGqWRX7od7y
4M4KD4bkfDLRVApFmQMrEIcohBaNMcL9yKiBM7IgmSzfx0Zrq+C7nC52X9YroOY1
c0TtBtljoZRnQlM1hl4jcYQ5DaNSLBZq5HgUTOvHYgD8+xH1loZ4frRmQKubnVBN
J7udnqMjxJYmZ75roqjL4iknQ7tWP+A3ZJT9akLcQkJV1nN6Ddd/lQGYJLaawiMR
hkqCu0vHTPjR3vPD3r/BG69fVpl9ca36952p1N7jnRwHluZp37PDMgglIChSG3y+
N2KTW0d+JQsv3YGWvx38HrONJERs6bqLorS9K1rjh3Qb54xNT04YZWXWwDkSlzu3
YwZ/5nMQJdDiCx5/WsvTMpLl92/KMgURWScG74p7LQrgt0SZEwJJgmJS757HdYq+
TVdiNfwiwMqhcQA63Xys+EiU/g8AAhS8ZwaA5Zdja2nePk5PxfrJGLwZbNfRbkiT
vcLI5v6C9ZTWEE4WL7tOcl6pa/byVQviLrnI/J9376bhza7Cxsw8JFhd8kC42+xD
IoYlt7z7/w8Cs4JzFrJ50yYhbvh49mKD8M9/Z1X37PN/B1ROBUmpBZJCX/HyWEiE
sjETR18PYWCSK4cJ3s7jHzZW6kCUcEE7uDRs7Z2Le9VVQUP696z6TMPvTGlvwkKf
52BB+D7yEdfPqkWq2hcpDjwv2YPbi9xTxP9N89jYsRmmh7mlja2XL5wt6fvnYWI5
OyiUlQaAQxopMt65UWCpgcpUeq3DnytKslHSP2VmZDwkuSnISQvCkbwMFHv/g591
Impipeuci3dM55aE3tl0wwTyF1nREwVm4fXNb1TsDPk3zO1Cj9MPZVU35Wm4ujDX
Jhlj1/7UTI/42WSwBlBEJKdC+76QPYfiphDcbWNjnPgcjrkD2T8D7+kEwPfPQsxx
gRNcgGSK8bJKbiecf2CsSXYbmQB26TIfeTsGpp+rHgoKm+r3PmPiMWHnz/mwvwuY
2nBZ2RIM38esGTnBbIIXLMqTIn4apbN9FoQ3DXt1sjEfCfjeXdfENCuDwGn1vL4X
zVToCkLGbFKOA8K+uZH2oKZPIQXFAv056/4G4FiMm33oKwZVD+w9XsUFvgwCucbW
cUdg+QUsuo4OJdlg3F11mn1Md444R33vaPjJ0E+7k40G5QyY1upBWyPu5g1JisOj
UwIOj4ZsC7c4c2NyozF/E5fR8gICblRGkd+KxhvMjEUY03QGbMlcm+MbQLafpXsb
m/EilBpwFe4/IssD7hQCzeFaLS9dW2JtFb5cLk48yqDsNzAriX2foS9fpRsvWKHu
wpiXO721d3r06ti0/NuZxFvvkpmScgfDeyF+GeG88rxKUO6NDx+65qMKRa+fM953
YreE1Emn7/11/Kh51w1UpaYnUWaoa/eafiz1N4Zdry4x2giUokRwZvO/OPPinu/V
p5FvP2l6y/Q76+fKQl2WQzc21gBnInjSr+s1202dgt84M+3UHPs+a2pann4MONMo
IdlUBBkc6A0hJUTj2upXXjwU2k4OtyZTNZK/nbQWwxphJzDB+JlSOiRv8IEF6Ycu
PifagjBy9ZhtmB+RCCOUuf4HVolhzbccNr+Z3QBOo/i8i4qEkCdxlPU+30z3ElH0
ojiK8t4Bm2DZQZXMiOSG9ICyDZ2Fj/UBlC6jtngToC5Iu8ctT80LeGjWdHjFMnPQ
7pv/XTHb7Dd74CMSPlTyi8Mi12XyEDOwA9HU8uMzocweJ3J7FGsRf2+DXsdiMHdM
vKtiMoOK+L4f/1ySd52qkkAWbVWcpp5uw3bcO6wDlKTsavILtrveYejbRYO6qxDu
gfvG3DqMeWgrVsWe0jIu0Xhao0Qq/wA61cxTjfOH1DNRqaQ7lZlz6GflXoqU4859
MxQm1HK3HNzjAeX6n4duVnkS4dhrKegFRCSEKFkEIw3APZpFjaXoIFDK2VxcjtnV
DRqNLLsN5vSZR4PQJpE3hGZeN9Ms4kK8WHVZDWtLDnku90NxXofAFWetwD5D4IDB
qxTjICMvs39a/f2UUs7tsRig39q6pKohAdFx9o6pVmkDVUPR4dO07t5a7umI7Fiu
5fohgpJ45dwGSNY8idfa9e1s8A0UHDtWy2kCSRz0TJ2sFb6hq1pTe7fyZCDA75lS
FwFlOdgDQ87K0s2YHwTQvn4NxVYPNeKGpVZQKXDsJoomIQ0YtSUAFOBCixWjjNC2
x4R8b7JjHi5GaGQ/mAqnUvlAp4T1uy5uc4gU1daWql2XLOioeRYN9FXAI4t6jaax
CxyqA/byOgygd2uWv9diP6+uwFY8HPU2aPsJMhRilKL/bew5SvAxHbh6hxZqPqqy
7Do5co0HSzJSeU2gz2c6lloHJ4qUHgko0if0ICaHUBPpC97FX8cjHBauuoTgA1cB
68zHiVLHhTokJCb1SBdXtV0eIRnr0jg96sL7hsNCfO1U70AGhsSTlSD5EmVLqryt
pIjjd7j0hI9tR7WpMfhfgx0kPbW3gkn8tyauPS8GLr6Ktt2inKBoMEujyruo8gY+
1VfC6weSl6Iy6YPcMOxBQX2F29X0+8Jmj4OdsgyHFs+BhzFIbmnbfjcZgE+V0zoH
ucHjZWvGgIKODYfCFa6HEebYHkdtvodlFdZ1tVrUGVQfpRllnO0TvaOtfFZNAT8J
o/d1HA2qsWZscPUlAtXs2RKqEVwe64pdQxbKK4I5peioXYc9DDRHJVP3Cy4yq60c
5NEdBmZK5+QuPNeChFgpJPcZzEDmZ8U2Z9zbSWTxeoluV1anJPGNwLSE+5UvP+Fy
0O440ZO9en9A/HfMbKnt2hloh7XbCjJNPuBC7ha7hjc/qW0/eYqWdw5lyStN5ZgO
Bz/mOA8Lt0fn1joehJKGdeSASA10gda9eyKKDT4hao0ULKLgRM+NAgRh0lHJu11q
SnEIsHcFr/sNCXB4WFzWTPtiQkO3VarXeADIc94m2gbOU3RH2gF5C5E4omo5xqi9
qRVW/2B1Iubp760Ip/QrsA0nXtJ40phvE+xSlY+cD3X6rhEGKCyBadmzRo4JPB5Z
wzfKqahnzsqMibtodIjEAk/JM4Cr4aBeVADzaou9TpYA5armRfG/8rMnMHTQxsim
aAntBNPgLTL0TQ1x1qFnIlPeooK2fMlzI98ykB2s1SVXeLWixl4YSlG/zfCNgduI
V4Xj9qyQ7s2xBUo8Shc5+eeeORE4pHPcoUcM+ZBi1G7B0bfCPSYQd9QA85N6SZAv
wVLcMUpovKCo1j5gtj9PWUdcDy/ulrPb+ljjIa31ucRySyzmjmwiYi/Y1/+PgDwo
jPbNvJgSYL465lH8pVWhwQWgo4gr0Cd9s1iUYVX8R8nCgUNV29vv0nvJT1V8qKN9
E2Hap3fk2nQke2EpTEt94tttDMaxpLJizByjQLMP5OTtQTl6h0f38IVSVv8NaXqO
AxzO1nS9zkscpjRw6e+bkGlDhsSZbUxzBlVj8j7d0ALP7qj1OrT90NRlQGKhN7jl
OYWILDH02xKT1U2jEipVpzaqRQnm3DmgUlT5ZknglM2YckcZbsVnFeQRs5nKaEx1
AJ6A0axbA7UWWOu2ENHkoPSoJ2YRW7V67HROd/c1QFBE92LVIH7IZtof8BAuaWBt
fsdReEzrd/WxBhAjGSVpQAfE4O6FpTR+eTAT9dz06CvULCyUTM+2Mhq7j1wqWQHA
lO9Hq7BZJdeFFnqP6CkwdlIQCnqSzqR36P59BIGe6MN8r88DLhCAGqpvFUjk0Dr0
55l/EX5bS6RChUrBszhXZXuTW/2CbdfALiaVJPYFEpnfxNf0S5KQThWjrqZhiLnV
Z8tk2hl0mZuvUcQj7JhOezrNFPYwnVp/KBkQ87kGlKd2Uk6AQ5ozcGDa82pPwOEn
vqnEvfouR0gaa0b7YdfnGDhi55avtWLmtFw1BSdsT0GHU6AOqVqSJFHg+E8pmJIC
7wfoBqQgv/+T/2DkTSGU4orF/Ca0KJdIzXHxb7PO5eedFXh+cbdYCwD1L62OqjB1
R0xcHPQfYROO2zskRtJlvQPPqOe8bywpz+oGHigqx2IJIurylazoi9V7mf34BoMG
KPRqy2xsbAlC02Ki3S9LzDXZW3nGQtQP+6uc22aLjEJQZMUbkjYSiPEtZgSPMaMh
LsPDYDGL4aTlhUsk7WjGFFD9AQtE3yzlmCarJ+jkdIC5aVIh64ndvcGrvzY48Qxz
Kh+Bh6qxONsWlXerS7wCm1wjwdiphaD3pZgT74jjyf0zjiiySI0RkInDJjnCIOY/
nxveyvMdKz/wTwiYTQjzqnFKqgcBXb/lv/YJgedZ77BZBAIvdnWFeiuIxBR9cdG4
PoRTIEfY92nzAHnHATyHZJp7eVa+rgEf1HyqMre+8oLZRrDdIK+8gxb7OXyCofuc
44ugEiHxkOEUjhhAmwIlwUZo+lUx5X73BB434VOaEFT4bRz2kvEAxgJZSv7rIM7z
QTqKz/dWhXqVLHhbmEvnrAadm5FwnmTs1xs28Am/DZrkKa/2KzKlnzpUqbtj83sF
WQAgn8yAyu9nqnuoYlR4MnovlFJbtY6JHvy066M1wYbt1wT0S5XIkmhK/twBvFrs
/Ximmmv+OpC6yMsfC+zgGMIJ48qQDn4M1Jv7pauNxPVXJYkVR+7TUYMC/dlHGSKT
6phRLdeIWQ6h/EGfP4fIZn/jyCccquO09ila6PcMAPN8W5GZnWG56Cwh+zts81mE
s4YqH77dBQRvOlw4WAEiXJqjLCyrXfTQ6a4A9yLFfMigoP2GoSpADDIxET6MK6+J
PMMfWZV9aQpjmSpcmEfxIFiPwfLmiTEfbH/G2N1LTehJ2M90FmM1chUocZTl7BCs
xWTXTwyVLOEx/z8hI3f/j3gByA9/0hlxwvXtgP+iCh2Zhq7dW/xjLzH9dCmnNJ89
7BGI4V//C4VC27g0OM0Lljno9B+msMSlk/j5AuwaE0c4vcSseEyzqoXhj7eeGBYx
77Fj9mVik44FXW1+08AFRq5Y3ywl8Eyqy6FabdFQdtrGMtHuj15QJUAaHuwErLNd
Re/jdAWWvK6Z5m/9Pogqj6Vm/4kKWV+hh/4TGKB1bzFJQorcus//IIU23zds5N75
6Jn/nzksK/jWLWhpZ/b5vW78CHCjyxH3NZu7mUVktwU7eOAfkWVjElGFL+94coJ0
UN6sxKdEvpuvt3lU8MfKTheicj6mk5iFIXAv5/sw85eiP23vHCaHdTovC8c+DKKq
JrB+yB/oZt2uBFTwVtEPAB62BtXHeLM818gJUjnRt1NKr5CdOLoAR173/LJuJjIa
FATuAgBrtAsm3aPEqtZUX/Gigj2CzHTcHV6aeKr1QTj5zLNHXSBsJnS5KaSO2+7l
a3VSnVyu823EEVCTuZ1nY3AQqlynFH13msED9AKAA8ep4Rhg13e0k2OIGJPg9FRt
v62wYNwDvDiUyYPwsdcVhYEaZxUmmIrAIhTOPQtOfDRPu8LBf3NufGRMDDcLnkU1
md8cciKBwNZMWZcI0oKm5A5CXsifjO5Pi0NWjLGWEVCFcKQiYV8lIOiLcA90Xvht
ECKti1aZBZg/5pDG5Cf3GiIRy0C+0Dx2RNcbZT3qUs1yHFbjZQ8RBRzNOjo5HBLJ
ZlD3SpwcaTzcp64x2sWRaprcLC5v6B8TW4ELH3Zw6vSnSr0csBBiIeas/JJXpFVz
vCaRJJhTgbJZ/0gkA7ZJt0sQYk4GdGhyrP3viwojPnX1JyAgy2qF40Li63J2IECF
86VU1Jz7z52kmnkvuLFT+XuHnZil8OjNrmuVQYMEprELyV5VFopg6y677Whq5Wgd
ZrxGAgIXjJKvDGDN8/koV+6YXtURNiuK+cZWcMIQseNRFl6bwIxRrwkVhgAaI9W0
P5UjjWbfxt4Qso6xQlr8u8FiTMqC03BE8vlx1UsD45ko0xOtbiKo6vYQrneiYR6f
YPHMuytOZiKy/CDucuLIhRw0Z+efRLol0vYh1zeCQQvqZxdcZZ9vakeSn3tdsG/Y
NbM0sFE60c8joc2d3kDONRS9Y3uvB5kmLzZXVlcSzWekUqqbpY9F8jFNzHb6Z+BD
DL7dKRjJBaHI5FqZTisC2AIBdvCI35sPU0RokF5TNkX2EfQf+dZI2sSj2EDSOkCv
QtqjPVQcSGLA0UqPvzGQQujWig36+1bVWBUOqlxscUP9Sspg1pTwTQp9gMikCH1Z
5MN4JeeK72qFIbAMAJ1WO0C6u44q0S9JtqlyWnLzpned1P+e+Yxc6cvRQm+uZjZa
xPxKAT2R3FoIenr5KsSHJnBYWo9SMoY+UdCSm04CiTLQznx5+B5GO9c1VWkOoArZ
VG4ab8aE1K+5pEUPZ0eEPkQqJPi5QmciXkL6pkEYE+WU5CAcu1GLtIiADjU4oL4h
DToSBn008ECmtJMXywmF51a/IibHuTKBygfvf3G7TMzDyC+gQkBElviO6uSGD7Dn
bX+7JCctq7HhaKcYaeM4Fh2m5ta4Kgi1OwmbXKWqFFT+yzOwzVyMY1q3ywSaedjo
OCoctJPauLFwTA9YupsVgQ+3/nqhaQ2+0n077othLPceLuy8475CYVtEXVrGBnck
+00An9/QnUoymytUGVWMTeXczVPh4oRntk7gi6iiibuXLtx48bIHukrc8dpVuWQE
MjGX9L+Vk4tXRLFb5njOK8VzG4DitO4hhSGZoHN8bVUt2kV6a1OH+pczf9YCLUxQ
FFAstTGnuLGbsMs+upsKjxA5oncjuqYk13/C8kHBXkYOdF/0U4z5UPjrJrTZGENR
2cGiSwj0YcriVBwE3pdvyd4/FDqGws374e5KAhvbd4lrGOlp9UAtYQRVMEL+ruxo
gWvrWdZgvqbYpNYxJz6zrx+RWljCxJHy1dbDn001OyoPLNmrHY0UussQxmBtJx16
UYoEUOHI7ZGjCsA89bxd8+McF7Tos2330exuj0kf6e3aAOixizcF+zBLb8n8+DmM
sMi1lE19sTgUu812wkexaFqsKTPkZbiweBVVUWk/PiXL079Hbzo02G+FxZblAQP7
BTsefIRARxV3hikzvojxwm0YhhWOcyWE5Gpt51upIBcDceSyC+zEMQSMA6Ha81jg
O8N53GxnWYyqrsB7adJW/iZJ12Tes0yxRfNJCeWSmdKSbz0TeuEBvI67wf9oo5Jw
0PQUXK+o9RL8gc+iiWD0A7Sjs2QG4uvDei3TNm3RIMAnkW/4I74cd97ecFo7VUa4
zlgMVL4NvkBOxCSQ1oQ9pXj3r7M7v8p7g3xdH9z35DQei3D5cDAmBojXMK4whdyz
rgmP5bfG/NED9CYcnEJeFcklgdlBT2RPjzTedT870Q5lSa2VRQtZVYlttWZZm8ib
uLg/4ly485Ys+ribqSTTg1IXSCHyMET+Co5firnZM/74MNw/gsT8ytLUlFYQ+Nwq
kld7OlTl1J8XvGoC4MWnr/QoYJ0RlW4A/uZlSN8DIX/QTToNUGWv9fPQDK0Tu+bJ
Qnnyu7DK8u2KU21ZA9EtQCbo8Tjtt6cbuWay5J6MGUnXC2s1rr7+DD1od+Gah12T
vdXUY6Gkiix409KrgbFG7re3yS9TjsAyjQSR7Z9nIozmfT8YFZz24cSiZENh6W1V
q/B802eZSbWMNS87VSrp74/aLkUsYUy9w7VTPXLhR2TGvmrMEXTjPtJJPj5yaTjY
Wh6daDz2gPGYpxg1ztPHoA/334D/GTimZQNq8ahp4JhGGm87YuesF/lZ+9Wpy76s
madE4exH9qS8wOnpHJOJa009+zoT+Dp1YVj0/xikHPke6HEXOIv9/uhgFE5gsufy
IizDKTbj3zWK5KbCeakFXpB3FKt36iy3p5xH5UJleDmWXuL6gCVJl9g3rrokFG3D
g287fHI4uf+WFr/iK3l1vjeExFL3STBtmY9OGyCJgmtLW1RtHNWt0fESVyX/Kz80
k0iRlWdKwKKA0nHLyRHO18nwdmeZTSOF2Ss2YfZIuXvNt7LIXbovGb1xLLD3Ut2/
h3JO7geXd5TRxs6YufI4a3EhoajRKwedkcciRgxHo0kucsakYbO86iuZF+gor5Ro
xgO6KCyCDCB3mHV6yTH3ES1xJF2+8mRE2f3lFOhOJFN5xycRnvUcNzMq1U67kOaz
IqmRcwdk9Oiygas7htp4aOcdHzv3jyfegVTAhbtJ/2dArRh9oZnUiERxL28fN740
g2pem4ArBS2AR+ocBBlDl2Z9qStLBfrWa26lFLoBjEpsQfikcl7aku7DGBvrRNlz
9c5N85vv2K9R7twd2r+hEGhRzYZUhqhJLKbmga57Bly09NXV0zR5lJrHfH5r+Rex
9JTF2xNMxbAsX/c4JHVJJjh925suEYA4Xzww1O3WWvdH2qGtTeU2/7EG91jp0H8H
vwlb3em1sotBCSZGqsUFw7QAIRNdhrf8/DjXmDXrOqHHv6So3IgoYy1uaGphB8Yt
tiVnWfZalsz64IoBMnmALTvVX+ZkULRrX9/TUk2MzTbtrjPO5Jq+gR1TZddd6Ykf
xmaUqj0nT7sDnVNr1EnwwzYTAh1U188MeLgKpm63DwnMnVP+LohPsudiXRjY8Y3W
/YiYQDHZ6hNj8t9ijvB3bSB+f+GzgUt0ET/hUdq5JDEDBqMWFgoxrmvP2X9mTzcr
yDObMLfel0mCPfiLFgmpgjC50FogmrpPBqXqTPUopDZCf4pyccCBM9hmc6EmHc9O
12q1pVhidn7J9gffJvOcmSzTXkoEYahgNvRfzSQQjjzKwOqrN7wyoeWZOpfg+n0s
1wreDGEGLGGKrxrBETVJSP5wd6epaFg4KOBP3pS0AMguIpjiXt1pxA2zQVrbyrFo
ubciqg3i8/8I1iqkBW//67ZrgBcbHfPFGHYU3eOpUbyb7Zznj2GnR6dpXYhZ86Fk
9KD4wj2h5+thqQJ3PqlV619/60qpcm4MDK1/YmW1Zi/QDq4/6fXSh8z9tb5EBcYL
Rr5tXVO5FpichZgMQqRZMuR8cBY5iJubf/OPWPR+A8iyf+L3n+CMPYXJMLPVjwiT
K+IFuSHKlTgvihMsJv+VReD9GZnHwuXt/vTjDu1Lqce3urVuGqIHx8YP/+FWs8UC
0z/yg2ZSajoY9pAQ7PM5cUt1sTeC1cXjsKFqWm5GzQ4bX5nfuRDFCbhL4seadCIo
BsAF9Q3T1wRbexg3a6kFntm3irO+09m1ibpSi+jfsL/wkYXsXSsAphXnsipn+6UM
eezA0nHTZgK2N/AKZoBs2NEC23iSZeoaKHzoQwvb5Xy5/2NPkVwUdqA2UR5XZ2Li
J3WoacOkpe+8jyG4X5VPdOLtmal1ysdOvluvRToYFUv0ua0AIKS3rzjP+jkIxEEY
mHF1u+x6CuReYicBY4NLPXrD/1VEPj3h7ZJ/M3VIW6SF0HEEIz7v2xYYnhXds40z
/nPKoUd9pva3RWRwOHXTUJs08qSI23fe3IZ2IO47MVp6P8Vc4V5XQPK5IlltUTQp
Ya07VGPQ8BeZnK0x3B/ogm4Nc+Zlx9e3Fijiw8xStzmxNklNTtJsSm5hTKfk45nx
4Hn4leyR9rv+YEs0s30BWHX8MBGkQPEMpOEyKLt81ELzIx5gK9PO5cXr027fNoFp
G6TQE4fuQpZNb6AF9NI6HVypbJDmx2SSi5KM5FxZsTwcqsSDa1LQATd2o3or9q4v
SlPx7DlMEGgXUK4ttvIYs/FQPmIZw1/jfBqGJ981zw2oRHeQAHM971xCPc4TJPW8
VhyWLnS3QmGU1J6K3ag6khpEI6cJxtGuMc6yXEZN3WwCg0olrI4UsImQdsqCstGD
hM2eK/9da5XpbDlh/+a+cRKoyKTmi4+lyJhlP0YHsT9JAmQ3xaV4DwX3tJdB5BVc
88RmtHiM6HR1Llk4uRk1dKHXYz2RrU1FGvSZYZd25aFqVvIpXb3px0WSXbqpFJ31
YE211zWgaPUL5NFVp28um6haFP5hHcqa8TKBUtlwMJ6HTm++RvTQRELi3pyQFZAG
lK2QYI4LxBrS8Sy/ZXa5vQQJoZiNlrCad0q0Sx15wHKLukrjPO5p/UNSEOQUXI/T
za5SGY3F62rLw3XubHhUplNtwYxpEHxShl2tMJGtiU8fRgnxTAQxlBv5LMk9KBIH
d7FkyXgGbc9OJUR5N2n+A9xPiQHfksyTRQwVGexuN++ikcK/2nn5kv0KYpos0OPE
2ScZnKzC+qgCIP25TQqtBdAdcWMiX+MX6sf/GwAP7SI0rC6LcXAKCX5JBbeaz44L
z/vBKXpChIR4rVOq3aSeeAuHb10GqhILaUlHtQl7M5YXVsASLkKjwng/+gnRVT+a
wfFJ5ihAnDHuhc403I5p4DjfHCNpPVvX9Tz9s4z55fi0U5HE0cecOeOXRiqZXXxx
pjGfgpKx9KTriFy0GTxNUy168DGCECrqACebx7+FtTgRDD4LlcILhZrTXhl1iH+a
03PC1mPzN0wnDFvqIrw/EbZ4QNXUriXFqE9KwVhvpByQ6WKkUn7eq2g4JHMxyBqf
VtRq/5xrrC7nHck5mVBa+22uQGPU0ThcZ3eTRWb9LGZ/V7TM9cBYTLQyF111fFBn
7oi/SI/WDSbZKXSLz5eRW921np2CHlNefIguTJZUIQHUioghChXbvzwZPIcFNrRH
YYcP2DK7xwyeH08tpwHqNZhxhoTPvpgJbqAzii92KVolZZfVJXAEzTkttERbwhIq
T8HT1EaZYt3u57ZxO2UIpM/MBb2UdC438zCWin54m8H1RjAGoaojBOPu3fFAXRun
IjRc2HsMkijIlt3Ln4BmhbqJQYIpBdJ/aM5xrKqYIBbKVGogwx5LOIjUFseVkqZh
0+gdIZVG2RJ9MTMkxKy56ODorpRvcEcaLy0NwPd24JvY5ktAHJi2EdRq4hMKuVdE
0s3ot7VdXwXErJ5ZhaHeKTSAph/o9y448HfhPhI0Siqb0yY5AfD/yhLTPhhU66Fy
5fZh7N5YgtroSQb1d22e8NcutXOiAW6/WZzTnRQpR/J0XPRAA7yP61Da2FLCcTaC
W4WbcnQo0VFLxd4Zw1LetPmNVjnFvVVRuEygWDZvShw3B/b89ffpbpzcI0/z1JU0
9TBzNsPKC/T2ztw0XWtU/Q3OsyNQ1sscCHq/NFKbCaJctuCGbl91a0ySOQlt0pHB
l7GFtMKdZSUQF5QMGNr7004lcLyW/uV+LlB0aNtdHFMFfzmH9J6dxpdwfN1zBr2V
F9a/hIplgNnLxd3w0ekfiT2Xw0ON49fY2dtyIwZyXhSSznCKI7tRnHA7qWVRsOxk
qdJJ4R4XcirOTvazdHYE4MPDt+fnJVNAmhz6i9KApx6nVSlohTBhvF+dNLOt2ydP
lPfZfly1pclrAjkWCXy+ZNvBf94Afv8YdCWLIUqYU0stpsF4bni6e/V5zDM7lSeM
vaa33I+qHZ/uhy1F6yDxGVaX4W8Dw8j7oHCA4++ibGo19+RJkzw9NxFb6mT7cFfb
qgmfVSJXMPEsn1fyD2sPmo9ZFHiEaYC7uKP89KM6dOD8zw4xwM18AHWY45IUTEQd
T773lX8nJA/tmCjOosKdP/1jKkl8UkdNUeH4WsZq1d8oi/OvMVQsSVcHnAvuJkQ1
VkRCQswUlob0Y4FovUqaKlMtLWbM9HoXgcNfzw/4WHLMFh06+6PPgIbxxqbUwbXE
nYVa3j/WeqFN/0Lj7PaVJ58AfUoZ2TULytWTtyVIk5HI0/hEuRz9EyH0lF6GLmpO
gUwTHII+JXfG8gHsVzC8LpnSETVYWj02QK108rka9t41AohH/rHaFTKH42jqU1AP
5kPb2X01WZ4VDXNms8vlKQPQDujNdLTyg4WqGREAA1l68Te3+QOr2S7GUOX7vdEK
XMXTUjmvlyA/fxGMdXBVFZwqMgXydlTkMnzERwWZE4tTCfqs/4pldC/UT4UFG9+d
rBQZs6EmuXTGoJ3P1ZYbLqNqqwWg9zhPRWIH4ZYXpyGtz6OxDrGA1WqxCNhnxYaO
syk1vM0FhMRIQRGX7JTVJ48mYnOrcrMNQ8rNH13CHztBXtbWjG+b3iTD7fzKNuLE
V9d80v17pNFfPpol4G/vnpG/gOGEIBMe5vAFtEX1YG7C+LuvSV5tPhTH8XR5cNWf
P3QfBdLZfmHRm/es50CILIG8N2vSccREKsUoQq3zzd54MthuuS+6E7jB+sX65Oc0
YJLWUp4lAv9xZr9zyVRYvfCvMCmLq1YA1qdywzM9s2HhmIJdh+MRGMyLRQY6+1AJ
f1GpIBK4P/wIGRVsG2E8/bqN40jwvTgaEfNic9VODl3hvSMZcdC3gzJc/ISXJ1tu
92iPBTdSHDaWCb5pW2y3YHb/mkC8f6aVUZh+SC73huZvoQwtjqvpMAl42gIx9Vwc
v3RSccUvcYEe5U0ZRGQ7rmqIlhwcmDaepeXhXs8JeWnmlkcrsyFddUV2LEVM9jP2
EPv1GlhQ3EposEZS9MiPSvt63eiXN6k2eajIsYNMfCHlrv9ynZQ2U9jW/CCYDO/h
Jy+6hQskNxMXA570frcxlo0//B3lZeJ1eJ7PcFuD0lDOeX2g9IpLmGGLy2LvucFn
USKKc2ehybu8L7WTBB+NKeiw7++8qldyad/KDXuIABtUeF3ewFkYupYePrr07ODq
Bu/ZduB3T34QHTUnnGKhpvvtVUdI7aTk6nak79mMIwsvPJfSTaVEwATJEWHrcoYA
D+IUjV0wMINfZLHxrfP4bUQSo+ZcmL9WELFaHKVBvWEeuMb/AP94rX3ruoW9q6em
bTmg6kjvfuTbtXsJQ1lDNLbV5S1jvTXHANDEn2ODPy9Srnj87ndpHpn6v9t8WGJh
NBVF52laIxErUQikmskvso7FAOnqwHani5FqzGkrk6fh34Dsd+Uymb9DLCessW5V
ehKVYIOgVkA3ypv2oMKRdDR2B1um+K7oTBjlUtuKCeiI9Rmtzc74girVIj382QWz
z3I/AJqXq5rRF0k+ZQEguTuCdWF6m/eGF+bADe8THAd+Y4B0CAg543dVJrhc9RQx
w78xb+ueTZIG/haImeIqVHldaFjcBkoJ9RP5eyJ8EqLvhEomEEzRfNwFhK/RX94Y
PZxwpvkMdQOR7dgkEJpX0ayUmU8WdIjngP582cXgZCcrXrXZMNz9sQNQa3qup710
SVvaKZlfkLpXzq/NthrJyrSEAvOEUAnZEp9z6Q6aEGBv0O7Cs9MT1s/iQEZOK+GF
QtAhXbTlkFJiacMuMBpv+eBpvWFnreVHSbBLXoeIV90rK3lSnvIaJfYC5cHeFMvm
8RGkuMTtyJJMA5fG/R4WzKPS85ja9eDng6BF3ADXVyKm50ZXfPDosU+jJL8mlbA8
DvSx0Vc2KfPsRG91fGKMvphWG6mpE8tqKLyx8X7oq6mQ3HZFhemLKI7pua0uIG5g
PaLDb2lf9BnSmhWo1Bv/7QosdJxNJBD/fuII+FaQgKvEQF+7BsU9YDVoGb+p+1Qq
ZziIOJbc0DD3GUjIJ2gFp64FSWMafvwAURCdTrTZEIy5cViw0yqKPtufzsEXD6HO
+sjLOluL76DDjdaaAa9zab0ZK71iSzJPBzoVNR5H8Ln7IcdIRpn4T1/2/Vxs9N0E
bh0p4dz0GA+BJz71lL2lbZVcJI4E3DNWL+mOtXGyPat01m5zlA427kl8qciRbr/O
0y8BiqXXp5dgXGbCQd87dbWcx6C8Aaoxf7fVpUpfWLxufuqMriXx7RgPh7j2r3WP
4aTgb/BDUk5z5bn2pLUK/4XVXd4XyMiN2UNOhDTUXfV6BaPOEjcfbXOr+icYSacj
NjXrP8VkbKpUA4rGdMqJtyahSGQEvLNXNrQVxt9kppGVMmoenMEQFqljzhKG5XiM
lp6PoiO/hfz9dw/lqW3E7/CPRR+QYAx0gLQx6zKyovkfv8rr7P60Rrj6uVIbZyoX
9HtGOWKhD3msh7HvzG37UnierwETJl9ZHyQcPdPhyw3NU01BlCPR0CsPz/thUcHa
EClzs0ZXpSBqycjXGBuiCzZWjLkV2EJjlMmzxYVi7hvnh6BbUDf/e9u8nswDm+wq
SbpXVJVceQ2ZpvgI2d7yO2PYH6pOHLnoIKF5/YlsaB1gceXu5RbPhks+64dO/jsL
Hpk+MaMY1BEGLVrzjrsZYj07FJ1jFQhTTaopsFl7S2k50za91wOt4sob4EhiuAQs
tFjDquvOFcY7liP9m0nB00T/fIvb9j4B0t5ClrrrbSP7sgUE9ER/6rC4PbOkZWoC
O3CB0HwEF+dE8Uu4VISmUVGqLASvEuRHHFubzeZ77rk5izNHdzh9RTD8rMNn9gfM
L3yNUBGH0JOj3LxNIQlddcdHmc5cnUBp1kBA1OIDLG2r6XpGqjIAX0hfLS1qQm2o
5D9OKMUt+NZCA62r9TPxXtIBKvDT5lVn1DVBHoHZE5dwv0zpmv8hQRDYy/5J8JyJ
ORouayRojHmwkdVrLDvgax8Nt5bC0Y4pecPa3QLi/p76EE6jyZc5e1dFRkp+i2TJ
sclrSC2SJqeWBWOtzhxUyki7wbwJRvNXZZihpbuz0hRPdsRALyZ/oILfiHOj0gvY
RWAH5Jv7KQBRHyyr/yfeodCpjVTxrJWC5GImGb5tufC8wUT8Bq8D8UNFgz+i2hu6
/opPzcXScQEzYc8mZeBJ/djrLImspMSXoE1+S9PhTM5uHi/0bgnNRIsFwTNcF93k
OWr+fCQDnSiI38OwwmqFcALrrK/AC0oED8Emu1a9IlSJRo2OiqrdGsK2qle/gdeZ
Q7HH11hURA0qVcXgS8GpEI18m6HD90FtlOcEEk4CnKS6VaWrysPCMpr2W9G4Dz6l
s82yDuD9Kw3c+vmvhjTvuD5k2wkz4KckuzKS3CY73IVxYRb/3d570C5Z+/WEqfOS
EG9YNDWloCTDc56NGmqW3zwDSnYOYb1Rk2wE3r3IJWxzFiPWUFzb2qH5A88BRoS2
NziHL7UEFb6iZDiimb0cYE5zOzynTgnASbY/ZfN+njvbq5/qWAz6xhRk70hgselr
X0HreAD7IlmVvVZhwcADxGZVyDJku33uqmcuTBQlJEhpWkq9m5Ege5AYPD+iCeMn
IL9DQtg5X2/QU8CZ+pIsQzySq0Hued6rN0gNN8Bz2BTcx1/YXSYpcUUyolRqBnXw
VXRBrNHG6z61BrDERHhseO6daflOTH9cZPjWnibMv5ROtdIz/J1bCJElokcEj2E2
rOiDS2a6fXnkWYb81QaNFRc6R0xKnj/CqAZBWyaBLWJVCivbCDjAxSWgBuzU3gMA
VtXC9g/Ua6VdjQkqXYraJlSreoSd/3hlleMYXaakj1DKv5ctjHfYQzPGoy7xrF72
dIxdznayrYJWmxUhT+tk4OGcIe4c7dL6e6ISlib4BSYmrvucYbc+ierSGZx/mkK+
KDSDTIFMG01rFw4zbKHi5tZfpZgQRVvsz0c6DUrYsAj9KgSn2DZ+Z23NUJPnpnqz
aa6a78xsvZvnLKjG/CgcMOu4jwW8AAGyD/kkKDfqGfJxhwrr4uItJprQJe4FiNVt
Djjvmz9UqykVHQzCyBfqCZBINYZhZjAaKrQhy5B71TuZvkgQHMXbJ+EmWaVzsb16
IoAyawvy8n7p5IODUu7o797MGNfng11HVNpz+MmPh21/KoZGgqMhEYnDTTPg67GI
NRJtnzU9AqMQVcVE3fYtAxABeoX/FvZMUryvyj3WtoTTTjTSEhQZ++6qSwvK/Aia
Jjp/j6IbdId7n+lLEqj37gnrUYHL1f8gu96tltDhLUYePgjRBQqCibtcxKW1sL27
vvpG14NaUiEs95r/vd5Syqrt7ulu/0UoeZWcf5IQCbqPCWErnNQL9WmwnAPjLII4
K2dflajnTWWzBVOQPRCFl1K4yOqLKhpANSvH5iKecwRuY+1HvYHbYX/AkbYNi4VR
4Vpph9irenSJ4nP6Fj/kUZgAZFPyottOS3PV3ppIHN0f1JXoBRede8GTMvDxk8mT
ynywUL118bg3ECRKy5PXkCG9AWA3sepBsm3HAN/G/lFBTb0bPgHC9Rc3RbAyMUkw
K83OSgDvQvCAARu3L4r808rZVRJ2YqEciNrB/fDXpvY+k1yuNHs0YU7wep+k0njE
sSNCxyzGfwny4WZeVzNzrgeRY+IVPJ6O7HieIBzx6z742fGrwe7hZuBXbfV6JMGr
hixEY2TQ+5JuoFbi6aI8xZfmGKLZVA17nhBORXDK3wcKC2SfJe4TbPHlVL3FagBj
Lrc7nR3Qc2LSos/ylBlPmy0j1aTJuxIdVVK3Ny1FFOtz17CEefyRLinwCR3bdoFr
MVHzJW1fQRzzI59/7sNxX2tZObCaHsp2yU98u6CPtY+EXo88fHSFbYdi8tTcGBcu
+5sPd9uHQQ5LJoqJx24ElffP1zjDNk/uNd0xgR0O9su9waIqKTwxNlk7WCAVfeXw
Uj3FGM5Dp0rndhxPk4lqg9k7+5g3M02DZ79TwYRS1CYJREG+t8RNDvj/cMM6Ltnm
wWMPrB1TimBvN3I65rRcfPPzO/y9nnpYpZ/hiF9WdsBxfo29X+UVGtkC5322v8uf
pbfC7AMKFHqgmMwmvtztIsuX7pDgEjZX70SXXymJhKfvegi/VBX4DjLjrAJmo2u0
h8geFo+k1zG8u656twIP3O31RWnQYFNMGL8lNwMPPAISbd+zi4lb3KT3XMlVb0SG
S9ySqmyrFqETUBvuPxC0CqeF/t1gBtSv/pnAyTOrPka3yXulrG4giAZV2sIGG3nr
TgBv8a8OgglhX1AnLCrsfVuLyAHyD3pMTG4QGrbnX5TOcJls8apm00k6gJ9hpBV2
AbgxszGI+jUxEPO3SlUjLnuFY/+oQ8jX7qY/bo9CK4vyVJcX+7jcQtJed61GTr5s
7POL6bBPv4izBkzVj8+/bZ+VUjjdLrdn1omVJFzcM4HIcNfqoW3Po7uj/A2OycxF
Wk6POdaiLS/XlllUVNbgsMgcJR2rjuaU7QRw26+PhpjxogkDpRYzFHtALXVVwnjO
LTF3wRobRFsWL2uJLQMv+bfZWyB9qC+e88yKeLVYVRmnMWrsoy0uYbAXLkHNAhsK
r7i3RZOzpzjq67Em19l7WW/Hwo1+41TIR5l8giuwg8qRQbgyRM6lPAUhQfTn6tSv
iA19p2eor++jOB7ADiZ/A43YxYKuBOoDylI0ppSo9EZ/rPK5brvuJWLvdbMVheFs
t+HjT/3ZEVuhJtrSrMjmsn47v915r5H42YGPrdghqAOVuBnbjuLKQzozhp/2LV0b
E965bjqDgjr87eCSYY15uxySmM588hToi+6lNiUXxZYPYjVfdGoRE2V2mZYPbmxd
kmpRlXbejzUdX75I/B0cvhWHPkLw81XUPHsxUH/xdW7CeiNCa5Q6hd8pPfONP3pM
Vf+1LPY1wKk8qQwWWygybOJq5nPrXEEd4cgCVCVPxRRbJBdzH1MBKs7gZci7diwp
72abYLSz7xlsAQknshTBJXL8wL8jeIh69VUatyrbre64c9cYBsudwHmb1WYNd8Yn
dlxFr8EkxtTW4ljFM/ZY/8QDlPa1FkyYZCvXV5CZ2giVaKhC2rAOPQiAK/ng22V4
yTZ7HPaL1EHLrlYPucXL+3bnH+IZhASX8rERFMOvYSqZpkePQ/AdBFe6LPsPlsIg
JPxAGl8d0yIaorkQ8+PPU0HT8kdAM9Xrk2YWr1rvDQ95/t9wehihra+d8tvFQWMZ
Cl6K9Ew86xBB2U0I3oMPsWydj5D0tSMqHb2+Fwl1WUdgPVcWqIm8tScoIAi0YaA4
yEuDbAdcya+jAS8XBGyKatW+IhaBteMO7+CcWZMWcxyG0kM5i9QEyT1F29LIxVk4
jRPdqQN33J5ixPBRJZT2VlgcNQ4XdthJaOCb3diQdVqoLfAJ1+/DkxjU7SkdyOS0
muA7iWZvio0G/OaW4m0A87NOhLOwGFjhXlwVIOq9MP4vha63ji942cYkE6oZ2KyQ
ISBiNFK25GL9umQHcLwAsi7/m7OhYRaKj3FSh/uVAzG1kXXE49ljtlrEkCqc0A98
xAGWQho2B1pm/CV70tWjcYmD+5x+lyfqD1Va0vy4VUfzT1ZySSyopt+9vhQYPqvn
TrpR+whuySCYXtR32I6LW13RYzSIxoJaxnzuQS1VXVA8dQ2PFZggMDg1F6iiJuz9
t9ezYd0HRGImpz/kE5dq9BZoOABwvTsi7Q117Sarb72UIf0xdztSIytKhGFcIl+e
J+RLgH/rl+/g2c4Y303osB6LVD4JJcAv2u86QFg0OxLQOgn4joxUJjzR4e2zjKme
KLqTQ9681WE0pheihJTTgDJ3gXvINLkRhd0cXtfJ690QAwEl0ZMPenuXBBFYv8Tw
+SDISDOvmsf/Z0Q9gWeQcK47DMoV7Geez/GpWuDKRFKjmTC/976zHATzQa5iGR9V
PPJeJ1UuneZl1rlGRWFSnjnVO0rjY1LSbdV8cQ6+mwO43D5QW8jNUSDErwzLh9Vz
KOz9JD2DE1jyvceVPL5b/XY0J/Z2C/1T4ABLqU275B8OI2o2Xi3TGaQxz56Qzf7q
S296VHezgwfCouwsq8Uc2K3UJXbqCZFlgBXh4XurTfPGH8jzl141Q3PWL2LU0Xtq
iuQmvqj3FSlrJ0SdzijhlVBKNDiRwjc9i8BqLWi3baWVaUxOmXIN63WlkfUnJVIW
80Qsn1i+QdyRo9hKYGXSMzSwA/3hkISUabXtJHqbdfNqPML9ebST5APIesYyyKtA
H4l300xNux0hvmzNeTCzd9CilBsqA7aSpWTRz0xYU1D1VWW4vl53R9o5G3jTqbw4
y9Xdc7oxCKwWmVJ3uJJRgTUK1heCcodTYCLRY2CrgyKqUxoPQpgVfaSGEsz8vqJm
eIi/XO65Tqj7dQiSMZZGRIbUvgjWivrqH8uQApsJjPtkJGQI1jgLe+7Ic5SNtFb8
zjNSkcV5XV2IOG4Y8ALqWZ1o5PxzRFqlPew2m1WfF32FvOjog8bYJSX6xYt+WkWJ
W+CuFNB1gFobzv5dP/qtRW29Q4v9rpmgfig1z9FR8Whu9LU/PQMCAejV65DOppVL
fymi/HMLKzBfQ2N4lZbeBhGFTFzFHOMZ87ci2f0P/NzcoRhlNb7iHx5bKK2md+7V
ylGOzwgJ7hj0MBglA6r1m79XAuT706rzoHNCealGzFKPNyqjTfigqBDZeQyWfhLU
PIv0a9/qeOCXqcZF7wcWSe8YiXYpOKhkK1h7pS3FDGdHDqPvqV+imKp+bVMlqO+d
SEuUOfSjnBdYyE6vG8wPgIG9iaS8sic+shT/4IYLNGLKK/T4SA+vmRiw6jplzUDo
paPTocRm9v683+oTskMgCjmYerErGTFvKm8R558kNMuB0L9TiieQvvZPUOIhmDeo
gQgvmRfhbLIW59pBNn9DFOKVDkZCZZe2tERON1Sv/8pdipg2/KXHxI58w+BvaLpI
eipyloHObYROM/ceLbF6+iAkKQ2w+SNLsW2LSSOQ4M5iVYfqUlhcmhqNDDCBlfBL
5MfMNWAOpWxog98hllm3Q5Svjh47W7KhqJ+/GIo//3L7zRrpN9x1GfRJwdnxgFHL
I4q+WVb30A49yvD/YwNBeiC6XAk0Plq4e6lFkJuq3/1WzTq8NhEYwjQunOtm93SQ
qJzWkmU3qZ+if+I56LU+AENT/T8YgTvEJCC3UBe6MVsiTuuTCY5ZczYjsVcLLutP
vXnvpDsY+J5qfZL5kMQOTjFD9x5ycn11YbVE2907lBEStcavz7fXk/bVBky9xH1m
JjWOrfUEuR4UXXPsWq6RiA7GJx0bmHdhloBF7Q7mubhi9W15BD948THB1jP1Et2v
QqSHTsCfuCWxkpR1zo10gGaCORYKvvQWla36Ql+RcvMstHc14JvzaoKxawOBxr76
kCExehjhWyXXWRpa1ASi4KlBl0TA5qR+SJPlXwCPBOBaTCJEmlvxibWgDqqDYYvS
32JWqUdQNng3KIZ/hDBdaI/b3j5b4X6RHLd+dtAf3S24nJH96sPmBZ/oEqGbhPZW
Np0/xH162QdaFyEEEwgqYu7DS09MmEPQ7nL7NAD0J30FSpHWwOKKlTBndjVBG7ry
RDaNVg4mw9je+BDbn6N01bnlRvCM6nxMSO/spr4zsvaxLajBrN55ssVFnVUjWVs/
QgCdgCj5eYDjW+5DXngPlWlTzW+ctlkbjDoHS/epk5Gr7q0lkFSMhQmA/Vbr/J2m
K2Zdgx2kZOlMubQzRedFLUHLPubQpZCTp2dk/+KKA4OSJesx42o+Mp0fcsP92bPy
yovvI9Lyjuzb9B2IUtNWKi9ZjQM6+O8f8H7aiD6gnEg4u18hJHBucEM/j2kfYjW8
A9dhcwRE9ZVVY9/hL7mzydh1CZn0QO3A41/lxgaByI8MmwVqsTtxBMYfEbMArkk2
nDrK4Kw8ffbw7cVePUma4XZk0GqZoyIcGrI5LRbRO3UfG3Q4pzYZlSnpNyJz4xat
uNeVIMRlhauo6YrB/KpgfDyHyTR0Y+b9Fxx1tvC0gONr+S7jOHaVsXTadTsQW46F
M3i7Gcqil7L+N/yrZJ944GivN7fcoanAa+Wr30rGYEI38qR1IFnBzO0bhry3HC7F
T7pC56wNk89UM9Ar29NkDfevutwPRPgkUW1YE7TMdzqsoc/WcN2T++jnFzmCo1gd
sOY8MVQmXNqTdeBKbthUTVgp+b8y0STp65n32GbGihMTHgVRSLOLNXEQCYW8c8Df
7dv7yIu85iS6xTnd46w3EoIgaa8BbFA32oIBS1Fym3HutLF5lpiPc07Ikr1rbscs
xRgYKEhu/tvfsv9IsHPn222tKtPuKipPQc9Hm3yjRsTgkhpq/hviKV54QuBpJi7q
zqiqT24DoGi0dmYagczD8s8iYNchnoB6NkLzEQGDvR0iGBgQvDcWLjeahbfZQyIW
6o0PI+zcnqHeFR4RtuygBieEgiJL8tC/Fx6gfmJ+XODFtd91wkHMdrm4adB7LcPz
W8e75AaR28FCfJjATECwyqxLQ2xEf1g0oBisxstgLJPZZwhU+APujRlpezISnlEb
s0XYb5+T0qqO4TYvnla6+lhEVkc/SWhj6/I0tHPS/SAlmijtbc9/Nmu3DVOHoHWD
IlXul83PjC9K5/QtkSDd3RucSniNrhKszfCRETN8kACiaEbxZfUQKFU7J/+JdkOA
l3ebvhMzWLtzg4EMpQixKyM412WS5sUsF1x+P0YgxW8JTROlMwmtGGsuZn4RPZBv
62dWLQELUbsKzUnzKr4QTBFHTBt86jgVCD3c7WgKgfUXpm/PmRS2lKjlouDD48pt
HH6BF+qpYqRIyl8Zv6Vt8eu9StTgyDeD+dSUsGAuL7ayePA+rVQHn3Y08MUrCiNz
zVBAsgXFZk6SIDnNIv9SCcewdnc/dnv1OH+gDAD9i5K+Qz/nZWEtIcPF3Ev3uGIE
utdMa4shQqd9lGZjXxFlirMwkoMzaBYbFkAw5T06mAi/oLssovzXlWZJP5gXpa7z
Ia9QTE17EGStSOfBuOOka7S3zFbCusBV2xA2jnaQ3C8yvSJ3x+WJd6XxepfEFCul
ihOz+L8WQG+sQLv29VXh7xETdTZYGQc3eW+XCP1QfVzaYkKZWqtmHCwduWpLv+2R
DFWWcKqume55ObNBCT7V7rl727LtwasCq0jy+SRau6cjjnnzoDscfDLMgX/iOGBT
4C/PLQpGLaDpWUKvMmFzXDzBEp9NRHr6fFc6gn5Mxa7LWdmObwr+AANv59QVZg5B
CRPShZl5JWESo+VysKlX1lIDBgYd130NKzemybHBf/BsMZg0k2aC4NVTLk0bf9B9
GtTd+YElpRJLAbUnnUJy7Mym/ySgeQDgXhcFdfFXUELe4c9DN8QJtel7JW/mosGZ
H50ubekSgOQmXadl8/b6gNilPNDZzJWSKtps5ERLYAf0bFy0Yg/Ms8GolAxCOttI
BafbPIrMBDXimxvb2JS2U5vYcaTc/hPi9Rb5RpN3fn4VvV9Qw5yFOwqsU8x9/Ij4
YGRLzMeUBDGdoD4gsTtrYEPXRce9oYmrwea9Ub6diNESJ2yeofKwglJTRgZyGLxF
oe+9Y5dp1cC6q2H4ijp830lpNcLaCbrNg2iNxid68N45R/IcOPigBCq8Id2Mhumm
c4evEU1/Jd9NpdSr4YBraBIDu5EWyn0ofHcTGnBE263ogi2NuCxm0tXvg8hB2F72
1K3S3wN6netEd4m66AvwwysexoJa4jERMZ08oLH/500PQLEX/+yTCAU2lox+RDza
0cCM2MPdpuT3MA0TYsOAR9zf4BuOrKE8n9U5LfFibDUzk+Hv2MHvH/RcYBQycZbN
SuqcX0jUqFq2EsD+pX2IeAU5Dbrjxn40aBJaMRFPe8rZWA8yUB+MHPBo6J6LoSai
DsaEOSoDBTQvg8rfgpDHipGJ/Jo8YQ2Boi5AxW4y5zpYIB7rFhLKUQdLtjd2RAx/
j1d/HD2WjPYdB6rHtVewCLRxaSX9smXXkHBbJdqJaBhZ26olDlO2pZpLoqmzQP1+
uUayn2g6DeJW9LBxrwKbjiHaOFX/4icQ7n/3XvBw72prrqs8mWROTgh+1jDiQZmX
FlvUPxEwDcwgY64GaKQVq5+bTmzzOuCfz/lcot2j/BV4NMebiRkQZ0CrBp8mwv0/
TasGhmINy4BLZ2LTH1MjGKnAjaaaQrn5R/LHNTtJarE/MuTUqHsu+rR8MaTn+KzI
eZGAcGv3MiEFiJNBdc+GMOW6NZi9eDafzsvhZyCnNYeyN3otBtjBTn9tz1TE93Ad
XqD7PeJ8740nv8dTuvMTx4OoYQ2K40oKlTyug89lbTyKHMRohejA6X1EtIkc7sis
OUVz8V4fQD47bLINOf5j054yinrqYnG0jxjpMIiXxif5VfjLVdjuBTfoUrBnqmL9
ec69NLyZmuiYxz6u8UWGwAYadL4g1dwcGoRB92+/6HK3Jr5qcFtdPETyt3qX+3AC
mfPQgE//4V+XJGvYIZTRwRm6+c+ksKpYOcQOzCfk4GFZYODnr6y9SXYGxLUmCjE1
foX9mL/jMCEM3LYp8A837oAkPZRhW0HbiIsRbxe10GjqlqfbgCGuT2vXs3aqOGsk
3rffnM6cloj+zH4xubDExpWS/sxjzPZHzycJBhtBXXMra4xf461zscADrZj+e6ux
AsUBM2iM84LQOh/EQ1FaW7AMAvKW4ypfsUhDzEne2Uy35I81SrgJWZJOTRIpZ//z
+afCtxbGXO7Iz152DokwePEGnOyQ/f8qufkLDqhIqKEEV+/x3s19rV19FFDFbToP
Nm9GcVrdDnYqwf/c8pA8oe7WocD24thoUMawCuS/O/amHhsiEyaaFTWp4PPa6u1I
fCuid/VMelXKiB3/a2iXH68B9EawNdOMaVkLcNNs2g478IYfbp7w9t5ORupWa3z0
m02ITPoHmFKLAq28HS/loQy2jnkzAWP+Jg/T8z2x3bbY7mFAD064A7z+PMgzuq7m
yZ3PpX143HL5/0ZB2odTWYQNqL1Lkhuth8dr7rV57/51dlD2QUP02Uzy+BdVn91x
CiokQRngl06YyKG/zs8KXV7JX91YHdLDycM11tSyyLvnv8mhN8UCPbXgh80WF0K5
TCKE48Ks1aNTeA2psATgRL9cj+wcoFx1KRTlmHi5K96LbdHEz6zX0ePObUTphe8m
4W1phPssOcO2zbIOS3Fxk/KdoLajLd32ziZOSD8PlVzHVaPWaF0gmmQaocXKyP0u
YpZa7Un8cA4iiWPW8nqmnX26vc5Hou7/u2i7HBAuj3xdBhTbEM3IiVOoL9phG2Bc
zZWspYQj7tZZQiQESwP7YzAU+vw3Q5l+ytFlcvhIEFDEiU2VMw8OfUnYeHB0gHja
YBdIExXrn07gH46QU/P4/R0mHBIOmnyqYKDq0Jojbv/pMkwPb6AyaLgXaRcbpVq8
fUbh0XkgX9jiGOBTLYoEqDhTh8GsTNOEnfNqwUap0GqT1iatmUfmpxii1XoWHxL3
MBxqHm2FNLPvUlMTz33NbC+SLZLZ7z2ASziUHOw2ZpgHhNXDHKykzXHs0jlN1jzJ
R1a5pkOyTl/7zgmtC0MnI7hRf5ugM3O7OVQ0q1yd+BFyaiLBs9ky27WomACYKey/
eg3hPGiy7UmBr55Cp0VxZfBFnr3BYmVCRQnrEPEUyB21cN/cvyY6EmMmKjULmMRu
ATk935pB9iQC1AmR64d9eSSRYYAGppspAOJ53XPxiDHrzKEAqRsaYq/nS67asYrg
ZXcA8NM5YKH7NguKrvC1xia6Bn1iR3FPG2oho0sm3v7CVOzSOetzEQsb+10thoaV
egQ8dfwaZK8OeaILqjYvGGltdVOcMh2PrB5UjCpIxbEum9ghi9Vlxkh9JMQOziZk
j+BFirSmUxr6O70mtQ23oeEwMvScimtIqwSuyOvHa1h2tx6nSZV1LgA2Uc8YY9/K
p52ktDWXQ6b2A6bW7rdEEfCNb2KQ+wVOyTokCN3OgSNLe5dCfgAe7ZDBbItDhk4l
Ol/88i2siW847thSzuVLI0sUvLSY1fQQrR6X5flvYpCfYRwJ2isC0d928zzicFW5
GWaCgg/J3oXbAQaks1f6RTz9MDyca3XUozojLgbvIuATVkmdSl45DRUhkNM4w+1A
9rtJI/PW3cfOrsbL6DYkgO4kDLtuXhTXmxO2qhxfRAS/O7v+Bv8TBeu4YepmSBCD
KP78TDSSsxknRmWjk9+AHaNdr/2fYiFdbUyzm7bYzlZ11hZB1lO93ZA18Ifq0uPY
sBSAyzKVNmClQaY8mDtkCzwTiEjN8XwMVK43SZtlLT6hvII+m5D/gxNvYkUYTyNc
9jgRIiLFhIF/Q85FRU/Mmz7ay/WI7A2vOGwFzDSx6K0EdtaVnrywMkjHkoU4zwYr
ZMj+Ev3g2XwJx3jx2rt6PMyyCxuPgXQmrrglwGmQKAo4O7Bl7WyrnUQZycP54jrU
Yva3HqIblFdz1+pCn5yGDoNEXm5XTgVx0MApNJ5pGM0oH9oNasUnuKc/2MdKkIpn
5p03HJUZ7L0ps6CJyilEtXPYNtI7B3nGwpbGOKczAhDwdQ9WTs+neJzXIXgCByFG
tcBfJevlWr89QjWFuFyr8umC76fqygndgXXTbAWchpA5MROUJLnHu+H+oRWe8R3g
NS5fDTUESkICz/PzXgEB7MItmjwKHgNgyL3kFUBHwnORs77p4eLOivAnk+mOHI2o
mcXttUFlgGdMYJp+hM1YcpXanj28ZfCjugFLduiOTQMqYJjO3rTbAbUa/Iee34Sh
LSooT6XH/g9s71WaIBAuMejYmHxCVzzKDijb8yiHQ6FcPgBmkeTarnsp7HlGqcq7
J8NKqxFzQgoO6vry2gH/jLfMCfYYxZtK8tI5xNmini192sIV3odI0NJ/wVYgsUJ8
zV5q+z67+LMGfVRtIyE/bz2SE+tf4iNpDb7NO5dZd15JtLldoQsA3tbzb7OaRxr/
Abs00FN8pvzN9wiQki0cBQuQdbJnPCfc59wMEqeoiCGnV8GjgOm4xdE2BJ9M99E7
mgPQKm1X+IfSQKgzWsaVK27gHDkJJNIzcGKGA/0W+ozO3aedpvnHAVOutVncCIx0
RnVh7VsEhr2Cf3suGt+Q/bbY0dze/zatKvuKG3kMiUgC7vJiYtYrTs3teIcLSF0w
3tCZtq0iWDqyYMSNms7Rmb079TJn68eNsYR2PrIeLAl44ucywNZS+/a/0OPLWoyD
+MPOxyS2dXU+laG8qWPTkBxBFfV/7gC+d5TgB0tF+/zF/W6E8Z9zHRn7hLSWyPRS
GmvQQ+Xrfo2K13Y6JP0+iBZNl6+blA96OU/10alwybvkE865cZNUTP5Hc0esOVgr
RRA6Z+6dfW77htyFTSmyJZMyBdNQfnVlh7+VDnt5TaH+HnciAqCxCpMd7N0Nx9g4
Vt5CnAOyC2XTgxefypNjlBEgVHd9rG5GD2flblMhlNZyJB513AcFdB+M2KzsOla3
rYJoezibk2UlQzBkE6Ly5wlLb5sWlTe6An0CxFofpcU9L+ppXycSUGJ2OXfOL+05
jfiQmh9foZdvQ3xh9XxZ+TdHK2SDdjHDy1xet9iOrP/B+HkcnpBPdTuy/tiAxjss
cirRaaMnrxa7o9kGBtELKhMqYiOz97cffa9lqYYKC/6n0AyWRIa/0/LsbOMXlbTt
BqERbKy0CXB8EhbNdMJWYVRI6ZzU+e8CegLYwhNmqB7sEK/cAlfdKfytXxlLEsPi
UxzGXYloASTr6kdylFGIWO7Y1C8WWw5bJA3o7HCZzMjI/1TaRa0iUwbl93E2WKgV
+fzQXJyCryY5zcv9NWORplqL0YUW/yWWf81Cuk256pE+yj/hEbDhAfxqQCDdJBMN
yQBo5jUsMtSwCxuC5PiUZXdtw/pKaG9wwzzsv9w1kxx5nb9Mo9yfZXctNeFNPDcf
qA4SEmoAsX1MXbkfVc9cld0OlCIwu8GoLq+9X7+4xEn3laSvFk0rTnnPXHF9Kce3
6182fC5OWczZieViZ6hTovUgZKq68Y6mbZWmHNr9xA3h8XpO08IDIA47wrOd3ik1
q/Kzxqs+p+17WaLkbjePW+/uXjbllqMSnkJbKCbwj7wBNsMCUKvTlwk4xc6nfA+z
JkZ8Bv7VF2BnlEMCI9gWbO8QEPtBIGFRZWPw8NXO5My/jEJQmqUF9V96jfZEYL1p
gTihoGyeMpoJ203BP8g/9cFBlGZFbQISuTMRLHah2srnPnZ3B88tCKAlMmrqSJEL
Q+6JH6dh4amLsiV6JHUyo/6SiJPvsG34U+rEXI3vuLaY9qUC/rWf7NzWb1e5xk+w
IWTD20OtB8AunLBtmytH1bIpZENXI3lz7xVZh7Fxa1n0EImQRH/QfcohF2Ovfdqc
RRoXs1u1G90Gzqnx9D9+US5qTClWTTPX5yEFGsO/I8RGpeNVudpzNzDDyx1yFGq3
rqHoRgbh+UKeZ88Q8+dY9UYYRPNY+9R8oiBvCtYUaAVUwy4vyRWFtGBU7F1a3Ps0
WBNPTTkpHfAW5cEU+9bkgwbG1plqNrOBlf9ZZdXUHAcapKS2LD8qDmCwyLPIh+GX
FrQlBoqDWF9Nn3owqCIcMo5JNmSbvrs2l99NXOpAlv07fG16wHIZEv5LXgDQq8sY
76q776+l4EsSFbsDQKF+3C6igvXNUowoRu3wqBVX4J663mXFUAb2RLvW2PH5DC+F
D6Eo2rcBf5skI2YmgHCgIRETYshEhOfcM9Dcqek03cl8u1FVu4eYbRTJ9ZieySmy
XcRG/dKTcWNkdWGeKfZeOj5i2/0sNGVvOUm+lU9V/8gDHcHOlDAHlnjeWCDiwJBC
VkGObh0mAMJMH/vcN4uBcFwUtINjcvNX1D3Ynlq5xxDUukLuR/WbOQhSILNsousg
xCjN8QsXcxBcKVry6K5YFi6w+JoQgU1U7yS8Ut79RxRApC/Bbi72NnhxQ2Dljdgs
Nigws8d59oKrNExjvWBWSCUipUjm3ijE8ZDiBxYgtmHtdqGUoniSULWqO07a0zim
jumA4eodIN/+d+fnegflPQF5VPk1bYB/DUVEpwiCXewOTfj1Biuy6Swyikx/7lMO
uefoi5/4vnOkgfqCGtmD8qchtaMTqiOkgn1SBpn51WxL8N8v5X5WfcGr5v8GHgBd
3nz0C6HdKPDtqDIiFubfFC4Q1PmgO9Sgw/XsxhtSwSxRabt3It0vFZKV21WfU4YS
4yRafrZa9SyYgTPfbAdKcv+jxWtfjXZwTSgplUmrT6yUeMoMgKGEH5itUi6aV/pH
Oxiv8PpoBgle9WIbeimuN+DDmdJ8L7hIlSJ1ZO3qj+2Olh1jxQ49swHLIYlsgfjN
4RhyX69TXxPNy4HeYDwMCBEQm37mBFn0KGrec/UkUM4gnuR35RpoybTNiRe81RHT
g71twtozS1gEuVxKMxLGy85q+Jqxv8xwZXKLJYVd8gIvx2FlLaPWk5piP3BFgsok
mImspjQH1yl67vdvnSq2WZgg9TOtWZrKli/Cy0LFZlmV75HwqeXU4W3RV3JIxUUr
P6mr7K5Yp9AAr1yy4Ta7aX664xsclM6Y15PG83KMGHoH1D9PU8Okivt45qaYVaGS
SdpNfYhDWtzq38PeMqYbc6m3wfOD42BBo+Ch+wUyWNyxM7lC7tPBhY9ucOtl895W
Q+kxx0D+z+U6hhYIndYfSUNRpZTTOlW24/XMnq6FatOAtQngTwZu1HP/F8Flq9mr
S6q6e2oc/BQWB5V4ytGB09T8V2Vuk76EPNT35kAyuUNCtblm7E+hMcdWQZ/DE1cz
N5l8x7zA51fpRiouBkghrU9BsFziek2LlaTYDV8jHm7h/iJLQjWg76uAptlIFI22
zGiDV8+RyQduMCrq6GsafGG2V/4UXdloRwr0Hx5G8S26/9bEZwvZRVcg+ovon9ci
W4HDL9emm/tzRBun19NGUPuV0+pat2eTpMt4k9os7uQ3rVpnvNwuvNX2TOAUEVfD
J1ajo/qhlLzWn+eXCS8UuAdXnma0QDyc9I6vrUNiOQZ2CuwDjYdS7RG52tiikeye
G03GwDNZc94IAgSaLNVbYtzb5uRmag1ADjW/i8mOoy2gnTgi+Ace+nR73BRX2c6e
RxIF0qAY8S42ElOVEObKOpKrBxrfgykZKe+yoKcx8qPvVv+70QuAXExJC/460w2Q
YvXk0vDgAs6i8NqOVDFiEw4x9wj+1AzrL5Iegxgn7d38ToCsuBXkhY8u4jqtgVcv
AcQApi4LXwW/jtXVT7vWaDKz4gjb64xARsFOt3jEg5yduAQFU6lWRG+g7oN++lzL
4zKREHRyMolJ/vd9lbGu4ixJtjZH5B+RBkG5hmT3BW087aKTqYi+iATmhpI+64Mh
pnHp+PEFM0OiAjiobRunRzaLwUlD0LFTYDL36Uz7cM3O5A8vQzegjSsvB1S7uBT0
G8w98Xua0doohqZSLwY8V7bUyUiwozs1+Bbb9/JVJvpO00AzkB/yOYSeQIP7zlmw
wIma7J3L1XQhWVQrNosWhnYjWeDkfwLwhzk2Lv2vvdpd80rsoKcB3hNcX1ilTGbE
/yZZsuRbS75ASUle+AXm51q3QvcuymdHxErlJcMpEQ2KD1gyKSjlbhbM1cdU5U2K
XaVe3ZI501YGkAuMkZrFfu8QHW2lCxM2BDJ34BN3RD8pZ2N1iMuMz9MNeeO/P2jT
kcij/8tN4/Ex0n71ImlZbFD7C+SWQpO/83G+zVVjGA/yib3WOFlAHjz8knNnUOpT
rgAHhXhtNcebMKD7/r7WP7GapQjt7zwJ3bXbLcr8FC4tBpNyMo3uW+xuy8rMQamW
C4jQIFtD7yzoGOKQqeWIiRr8uwZxsBw1I+BFiRHkr5allEEZd4NWZBPTLa6HfF60
TD1bMKasbbL02djc2mjxtUAcO3VzHemy61hUQ/xGnUUClDgLxrCs71WzzpMddP8D
aF1M8gLyZaN2b8mEXJ4qtbjq2HFHSVZAvyuGyvGFo5zgFMVzPfdT1BXKvgj6mi8g
bcz98zL3D5FkhDdyVqR0TkHzg3o9o261oeCiO5napMtgJB9UI0lEZMkr/oQ4L4vB
qvPCdJTp4WWIXx6fC25egSk32Bp1oJC/CN/GpaNGvgZUcPjre0A/2wVO6ziOliba
76h5iP2QLofFdeBSBnVKSQTeKY2J20KzZZ3OKx0rdKCZd4pQUSEJTY73b8yP1PDw
072vNjSdYNLzbmwDdRibekqpNfFH7ECpo3r+HR3KZywzqzBBy7+OqByKy+12G4lr
2sR4I78P/NEmWdQuB/1faUjJHmiPl8tWM30s6X7xFh9ARL9NJpdmpgQ3mGU8C5+M
Oyqz22voOy1Jn8nWb7Iu+ARntYiP2sEOwr4BE2+QwjItUZ3fKssuAy0GjPOYFSS9
BYwD1HGnNK8XQyI6vGXFPHgL+uyWLmk3b+pz08S621R2bGWBzphRgVNyXeR0TO18
q7ohpoNNeYY2KfBDUFNAteSMyEnZ3FSNquoLorxwIigJ0S3kC19oEezeg+57ZZH+
JnMjtqo0yh+vtVPkFvf0c0Uz8hz7+baN0XeCSF7EjCXaxvCkeiWi1yXKXZg+gWZr
sV6wDKZ3VJQFEs6rNUQSi2mloTlvL3koo1GYw3PGJ8HDdlchF/Q3DTs9YXzJoUc5
IMuFWTPKy26FdBi45lk8XbHi/QOlItHg0DW8vH2QF2l7z+3rH/z0JtCdHB0B4jz4
fYicq1pYALbtzFHwvIjuCxwuBcedXbeH+Fvv+HTzrY22TBKlX4UBa0Rkjzpd4B/y
zPRJryLMbOACiLxbjKs2zPDomYqt7xVglKEcVDRf2GdTPsf2ymEgKmGeAEns+QFq
41k+4CUMtFJGNqcpdfijRJR2Y5QnESJhaJLzamxvGhGYPcF8kcf37F3R+eWWPR40
T7tQv2Azqbc7btkRdy65pLrK+jlkNZX6kFAg+TY3dIjqXbc1F4jyL0sc3jbT0sRv
fzEPXIQMi7Q7Dn9BJZJlsSvGPTzIHeKh1DwG8Rwhpo5J7DJAEu6NWK9NyOQUR4Y5
Bii7UUNJ86+cX8ZgQ+sVKkOw7u8pOxOeqRyCcLskKT1Nsi6zmvARGgSYhtnkCTLw
UKd2MMmgVOqFCb2v/26yWfWuD8O/Vh1gCxvb3tHGysrClnFwkrRl/ZOR14aLylB8
o4l3NlyHvMi7/MnxjRbOqMwyCUB4JCRTwkKAqX81lmDY1wZHrggJltNlhhmBD6ya
F1B5XZ/oYscySBg/WkkUVE8isWCzS//N6d8WBtOOr7wfCDaoeq5ApWt93a3XMbq1
kDQxS6bevTB/eNkTMpzg8kLwhQTN0xAh+apEbj7HNJDX2tz3x8533IPM6uCzZCa7
y/puP0vcbKFsdtHSyrTcQlcnTaO3M9hQE9MWC1uq5I30u0s6KcJ0rZ0p88igj2Oc
WrTEkWkBOHFKc8snWB0de4CAkoX5Qm8uPLuKc+WupLyDNB93YoXfwiaI/ly7jt39
Vo8ZDVGfrV5FA009ACb8zxgKfBIFIbJTwrt3JJQyejVHGZ7e3MftHX9lxouJlgG9
ylFlcAGcoFEKasD5FfvQcrS8jjL2h2PIrWpQ53nTtzSpIHT/ujkZ9jqVcuskYDzk
plekeHzCQ0Ew1R2WgFXkOaaVYZYxQgxOi+1BBw9n5SBcu7HZdc1OkA94e6LCxzJx
qwQhOoRXJQaRjrzTTVBnodN3NN2Elzkmj547EZ77d/FhMXQSZJoNpek9CWj8DVeo
7qz9zVhpSt0ofk0rhaNWc2uUgPlRUq63FtvMDosPzK23S7qXkBIgAENl5Jc2JD7D
GT1cjDxoXp/ecHjJfRoLUFr7gHMIF9YA5lXI/IuEaemRQp0VRVW1g6ItuXmidgIE
LyNi8Zc3F0obZSYSaJq9RjIo407Xdnih8OC+UnEneD0WZF05FI9Y1zo8upTCKLlz
0Hx8pPkqhUJGdPs1pbP2XTo5G6HXuvFmQh+FCWZ4Bt4SmGJW2Iz6b6ixpSChX3Ej
vDJDG736LYOsrJTyfp2S8okh/WxX90wcYc4AXFEF36RamJ6fKvohjMap+TJ306eN
6jJ3nSgGoiWWQJ0Ni2aMbW50MgE7xf97mke2Sbra3FpacwI4Hf/0dJm+XHDKjvaa
4R1bILEshyP4gKLUZsrUDuGITT2XObgZmUCaj1mBOezOOyaYp2iDu/KfZfNgRUtH
QnY1iB5xPvUAuuDmOJaCUqRD1vI1aDfjK8EUhw5gIWXZ8vP3q6Yne96wc7fuOhCX
0V4Hit2LZntttHMihugGCkvUIjlX7fZJ7a4H3JNKWdKGECJe8rYvuCeotFSSx6+P
0vFxmA5IXY1bMVDmIdlAXAikEto35n7K37oyBG2ipPC1lPcAaLVIZKeYNJglqGBG
fUVJzWwIhFi/WmLiUtZ9MDUUrdFUjOE0b8BIbAs7stRzDRiNz8zBWNAWHFu4g2uf
WHlu98LASY0UjNCgDr2lMXFsruZxq6PGnoG7FBVwFT35ztN9jVNI1GuqUrOns4ED
uUhAaOfmTBqRAim4L+w+MQNI3f2uwMswvbTMRkJ1DgaZBq/oin4MR4ZeOKyOdbhc
vYepR6KU/K+hWMPZR34j1iSDe+JJXpaYST7+3WTXGSvtYlYv22cdZ4IF0a/COKhQ
Di5CAiui397KE3lEMJORhiNNH/a/nJsaKtbUN6OV+kMdagksCZV+RzyMInCt8LUq
5n0NFnUdP0eHt902nPmQT2ynzc6pavEvnuf5TafzSfkiLfPxEUnLjwRz0IdNKIjo
iRcMINMXNOtrsZKBnJXEJK3l89krU0PZMfZO6nV2IBjxgsG4z3xR+EbR/IqOY+sA
fcSukVcm3YzEVHCuzFLzG7nTbucTU4546/nXbZscH85V4bQ4+N3vgni6x1Erkyzc
D/nuNsEXihIQlYG5ArWvPKsH/5yKN0Qmv9O2VWnH+a9SuxsZpb/7qlVK8m89cJhX
YdcjmHvuARG42zFcYbzIPUMrQSnJMEV7QhD2aVCBawxjpY/CGztHnQV67XhRY7lR
hOwFIjM8sL4Dw6PSzWDVOfM/9YpGT5cjXUj0hTBX6Qm0r3wU0QQLpJJRDuuNETx8
+tylILvTCT85moxNapF7x84FpBxUCSax3QFjtuMbn+v7LYcSKr3TxaqPoFWQ9Icj
pcGmMTXHYbaEGldJnjMDCIvzYBo3baoUj0mbK1Kd0t5on6eGnejo3zZYE/BYzaSQ
cYAfRhPTt64uVlW4adJow4+a1D1Lk2035JdvTxikH+fBU9woaCwwNdNcf8Iuu9EH
maoCGhrab33z60p+KqGXGuH6nEwu7m1YF1IIQrkQYez47DvH+xcQtEzufwmli0RX
sEjB8uEpceKYdN4aWYUfsLv4K3kiZl9AWfeMly+Uj0eUgr4KYoWh6oqFb3VnjUTs
wA3D61O4ciEYzbAbWXVOggQEdibltP/IHfcqdv3ama8z8k2jtma94SWjduFFxiV9
Pu+XBFWHG3ShdPgZZ0+QZZGBOYnDHNud73XyFuAKngjaOnvB7zgPWBc5LU4gHCtU
Z1nxs0Jtll5XpDOx1J8fxJhjLxbaIZv80jGjpP4Lb9RcBX+OZUR4LH18OwCU3DIH
ARGsxmKclhFOFVfBGwWXemVJpLU8yJSW09yyzTKYy+uEUhfr9YN8kEygO8MTTReU
C7EVTIYh/pmD8t2NA7jo4IeAHFOo01MyO+uvI+Hhm88FrcDT+DQL4QkG/37Nhvzv
89SlN3yAyDC5XJ6lficpKkGqRV1rh83kaT0IdTrRvTw9gml4AwW0NCLRw6EgYe4+
mJxmTG64I3OXa6dwcjJQQJPnRVfauLa+JwjMbnt9zHOwO+epVLHaKtB09yRgUSa+
QpMEs7uolMXH9jhPHm4fuV5tjOJvKS/Q9VN9xLJ+BNmmRsLs3YcwH0Yrqj6iGiNo
wckJ0dutNj28zTGGzng5f3Vv04pEiNloDhCejmhQlkxGObA7amu28OTdwEuw63ei
9GLbJRd2nB4V8rVoIvOySkxzU7AK6jnEqFiOYkjUZswCjqaiUrkiPbUOAeS/oMOr
7K63IlfUM/QcGIqEBfojm1flaWW7vZlDSG3vhpKMb2dbOKbdxtapQgG8+mgSrALh
nRSebDTqyKVd5Dh/8+RHCR98TECTMwfDEDTZ48h0+FMQmycDZ2F7DU6LRHVcxa+g
GmuFDGPhdKW+1t21sMrGh1JalCmdhwkbbuG9zw7dEHsQttgUwb0QbfKa37vR9LQx
+Hw0Z/7xEgcWs89XEwaxRwJUrFSR6uxl0bofShg9HyXa5bLWrjHCD/l5/z7nh1Wz
K8ll0t1sZ2c2HzgsQAvqTb4GA4N9Ca4TaV9t3qVILIKGlQacXblf3+S3u/LPRaQ7
by9EHm9j9TTsHwZ9um59tpVIMBo+2oJ594PJCns/LGA+vc51E51aJKTZpiSqSXqD
lYzJqFj0sMyeHVOjrje86nEZ8Ic5pI4cP4UkCCYCjZKyz8LN6efbH2j0avnc9xn3
jD/qn5AVcHpLRB2YdcR7q99XTA6+3oLHw4wE1TPGmW6YvsBz3YfeHDE2OMvVNdEf
9xtlPjjVhi0DHV0cAkl1A/az2oaMNhWfHiS2yVJp4Pop3s91vbZN6tjD7anhDVMr
T0iSHvqYb6Zrtopwn3TqtEjwhUiqB0PG+7aJrWpyPkMskbgjwrGhrTFD9wj8Ni/P
K+y9FpdG5NvEw2gVWC7VVPcmjSoX3fm810OHS2BnfmciD3o8JzPT4omznQ7w1feS
0Jd0Ufe5vCa+y19DObf+GKq9Ebqvd7eOrhKMWWD6D9epjiBUW/LuRa/hWUz426+D
nRhFgeoXArOIUqppg+fy06zXIuntP25kc44feJGanPfZ6cV8x5DaLvIfQFszULN4
WGR8ReGn1A1RvtonQHYF9yRQaIVUJomRlIUPvp+fDEkottXdR6CGciGnN4URQVVI
1Z5hcKd/dgU8rr1O9iD8J0otH2KMuAaG4DDE62Oh/KPp+cfgBlAGBTXymFkneJkP
HTprxbxZjc61a/9l+0Cugy4Vug1+vm/L97pc7tKAsAiXV+mF8DsQbETvSmeDAzLQ
ifx24NSNS6okQ0AAm4INNFO5oAeDUkDTT7BhYJBm4hJ+/2zzwzTi7UP2mm3spSlD
hsY9kpSbTdGxxGQMiQj9+28lqzk/ZkFnsRsZkPhogiWiKlxI/u1CgJjEx6Rkc5pQ
7VrRz2nqCQzVLosS5kwlArnKWPKFFxUUUKp9pK3eTm2oJE1FRMfa9IlBLaSg0Ltk
oaSBPOgilQjFOgcX0TulhjxH2ZOSrMPP6flq5+N3sOnRt65UJXx/jIUWZPAAWHr3
EInlIz8IBOSKx3idOcylrUmX9XENDXyYD4cjP48lxK9QuftB3Px28yROAO8t5Jgd
FXPSnRCDV7Cx9Zsr5ww1BPgoLbAItbZ5kYcwTpfpSQote/IF8azBrChXdHHKgCwk
0yj4cZBrstqOBr/38E2cVhDt2XZY1e+TkoD9F7mS1BRQOvSXQIUQw8T6+icrgHP9
cYUKWHxdZS45ZeLW58YA2fDqquwsTmQQr3msIk8iPs/PoqqO/dF5PmuzFJJ4JG+p
er/9/ecaAr4OxLwrM4P/LQFRgelKWYEbncNf1GBI86cqcgW3Y0CEqnY5Fw14PRAi
Bp4PWwdZukS+voKw85z11R5jsheEkh4X+YEqgVUhFqEH5QCqWNtF/jAgKh6CWumV
hWjV0HNMpY4xCKfYEPfmOi4GuTQwQ/+U/VZYCeV6ncOhOdOVhpMx0GTL8nAcMyWn
VNX7pH9a3/giopSj3CGcgISUuRrKIZM9It4uWsnVG/7eZKhiA17ciHIJd9jZo4UP
EnpfCkv7WRazToXuZk8BLSM7FAvdCGVq3uL1DSRu4EsE8XSvdh6SkwvleZTcj84Y
JyS/BtZrvmLWhkuqy62qBgAlICWl/M/J91yMA/5zFBHQOBArZcSRbWWPj1YLzqWw
Sapk5DK/7168QalKhWRKQ0xQSuDjgFgdbX7a2ciMUg31KW+8BOXv8wrtEuAgZ/LY
vRY2zSKirWQNwXzC3YQOC4kwAU1h48nPQutxJdtg7/FEShf0CSi7da1fRK1ON55V
fGAFgiGz5SzPw7BUxN6K4kFMF8AH/NtGFOiwkWG6HlEllmGq5bHSAtB1lqNyLFiF
3KxBsecfW7bFfHMqw7NJ2cPSuogxXkJTYjYcN2vgSPweLPlvcw/pLuJrtVvJF9ED
ZfCgP6DNcv09N9EqMmhjDcYzYasoZWeVkl6IPns5nSpplfbeU+jn/HleY8SqP5Kj
+EEBjTsJuvxROnkZQuVNhnH7UzXXuRfBqpfH/M70VsMjJviS2XUIoN+OuW9LtgJ/
FQz93LWhSGUM/Y+EVEYQq2MKFRuy3nqCrGOc5wTvIhdK3bLfPzfIekxfNLsgCtiV
tjWIKfeKzFlM987v2S759scu0AglM/Ud+bIPI0g7zBtRCsXxE4V2V/jSmUx5nuED
wsMWLL9QfhgaBvHhAoG9xYMr30M4adLy9/oanXlq89BFlQaVHha2UtfpfF3KSvHA
5+mhYHrKDjrxf1iPFLbgIMsf4k7a5IyNc8eJ7gXCcbwHijEC4CHKxxWowkJSZZJ+
IQB+Yo93w1eNfUI6tGXAiXwK1ZmDb52iDP/vpMeLnHW/L1b2TdOuarWiHI9T/u2W
nJ3Zri5GrcSgPqCn5r2+pd0sqKx7uvb+7Anz9vGhoPHw7iLivEQNSTOk5BI+VAe3
/oPz/LY7Nb8qWELE/UUxCxBLtoGoEXVSMNJqcJXi1zN8PtLqQusfWkQ50+IT/l0x
zY+CayxKBhhucsHrB0DJPdTxogB5X8V3ZlD6glNOjpcQNUGJT566ghfLP/1S17zp
Oi2ddt78XVyNvLWUeloAvvI09mIhk7V6eyV5HJJoQLuadjWDH+VN35y4XM3C87U2
WAtiPFum+BDmu+/c0Y7TV6+gQI9apGfx0dD7r4NpPmhPcpzoqSuQqmc3jzuFilMA
lPUpC4B5VmzKW3IdAeYwgvzvE1ciPcd4Lnlxpvo2vwQMUYxj4CfuHaLGhy2S0MJ7
w7KPh3b4AQ5Pr3rWI8S66A43tsuk1yO6++QlRnrqb6r7YjQokjj6r4ESwWOO9rzO
3sgL//yq0tie3139eU4nwN/WLfBltGQAI5DbQtpmPj9cp03vZe0PmfsOJHkocd7N
bcA1EojqC3T7NdYCP2MGiw+Nc95sZf5u+d3nhDQQm+xW4sK+pdMUIdEknsgDKP8J
ZTSRafYrIHTsZZJKQW+9oC9D/BXr2vCVzOdnIXGrXCgrZRGM8OGzUz+odDja/R6G
HLE7kBj/fnOZYRpFGY6lvBzwG+mgED5shBQIG48I3pLf9Yp98yFOyXPpE9QKF9lx
97ApJQ59/S9QWciZxjzVCOXcpe2Itldmy+hQIjS8ogTSgIL0fnr9WgEiK3ByEafc
jIX1d8b91htoBN0I+yH1UJYupThetCkIkhvI+ZkqwmcYtrI9fQ0r9g5mHbYBpnNU
3hm71duVnuIxs83pTM+gZVXAg+OEn2QrYwZgsXFjUPHs6dfkr/9EqaDci3FmOLS2
D3QXbSXyMH6ER45XEFL0fbUDMAblVOaS4PjJcb69xifnSAQ7YOjy0+6lsnByWvLV
edMFqAswxiM1ATBIh4r6J3GzckriMlsVQBChl2DoT4IaSdBt4NUbLIEIcvV2zQsu
hOIoep7UT9zZvbQb2V6ctpEgVQpkdj09Le4FqD+W3VvMYuPBkr2Qzl6FocTj8f71
xJ5mfzi66zeb1wF/JXAxX70pn9ImQQUM79w0KXqNIT9DHtV4TH3R5lpQNG7SCG/L
Tt3TecS6pniUVZOY76X2kRFADwMKeMpjzcCYqwHvbZ550MHzuoLMKRNYl4j7zIuN
kwpFl17zsxsLXn5aVl1kitt2lzqORVjuQs6TzKAjgUcleai7debtdLQAW9wdwKb6
+jTI6q/wbsODyaEqyDPnNPei4rp+SdJROQp+So8Ifi+kO+NZQTNCARo2DX26qXPW
1vANVSKD2OD0S8w8n95EWugU9/2jPRQ4K7tAuE784xD7/FLXyZL3TaehhYycTvsH
co1t1N+gDgujbntmnstbsjgYDDQ96R1qaIhB0l/jeS7PwiSK2MHix1aqi5G8/d3s
Z81MhbhWou47MbgzFR0AttjTJ5iZwLfsPv+zYVwIhusNCjbxJ9gIqQKbDFNN/3SQ
TurRA7I6ohCGidZEN1M6/TTj0iYlEEHa9cBcljWWX/GrdjkqMk1GwykwAzvZpUGn
KMyVhA5s6gZ3wsDGrSpdCy4e1AaV1nYmOi+p65VbK6sfQM7XdsXsFwOB6YKZ1s2R
tBB4h5GEldfR4A1g9/VmSPOV5Lr61plR7rE11Wea3RoNPgbPavPTJls1Y6v/vEiZ
S4mSIcaRdwV5q9V6ZFlNJg3NoHts3STnipmlsrfY17XVdrWbYUtRdpEnf6HZuFRx
zyeHnThkSjDcuy8oOKcFg7ri27IBenX3JXd92xOks++hFyAw/N0dTniHiruSsx5v
s2s9Q5wADqmwBgj9A+slkYpbqN96AkAwBcfnQ8cwex4GVeA58Ib1FCKMKN3yS8k3
RqgYR9TuBFliLdtHZSheMebl+7NO0pyRKMcaen69tbMXF/jZe5hFwb754hLq+LAg
bCGAYgDwAYN0KCyE9JyGfulalIH7OiDMoAajXL3ugIM+F/kMsdidpNzWvvbz9OJ1
GVyrfdNLo9w5UlICS+G6z33GbF5mA8zToWIJQKoj9x2IgWvznXRckh2Y0p8cWRcw
tPJy0MdnrULyss3EuxNX/2vkZx4/ktmie2OMCb1bPz2bya7HtYnkREPjWtjHwuoW
tfImXJONSTsP5OJ3Rs71PqxXj8v3FTvmQ71cIDYTxF1U+4wuL3gvT5bfPrpWi/H8
aNEGlxk8T10aYGBNw+0zkBTofqvBCAHQSoS/anr2kQ7GmO7VkF1OlvvFR1dua6Zd
W5uVXiiFNK4ezlKxWv8HAvlKBRAYEWvnMmaHKorvbiZxxmR1fv4K7IHE6OUscAAc
Ar8ir9VeT4hp9Xs6dqzNtV+5I1pKYYMqPMJgmwdBnt3N7SKkAQyWEjON74KPy+jR
kobon10wtue3h1KPtggrrVZbOXUQfAiCo84kFBw584USftDDKihbWXmHvG2c0pN7
F+EWhInmH5ckjBaQDyeewcyN/SSJhFYgOKe8e8/Z76i1mMiPjlo6gxhkfNyfxnsq
mgfE570eNVSE6G0C6+R1duT+E8uHJt00UAiZ1Yb6WN6dT2HKzhLVXTkUbFSLKSCp
OkWkkJt00AIWQmSoucB1yoOa9GVKZSIvF+ta+efF2+wzvCwYOOfGVzeI2NNtPbg8
Wuu9mYE+0cBJ8CNj2upd4HfaipopZWeNO/X4ynFNKopXYIxq9LoSLI+zuKX48XFw
LkK819dtJfXkIpl9WQBykOExG/cLhjy3BuJb3ChMdjl0MB39n1P+sJn7vyv1OX23
InAkliIXFcYYcEhtqFnr5ddQduf4ZXm2KRQZwrltOFu6x2LffWH8I0+HIwefND85
37H4YK+vfSYnlt9W3PBZaAXkIl/FFUEhVrtGM/QGwzTgGvFosDT8fVTkUh5PSHw9
LCxT0TerxxqluodD+gG2CEMAsT/hLSJNlRAA5Jnpq8mdFoz8k6LIgKZ0jA0fQIOD
K+TwuJU/30nSO1/wOY2NSFNV1//2aMMZoxc8+mkUW3XfXyeJDvkZJarfo6FDZr5Y
Cmt/6EFYPPoYHyQ43O2DJcUJfJAS8fbzY351lEMwec3YE3KNF3SOC+b7DUfs7Kh3
F90pvFE5b/ignG96eKGAZc1Zs/FFtVNhfq7gdF+wZ3NaqpMUK48R3QK8+S53Nebp
AZZTb4iSjPwdZSXlUlUrRsqwtIYfd3AVpmPA8QyLIYpCpv9j6utWUnBGWQ+vOxVR
g02nKesNnehOHAio3VyABDLGL4xsf8UTlFXFJIvOAdMIfysGEvV9x4QgbKFL03eN
Wt5BAhG2z7GIXokdN91LSdhJYPNdcF4jkjzolZx3/plEHoD9xDVkBvDDcECN608U
kcbDaypL8i3KuRjXQeKHRo6Srs86qU5Jqso0NiXjVIEaYJPF1piEtGJW7ogrVLZx
qVuwJLDNu7fEkj+K6A/7WCkDFIB8VPfVRqmXdriEw7VPPTI0ySD4g1p/1OHOQrki
6Fkjg/MTYQWLnO+xx10q///TMRmnE6+A8GPLp8Zn0hwGwIdfMwgYIO6GCL+kcfq4
BqbxV9AShJg3Gfw6b+pPmipazZLnmV9yIiIBicAoE1WG9r+glMYAbHVPb6aHfbdu
DLwMP0zqgvwpCPb/jFiGOZv5E55pbGNxct5wJKe2O1iYeGAxJBc24iMpAJGHh/4I
8lshfA4FFaLHhq2hEETifv8TUYy9oQ2DqpquESjYDl4UgW4eZ5EXEXtDJYZ7IbFB
tjwoMx+1dIDvXEj0/rVeSwQBFTYlmGujqm4NjYIiRZLiHVKhhn2ZuA7YtVHd5hua
tSrTO2fInFPgvAvsFc/3ab7Y+gi1vSAcIXagkayPvA0OfA5P1Q+RqDsfWy6yvcVF
jXMnaH2zMN+d/djXzl1nE2vkiXExHSfoBQszfEb5n1rB5LT1DreTePPznspgByIF
r7lfvZXTpsW84kfnCxJGwuucpB0j3g6fGFTESzJ+4GMYgoiyISkg45JiW4k+Y6Fp
7bl2cYg3piIDdb1jX2/e/t+MTS7vCOj+Ip/n+Qc1MecNy0d1s91gpopiSFjKP3aD
FHtKDDLgFz0XQkdiQqn+6GMv7Cb4vhY2+0yBnInf7aEE5XsbJRqU1hn2JE9FdnTc
lzKdMSs+X6unOcNevU/eCeqXXv2Ti5e+OP1+DdAGTdC6mM1XFn/wamoq1bpElTIz
5IpSJ/nE0DnsJd6RJZaVpxhtKCJEEkTQKBZT/zJdMITyFJiaYNPoYBU86iMfP3TD
Wd5p4gH+1GUOFhOFtlRL6fusWQ/1ckaKYJg/N7Fh+L+A8n3njAVjYVc0uB4N4YJ/
hGvs8Ikh0bhjl14wDcaqR5LM8Xzq0P6xM2XNCm9uiA0//w+PcAequ8/wPiEruQYA
oRDqKFT2GYhSWPsf9kjKlHo1N5FU5+q6RBxqI3hJktwOYLy0inIHseCbyqXc2XKA
cGndvkhdoAPYe4qHAl0mafA0ailLO8tZO+rGgazSsHpXp6RHpphHs63LCN68g/hd
dtf8wlykw5EScvWGfSDlDnwnTuypm/NV58VYTr7YFrnD6GFDMj7/K0yJbxDCP1Ue
07H2FgJDcmLKED73s4H8qiKaIJ3TCObQUHKrvNzlww1qB+cwVg5wlYvnFBRy6iNS
Xn09UvvKp7zHsi7cX6anw0hMmAQ+pJ28NxJkFeYfIryYre87P0KhH+IIuZAEfiAW
tT1q4k6ojxkZyhsz1ame8wYm5Haao5s4JfpU/X3YALgWI3Uq8hpEcvzfjYUcLiSW
6NAC/Vq8UJrkTYkC8fRoFjPRVmzlsHjEckpYf1I2QKDfeLWJSPxyQmWwu24dOuPX
6aTzabzalPQRTkNFamQ09VBrrSyGznc0DAZVK6JNd//YGs/LsN4CZJUb7RJc9yZ8
ZX7VUMks/eDN9iT5/BU7WWYDRDenNxf9lGjahvHAG/QiyIsBDjiZq+Om9qmOqiHP
RHFatlpNIpYrsOCzdkbMmbQ5+4IaCp2kEzH2SZ3aLM7XTEKjIERcYY2kuIYXiuh9
T8KdGnvtoalZjs9FVtoQzEgjHJdRa3r+kbYPqSfoOoOA6TviOCDhHjk9GEbpgeH8
zJ/Ay2ex8biHofyKNqv9WazNpun/g3n1+xatrgdGJyPwxDIKIayTtaPEgXpurnPc
kqrSsubmzOp3SDQ78UGQSvQHEOGx+c2aQUJMzFVjuGE9LPU2Wzr4HewhTLnoLRL8
RKCaKp+cmlpnyP6UP4MIfDNKou5mxHdK4Xw+x8U8Xi7o9rUEphjWVXEqOrmphyh3
a9tstIlBn9UGl/o6qfBYPv+vjN6rJG5bI4xQZiUXAlaa7cdSfxw1hzyz6XShfv1c
Y2ife1+oKkVsjFtmNK9/oFFNgmeIkpqiRa3heS1EzJhntqyVyCkO9FzH501Psyff
6cJPoIkp3OvKK/HRP2pI/kuXBH3CgB48K+HYgv0EEtTU+aLVuFiuHry/mRaOu7Ki
2iLyCcJWpNX1DT6EyuSK74hGC0VdilkRNBNPsppjyLijzI8wygsQqaQk0iEhZfaQ
dnXu02ZaGtzwbG131D++a+JXTRLVZUUZkMsrJBcE/+wttJbBZFBZfLfZh+hrw7aY
8G/weuI3sXrDiszZocVLHHV3mtitSGduHGLDgu+wD1V9KDd8a8xZHX4QhYsC51+Q
s6ayhXWS0LnC8aVDiLVZcDqHzxCXKCOGdrvr2nIvf7f/aJBmKHtv/mcDv5vG04zQ
G2yBdY8/o5h3she8ol0/k4wliQFEkA5k675PHx5X/ZcI8C1s/yd4pN43EOzF8sgv
25j6U6Lbsitl+x5CvJ7rpJu5K350s8hQmUlv1ZMm/yZg7PgiwjqbqHzv/4a34DgT
Usldyfz0S4pL3VrV0UnmZ9LuBxdAiAmR5wB2dr7k+kOHj/uVYVSkawGH8V/Mme2h
2mGefl1o8kYarL6+gjcRBvO2Xv5v6kUY4D5thvZ74AutwScPQvyHCmJYi4cyTDCy
rcnMDqPl5PYPXvlgvOB76dEpYAiOfsLNBgMyLx/F74xmeV/DHr4yIeAm5DrfmZOk
CPli2+O+171e+9uZ0lmUSnn6p87I+Blk+VVQvKHJH1KiUukSuSXVbLdwoFGLNZ8z
BAmY40G7ta0K/y3e5aUMlpaDgPRClci/eTXjOTG+dNUj4xVjyuwo5G0eVs0dRAWK
e019HtjV0c54/I4vA7bzVb6G2XGaaZChMr/jwYeklwQzCgsTBbUM3R8qn+FXOgbK
GLQrSp6VsirizIrDkWXlhqQDu09SHTS6SY9TisxustxFSZ0Yj7z8Fg9tslxk6DHk
XBihIBrM9IoS5F77ePQ1MFeThPMYHCgjzR3SNCU/Vir9okJtthzVt5XGrLCdBOmn
9VGlHcMO8jPdFgi2iWNheinU3VB4tJoamW05BNP2zREG2jZ9M/msBXKeoUpr1Ah4
dEyUMdRn5cflt9gDByb6EWxZmpNfmcMlNDghOWYEBYzb8WlhZb35YdIzQgnmXkA6
l03FrdugM91Gf5LHYokJZILwg+7WkcjPqpfUMRCA/GplVI1T+KZq0/JaCE8HomiZ
xvxILrE2fq/wD6CLoiTdc5PaBO9V4+orW8nO0J6yj4vkJXlgLRRaotpJAcO89pbd
bHHXKxczEfR/ItUTJNEcn2X5EySxqrjYAu+QjSVe/zLPiSmiMcp+nQJCn18LhmCz
Ir1yTQVPLaN0HvnYGHLcuGtJVx3S4Pb11hDD1D5ZndrDbe4wKYrqxLRcVfwprAaw
vmNtvmnBE8PpOrli/fWieqzhYQbrXeb7NT7gR/MNc6X/MD/oWobgAc/QA8PqW0yc
Ty3HBqJOLKDk7Muwa5BfBPZToc7TRI7X+gK/XM7rxGdltbcOQgnrjd4+vLZuOFKy
aCk81LIGrTe1hUEy7zu9Pgt0jLUXKirKsXp6Fs+TQm9+uuRXJ0TyJe8ukKh8H9UK
VqoOPZk9JIIMBoC89HgNJ19Gbe3X2DEOKIT25s5ysw/CEhn8aPgG/Ne5IFW0rW/I
kWSf1FZEmMZAlf3FPO27/k7XeGCy69f4AmsPBRY7ynYiUgs9ZuYlLmdZmiDnxGQx
mFMehF/RUjp6K5bjHC1iCtWLZGKAvwfgVkCCVSuGYf/Q7NtpR4OvC8JV47ZMUPin
BC8Nr43rE8jR14y34vRJRSuy7dJiZ+MGwyCT4CcCTF8aWAke7Ub1rUD9xVHXyhf+
853o9f+7ncfQq/xDFczoj9hcnPRmUDTOVKBMh7ZsWmA11ijtswqvCXILFmBlXzGK
FjXmX8P8wzZQFPZYWLlgs8XpwheB2/Knl6OmMt4NovcOQejKoq5x7j50gsBiVcAY
ka5t9r3iFZnT3vHYb/P31ao5dDio8vRCI1+dzaZfr9Xfpp+OEFmCS5QDfKuaezjS
w7NhOJZI9ZbLSfHraQCAL2W6HytXVpjv+tXmgk0CBa/9JHoNPv9USLSI6y7cBczA
PL290R1NGbUVBU4TSkZpJRZok20pkAa41C5bbNqPCifaRKCrEXu/bmpjgthl8Nqg
Eniei3j0EThjauctLR3HQ7/PlgG9CW/3WcqKhVz0qhie7GHVJ+gXeHZALiS5W+4n
8tixeTpBA1wCctcGBG7DGC3KVxuSBAsYxBDFz+pWigeO24CyGjm7+SHOF5FU96NK
7qCozJpLuow+GotIUg3aHwDOYldi+obZIlW0IGxl4HkHT8HVGErs73yjQxJHa6Pa
c7FccINYL0LWhnHpBN23gSMtOM/B+eHgoSFIQbSm7mabfWTR6kQRCJ5wgbPiPNQi
WoZMyUEENBau156xTci+AvrODdd/W1ZeFDy8zOrPFvnPsJbA3ufq8XYsKlWR7ITZ
tmAli8RkeKEqyOFR3+LbkZalecp4Fm55UTqzBpclz8tlbFb6/ynmhliqd3wcmLbx
zIc0C9i5FLB/xgT/Sd+e/S0x4u9T+p7Wb6gVlnUk86zGA2rG4FfBD2uHYCnp0WnB
kRXE+dtPb+K4pVjypq69VSwpVnw9GkBtf15xHLXKQWsRpl0paHSbePemCXq6pwiU
Y5DznpOIfb07LtBGLzeVnJD+iTD+M5l/xee0a1pvN+hRbcYVgMcqSGtMnR0+LWoF
PNmrmoshcU+QUAofuNgHFCeaj8QLgKnpUqTgjvMEdDcT992G6tLVjRgcdyP0eIbs
GopYCcaxszVUDHQmjmiX+Zvxcg4wH+1W9kWiHHDrcctKq8DuUe6lfGWJlN/JAQhQ
U4EtL7ZPqLS9PrQbKF/fu7DYZnKDGSieM/CW5sAnNwVIXGdhneODln91CfwPDYM9
Pbi84bn+cNDi7UtKkDZW2Y572tWcFlrJy+USTW9o5116R5bRfVAgsrgOnfhK4lPs
q++7MRGhXXoIL1zq94HzQhSDJ0BnCU3kGkSWpPB8kIsaSC2DrQGUeAINWtYe5xq8
P6BndmnDuw3fJo1MZWanN7Qa2mjsVDzPc6ilM7QOLDLUlvSx187oa2v16uLXDZRb
QhWXs68fS2m32CeAhmujXljiCOgtrkVoH0Yf0l9pqa/dCmz1RIzLWiVp42sjW0kS
joSJrppT4FAkmxgTJhP4QS3+TRCfnvnIUWgkeT6iALFJQEeBZmGNVA5Vc3q1xDvX
UOX+F1AYSkOwoy3nqYnpP9HKKUSHv6E9SQF1gJ8lG0a/ExQ3q8GmpUjj0sfmuFsb
s4/pENDFind4yJpO8yN/dT0BszbFHOXPebrYUl0VJGZ4wjXzeZtE16su8PLP3kDo
LLj9pROc+r8shubu+bkxDPCzNosiURAwBpkkFHuKqe5vWhRg5OZcd+jfv9chpGDG
JoMrTGZ6Mv4mm3pPGNHWf0JR8ibjjbTFo7AZAa5g8+TU8hAm8RFkjuuDgHIU/PJe
ZU1iGvDgCs2BqMujrhG+rBh1zrNyMKeWVzQHntemBTGas2CWGEGMfu6svEX8f9Xq
06yyhJXPB+ZsPwfMTQ41MU5Ck/6Tt1AObInPveT05gwm1qA5Y2A/42mpGZnOWFbq
JL+kdDS7S/yFu3O/MCUkv3G+r6m8VaZyGl4VtNkVncwGVv4BXd2C2mzyFxBY7nVc
jWXB4tHv4b/M/kxoTnGVtB6Ab11B5m7aWzUbXdtHs4qv8+SoTyhP1+7P1Xq4sGHn
3DnuWlMrhN9CG80bjqvvNa/+HUg4Zh1+05duL1GnZ+HpWmC0ZU2FAA9KNHHQFijj
VbuTqLN3560GDOXxJWawPvqYWSVP73W5MbOZbYQ5GeAcQBsyyIITlRZcRMTLCgqF
GqqalATxSjWRplK+SWaK5c4yQSsFOTN3j2DmvRY7SoGGx4F+laN1wEZuAzLjZMe6
uVpGl+TEuAnJPFs1YT7j6NY5s8yu5NY9kemZHei+R2cpGfx2tPpCYnQATF28+KFI
iyFric3yCl3GiDZH+qohZ8Iw+3yeflZER4Jlmzu9ubvYf6wEE/hjF7Zp0/c752oA
QYmNmlIKesITpMow6mo8MmT3W1HOuegbxc5iqjGLWCLMgfXrG1AqFKoeQU7Nx+7e
PNBkzIv5IYdbKjyhsLbmNoLX7kkJatUQKKCcTJFHMQtUuVxiBs1Gg8suZDzD3t84
ra+vQopF1TWt0t94+Te47EEZHRWTeQ9crW1+5RpcFkDv8mPGgDTl9kO+yvMYP7GY
6ZXtYoEgxk3SPok0kA8lS5FwmH6PAUipFaq2KQu0WuGVUO5MSBLsUz2GTpc/7Zyj
+EaEzlqqSa5Zc+7v0jER7Sy6VSoEhqycntgD9BGNX4/gU8gQn0JS9hLi7F5CJIZa
11AaWpzq7jeMUikQl1WCj/DyYsltcdZxkiCMQkrwtX5ICJZblCtO2NlN8nGCT9iT
mcsQFyPQyBHy9TkGowXXZ6ilU4dLav45CEpxS9p9OlOmkNQRM3Qztkpj6tKG+EcK
C5JukYt+8bn57JhkR0CtpYxCCSsXmIlGb2BhFb/0fCHNxmKQkTQ567lGqnJdB0vx
rKRIzoMfkht5nVg4zQFRo6YgwUAp4koiBWsoEgSMv+uD1Rs86mpDtMwUgbDq1rxw
4Re6TGuhZ4dilD9GXNGxQcCXqlx0QQk8Gphc9+Z2d2MZlwD/CEzqk6kqOxrsVSxt
L5F+dLqvFkkEdYR//EqmWT0/PZs0r1om+tLYOTCcMrXocT3+MNGvU1Ot2f7c8j54
qngZcXl+p+ydFC9dDW7y24zBUhhXVyiDSx6lDR/TZKh21424MnSupk43O9y5+f2K
D3GJS2pKYL5nk3EHuLJaa3e8a6+dJwd/077FDEWJ6kHfilRN/r57z0nRuUp4VOUO
WL9tM04bo6Ev3xMeqdZnTL4ktGarNWNdZG/PC/yDcIMLEnfevU2jnk2RZAW9Go4m
P/58kJk4SgFd1pGUCSjfcQe8mP0+s65MxuTcH5Mub4WlrBS9X4OEJuWnZSUqsNkO
Ya6NZ0itgPyYil0UM1kYq8JnxguiGRHcVeAQTiiW1EEI9HCaqQ7zOwv8ClBMYtnV
P/92VU+UI5Hpoo3kIvgj3xllxVWcj4brF7fOLvAydaz7Qhy/3PwdvyfV5h7ED7d3
VV0Gx9x8riTrvTE9hSytH8oqgR0IJBpAim/Xf7qMoRQn7W0/gY2YLt1u4g0AiEjs
8quYXjZXqgNvRyLdJfwWwsKwVvcJfP2vbHzym7V5eYs39/h7pyf6317a1R3ovvgm
vMBpN1dzQVuBFwWqrHSdSouEc6ciNIFSzeJrzLBKzmueMxIMEIcj7sEsuqX1tr6H
fMHBA+9HoAMtufwHXN8c8lAsA2sn/Rw9ROF+Fyokp5VrNTTOMeIWPuwvwnAXCKtI
TLD+sF1C4NuqSZeif99KGEIryQyqFt7w3me4WVypV+mNR+4CRVkVJ7avO0POuw1e
Wls3zPhNF5e3UoiRI7p8Cqz7KxlF9+tnwuNgR6peiSc641FhtaYpFzvrBuk6YTGR
BMnw6R3GyN9lFhPaZLdWzgwACTkJtd+3BljYOI/gBwuxxZ+bMj0mq37qWkK7PZ7i
H8Tqyr3Bm8+F/6xv6qDXZiadEh5Bswp+1b4d81zkYWbUq7Ltdg4vxvkNJ759pv4F
5Aqrq8mbVbcCnKMwueO/0D8xoL5RV/ti9ZmnzHQ34Xe5vNXnZaJ7TRAH0nuTNGlr
HnMguzBufT0tsCpAZXHYypj4zkUB2GlnfL7+7FMep3NgvKvoCCNXXDGrGSohEefh
iFvEOOe+ArFjkvQd/9xTlJ9v7jPGaP/8eIZObYnLetLU2WvgWQfggHzAihs1KRhS
yP7DKiaxpabRnU14BdYTwmfgbd0jZFM19VLjFkxRndeQdyLAny2midmPETVRCdmY
eNXgpyH72olFBgS57K513pOKsxUYSuEK/ypsirRyP2iCWmBcmf3onuyC9FQvjt2c
mW6F2u6QHSM55v5rw84F+nq5fj2KCqX4MWpgEQJmwBQ5WnbFj/2QV/RJFmYXQ5R9
kolutQQyzHdO9O650cuqR16N/FeJigejjzC7rd0bE2fcm9Z1hHfbisQ5zGpRHjtj
j4jwI32pxgUyzdnUMtBDAhQnOAtC9zw75q9D6SzXeiH7h4Zi1t8/ZTZylUlkZVR3
leSKBi1in3WYedb3djgs1KwDRr5BTkzQrr2kqh+Xes9tf95hd96pR7UDLjML6AQo
VF+cB5N7Kg6xDTLkkRvzIoVKKTh+tSRlZ9z5EdM398Ug9hRvUnigoiSXhZfXFqXQ
HITsBv5m9LuNzZmSAnJEyP3krr+vN7jOOzibkk1Nqn7whK+wtTG93Iv0tBmC9ofn
ji6Sirw1xPm9A2vx9PeSWeeIwpRuBAawMSiJ3PQ/y8RVfw0C+bXTS2YHyCF/YH4i
aFQzPzGfmHZqMPWoTc1eJjJy1+U2sJ/PZt2JlE44ugXwLR3h7NGckvkGgHOqQyHc
2gJLmuRVp2NQP8JCnf6rY6lYmi79b4a7SdrKW/JwFWB/ugYxNG7XMk6cVEy/0cap
EVInw9B8cZZbK+z2gzcWiqcaK4I5WvGPR7hnduOYhb+Nq5LO5NHYslvrA0EGAo2z
Y9F3P9TYloKd969q5S0OAxBaKxgSSQLSwMsZG4qD0oR8nF45N+qaF2FcaQ3ZXsOj
UvshomfZd9QetnsoDn6izkpSiri/cqEcnGiZNYPPa4IBWigqtDcv2j/xkl2f/csa
AFPzcV0dLt+9SFb7wCizKyZ7fV2wQTPKtXKr1R96cC/tFg1uwdETeZtmqpYHhB63
sZ/Vnau3swrH8ebolZW5soBAtNHoSaApmcLry8k+zDZdMxCT0XV57tmAP+8hA0Zw
aixNWtLhaYv5BZCpUG6QJ4xk35qebeCNXc7qeIPDisthQDniwocHgJiIThKopoNl
c5OqSFRBWB+MuMnhP7Dy2sQpReq/UbnM5lBUa7C3enSuw06fF60reAdbEPmqUSTU
bk4UcaOynWbZW8ET/Xs9PzyhWEJ2lVo1J97H2QvMn9Tkn4l5vRU+d6CjxItFjPNV
YGMlf2VexWLCVLs/4V2Kj4d8NGc9VxEFPRwUlUhndnIYTUsYdFvW8sPCHzPROBPs
hH15QHNv/JcgFnfDTbp+e3kWUx6HMGp7UMEDVrg9FXrdvikNooSd3aI8HjKO+E+m
qEYNNJiJ7iDgkW1QQP3RPsIbLHF1cGllNRExVMwDISfcXUfQ6yr6i94IfUXQU5B2
RR1wuV7Z2iRmZWqVa326r5TQMxg5qc80P8cShHUwvACO8vqz1AbrNMQkMb9nv89F
Ftj35yY1Fn9+jXPKB/mlJa/k/55p+umUzuYDF63YGaOV7BuWHOKyyktiFWfeIMI8
fbx3WVAngmI9DOLn4mi3ArRhKISXs1CDUubcGEctbW9jt7NLUxEo6Zro4ZA2rdFi
OAEeGPFjvBWTbzd+zSYXRVOpu+dfX7XnnpEI+2+6qDosko8gctxm8fJ3y1Efzuaf
zatWNFywTjwqsb96KVgjQlCTy0jzyM+KxlaM1bew6cOqz5Uhm+bDneRfq1Y1dpRz
2xEaGUSgFNyMk3PUPY6mMyqGfaT1QAzZTxr1hqigfvcZjRRFNyLTq0eg9gxD1/UN
l/9hEUaEZMgewTu3QRlAU52hLLrxZwYbKZRXltafxI4C7E+WxX8IvEPXRMopqjRB
3o9B3tM830uehbNby/hINCExFlkAULQc0R98ZVwrIleerL5TpGZqbVFjR2OXdCwj
7m9aTB3/pMm9a78erlzNXAt6tqROrk5XC8ulUA8EyQU8EdF8NIthAdP5OCkY5ZQa
UkjfgLAPkrt3AYXQ6VockX/OfH7VzRtKEjGARYS3sqwU9maNHDuebOUcsWTOxZOY
CLaOQMvXHntopa3oZUspoPF5nZjxPzzZcX/8hEqxLLJF3bYuHubxjFCtBkzkAeve
dBV3upOVfsqdcWsoAZ1rs4xlUQLjb0yJkJYqTspqyLttbkgNvm9w1PKmOOMI3lqu
pBBIATi378igVq3R7tMOdeTmfq+hjpvqOsMZ4LaKP5XhycqbL1iB8ogiJSUGmszC
KR5g96dSMQgAJeREr02fKaAtwjuVfVPpb07GeQk9acJEFQVH6EgYvZ2o7GkzPS4n
9hVZlOsMObHAxkXr2UyW+MDhyiHAz/77lCplArAGiGAd1WVtSX8R/JeuZ7PlumxV
IyQY+WyXkZ94z8TznWuAlqYd3ixwXxg4aXu1AWXSWirflmoJDrhSU0utgbPhpPyt
r36rDPoS5IQ/nDAhgkKQ0yGVwYvVILm4ckrAVVDhV+5614HyV0P1Zkg5+AD3Rm17
mi7qjQeQuH4OpnYnXsaXaGjmEubKIDEwqIKOHpYZ6Hk3elVc6FK5MvstJi8G/+Cd
aghyZ/O/5DtvH7KWWhpSngFokkrA7y1Rc3fhPll/0XzV83mEEqgvMhjuKAzbK7Dk
f14vZ/Dhc+bQohuWm4s7KP3LRcHOLlD9tybS1rkA9xZyfyAOsHeDy0Qx+VJFTMLW
Hhrdyfb9oMiu5TMPmjc3J9ElG3oZ/2cr3b9Iw8RJJ/ax66GCfx0so0S62SQ+deEU
DGU28FpH3VWvsbeW1XNkHE1a+FAkhLCmIcV0QNggaEOwQMG8oVVY59c46VHIpZz+
P0DxnWZHYBKT89J6Sfjs1cRc/8DDHlfhnkm1Hy+K0SZi+6TCp79BrwJ1y/3GXbQR
yTTMzkNCwj9XZKt98yN3C+iYTHvtU1eaANRD90j2w4aA5q/mOWqaJq7/u3gPDqnD
fSuXYU6a2CJf0CKJ4+XMWaeJrP3g1sMc1hcMPfQksMHy7OuwNIVeQYmg7LouDgM2
KExgakdilkLt9vhcG5aqF6vjveBc7vSk1idXaSoHlyiMe0PhSEzVIgvED0hoID17
chwS3qJ709MbfekgR6QiNvl0wR5XjZpbRaaPRDT215R4RCkhFkH+RjV8W/tEGbTb
nWRizjMALCTGX2t4vuQIy+VlSunhBLIQzib4t8KaW/ic5cYSKskT4bgp0zkFxkpm
kZe2nkej1/R9Z3eJmrAwQSZG9PiHLLgRunzMapur4WzQibUOYhvfbzqNeP/K4RXI
IT9ZxmhMEMlAM9ka38HO/3eYpH6Z9mKAP9rEgSn7ht99U2lOjz8zwpkY3PHEf9aP
yOH5jAKQzxlBrbI50xSNPgfy9fmuzHhFtvd41K4Jq+fpqfM88FFhWXgzSkZhD+c2
ZNPScZqwLZY46xDIH4vuBc42pR0A56jDlYsrMx9ZmV1kiX7KjnZR27cpMkVMIUB3
P45ZG1MvHGWubVZH3TB0lNEF9reALy2YAOAtRwh0WiTa5HGT94KRwsw2VkDygckM
qGd87c9+jaSKxxy75BDocJHzkMwz6cFLVtv/qGp7YIq+rr0VJJAWzcwUS35vokGJ
i3l3elfd8qljZykWLWpH/DvtvU62OKZ/blc89ISImeH6XDwQue4DTLGeJ+Na9bEN
WPC1SUaRl/m1hAH5B8B37SfcOqbDL2NIaJazSBj3SWuG3EKb/Bk6Mi3QRPpZW40w
eXpkF3EqiN72QcjGnt1iP0zmW76VsB+p4wqwf3xPKe2SUk2uQSODA/OPgX4UGci6
vdZW/XgxYnYNO4J45hGhZOkxDQ4vahoebK8gdKIbPXs5v8l0hCaU47GYD800TIni
b6pxl2keeGA44lKy1I1+b4ORLaNsuztViUbH+syLpWC8OjgnKvWpgzPfuxD5oWue
k1mq8eSeln3R1qeGPPtQvgy9r+BvA7jFJLSoZLlU9nmrBz0G+M/QLW8P390sHUPA
jn4kdnAKHtpUT8TPw1k3Z4lApdFdNxuaWghyf2ILRUn875ELCFGOwizTIrZSU9lb
cDMobd7Htpyv+NZ77O7VsiNZfN1pMqX1gVixitMb19B3EQ3DWe7H4ssPptqjBG9K
2dP1iRC3QcHg/YrA86tP105F3GVi23FDmo3OJgKlA9T8dYxrSa+4dJKziD+VF8DY
xoqxfVhY97dgVrnWNjrkfRMs3rqY6vADUmyWOtZxS7jttSCs8/7Z3/Tfgr7xvZtv
0uVsYmLQnBRWqdEFOubjWPSGK518n2h0YUEqn58SQMlmXQfvFEvZkM22R/iJNZjg
Nt3pPwptfRmxHDbNmDPwMfNdj/Ro3oeV00yXlkjeFs70OZiWdiL/FKLZwm1ssZ52
a/Ek539TECVZwBiju6uC7qgleG6jDVmVfx89ZmylwpGHNRLumyHFyG/b47TWGJAX
yxAoqqLoO/L6T1WmldZzEJWySO4zmNWvhqXG4NqPqad8Q7YVWVPci0CWqKbaHvNH
U5z7kgujAABBVOzQ8I7dg3OdsrRuHkSgRlCqs09A16/ZdnHOrcJ9A0kpLcd8lXP9
NCSb+X1nXU0VqEiav1P55jpEiLN6Tj6T9RP+P7pRtK+HLlHH1QHasQd/k0vejyBW
LIVrivqaZxLj1lCMV7JAcM0b3DIW9dZ12EhqjkvfOYWwXEFiXgloNbBA03gYAJgg
ak8CNEPq3Z4aScw33PnI+rf8YaJn6fv0W1B8kdOufsk79APsiiACUs09TWzXzJXq
seDlEH6xP+T5DIOfVVSVpq0YEF3d7rVjQWPUimsABGIMLCMYNhDP4OqAkMSRoGpD
XDgivhM2YbieR8PqDZQOMEexfdk2LK8qumwI6Q7J6Urnm7N6ivCkNPEYbfgchnf7
JuM+gtXFrQvFSmNUbvDhGbwTKkeHm0OcHSghSa4cphnpUytsM54i8gyaZ7dLSKr6
R+iUs+SJzwzpQ2M+V+8mnjULxLP0HACY3sriSWbGGeJIGXQH7N/jEReN8AUWGv5H
8c5RdbQRW9c5xzhYYzxpYZY3XH+hPwOR0LfiATkHNmDkQtGELBzwv5M+8ypU6IRt
o8qRHVmMfF22v9BqAdcV9uNdUHrnzTyyw2R6UyKKIIzJTCpJCaEd+W4Z2rLtQBbt
9nc46Q0N264L5A3gdczkq7f2G5xMDXCZd3yiLv4ILRVa/aZxqxM7M1bhEdav+hal
VJ1IGizjInZ+4T7prMspyi1mHMcVmeLcQ+bKt4Nm0Rhphv8jUIjF1FvOnId9zh7X
MSxQWcioEfCLrCwQ3cY8C+J3i9G8pUf8LIMA71iuLyscP9HtL3gvz3RqIePeiBOc
fziCMAeAEDg4ryrIw/ZLCvnYTY6VNehBIoBLCQ1JxPWKIrHebVTwuvQ36ZWUv/dO
jxjyB6qQiAxszFDYNdJwDi24JXomL8PayfI0d6RW5lXr2mFC4/91gGUtmYa4ilWN
ckniqzcXgYmc0IZPSXrgb1iaBeRrrHRWy1Yt/lckkDpWNiDJ2wSgQZg9wCpDK3NV
/ymojOilD+d/ji9RDqmSu//b9uIWHlObezzeVKY6IOLmnSNu6wT2beTjEpm+j2BN
URPldBfWWc/D9ZIzgsligo5pTzCKZfXOLZ42sin/08/JD1/NjZgmJO/aarqXwV61
5TPJD/zCyBSTlRKx8+YHHIi8hfJyMZNpcubBr7i9deXh6pdXjLBcX3dcWihmKQeb
Y/SSBRssXWc5HCqIkXnxqjjhjrwqP6QNAnNSIxL+OlS+4+KJOg2OnMxk7fy6vOEs
ug93uBEX/wnat2YiX/osyA9NpEhc/QsmgqPJQgV4Pqeh+6aUK+19d5uGL3cUCn8S
RdynjBCuB07VfWf6kbOmuDyDQw0J01VkENKGS9YTG9od+eCwiLlHFuPReidROHoV
AfwbZB5cgUNG8fqycmMb+7hvP6//FbPHk3fBfO0zKT5QmG22XYixu2eA63ZS1sCj
MCYP/ML4yM70JSy/NQEz8eVA6w0fVSQCFaCX77cCZukVjI6y1vxmCeQ3jI3SYPQi
NjCZjM1+Ca75NDBT1IKyrMmeXp9qlDY+8Ne+XVn/cD4S4OtnuBCkBachHplOPS60
aU6j4iJNOY8PPtzsMZ0Q37hO0duwtwuQ/HauaPGjc8FZOMXyKZssrXJoUFyWHwvi
hwVKg4flzForsLvbYnXhz9rXegDcaD0UB+T6tGzZNJ8OEhgX/85nz/wUFIotWJuD
ysz5j5hUtCm78qPk6DtQqqoScicdrcds9WvhQ1JZCatf/NML+TbtdvKSS/NHq1V3
gALVvh6ZPBGtbx5LELcb/DaFjCPXMLLLc6dMnclpRwlmaGXo2gKj2MWGK2qSRrTn
4oHrf+mu2jdm6w43aKwsyxbSLJPGP77YA45N1XEqZC1tZS9IWOX8X3P950miCX++
8xXIZTmT8iiW8nXv8W/If74pHyvu3Ac18KLRc6sMkKyMwshHG/CTHN7iwaHEX+0E
6Qn3jpwvk2O1JB3ioAGDHwetknQMbi3WBuwYeNS5sU6jf8T+xXtjBqQI0wB6ZRdL
gfCeqy0TtW5EPuESG1BDcBFTDnwC7HKg83HkXyjCJlAi+ESTYuW06TrNhfMtOZ8U
ppIzG5Flp25otyCxIK3ys9X/gn9cwe92C8nhd3JR26ia/70OZonH6jhfjTbYl+z7
QcZzCggdir0VTObMexPG7Jvg8O00eQMfTgD0D4oEUDBmwfvhlIhWi+zPZehc23wK
tskagDwrubFSdfiVxqlxn+L5GP559bTllSuEZQPw0AUZ+fo//djqzy5ltmB8eXB2
LhVZ6O+sibBJUWuASL8ldXdj3rK2e1xEdSPJt48CFZQM11LKAQ+oDo477r/szEjm
NsfupEmm+4+Hny/Sc47ji0G8Xgxy/bR8d4HEiI1RGGlmsIUNFMM0WixbfY1behdH
Es9lH9+wGs6NljuRYeA1mN7094mAvf0moM6eOZ0QKBvYONxtUxGvM87uo1wwThX4
mTDWAkEv+A3tK3/4xcBaCc2o3b2IJVa+OqjzzUeGZe4mqzLVsMiF6ZxQcI5ucYbY
ncn/hpRZszzPGMvX8VL2t7VNWEP5Ne2cnfVEAYXOl4BhErILfTEKWG1CQyw1TRmm
7XiaaVFFQ+CUf6QJHyyl64bivRtjmgO0Qps0muDY8nC/adt2Ecv2ovybqz2uVZW5
OqtyDQ/N038TBVCqgTYle+Our/mXqLLVCS47nLot7VTXTVDMHHjmEQweosp4oN8o
KIsnIqNn+oY03HsllbMUqc8a79giKsTz71IoPJaXxcyKo7/TWjq71bX6dV4iXTqK
p1E4IWzWgotep1IMRXXbfAOunYkK19KcSgICh06QhgXfva4uoD0CT+cJ9HLt5+Vj
N0ENHv1jlGXpY0oL76ggCZ1LhS7EkdKuHVHEQuPXUbc3ep5dJt/MOA8wHDIjLViF
rcDI36Qm8u8v9tP3dBFOhzGDBsFXbYPj9fk7YAXJh6JfOy9uJfJdxrlaVVPFDwcD
ZgKo/95OJ4PlYxwh0Kp2DPN0LI9tLst2RDwHIZeDa7uBd5hCxuXkOOm771aK1yd7
5kDpL7vvDnCayKtHAFjFe/FwlnGl6NrprVJKInBw16l2RnbsBNDj+Bj7KzLTiqtQ
vSILASJMyZ6S0G4SplJgp9fcjHHUrw55+6qG2r8Eg9VNkedHCcnSBbGm6GcuD+jA
ozOlasnutU3FgUDy/GUoeA1J7NbSUYlQNTybituxki0eGqBFEufJOAUDSC+OWs6s
XOrkPRUP1I2rw08NrHPaZ7xDezYyp3WCVDLPIrDNL3feR2FP+8NRz5fK0icaicoI
u2EN1iuKgla462HwafiOFnnI74KaUj8F4/N9/LwnZiwGtBlQ+QbySDP9lFwRwwVy
NeQHKnt+DALRjnw0oQSg2uoq3pwQHimiJwa0G5AzJ3kGMXh8TJ5TvOlGE+e/xDfc
fq1N62lyQW786Cr5bk0Gw+6sawME+HKmPWPCXVMZnGJ8nay0RauPB2zTcRf1z5GO
Hj+c+6cswA+TaeFZCMoN5lLK/1UBBFs93SUHEyrmrXuhfTvs5CwnP9r0dmr0HMkH
g2KUFXPRD7QYQLMUv0TtfnZ88aj8FkHxrWSwxMQPmh+wOyoiPilIO5XefPJCztws
H++5ycXoW16tFIH5RznM6g+Zb8lCUiC+OTeBMd56aqRX4WC/i/Yt76Ut1EGbCKe9
QbqgSULaV+uBzm5KM3SB+RJVaIUoB3AtoXNEBZKSgyuoI4Dw0k2gZzd+db7DQo/z
vZf5GxVX4t5TxZO/jMVIeQtgKkzQ8ZrruwDRhlCZ2Jgb3pXl2szIuapvBK+p+fPH
4RYRNZW7PrMcR8Dz1Yz7vFHmSL1riO7JZeFqctvWFWEtOThjaNooBdQfbKU7rZI3
XkkhCQt6nK5FpW9VY/9esF0A7ByRasSmVKr9xgZkgcoegDP4aG112HqXZ64aXOrp
L8zgGRVxw6+q5Ne9fTIinUuRybFjryceReU8YZoB5OT9fiRqNheOaTKY5FthwY6m
xC4uFYsSbB9/nd1bPE6yaaUqpKH3p4h5ZchE5YFIuMWFmkNom3vbQ/jMejYYYepo
aR7rDQD4otcSuBpbGXhoJHVHDSnKrrDcWHx3X1goJKr6UnSQ2UTqnDKhB6ubAd/U
rucdaGhMPXZv5AygDSNgQkqe+aasF6uX8XDoUKyurdkJXMkYCeBhRsvG1zcMuOo2
ROnr5v/dx6+Px4FHz8KwO83H9Tj5o8hMDGtd8hGEA0/rVeXfHelJeQ9O1EYSb+IP
FMy+lLlURHnc1zBif0X4F4lHc0L2pC6xWJUxq/GbaoiDtmiVUPkTWFAV425EiAcP
T4v0DagRpttlyg6La+BiIB529/ZdeSKIFzW5LzBc0FXYlzs3TK60KdSAqHl8nW4m
LQ6zWa0/+f9BA28h7+e0lI5vpUqRGbAJSymrMAmY9vnJPux1YFScjXkRP5KGHrn5
efGX1nxwM27FP3xhMqyZKoJfRy5TSIXC1YHUEVkK+ExP/SymeD933GwdywjRO1lr
KqrNEO4c977zUwgGHMsj1yWU0Lbj7E0vsYr4raZs4kJmFG0AKUcHu1DZtvhRZACN
SgU8NMSkZBTOldKRerOdqHKWOhf7C0dr6n7K/DWN/ZKn29APaSQLLrbsmU3l0kBW
tjk4GkwN2f6C+1I/zdo8UQQq3B6iofw2y0KQtSPfy/jTHrdkenzs6nRML0Vd7V6+
M8huGN95hKqXBFgwHu97rYJPc5bjLE1ZjKzfnwutq6nuYkqhGsPuV9BjN2R06w8Z
nv2YiT0bdhrs665OWLiYn+8QsxE8I7RrizhqnzucMreUxBt3HguGlo2V9zTfNoQH
kHUIW89BVgp2RKLTPihCVaNQ2p5KiNIiEMJSd4PdBvQ3usegAgZN7H/vrD38BrVs
BknZaH4+ow+hqL2gZXwxcfECWqRxKBQcoD4Bd+GFm0mEgvJpk33jkD5CE1cOFNJC
RTRenLC/QhCW2BZGNNtGwkEureT+Wag8HGKtTaR6gPXm7J9imufSCWsIh9Mr1EDe
96RlVjlF70QMrYt8EK0EvmOVPG+kFl64V2FR3y46yz1aK23/Xr60fNaL7NyMmXNB
IU5bcRqvlFI0sNwMrNMcEzOOt/uXoFmmdrpdRJe65IwjW4SKGw8APAOthALLWGKM
B++5my8oI5TNae/2YSf7+kEp3Q7W7wCrgrR7eqto/Ukek+IBleFYGzNvo73SqwwI
8twlXnE4tcUcEH0c4iNE2L9LkNK9msJ5oSslL+YVYj6vwHgGmKbcDMYQPv8fZSYG
dxI8Yxpb3l52RaRN04uP873Brad9g1JS8xo0nzuHO4F7Cv15QPtZeYJ5P7aj6jDh
FymItt/4djqJZliNddyPAdYaV1Nta0b08iNOIxpYgOTlFUDnYPNg1bjVHyMcaM86
D8X4A2brMv11799gZsdrvwQE3etEjtDV3DzQwcsRlp11BArBbYPr/BSU7Y6TXASv
BHOl+HOLdJkvmDQNEHjVGwGRhhfR7GY7T6nKulJGVChdNqMAxxGOHWxPxkE1AlfS
SEZWOAUOrNh83hnuQVeptPQaua/4EYVI5pXT/qO06ZVTxQZIvExLb551dnzuW5r7
VeUWOdduxJlii1EHZ15TzroiMvtIP8zeV6+xi/SHzjoPuJcRjH4gEkr6b0VBK3qM
IQrllooM3tzpXg9st+2WO7dH1HVaiefS9aviyfqY3e2dju/GBNjP+qQKOFetiyk1
/rZ4NrX+kGim//Gi5dsvQO1Flz179uZRJZuy3hPzW06hbTxaw6ap8AZAkOYY2Ks1
O70b2Z12W3YqnCWMsTDnI//+27Y1lgLOOHXK/nhhTHiRfKxdMZZkCt15fsoY3lpW
HHl7TWNTAQYf2d6yiUpxZXacCSdT5sdhPdd23QjNSPxkmHjCnTRslYpxVg+3wKyA
DSev+DDj8gm/ER4m8BuSQNGtjK4sOJgHdSldkZYldyZs+024aCYny72VkLYzLo+y
PHGxqJxFOl7NUiakCp1+sZpn1Ks8ICVLr9bgVUFGAqJsCXQ0P3rdQkBEoQ/r2X+w
f69TOJI0ebRL9FB7542u2TLxrxinSN3FSL5zWMISbgxGPs7DeCMRU6Cz9J4mghnI
SmydnHwXbNNX8LYlgS7m5f9ipHh/4HTSo3MfDgkEugkuJylLR6WDI/RetiqRs6Ap
8OLwFzBrtybxe8vScDK/vIks8AO9TQhlDufnVAVVK93exzWL1NME4xpo8Ss8VeTQ
nO34ZehU+XSqYGUcK0CiEdcXqtdBMvqMoR+Z168hEYu4GQQ/bB3hiBSn9jIbWifw
5XisabzTFj3fmtA8xK/2rLNjrup30CXhDw7oKzjbKmw4nC2sjIXzYOO6UkhWWXOu
Lh4OkM9Xr4wLAOxqM9t9LG41y8bayoeCwJJD3UnDy1n4rYsJby4K6hhbGJJY9oMN
o/ofvgBa+6DXaQSQBmJuXRRCIupYQQOL400i14NWKH7bkCZlyj+B2Q00zhNuqnfR
BQQl2WBZWi3ErbAVPR8RCEbHchZkHJM8I+OE+W3vwi3tuMPQ/zj5VWRS3Mu/omIZ
ZZeX8llAwLo/ZY5cBtYFXq6dMyaWfVW6vIc2RwrWD0o5fpD9vq9IgR2HRNpUIXZj
tsOyCd01XIxv9m9VxLVV6QlOyDf6xu1eh0V5JkcAHiGyutli6g/WC4+xMYlaYnQZ
Yb3nCLAgB6HD3Sfswysie5UznjhsfoX3rVlFTyEHkx11IJZQ8Qh436NrkWqmzeq8
D/QtTiKDHTA/C9wsjfzxPW8fSVoxqfVRzRLQRj1cmWrmSfoEPS3OdcDD5qHJXo50
qwQrcHhFRFQfNBJJtUkDACcIxcRDL068Gq+NzV+QRQrk8N//wYpVTRwUtGDwMJtt
RvD6zmZuxUvaLOsCjaQ8eOlnxNC6sg7G5uv8jDCw1kQ0Di9I0rnG+fjaZiQv02Wq
PVpF/dXsgdBLB71EtS+2lq6Rjq0fIm2l7+YpPDpodVfPhhKA3ZJduMLbCR4JACZr
xqpFM+JpzZlPU3CtUS3IVbVR+fMTxKXQk8YqSPWGl2b3tmaKIO/2W1Zuj9CWwGyy
Qbeos46br6rFfztmMzXzQtmNQf96GGdup/GpIuqxJuSATP8Zo9VOgzlLaORjCsxC
pg1LrnNYf5qUiDiVSFbddMcDkJfESB+VoTzBjaUl/DXVmomwsjZyVwVui7LZW7iL
D78DoyIvPkkQCKxGbnZwBVs5jVnFPUlOgEFdueNzpRDqQOnmld45+cBlmJr5vMe9
IzT51o8/E0ZzXgM8UqZHF7SAFc7ToA5fz72wJTQCs8+9fCGGBjpGEwtBlnRbzcT7
4MQhvCC6BJvz+/gimvdO26ecjB3WHsBy5cSU+QdHXnHzgmux1wyxR4oPXFpwz49H
NAQ2UngSRpRXPNbuTgvBbq0Q8e5f2ZU1py/H7sZEBO0pT0qxzPAAKU3+IpprX4mG
GVHnDLu3ovJW02t/1doFaZEIwhZdipWWR8L8KOy1ts8C2OEecb5dN50Eur8TfSOH
FMP7M/nX4jQU/6O6bf4445WihIaBkFnhl493Kwth8KTK8vFLsxQ3l0fHqCH9fiQo
0zvu1oyiK6+5/UIca848qk6DCK3b++kto8TcXNo1gpwDRnBVmAwC4SrqtpMGrLWf
VbqUz8ey3FE90ttWE31xhY/R50QDFlah0jNuBr53oD9yQLlo51PQfAd9Rdt6stlZ
yzDxod6QkU5CWcnHSpsZO4igu/libAKMsGqadCO+FIQwwsSFN113+Am0R9TWV66d
9fUh3yAvQOVbon2oJc5lLRPk61bS8EqHB4EW3KjkejlKRqTo4ni9s++cPqITgRmc
TQqNI5UXkOX+4fjjEwknkBoeONxouXY30tyK6FHsqhUkMmWh0V7FZs+KpyDgsaqO
pbaw19YkNBZsYparpx2sPeYzg7oc3iQnkc7SJ8v7rdYUv6VKYJuNBx6kMO/C5szg
mcBaA0abkC3Z1qHbwadKsRUlLkL/uzhBKqLnaw8zgd/11wAXsgSECQaCZEpZ/S8o
e67/fu6QuiW84GJJLUBeQkTfSI7iliCRrLJOCpAnh2p0/PG8VzqHqaSO7sXHzewc
+78679JBX0ayBsww+uHq2tLpJA/vxuIBpwuMuthXia6s+LNpeuUpe/RSIi5UN7tH
KUebDQ6AVo66VhrOh642m/T8Emwj1AusG9D1Ica/KN55IU4wrPyP2naFtVgPHFrg
/Hv6c2gw0dr+tmavpvbNUvLIISBk7I/GXxbnBE8xqotlq8Yz/MolYKTDLsv6JjYW
g9KS/LHHFWRBinuLmgxdHuZAvef1u7zbiOJ3pG6lP4IYQKLWD7dYULJj3+vehB0k
cxbbAZFZ25vR4zPtr5IJN8qICFKf/SzJtRXK2FkJFp928TZvLqhFdfNIOhJA09AA
m6z1yQvrILoWwIHl0qsmAs8pnsFWDmvRLCB2IAV4UXcIRIMIqN15mJh3ghbad7tZ
jta/5yD6kIHGqaMBHSHRPdZ3JmJR5UQ5aKr9TNYlcBFc//kc66qASqCngKkbwrld
Vo4dtk06ZNkXK2L70T4HPEq2dBZvOueo4L2fXyQ9x/JkSjrE6w6wjdwflzhWrHhQ
mky2+oT0sxNsQRnX4EuvPmpRyaLlEwy5vrcK/jTlkYl+iX3JtsMbiQK2o08S9FKA
ev2EqoLsN+EDjBCAxS15aQPt1+Gy5J/YRfyxxKY90cD0O5ztWJ9Zt0ukCVj87WE2
io22SGf5bCr5NX+mv2rEv8AGlScobFxel3SVtDwA9sYWrpdGzB0NqQJn6GtGR0m1
9xKTHcivLdg/ociFDuPqC0CbLrR4WrSjwJ3kFMtbiHfN9Uex+IAwSDTJE1JlghvA
8Z/I8VK27qzwTDyAwSddk+u1djG1AE4rReGHH2qIi0O7613gvKwCp7j8F+cFp9ls
sidgOKkwWk0ezHR54gWTz5/AJhS6UXg0AeRLrOtZWA9EjzIBGvEgiQRVBH9VJ9rr
YxcYvB3WVLIgJb8QNT41kXk4gf+jq1RhFPQlWYyORRDesJYn3jaXSyghpB5mTN6a
7x2Q7llZZQu21XkzqZz5+ELHZ+5E/mtyWjyXhIGxYo1yPlhDtZV/IubPgj3cWHCV
mtPkF8BV+UIxGexpYcWB9EOTHlCzj5nU+QXfb+/s3qZEnQr4HDTsntsKRoJ2lr89
R+cJK111t915AWZwE4s5ZpmnppTy73pxenkzoJj+Pmm7Mfim2Vo1GX/fcOFHTCbV
gzRf5VOSW/EJcgoQy0mS9B5s2SbmKt+1Kmfc7kxZtGWin27MuIhH2Xgx6LJN0Fn9
YpPMSvCCXewBG7t7OnmYZtCX4pfLfj9tJgSFy16QmMESQ0NlOfQIPsIYWgU1MY8w
cL8tyQcJRkQcJVTHfVq0dVMr/bBS7uubXK+lbYmGbmIJqvPL/Kgr46UlcKEAmvy8
EwolmYOfzX0Lm8de/gpxeDV/XvqTkqdl8D8VQltm0BuZVKQjgESEtL86jgptvBwj
0gglW9+UR279h2aSKKVtIFy9cwAKQExRFhRVrE1Ov/zWolZ/1aSOqu4g1oy7NfQP
o8iD3JWYZsHB0s3aP/tynHKACSXD80lyMSRr8/ugQi3/NEvrqmxvT3yBaqnHqilz
XiOpjF4oe74xwsGNIO8LG7NXDoAqB7v4GoOkvkfn1pjtWEXGtRW7XrBwcDrb7a7M
d5m4POvDijGITHv3eGnqrA0PcmZbUj2s2WC8211mNFiReYoQMHDo8VjnLaLIEXOQ
zaeNjj0u9vdokfJCGH837sMnrwNONQ61oqLe5aCrSzXmA2HeEWPV9H53I6DZ301r
ZHDf+yDcv1Emh5WEtWGSdedoeAi47/poBlBKxS3RIFuhit+Wg11sTx8j2HPsHOq2
OXD/nbk1aQxnkSpADJux/5ho9fTDk5rIemq8nbbWhUEYnZ1On7zqKVV2bv3F5rZY
DXM9nDMft0RbpR5u9Glkrff+3LroqYgv7K2+niDTyHppS3UwSG3piAdbJySv4vRW
TjhcJZvss9U4wMH/tm9CjWDuAov/I+qff+oWrZeIbaNty2DLM4cnTkTqvh4EsLOM
wH1C2WTDETw6CaLmuDjNCtfFBesfUbWJ9bkcTz5GTvD6g6AUQypvdoLJIVIwRroL
zu7RdSjsKqyYEBCwMLTYiDDBgb9BEEG8IG8DWPeqLfWV2pivZcbmbGtst1cGuT1a
svWDaLFDgx2bsaUc0AP56TyH9gJqOTRny8GGnfQ/ELlT2uUE14dHKxfjtAFcePp9
qG+DITffSobeDjfxtT4xl0p6gOdbGbs4wP/2enU+j9+Ouvn1vaFIQCQ+d4oHUmyM
eJKIWfVzPQDLgWElELPwwCCeoY7nbpt0UL5/zyvZZqdZ6lGRbm238CSwUW7VztRE
m2PjSi76quaz7uOfrPkKz06COets4XrsgmtcHmUHJ9vgxGVBcTxUf2yKyfk/ASCi
3nprIwPnH8WvbdxzKcaAKrcnJdhl1XrWfzF6/kSa6dD8WT1g5M0CctVO2GY4xN/g
veRZEeLdJ82m/xafyMMbbUwXyxJjEjMnT4agSP4Mc3fc/GyERieSEgmm5sSXZ0ph
EX5ZZlqOyYuiacKPQtQKm4nIEeLGSBB43YVK9uaacELS0gpDnQrd8XmHC7tlRIlL
HaHrhzM8raWd8gZmVBZgkO00z0tczL42mGvxwS4GuW2RoL7jJpYRQ6+e/c5uXOtI
ChapYSyMP9Y6W7jn1yfSJ/CIIPrUO13ethApPzx8z9ru5VbWzctE4pwd56FnSNh9
FxoZlc3yKAxfzmNNeOt9FiEUQ9hbYzhXjS0Z/FmA/lJDsmPkc9LxIDboVytUpzjc
MjQfUy59Xk+3YGRzVQe2hmUIhLTQibYe95HrCR34mgWn6JIGA2dS0zm+nhEcE5tn
wxwbv5DqLpNG0rdIjTQMLynfot1G9Ydy2FZcFZd1s5jQytzTgEekJMeuZY453ofa
NcHiYywb2Sa4gaDrK9/9eohMq8xi5VBCDwksEjAaGX4bGvOGWpZQNGoILZbBOdnH
ao6auq69zCDqj/hVFjF1tmIwaiH9PkY7m9xN5MJ003zX5A9K70KjJ3Y3LmCVv/bI
OMwL4iVDVX5GivQRGHLxuwPrS18G6tnenOv9kVcUxNkQc8rnE/4DHPV/lFQQ6eo7
Hjm3CNG9gbOw9dl+XwqQGuSbvueEe0hBX+cY90yb+y+AwiWx0X8tVSQ/UDYhhKk1
LG9qG8mdi8JP4SQ1xP751yrV81q8wFEiaBqbr2yYbTeEBu5uijbCRSoOYTHYFxtR
qBAskHt6ZTAD/LXorejEF/AqtpoZAWwRXhNXvWi2GFIK7DbZPvGOM8iO2LKjg5xm
fo7NqpKU9KUP1J/+nDz+hyUPsSSOCWY4KTSvYobkuverOHBuHx80fd7YvbZunQH8
9KrhJRNSrHnqTU6GzVholkiFaOek6BSlBIMkqAddyUSkMcQ0XH0R5nXrycUs+XKy
Z6RrzK4tv+iYa9Ci7+rHPtsrTcIe07cHtiZ3jpSVBW5+Z95b7DgvoJhD4fqCbS5S
cnVbPzY5UWZ1JJ/MchPSrVWOvuEdW9/EITgxB67LQo2RS9+cB1qg7/lI+j/fRS2u
tpLwZoItTiX4A5fJISCGJtCJvu5RMw0mTRm8F8iC84dzmQFjSVVfi4uGFff9You5
SNXn0/tbRA6L6NfYlNIcGcBzBJVbW7gv37yyvnscy0qFnR5Cz5b2CKm252lFfB1z
KjR8mN6FOwtaG8N8/PzausSm5OHmjOGbLCG64UGP+YuS7VMlAioeZd1PcDYE2f2c
W2nIkxiHEiC20+JTqxqCfeZkDyx3JYUZqNEYLHl/W0ir9qWxiY0xK32qODudMyGp
TSVIrekxXsrBApmHiNvhdxzv3nEhdZjMkk9GzqW/brF6gKPCw6vDHA4lVcQhhTv4
a75rL4hmeDSG+GkGLyCDrJKr/P04O9rL4iWtBMNBx5ryctb+sTR8gJgRkmlhtiVd
Uy8hJvXZhR/+8jvCewZUbgt+ViZ7oi/SKoBYMnhzYw2DXr8ZlMqEoPZutNic0Ttc
tlo9eUispARhGPwqwYD96EXe/7I4sP7FOOkIgrr7o9TzS+To4B1bpa7k32cPu676
QhNWW0mxg9mBgMUYvJz6p9JQlHCoxQOqH+F1Omv8sLZbg6oOdsCvo3TQg2RcRP06
r29exeJC2/g50NdxlzcCJbu9Lt2X/zA46t13OjKrACd9Pe0pKm81h3KzbvcBgB1m
mPjaF/OZcjMHtWLqWVWN3KsPD1W+nv1Aergilf9pXt16kFhC0OOfTr0/kPjOOzxg
vRGgt4+ApQv33nqq39IvVeBZgvtaezm28d5G4JK5+1o872C48rn6xLLB0jsR+36W
xkBMteuYXb5XA5/5gLdZQzTZJ+UsXPnYxZtKXLrbNjZxvFEf5PYg1nMM/dYij2dA
hUrUwUQNQZA9WDTMdcaTmvNmn2i1soP8ocOT8O202fWblADHCXlR/vLB0a7kbtEP
MHWaaWBsJs/mRFFZB+8OoUnQWr0gKpREz6VOnd+3MXV1nA22Gs6cJ4oHoFFw5UOq
QtAmh4JnSpzCTglAgOkF9w3YCqmuOL5ia5pndkFQ/AuehelgMYeoewtU30WAKjyl
U7AaeksAw03dEKWg1pT6kURchNjL8yRRaeiSMFOieX6Ec9iqVw6A8K9sySJndDf6
celz26NShNt0Ri7Dc6kQn5NcKvv4jwLKAFAmlzNibbCBULyjLYfu0gYS9q7wQJ8Q
LYoXhi6q0e/4BZXGIEwf5PJF8ADXBGG0BEKw5eZ3bpZ4WUxKCUKeLznOE8VAkIkO
b4YQzmxJNJS+2rjsRcvWqZwUpBD0wKzDYEM6VmYA+IgFcLHKtwSFLHrgeju+mift
oIN3+CTaOuHgUbuIoz/0v/+1bBSf1Z74Toi1LEEmTRMaJ6CvCQPBrEhE67x8ir7k
`protect END_PROTECTED
