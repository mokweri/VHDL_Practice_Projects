`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNIBhJW1bS1+0tYqCyM4M6yIamYxWhNRYpmC/cmvmqbJYaaJQgh0mUgYAqla5BQn
wGVFCT9BALogYvztIqyQlFbgjN7GyGoFTKT4rm3MB22+N3AMDpSiHBTo/e4aXES5
V8/X5rPyfA2+jfd9Rk1MqcuqeqcCeLAzQrt6W+hARaLw33wT/HaFcGxr2+UxLr42
K3C2eEzfqUoW1vUM+ZJtRZNIZXJDMWRTiUSnXSZbmGojbtSfmXpsXlAMU8bCZXb7
KxMHFF4pykxjFQO3cxTWP576H4/t+5qGRMaVobRb7e7vDsLbHXMvSFKXM0QrI6lc
+3ZlVHCOKAGahhocVY/gt6PLoZchmgHPoYY5FHAty6HPCr+LTI0jkOtakZBjna6g
6mPpf5PFu0f4zthBE5TDbcYbFdwZG9XWO1IQZP3RAD/ZXYXmhHuyp5pG9GcoY0zo
Fwa2/xi4BCXYeHZelN8e2CtAVrh+qSgXDW2ilpYcIs5mbwOR5ICaQZnuE9jERyo+
T0oOOYljibXjOyqSVNpKrO3ECIs8ZY3vX1/cB9owNIFYUd1gzkQxgPrlABsQ4nuc
tBcfrSdo9UB6nBN2vxF5acuPZ3sl/0ZdgQaTRyrAsGnombVjzPaiCJrGEpsiGUp8
OsfSWFyjVntGsSIg3d1WBmLk8v6+ZRM60IPVCTnKgHm+0Bh8KAo6WvQau1+iULvc
PPN2YGtcOliQ+n6PKN262zZbxrWTP+TZ4kIgD+GxMjIYamqOcPOUa6d+b5WRdFN5
PlALzo55CV7id58/SDnIuzW4grlmBa8uiCmu3AD1lR5RJRr03wA/4BWMuzTScbVM
xxVRYptw1DvkEoeOp8sIXJb41bTlYlzgZ6mAaxvtIVZW8FmzYI/tZx9gVvnBRL96
PJwyhnhen6PIJP7PKm9C7do9L2HHQmM3eAOAZFDEEpGe0h1y612Jizn09d9/Azwz
nOoFUv3eJhWOuhy961OI+GfdGWN/wSH6VbbJTC3Dxcr+7dQyhqq9WVl2734y3bXv
V3g82jaAtUzjFPaRh2pvqvypHGFQJlzhfw0I+GFj5vtOgSpEI5/QPC24C7F3A86F
ILw598MV3e7aeLlMkXorj21CAo9MuAXjy5uBAfanvJcOn3KYWf7eCWlgAWBMm1hc
wD+VPdh9cMpTPjFAhHNkV90EuIMncckK4pyKSaqIN6WExnyuwXrQe+cLugqvwclI
x1Aq+m65jQkniaaBfc0rVq9STJXH/CuZC0Y2qUhkJuzieZR2fqziaXOhZeinsTWK
LL9+/vkRAzXNhKAGHQKuQRYpsmynLOKRwMg7ZFU1TjFcVXBRAZbNEpmL7NbB0phF
0xNOV7e94odENL4i/borbkfYZZASQ8LUu/6PShWkvqz/K2e+zhz02QnbsaYRAIC9
HA1aCQUe82vcOqv5ppa48e341/6gVHRT3oi22TBH3QswT6q2qLerEhrJW+5NVKEh
`protect END_PROTECTED
