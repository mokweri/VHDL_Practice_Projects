`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHGGnmmbvfJd+RiGsQItoUCpKhXj2S9iRLskzLl2+WLX2FsJOcRqSzeMNRY2LgRg
TFP1iwBjyaigRRRFGQPoWJxo/3493sWgAm9QJhBnXAJjzl+k/smYSk3MBTipgLfU
pwvHCsb9f798CtEakAdYSnM/knxQgQosm13FVRo04G/PjOjKfumeecnko0yRgfKo
FgUMWgKNK8rwheZA32h8ZS9OtFZPAPnkx2ajkM4OUlgWW6TMZfCbJlaonnbqADIV
Und3Ti4qV9QfBcUCVXEdsctaml8iZ8GtST3AHtiVSWoXL2XqZQ0vqSvak7l2xKT6
rrPfIuc/tabb86nE2Z4i1ip+T/Uw5h8vdw/HqzPpvscK6DlwAtt6noE9xpsigex1
IayX44aH5XCyqR3yGnSHPu6rhiDxb48WWI+ytNVcHLqVNDDrEDyajgQf51AzXjxj
uENubHrVdfm0tT+bnKdqwL6rb+gbYYCpLe0vMe38xK7m7EhhvSSJo63tjqrWwGpp
Em6rhLmZ8ejVfZJ3WsRWOHUVGJAOp8SLkfAxgkz5/OmnJRNrA2MOXXf2RvmlX83d
nUlLn4Hu5jpTvBDy8yqzQQUAMRBAeceJZWblfTTPru3kUwyNxouQf9ecDXZ8eKND
gIcJUwe0erg0XxNOjcsE8TPKeaF/3EX5zbuhc0JFLoDIMsy7EMDiBVaNYUgjwx5y
pnlkDoaiwsuLIEAPXspuwJTnXwzjJ9PZCgVilgvPw3Jf1nppidh+EOCv73bT/bBR
g0i5Xag7ubhy/vhBEeA4RzU1RdokdmPgows9I3pA/7+6FZITzt4i9V/QLWxGFRuk
xcLfQrIhF9UgEwJTuSbKo/QChiW8T7wPxqv28ZnNDBs=
`protect END_PROTECTED
