`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sO7r+6Dly7VdLkKzHwrqfGeIqZ0Shg32CVSjBPGnyrXR4thk58uvrfb51DoVJuBc
SyAin1g2SA3qd3OPaiQJM9N3vnZq9JeJjgu4L2cL3+WmeVx/QWk4jVtTgTYyqqYj
JHpcIilAFexoxCZMC4eKC6p7JB7pSpRBPYMUQwR1G0ZoZvR8ePN+bS4V/Qhi1iAU
Y6Q3brk5XhP4YzivzJCoOF/zLpowRUw0wRScUVobuQ/EL2YxJFZei4Vk4j5/RAxT
jAoxaoNRloa/0gnwNXp452n/qV8WjYPYfciYQDSISHo+KafU0PVyJpTrs4WD3XAy
sBUn8RObefYQUNu1KMIE0TCTxF3pmFLAttvBRPmN6Ppvo4t9AkU/0ujSmJRtwwvJ
CPRIa1+u48ZGarm3IAf0sk837RJHqnfanUb3+26zSQsbnXLpqiO1UstUMiBLGs0B
7X6RdhaCGLidIG7wsa4pR0FvHWzn6cWd9o/vn+e6+2jN8BNULgEKviuDrRZlf3j9
klqAfIzUQw84t1L9TjozJ3ZMZQZmMF/JNmK2mr92Rfz58QpK2eOqy246saT68oj7
yaxiKhcExNfd2KldH0oXDcip7w/tvDCDMbKhsitaILJRWpGzvGGNLu8/JxVe893n
l0UrPmZ1naFmWW6LD4clbN3FBSbWtXIuS1oVyZFhUlSX4A/cwG66Fy1V1qHlijQ6
VQz0Fspq0Z5MWcWckSDW+oYCDQmhI8doCO4DvXMAlsZbzEt0B7nwsH0ZKfpISmLJ
ZHmKYR7vCdMVVL4pBqgL2e+8j0byuEwJbMTbgxP08V6HmPdIQclrJHALCfXS8CKs
rd2oS+X1K6RZ2NNfK9Q5RA==
`protect END_PROTECTED
