`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/RYfDGaTJ1YYFoZhoKwHnlgwBUSbQyvqSoWrcQpHAJeZdiRqERjQWmiIEtSfG0Z
tsF0hemF0cYznsN8dTGeVDvdGAbQKqaDXyXWsmqlXr02rsnoN34F2Ky/saR8lxkn
gi7MthlpQWmCjmf8iCAV8P240BEnepw45vChe4iQ6ToSylCzv3/EsPyI3hfQwl8t
Y88oSk/0ch+OK8597LYrZndFH5hQtcJpM7eyQEIRjApvewE0X7XBEbi8SxtLOfkl
r9dLS9hO4/jHQGhLGdI5sxGkRXp8WSyU1C/vrnyu3mi68Kib6rN7K8kk+vG2EFoI
b3HPl5VHDzZPvUyv2eeuFjNVjdBbE7Y9yLwWGH5Y7vTObpg89GcoT1xseMkfRatX
fU6+EbQkdI9HK1Pv/dnwpc38TDg1A5eORPHHlZ2V08pwmp7D3ZTeTYOJD+aWkQ2O
8NSba1gcH7w6R/xqIQOXNiEFa4X6V9gJmq73faKO3ax+Q0HcXhbxwlOOlBQU2drK
uZ0FirOpR+BGlSCfgMqZpFb8j0jYA5LjZgZLC6n0tuoT66hqjw899I+oqqIchSgR
k/go5suxtpdLhDWr7FVum5MZ+CkKBLBNLHYyuNynJo7fdi5LYmxeY5gq4trx1cPF
GSe+ls8LzJg1YcI7QRQyNti54v3Fznc1gXIQuDaJLXfRzwtf43Wc5ZZ3KL48iY48
Mb3Z/5SZMgDcNrcS28B7DUwgEtlVkWsvrMl8uX8xz4i0w4E53jnHdtZa6UstHZH5
0yucb1n+ZEqRkavu3gXmP0bPJt8l//8WE3v/x8lIh34uZpRc8naQb6Fh4Od7LHHn
ThlC/6k8xC0cT8VL7RZBZpBNywJPXCXtGAmFYH7NVj11W4j/Om4TBcOAZtlIaTU9
cx9RHaY5a9ZtiSBml1ZbEe1VVzGvTgez9sjlT6TInmBlLq6KvG5gt6tjHHYj+qrA
ChuoiPmdTVV23EHnv5QXXrLgBDhFrgteU7SfRPaLvrRNQBCHXYNt+LUZ14nl66+4
cCMDfQh4RfBRJCNGIUsqpaL63FjR2iDejYVvekiaqosAEsBqdUiscwMaCdxAjr5M
oxmPfsUND0hH+s0NB7noSl03v5HWkuMxAPiebIUzMWRgPktLDoAwvnhv4XkT0vyf
jCHo/vdLQvbc4du9x1yXIAngWIuvrq3ghAD6aafQcfEHl2AO2VQ27aekGhWRkU2t
SiA+MjHAyhCIfofKt/B8HDX3wgQvmXDJCNHft9BUqsarPEWV1VwURMX7Ih3COshr
MaGegcXgKn1bPCnUNWyRdmI+6Rp+4LPT+jVAGBtKJuJeNfTAgoR0clJHzTK6GXLg
TjpAPCNyX9xgjDoGxzfn8jNqE95Dt9b89+ZHm0fDXU6vne8u9r6KhOzcGM5ZDe9l
WlkDBV7Wc49CDQf3E8qgPYdIokfufWenYcsu+7xIVp0h5ixqN1gz4h+j6V8+g4jh
n7y8sLl42LNL8srE2dFN9Fg/OfjDziL4Nekiems000GdWwBYvNH7Mw0U+g/vbDXj
yin876d+aJjl3SxsBnNdiQsQ1rMZw1zOmsFjJz1sowIfshzJNxx+hroy7yQD6hUb
+geGadMpCp0mBu40X4I9x4JJ0KJtpipfR/LYFHYhBiV+ujDSDG8rJTu+ht61GrqJ
lI5MzfcpYZoUKt9m4RgxYZIBIdigJVGOeAJMAQNlWNgCk3zOSTMmwqnUDdnIag9b
hdqxo79CgQKHdIjnkl+I7OqCtnc7BCLxMINd8UplTopGSpGHBYQ9hSs4VvdVSwc0
3WdbI4E6m+n+JdlnsR5xwa29NwBExgHQLCE2We2WveXb6ZeNoB/hkYHe03Lc5a8N
OJP1HQ57ZEuCOYVTYvlCCbtoWq9xaLYSrf5wFEFX+/AkodOdTvdsWerMHJhMIh8o
D2pbLQ7L4jo3mp1KX6fWTOw1UBxZbDP3CshzlWR12DQ6xj2gyePENb0MTY6ky+BU
SGEe4BG1v4O39tX0/zYS7p6f4C+tvkmqI0TootMyPGfCdKoDGakv/dsbplp/VuC9
jRa7agba+nZ12Ucv5QRFAoIvh+FHFwKPg5ofUd1E+mOuyyOjFyNiEXQwPm/8WezO
5B/YFcoFpznUyI2xPyyuLJCdhLVoozdCUdg19RuuHvVvOR6c07XwS+DTs9kbyc2k
IQvlpMi+QWic7Kat/rX2Txjwc4j6wFu6H8F0AiHkc4Ibg4/lYi/PlA3pYdLIkVG+
xW0uTuIEC8n8NmiM0FCNOR9ipYYBLQzz3UhO5AtECwwXKo8O91o8Ez8vf9oAB1zE
YGLn41e4mj7qo3Gbb7JF5Cpg0BfewvQtgUUN91ckZyXq9KkYClTZzxiJ/AyYdsD1
bk7hY14wHUTGYcGuqKu7g+bEAzLTqJ3gvyp3PcZsTMPSL32v/kImI0+gVWs0nJRt
BdG6y67DBpf8msFwPhpCaD2ThMWMTvgyRoX0lkUBtW8ekosFMH+JiM2AfD6ynQJU
YESpOMPuyaXqz5Sq0g5GMIG6X4wVUaaxLYNIRSR6v5Ae1LwPmyaSGPOkCm9KYniu
4rN/B//LLpRuLhYdTUFqLb+hIL0Ctj8umkba25GcFeTcv8Cm59HVYxm6h62KtHhN
++sTXQq7H8KcDu6DRJSnziOJm/SJDlsgrAQI0ypIpxze/R/A2Vuv48Wbl4LzYEjX
5PAug5kS7etjG2DloAwbVHqWIcEV+doJMedNCuEg/CGQt2MQNRlpIEpOzPOYPM06
yY++PhXAs82aLbMCquSNGOoM6atxNdt18MoQ2PTsah0lDGWIAKRkEOUrQsGMackb
NSj2X8KrkGV1FoCG08V6T2MhUrIhno3fKAoAi2RqU385iHPNdza24wkpJtmKCodZ
KTMX6B5MjZfcfL8PwLZqSyFC4WZPDqob8L6Iol62KkAGf4NQq6XYDgh7+P/3+E4N
4YHW7yD+SC4NRetyBW6u0ZLZLU/G2B2kztXYMoXakPZtO1Zmajb8PuWVVFxI/9di
qV2+D3iVdTCCoePVdEFZaWAwN2qXH308wnUmipexQndZTN/IiEWEhbCq7XSh7QFv
/d0PE3Cmmwlhi1tEB59UjoRmIzRB5OXWy4lOE31N8Pt3XfTdc2SQsTKC3veECmsL
54qg/aVbuDwRTttYD1xqzRXn6xOgsu0RL3JMLofpFFp8I4UDeZcIEj5+M+UC5Ijc
YHGufhAlHgHcA2W0Cu3UmkpLW61qj/OgmRyNsxO71kNkyzsa7BcCFwtuH+CxRhFn
EV+GnowIQoMxk4Pk6KLDDMlcAKyHMJxGfBUW2gxhSp0chW0duwFIGapKEhS0DpJ/
sCxsfONbDZSLsEdKM8grQOBuLEWffgLoblbcKBZhVHVd4hm5bj54vgUGIHs4Atla
8Guy5E466wXpx3fBASVBazM6RtO40v0uVKiRoZQa4Ig1Ffdtj7QS7nphUHYHZ7Cb
9BDq+crI3Q3CgZIFi8kxDyUzQUk3410gPr9ERWqpvRDwd40aNpmGpyyrOtglyXJt
pvIb/P8XW/P/OlCwOSxGkg5OgSBHAE3loUmzREOlA0lhRxOWrIeDAtlobA61Vu02
3wI15xgP077UDXsVXg/1wP6/FM6+tV8dstyLskeKld1e8l9Rvjq8p4FHsE0WD9nn
QApF21c6j1xkn5SbafWu37VjrfFqw5oEN9BX43PpCkoSc1hKk6rjWKsdNQfBUcMJ
ki2c7qfxeTe+lBBfbz4OK4FVkbfy5wSIxNa+a6Kd0vp4EyG7yLVO/HQ7LbUx5nbK
2TF78mNbCs0eN7pGkB8aBb1WlSTASQ+vRRs6dpa5x772ri3CJ4vAnWMJ5Oazb/ci
HhmX69gsOnyI9D4+VptsL3w5qVFkrL0OFuMTogCaYIdKWDI5FJbq+810XdOytnxg
U6/x+x80XfCRs2hncUtj31IlZcDJaHConSj0xj2YzpI01vGJHebvAWx/cLrH8Y0G
uzvmHMX/h+Rde74C0iaBKbjew8h72KpTtT4cmg40yE7KzvO45cnaz2TM8Ez/P2si
bB+vnW9pEyS0RK4eX/nlLbnHy6HhayxB4VTEZfSYlAtO91imaDE5CSt1jHrh3xfz
IFK4uYWCjppYxqBjEsW3vJua6R+u8EzZ+F4O4G6hHMsGQwnAxQoJQFcJpf5sADrq
MTDTstY7f58dRbBdSKU4R9zEwCevrRwoGxUIPPcaKAdxkLzoxzenSylvwie8PyLE
1Cu5IiBtol4UDX4QbuoUD2dW+DbQJ2lTtJl6owMLCQ1CVL2AYuzNYe4aKpejDwqe
uKN4+Mpo1rnR7129xFMvfXVhtrBPt9W+pwXAYbJeGZ3LVoaVp9LhFBUvkQFHWnrD
CJTopvVaEOsNk8fOxaTCCOTKOosUS2+W6zf97WA049ugWz4NdCpu6XBMM75r27SX
zwR+Ot2vgJkxr5MOhkLzGTNceTdREdHKr1SaQXZbKkuwd38mvsCiG6W9hSPdyWRo
WuHUf440jZbYk8exy1MG85NcSGqkxdzte81MWvFvDEHygtjnYkocLSCv679B2sXD
1/1mCCMu/dg5HJ+9O5NJpw+C9g6lE7H/ylsgENJTZY8xW8z6uLsjNDMvKEF1yGIY
`protect END_PROTECTED
