`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gPqvvaTtaQiUX0hVj5yt7m7+sYdqRtuDpKdg3ngYBo5lU9/wnpBGiOtrrRrS1lVs
WBKunt0JfayGZIysnohaS9NOkVVzOJz5yBxYB3QJKkmXDDyQ/Qu+wVWye4mZPb9t
vHsrQE9oTedVcTkz4xfLyMJEoRqGPX+m/OfyQuY2IUyKxmqDdsjukgbqHxosaH6Z
PQY5DFjh5YpopcWhSU4WoH1MlJ4t5vm1cKwlqP6q/19r6DT8DIaEu3AJsVnxCkVQ
Cae18z5KyFoGiAeqTB/wMLq8Q0bZFnwhDjBJnB4IIFX28W9VQmpcrEQXBgLs1Qk9
RjFo3mVdw0wz5s/1bnZBY9Rs5RtO5PsjYtUyS8EEy8SAPvqZuUEua0lIONoQfyS0
NIwdYTwlnwdkjBj79EIpeNi7ZXNqqNjem8Ie0DkVkuz/qLAMabq+zqf8ACHXYiP1
6d29tmrMMVpbwghuoJb8+E8JFt05byLgjk+qnmBYcguj3wUqoCVTTQS6SwianUNM
TN79aJLgvl48OLjYDtZCqGAg/3St/klJtkTbFHrmwELJ02111kpbUHLesmteTx49
RUAtavvbLfQ1Pgi5NFD7xwsQflrQQGc9uaHrdO8UIWA4+nuZQ1UqvUO+EaSTfZvX
h2KmgZ3WO9HFVL7trRqF9/KO62ADpB+lG7gLcl0lZyhXRtKu9bxGM+K5U58skfWK
hEvnuPOzJvmijd5kS+XnvuaQWVlcfYyADaP7IbLPZhUC3gtLL+fnmaFCFm0b4Eng
b7QAtKUir8HWOU1hwHkTZXCuXQE41ZL5Ni3A+RpLk34QBJ8xFMQ/s+/fqVvUM9Z5
uOjR3b1v4swmyf6QgU0esXkn0PpPywVFExySk/vJKcV8H5Lh16AQNFRLRZwqXy4b
D5iA9KT7yacJmAW4oSlEchCMS71QgDxbHjOSE5ZMktugvwyuAK9WiNgztCx3Qfqs
Y92nEO7/Bqa5ZyzVZgTyQCehwWWssFVFmlLSFKQOvDkdT5Uhlj+iM+j+iHxSPyJC
A862aTVTPHl+TFkf4mNDNiIQfrM+8xmxZbg2ZWEENs0O2DbeOmCd7CHxs1fKX2CX
`protect END_PROTECTED
