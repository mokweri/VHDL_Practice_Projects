`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hT1NzzRlw6o7SDtiRshd5/FHUqFLeOFXPG3maMDYReaQgCj+v3hIexZMcZCooL7q
V6fJJAAfo1C9OD6MF3B0IE6yZknr0TgN7fJOxRuEZQdrgyN1Y29mVYMHJecw+xUC
FJb/C7w0ALCPOxotj6iDXdKgTdqmAIUWGWrPIMvdclfY47hR9aOniPgUww4CRJ2P
EAhlvjhLAEaGnaWF4MAkLGJI0u0KtvimjBeKNJxe1qMFSCWJ7DgwtN+aRBr8+I8v
IXtlNcZlA83ZdHMz+VrXnLwpzphsRpI1w0caXgRGW2beUEn7M/H72yDuMgkMb8Nt
ruSjJqxctJ2MRlKFCy5lwrxsUcjS7JO7/2tz/zC01YUPNjtoW8Fnf3LxZltcdsCM
dnKJIdoD8BZ8T+WNohkfAWjrS5ek9G2akxTWO3N+hNXdnW2oocvTofE3U3nx8day
8lfAcYiI64WgbhR9l4CtfDnXlPDwpkeLuMfUOLZ/NbhCzNxGEq+/54G3net6YwIf
w5UklmqZwmG3RyAtp/DyfuMhsf6qjwNvJttompw7pxyB0rlpKbJhuJUTwEUn70FV
n1GfHp42aCL3fc22gdFjoi5l1PqwTYUBiYBSXoWoxq7OF8uUGIPqJlDJ5yMvyV42
C+yzgEY76wQZkz4EWGJNFV2WsbmPk2ZmSBDoM7xPEqTmgD4aBUc9txs7k3liNF3F
cyQDFYzvTR0W+EjHW351O5o6jWtpyaNhUSlUwGnmylyAawW7yYNvmdo3MMJAUBl3
zRKUVOLLEQyjlM9N/1q1GrTMW8mnobcu2xYZHBw6GkidIEloWyRMxpSP3NEaiE8Q
vONs8AD06fD1Y906W7Gh5KTU7Lf1qW7dV2IzSMz7DEgTyUzOSQFWo4RMw2H8MEW+
tCx7jE5BTs2KYwBQ4cMu++a7g4sV8fHN/GcU3P/hQ69XF5Ak5M8/2q/tviy7bhd8
a0ktniUm7TYhfwteM/W6guDjEK3ScFIt3Xnm8APhL3xHJ5hfuqWStUFfGbOP0HRV
2tsp/qDSUEtxoW/MwpoTknfClspg6GJZ+YGYDmpe/nw=
`protect END_PROTECTED
