`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GPX0xmpgRnkrPG+l2E+83+uwOGdclTA3qg1VTrGD88fEWSuYayZPgHyEU+3eQyAd
6+65wLvmBhDrUHP6RKSrfsF+hZE7GmZZMEgePqhmU/bHsYyfdy5uXN3gZATcQI/4
Td+LXf6m0gityTbDVi8wdQYv/FdVlmXrq0Rp+j0mcm4hYbleLN8HRc2YbvH2KGOM
rJCktUh9XypbobDIHAqPiNoqLf5u4N1iltKay/muN0EwC3xnBA78PsuvcfQvO4ct
cOWlUWRQptUKGCPljmFggiW68qiFYogb9ZqM/C6zdrS1QyM/2pVkzkd2/YvtG5yO
Pj/+fm1CiEjtx/dUNe2VPNlk7zgLiJ6yz6fItEvcM4+GLD3A654jRFZhrITLg5nj
SVA8o4UHrUYKqW4GJPZixdKgRti6w955n1rl3QwkgUHR1k+3Fj2OpKPLKBr64hMk
nUWkmVbYt8dhlmDIJLCPuHn+V8QCnkbci/JPcqzztocWuJtDfVSVVgMc84fp2m3d
AJfcft8vTa0ABXV6LAOB+8UAsCpynGu13IbcxxG+5aK3p6UADPeqLdIyS0L6Ix58
hdvHNoNdg7nNmhr2rAsQ34iL1TWGhk1c6eUTwfDeq0K2w+Yg5YOtb6rayXBQBBiI
hu6f9J/1lV3FNMrqPl9hZnlVr6ZsNJgvWp4TH7THchEOtsmD0MBWwr4wRdjUWByO
bwUbMcj70Y6M6OJ6rgbrSRe8mfaJDz6sb+f3SL1Ms6+mPLF5ZJeJB0FHLMjWQOWQ
ev+aIk09ZNOHt5200jQeD6KxyZ4q4q9aZXZrOppfQ9GBz0anyJt2YD0BTD7+yLZJ
`protect END_PROTECTED
