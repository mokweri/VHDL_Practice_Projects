`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KJC+P8LkRDNxuiJ8u9sLLNjQVwlvg36z//6HDzXIfAwAD6YRNVdKXeMgPC99Net
92cpnVusYEHvwTgTiJsGNJ3G83rYb2UdiW0PvIYVd+OX0RaYpBM0Y5hhI+lPIJvM
GVx9AgY2wYwkqa878KWnf24BrAFhKwGuesi8Zz3nDcukwkOL1H+ghnqO03fSoLnB
LJ+9RzffaT8OKYi5Q3H4IJXrlimQL/pHgXnftv9ILw/cVodgFxbJFSL0gdImRby1
GaYoJGZ+z/HJAKJw7vpwNq5qOcufaqwXG6fkoSbV3IK8mGjUf/Dy8hZdhvD7wvfI
eJ1ThGOVL+G5AhxCboK66C9NaJ5qomI3uFD9Cwkx+Vu8kvHli1LRNT6/N6xeoBtj
36Jw9HDu97SSJaPfXBVYCkUI/lKU7o0MJ2D2KVICkDyb5/R3DNKWW35P/hQzG6ql
mlmfMxjHdQV6lpRMWVswkwzqRnnFfJsvp16qV7HXQwMEsPGa6JwIhlwVLJmQuVMU
2qw/wsehoepIZWjBiQ+webgVmFgtJ4MwLhWCO6A6d5fCR/qdFc8QsX9XYeNeWN/b
UR1uVHnMXmw5Q584Pe2H3ZxsQcVS3Ufc31qrPNbOBj2zQP3zvA0zTCYwBE4ROJb9
vc5wEWy9cXs6e2Llo4IP1faVjT5Q426u8E7nasWLd3qx/A+sExhmhW3kVll8lQQN
PV5OszNGgAAgxkUR82pBl1sStADRtBbbzUQwjSPjTmkBKPiSQSlsAppEQcSdLvQJ
KeLnL1EA6QtIxU/uTZBh3w==
`protect END_PROTECTED
