`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrCCsBHj7eGQZRxOzw4ySBbQYgYI/QxMg2g7CIvMLb4YfNyujIFdVo/5PtAjjUtQ
HS4p2EZak3ldT24vaNO2Br2hR/iOR4x8l8AHVMEpZNtpajFjHJUHJKbFP1oxl7zV
/qR85PirocJ3haWLG+gSW/yioDfzgWyZcvAkWafqkdY2a8hf86mI1WvcPCWxeGDa
5DCLTBUMkgVQqPnX5sE53KwCqkI/QR1DRIUtTh8vtcjKG181njbzkPtOeKe8ZuIj
eeZxETYfQLugB8XBeNSUmwJBnvh8Ctf+TYQj7uk71SJze3cJXcrJNtNX4GtUtsxx
tXiN8BPdg56PL3038Laq+yZoej8wHKvOXrzQ0gKEYXCjiCKyrODblB3Ny7NHNQXL
yo0l/VDK/ofnsSrRHBc1feHJbZlrJMqgcIl+dN+J04XMlvsSSWCVn2f8WMisE0qZ
6b9qFrCVbyxmKltnlEUbqU9ygpXlx5DWJ6YyM59sZuyZYGzNnVmCrtiBDWW3RMS3
5QQe0MFQXeJ8L+n+1xfm/rWNEBJKSBsppKkv5xG1tE8Fca0Udokkm2WJpMvLyWXh
mOk63poZFmxgxu47Qo7SfCw+zMqLlJMFzxeQc+s7bEBoQIaaWQgpeN6hoa0Qk9u/
VvIuU4q7kiY1C0Hr25CUjySXeZXq66LTkFybo9YcWcU4cuiYN+lOwsJrGL4/pVZy
CwffrL3fbcNLzVsCVkwZfksP56tf3+H1xKc4ZP7Oy+RnvaQbML1Fo0gQ8gqbfQAn
6xQIpy52brXoxZpOqygZNWeKy+nrWbAhXPQEfAhyxWdhmFKNYavkvvxxFoxpbrVP
kGUoV/9akbkQAxxQ/9uh+GV57N+TnBHnzRyx2arba97il4idb2jjz9/m+oquOnHJ
02Dm4+nuRKufpzZdDSQkQOzuQwxzIf3Bn0frKPS0nM5tjZMSf+mtBooOO7/Y/s3B
7booui/6Q2+6eg15kek/ZO1xK/QYfmLidWgVYxJ3t1XYeDDst+mezlR7Zj5qB5GX
mkFviTuIIlEQoGCubwiVWjgpmRXl4GDUKoQQEr/oYr+uzTivxB0Y4dqp4b45U4IP
XcI6HKHm+xviIrSb+vdf475Vj0oxReJ1wkWq2Zb734CIjG1M40DkYZjjzk+kkwvs
uqHZC+fT1YViD5jmGSwarSFhVb6dak1X6S3X0Y/4tkO3AsrdVTc5yui2Uii/7PCS
xoYX8Rv34tbRHxIwI+75YRtDWtN7uC+br3TeyHZCYg4xHE4KtKBL9/aYSga2XboT
n4BDS/akq/HFEy21ndqJd/6rBaNo7KItDs3SgBqoPBlOKj7oGYTx+bsGUVBPCLQC
l+xgmxqDp06bMDd/jjcQFOTtIMb4Oc57YvG2r6xsd9F5FVdx9PhBj/fvY8H/+C2a
w0E+xnuW0eYGACc8MnVzkOPdOj5K77RWO5xwfNg9k21S+KJ367H1KdybK69mLOoZ
zopOrPwqdKEQug+U0m48hL7ZwQT7NbjyN0+P2giuOT9DAMdRjdjVKdlqARg12OFa
K+T6mZ95o9x5LYK5r+EPD+4Ft4MxJDp1CY2v1sRhJI0iZaF1/CLFfjdH2Mtii/ov
8F4qsuIKqWD8PH/vC+CNlXvWpw0H7uk1gVdRzc6fPz1PWcnpMhMNneqrbQQqPmMA
LjXgCbL7RpWeBX5Sv6T1fMl/cYsouYB8fyZdyBlRKU2oh4FSCIJZWY1BAxXmUnpT
xNJiAzsdIIInpvsX9ELvMxcy/gonDQhYm0JfID+3IxogK59aL6XP/2iITvmGSvLR
aJx0tm7ElousRj97f/Cej3nRHvKoiBNiJa1tV2mCmuAL4yyy1DggojSU2i54lD8r
RISIwp8XIwI/N4mlf5ESQRKT/Y0LBpIK5k91nVFPHN+llYtSaUiuS9/HEdK9AD/1
wPB0xsCRpMseJ9CjHsq8WUAtv45EMM3Uo5KJlVasxpng7UZ6/T/z4MdBN3Cu/v8u
DGBlFdLMT3XH66r/ANkQo32NScrn+33nOKaW75zA+HWnJEjsF1I+IXNvV2V47/Ji
e4FAle7u6OZkS09bR76wHVgnGTPa4TkKbFBc639ao2rUoZnjhvCZrio2vYZefaUo
HJv4yAhaId3ZagH/YddeytS7G7fvW30fJ+9ODqtjnQ9DRzlfjFsUkOkus5ZkhDb+
AzauRjtwzb2cxdE+b1tFT6wv5ag2XRRiIX2NvdV97sALkNME78YFJKW+z+2wf06+
h0ENWbjlQ/5PmqQ7fIZDuNAxtNaCXyo71iYpzpKy1eSTgo5VDPJzJc+fJlawhEs7
eXyBPCzj5IZMS3/TuvNFId4z/NGHt6155MBqsiUhrhp2EU4Qx5HnVK2ve5mNdcWU
91ue5nhBJY/1EC/kExCALQ==
`protect END_PROTECTED
