`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0GWzdoLg9HbBLiG2eIDkKDEYhCaFIQI0cUtN6eSzotGfEHHIwDAgl/PEpTotKb6
IW28BaDJ87kD4mpkXlRKjeLPb+aTjNC23texeDHMt+slFOnoyvXBZ13hCEVr2uo7
S/uxAC45ZUhwOZ5zTTynEhJzxf1b23yLYClKYAsPIw7W8QByXVDE2+5yB0lV+9Q/
KKhjEaBrCgfTORG41UIwgmv+h7GATqUEUFAsEt81ba68arI0+1N7pWwMpFbWfJcz
bFDauoQ2hJj8Vdx6R1td0cUXGEwwUSV9+3q94FeIVi4rLASFyxydFMHmi3oi4hF9
ZFthbuhEmJZls9UtCsCGhQzieUmG8y+hQwjbcsseNi4FCPScIMmxJEVAdagmQCFw
ymc1X2lQKJsw4ySSvptvCsgelP1JchhsVcYTOAas8lmgQc15/tN79HPT6LK2TLr6
plmyeHH3iY2peOBSk8H+jVzpKUyIDPfCiLuq3HNDERW6Tav7xb1a8mor3+cGzTFS
myRw93edF3gy3867JP1p3U6/nXIFgoKpmk6bPBvRLip2iehkaBq3WtBY9sNxS2gs
bLAsSiNpSGLPBzNnLS+nTJOvhK1XHHrBaZvhzrjm6LzD2UPHaqpjrS33aFlpVpsX
X4ZgyyXZG1FqOaAefkQPwP5qiyUue7eJu23627AaLOo3ooORA6dplz0rpOqpRFbJ
9MJ23ilF69NjKtuj0HAZSOacF8mIIFZ7EfNj36cIliTQPQ7U0OICVnyaunjoqOCu
4NQYrGns0qF1buXxWz+YZYjZwbkf5Y4C2Un5PMGTKR/82NvpQv7eDczEzWydYjan
lJ//L6tDEFCeAHvvVQoeLXTO1Aw5hPebBvK2GDybC/yeDDSu6BVBRVRPuC/vehWa
+Xpi/nXn6yHvkDwafOF7BT8TEGjGzKvqOhDC758lxDMovDSkAt0QEQt2wud6kWJ1
svVDdkUbuYE5gyeBvc1G9I002HdnNXjch8BiUgSOJrWdSxWxSo0Ko0ktGYwaDlUd
wxfLzKY6PIdA5BaVWY//nta0Ej0OaG/IT4EjWZlitnFJeitdbefEtGm47Vy8q+li
EIHRrRFgbb8/yxkqdCl/lDePkKNnq0x+tc7YKBHgweQ=
`protect END_PROTECTED
