`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+rHDtSzCor5GwainaYwUhAZz53QYtipoJkwnJrd+z7V4HSIhd5cu5LEuKh6CHZv
UO37RvD2YmH0sH/4917iyqEanfWCEZZtalx4RfIaSj4cg8Kqa5OIA5qSngeYEXAw
+So9XyoTRTNNvkGu9lpyDgGw09LQHlo7TA1035UdsS4E4CG19B1JoNiUBmULC4yn
3uN1Yj/cZd3ccylSe0nhmhJUX7AD/+CozxQi4c7OfsXdH6zzF37bEFuyQt2kF9zh
7iimoqAweu0pKNIzINikyi9I6OY1fWbwKQo6jXzXCAa+nD+rIE+FhW6bwBZd/8sB
/ofoRAWENhcYWjPokEl0C6Mm2cnPKUYgWgdVwZYuH3jq16hFPFMaT2UtfUcHqk5J
nIjzyd9L9omAg8PEAr3I3n2rqGMYkvDrP05BmY3FZtj8Kysz8yqa7/cKWu1KEw10
dnfeGY1+LLy3ZW1RFDEZSJAqep3tK0K54WSclILy8FoX5fXR9guk4P/mf7lH1iUW
nsRYiIyDBBWSoil93HkSDGOZgMBrg3oXlLql3gScR/Hp+/NcBtdrf+ZMawlluzzP
gkFjMmvYJCIdrCeO6RvSBySByAG9tVGTnW55QrG5XgKZlP0qBK5EMx3hnaFnml6z
rEmFeRqjaZahnWAhJxKEtmSQwiiUGSMDXDm/nOo7GTlf13XPZHqmhqtKds0nPwow
3TdoNDMzdpE6wMjGqAbnk+XCDh0jr7DMspd5BeqxCNKLyD/FPXDe2NeqmcKc02N1
Pnxxi4azTrjqw/Wq607XoevTTqyKSCs9HMGe298BIYHS1eOd4HylXB8P6aNBByUn
fVq6w4atjuR75NsA4eTfS5a3nK9YoIHspQP/dTRHAXKocHnl0bpJb+bEcDxBFdIZ
DQ4mckIHBV9pF95vUhmt4qB84bVGvQ+dpIbn0d1E6RzCqQjpX4YWj3H0TRWVCLeG
8QbkcLc/f88GAQozYWaDCvMOwijWFhq10EWxkrr6YGj2cc1EAfvUJ53/lFeqemjm
2HgcsrV9sGK2KnGTa5FxmlgirBIzDz4vE38mB1PqwlC+j8OCAtLitjKRUuUiwoXx
38mI9zpFnAQjLdOOOxZ+wutk0gFogFtP1MV26XYVcwQV5e91LA6iGFPVJ1iZa99F
hC4eeRaKDY1KNpSpzyRtktnUf8wGXsCi7PiL1UtG95oVlVCtN5XGqqYL9aATn80m
L1baTTecD0HxCQmv+tW2Z4IzZn8FsI/1hBCG8Gl5l35fPaV3PSjHPIzbvGTPdXYH
xvlh1OduMpqKmK7xtpO7a1zEAxeD+85lH/Gfa7GEkILSzAamjMyBy2GxhZitowpj
qAxiQSJhuzLSnSdjcda44qKhIHofCNDkMQzNaCdgXUI=
`protect END_PROTECTED
