`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLCP+wiW8jrY0AnwNfH1rdOnQYkeq3XY6+ldFw6rnGlH4hoTzQmFQoHxIkMbATNy
/KUvaImRhw1yQzir8wcMMmVFLamc5W5QCpEXrCzSHv+Q1OHpwrCCG5ZgpD/I7DlK
icvZl3c742o7xzR4Dpwa2IlbqLx34e74GYYdLkQMaPwMJBPQTcvxam/uNUR5l5D9
UZNh3j09qJNjGl1xBT3UDwRRTJHhfV3DWWhL+rxTR5FccPbyahJO4MtxT7dZBuGI
KtvoKNbvpIZxjy4cAt+ox+obFzydDuovED4uV6YtOUpS4Zwo9rTU9rIkOgJKI8fG
8UXSrVeidD/HPkwAcw0KrpzjX2cK8/vJMOfAlOzWgffpOLIh211opjleZu1X3tAQ
5vSFLuE+E+cIw+5VN1pX7WJCDAorJIM6O6qKEm09hGAWpBR1kttYx8Aq332tG7te
HYwqEO3tywue9/EI17OQvz+MA3kuvMHeJ4fmbNcqSkSBh/sIg5K7WPnP11tWMk0b
y/+HgtlNGyby6mS/5NEXDtFO+0V5m7n7I42yrS+tuU1gQMK7JlkDvHa7bnzX5pQj
IY3ZmiD2RGK0J/w+CRvSIWjVihUvfeh3KhZOVZIgbDKeAILGYOK8GQOYOaz+T+HM
WeCTbEe944ki+3pJx0fwO5ize9iJaQh3OrlMcu/8Vi/c9Jl3qpSzSfVKVR6E7XF5
CwC6BkCINDEsTLCVhvstFuKzpH0VcXUferPU9Py8F+M=
`protect END_PROTECTED
