`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aikv7UULiLgQL/pa5c00Fn1d8DhqPrOSARa6Gpkc944Ll7gKWbcTwbVNXB0vHXlR
dzI2x4GvXvVPDxjIfBqeryrEcVnm2Ph4oiYKYsiv12IFUrq0tVJZRY9q/if+8ip3
A5OCOnT6rZHqnIB2nrS3lLpzP5dbBA5Kfh2YKUpvODm1pgvsvB5J+XhD03f2txt8
6b/8r+u7k9GQuCXpaq8N4HLn+L5k+FKhdQK83FmC9+WBm1DRPdLlmRjrWB4qiOle
A8k8KItas83vokRNskW2XguhC/gLFc8mKBi/nb6PxQXEFOHispEE4Srva8P2uIfx
FCcktGVtw+kywR1afRQoFys7II8d9gculYYwSHLdV5L+pNIhXwJatp9ngkCIGPpA
nxrLWAmpB7pJSmjtVfavebrDXea1ky2+C7oynafOxVNC3e75ZRyBDZAzemKB6hd8
vfIZPDgm8dKHzy/FLNhpb87jY0ycJPGb8L5KlAZ7d4g=
`protect END_PROTECTED
