`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zrNMJljjwKj6K1/YSq3QfCL0wQtbAHpX+eB+njXfTp5IOEfPxbXNcXnN6+/dWuFz
NC/uL4n/IUjIJGwtvqktAbDsqL6hc/rtrelUgj67AKUO9SeXqxHrkfJZtV9OyxU8
9N5u4x0GyYRUkHtOaCGQpmfDDxw81TAQJImhAUNXXyABphkOnoe68gs5WuL8zlg5
GpruaMn+MvK2yRSMhcJck3u0eh6IWPPnLsf2/Db4Sbz/UyX41YkM6V4femFDNv5F
mlJ1K97WDMYMUPWI4owS6Z7kMGhnjWlQe7U4jOQk/HTVqjU+v4dyzpL4iUkxBZ85
AKS4yIwwtr+Vgv4XgojQ9MjAv1hK8zxqd3BYJc2PzQGtGwyST7raH6iIzEppnjt7
Wn1TD1hx6ekHS0PuHb617ELpb69XQwS8eNbox/cucBkC55tTFBgdexqUFUO4avcV
a4p4xxSloQv1ejh40wK0bYiOVOXEUScn6WtUNhPy1TV3RxP3PzAHNquJ2XPpCfuw
ohXJaPzccw+4RloRO7bM4eEu3w79hYry2lGlxGBOckl7n9v6ADSb2nUKqbGJ1+Dr
dCPgiYgQeFAIcxxymcVXzCjYiJZXlbozBr2AYPoyKC3tDWfF8kArRIx+8OXbdZXM
4u6o2Q6ZyMfwuGGHdcJm57EX4RWpOfVPmMlVCwzwZZzYEcEhh03PyaSJ965GDL7+
uHi3UbHHHDVSS9r909i2VOkC4apwU+/Ws6MTZqXdnUSYQ21B7p880z2UlCJGXAbh
zU8tOQvMQQMULS3C7FwAj2+vMfteJRDNUdqOhhp4wvY=
`protect END_PROTECTED
