`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QKyFCML86mpfehDi7M/Yh7T6tseXoBPtDU+4K2mCwiSfQK8zAhrl0g9GnTcAz8D5
VU1KVdnpfBkJTvj+XTNI71EGT+Nf8s93y+h8xJuIfDJpEfN3RHQn3ieWwhV66Vlk
ycvFuKAUri+DgfzhgxmnJOAqMFBqepFAnQZ8u+cJcKsdzjEFrz/UYc9duye9nvcZ
egOkQR7lNSyck29cCONLJlvRMKjlZQV0LzE+5/yKu+bJWqkW4elghEzjNgzBqUnb
umRGkd21Prtbf7Ut9AhUqOOA88jHGcyc8Vk5nINiFHI803/JSz1/qGNXhMsNflxb
oNEDCpTWissN4hDYk4rtwxoimvJWsMC6eXlIxNdUpgETfII0S8HWIX2P6L0jCSqa
d0vlDT/GxgSk64Cb9vTq3tVRVQF+Cabff6fIbcnRJqacXS4DNXeXh4EiN8wb+Xl9
s+nXD5c46CinepXRqPHdRFy/F09ktruz8xQwg6hGehFyHIwo5iljWAxoFtGHGVTU
NBY0qH7WJXdDNBIllSG0uFrP1QvpcK/wZXSmx4nGncrOYDgoWLsEALTE//+SyQwk
sh32zmO9DJh7zNfPYuqMpxJJj6XN6fijjnLiUakWcWc8aFrD6lKZAolZZttJh0qQ
kZlkipJSZy4ImZ98ShBABFMCwR79W8AQFzTkKqlI+NTCsr5oWMqmOFJdqIUmFfWQ
`protect END_PROTECTED
