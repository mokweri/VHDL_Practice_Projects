`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tdQdpPkMAoiQKi+5iaTkS7P8rKgzgJtOfokyzhVJDW2MS5sBN/Uo0ZmTaUvIkc3
CjWfivm3yN+TkGGznbH3jIRak3vrJV9BmcX90WmuPv9C2Ljcuq+3ITEYtjLGo73r
fFRZxoqP3w+oLCv+Nil8AC1drr0W1EFRNRCffr2cdBTJ/I8m8QAuzvzkFGas/1qQ
e8VR4gpkPsRhg9FkTmM0iHJ8XpXQrqJrQ/OF9G/zaqMuLhUwqD3Zsp177bVzk60j
Oxcs1g+7exwSuWeTmtblPyoOEKTDvdpz+WBdt2VmXOEnU5FrDmReZYKSo5Y/8yas
uIk4CMnk033aCqtO2nsjxLQlcMKqDvmNbwKqpQjMAq3Vh9z8iB2DJIVPbOYVZPxx
QcllDXjuPo+nZkZE0ZBnIcdSwx9r2Ot2dQddCAYTfKc=
`protect END_PROTECTED
