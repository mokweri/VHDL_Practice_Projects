`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOZMmpNNrtkMXEM360JIWNEojbl8fx6A658F2WtTCH6xI2999vu59nzD44+f6lBi
jQSoo+ayOK9xSMA1+KWiV+PfiLaLz61G4U8c7vhIbL23HtMvV9gkllLzHGZAkRFA
W4xPhl5HAlPHkdWy2ZfYAWX0h7VLhlTONot1Ha7f4+vXOePC7gKhaAS5MX5AiXrG
UqHRhgoc7aap5+FUCPJ9yPYMx+BgoDhzdjV6pXYun9X4z0H+dezRPOSGJy7oj+6B
1OpyDepTWAz/ASqrx5aaaOnYgv3BT1gVDQvcZeTNfyT3N/8AhcYXFCScSJYvwd89
+6lCzVT4UWUfsMxjtz2SBksz95fab27OKG/BFHKaYhVNBVWwEUUo1WxSTeCtlusM
Z1ayyRhPOIPxMEcCSRFLZV17VeUK73dNtBPlg9niL7CLY0JrAYpj1U8DigA4+6Fd
uFPK4hZOaGmJDxyHA3xuOxBU1y6fpw4N88NiZ5Gtt9EL0veGN3FA7Dyf7A3G1SRw
`protect END_PROTECTED
