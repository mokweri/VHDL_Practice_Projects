`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPeKVVJNLX+FoGP0aUKMQksKhRZ/PQBLlVtU0EyiXh7Qpok2pMbC6BJOGbkvVQ/p
b1nKp3RlEgFBW3xtKlUrX252dQYMp3ncLB79vdpeBAEaUUGlV2yBMariSAZkTjFI
pc0AWr9jygCwlqJt8rFprhRaV/AW6/TMpXkTn1F74m7gFp2w8NsviXH2XRwaoDNx
PiR/ZvYKXo2EzjQ1KgXhngNhsZAJOLu4yL2S2/QdxdaijGCwvH/aW6WU+M4EjfdL
3x34lt6HSa9mc/bTi/X3tQodxcKi41Hged3V2Jt6rrTATIgmUKdR1xjLmOMXL+Rb
4SwrYXknPdwKe2cu/p9Tr0oFkxZQmID2Dbt3L/RNmAYl9ulmvb9d5pIzxtzBixBM
w2KGaS7HJDk2sN89hP0d3Pwk7F1FFFwWs3eqck0J7M5dTANVbM5JWhdn/2hwJ0Ce
Rpbjv7pqGtamnXPxdVhrTzdELhMVpHN4IpIaJGSm9WZ2xeJ5ba2SL4XVEpIUPngf
4Vs6uBfRzpjzxo1Ae8xWVZI6dSLuYN4ssSzf7J2HeDv1oY4LwXENyeFpHPnmOt0/
VpVyZkD9/5ndo8AzH7IOD22caD8/Jxc09pmOEo/2XUl3Vs+FWfB/DaguqwCCy9JE
n+vPfoXnuySNN7xGsxGabGlhKWg2ix8oa3S0VHCMJvF3CdT3E1jhLmMQ7AxCbrXh
QK/Gl1B7jcSw8BYHKkTVgFxOVwIIWbeAe3NEIfRbNd5wPgN+JpDrtRFO1vVQnRel
c7INCO7E0iNSeS3ThEZhly4qZrJyRB1Qk8zSkIEaOxWU0cxyhpLx2hpoiq24uaW8
HLMmfPaOqNRuK86fr6t0pZ73ejf3KpLTQW3Bp44Sh9d6/Mt/HQjyqVKECoa1e5xM
8+w0ONAmtO+HwDJBryoQ1VCSmQAioLjTtPDjqaDs/ScyaWHL1vDkVMVgeOPiX53y
AodfoiwEpb1JW8uKTq4YHmgFnsXSuR8WWlCdHDzLSdPHOD40CgehfHraJ8ASjR0W
8MrxRfKING13DS4sZTYnJDVtJgDaLg0tcSctYCNQ86KcvNChU80zv62VyQ1ApcKa
7AaFdXNTJ3jc0KGORZU/nvO/vUKiqZHui99K+vmCGyXPYMlKhtwreg8Fa49y5TNp
dyB0Fjdseca+3V3KTxjyrhFETGN3V19Mr/ZbmOVzo1AXqwwsFSZbYhnKiVuNYyVK
XZzNEMAcujFtIjM3CZyGZYYR9c0NWbrJU3vt7urt0pxhJFEsscwSEczSKEiZ7m1D
XPCLpyFdY17CuLRc1ILUW1OfCmVy/gbwoLL0wU10lXeKyItiMA1HWe04RNx4tXRg
GsenEdKkZB4v59wbpNWNgS1/0v+CSdykbKDvNPVmSHDt7iAky9n4VmCeCTPwoNW8
P5DQ7r6q20GSiysczMl6Gd/ktD2QOUyVAabYRAL7fW514t1Nw+hoHdzrPdnyOPtM
Ym01wbvwetez5FMXr28YPecaa5KpkfM7LdB/BtL4TL+m2/xBhHnOaYxg+JFDEinS
FpmepuHxS1VYpBAjbQmtD0/HAxC9Y7XRoXUQQc4TRIzS+df7+P81rHFNKHWB2nKl
f+t1ss64haXW+d3m89gUKRwAHDxqg4pbaUuYgw30SWSJXvLFFFKb8rf4u4EpSsLB
Kdyt/c9isldmoWzOBjeryNTEmkSixe9R+q3aNeRqbICo8VylluFQk+/lJqxqsUo1
1VWQposqj4uWJwrMvGwLrFVWU63yCYQprqI6S+L8LHFH3fnrvSb70St2+pNd/uNO
xz825b5z8oM0e/zDzL+Eclmk5l634kGZqbRqy9UPpQBkjj5vZ4KaaoKtYfeRF6P7
j96VfFzFzD+se+OGFMdTdwsfP40o8IMwF/Tqjy2f+/B1kxnIE33B5FaMdF0SXy2E
F1YqdwbvzG75DSAaTy9DCmd83kPx/An8qPukwDmgEmBchsDE1Q/vigzN+zsoa9l8
5HBuMft9oLTjJSJwPgA8bFQbbS0Bo+4rNsHUGfVEyLAurYc3hSt3raEWRPyus+EO
ybLtUot0e9nCVVAp1If8aYkHuVB63gvRx7Bq/JLDmkDNFhu5IvMugGif82coET6l
/d3T4sYNYTQoVfqZcDlcaR4dT0y8tmZ76Lt2yyfehSvgpbYrCHjl1kIFod+qc44V
6nMObntlcJOzFI3OLBGNzD7xlanCWrR3QMfI58i8Ly61QN7lI5NshRhAu80K91y3
gaDH+iWFzKw+zpX43oDd3YwFGdVBtRs3CmvkyZl3jCqXDQ6uFu9Rypk5DY+lzADS
0RGkYQVf2mPVa+2+KtFxHAOs4z4JcQhGIW4oQj+fSIg1JoaJTxmx9/CRMagSE1Cw
p++g8nVic/xAATwORqqeu+MOjHJNZO1gh57EyUHibELG8SccG8BthsjdVsc9+fGg
ScbpfBxm9rzt/Aim+Fl69g1Pv/uNemFUtS4V8MS0dResryFa9IDQ0t3VrcEycR85
UfimitbbsDcyREvuAn6MiIX6mvSDbp9I2o57EN8+1KCU+6Yl3qMrMI5Uyj8i4ov5
UwMGS1ARKLcyacs9C58DVWlIV0HWUleP7QxhJUG+CAEB+R1SnovJmXDycUuIlDU6
741o6DkadxFFb/5k6VYRapDGldbxD2pcP/E9JhUraIPfM0rMlFT+m2wLsGx6oxfi
HrpnD9bgaIebvc7NRZgrNKJodw1JPpVHRi7NlN8LMhXmbh12gsGabXFi2gqYFls9
aqSSpPPAvk9GIRB0H5TXAk06/UDJro9uczsWF09ZHw9x3/6gHSVns6/MpAdIFtMn
oK6Qeo85laCK26CnN3rnMVeP1KRYActydZ94Uk8WbrXyLE1wxeVJlVfj29kA2fK+
qoGFtiORH8BGLOu/0B5ypWSm4XgwOFHqbPk8Riy6Hmc8YZhEkW2DRXkbF+Nv8Bw7
foUO+FH6U36jFPKQzZ5LnFkAELmAqBv65EhNWtVme+jH4BidD53MFhTOBhk1/Db4
Nx2A2EjY0n0bbXie0Naj9nqSd2wA6MvVYqI93/75FzHsKsaPO40Umf2yHq8fgRYy
oYrtopWMsWQNPVpAqAOJo2fdHikovkF2NvVdtPew34CaC2AmcmCWoCV72SDveVGc
1O8XGnEhnkPDph+8EwQtCtG5o8GEF9tPOKx1tUWQkJGbQA5ktBnDDadVutfqBkMR
fXd/qMXUgb8tMJ4C5VpMfgleJhs2100tsfU0twDtlkEiHEpI4t64sNpwgcMr9S/Y
hamhR4VGopuGGNU1D9m7grg9EJqQ0D1Y+MD6b8k78E8vUUs3IiQN98t01+FoZedU
hN5E4nmC67DhTVG+UYlMECkkdVFm51IZh8TP31lfsgj272jgf1oB8iPYv64XfTpw
vGDwAZ4u9OCo9Vh7GeI4ZSYtAcSzdUBz28Q//EaJGQBMtc0B6L8+dfIy4pPPZD4a
IOCk8pVMwGmsX8DgO5EERlk4yJJ7KkY47qRPIhUoHwF891JId8Kjf0OV/Y+ldPoZ
Cm86a4nICpHyyGF1yCV9k1LPd59GG6O9qyLk7n3lJQvoc2A/XBCma6IpUtdPiBuK
PiNXpu6E4N5s/a/HohD7+qNN5T7tyXyMt4M7kuqSbB4BZqCAc8vO5EwsQvTZOBn+
7cJICYjz3vOUo1SXTjKaKfFonIs7ci/s8evHKUeBrdgqn9XVA2cJL8v2KPqsMVv/
lKPA6bkfNo4xtFqPuGS39Wjpq5Q39P5IJtDKgNpJWJEIknQqXFmUcu/+ihyb4D8l
Gy8K7EJSks6/+bwSP+IZUjRPyqdWq8Tg9WC3um4zlBH+cE06QEgTDvxIxu5RUrV7
oVRiLrUuUUDrcS7+vQrfT0qMw+rFwV/nnJhbo0j8M0BuKaWedR5gu/yCLZpGe8cb
rHO1P6H1BlK0wAyP9X0Ps43arb0yPfbu6Ph4nn2FEx9QVVhrJw+5CX9MHBbRo22s
sAyQ64G7QIcgtDkuskINypx7E4G+gDIeZ8B3+GSrquvaJIqbsDumhP0K/zV4EIxY
uP4OYqRDNsC8g7wI6PiY59ZUH2lSh3lprDz3B3YbYB8dr1if+SkEbo+dO1WKQp0W
6nIRiaGI6wpk5guqNZOe+8AJdOApd7FxpW+yU+Do+KqzLKQGsSrbX54p55kTmTm5
MqOkWO77myx0/0QCXayn4rrspXDlyA+HHoBzGc4XWE6yUcNNyCqc0CQ1uxhmb4iH
8Shmv5eIzUNNrwAjfJ4R3sCRLeDXRGQuZVtCZ7rEHkxemMRqSdhDoRibRrxUs+Qa
NUHWBXZPueRtIrZJOYZnlTkDaHMTwrl9kpip0CQC9kkpCU6Gmyq5LaxCuHa7WYo3
/IZeIOKF6ArnQVF11tCKFdGdVAJvmZfd3Bv5P1w+uSletqHVcBlTCdXitrqhXIEe
VrheUX5onkLq+EBb96oa2yulq6dCgWMEFoOwO5kqcNwCzUm9Wpapek0Y6/cu9Ivu
pdSQFkhFA+Vgjf7043ZIaXShppS2hqgSe28PFCaCPFm7Vr8/6axvxUHz/K0VP+q3
vq8JhqGdQRBfIiBAhQ2oVFadOhaquQkVP5Oh+g8t04cWIdj3oC6b9iJPWvMcYvsW
gFj/8Ij/rpC867uCdi6NFnGfhAbIcszmDUFokaYVO5/FrR0Mxsq+8cNnnGlNPrHc
REeBuWQdw6B23iit49JA/PKzZT/56rzYSRn35LwkQH2KM3zb02nW9STXXoU9BU1n
FMy0aeVbs9WE/s+QTcLT9VjGaDkziHuZwD3Do+EUmQphs4aa1klOWRVTEzCUSAdW
OJ1dGCACykuUgZM24bzI0ZtEitxs8qeGGQ2PaNXy6ITHpkXS5GAFKNJuuV20bm1F
+xEVs3qSaKvo0l7sDnsjQjWdkhdgJ6tbxwnKA8ycdFIIoF3sLyKRZNwn/Cc6elwE
1vuHwY0AXOF9DAfpwMKR7ARzaOP1kVmQp9vSB+YYdfKUT8PHxEiNFZj8p3mHyj8L
ddPJ6lKVYAn3+aknPGXLOshWuOgd4wFSYupKZezFsHpi4JuTUp+QbDvW9yjXLtqD
EXyl9DdDjNxeYhZaFQTjbeqdm93JwbfiKaoTS6JLBIuvOAQ2dariqXfZP/yNk8xh
ktpb/YXmw3qN9FHysl0DjaKsgc46IgG2hF23uHN3kdKdLX5b+2A60wLHrsj0Xrau
yyL7PzHY8f+Y9SOcSK3dsL1GEFPF7ELzC3UQd1y14YroibWl8goUvyjjHsMR4kMf
WwfxthDZ3fOYfNaHvXIhVmDjoG9IfCtHWmJc3cujddRgfXlP0nFZ9jgrP+LC2VD4
Ok+Nggx53EK/gck/G1WdshHU//P1+ja18QvBsJGs/CrAeGa/KWwOph/z/SEo9cpn
XsHcVpD78iQw+g5vcP4Ov3F0BDswibtpfkHyBV1ymebILibfOb+oCgNLzociKuzO
Fs8u0NvSEAr+NMmakE8a/rjZxHK25qMkIvjGoWWczLiqe1oy1aYlAbsmMezh5k3c
U17n3Mp/o7AitC7jB6RZM84ndAjpRUnVe2zHsXjuRtgHXlWiFO1a6H/n3xwKbUFx
mYseAtU39dcP3ByNB83WlHhl8wLFjJvmpzkbZwB+6nvi55Mk/GHCtVq/PqwNhFHt
Wg8Jc7663JtlL0foxUJembAiuWqwkBLFA9WRXGA5r9ySIa4LnLFSlaY2fafoAGXM
pQybitZ+rGT8NXTapLp5zgvdSL/DTvz9A6oV65UHNZk9P/WN6VBzoSOPHEhG1DX4
tTB99Xou1T+60vU1o2etUvnUz8YdkeSSNjv5K21w5svpKhzp5+PqG/JmKbDE9PaU
DKguntdihqQZddXfjiDG6/EVSEMkcuwobKl+riTJ4ZQJFWIh7PkRXCArMwmOPFQi
7vH5OtzeoMyrl2LtDm1VaZGtlCNI1bOfYqphACgcKx4Apd4saBVEjnazjgMJf8Pf
o+MzKyo45dvA0fax49FLEbT6HUIAG2HknNZnGCLekOFi21VVAbiBq30BvOZ7B+vu
FdA2lnUd8szJHb6zZo20t9peACUobibJqKENmucAsgvLA8b9nr7yF3E9rZyd04Ng
kK8tvsx0IptjZPS/hEfsObLaRTtVjqFlDV+C/8jfFcL1uvhYOB3b+k8NyOFgsWyt
IM5N+jj1ARNN9tbSJ16q5WSuQylKD4kVwOWNtZTK2R3Rba9i2TWNHt9tIudFqyT3
8pwiJDnNHuMMGPi+wePN8M3t87ZSJHIhQUpZFh0pbeKeGkIsN8tnuiL7BC9akZTr
K2qY/co+uqhacQ+uu42O/iWecf738Kx0TpGxwPE57ty3wGfH4YKNIsfz7PRzR+SL
mZrRVk5z41KfRwciBYbwGlPhBtriZfL99/pVVmZzmQObRhVhrUpPAP4L+DrnaSVq
QExvDfZKRI4nRAn2xikLzvoWCL7eSga3d41+25NSzvlkB0g0ZxTzPD9vrdIYVXdK
K/wziKu3jx6D6TDCYWFBru+IJXMoB5KkeedCRYAh/rYHpjtJ4UEuNzjs4wgBq8nN
fJmMVDNJdeeTzCjPGH/SQNgOKy+OLmSw38rniOSj7dCVfWz81baPR9soDUBJm4JI
Vb3i2SPkw9mgiaiMLIf3oPMi5uvKa1qUb9r4+/0xbNdNpV4CFg0XTf5cyg0xw5xD
Xnu+ZoPULdmYe0IlAqNsdEmt4b30SmMv7sHKG7iqdUAmIUVVvlmyMDbb8ILqa3js
DlaKdbAJdSfxBrH1zThqQgxBu8x64VuvYyTmaU3yVgQUw8ZiPaMPr0pXf6PjRlU1
Pcs39p4gVPiCRPUYWFxorhGWpQVulgwMlroK/oE4yTm3ncLR1H/QT4H1H4H4q8GP
usTZtMWzVHNyAHNgzRgSSfhG2omjAsyqUjdaWsn48d82bsx6cQOUH2v7ndPCYkwI
4GL6o0HmyijyzJ8FW998JW00LJc03H5+En9hD0un4qWEuRBD7csiLyD5qukfD5zY
SyHOgXxzU22pPlzwoAcRxPMapCwxtW1i6IFmGguhSslxzRxBu3T36eITafrTQ6DW
g+bkcmnoRFVIdO995O14FPAyT6+nJQhLd3mkoT4IKfhv8XYA98OVSXxPAYqhLdLt
3UDBTNeQ7aIIqepZ18SyW3rEysfHC08phQOIq9+z1gkzL3lu23+W7zrs/HHYru+1
KUapoLiPFJ8xSEJnpRa6Te8XgDF/rF1ogia3LlXd3+rqvTSobN03s5LF39hkdV8b
9LI0eEpyAX35c+v74fjLQA4ZZiV1eI4gCvLiEYI8ySEQFTC4i6J379NT2wtkKexG
ct7WKnzfFSNeOjxdnkRkLGb1Rw+L4gNfph0Lf8bj+W4+eOTi3FbR140Q+dL0YhbV
E4W2nLePwB7a25u+2TDDKtFNnM1VOiBCSgLsEML/bXB1pyPvW4knYDjXKqWQLARL
Z2QMviEz38DSpIuujJKnzVxwJYZfqoIcuTNwH++sCJT0jfvSaM6fmj7H4OgLxel7
0+ujninZ7uLQRcXlDAUKOuVrfRWWqPMOLWUipY/PwqvSoytFevv1isaRXLBdSUnf
Q6j1+JgXThrKMo3tBX1wpH5Cd8ADeG9vZ7SiD+5ACoMOan4O3JgHbJSr6GrcilEm
DQomOq5ecuXgyQqjJhSh7n0C8v8T3UyMWOS5lDyEWOSELOXFDFVDRGIp8yy9mfI5
3dzcIzRafJRqrfr4+wfjdzN2w8hF5ZuHC6mY9iofkYTT4gw0aLu3e1p/+8MzW/I0
XyI4y4opG3OCa42gptjpL8tST6/19BgnDs3p9CFlqvHQbNPwW7jWKe5AO3I9/seM
WgHYwba6pg/w36YCW7acLQKH6OWoSYzIzery+7mOTr/NWYB1gxL/92fGnNEyWNLM
8SrOUwDrGepzoaEaRoQ148Gqzj3aOrT1vQfJ/JsSID7XUOwccL6DpjInFJhqONLD
Yba9GF14ud0anod7UUeaSQYgMH1Px3s7lpAuETCA/ttOmUmsTvcIDmAtef42zaFn
K92RogG+jLUwIcSVYUm5hIK0jw7PUPSZe8m1yhLLHRnnfU2QkQr/9MRb1AQ1zl0I
08U0eodpvaGPzOZBvsmkyOqaaA+fk6544bpnNr30h0kYMuPUHOBzdeA3Q0rQweZA
p+KZgBLQX7MeC284dDwXdFwbnqJbtz6jDDvjQFf2pWULicjR+3ruELBC8VTj70k4
ha/gAhtB899vCrWKu2lsPbQnt6QsAl5Jy/70J5TyJ69nKMt+PrFCzT7QiA9K9tib
fRe+hJIGLrbISxssl+/1XpfRcMxR/lE7Cm5LT9lBl0LOe/icQkoASH3AYb3jAym6
TrxiPaUKcbQBarAmdqx7lWrGqWxzWDZ0NTtXkN1SDayFkM6RTnh06nXEXsqac+KR
2m/NvLKGyhLKPtDmdgF8NkgcKO1ZcAr6jsT/1QFA3FJHQHGkl0Xm5gDP94sDNts0
WJ6eA22qqwKFWqPLYDwbK2CBUu26euf862itIGS6MyzeBGXzT3gmmNZl1YIsHciZ
qa2kOqdsCjPbLNjXQlFp/XegLleLo+ZfJMODcb+vmrewa7ccpNaSDUv2hZmw5eSP
U5uivsUdazncw/vD/Wnp3Jrj4vNQ1T7I56QajWVsTTBjlsSWZmwn5+o/68TJwar5
4TEzWXJR1ZIkLU+JkWOX0qFldgzzd6FRMkN0GoeTV7YDvGemsSdlY8mehFmM4+Jf
pJ5DXeGEf6fyl2CwZbCbgSPbSJLnt1gXiamRRbbkTgl+RlFl2N0DXPJVNnfPY/r3
luucfhuijYIFCUlZDa+fBtSvWUdpJnqNDBgx9O6Mt7v3z1uyA3fgyXLDNTPBFSdU
RBcVDOzmJNTiy1cfhCbLy7XVv/halu69z2gQ4fxuCgN9mS2btApLI26kB/Iy6xMf
tO2hgGnIDnBIZW4OS1wCHcWQGoNGF5+rT/K4JtmIDaeILO+mc4fTCmRjNoQ5I+lY
hMaLDn0+eQuwO582VUPB4YWWAsRaZAnB+4xP14ghLFdqXEzgdg4clJU04PZXjCaJ
/FYh+STHBEs8Dp+7W0L7gi0AVjH4Uw/Dt19ER4Y/mhm3DCsqa/9oMqdFFuTLXfQ4
5BfWLLv/vYdJrlpsn1iBa4uz26p7U9Cj8VyW2P4Z9zrsA6EcLa7Zo2/XuZh6uXBh
jySRybPePmirYWlP3s6SEOLGJ1X9tIt4+xCvL5s874rcodXdbEgheo3PRXDJNLnC
eWH+uXSw7cqKvR6rhxOFzObyRFFFoN8PwvYluoJDxqD5N5s3w8EqzZe6pIWqDktU
NPZCMHoCCT0J1RPcLib48gr1IenQSGcEWs6yvCEhForpPUgBqtS1KGx0UMa2qo2H
CtLCmOjVzQRqRYg5qPQTlzRtao/oQPX9ofgkWEOgY9ckRwdhtksjqnX1DqKUKYts
HtvcwI5WOIfF5OBxIJ1W/ASikkOlhiBQphCzt6VXi/KXsz7G8yOboPyIfzn0J+OA
wNgQoF5w4JMtq+iUGvwvLDhcKoYEhZuOGXNwtUbJ93oOmmTJfkFVB3LP6kiRiCnn
iWsr/t54Eac8+eRbzbtWOLbj4bJ4byNvgrG3xqsRwF2lcbx7K5GJCyRJ8D+gsfoM
le6N2PC1zlzilGykguMOP3i3yL25UOUhT2lrnB3knAC7pHaVvVf8h/Nx2R9izLtp
U5Ppa5YkmA3rtsOfYojucH9zIscxRVkMMjzspxRSM1gzNebMGFxFrY5gPOkWmbGL
WXsc/35Une7+An2XbknlYn+XryhAnELGnNrFdzJETrVaG3dMCujNad/9g13NSKjW
TVD6EId0FNyfI1nksk40APKcePemLOZm6lQQWi8ny2Dj70lSb9PmjbUckX6kba+t
NPuBK04GeGTSysdHJ1sQZv9VoULfLc5xklVt2ao65bT3OR2fMzDu0jzlRIwK8IaS
du4SllgWGCtzRbvVjQSp7peU/Y4eTsRqUEdccqurDbZaFXczlKkaHwkh3hU+8cTM
nC9BrHBofpRTHFO41tqHGW5hDuAWnTI9PBshgY9J74mnX8vqrZ3B/ZaZck2nmRtP
ZTTMKoWSOCMWz6MyB/L2Z8CLdc28JiqqZMl3LfShn/ZwpMeysze3cpV0o5cjiCeF
ZpUsPJHx31gw3kfBLkZkvq4hlQA0l1lXYLqsFS1KgHFC5urbH3NHz5INRBVWLbdh
VNPeXH3EG4JWoo8RQng0zxB6XuNfeZMN9ouQNhQ8nUgv8WNQPy7X3NROnv+sbrcZ
WTHiCS6BVLQaRKEJuaxH4DoKKwJI7JY+tWUCzYM92HKnksjlLkDTSVFhxZcOW0nJ
s1umOXrps1aFQmzCCqYUbXxorjhmeNXJRI9VLdfd0fQB6KHHRKkslp7UeIL8IyIv
4KjALi3hXAEKPfOWEfQQMS3l7gBF3S/oLBbnUygjRVR4jmuergmD8+3F+rQy/xGa
2wmcFtC7Ki5B5d8AR8A12IqoULiCO+a8lAEq/EK35g48IU00MwMS3nuuxBVOUhVM
PLjQq4+7SZI6uuZzKyS32A6C5IUEm8tWKO+Z9QXGy+2U/AZQhuLiVWmJrumA2c5n
aIFvm8qrZexNR7jBq8uvhE00YdLNeNGuCQHlbc2KlzDKYViePcC9dptH6+xA3HVe
S3xbQhNZdbJ7KICSVFDPu+VhZWQJ1kteJizZ3YTsgYhr45HBf1yTzx5UEUX2MqQr
FnH6vv3L5fKzoueXFVHtDq3MLxFaQPe2r4HccN8+HuTvMZU7+Bu6iMzXg165NIt5
CIfhW7U2tHWtno8nlN4WwUyO/A7ntbeFVRTOauNY0ScgKxSLACg+FTU/MsNA5PnO
qXW1yc3NPTfJ5FSC5BJ0HARAa/Im5IL0fut0A1IpBbxInYHc3+jUXvSC1xTs5SGs
C2LK3Y8kywAw+NMhtOj2YhLc2xd12xJs63qZuHwqD+Zoh6MOpQoeaqeAgICrQ3Jo
bnB3iCDToYIhoKG8uB1J/ZTXEwe+arUDy8wRF98HRHLeLOfwpPxyMujz35eKNRMv
aZryUSL2BPghCb9JK6trui5pztUIxLBaNd6rRGAKulRpA+nFzyXgvbgZnGgvsR7r
WUlgEHWWS0QMabUVmE8wkKG52HMqOoHfwWUNkv/4y81OnrdDD+j3UfUFfoIADbdp
e2U255wSVEpyWqratq6cGFJBU2OSYLMxZnpE6TBF9LWbNOzOUWBHO9llI8usvPbU
3Wvsu6AsD0Mjm0ruJ4jNrgA/wxvpFFPixRbBLL2L4rkRCM9tHeqQPGxYK84D0Sq3
V1fNhWS5mTIXMn6/7woLxdxM3of346x00CmdTwSSiwZ2voxUkht8+kDkWQIyo7WH
HM+AAgqNPqJVY12+aguPvdWPnexS+FoiR3sHecBu0VJlqr98KwEIfRShiPSkNh16
ABRpvxbEvmiNrqpQ9I7VrI3XuVbz8YckopJ2eUo4w+usQhY9MQ8nCF/SW6lpl0nG
ux2+J2Z5RZcF0u+XZaB8auBjTA1Ksr5YQ7VUBrw/BbqKx4L9NOJ1osyGNPjPLEuH
QXXcIh3BzbFugnyPKdEdkJysHrwNW7Go1jlDwi2MI9wBVxEQ3Lj92tHRYLHd23oJ
kXHLA4PbgmlY7MQ1N1KNmYPm7DyUl+mGQHSnqDJFuGXdXr2WidyOb/6xJh1zFCsc
s0j4VNOOZDtkecM2MV2C43YmeuLM9DW3B7mfJ+qbS3F0a4OaV08tzOGGDyZ7gWX4
dZzeIyU2a8P+vzoyHYRcqtxAeYvxkPn7qdzdFPeR0KtStfPKV/yr/4a0Nzy4yZbC
7ktMTy8fFGR7rc7DiSGyaD6go4e+hzlAfGR89XAEHeJSgwowdTSyjXOOwNhwAK64
nQjyGLgtlhWmu+5EWsJupp+TcpbXQNbmXVV97F4CCPzB+hGtV65B+Des8SmOZpiL
j4xy2+1FVRGIbk54wuAKHJD6b3aKwtLPcGJQG85Wq3ExsgBvX0MROGk7qLG5W/pR
LF9wgscQGWzfWC+x9qwB9N3sUFMQO0qYKByB56ESdADcaYeiJQR+jhJsDBzmHBrh
1enWblDP0++Shl0LwIWr+jwjWzbf8zsewptGxGCvFi8IE4m5VgwHqyouosF9+TmH
H4fMuOMQ6Qy3eejAbkkmbKjOzx/gGz8DiP5PLjbtRycy5PT49bxlg6jyQOtX180d
AZA1Q5FhW9sSbrVRK8/JRSaAl8FyJW/SUHXmHN+3E1mE+8IYeLa+pYwkyl0HWkoc
nzPn+CYNK+thoyOHCeQ+0PD7unuoZ+fzWFvYCQuFHqPM+kZ2+b6D7pC44pBwvcX5
+C9pHIUM5dJ7pu2eahwArWvzxhVNsocDcDXFTIoLFQTRdwHMZGsM/O7l7S33CU1V
dluzql8PyK3f68Tw3YucsuW3ucjHHAP/WzHROA9UA3AFe74jXT/hR8lbCgtou5TL
7l2U4CagOk1HsZdtdXWBaIRqo4vcxKkuCZNHQH8JzoZCA0fBNfQuu3XES5yLy1wC
C92b+pG36eDbIJCVzQu1gVtq6sLSzeDH8HSUJARG8JAXHkGa4fgELgYXjA9YeRa4
5nt8wEfHOOp8FPM8uJq5Q84Gw4Nz1ysfHD1Gr7UZaUSnqL/PT+AMy6wOzSlCEkAP
vmv/x15S/4pktZOjDiukHFhztrF4crMeMI408KpB716/brTRNSNk4/bxa+/x397n
ALb3sKoObUc6emfTUdpJkIU8wLnXIaZ3D4/hU+Pfi+6xFXDYHIq3CGhn4nrhz5Gs
MlEeDdX4hzE12tZRHc5tjLpsrKKYSwaH1llOeMuy4gwwXTmMQpg/HtGvHjgdYiwf
LM7hNDupR075WCKQwyFmBYa0YdfFWwSsKrCj53r/1Arx2BfYXtFzoW9s55bSbZQj
8Nnze1LFG+/Zw9FVfy3gxuzXb4nhov+bT84EjR+5UItA8Ths4FK8JK4Ep37DMbkB
GYpjF4RHdHMyBgKtx/juvCnzix45yuvD4ci3MqX4V1WRKyYAO7k1og82RZG8nXHv
QQu8wf84srAtOJa/A6Ucb7IDVyDQllkqc1bfd9axOnFKR5pPyunP+VYeXwFpbR8u
1bcDzBfl1q0wS2EujTYTXNNwnqu0Gq1DImgiyjlNNgYIJPHfCaWJUHWx0rjq0jy1
zJPZhkfu1QvnB0eMy8VnMFx8S166yrl2Suux7gTfkpPs2bnHKJjA2q3ea+4i7wCZ
+15H2Us8PelxC5kndjeZ1ylDJQ4fVrQxmLPOXmkqZKxAUuCVxbIxtBCSy4lvWT68
vquhnEIO0nt1doAiSyWeaBaTnO7ZnmnV+gINOnst6/5Fdh5GTGzepOUSjDiF6Pd7
Ot1waKQFrlc/TCKkti50T9A8V2l+WPVl9/nhV+ZblsL0y4zS9ooGfMC0S8uAhcYT
6FVMyOu6YS4KtdBXURSFAP1FmtsGqT/RAHpaH6anmLyjmKkvZ7i7JumQ0JP11ups
TGlWYOAg5aB3qKvvIiYQnvSU7yTJk8oivxIjMAQ3SyoqryxP503pN7D2TUZGY67D
KY2ozCcHi+0oAE86Cg7yR947IGJhYEMuKfC5mN0N8Q/z3Xzwh60wG9TboYeZtVQi
PwaMQUdn5p0/1RjcdOMq5XAMAMlzlJu5FqrUoXkOQdb6czGwXkRZgtur7OacAo6Z
3KYD0RJviVc4MZ1qMiTySJgUk/bby+WbBn52bYmOeVc/Ia2ByYAAQKGkKqribZ4T
+wWSbMdq9JQ3gMAEf2QC/XjRI60VSj8GWGwzchilnnMWX/PSKYJM00w26P/RIba9
2tUToyKp78p8oElgNFjPZKxI84MqZ8AuoP6MQCKCVbDE6NaKkgOMonb+0Js6fAMZ
GZEvdkof9CXQwnC1oJ2imxrn1RhBfByxQFkWet8X9d0qSn53UwYfdNuJazRZmuQH
Yz6SMEpyn2Jt90BZqU2eG1mllzzP9uxD2JlgWR7BbG4ZTIHWQQjxiTP9Zfp9KRBJ
/yRxIfqhoLfrcrKIMenOBwaZvQUq4d+xzZFgwxXlHT7xqSh6XkAdOT70ZX7sGoyt
y50/j/nhjCG1H8f+OylQVvR4YE9BJ716HfZI27U3PiybAY9jqoHAcjvnNHNq99oi
noQ3Yli/hE86U5t+Gk02DEFj6CvH6xBxKpt85eC5GObH4lO0CdgMJn0PUTx90FnH
9RuLZ43SbP3IlaQIStrX9k0pi2Vv5wCoLYeh5MVfxxGBPCaKaLP4ffa6MDJUDgXa
4GgjxREILCb0sdyevV7oGnGVzEm+Nao0VVqG3dWSfkzEJCdIR0v7Fb00kGwjY1P4
ksbOQYAxqZSvEhKDxP7B/CS8IfZzXSAt10/DrYmjHjxaIhgo/CFYoLn3JMEVQXd+
+V40qUhOtreBUwa0rmWenPsDvuczcLyjXnHmU5OT/mkqDtH6KoG0DQbqDRzeqpeP
fqS2H/AwdUMQg1dCp++bogreL8NSIY0sZPnkBIpIJPMi5f69Ur7l1gIcnRVtV8cB
FwFiLojeJjWNyRYQ7MPpeUa8bgJzQ378Cq+uO1v28iBED3zk7rk02oBkmlT5FrzK
Ruq/G94imzy/jDUqW1Hjlqw1k6nfqDIdjgDrsJ8vMuSpp4ZCvqXDDzZHq3pZziUG
wNYGKyZ0TVtyds4gpzLPJJTqNaWKPJNY6peU7zFoFtQYBy3v4bpb1hRb04ordDHa
0UcvAbAwVMGKX4CtnX8MT5IUHs1ij5+hUI6J4aCPXp0iV9hfTtocSsJg26Kn38Qr
E3ePpO2hbM3xFZp9aShfimVkJ+ASjUNxIqB4JZU7qzSD5OrIYPJeDkoQG0LzqfR1
SUljNHDUW8GYgDn3dyMlM7uJBx4jXGrHmx1kDQo1jMbabTxBVQ9jjXnFlEWCLyKk
AsOPJLJA2Ze4eBU7hEmVk+NEQYlyqzeCABHhmRCo/BQO2kSV5EfAxFAyz5elZYrU
otoCPae8BOZReJbXTxVOHmsHDyBiZ1Qd+rqVd+9i1BJQ3Uti68ZwQ+mVp9SFeh0f
ZM/0qNMZF0tRVnE0qOZVHliT9pDhm2yY/JlmCCBUrtM+gV7J36jOzZaImflIYbPD
mnZ1W4RrwglFd0QVENQKY4J4yQiRSMWmSYNMXuk7LN4l8Ry0DqRICmLqGVsiIQqt
Hnm/L80lVV2QvuGGCEwfoWMUy5bHtDCVyQOQU+BEml0dP3DzPTlbO8029wL2M/du
Of9x4qqgcbbV3vvVCt2Ucgrys1BqkFhkG3t/ix1j+7gp10xMIc7DOdTTZAP62Af1
30jcwxHxAqPyyAzhPtxqq0TthNr+6QgTtflG//4XRxmCEfhYyDqO/UqH20Lw5/uT
ZN2pcVQez2DQG1xlXrpAETBXuznFv5RJ7a5VHMs5Q9+wAU5lGQUXxIle87/1VzA9
laMgKYrvEbHYW00C7e3o+BrNTR2oF3+e7IxZZd74u6QorNL8lhg9iTxzmTSjUMvI
N9Zv3GQSpaEXBqOIpKWqXAlXHpQZr9mD+c3ijysugWJIse+Uiy+5dYBlmNqu7V03
AAp6iKVSGps/YRtOHYe6wTQZyMnS/BcsFtuKQKEINjRhXMlvaQoQT/QWURqhDvCJ
Df6hp5TrvOp9VfxB7B3bIh/aTx93pCayve+2K4sUcPJy01dsqsi02qTSANFvvyBO
WGPYGl+jrbad/4iLsz53K796/oCxmvGGw59AdnIjfM4u5JjOuBqMyQETi8C6rMjK
C84PyuzyjEGciJDtcNrphKVqpiiyTEv16ECOWxQoKYhT7BDeCr72YyVt0CqQd8v9
yjPI67pPTkrG6cbvMaEw01qWAx351q+/ngN0zFlCR04Sjec30tG6CLkKm8w9dTaZ
2FnE6ze7I92Uvp9hYPKUeQsxvoi0YFUJ7v8N0vXIHRiQfbxuOup1FBp3qI9YTums
FXjPT0K3g003/PCzvEK8YggILN4lEyhHEmjLbuO1CU+QrSoFDCJdIR01r3XLZe8n
G/NoHJQZvI+UPMS9nl+87Z/26Rfb9cG2Iv9DHhf7RIyqL8q7TDCStzYnhmrzsF1M
xQ7oe+Hbrk0ahv9N1v+jTiO/YIqDXWSIK4eIxOr1mR3wxIe3mPkZbcPUYUbZZJ9i
TYQWsdnIIEWhyw1SZan4ECl6iJbmIKCAkpzaGKx1rxfM0UPeZpBDezye0U4p9F38
kcl3+WH0GZbfMssIFrZb2bKcn+9Z+M32KTgX/0IJ+RHq54N+4JjMie67jiwsS4MU
YWpl+MEIjkNGBYCyHw396Hveg+SBCVJvZpdwjTGT0CTMdcauObWPvhb7pE1VrwiX
fZoXovq1hCjTB2Ud7hZboO4nwgvWz0fxvbrneqT3WO8ivtPpkdqg5edtwgb/9ovJ
gtOxSbHs5rbCloI8vWX0M39ICnpGh5p9UrNtdr7zoGMTpFII12rzVhZOVVDK3TxX
LvVtKPOqXP8tIC76F0kL5a+Rq+1LEQSBwNXAs0tK5o/MAd+8JTfLpal1C4PBhgyX
38Pcv6o14fgMqmedp/IAs1yxHgA2aJzGyI6uZn9VoMhfrTp3jUazfMKegmeEszoD
9eqYeuZw+8lKmdgGkY3LdBjZJueRfu6GD9fLvr636HW1YhhHNQKPNxd4DOr0jPgi
vGRqtLpmB6gg8OMOm61zJmJruTsV1pJoetlAx0MB02J1b4vq7p2ncULzb8kTd1NI
kz4g9NjdTWMELeqyqtwXrpvglKx559M+tFumUF5WUWjstUp2hj/hdE8/Ir0Qb/RU
kyLuvd+czSuTrfOt9KmGiTOfEfrgoFlfAaghKh0hmc1Ajbq8mL9KHi1EaHx6dalT
daofUyJCLsyh5M1+/HhWuRe1RY7eMZwp2Mt7dGATEYfxV4E8XwoiKpQGDy5YzkCl
ypwmf57LVyOYcvauV+iN1QTI7d4GC4DatykMAdJFXjmhPbSigsmx3qnhDRjN3aua
+HjlgySMubKoKqZa0xRw9ISzH3+lrVOlLi+RzKVoK7713mW5vnJ11lxfEjmm75lZ
lOJIeaXQOhBGBA7T6McL61wiLP5Q26U40SsTX650Or2PZaGp1AGMB5E0yn67dico
xvq+afzl4Ltppc8DeDPTkTqAM/iy1Taf4JTUQjqZB41btfv07HtTfE9XEOHCHYMC
YqiD1vU/NOHjRYoc4zQfTbU4yb4/w4Enn75lUAqjq9EFsXZ2rthhZdC4XCli5UOl
eWxbNt1yA6dGFCf9dwtI3eWnMujtkFS2iZ2y1sch8hRIYqlcip7N9SIQ1q7bWYEa
M0Dq+Nj1vpnGDHjOR3JnBQSaOUmq3D/1nAFVhhCtuLmqe3T2Hmzv4JCuDy2jDC1b
K9LPN8ccIm/ATqGWpsAR5Ry5pb+N3WqQSPtYl5Tm9YZBRU6ywASXW8z1Cr2tNmlb
gAD7L2ATkO8yG0mlxhjkNIZ2bEU5z4VvAg/BapoZeC5mE0ie7RKfrVlrm8QMoeH3
A/zIg0JOvwwllmDRZ5i54sFOSRxGdYLvCeFdmMwB59/6A8YQuzDxuDfxrOtAxq3A
BhIg0wHRZ7rJawB0fzq0YaC1IZRmZ/voMi+4r9fdylcFLbd+KNYh0JZH7Sjxl6yz
H+IA3Z/xFf+RNLcbpxoKhX50dSWECTQOj8meBn3HCORLsh2LFoCisM3nqZhA/Ze6
i7xH0SFgzuOWtXjWU65kkjcyeMHltwhHo0m9ofhigeHlIaUjYOcCi83el7d5HA5d
XeI6fFavmbNDhxtndA96eaUKcDoFzkwd1fi1TZAOz0sMvv82ZpesgPpe3Y8uajyJ
jqSK821eaySyOVFogu0DSLDLBq+7mPfDC54U71Lx8jKCJdA0h5GB5h1iGivRahs7
clKZza5FCNeR3lFQAiQ3s7csnZjSa0DnXKpxPVlri5oAw63OfxtBbC/LcaLwkHXu
hrQCKNYa3WL7hBDQiUhuJzmKFgAL5VM8fDHv25fd/ezyCWmcny0ATDy6oLy3oGn6
H/0CnsWTzViXY4E8n9de//HEqEPslX6KtPS9PDx/tmJ6vXpDTuA1naqWAfseoRoG
bvZPLNoKIOg0MSvAsYwuWthYu4WuaA8d+tadAI1NOJIqhnMvDYqm6rZYMCO7eRPn
6UixYDfh3rPI9BBymSEX8g9FiLM08OwhjM5D5smssxj/Cz9BuZXH51gS/RihscNd
qOIklGPZfVCfjMGC9p992Calpmd/b8hSUDYXmVj81T2K3zO/4ZWoFH51d4NMSVyJ
MUvfrUB4k/UfnpUvFSDQdGi8AZlU/gmDKX0TS0SBs0pnA97ASSv5GIwbRKLspy/m
AWa6RTILklS5aq3dnVb1W6dom+uinC8WVfdEurRsssOe9s5Whc2Rv0j4hvssoxI/
xgld/dilPSc3zS+ffpxxG+A1mNst5aKJ4CIRwwiDYWm/DWD5hGTViWEcXpZR58kM
ZXJOg+ee+xWoyEgonaQVLDAtI9PlHJaN5BbW+Df1rlXJjEuflS82BcsJAPmYr+aW
QFD3M+sVPPTWWpEO+sCw7fgO0xM1kjyfSMuQjOfSAZl8huogtVxXKJj4YyQ2t/Cg
T0n7/i337S9HuXwpJyKfNcNCXXYOp4n7crd5C6hIp5/BHJNZgcGowRDlmQufyyQA
3eLygJDV9I54Y46yINdOuCATXLSzBfOoyoKZZYopwHmtAyh7CP4N03Xw6pAuOlgk
cRUMp40Jjhrprwx6sZmhdynXx1SQc9t3s58FAqbsK36SJvd0Ow83JFOnrkoQrY13
rH4QaGslmmQlwTzxu9EIGuGsv//pqrQAh/BP/GyQMYg2qQZyU7xiC+7TGrUz8t5l
hM6Kvyg5t0X6hV/VO1WYh/kdVHSuK1Hv9gL+WJCQSmdoVqcpHW2O2IDxkGAWT0/r
EDN89CaQCV6I6HF7U66SLzDPLjEQ68ENc2KHCCY7VcDaG8vGIsL2e0BlzrLw1jkO
W/aC6TWUkkLISkhJe8T7N9/FKAKGw+nPX7mZBEzlFVDwjd5czsFdpTO/IbL03g9J
PxrCloVMjIwuUJ/VPrMQ1Ixl8CGtAajW3afFbmgVCShqfNJR71b/HmyNr9kuh89m
/Gu4rc+/w3wSleKAaIQOr+NkwUGaRuTOAirilDeq+as4FfpnS05LwU5rHzM+itjY
Q0y3N1rXZKe8Pcu0/iSjne2Kl7D8hWmfWr+Gqs10SfzKjN+N2wKOxbePuZdRvFyS
NFRCiGjHlBpqZAzQXle7LiWtjXgq0sG5CVTvyZwpWIHQZ5B30tduqw5nBUer+ccH
c2JFXrghZocPfigB44Iild8jGhpjUhjt01iZpREdahmRQuLPlUraTiAtYUDwf2Ao
hbzeOB66wPsZbFSl7Mx1Jj4g+/quDIV27/29AZH5RQd2H/iHAfjCIjVr9WFmf5XV
KuobOTk5I4WomG4UpfxH9A6H0e3Zt5HuMJ9qii/Z9rk69PjsDteZHGjIzTLhE8M8
rVDFCCE9n/2zRzeniYiWkJ/ifA+MV4MW9U3I1ASeCTY9Pq+6tsJ6cvGF03oVsp9H
4qhi9HLzLVhJBnmpj7Ah5P8A62SVF7MzeFP2oQ+5AHv+Zc1d8CHMGiRgN4jS/SRh
Ysx8td/quM3379Ho7Jp7PCUpHEToPIKG1kP5s3QNHGgikkPJea/jBZEQ5di4qDuG
oSylL7ylfeU8buPf3zD9lHdHgb49wKmUVU3QlTWUenYHCYS8dBzeB6VA2qyL/B3s
GWmDsgIAfLldf20inHMlJNKG3KGUcR73p/3BWVks1DkQvyOugkPtuwMggz5VuHwa
Ya2aDYS+d5DQ2V/a6u2EHI0/JEy9RUapUwqQNQSebrJCCCWlhNkR8wOmPbtAvLxu
0hU7c0gkq1FOAG7AAHicCt8tJNkgAWz87HG8vZn7Voa96MqnuCJ+4dfgFUmM91lF
F4+qrYy9vaixreIzmwjtbvEqJYu+ms48mgokyfjoj2KCdlTL8OH4DoYc322QS03L
XXj3kpDkBNC8ypRDwWN67yG3At0SxzC+2UWjUmFvv+4w42mfAyjB7OdM+UwDtUxC
oa52hO8AxhLumiaooig+T4+Q/9uVPfU76ZDM9Ba9vtGl80FwbJJLksljxmuF9ui4
H4UuDLZvIdIy0S2XGBeyIEL+v5JGNxiDJRYJOiO+8jh4/sxBh9JCRsFnAnDiDlkg
EnKxWqV4SXWdzyI9VWyt4IcKMPiqkjmIJuuBHTIiFN7CpEY1buCdXNwWLyI+HUQx
immHicu/KvKAzmWI3uD9QG9Z1EOuCHkZ9fzfgpsSQKW49BJC5n69q6oZvc2wXvck
ACaVcE07goWa+VyK+292RKZl3M2p3lKICNlkqcYn97Z17Mztq6k23u7N8Nz5iwgB
b5rAOe25ifADbWNPDV6EP4c8MHLLFUGEF1Jp/zYgXfezcpxDX2eBbPRJz+JLbJKn
tDJtLiHbzSNnwjaswgjSIzGvQRwPH32AQUWiPs/DK9fweWNC5aKvSxeFncfM/V0y
Nnw3rsh/rFUEWBg9a0Kcxsvf4gnOattdjQvDXBQLQ7NBRUbcZWvGcRn8YNc8/CPD
fW9/kzkHsmsR8rlCEJc4GQPuDePxXwZdeu4IRlb+HegDVDF3UZ7BAFyxmWd/55sr
AUwzxycYymrZt/qX+oMwsDFUxvZfKGVe8kA7EaqNh5iJRyEgScvPEcXVip7agvFM
iaQHUpW78AK4i9Mi5ruKaQMsT0Ua5jIPBUvPl4ffzSHmvyZmg5Yj+OlOHP8CqenQ
aHsBwOrSFEVkth3Y8K2Dij+XYXmuvthnFlJ9y0IIKeaODSv0/cpsbigHrghpHN9f
YDTnzcfwn2H8DpzqCgY+YRG2QKFQn9cxog2on5J3a5LqQbtbeKj6dE8gfj6jeTIr
OYp0V7ZOoKabVmiHgAviml2AsOvB+N0G33psqviw8B/dHQIlP6P+DSkQE6SslVJu
NfdO4/Z9Wma3FtJbPD152WHvRZVzmW03mmfBgPKTWojtukStGd0buIe5NrZnV0+F
2epZIjFZDFpI1l6qyon2bJxOrCGcUlVJ5kyGe6RJ8zTjV7f1oHAi7r2VIdtc3MXY
dVz8lefiYqqBXDMtLApK8SAu9rnKf41KHBvR8UFVt1t1IGtVTME9je5CGvsX4Xcp
nHl4mQMlAQlY+9gd8pzE3NG41kRFqlvyoEvqPDUqTw1Bp5qfH6ttWb1Sdq0EnQn+
KN0OzjIf9Cigy04q9UJe3QTQJ2IKFckUkuvButc5ibAJK7KnFlp+k4KxX3uEbHO+
25QpTV8cdBpPPPnxAtdtg/hkfVwcHHI9454RoywHQ1QUfclo3dbtfFnjJrY4jMEF
m2v37h+mPvyO2WYwwrXbTOBTVc7ROc+FwwmpVkxQewbZGkGl5HlP3sRWxrleI4xq
Xrz6L9S3zC0xr+WRGI//51dDHVUNxJZHHjy8fTCy48ztP/TxzgJCLAiZNxAQuLBp
KnhCtiE7Nm4P7obyKVhH0eH65qxFoYPXux6fXOy2L9mcVYb2ZbpKlPvSCng9nV7x
Hhrxb3bIzSSbxIVFqj2JIF9gQWdDM8ARRdu2b8MyPxVtYiiHeamCdaQUWl52aBTQ
ymcdEEHYunFT5Yl6jdnIrLry6nFUSerOO/blMO78RT5xKr0eX3XKsu8C/ugeMleN
h+pvnyJSDRLsi6vCYpPcGyzeOBASmT93G8IbbHDfLynwHHwsaRkjoekkVmNSmtmK
icVLxZ1541zTiynQ9ETdsbagA5ZLlKI0Dgnqq229gmIzDtce2VK9d1HnsWLGiySc
HZsgRZk53e5cY6FrcWIdvhhdjHZiuSl/8MZpbOlgkSKwua1zZPrA7QWiA9Z3v98y
IyuBWfPnbp0YJXde6VF3cMc/PVGxODg3QIVIjDddSlx/xREoyOYnPiMBEIpjgFQ4
YbaZxzMLl3YFeTpju6qIBfZ5sTzB+hAlNxj40R2nyqJ4EmBLqcKG2TdJv9+s8ugc
iwAboM1XfNIv6gLYUoiRrMuuod38g9UauReA6LnibYwJEWe24v3zCu2K8b0O4pBd
e/5suRGfOMx1npsqgLQUU10glNTAh1aPTCTw1BfaqX1TsbMcQzgn++iacNFAvKKG
UnnO2FRpE2eZqlis7EZ6ccg6sOYYbD5ORGrgaRR89Abkcj1k8VNFI87fTMIgWQJA
Xqf9S1TYg2gCL1KLCPXBGQmSLB7kRShEdnqZQgWH6kbHNABtl/6ycFPyM9Y6wHi6
oc5HGeOFkphZHesCIAJrKeIiLLklgk9IyZLosbTNauB9QvmfCuSrMnpB4PgYo2Of
sAsCo3jn6l748B3vPxO88ibTap475BJ9asEb0t5YYJZ3ZxHQJdyBwGi08fbZV1RJ
wsz9wZo3AwtvCrZ1DLqdGL0AX+W/8ekiwaDgCanfKipPhVIEPH21WXRCdqUNZhoD
NSrp8nCShv4nXzEX7AY3hNEQNFK6Dmua+ID40O6bDrPsQvvMSnFQ4MN/YVsV3yAi
bg9ILXyH08aBeiMd9FNNvfZfpTybYSp/vwaNAb0MFnacavepFIr78vUF54MmQCpQ
nucrWpY5x440KoQLN2XSv4azSDI5JXBGS0J9nkNGzT1STyCmzrXTkz17GziLsmkw
mBnze4Y2aKhJ8p5t/eprOcwPdObeG/qOyY2FnScfsG+gLa+bJDr16HLPOFeBYN2h
bqScjft5aNpwbYbvI5kqRuhv5u804/FCIoVLDTyx6E8qzbFsxEvbvrr1KF7GbJ7K
MrBG/OsLPF37bl9PWrKzkCXtWsImxnj+3/Q8JZDKAmKzHGt0oquPrFpt3GZFzf/j
er7/b5UHfd5qPSKRKFiRHZcrfU9UcvI/GgXF9Fy2sO3gYmHPIlHWIZZ0xsmx/WOl
J00TUvRRiKeeJjgEPzO78WCPNvAgTlY3QCqipDlXA2x9EjQnbRv+RhkcQ/HW5rFO
Qhj+FApMU/Bw0dUZR0Fea2T2woOpuN3C6XRUAFPBNjV6KJcG5OpZ7LWmwnHFiPSw
2gEU1vUhXmtS883+1Joox95ktYrMrWNnO1cgr4JRXIPoY0csk7JJFjUOgrPZ6g1O
ixY0Ac97ZIIJn5kp3b+X/0Tz9hO/9icFeAt2EMDWiaT/N2nnJFkfYOnFFBLt0eVV
/TiGwpy5fbnOCr62S87zxgbQeT56g93921yREn/CaQwJgVYp32sIECruxVuMAZl+
BM8Nc6npFnkwZnSY6DSzS1RGsgoRUIhjbNtDsHNVK+J2A/omyjWyg+/HWQioH40y
US9fXNqpD8/uZ3xvrZU90+/c9W6uIL1oLNgZkzxm8weXe6Nr2omzKvd68RNTIN82
6QOUkd5jyJ5qph/JHiqCEUCF/qbMsBIgp4wuOTNDVqn18RMt97GEBNn9W1/jwKPM
M3LYY+7lAapNJHWfv28gJL2Z17QAMcWUU6r6UInfZ08PyN5VkjHd0vAkjvQChok4
e9yci2YoYY42lqh4wDohaNlBsnBM8EW8azw+zLgcyadpVq8L4Sar7Yjyzr9Sj6zO
vNLxDAefxEP06lEo20O1L+EnLpB2o9FNk730eoHTSIox4Hksyb7dQtBw92iCuNmf
hhQMg2e7JcduOyOoORBiXEtIn2nTwM+krkb9MgZAUir+zev5GxCpYCQ72oeZaA6v
A3EYhgxfouuKWG0fOrekYL63/Jf5lf0txniBMS5MP/AVXxGyJoLDrnSD+MNAxTGe
7tOPZlO9Rs3LbhDchuf66YJzre84Jg7hRfE7FAmv2VchMx+2dyeLWOz2uP2+HSmE
FHSEn0buxzzVN6GYvSVmUXEGE2QcwmgZF2bkEl814IEjkyr9SU56fvTYSOIZ5Da1
dpT2Y+kZ0upb77M8Pud1FNkRmH8D3aTM0Li54ulVCHQpFJ5kUj0LzRYw3yHCreOF
bDo0AXRI/V2PVBhX8cjM13+3uQV8dwAXY9C3kOduYy7OkuuUiB5GLnP6eJxATDPZ
BOpVDC+fiPkdp/as4XDNCiDfQct4rM4+z7KX2veQ3/Q43ENXlSqgEaoF9b4iwjKP
MHBUvo7peac+fLkb4xe6qVUFrlRbvENSuexJBWeJRycfsVd+36iZ7Ox1M2A8MyE4
jpROcxYzhDJB6+hREnY5uEiIVb3/z8V4OoqxYTWe5ft2mI1Bhf6Do7CYx5CUN2ks
oIy+YPLF9kOwqPV0eCjQJHT+lYXNzIpYt4nyxKpvvxUJziAiPseOZpIQd2hpj9KD
ZEitd/Dr1sEmqPrOO8ZuzBMNabl61pBpsSIj8FeHQCZB5YbYszsebIBjyR5jtP/0
ONnq47/ygzEi6WElrog4qvveyLfyER3XF7xLQcf7OXkRBpCJVqTXBZIbZ+PUv8QG
G5Fub75YT53Fy0AROHcNB7p8L1xcN9gF545ELuIyG1960+sq+/W240EiquPgp1gC
JSbomFuPTnPuR5PNjELOzCgbcqaYBYBsZZmqsvBWavpXzetQNiZ3U2uThxa74Qbx
UskbagG6Fn9kE1IpLthugvx/K7p4dDpq6J4qnsvzYXJLEiwY5Bk1iylKuH/rIBK9
LT5DZ9IfQyrVBU+Ji/gHVLX30lAy39BuhdRbiGjeItQ4tnyOZdLm58n4huSBX+bS
I1O/Pfs4SzX40sQUTpdBna8GetHTKvMW6+yxUTO5yvM=
`protect END_PROTECTED
