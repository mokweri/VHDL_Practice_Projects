`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f0OnDgNbter34YBcXzWwzpxVCgBaf4s0AIjspT6Re6koRMIbQ5dEK2dJesdp+SzR
lMUTuTHAAdY+sCglRTaRjaqSb7FgSzFsPu1VwPtzfl2FdRPXAfpSe6uNd+w/tVAj
Eh9NWHZKlAMoX/kdaWdXykbFNZHqOhWaKtdWZo5PHQ3sZ4aWrV3GL9g8zFFEIs21
ydC+7ElpH+HZv6se0lh314c4mhbm9s2xetxFpKCSfTT4B8zjL+Cf6LHcMqMPXR4a
MbgaMwsjV+RNnA0L9Pee7ysoU1kQZ8kZDK1fiQKfFYCCJkPrwQxELa5NJ5nyzgvV
PbOLZw8vLqUC4SpfDNwfU1grmzxo4CMWnIpCie7nfcA4jdZ1Yc0Wq9WaawLjPrLq
`protect END_PROTECTED
