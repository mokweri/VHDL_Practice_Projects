`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9cpzVlAjvjHMDJjvZBEQS989hh+Q0foBscOQdRV+MbI1NGr7jplRLUrVCDJnK7N
qFIG1OrRiBbnMQukJggPLIOcIChWuU60jt3wT21ZOTHkxpdOdnv02DO519yxphA8
qzkJ28seW+zYA5OX4T34p0C+EeYPRLeuFh9K2+BSHsFoGQ3BxdDhJMQqU8R7mgGV
RqkZdTVwJNjlV9qRCsSzwVFgpH9XdRZLeWOFNFsBa50EsHd8xKOyj7QMl910u1eE
59iVqF2SaUodzRl4V8A2G82mDwK/Ms4iYokoxWlsZbee/D2pIA5agqmlqlP8VoF3
Kbya3Pe9LxvCpOQjgYk89SZ47iAVtxtQZRbSV5yqu5wL8LVDld1CjCfMVFOVf1BH
X7tM8vo/aOGPiCVTIj0WRB2kh0r1BVVEEqiWg+Hp6Uzkd0sHJIHMcpBom7nr/v6d
`protect END_PROTECTED
