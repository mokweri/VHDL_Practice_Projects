`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCkrDJ0CEeRGQs61otNYM+8v5BWUSw/zp7fOWfmAlgrTAcueyWw4RZ8fKhGBRgts
MJp/1ehjO0SqMVMZEXgTL0xVQevnc/ufmdOMd1sMqnDkBpnrwRE3PrAF+I72ySIj
HEJKy6r5i6YGv7m34APh4UG+CzGdQfjevwa7t5+0PYDGkoAfhnPbB2fWUNXiliMw
0VkqugWJDnePW7X7V3HzUPIJTEMFjSTTz3KyBIlDasSsNTBM2+4Cr2ARh8UgApD5
b9RRxwAL75wNRRqh5kugnLM7AJG/12m6Dj8gJYBc/iwGA2Zn3UitLzBDJhza3Zwz
1UNBeAx9cI9aeRc424e9jN3QDx8M2Tnt2eqSjTwfQ9Q5XgoTTxose095MliDXkF9
MnsJLu8LZhS6Ags54HvxVBbCcbu8s5hxhGnBi62hLSDWFdV79GWS0zRdYbbYwpGQ
z1hyXTwirlU+J/VXKWc2V3QrJxqg96sfSJylcu3WxwAj2oevdxUwMJ09KK41dm4T
YjxFN+9l6dvwEcUjq+WX+leqr+UwzuwfG/YyWwrJPVUqMS5GJftHdcWnZUzCQI6b
QhikIpgPyFIDGXqNLG9wDqq7RP4JFHcNNyT+8bmV7yw33b0LhuKRCtCaw8lJhFgt
cOCCEkYx1/Bx2AFlyhXq/a6CAkYMjr+B/hu2TcPor6bG6Q3XNbe4pKDuac4WTe+J
ZbI4prMkOOm9Va6C1LxQwGSYtdI0Hz8KRprpaFYVdm8RjpS0YU4Lg8W8kjtGGw4q
en4bf8cKv1eRQFFXTjONxzNacOhxO5u8NJuq+wfjfAVJz4Pz+EG7hIMzaMIo8nwM
rWrRc9HpnYd5aDpRv3et6NaEeTBageRwFb+6om6dPixlflqEcG441haQd4FT0WIr
IMzE1DL2E/uINAerHn8aYqYrCKjPZGROCN9jtZbUUW7usqQTY0aM5uKlImlnnu2q
h3wSL6et4MY+ItvmOEFoPkogi/x8sFCGp7eQij8EMaD4WhOFj9/0XtXHdJlw7R/a
q03J7LEGQujQBZZJAwaQbZ1qUbsHoCvZxMrgcpFbVpVEauOEGZWyLtP65U6c95l5
N+E9ABl66rR+mERchc6cHWG/inXdUUUbB7v78dQBJb/bLBEMVBmsBiag7rSllnD4
OMgTRSDSvmVgep21o+D2Cvy05f+4GGQo9I+ytO7/d/U1MW0GphS39BylqPLlpToE
ynsro+15nRiGOY7wOgQss18ZlhX+9pwqfZo5DS+OVwtOAGMaXotY8xb0eGvGrvEe
P0EaxhNOiNCU4PNECXY8ypiKvjxRZtsWubie91BgHP3vNz320dUyioWsLJQohIcT
opf4x+eJilkFjct/wj3cJLViQ+xoYwnfBG2ppD/xILFN1rkk/+VGhpczVnn7ZC8c
Ra4McHKjdr/Ef46c7s6K+DM9Koqm7M4/fS9Fm8xem+Y7jWhnpTlAs4qEFu57iOBZ
CETtpWRmDMAYvE6+BHX0YREp7yz+kTcSjLnLf00YHk/gGB6laiTmJRb0xHbDTkoe
w45ty9jIVzHape1rGbUp06L/Qtm50f+/i7R4gsgqnAS9xxmW0Y6BQAa/Jv1EXtiR
VP60JnIovyI9gv6u5QV8U2GnSH6jjzGtNK1aux9XMGyiS9YEyG6JtBLypSyNzfax
C+p1VhuhJgKC7LkgsMuBS7OHySmXhisxB0UtZmYLT3Rzk+8MPWQ7cL8lhkilMs7m
yKCzaHJPtd9at7BBq8hfxul33brIEJBtSF4BqGBwqR2Bc08ZEJYeXGn9HT5QVnTs
W/JP1TZcuHKHQSSntzNE5zyPFwbiCzXvZV4yGARfrFxEhNbLugk6O3CDcHaF2h4K
bnuxBcou544oCQuzNezL7J14ia1zA6b98uynXKO7pYSOyn5cPg+sk9KaV9Pn9hx5
PKHTio2StrI5aLLw4hlVt6tZbEJGBLqhqlaxHFZPRnNocZrUjkTGR62ArFOCIrFJ
UWaAvimciHhDmcimvExypmuyWpHCa3x2vR+Uc4ckaUK6MmIa+kSGJ5Hk7Ew0o0I2
urmJLVFiDae9395bTM3IKG1YghqAUfkyfH19rTmbwOudavhSguLK+tZtj/xOgCFc
oxyoxhy68SJDBN4GsPCY3EF1SC31TxYdQ1p0zgWZjnzFdiia74FmKhYPE1Jikq7t
NAwt1LBC12uHpxeCyQiOF/ADtQP7EgSi6EuUy2SiD7hordO2F/cYV9QGbOnxcuJq
3sbxdOIhAU20U2mOqtNdeK247W/Ft4bjJvh2258r/CNYhM+g1xBYcz+dGImYa3Jn
LSLxmiwJLxdsUec3Zdv4h9IAE6jNPyeDSRjsBvakTgWZRI3V4DFB0OjAgWLoQOcY
KE4HZY5/IAigiy7HmUPeKFJYReHOfwMISNQlM6stKVGHhltPCoFbPeMFd65wsB47
MPFHm8/fY+iUcyGGfkGq5c2CZVBCIqXq67ELyDr44YuSjR/DYdfNojOqO8tUSWR4
vVeH5+SPmUP9c+ZcLncv36lf3i8JCk7V8wXj7WM/tDm6lDJ7KIyH1wIxXBEZEWtQ
PbW8hNDj8ALYd5AmUGCe+K7m4RM6/5Z1i1v9sUifR6uLehw/30YYncx5jiPwlr2j
0ALzQbb10wLFLP54lrI1yH6BbFuKC8gyAm5EVnYvn3wd9C/BmMpefqTozJCX0SKB
FTm8UV+LW3w6uTNLHoRfznxX6yNUK8vwxEHdNp6u9oO6iP1TsQFr7bDURW9h/upA
`protect END_PROTECTED
