`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jPJS67Uzc2TQzU1nOK6O5yZ/d32KriGhDRgz3jq/3JfBqpU+pYWjcp0LjXQfpCDb
ngNQ2o0+LBDo3yPD9T/q+mFsGSfGt+7o3AgfWPlRRKW3KrydzObjF07b7BVIg2SG
q8AZwqo34RDdGiLEH2J1tLUOdclgkrEKapeuK2f5wuMFt+4L4RaAh3s5g6HstFrA
yLSRIDlOvs4One5UcrSq8KslpcfWKz+m9Llf6v3rCIPG+sQHf9Q8w5266ziDZfRX
T8z3A02V1Ij8LR1b54hhcx3efzDrGMdV17sF13KgGSIVTMbfm2H0c4zgFC2MkMP0
WJ6f8EqgZdiGtCPlZNkMS+ANaTEtFjrJyktnnzeGxsvB3hjw16p+TE9qwxMWX1yJ
IKVPpL+/GfqXcO5zqvMWzncbTwWFL6/GkIWG2O8q2dJoiPKs1mucc58Hf1P6LUWz
kuDl1qaBpGutdGOO2TtKWFuNfFcpkGllsFAqVbFtM4v3KdTgmebTCbxOAsfXvYNF
X8zXopxS8kBbneANommNkF7usSMPiM9ldROycMDGbOpHmON5lfqTcaFqDOa6iibl
PG6X2+bbXKNIS9LoCzKGZB4knW7aoEll+H/KBJFG2HRR0CdOaL/kL6/vPV4M1GKL
WUJXBqOHfk6wz+m1bBGDkxWRjsMOPYnOeullDyQc2Te3XC85Bw3U5VuYCVhLef+l
NlRt9DlQS02Xd8D1QwQPujem/FB2CAyBJqHOGW9uXPxLDULig1z86+GYeKEYFmcd
5JMd2kPQf0SwOs+E8CYsdUr4gZmBSAwwkXlo0IFZqgKfRs0QoTul5CkAKNyg4mSB
pv/R8OgncUfcWUvV7XB+ViEPguSRzBMW39dDB0WQm6N/cZNO+ujVkvsYY+JKGrN4
qM7OUlxrUS39c1HaC5reqteEYz37F05ugdPlWtinKGDsOF1wNFQdQqtehvl3+Dft
xLXt4p5q+gm61+jkPinFx1BYQQDwR2i4uyD72J1LHAyhyNwcyFroKOaC9V2ttWo1
rwEWYjjjw1ifh8VEnzdxYk0wP58g1b0WcgDoECc369njR7A61JcYYs8d0r6hnZ/4
Rgz96AK5A459DccfpgBgzqa4IgbzX4pt28g/seGOWfPo60ZAZ9Iv653TxukJvK30
cMYC6LT7VF5AS0yFx/kZ9a+yVzusCHD+nOYuuVgmfPu7ZP+bgk0UoewttP8St9bB
Y39dfxPEsoP0jPCAiaPZVQHqJvM79AcJplwuIfqQUkbLZ3Go1QaIAjnb3gcaQ8J0
2T7c0/kuZy7RiRX8WQHii/5xE+God9bGJi34hv6zRM6P3bRG/jZzjdKBQKisMG0+
SiwmyS4hB29Wey+FlfL1y6T+ZRhXRZWbzHISzUc850N6UvdbyqaoT9nx5ehYarJW
m5q5wfTmxoCzfV1l4e3FdwNNkNbuLNgtWmq6cjhqgQXxWkPV2ViZod3el2qltUvL
zFAdDaJx3ji4dQ8RyThkpJ871mR5xpzlYMzVw8113sZveiMc0dKuv87kYygO/27x
jFtX1mVgOb3LyAVLFjX+6chaGnreYl5GQz4Aq07Gm8Trq636l5wUx4B7+C5027mh
Wx3eNRquM1p1uAk58oi5orrt3ZkABZN7J3Y9ipHP216aHBhWRW0nrGDFRCnJ1+MF
HSNNY+b2TBCfvTZlvM89gkU8B2A2D2OLP7pdUI2ICcnf2yUNS/mx3xaQRlarcnuy
CMwazCZetcdaJ0n+ykRUJ3wPynUHxzWWQLikxP8X9jmcmUDBCsNzBJcMOgGkiwMC
Ud5S1nR7vN3pTLbv0JHtV8L2azIhX6+2hgiHYkeeJzr3FBczEj3Ci40JwGEveOZv
6JmSUHHVCJC9MijXerZGyF1xxBmFniDUSF3mojXHOH2waiaqZdlnaFIArmzFQ5ax
bF30hAOeuYOractt/3QpA1p2hTtiCGEesUKWk7ECJWQsC7nvrRIOiRGM2XKsN288
8XiTZslPMNJiRldfKwvosdPbZsdnfUvupEaIfdm/v/MmLFMJ8//63Anz1i8L/jME
lEPlwXsRM6VrQu66A0sBzqGZZ7PvNsZ3qUwjUG19x4K5saU4CLe8JuFiI5G1ltRc
3CPN8vttQaUGs6gzz1+fELeSmQ+NXyUIfTON0ZNzKxHU0ST6kLAf0DpmKAgMmlFQ
3gzzPBY9KIfZcDytthuWRz1whJA7eo3vtitmSEMMYQas15ZOg141sszNfBHQZQP4
89gMUOPc3rvJAK1T4p6mw9DWdCP3Q8CdxGqPGGFuxgOTBtF4Ww0VsklvG9+tFI/u
spDY6I5q60Ead1qmv/mBn+CRMoiiY/t3jnoTplwvmv6EPPyXWTi8Q6lIaZA8p1FO
SVtoKqTCOJevSTpH3e/pDt98z4gNglc2jFVxBnY88zWog5lvZC/HIgYtshYEMSAT
O7ffXaLP5JnOYS5U9ru40PeaM0fixmTQGaRpM8haD7iizqtpOjf6XVpY0Zp0WeCs
00Ll13FVIS7teq4Ull/4IyDdpFSlxjgFSx4KRkefuwAg7eS+oC27R43SbjU0D3P4
JSA5DqhARVzQMCxVsc/mlJ1QSWLBqLqankOnOVhQvdGtFS6FevOo22P1gnKw4n2L
fttjbCds+5AuKHs37ru1tsjmXrY9iJKcKHVqT6c5jUb+MuXo0Ksb2XBieAhGNWzv
HXXSFPjLbW7xDLFg5qjdK4H4vEXiUR69mwSjvqaePR+LbDJzU8I4z6Qw+9y+8ZMg
BL5Z+9gceUvZwzwzwyMftJ5R4gjo1R0l3se9OEkThAYnzMjQK/KwC346EY60oj8G
g1QLIDTPjqw7WzT4iDWaQclzyGy9ANIJxOH/j1IfZim4NWCvblo4aULihFkqdXpC
D3jREZlYCrV54LsjWLsraTamXRjT5mtCjBAiiCRG3gtX8Uo4XOn+oGa5rlCFNaAA
aqaaYOCCTVs6qQ/xu+Q6Rrp2KNdfbuYz8JlKdx7vROulySwipl9MnUyS3dL8YGOz
+zzJMFEbU+Tzf1vQJngUC2SxYr5IoP+NiJt28t5frQehjMp26Un9IKz2lG3idgJy
jBFMR5Eb1nQYA0IOXJLaZWMNkpqnVu9jq3WHkd+B8bq53utkK8l37nepoPDJrQZb
wWmCesM5dXoOulgCbYLZs9aHBrWqpBnuf01XPHjiYKxKRq3rGhTWiafVYXDIIM5m
ypcK5gixRs+BLyZuV39eB/GD1w8zybHCAHV0JinhH2+sW3qUhQZNRNgzMv6ZLFIr
M0oOY6g/zHvwHGE5DjQ4IPmbMQIdyEF/1oGCwO9gDQMR0GV+KYwXip5ZGqNonjjT
ZlxZLAden6vUsUvI2o2SbR8sdwmLClgcVbAJrgqaOuzyQnwOpg2aqddWDg1TI3YH
EDSGy7W27VMVxgZGrgkexc/SQCFIgkS+lHuezyVzxSmTolFAMdU4MeYevC7deuQ0
PgPxJbeTbZ/2X+/54wtEnFB5DSaVm4Tnrmq04w9IoteHL2X2evqc5UDIbw0YF/kr
`protect END_PROTECTED
