`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hun1TMp1aaLkrjNaGwLpOzeNALf8VcdVM8/oU05oKs6f8DHII9aIaf4heStRkCyF
K4e8+TVMxROKR0RvUpKYO8TM10Nt4wGEHiSWM9IMXyGwxsf8DH2NHxoNgOESYWOh
RdoBi1hkp44jH3jbeM1L1rFYA0VLzrkfPgSPBdQ0AA4GkK4JKSZn4z9g52Scf0IY
uK0f+4RwAwyE7qZKipovI7IZrJ7EuC747b+jh6kcNYtGvU+9szlVh53AT48+u7VO
uUh98Inz9S8NOq1M4CYwfVWTd978SbXdc1xyHy9l2dX+8Lb0AXAZMKp6+lOZpFhm
Qi1RVDZ/vtauMxPMn+VAicysrVmR2fLAJSX+ORN83bdr2cSL84e0WX9wKmHEf7Gi
rj2sRpkeqAg1Dvo2gqmvYQTZRoVf+8AEJVllrXMWU+R+Sr8yJOOyTRxraKbP1ZJ5
jQt6CZjwwWZxymCipDUNFeWqbEyyt/oZ6Xn2VdoKykfg8J6xCyGIsoEuSvRhA/pY
AwG0m91nDW7p1Stbch3dxokOvkIWmjNnGYHJRRhbvDAOQMRYDBwspXHN+eX7goT/
ZUL8ClQOnZqtvlU0EZ6xlnYuBMwwGgM+Zi4p7fwQAy/cyaLRptjeQ6EW3I/MwxyC
ZpK5xG8xXiGG1cCEeJEuY1j0PFCyf98QDWH7Er/wrg/xmMCGrBZCDqQQy3lcgDYH
duBT1+Kc6FzAsQH7Eso/A8NfLEdMTxv5IsnRP4A2CosNIwmdahkQmoF5CkXkDAly
fa+RDziy7+fBZ4Sko8t3WDKe7dc9JHniNW1acvRhR/w+51vwrgmBZWrS3+VrAOG2
tSyT+UDMvhkD0tDZtQIzm1QVv66JZ4zDrQI4tYzD78CFP3Wb29WUFeLQqSow/3CB
Rtj8QvAmSd36xDkuLCTLOpmWCXGUCzeiufzjj2j5pOqonhIZWqZichKz8K0+Zp+j
zran3pnbM/WrrjYDtFzxa/G0eSSoooUBhjE5rtciOzqeqQKFpCzSvUdHWBd/wV2B
7PWK4/rWd/59lleQlM7i33SytkZ+XYXoIvfTiogjGlSxYuaeyXqCLTIqXS6cK59e
DwySM+SToDMy3NKKGE8C2hnKH1TnaCs2AtOxtOIpbUR2ZcDugj0duwm3gLaVLkle
sYHuTTF7g47Bc8HcZmgY0A==
`protect END_PROTECTED
