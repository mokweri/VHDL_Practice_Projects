`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qhb2MfoAw0IBWKv3ifC1gGRgPyBXIbi94y0qC2AuNlYG+K3czCHbxSW0ZPVBTo3P
XO5PpVg3+APGsi2Q6j8qMuUzlmoZAo9f4omWNoGXrgBj0wftKRIiyoZuBip2+grO
2g3cUuGL5biiA0q6CKmvAoamYN7WEHy/fDYqAb/lgf7cQXb36hLzTvOwS3+px7km
N+Ssf2PQP0L4bF7tYnYictbc8k56muHpG5qf7Djsao+t62/pOwuPTzaigla+FsQV
hwWZukK3dFToxs5+aqGAIkZJXHc0OxpRuWagDhikeI3qw9E1Glhs/ouHwWAupz6L
ZSt6bTubPZyQPiIGbC8lV8dbsGWf0dOgp29fLt6SAojvR9NootJoyD2uh+6zrR1E
7Xejq+yBrm/KQYDNFiTNcyrk6yM1ae5rl6nieX/kZFxy4zIH4DDmaWkycbLX5XIe
ETLc4waooynaYK0ICrbWFgAFzoqleRT+n/benddt/AtxZ6racL0kLU4u9xKbNPc/
F0ElaI0ZCQ4lgRw4Nh9mStBbqIDRrc8dTgYGAqPSSukMLBaTiORj6tt8XUYPIb6I
qe82h1Eej+XgVWO8+1P42A8EMniZHZYU0d7DQTo9ZYDHhOZOdwV2Tql81hZNXHAh
zfd5AWIOU9+RsM6Z2UFaW+1UhDN6gDamHaFeT1PaAN4VuZArFdf3aAHC/XG2PLji
YbZb2HtSem4UtKIphJ7luRrgwFQICJ6zA1E8m4LNXI5mq0hx37ofEfmG7FA6lfb6
wxrD4ku8SA0sN4PaaVzLTMRZPAuHbxUp1UJWkUb9OQMAbide0LnbaMC/fyT0rVjL
Hvvyy9hjLfK8ifkCqqxUti0tie3v2NM4YdxMMgTkKBCZQdhTXEZPlrzC2ndGF0M3
8qdohJ82vW+WfGc35F7LZKi3LKsPM547d6cheLUv4zJAFc7W7pSaGCpAeheBavGw
rE79RArYJq5DPJfDJ3z96gjS3FdCMa6FRmqHtTg+tvRciJcHJKn+Tek9Db/I99dM
FjP2kTF0Spe8FI48jR5/fYCyqYUkvxL9nfUHhg35iFB+B1zjYQY0okuoofKyd8Ga
lAZzbryAzx615j4E30/wlOf8weggO8SCMIJaoqBjLNx0Uy1bofeztrECoODOzXUA
rX1n8Re2zcLyPWYCEf+axNe/UzhVkYukTLbO0YVes6JEQ6wMvraKAiJ4ohBw/1ry
XVEBFtSG1Fi6mMrNCcKbI2Si19yMmEc+Z7r0Xk9ZDLmWtAyl77TzQCQ9c9BWMwZy
mTFHxn8yO0kr5EWojmyIbGipIlRHmGCbGJGubwX2bQhic/Pi6nzHal2zEf7CYm6c
BjoQP6cd5ji+mg10YHmvdUkCoQqLSYZEEWgNW3tJrr6zkR8X+QhfijybXS4rwdAw
5iY8XW/TUw1MtJi9TcHlkwK1U1r9rnNOF/UVyvTnP5Yf7uncmzzgtgSlQQ57/Ci3
PId4SSnOJhJZIvmXCAvPqcqoy/L+ubGY+JZztqewburMVB0308ael+/t0Ou/4B/j
2BrP+yV7HyIKzHCjbqnnBVuomJoZikJP5KUJRQjKIlvCdiQxbhBjl9ogj0y5cHlP
Jg5bq79Tenn+2CcPM9lddcCfkMZzYIiO0LPqQoPuqsCgO22J9DEUJk23DIUht9fx
pe6ljmhmWnMEuNP3oK2Brpxk8f4Hn/Sc1wXA32WVkDa2vv/xDdNDY2612o3JeKzi
5s5Jk2z7pBrZaf4d1A+nczTh7Nxln1wvD9xXM2eWbTlzGKMt6utibIsCqTT/B117
nmRsfY13mn/R1dhNiPUhaSjtTT6CF5OUSJtmCpsJu2HW4G4r2LXasMnbEgwFZUP7
uxpMX3QI8fNr9EXbZN3FYRfyRX3P5cumaNB8IxkfgtTDlnm5ldZfSfsZow4xlFDH
VA0Wk5Z4bJThRGx56wZiPPUpYGKHYvK1ZYnshXyXLoGGWNmRmBFGJxEBN0S8cqZj
jSC8LJSZ3h/WfsbMHdnHTZxFIupb84KOzgCfGoc53aGSKXJQma91Sj+9Se6VEGt3
WhuHUoLn3KEjHPFTxW2ojflouonM4EpO3aUPoFPyE8nBioUNxtWGlEK5cqa1VenI
Dqs/qhMnJcCmOBnM9liLkTDR3dUtyhg1ZAzbxQSLFCv6QAObfif1Is7UV6ZvdxOs
u8mw5eUsvGZqlfsvZhYhEg/cADHKArpd+fe/zn1/KTFslBsd45C0BB/hIK82pbtk
TVmixsbtA9F39RvB0G0JMny+7SlhvVmHK69jeIvugNRUJlFztUIizIWNDWSV7MMS
wY2/Z7/t+RokgIttuVm7pBgZAWLXwNPisWPC7NozTFT1lzB/qRB9IcjoxIHARNxN
NntR8dTdr+NqrZYtPqqeD2TEIL46lDVy62aR0HozItm5yTvzAFr4aQwwF4C+GgKm
hTshy2py8dSXnZkeacrqPFhz++o1gM1zgyixbN6UTJKmuuQ298Jwfnc/NPVVrsC1
W7Kc0wH65l+IlEgB9zcepdr+cHfGngDJw94Ugs4o5wKsCJ2FvjMJgDUBVGF+VQ9w
oK3a4mGLlkijYRVpbLkwyVjezLv393G/UTTTrJdc2wLhvjQPP8GEgGzmHnkvuLAR
y/bVc6jAeopuDROxPrT7CC358581HCoJR5mOZFMyhlMLsyr7TV7FvGkKuQG09Rwn
RZksDLHFc1XYSCy7EunExcSyNPQdvHTy+3DwwIDLgcw+vacvJoPWDSVkWtuV5nZs
/jBd2rlebEbGepx8dw3LoYOfw5wFKcXo9ZZdF0/ElfEuhShGJ8xCcOybqMeFRtdi
YWMKi9y6a+VQta8C3u7PhxTa0hqVo8CYLOeNYdwlv8FoWw/12cNg2Nf+BaE+DSxt
QfHdOuZZz00xwPalZq/YNRYiKqO7uAG2z0aPGBRBhjYd5+3QJ43u/enPO2de2Z+/
WZ2kB2xvlydXdIREbK9z9ySWyXjixcoYuZ4FbdBqZdHzvE7pjuXsBMmlWI78G4/G
4+lcLWtSh2OAxORryiUJd8Arz687GsfarhvSthB+4yjZcFg6/JnxLTk/K2gaf1zh
lnbgsZvNxvSHZXG4SAjDLdHxk1NzaLSAUfucZtisN2MZX8uWMPqe8qr7vUI1bzV/
chn7GchwzcGzjmH5BIZU/NnngexR4fCUB/8Bw2hw4DehX7Tk9JiAQx26dPKZGR1u
5ZBe91riDQmLs2AaHjAhNgVi2ZBxe2J/LQYDAxuW/hRT9o4n5g6U94Kf2TdWbwau
HKYd8cJpzOpl3bxANqcajeeS2BnayKt9RSzqPlxWSi0QFcRAAiNmtK0pAo9vKWDh
6WbodQhXPhqmdPneSSLMSc3Zobwz12Duwqf/GCdEt8Q+BOOdYWAGmHeoYHSlQKZ9
BL2JeDiKLy5YjyFUAeSNebH5wTCYJDcbW18JVICS1WNgbQNe4f7uRdBWj7zsv4vS
+3y94e+9eLQP2AZip3HpBjWQpcQ8Pm5cv1xOiE0f0Mx8HbSYozCRnCl2Y4pzTZM2
QTc7zUrIOmstvz76xFQlVrpQ3esPKYM8PqLT2RvvlMuCyfKankM6PR5Jo5gEgi7+
+mhLT4s/ZyDp0OE4Ma+7IFBx/r8/NB4cOVTO+QsV4UWHT3u1tDNBmszYUi1OHcdq
fBGvopnYRute6C6UENsAswSJtzcG1LmJFVpSf44NlOB/EzpIshKAQSm3+heK3U1D
4JEmgPl03tuWlfndPtUQKgnhfe2mLirwJICMaGvOP+Tji0Yam/m5Hcu+GFZk+EiD
+xDDwtpabGISWVuDl37qOsyS/gmmNgfJQ27DVYg6X5//Gvk636rRmAArGfHZaUAd
I1eDk59tDfVgLEUneXFiyQ9fhYMB6IrUkVGgQTnBNm40RB8A8STzrPbObXd+YcWR
hLDZiv3Lw89lZWko1+rlsDFmou3Vp4DP1/Ojpyhi/5VwRXw8NXS/JDZoh3CBPw56
uc+Dk8a0MI9FLDShQkMz646XVLN+kiDeBmd33VZKxmoNvvmYL7Lp14EeQ/+l6e8d
NoZWh4bBJgF5ow056ZRtbrM8wiK5VXfNgJNmEyC8R/rnQKBBmZWApdsyKh0ZhNbq
3XNIrRLDTyPvNg8aoPBB1rJYQh/CrEXrcWC59ARRMyZ9Q+dbGQOQuvK5rbHM5q2x
/zx/fqzMJ5hthAi8ww5y3D8IWUklIOWmJaWb+knz5YA/IhKNezViG45ZfdlpMOii
BtJnAomPmzbA969pFwOSRE8/21aMVOjN1fFJjOcc22RSiqjpG/qCjGrNFnkHfjVV
Pnt3V6UZI5cpCd2chq3/Dni0CGHy65BrOWF63soL55s8THcYG9OlRNzrL91cqdq2
YPGQoEMYXCQ1gPifn20b6GQ6n7yABmBOuBwb3lV+NsrbPNY6X+tJOW61cWOMUZoy
Hcaqh0q5i4daENApDu5/vHrlX4J+YLPJ7pJdx/vDiPmy65tfEfjmBq/KXprp57eo
4qFBDRMMNOkXCmrYFOIK9kYg74zCKp/0fRVfmGJVjdMg6MwmKHdvA3eErH42LViN
yEc3dVDTExme5cQuAsfOpHGoU1cDFLTwdpbf1TS+0iofyVDHNMDaGxCdfJkSm2Ei
g3k7iNBgtg+DNAlfCgAcB/0rUzFPm1BopvXeYft2caR7kZVy5eliv/3Pt2zGUZU6
6tFu2PjezYtnlv6W9s/pzQUgz8/CgGj1H0V0khPoh3oJ4gk5mtJq98eFC32R9cxT
jjjChU+ZSz36jEjIPnqyQrbwBpKrGaNHcxVk0wsM3afF93kWMaPctw/DxgGS8BW9
jEYy4O8O8zXIyGLJLYtxZVHkWfRi0uu0saoPAiLSDBvVI6UZCgjd1/AP5WK0f/d1
7ekNo9VF6R+llhhVRT5lNVrWvnlp9LoDqdrPk0lo0CTC4AmAmlprV+x0bwakZMT9
ddHDGWiJZ8M+0wX00uaa8JBqt91/O8NKZJ4T4OnHf9u8tfvThAkut1jwP4ZGqDcN
35ZnQ4piJ1XjsUoRotn5N5EzdYDwNJDLyw2vyIuQftRO3cQx8tuKzUhpn/hNksHN
BPqdfIpMWZCh0H56Er8G0NqfeXxrbwGRp2hgSTf2Fjt2FyzwD2Bp4sbkqcDLjvGW
mQZ/GvrUIMwh+lcsE/5EeMchx3yGuNwguYZ2Zqkzj+Y/bGc7WKDO1Hc9ZcLVxtON
vtfH97IxmvmQ717kpn5ZHSqzvIFqa+FKnUEs9t0zX6po7Gmc9uuWwuVv2vYPjo05
QXRxhj1nPnPBkR/oB1QXv5q/GYIS/fsr2MMfowalAiV2oQyL1Ugdp7Ll4S/waSqW
dtFKYafgLD0QQil81UqIOdikggCprfDHCq+Shw73YrEt7dP/kTXXQx0Q2uW98hsd
0en5HW8Pil0T8FgFTdZSEgONCuh+q+78rrh7vf72QDbf8IxP1eq06muBtfSpIrLj
jqskKve3Dn/aeb6MlElkyLuIYx1OQOQJiO/jr55/IlQKcUphOpA7RBZpxDq1ktDy
scqOOA0Sh3D/VUZnZF5wWmi2zH0WHNzPecdaBwK1il/obrgu0ErBjLbpcglofZ2v
FQseNsuJZlJi8opzGh/n7O5VXLId/W2we3EBVkOsUMqp10eaF6ZadLMubePdZz7S
n3JMOV5o5Vj8Iqt+AAiwFPGE+2S6va8X2HKpdjNMTB8PYHdIgQo2H+Ks5fBsppGE
zauILesHBkHOrOBLg6ghKTKJn9dxqs5Kc4OAp0XAdhzUa2mUo6ebyK98RRQBF2HC
ndHRdkUA3Lhxni3ttKlQWo2lyNRYw3jfB4h69bakUby+EE1huITIHOMy4fqDaeFJ
syo2sK0MPESW9bD4qlft+IoQ9nbi7D4O4SElGGr1WWq25P2AEcKLtcyKgAglUTt6
a5/kZnJWmN0ceGFJ7AZ9dr9DHnf2g4FJIJL8Z7JmPpqu/hXUU261naTcCJACffMx
2QPNaBRDkUZZ39LQRgBdDReorrbRaHXyN2x9imqlh0VXbhzfAK6ZpguzqDEy+KN1
uiEBsLrjc8imODoLAL82CCu5DeTJpbKIh8+xgdjQns6rrBM7bjvVks+FjfPOVA1U
oDte3B98YqYOwATuwAm0pcFJmGy/6e4AXTndxbV+VDsudvdaSGDidgqz6wv72Zry
47PHvrcMfS1fbqnbYbOSXyhbieVBBScvF/dnzaeDnMIb6iPfz0Y2KKN3qnm9cumv
VxHorbowMZqTGvKP5XEOdkSfleGg8yL3zhF6akEAnc0iJIG+RtVTxvtqNw2ku9GF
KHpvna01eaPy0MKQnJjGdPFFs5SJb40ZEGDsOC2LJdXmr+wEznB4S41enzNt0egp
FVN1oAL3fZirvte153S9UA==
`protect END_PROTECTED
