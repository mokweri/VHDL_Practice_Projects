`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyEZjEHX9lrhdLgxXwSeev0sX4EdVbby6VvedNLYz5KAH9oorU5uwXcDYA9U+3Ri
xTSVQwXCqkfEZ2IaxU29KYpYluTVihCmJrLLEQsuihCl3D+zdB+bT3+e1w+W0z3F
betLmPYm64YG+PbZmdCCgDrqDsPwORPDGawLfYKP4rRejONTKljubC/wJw5f1Kvh
fb/kgHlYmmqC5MJd0dRxcgWS9WsK5UAd/epg/P5kOKV3Da1RhTIQUFPmYF/82DEM
iCIaOv8Sd0FRk7Iap5zpLq2T0TrM96yRcGbS1tkGOOmvNOIQ8MElOcGA8Foa1usq
Cg8z84ixWQBOWWXjk4HCLQBff5oR9glKODwXsxLrp8oVX4zQrR3wOQtZI84B2MwP
D/h2j9ZKekh1ehhKgL9SytKmG+hWuYbko0tP59lr+ZFh7idQo8TSC1TAr7fAEc2N
ImecrYJrSvu17gvVJNhFEOyYuubOwIpXLzPdAvoj5ZmD9dAErj9dh20ggOlyEBEp
Sg3Sfv1Jnt4Gm5wc/1ljieOeYSeFofPrc+NTU2z+yLmflkR/8jZUoXtVQMlrmAVp
z5Iqc7dtKdIY+E4vT2X2oilgmfmRp6E66yQvNqGdS4RA6QZ4WCeVTzAnWRrKRQ6h
BQsf+CUYFF7ionQ856g0+/aHdjejGeOv7ObWLtQIGXqx1Vp42G9zmH+bGlBfAJ4Q
gbB7zcQE3AmhbTAMJc2JRcheCuNDUqQR0hipH6Gg2XVcHwSx/ux06+Bqa8VXlrN4
gQgt8P59qHJd5DArIBAxHzAnWpjel+NFKU+DuNwsF2OKDygTUVBpBCvg5EFNMDDG
zPCw8Zb0MxkWZbaZQBmcJnO6eZh1I8c09eHrt4zGKL/gMqn2+PrFHFfEpsDI+zj8
LG1X1pJWKM5yqrbeXs9uLqLmHBA9ShTZ1atCbL0mxrE279h1BlQWcT9A79Or39Sw
3im5BB/ABfE+2bTTKJk/VZ+hMpi4KoCk15hmCjQUV790dOgaQ1asNVhiXjZtGVmT
INf8mZVka/+heSBXxIO9hhGVSVKbxwL4QFTRiEGmaPhpP5sdYUYQTHFMgn6oP7FN
NZerwwwfN+mYZAcLN+TxLPlxSdV+Kvl2u9z9fjE/ldUA+OYcegQH6hzeeJDYRsUA
EN3pFFgZpA4/v08amCGzLt9x15GqATwG8fqK2noxlMl+n7cGyqLz0Td7v3dRSjeK
6aPOiH3JUV17lnLCJ2hLaFCWOq+aJ8zp6K9Gib+Gr1/o6gObvSpSeUmlvEGfdvwm
TGim2nWmjvS1v6HBYmT6wcLipiq+UIYMHgDUN8V/Hcslpdn1NPzMhwYbsNe0YD8/
OLufChmZyxp/QSmtwQ1NOLlpy7GUoLGJQ9CmgnHGVkg1ARSKeuMFveqj+iDXgOal
Ag/acoqm9wOO7vEwhpokeCl9sFKWu0b42AynHU2ewQJEwWDOXu2QxNlhK6/b6VNz
HQkRITtLvKvJ2umxD3gg8yrOhdGPj2WOw3fULk9YA/KESn6ix2vBKqBo1NlLqlsH
Y0LhMy4ZVm1ToGDSJ7YBoPvxODhevwxQkFYPerv7W0kzsv2qgs20cICw9cKgBsyW
jGBRuusFVqZI/xgyVcXZv12RMiJ3FStg0L+NZ2lHlRUF3o0CThLuPzP+VMw1p79l
3F0heJ1kF/AT3I7bWb+p+3hBUlTovuseifc01EHWPuShizP0aIIWJ4OwUYGw0cwD
EArEMz7X12QR9Q4hJwpWeFSweUSE4M/VNDyP8qAn+VTaKIeNk3ZSBE/f07MkN11y
HFsKJ5cqy/UaQhK0lAeFBJZooodJYtNqu5DiXAOpyfbdYGZsuZRZN1A31DWD4lzm
4N1Adr/rARZxwdt4p67+932QDy9FsQdhuRKElNNC1DU/JQrNAMCFloL9BjOGbj74
CYbulYzGDCm9l6BeIlPtyR8izUOX0fYFh15fYSweX3r2qGDDf3CwKKkg4n5DCqBg
ewR8onOVUVZGUAfM9VihPw23QovE810wHQOH81TPHSFTbXIpa/Ny8wnhQIBNVbMm
xd9XjCW7kUUaP7127q0iu46YzM8E8YK/NEfk8T8+JuUfVTzNRgV3ZIHoZuvM8/B4
xdTMc0C8D3gEyiSNACj7ZOHZLJMrbSR+D+B21VRdC396sVo7Ccj+espmSrU58PGu
mX1kRvIloUZwGvJkZ2JDp+3K5KoOhTpI6rXwMFHTWosdDAvLuaB9vJsYcP675xeA
FgfaE03DhXcIzwg8yEiyUA71HNITWqa/aaTM77giftMlR34H045kDNHrptzTllus
SRfCqdeq+ev0+MBiKTIYpCnqi+CS0XrxtgLX1TyrWldkMPPR/wFNufZZsYdi4VTr
TjOxsPO9WZw44TK40p4tCH51hnAr/mL/msec90jBUPaxIjee+cZ8UDfTSrtW0NkT
+5gW2Nm40JwSnHHEm3ES0m12WgfHBHap/NotemSjzPd7S58orNtyIMv260zsQ3/y
Uo8+s7V9DMzTVGgK2yCYsqI/zUBPN7MqRNa63hX5ZntKJtcCQ+FyURjV/ukuJtwC
nm04Qhja4gTeq9r5BaVCcEmmcpu3164cDCyD8Oj/2N1kv/2Y/iWoI8uKQVtMoEqN
dpZAt2vlI1EiCKcIN9ZvlOdwtkpMTVv0RgJ1fMV9suFuG46wsTaQiN/d3900bYWD
Za0VpUb2ffT4rodBNwWro8tacFZaG9O0/AdbZ3rZjsx08kTauXlhClv/lHcwmCnY
QRDywzNTp+QMf5lu6rhfe8DGm7fUNyBzRie+/rsTw5LqZwgtYp9hrto0iTUzxELh
DLo3IeVp1VNA31cD1In9p62ENPcT8ZiJ3nZ8ogR9psjloWmpwDzfbFecSDKJ4JMj
s0BVaSg7AlDnLasg1vIY+uD0/n3Y2FPO2WzE27ZUqi8Any5jelYWgy9TNA8+BUgQ
MOys9wGZ2X04LLQ8/qi3ysYeEdW2HaVZjR7BOmUqO8LEQ8b93hCrjNn19rNHQLVr
YWuLIiRBqHz8els40rcAntt6wtZrZjXxjBCBVZnxHGPxjWoY/k6Kh4c4QyNn4/Xl
9BjGvqUf8EuTAfZYSv2iR17uEucP3fv0Ni/CXvtP6m4D0nNhB981BaF+/+RnbOkZ
LEtVk55iDtl/lHnjtJaYuu6vQYl/LOpFbqO+tFEVdQVbzfs2OU5/T6yLpp38SbjE
H+oBS7MTRpRX91x/NQXt2k7mLUbBbJ3lLEGMy7vwL1YOaJzGhZCWAr0j2/wsMtxv
VHxhsjq8oQayO1YeTQaGOI5GwcZ1VlFmYuJMebn0S+9rfKTWJAVfsu725E1GdsWt
UmFUYHZ+b8NiPyL+XtXENR64Gaz34NngBoO3hn84qUiQo6PxM/i6O/5HsYRrVPlg
E1Q0rXPuCIb794Rpv4ZXu7j8GOXmFqrxyt2arTjnjBf4K0bAWgSNKoOXNYa/uBg1
SXX/Dm6IjeKSbOlhNruWS9oVyatZfVTgG9JCS+5ohenRUjYWlUtJF5derMx6pi3K
JPDs3uITe+hfO1l/OQbt00pJU8keA8Tmz9/UJ7h0C9Y+7ErUix3tCAa1rj0oaseV
WCqdL113z548mRHvTN8QnPf/SvJdxIirIg7jXSTGP9vfJIFZ3A82FUY9YGw91E6J
9mt6w8ug429BBClspobKSVGmKpV7VzXmOidRasp/AaMP3NlvebeUfudu3SGqk6tR
D1jkl17aBQX4kXVSKyatAznUitAx9wBlij1CqOzSGUPExubMJOpDHWhGz0hwLsMh
luxC8P5f7/GQ5KDd/Tjj2NX09WnX6maQxh39GjirxSEK8vDaGVOjrlf74xGL9Y2Z
yFAPF6M+hbLVE8IERkmlekd6Bn/FDAvcRjG71uGONXcS9lyYbhG9YrFcq//u9rhf
+Nm3h4gcMA9KzK1H9chu+wPz1aWAUtQzM8g0Q93e5zcVSkq2fewdyviBHRRgvduq
XZhZA2iJ1EM80BaFW/j/W5fcieiAVxWTZ9MakmH9oj8b1MCSSDurXNtLKG/Iywwy
WAbQOrcrCjT/edBobBN3SRZWIGjGdc+neQu0u1+ICk56rxJ41phEymcjgITJrSZ5
hznyO9qK65NmO8MVK1M2QOH2aYX1BS3/KBn0UnFh44JUNCUR51aLlxjQJV73iLiE
lVABpOQGCsEn1vZkoeajJWSNq0AsG5vvoeskbZ36uqYmsh6qn1EnYpW1cx1N3l8R
9kZ8WGsdKSpuy1qOuqzeMkB6F9qUx/0rIVUk3C87qYjutTfYSyTdxJZregH/8OV6
TGOgMl8c5+lMRGimHkdjjw5ySsaO/ZynfyNzQH6C/ZIiKUWr32NAPgTZlRPlDLMR
SFQd12tRKIzK89nxk3vJHVJHRbMZCeRwNqujDUKLUtCnlWqA5ricm5dlUIIKcO9y
UO/ZH7Pid68Q3Ljv+p9KlnzQ+Fw6NTQeEnbF6LCdfCwscp6ua0F8Zz24SAuDjDuJ
F4U/v3LE/LRTl06I8qtc/QFwqpIGGcS2tsLEAYM/D7cGVq/ukcPgTcQTAH0Ly+fd
EKyFLNAuS16cZIBXz9r3KONns1x6WRIglq9WAZnFJEeHEz8Nnn/foUjJooP8bpgR
Ndz63qF7L0xeLCY+cC7TcVTRw91l4aszc20OJ8IIg6NqfitFcAAjZoGpaTWr8iX0
sty34ItuPIuj7wVvRUw1Q0ATIfe4QgI24SeXtMSwHCOCLWgY3UEao1Mr02mz/8qT
X78mDH8IN6TSvBqdNsXF+wZHeuPGMkfnQ5yHHwP3HTyADYH3o6HA+uNckhAynpYo
Yttst9RtStnHn+yQJWDd+3nKaQKD0x1eRC4Djxdx3Zn/9vsm3KXECbiepiS36FZA
+4n6QwjH8wxwL8BNwX1aEbOdZjPjXdRIESlJ/CnK8z+U69fVJa3+4LVBV/iNtUGs
rdWdeIz3c16r91XYN+LykrNE+n8EAcCcYv5YKG4rwRJ8hXO05aLp9Tndjgsb9VKK
e+FA4/NZ9cou9LIjJbse7B9GGts3KWSt3LWGGlVC7kbRlXYPUmU31cDyC30ueqcX
NPbwBCn4YKuyIGW2pnV9AZ/P7y05ZxVVzdIJz6mJNEYaB2RA3JrDtyuEaqqWtErl
DOZ9wQsabcN1aAKO7aDnh6D3MFYH1K91wDVVwQEEFUQzYtoG8SM2GzDpfmftCsI7
FWJL9+CHWDLhd/7kQ/0Ne3mtNpdt0n8Hd2NhXMTSGK5p6KA3loYZJRLJGVXTd67m
BZSvyONO5V5sGIoktR2+n4MV9VdbRNjOzgO4aQ8zlUFku6z8A/eHILGQLt+0b1cC
KKxX2TSSgHmEyDgWuoYztKfHiSlDdh1uhPXJaB2YN9RWLw0v0jxm1vradsLBt3kI
b0KynJV1M7kf4MoMhJzDfDcuz/5aX8beDrj+opyVt+pTc0Kx8JgHVIPGVYYDRx2Q
/u91drrOKc+zWfLLqK2uPdE9wup1MO6BzuQ8YPcEiJ4WjCSWNGA5IHQTy1XgD2vV
HS6fLYWWwf5II2Gwzo0Admg0NFKP9jpZRu/VE9WG1FGRMM+zK9EalQD06wn1ChU9
Fg272yTuBHxfO1SEh8nk+AXNmmDbO5of2iF+atnKpIzGvLpL3cF0mmAf75Cn2ExO
dSuWjRzUOkTggtEA+RZoaGhjwOnONl7aF0v2+f8BwmvIdhsHrU9QaQp2hLKmbRN7
Uds9kaNHbVi/83YuGgz7nJ3eHtytlUNm4uQorV/3PUGW74pvtN6IY2ZyULRjMLDR
RW5dNm87ByAvjVbisCC3xkRvmFFNkyK8j7hHUwVeR9R8CAWllW9eQeZOjnXJoOTh
4rPgcZ95whtPoX5USMRHU3xgcBNnofYwToY4RVIDG3RUsY/4VZSsL/kIJs+RkSF4
nnN9yOa07NFn8aKUQZ4zVf6P6mabw+W1qKWK26oc/IY1flwxq5Yuq88swSm6R4B+
CtOaIA9gryA6D2SlEcQo3FtLbs0IYoi3051jFJCWd50cdfuh1O/vwR3SbDcaND9W
0C70P5Twh4eoJYGLXINx4OnxBJbCW+7weLZx3if43CwlUgaLzZ1rbqv8QLPkOPLc
/xYcTjBmXATn6EfpeHgIrjpHFWaSnhoRZYV6FKXU4IaQlQ02VovfG36EpPjUagjR
o585UmLVN1uLz1TVqWQ8hPjBu2emomjfV8xKJsuC412ZzoVQ1Uda7MO7o3JdKGdQ
aLKLkyndh/wuWr784Zb6mAO/BwbiKkFsa/ZFdSuMFKsFsioIlzypHoCevhqd/Wn6
GwJT7eqb82c5NWASo75vMzOI+DheQAM7ScAHxBs+phiPkSgHoagIVMbwQbFw3fkR
WclCoH5I063GEn9p4WGhy+fvB5fz9jHgtrz+rnDvxfkKIkrR7C8zpI6an0LPTa+o
PgFb+RH35LDjBSxYOnw/nLeVz2+g0nQhNqqNn3DU/xRIl/IHnUAiMB4V6DMP87wS
GhhRr3n4ITZoVys+wmUY+R8hysI4fTkSetlx8gnh1AifmaCfVzzsb2LP8qjJ/5IJ
vzeyRYtLRsLMoV/apvb+Fe1hWcUAlh86nHP4Ou78xkG6yec3/gsI9VgDLp82z3O+
TnGpLhtp6OPTCffhcMEv+XRodrArt5r1Qeb9teXYXYcPfLsCiqABhtunU4iaa4Xv
hMeqva1Ergv94hdMCtFYbJLIzUavxPB2ok5ABKu6YbLd1fY2EiXZeIzPK7JJRVWq
/AZQkxhTYh3bxz+lJHMFP6dRi7oZPPIb5fNGxzesYLLbEUkB2c7v4ApIWJrTdjZy
k8QWy3sN64AJeja+6whtDxb8Uc3N1YEZZiM9d6S6PIamgJhK3IsJMgsk3CR6NzG3
JPjiywIPwuY8N366qOXaX8kNNpw5jQzuQ6hV5yIxzGzEePHYA9e7CaN1XtBnQM79
Ay0oMgOT+xdMfElLedB1eTe/6VCVfVhVydYidIcqRmu8OrQOmJ9b7noKumMneHHQ
3b5bMPyhFLZsEOi82LlfEqGsQ9+iD6VxQJrPGdOXwCKL2hPvzUG0BN7vbjZYMVUY
jqPY3hbjxiogAUIaoHCReiIpwUSzR0awFxEGum2ivIXWwEZdMvZRX3Of+1Ed9GD9
tnkVS4Y2A1xlMPbI6i+hhEB7UhWWTveD9eaHkF0qNam0HD5A3BCKTz0I7xAtgTdW
Yrzr5G/pVMMaHte6LgN0QzHWPzNUgrP+5O7AH+VAYCkGv3UwDQWVIO3RGlScWLIR
9KhL41eh+vzOdP2nXAQBbvCRM/erA2bhY7afDgsP09aBIva8Kc16F/jJ4PYQ3ZzH
lZCxlLSRqzg+8lwZdwiRC0/Qe3ucrm3zA2rbIeZGmfQykoNx3BwJEs5gZzW60UfY
+1Ne5w/i4gOdNKL1+OJR6VlvKgvEvTocBJICSt/CYkmjTIOedomXFGG95WO5oRbS
HRL/WmYBakgLiUe/3jk3wy3otFVFqD3EZugFQkQCSvvPlClVxaJBcT0XsDr3g46K
Zz+VP+CGAjovv/N4DLrjfcjeEQk92g+p/vDbjvzng1kartiR9dphKPYdSnU0kNcE
41+Xt3lKH6ORa7FU7YNGY8VvWPk4qXeoDk6vnH8JCN22atW82ajkrMB6qjeiBjmz
bfVvawH1rNeaSFj2NkXsqbwlugGxb+2ZOlz2/Iag72rvvGjsCCQghcpkanc2VAWq
RiMig996aZY7qYCEwhIP5vAu3M7hcqWcwLd8CzgvfC5alBJGEa5tneMWuOBl4T3j
zXsaVk5zcnalIchzXyYj9TaRl8o5lSPgaYYvMDDyFHaEeG4ZCxZwSQYIP9lPhUxP
f3VKT3+EX8ubZEZs94BxP/mJxmVQOq/cRj+mqrIU4qLJUpBaWkyQub+m1GCfdKtJ
cctjzReA1x/V5mudTxQj1F7mZuVjIS5APDDvBZjv9RhvidRrvVEdk0WNnfgY3Jpw
PhAWV9souNE67XMph0o4N81CFlZTSF/q96S9uq/CkH2y3z3hSEg60fVylW0dpCKT
DxJGB/m7gijZWRh2ZALkJyeqcTHrEzs8PULvs6SU+sRnSpBA6Iil72X5eX4UKcDj
y7haxF9xTpMJqslQb7A2gnaKlRXKgfcc+RtP0wDCO+VKCg7STAsyf1cnHYSKxDqV
zqrgIWEsGacxzkuqHk228b4Zvj0e8cHlrG1b2Nxi4PXvya9UReRLdQxsLIYhWgZU
i5KbYR20zlrll0luvsckuD8pEdXpYgOG+bqncdIjXYJSPKVTWV8JIZvviiXcr+/t
9H2W4a35YLpr+IZA1reYoDvP9OOJ7AIUVzOq3MAlt62gEItkAW+2oigtPXZbeFqF
zgLzbe9BAkDmCcENBN6ouvEr18J4JrUNq9eyFjqdreyx3xzgZCgTjrhmAxkSdiXJ
t3MZSealShfmLYX0Jh5EWw31xpb7c9BM4DAGuKF9a4RDw/ZbLjzfd5tXLiwJR9PM
TWA3ZQVNbgrQSxxXOXEEngxzDW41FJPV/M0kW3JQL1a3XlihF1cH0yDk/OJQhrr4
hh5bXOiT9PWVlfi55eaZG7hw6hDSaPZBlzJdli/dq0/i/O7DC24juNRrDL9dDzFK
pQbW665cF/aumR+b3BPkNIkZ/QxqV64qnlikrPXhAk+I2zQKBx2edq6fVT3NgwX8
2jacmkZmYl/Jcbfj1iKJ0DGtf5m7+2QzCJewCaBOnF+HRft2ye467dE23/k4XcIm
yTEePhXGDxrINgFKjOc0IZqjDR8gEXmE2V1+KWH1ZrQAYlOpS/XO5DYOXuYD4zyp
v2FEZ1HAqPMCrqyq4eF5BgCeErcRcoW/Q7Gc9yX6uqoPRXAkyY+Zd0CGJrE1ZcFT
VOzUBF0+hEmd+eGCV/Hlcu1pMEEWCZICPzbJQL5rWPShEaQTyXqaH6prCNPod9lh
z8nUusyKrI82myEVnrJttwW2txlwFpiAv1YVXWom+rBDnJQFm/ynKcQx8mUdqFGx
nyFkjIylMjI0fR0NWh8DmBwVPe8Duq/bUWsuZk4oBZaE6hUo+BGY4e7Oiz6fZmUy
A8UvEMuzXsXB8/P0AUuFkC+nbSe6m8awXJyv97z/rzCAUXeXgq7ud1VGf5bIBFed
UacTcUXs9pdQTI7k3i1ua1krGVjWAXgCZ03tvaqhDDjSL99OkHYxdwn5bVW8CLzg
aItfHzNASQw+cw3uI1+u+duBy03AdI76GB1GunnhBV+h6fLyF+k4GpA5VgswxwrG
+aAbZU0fxm1sfjVxb9zALc+a3AWl/598mHDWidy1lR3G5pXJ1WHDoTjoIJOd/2Gl
fCS4ZxC7cCWQmGiLinhrf7C3COn6unueJ8YPNcusr+4fBxiT3Nl65l6B+oDS4Qjq
o5/1c+VvAxsJAVW+P0JX5KwIhEkzoM33jHqrQyBMdK8Kon0elzHixCKkKmLXyqEY
4S8KlxLH+0/hY3q/hux/2+7oyaTl5RmpbgtgWtcMaSGe6gwiynGPPDS2XuLxNcb8
U5kJFbGws10qWyYqqrW32hrdHiGTlTpmqcTfepsi5U2/LmTexSGZatdWwTxwO9Z7
+v5jLFVVL9Q1J13rK5XA3qwSt9bAkHblXjsHsM5V5Mo2/HdwJ3qdDyJ0UEWkFpeT
CIgPu5pD/isKVhV1GiR/3Y9dlrj8WZd0Wi98dHJyOPGv3oWy3UkwD/h3zFEGzJ+Z
3pRZUxikJlnnIPdQuX7z8iiANDVxGNEb6PST88JMn96j+qKdjwPt+HKtYvypj/qe
0NZcm39ikc48RO/KHyGYneffYIi+NvCbDJpB+u4pznjdr0LUwvUH1nianPatVxF7
E7kxHq4Re1P2zA+zYDSG9RHoCbeBWQytAkWTC5G3G8rA9tEKXR7uxJ+hS8G6aqCV
9bKkjZg28dx394pkcuLzCmfLvDYHQKS841FXnE9nSuEPAHu5FidH3jWgoaeI88eC
JnBrwaj6gMC+TkXfNKlOUdU6TNjsUaPs34Th29SuCPkJf9Gz+zWMlTTZ5zBz06yY
rJa3vThLjHVk+dYh7ejtjAZnNVyeCFzBCejry+nwZ4snWTGEWOrfTc3BhtXDSETs
WLQdc1uxX0hrFKdOVP4fpnS+nqjwvO9Bg57IATR7DpL/Dohb/241rKS45x1uLO/s
GTbjX9JMGEsEwYqBlP10Cw5A/NtBY3ihJEPpN/Fb/fLCe7VnnEJJ2JYyfJIY2MRM
UFXT0ERYoDLau6eCaUr0R4jnxM70MxvRTQhidFZaPZVuBelmI2oBn6W+yOHT9Jnr
hAmub0i4NuEEwkckulhUAvJLgxD1+uUGfQ8ahX+F7A25DIp7UJgIkf+RgRKyougb
dPgEPSMdM8z9IBHSOGvslGsM6EZFPmYK00K4SBwtuvNCgZB04z0T5yOA2CAl4rfE
5xRTFfxXVdRmmgP4u0yqdEarDBu/uUstfGX/CdHFHt7Hv3/M3d9M3meRRk3/X9x2
l7iTTEXTUyBpykwmEFJ6Q1tv+5Bqt2HuE7tcWQ1SvKEuawfVcDDD9O5tFvPpAeDE
BmYb9IHHUwp67oKRvvf+oyjB1SjzktVFL44r4yfXm+XQim+ZAVlV5Ddkki/JIm1m
u8WTUY35FJnSOzc2UIfl3T36ZupSRjF1IaW3lZ+ZQ30D99fIIw65O4N2Nae4uM2T
VFyxKPIDW7D97q+1AfKDaKKXxGKv32FF5u2/ZahGKwbgJfB2Jv+05ObsarE8NZwP
Y3xW5N8ViKpFtJFJSaq4uguQut3BdLhu9aR5ZiCXbJXeZFZ2+O8gAdOMdfpJtr+H
Q9OJlbVp1vKdhyy9JHWkbIBSHhpa7k7Ys4JNA7w39h/nZ3nRgHjWllO0kK/Pv9bf
gdY0POd6ma+0Z7Egj2Bpk6dvFXmzLHdnJuIYqPkV2IRRg3IDt8+9k3nVRXSQTvJQ
xSD9iWXkiFuELG7/P1pOc4Y+4sXBiVpG6+YyWyvtjMGBkYKhuPguo6vaxsT5PFWL
+7keH4GAxw0u8jy+p+5sW/qFnRLv2skIFNAuVdafWQVQ9X9Fet+CA5XXM+tw29dP
pDSpobeV7I/dZufR+n3rTVxSIxwZ+b9iVTC1mIXlp71jHXIVz+mAQ1LnlTJ2zuZQ
Yo8QzqRpxbzA8fU0ocRy16rONw2yfeEHx+Z5CryRDuQS6WZ7a7WXswqgKnmmI6mr
qfrdaOkM1Vl5yfzk8lvcmYlAZtADeO461bIKm8ojeOBxINriBTvZj+UCzW42F8Ic
BO9gSygB84rvRHT0kHkqemAOYibrkVMTH5reFqwppqkPCF7Ajb23+GuwROqWjUJs
GpdypTA8mRdZf0Rn1Nj8yy6if5G7m3Au8E5Tv8Pro3shVsoXWKU/YTdRr+oI1EiG
DgQdqlyIThbCCU7sUx9pdSuSZPkC8porV5MFGBlQEDmJlDAORfX+vt92mcEdX4Y7
koxEb8YzmxiijgaMSYCbqMa77qXiTxRmPxz/DLRCjd+bH4gRBLMunjGrlkFe5xqT
id8lPlqCh2CYRvXgd15aOJ3531Hj+cg87zaH0mjK5lHIDfJeT+1rQSW1F0119hTp
ga9UOoU0Mq8I7nSwr7tFe0oBSmmGWZZU/lFGH/RSIaiVwluuLhAwUmX2hGWCmzU8
eCEZ//AnWF6wkkHWaAL2sTLyLignxpq9aBUzNbBGAFkr+k3nSlFOX5Vext7FMKLG
JZJHCzGfekIKxkncf6m09S8LdQODX6O2zeIyB0ZqLDf3oChK7HHGA/p2y8a5YYiH
PcCQzaS8zghDt15i8bVECZ9ubi3zRiam39J10ZibaCN+QDkY7xpHKcdTsL3/a1fF
BTBKxPC2o7IMpUoGyPXTzDykjk/almb2v5jC1D2aLjh0Y/lu5B9DolgFo28mj9h+
aY14y7CJFdpylE0WrViJvnGbk+l8eAAECooVmdR6++HKhTtutKYP259/BdxBBkQP
9LJUUZYG9dQhBc5U4uKe0f2eoa9MsJT0HcrArLlXfar1miFz+kr/fJt5XmMX9oXy
aR7zLlZNpbOMcPk+yl4L2ygIfJxK7w3Rm4CCEeyk9i8Tlt01xXGZKACp0f4/bX5i
VWOafgI5lo1hVr+TgLUQtiwXNKLqs1XrTd1F7N28P6Beunp7JboLy+RAvuMaL1Jr
yP+50oc2RY1OzXrnMc2//C9EJ+6cpvOHLFHgveFmdWdruaM3phsDJndw6RguMzrY
yVOHlGNDcaxA4rq4cNgis+GYpgbJ+eYMrBI2AxNyV2yJ1yi2nbHMaAoC/oFtQCYE
JcYg9Aq2zUzZwkEAXhc1jrcKWkz0zmmk3y2gpu90EJ1UxgPgdriLUxbrPnRW32ST
/a+pyGxt71ZQJBlB/k2pPvVsQLZ2kFtgvOKUluhSFN44Tq6V7irRGtTkej18qES6
o4KjuvlG65rFNopklZKtS5mFHftXk9u5TeOqCWIdGFaoe1pjiUFYI/Vhhh+EAms1
8JWdaDRJgATt7fZd+xAUBdbKbJTerjZnI6esX3RcrTek9h2kitLTlDUbKT4HVCeU
eVLvMPrnwA+Th19dVrW56Xoo7ei03UHDCXylS1AnT25KXmbpUyMo1r1+eQdY59Lw
s5ERwTl+dPuvvxW7uuPbl9MKX5zHAIpGplcOomr+XsRnaf5Nc6wA5Efw5ucd66Gg
ZLw1GbM4OxpFnXzctr5q5UWvc1oiWLx4sp/C4tzpfR0AK25GpQIKeMprWURGaH6P
u1jYwCg/k42Ce9t6C45AMRwdj+ZFZoQuUVzJZp7Ac/P+u7h/eiDFgO/KjDMc2dIb
rx6HlF3TYzQKblrMcjyl7njOUfY6vPGYdNf4Spv30imAN7BpthYOY0gb95yFPUh+
HUjc1OsfiRZmF0ToEgfCayMLW364S0gEpLYqRDj6y2bZz84zrLm3FU1Z5KUmLM1E
RW3/IuFeOUGyguAQu5quaVi7a8tXViugvgejOSvsEmbCL/NAIoqhs0OYCgSxhrza
Fknk2ohc/UHAdaUAtzx+wlstA9fwCuKlCzbjBSoL3ZVFH0cg9W4oxdMMtOuNr2P0
tfOcGqkQYTfgiqakHDJHrbf2kgpma4uX9o3yGywrk1KJ4KEhFoxG5cTOwIjDxx1A
J5L/15cNKyXliWrlDjKYnI88VjsdZ+fpaUPbHJU5R1bHH0UEGRz+RN/n1YyEX+tA
+WPT0qONp3fIPPQEq7+eBcRDn2BYdX8XSxkp4qPkxG84uLbd6Dl+Y7J/KLlIsSLv
bURaFOzN2qFWpTXR+ipXY1Nqt6t9dD7M+9G9BDohW+tkgBR6RKDFwAd7CkFE0yLu
KCO4UEbFalOHvZAETIOrolzOszdoNmcian9pSQqXwsRMmRAdCGiDUtEP4/pKVPib
ZEIumjRDZrsEU3tzfT35yUZm33ZzHBdsRoiDLDR1zuKKNK7zRgebaIs4BD0EYSyV
B9fRfzw/wCXHbI6/VRqkjzTLskh3sVyoWTgG/wPLAs2VmTMNsVHoxhrAhLo0wl47
DdMMYPcQbQcun2PqhQFLlG7u3to7zMCxWvbe+kFJLHkL0wIPmIR2StmAdaoO3m5B
yRfMaXriKNWr4RremN3ynuYkyyhq4AW71CFIq42dm3unNwwVAP91YgfXzLlIwkMM
GmBZifeo4aFin5+6ik9066T/3uil811vG2o5LGvro4qc1CbufttuelX7Sb+LAbYo
ZA//qQkhmoDGVrvI62Pqt0kIZabg05hrYjRLz0t7uFdBcHRpcPLgPpzmKsfnXwC4
qgecdp0kiDN8dKP7jgCpd53+lNHgAe+y55iUlZvFV8srUZspwG/vRMTRrleuKtBp
/yUcVB658SSRU80+YEPcIdzXLw7aESv4KwzIeN0N2GuwXXoaE76P3YJdVScgXsmd
Lm3g0aTutfeFwZYldob4T+Mbzb4wGf90Mso7amK65md+XldfT+EP0RjlW0oaANYg
ObAD0pJ/CMvYWmDQp1h7BeH/Bv6yCZJxeJ2yaHbdRwClE5RaO6MRM8TSKLkiuWVl
pCUp2vZ0TWzR8gY1MHu+siGqM+8J0SpHvjoNwnTPwIeoWHrctnwIVqc/6sL37CVv
x0CH1tdB7J95nvrFuqQKEMCCch7YgASyCgr2o/6fKKN9g1hwIXoWQEhdxk4lMbiE
4NLYbRjhdSl9iz67dNDF0ZSszdDnvPhgLzk+nZ8fs6jInNQmrGJu7wz43ykuAa0s
9lvBeEoi8Z2mA5q1c8wIxahqncKDGDhsS2DVvERnPgPgba02vQGDOPQnoQ+zDCUb
4LGZn4vsXtVjsdBShfxmCvPpiYifd0hP/dnnURovjUypPqyq1xE6VpV1Gft4AziW
`protect END_PROTECTED
