`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dqBODdl1q6p2jXgdpajWEUGPNCZI4vInJSZXJNM/vdYbwo35eEil3eFaRkS6agGr
PwFBpcmzvtJJ1G5X0dGTCJtXx5OyG4gjIHvp2pNlRfLcC6sxkYYT0Fw14FAy2U+a
QSNmdk9u/6mMUYL8QvVzJQwYZuR4VG4p0gf1BTD1laa1h1+keyVCQ7DYIzMUi8eq
TeztSIZOmHBOTjhf9OEswcZ1mSRace8lNB05K01CNYAopyl7dECDUFxOvKtqjYAE
/5Vf+eger0WJFcliGjEVzVcsI57f9CONWTOTcKyrnlu+a/FM1paz/atnhaGdMhtf
m8+Vw2X18Q01S1U6unkXcLqQuKYNyymMfuCtqy8mfZ4o7f8fW6vOvyXo4FjNREqF
cFlNk8S1NVeLKCO54FVGpWdh1+MGtzuz4WoaaGYjPPr79ynxY5+kk1I+aUFkmH3/
dCXNM2hL8TpFUpeZO2RtC2YVc1UgybQ0P+TUbRmQQYKciyZMUgtYCjZwBm4DibLr
TfnuF7TWv1qmwKRCJK49MT+ayLXyo0YO7NDj+QI0dEPoUy0jmU2Pc3DfovI8gUfC
/Eh9zUv49mDt9okj/O8FRsBb6rREPJdvKJueZ5EhrI8HkTET64/oDJ8cgYpGu88K
hNnFnA3YiaiODxLmcqpbmeqMjSdzkXOznz33QWXTA0t6mzElVsD4OlnFWhmZRmN0
Zq0ZVmMSDL3EmSj8xw5vW56fBK+uHMGfWYhlafx3AzU=
`protect END_PROTECTED
