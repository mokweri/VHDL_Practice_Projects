`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nlzqmZSvsaDblYzTv75buHDrjRLanxvwT4iUFnAnGieK6Jf4FwQMypKyZQVH2iC
VS8CG/38CgwiLs8UmMMokAXsqzezGALNuxti19oLwtc1NpzrvhCathvcoYI1ZYRT
y+2Fe8ateexRcHdMQsyFrdxUGM4D3yMXqEECoVXAalbepc2lQjhQQHHeoqklmFBN
D1Gl5dJLGMTIe196It7mf4AxatRVOi5cSUx8ofEUyGxMGB5aR8+JInns0cR3exzq
6/nBg6KnvW93ct+Mt0KLpGhcqVXacEyHNxICYi9GKTL+0vFT4vPmosi69IBUAD0z
+EZMbS5GKfrj3szaEGzSOeLyZwORliS1XXsZy308z9jtQ1zdM00O+k7oQccDFQ8K
ORCaS1I9jO1ugaYjmQWXtV5uwXMbnYTCRr4oyyY+GSJQasN6RNwdDoBMDE+KgTCD
f1QjOOd5zzAUyiyvSCqMiyJ+weL0Qggm6kHHF4QBaM22XjkducavpPPjybY5MwDP
N1ngxVbTkZz9A0vCFJnctu/ccpGcA3eks8604+3v6EayCcWDxH0ETfna1CX2AG2M
IpPZtDp1zNvfvyKyAiboaNn2OGPKQKtHD6t5O63MFGION1+D5R5/+GWBbM1FI3F6
NzPMnJlWfawOuKNHnZythAqCMi4b47tGoQLaKlben0hZ3607JX4Bjlii1fjYYedp
bzqAA+qj5rXO7Lf5fgupYNbtrWCaqxVQoL0z+DG7dv0WmyV8usnWZuP527mvytd6
7qJ2/SnoCFkNii60jwvzAwG35HhB4LMUitPPziMhTdMvkwmGYT+ubgaRnlW/UtJp
zGFOlGUeOusOMLfbycIyurA41XsK0R+MQ69so0BSomvouSu1+cVC7M93mRo0s0mS
snnOTt8KBDFAvZjbLujtoiGBXvbD9FjESj+ZC+WRzN/Ef/r4gzKh8v/dI2+y+/0Z
If2WR9Zd3kD4MWrCKq+kT6GsU/JRRy9PUUi/HRqd9LSwKVN2lFAooHxrfrNPGH9c
bvyaNobWs/tqDOawiIofGotezfMbMdUs78X/KVqPK2H2/3FApBqRMYeKqD29iiv6
JaF1Amz/9UXd7mRAyi19Hff9HWJmSY31yxRh49WHRxmM9Y7HzdcTPmgikek2W31X
wvpIWsjjCWOHIx8U9btLqlcc6qHQ9TdZ9COUP4bzyBYcErKR53PSufhDcEyu3aG4
471HFJk5y3JpurQLX5n2P4VXuWyS3/9F/7E9wDUR5tJ4VfhxqFpedUZ/HMS6ABw5
Uq84noC1+TEHS64mDJDpdtmo7xN2giotEqxyBd5E/wwGi9Qi6p+jX64FYuroyiD1
e1G+KcU/Glgp4KmBDnYJwcFuPn961ncRQWYpMnhnJBg9h1OX19ICd0aAsdoE2AsM
9HAPo3/5kfIOEV2gDNzqU4IFMFYNQpXwgQpTRFDFP8ZPn65BgEvVmTAEqKKzowc1
0xIpxJd/eGyCQbjiC8jpy4wrvYf85ly1sRrsMW69jiDZeGPjjl8EBTFwxqFitVha
TSa24Ga0vwIlhL2NxTR3GbNShtzoRlCiMx8pXdDABdWqPPEcxuCetPjQd18zbLix
77mEbtWxWF0+Nz2/nukVH6WFM4lpx3KtyJENRstvyB4=
`protect END_PROTECTED
