`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVq30gvGC9qRxLHTPwy9mU6Gmk3ie+6bc8AJDqFOfHymbSMdvTr3ba2TsVkzPiWI
dYrrd4qsSqmmoyYVc7+Tcp0JqBg6me7hY8fcnv6r45CCSrVdefP42mG30HErerJv
s66z8R5S2+HxJeupGkPzTv39i58JoI4p47sG5oW6CKiI6f39WIlah8eTFMakoSe0
P/vKcyIWSGKwwkOp48HDiFB1DcleNUZeqzSDoLDVi2cv0sVtrXrzr2xESVtLMX7V
PBdvCTOXc1/prsBW3g/FmHAoVKaxzkTjy1z/11MnR8Pc/SiyiVlYS5cYK2GIV4WU
OniDcsHXbHM+c4BO7zegm7EgdDuU0TQfX32IAy9h+x2hBEczHpltYzgqH52NVriz
5bfKIdB+zMkCHarUPFBObZfIIexlqEC6oZrLwGLWy+IusnRx0s0agXRWVzRVRWrW
hbqtlzH/sJQ8oj/jJPZxUgpDTFyfDP7duRaLyOrRrejXirHI6nHNhlTuUjNK001D
aqs6+SXduCIwzfQlxW6W4F+Nyo3NBN/rhsl5PDuk+hRP/TbBPIo+bFGWxxJqFrX8
cqRcwE95sttr24d6cWfHBgf024R+UL9QdoKStdRN8CxjuFFT3a8q2a5LhmAwaZIW
Vx8TrRmP3TLCnuOf2l3uSTPvpMSbwlTvb04l6gskfpdhUapPzb73+1raop1F3EaY
7/DtRB+GYY8i1j6bJOR2iwyXypBCiqlQuYYlDZC8iVtxVwnCqxzNduq0X27qYxW6
WMP9AOjAY3sNl9PmTdGy3lT7ztDClL8TpuyNCA/zkoUU5SdTIL89c5Rd1PfGSvwK
Ax0j0navt7BCy3DDPbgFb9vg5VmLRFMk5IcUOW7m1xnkKz5qAK9hMOHKe3KGod+U
/gv4u4AH9AKzvjMa75c7eI5KYnxj1pouooYx33dazQ0eH0D9bO7tGNNp0SfHiGI8
O2rO+7U3sp1szxRMD+SVOjw4SMpCs1WIltjXe2cL04VwP+6Qknx4zXrfhMhUazNA
nk44QVAJcBXsg45dQT8lBK9Xle+WzNnPSfDdb+JtwSXfPVA0ffk3Nzx34csaliEO
`protect END_PROTECTED
