`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kOvhlRRMc9zWBwQfX4rT6lzWr0t/hO9Nuf5V8eOpU6ryn9XR+oppGKopfH/H0TB/
ZIUbSOVTaCaXnrGpG1F9Lo8VSQ/cZ4qeVgHFesShUhUdx0c2NyTkvxKMZlHmzQxF
tmZzqK2tFJkPfG55Pn/MPmUed07tmQBwHtQrzDzwjf3fYZ4uYydMzeDvvnVLtBHA
B+MPVMlUFx4p095BOA4qRT2lEqpr66h6u50qzBICcLA+gryqZMrw/zEBMm+2flpE
LbCkXaROfEf2M9A7NR3skZGqRwyy4lZ1zPEFBHxreeCLrpzt/dWAkE9A/oc4hFcx
v90PSiWtn2f9Eg1l3fakiIoh96zbpgVht0iFz8sGcMYzC0ycY2LCvTpp0cfBlFIl
8s5Lq4O4wCGv0HkSfcvFTb6ft3rmAuH3z+BRKmnyBmZzY3rXXIFcauNIcVGjG/fr
6oktOijM7eHbkSLqX0sVvEkSAnSsPihIUm/cN9hLa2vJgpEPZe6UNBpcHiqUhUhd
Qm4aRWlkoc1tbL3uhmKUev+8FKgmSP3UVPHL24aNhJY9HIVCh6Dn7U22XIin7YIV
v2/itYUVGmYA1jd4UErepP+MS9weQ4EwlErO76ZDut/pgmgq5HwmrMqT6BXyY7Ai
kuKcqODr4aezgWSYr+lwyiNMX1oMqvoVFEtCO3GM/zkbaZRo4yW0Egnep40Jy7wZ
SeqCZQLGOlZIe/Fe8GcYs6TscsLCTzIJc3RlitkpMkCf4E+lD0Lh+jZBxT61r7YD
QZ3f+CZfweXkSoM4VMdEiUrrK97/AqiKOjaA29gGsmFXItUuC+dSEQCCO4RPJqQf
PF3lKoWLdhGP3bavb050wQAq7MDNG0JiK5HsNSx34nMy/kZRz3S7zxWaauLp2YAm
jvJ0yQhfBaL9zmtGnfxjWc5Zi9mGkQ91HA0Bn3rgL2CsoPIDJy+5wRh39W2WfEkf
UU7ZEk5JDwmz8DRcWhfEr7x8IJgWpqbGgbeyB/9aYQ+INznFemnV0DfVhSwRQuvg
MxKGUqXYnLmiMysrsSJsl9ErYsiNbCLazSk9YUU9x+16N7NS5xbXLNveV8NK09vr
MmqTHi9XztzkAp1YP5zBhw==
`protect END_PROTECTED
