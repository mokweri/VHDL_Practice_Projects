`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PJ7p79snYygRQ/bo5E4tCUrvYsGCN7rCEEXJSWx6D3kEJ9kHpJGn+uLZ65tGU8nC
+6TCT4821mFQpLKsPt5pLMHGg3xBrS/2QzLEST9o5WbyyRSkO5AELYYBFst/M3+K
s21zowzhaiupMYpGdv7TEIbxWSG7xSVKB+kAhhL2wNKitvxfryPqLOBMtPs31HhC
wdWv+MQlejne8QP8IvXkrqW9iVLF+qw6Yg6LUNn8tHZEKqSjmuubQc4S+HItC+9H
JK+3+qSWra3EELnvNT/xoVBSDPYLhQox7rKcxveEZk+lvuwubHBYNChiTVSoc823
tfr6nrK1tLi6cTEHVrdEW3LrC/iuNN1pf0gS0oqmgLMKk3ibheZ6qH2C2BT/7fwp
Zh9GacvzZPfJiZdHFnJIDCDkaAN2fp0n0QElOEoapHy5/bXlFl6Ul3nuP876ZZK9
sXO9hpSZCoxFucInEsutZUOfZpbVBswhLR0HrkCWFRGMTxpzUobxmvJTPNgP3Irh
Az19EHwV/t95v2jMtGjzSkpkDgINPfysLQnS+GedDjO/cDmwvIqi10CZ8dWftIBb
dj4w4gfgV7aiGCiFl5IgboMUEa1aLMHlmXrCAYp54xxyepcfs1MqUIxCx+4qGrmc
jhOYhk1kvge3YR7eV7eq9WF4JFb4BPXRcilXXaEncxwCY1gpkYhUfPwFxTndOrV3
RRHjph+qBDicHenDXHAyk0b8HpUybq5UAx+2vObHT2BW8OQxkgfFhZH5wCr57s4u
0L5mFM/UKkrl+Ar9JqxM2sAbGEeC1wdGwGvDbCSZ3PwOX+jpDssdi0d2f/Zak6Wi
TbLP9vqiO9TPhNYwwT6SXvc47YtE0vvXgf7h2dvKDc/HtTUz99mE+Vrh0ctSvcXA
FtRKvJ0DO9dhBrhf4aG+JO3/05vASsfd8luXdcQo1s9Bj68omMQYUkVcSalzcG0U
Qfw0YStuNZEYs0DKRYAQZs84kQHE1Zsw6xMM4GBikXUJR9znraIOH3uCGWTm5hWe
I0seMS+5xnl1MRlHPH+vKSbjOIYV7LzQzY29Df7aTY3y3WDc5sd7bwBRlr6KxeOv
BkT/fn+yU4IQrjJcs8O7BFZWs8LFD3QCT6LdhOuKpt62T3Fm6PL34ZD1CsTgQBMK
2+EUOYHlYs596wXoKBeTbmhsn1DVZ0k42GrAvUYpqdZnbtAu3NS+M3MJWPZ2C+ll
lBfZOq5XcXB6iGmQs8XF+o2u78zOrN63A8b6WLV1R33JEkb+EmfIQCEfZN04DWUA
IIadn0HAYXcf1LR3WhD0LwbvnpuRE810RMMb2SofDvnAOIYE49hXhVpkx+kUn0QX
Hp5fLWtJYOX7RrADf5wfRwNMYv0zQ9T2VakRe/QkJgsSih8jKcZ/qKv6CGKCg+2c
TPRM5lnz2dY4iUjuLX1wpTJNnXWjwbX/cn6pCHfajVwgyV7CXCh/J1TrnH05eUPu
Z5q5/fFa2N3b/z1/xTeBflZA8nOZ4tn3pTsSkMODxAyU1GY+NPNd0SQFhKZLuNIy
LzEThIGJdlDp8+Zt6xqatUxy7x6eQCvNPsfUQfrVFgWEIRS9g1Y51YTXkH9d3ubd
h8uULnbliaX4YhShh6jQtLP0Qcu+5qiX7rKSXrGCwVTrNKr3AlyaUT9kpvrMG2vs
slEY2GxIbL0PFQGO9Ue2qaLxqlpjxHRe7Iy4qdhtPkAxXD9Jy5kpWxVQlwFgQLb4
PVcNo3qNCOOZ/rt+zgORTY4H8xE4/zr3TFmohBhtYIovj+/7mx61Hiz5Of1ISi3F
wbK4AhNKrMGC4HEhNzrFcf+h7M9EXbDRgFVyynUHM6c=
`protect END_PROTECTED
