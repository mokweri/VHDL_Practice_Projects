`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dCivC+MFicjubpj6W0qQ6MFrYJmuNEBuipuy16iIWGz0m7NOzPc2XAl0wQBXkq2c
AKIh/nmyazRGtpDIXeQ8Ls/SzFJJU3n3OS87hjEZq80/i3cgmxIhHVKcjwIe5kog
FONMQS2W7xaue0yEBQw8gEYjmFGiiUbTrXR5P395KC49vsFn/Vf5y70q8QeOS6H4
MA1rKNdkW+1kPGpjAPnVc2rLT5C5t3uEm07RD5vHg5Os1uC5DpAoJ2N0ABlHJZak
y/AKf6n9NeNTyeEDHDdmbPitydmmAQXhN77mLD+dkWDS50issyzDBgEO52aGZtRA
pZL/mDWAYRI1LEcsiAGIKooj/LXq/aOd+NSXg/c5O1NatXCoutLzYSBuq27Ocrou
Q7XSZOs8AuFU+FYZqmB+25sQ7DBQTo+7wrCV0IaxAJV1vJsrp3DrdQej5rScdm4M
LfMaqv1m1sP7sxTUvTFUKrYNW7qS6uYDuEil+29sB090/hr8WHmNbM7WwHBGa174
4hVPmFTBQAEYctr4mtWozy+foDOqyYGEN5mH67Vtu2GzWDXtsLpisHxObjQyLdRl
iJ3+i1VQYai3EE14vLdZN3MWz8EQe3mNyWlriQIEqhAiHou4/UHokPs6Ab2GZcsB
LSHQZwpdbFn9DHNS1tz62NXjkUOwfHc1LdrgwWTN8Zw1ysT7Yaw7Em7inV6m1r8Y
H9E+QVjWOTsvZlLC9rIr0F1TmNIqDJalo424ZYRocLg1do7mplrE78Pupx1l5pgn
OpJFc/OKS6OjprcuNNDdChpU3X6t1ab4nSd4zKsdk7jJRf3TowAQ7Cz8lQu1EtDP
8CfkHtyoPUz+DsdVdFRH7G8MFghRZNktFDHP4cHorIiXoGgETGxuOfg31okm0k2G
ofSubf3cnnF1hoYWVEQmfcuiosOr3qV1iOlAMwZXF+RWtNWcyD3K0tEFlhL42ltF
Y7JqdAk4CSdlcr2Mdsyt8ybksXgwRa5kCEnOFAz9H0W3J3+Wq0BWnWM5PV+wW8Tp
DJmmbxcGHRXWSFYMnQiv2HDezsnQiKtG1CdlFQeMXJz0XNDNXVyYAWEGEtgy/Yv5
2I8j6QJiF8dXrmEnrj5xjDz7mgIqoM78snn8roJecR1yFBkj6+hBe5iI0d+VSbNm
bsdYyKvvJqiQ3zmXYV7Gl9yQrsHCvyEnBMFTq4PGv1sB5Yws+GWxKRod6F2ST3DE
LWiccuJ0adAhsJcobBJHK1bt/k2TMVE52vuWbjbX9tA7/1gIqnKBAyE51GuOkEaM
uL56RMTFZ9g2+i80ErrZsPjePZnUvk7bsegWHwKlU8apSPqW9sIjlP6JYskwkki3
wxxoPThcD+KWFmQzEaT1CpZKsh8vNVijydPH6ycJGZk9CPnPxb4L3lnKLWLgs5ii
mkgHdRYOsQNN96Fa7b3b/+lzvHlWnYSdLMyZNNw14aGlnRvZpOppjlW4CdlMjbl6
k10E+tQjxl6Qd+XAzwmiojcKYz3woyjcqCZ+QFg/+4Or+rircQP69nruk1y0gt/Y
M3fBBadQ+gXAnSZueGicC2ICWnz7y3hVEWjxZiYkHX59pmXMYDMN9432Mkfpgz6s
RK8SgBbLe3Dxid6RKT84sTUXKKpTVHBcy0ioA1HslwyWUjM3VFxjvdXAanxYKNHR
ccfxyeEG0CDB0/uPKM1SlTIACQVsfLeqDuHbSsNUV1JnU7VC9pvbXjwC2leGC1l0
iOi5mKqh0v0PXnrOGN4CRtQxzJOZVxlrui9ItUlAQHrO/D37SORLAQT91BKhxBEE
HbAu/DlljU7LkBxFFrhrdZf+YKye7jmnh9KQ8+XbKcwqnb1MfGLcdjAc7O1YOxwh
l5qC1lxOBMOL2qQoRwLsl00cqeSafjrpZ+2LpgR9Wt3Rb2mcxoWqDv91lLzNFsLj
hPH0LdKUrA80wptZlACmT8dYQkJOwKZI2OltB//7iD3v/83UY4+oCt85Iscywi+A
CUzxGAq4+BF8iaG/lZJe3NtXSnoHQhowVSWggp4ELAGARF6BOhAuE+hFmLa0NBUE
xwRKMxV8nJXLgL2NuoRMhWpm3mYk0qcRpqlEtTPYgz9NURrE8Gyj45eMSC0SADpb
t2Afhd2V2qWPtvBqBtP96KDydd5Lvatrhzal66FI/S3R69t2/yy86YjSAM4zRaUu
78mKQvMsq1CeMDUL+DrBJoot8X0EmwdO5ihnqpr8+MlYEnQXpY/uIyBMcKFc3GWL
EKg22NgbhewC3et9l6iwH9ffacznMXyRzrwX3vikD+xsrOcCUVNWmDSoUnqjT+Zk
3KPs8bk/WNZkeXY0zBLD/S+6OIjbSUgIKxJuOkHUfUyBEzWr6QIbawoeotfD10YA
nz3B1BXtO87L2w67x32W8Y77Moq9oLTAPBvoWePsk4C6tUyhZ0jsMXJwpnOk4vbY
dqpkzXSFppa+4K59xGyyiaummTEa8DLVhamwsqGc9387a9+hsivhhV0VbtcmOgLS
KltyW6/6g2xlT6ZJo85qf/JTHsVJY6dyPHvYGF6uDJfqJ7d8KdFPxyznnI8KH00i
SnPZkjxO4nWDJhqmwQK9sRMmjMtbJYu3pJDGHIppsrNJr9BiYWnvYCGvxw+0M76C
2q+4AtQvKcSzKH8OhCmYvsRJwHZnItxSEZEaHbyx+fyPzpOTX2/azOAMJ8C56R/j
iScqayG6WOoipVbE3vNj62wPvNjiKxVgsNeW+BFfJnjHalUQeaR8kqslsA3VRjIN
M/WxjAkToTNoV+xgceG2CY1/8ecuuDFNK2Q+Sb+KYzh87IJGtaob8ifOANRnIz1h
PNMUDi0+tTpECZxBmIIg/os480ZRIElUuVKxf5dTo4e5Lx5XCftEeElul1ZZq6xm
SBHsGLcQytDRl8iWOmuPwsbiP08RWigGFIhTDO9GtyRibb38xG2TrWgajiv3W7sf
l8Q6zf2MhCHVhaZ0jfuJFxC9LbWvu2LcHh/f1QpAo5xaVjx4nA/pagiuDNqQqKlf
wVyFxpA0BhZ0fKKzvdbKcQQCUbCuHQRLXWqgH///fvCMlYKvx4c6cqV8YsgBYuVN
cDKX+etYW4RnDeJFsHJYh7KUOxq2uuVPhDEWqtLy606YpbFb9sRUkHtVeWKMrB0U
s393mnar22PzN/BCMmy4qRLSuW1lA2KIHQEispbkqd+JEUAsPVjsiu4i84NBZo15
IO6e7UQE1mHhyKspSTjbG62BQvIiyRo4nq2S7LphXVeTyoNf85GaZ/MLRcVjHPK/
b0+QnQPln7js2jSEHsm6QvKdi89pT8Y20C4TRPFwjgnr2sgNNNVXqj//6zUMWe/G
DXRkdicqfAxq+wTMo2//fui7spzQ8elxSQmcmouEIPJt5HkphKnGNTgYAUqzj2Nq
NXm1wpSLNYCcgzDVAOsRjK78y+CQ5kPPV1N7i1lLfBMbM48RLgiJOLrGrejEOvxf
xfasIbv1iPF5yjWzXotvLIypMFboa3Oq0EPu8mOxGtafQhE7Hretv7VptEoqF6a+
q6V8do+5i2u3G142OexRARix2SanuBxJn94dDfLY0FOOunPz3vOGvIt/zEy+se9p
vv5fBZH7JPtRNRNwULfniPBYIDjQIB6PE3IvBdotQ1MaHfd8u9EOeItdhXegNDFw
7/2S89XJkd3sdGM6niX29dJw+3HsJdhUlTcbSLmaKHeJ+GiDCXfeXqxSFoF0rCDH
fueZ1Kl53YcK70rhQVbWDuSCRp29Zm+A6CQL7tZg98zBQFasI08dnFIqi7dLmjlk
RbJ4JbpMp7JLqTVPwhXkwrWHBuuofSOvkZOH59wYZC28q9D85ocBMmIf+0IY2nRg
l2WoBS6GpLhiLRZu7/tOmWt9EVX5E38bdmQ3hSJobSqQV8qCSCPap3RxCMwXoSH0
x9Vc5q2L4YTXwbz5m55IJMaCfx7pYqP9n+kXYN218edDMKWZ0Jj023CS8FvPLd7+
Ib+8SKTEj8MKTBmN1+gxHpicQrzguZBKQbCqHYQZgnUUUFsdJYo8zNyERxcflfES
8ptOAuOzOqm/KA4w88eiIUVUjRj6BJl+NgUwiw6uPLBvK9o7pQs9d00sfvas+nRE
ha1LktO3M+Me2c1ZWnYWWIkHxCxDG5//em177+kyVEonYFPGBWNjaMZCu9hNycwT
wJTZKGdxpVZNSQfySI51G0vQcqsttMUdYUoFvQjoqx5SBmJqrqd9SEuf1Kmly+gl
uDzm4j6NhmNtIBVr5jL3Nau1dAERCyFe3NJJNGEAcTzCp5B5UWLEjR/CGd8lH+p/
7xdDqchVeUyuKncotSqhASqH4gm1b5uKbpOIjBlZtYS/xc74QSAKbeRJ2uuX2X1C
mxxY52jRIpO8d4E4fPPOBWCOKBqm0HZKAcGwhZ2ZvrXb5tu4XVEMUrwbTE4qCkLH
IMpiT1sHgPVNb7tFIXtUtykqvxviUmY3Pz/qGrwp6bcwxgsdxqzrXShV4AWG/H2k
D46qBZHpYvIOkMgTJNZ4rC0A0HinoHfnx1Ancz7QS9NhD/3+zWSETRjpWgKXLtF0
LRZCJsdvL7+WjrCmy0Mu9IFO34q5K0U6OTzZOeQgYe4vdAWSfelgXKmKZAwiMw+Y
UJ27VNwWi0/wQFsK3Cw4iPcdpgA6AaP0KXHBvzsC8WdofcTzK17X+SatT6GeQNgo
tlhEa4Ws9EI68W5AgBQDKf21+9p+WTXzuagzOFHkybQco7UPxnFeWRjSAuEG3Ohc
K6kUR44GkbTY0xhZJ03kAD9KVKQB6umuWkaGfwKM/qP+2r2P3Ausxs5CGLoq2iki
cXcIAmn6Tz1h/OG2tls7YWPDTLaN4dq+lsruDnP+QOrGZev5jK5JdUvr++5EW6+v
OQfwjz8tr7ik7oyqGBsuCSQIBa/sFOnB9bmMDkmqQU8P/wJlnyUjVmy949e4/NDH
6PTlg1umrnIQ70zvAqVy3mXHA5JEfgh9SCNOzU6JOZzw7pBMOEd/Cdl7bfrlMhzJ
ppTrE9O3xa7ufwfa6rK1yhVbeuEFws2LXImUnmJM0bXYFNBZaSFaPcUew667lK3b
d+ZyBukcfVOBny7rTfr0mdn9oPPDFAjFrXmy2rEDCUfTZjnv3/q4r7icp9KBuwqf
I4DQUqCW/IAt5S5DqDDinU9EDaCCt+1ixoM+euoDcd0bQkQ2akZp7dCygPogLkfK
erRMRzk0zf+RY3UkoDwsrW+Yq2jesmAqjlueivzZ2+CbDtnHwnpx8aPqYA32mjpQ
louClijhb9PCkbqa7rk43bOfZEo7KYwwsi2jyFvws0LkppbRdJKOayc6j15tPNkk
D7Q3T3/m77H4soS15di6CpLtb3hAHJ1f0Oww41Gu0wiD1mxu5lOQoq6B05ciaHNu
XV1zLJDV+d/y+cLcPLxh8N4XbQvINzf6ix1dQXCdLa10SGrlURchWq061oBuZHxO
UYTUr6F/uLVR7M1OseQhQ9IGBPNvO5cqcveK+zxdqGmjads/GAt9JbTyu8RC7yl5
Fqx1AQ2tsfUcDxfp3rytaJtz8+KAqCbIrOBNedbAPL15DV1LW5QLtISOGrBHOfWV
2rRcC9zvcTQ5Rh6d/IkbkSeus3mjnIOlnX5XosKKItIneGPZP6ckYIHlFkfp+jRE
iMCAvb/kYwg8HcW1swoAk2gBNLk6c2EHgnQnIYpyrvJB1cQuep4vR1NPjq0E5Ir0
L8CL7BsQN9iUuF+ODVDlerJh8gV7ZXwPzl/IBnruZxod5GYxENm/gEfpZaS8nDeB
+2xbTkP/NVDIoMWgw+s/lU/veHM9Dt9NdeiX6Rd2zj/LPZxPWYPs5n+NUlica/7u
YswlqqmTDx3KU0DPiHrGgwpbfR5BoYxVWrxQSmtAJW15hzXTE1HKO7it3uxiswxv
qHo8mzkJw4dt1ZJImt2PgVMOyjuYOedOihzSAECQ3irvogPQg55dAHkhTWJkG428
zdWs524wFHzjsUqNefO4sd3KLP48mockLhMA/sdGfI7OO38eG26wjDEDDlpqVW9e
7K+ljsxJpUgwc/vwIAC6IPGgeyEaA3WBZT3sp6h6HoZsU6bP9EpFuns+LJu0vXO5
kd3Ik8zfEtV3boqekDqUygu/5IuV2EMoSE+8eYyejte7iYdXt0ncBMWloG3+qqxM
e1Kcfs71b90c++RXS90upYRO6hk9rWQHG2Rkrw2c0s05xJqonJQkePduwtNlqpiz
v817S5FLuGTKB6hhRugpDOI83sNO/tsqwX5hn6aYzophFJw2tw1B+9TzARcbGoBx
cqi5rMYUU4nl7S8x96TFMdghO1kTYnLElYwuWo3durW9hm3B+XgBKGtYIhyLKCFW
XZLph/onERg1YDY/7i0PhyRUivD0ZetegaglYAe8DVIT3HI17bB2UNcDagsjxHo7
84gruTB1sXyhGsrWJgAEAWRcnXJ0i/UfJ2WPKWukeE9gVHIv+ug5Qtk8Qvw1xbwI
RRRs5AcJWmZJ5YH1/nmRBsuy6dg2tuBXlb7BIIibA57NI6pmDE/joZ8s0wxudxpu
07vM5NrIVXg8DCVJ5N+wv5X15nvZv5R27qc1lNBZJ69Hhlzad2umqaulZR5KHUHX
uNHV8u97Y+pb7lYQltyiKR4ts0r3rExr9keIvF4qTW3PfUigKOFq5OPiYZNrbUYc
P/ggxKWvVqeYSYyeA22cBPbrH6m68EoNqQ5TnhhE/z8uFWxfw1S/jUxe7CUMZv2c
73jqNz7psTMOPt14j77Tv1W7iJwl8QKDiHIuNVl0sEo12NFo9/PBToFyAg9Y0Wo2
a9dOC0MWKSRhjiFCcoLN1LMLxxMcmBhez6yFWiHw9Pv2s+DJPLFC80VC+J2uxTli
9Ro6LrRYYT1evDntnOMUi20sqYTMyeOnm3CiDiA4ACw2aVBwcDb074wbgXc9vp9s
paGMAEXC3KsOZXqHyNCMi1fAHNTj9zoOYkg0gbzzCnkGLD/bPM/KHNkDZcorzVZS
B04XFZ0PzXmS5l4SdPMNjhqdxPldzoXhBZuFHIEXu/9FkZ+R8T9jacJFfERtOgle
UlR+3J7osNtHK+masQRgxH49gjKwJ7K6rDdrdh/CONsfQMEsSTxmrn9iDtcKOcbH
r+X9Qm3vSD+apO+b6Nhb1cYbLzHr665jVq6L++AzaatY55WXLfC/9l4GZgVgJG4h
ScmDitNEBn2XE0sa3rtJrQbxULvcxiQihd/ROQAbj+RSHlMsmrfQIYvNj9C4yMNl
bVRz8xKgI5cAZ5+tNxbaJCY4nvDpriOv91kljy40m2uZryLKoeh8cLHK0TtmDF6i
nJ9s+jNl8fSLeI3WHZf866xSZPCQfSmVA0VKcZuXHRMtc48tf2O8bKzsPcslSo1b
a/v2b22TPRXbUmNQ009yrtJB8s18ThdeWq9JOxkCYNnHIiLZvW7JrtVzLMxh5aYn
5S1LBefOVAFBpFizCMMmFQXkRh4XIAV6LXthr6CzuLdDYQLUH4AyeTTTE0DRiIJ4
mlSzLhN+NnhjQBU0SnLk7t++JrZvcMIXl8+q7AYUyglliW+l8GOa6Y7AQPnoZ6fn
6fLKuFNRIv/H92hldMApkRCHDOaWDQfKyv1amx5nSJKc8NS8M6vpOye8Vzy4CW0w
fdudG+QcT005Fjq3y6GA/bZyZVn89MN78cSkNyPLxNCgzIxWkdMNYo3fiTTYV3OX
UmAZXseasTxpRF+5rqSH7MCMOTqRSS41/zLplhyukN91/OJfofYnjNa8/MbbMQj+
WW+WAa6QVYRbJwlk4uneuZipqcgwgLKEj1abWgy2uDfDvW9zOtFCO79F8EJvXFzx
qvmPZrw94FnAviacSOxdWoKXodROdgZ4vmU/jaLAr+K1TdW3qzKSqi/kX6R3QLrQ
x1J9ARW3/NHzS01bfPR6ZuBOXMZdjXblz7vByvgujlAbswX20ioSeIWp73h46KOX
7SwuNjM3dMEhed+9XRT4XHMd/3+fSZEaHPoUDi5OTJjtdjjfopHIBQAOCmeHBXrw
hR03PjzZqQzmu8qeBLnA1XDdaBBmLebuAXOT51bcyLxk2pFZmeJZUIWiY9EpxARM
LHi9np/teDaDUEAOjfhyNQ28CNRryi4Syx6m82qoX3WVjInDziaRa3PFQN2V6pUi
idqJjp1cQ0P249OE43Gv28SCl6b2OrEUzjQQgo6f3mU8TgVVXyhQUf6E2rrcZ00n
xMNWEKhHGcYPQdIMA1U9yolOrCshqCfZcvAnO89VsXa1d8xBTpINKMYvHUsCOkm7
OyEGxYAYiJQsGSHInOR1LAx47HSQWgh4y7q++3wsb3UD80Crl4Er1AGljXbJCFCR
ay+kd4W3ZsQmveWHE0MBTEgGbqayfhAx2i0itD+LsZbhX2lroNz7ipUkHrZFC1Bx
F1mhbiBV1uAja1Za6C0dgWe6uErUPr7ij8EzH8Ay6piL2yNyTW/dp9ycc2n7/G7p
OykV45gtzR4umcnpTNst0MhZG8NGSBEnJ8ski0o30eWJbqlpCDcIwPUbOXePY/mT
Vuko85dRcpUOjKtaXsIG9xSJco9c1Tg8R6ze9J50LqxNs4km3PpXZJv/HhkF1QfR
CazpigLBxda+S2LwdbYqtRyFeLmuGf2ZcZWJf8+gbbLf7PheeA4Gy8TTjUyDGS4Y
qiCrb/fr35JRcm28XiyXrJxzMKe9H9vWHTmah/yoxecC0sf6BfjuDU48i2dLBFsX
Rb5ptb3QJZD4d96yswT9xP+bYDFn0ubp3S3Y/Q+o/eA/0Jd6vEPv4k+nemryUxW9
N+wFxzq4JA05Mul6LzbHWY3StZjDt1BFCQoffVgBTvrQeamcgShXVPQe+WSdSBo5
+bRg/Fgpjz0c90M2tsByS7gv9PSNK/1X5L/+Vw/25bg6Vl4QeIAujYKZYv0AozUk
LpFdiGxdUL1hsYvlOjlg2kAFcCSMaQvZpyKKJg0ZE3RcL5XDsLnsnALhq/g/rmWf
MGuUfCvJcroVIIYg7D0BgLNUZSJ8lv4aRCl87lyUq+aZRKnvGbrt3geYH3OhjyWV
JXY0CFg0EbEe8dHTnsEAG+ug3hSfiJUoFAO2Rs7ei+2wJVOtdsA2aUHihNRxdzwP
8DqdSQRT0s0sDIOvG5WATt+rXm/WkUuqFZBlEEeuy6gEzD8PYOQ9E3J+aZVRGMot
5K/Ry/fmmeG1PKw+fQmWwLdEQSA0StngvdcPeN0gDoJ3SvlD8/Ahxf04C7IOApu8
XNUjfhww2Yx3mPWKtD9ZUXrN0P547j8hpdXDFm0WMWee7eO+Uk7YetwxLTomnqzQ
OZunIE5kx3t1tnnC3q4jG/uMmORxdQv+35F7pNmGd3dvKn6t9qQ/grvNwM2wFbOw
0D1tU/qgjrqT+Cvp9FAiIlwjjrHjXcX2yXESNGJ+Bw3MPtXd62lYsuU8qVdlQY/q
N3qpcVUaC4btm4IM2iQMH7acWUsG/QFPTAlCnUe2ZialAtVU1U39nG66SeiIDkqa
KHVDT01Zow92HK3qYICIXELVzuuFoOO5SrBaK4/IVUnlqY9Nd/Skr1yW5by6xdFT
PZTd8tq94I2F6dRY/7ipxRq//ODD5j1Arj1QUfUfvWWiqv3Rw0u9ADJxFDwe4ciI
/A/hhfhQHTaCI2FSfB2IcHiKweVi10h9DUzF20ZlETD5BPk79fmmHS06AYiSGQJm
htcQrqEs7IXSQxmtAunmSW9kqAXWf+82ZGHO3S0rwEfyHHX1MIlfVHxeYkVoxvV+
zPlCvcKb/58DvKRi/yExzixFqgp+IankkCvPgpxtmSYFID8hqNKK/8j2I7DACkBt
VVlqTAtfkG9FmGXoiGpASptUhzufiblRPZ+k8m613EjIPvSzg7InT+AxwlGGBi5w
fsT77Cd+OUh9sLarob16l6uGvKq5z5Z2F5i0gQNbgKmOji8dxmjk59xyzklF3W7f
OoDxn6MM9IsXAcJOK935z+XRQX9KRisum63zFLpevOCZ5xr1Ny2rUBnMPQL/8dgQ
Nry6ffr+g5+elL8VRK4Dw2KaVwfqJF9BCr2PumzP8dzDH3OLGfmrgisujheazvE+
dowaVmt7COZ4Mset22wtEeJXRHZ0U+LrgDVeJoQh0CD/7r7s21NaDb1GuG+BjOvs
5Rk2hb2bil6p4rCVCuQjyBYBnsRCS6ycl4tXuj9WEICHuhG++kGctX0YerjcrpzN
SjxB42FIyTDpD9c8RhEJJPHcS15q8IardvsKY5R2Y58IP/E5/wUCORWlrGtp2YCS
u2QwBBLf3TtYbuWi6UnJgHk/AAnrlbH6r3g8jjuUZ1y3S56r98REyWlt/VoH9IlN
RblvY93BDWIxMwN+9D0Mhgd/jiAa5JmRGROiNaQFuPfHEibjuwChUE4O86jQtYtC
zWTAlMDm5nGzBIKdqIKL5u9/B4lr1cU0QYH9bdnflIxWxGpEnESQRar5k1uBYRjb
Hqy/NBASbvO9AWVswk7usbDntq1Bh579Cpn8SmGKV3ogov59qFxI+2g3PZC+0jNV
RODuOo63WMs5qVh0XWKYndWwbfmVUzRwt4Hk6GCpvDSXp/JSUSwzBAQLw1NRfX2B
mlQvOPd6taFLO80XO/svnVjlnhr3j+upuBdeoQ27po+Alxr8tbDPs4LUmyIb3OuB
/B886nku+oV6Q+ToHKNMXZfvcmH0+aKgW/9LEDEvpcg1YzzV6T8Bk94j4nh57kij
VQMV9KFVd0Bah0o/qZUJZ7pti8Kod+f4GR3rbyqge23AuM9PUtOGfSn4PSPobMPv
vcLJSF3jV/N0puJLEbyAUyO1UO51TTkgxLEOF7px+sxTDCPnWG33zjltTaOKSpfj
NaEqyJx2oKdc4dDqhl1pu+ld0irMLpKMp7ll4tua8C/UuQjm0kBYPbf3cslcCJj/
AWULSOD/NxUjv/0Sosf1NZBMh1DoiFzaaYcNpAoMc99FEC1o4Y7RJNePPUAWAlKn
lcwxp6TXyMLh36VLeGoCvGsWo0pWifdGTkoptL7z70bBmSWO1oXz33fsXyD9umJV
6Egz/uRC3z4+r3och9lB9tc+wLwK3+t8iFE7e505e2+95Q0CrE4cz8sSNo1uJ/jD
D7a04VRlqoC8NrgSVa9aKpBsB69Rve+kidnuGpSHyYcDU0Avcq9AjjT1gNyT7P40
7l+XDAuY4hFKjU0j6qlNSu3uEMvBm39Zpyczy92UN5pK2TQA+lQU10YcKtXXCqNQ
jSevPk2aw1OoY+RgOmm98DG1sxoPBK/pwpB10WZ/x01GJpaC178bnZmI2/8FgDmM
ZmKMp52PNWbB8wb4m+sEj6gsDh0ZagDlHleYlcR0q0BvVYLUi2zykoBn/PX0tdz6
YBrkRxFGFlrpck/pJobSR1eMvYgJ/+R2bkvgtsHcZK6lPEix1VBIMAex8Lk/urES
nCkJbm0bC2SGbb9xCVGxDXR0GpygcWLSV6++kjUcSUJPTSkNLt3HOlW/SD5UWVUY
kuy8U7qeLFvEM+TLxYo6VqN0z/8VZN0HU2vFa65xEBkh2d3COu625f67wVhwgMCO
m6uAHo+JOi7hy+f8JPbgsaQ2WQU0jR4Rn524P+X7aaWIz7MvlACKpLMXbc6AVkLa
3zBkSPIWfEFM0uX1FV9X7lebkxGARImEeZ7WT08W/wTU7Vk6yQMoTJPNI+C8Rl9C
9tE3uKCyyhBJhJtlGv6qYCgSaYoN9xbRk2EhRaVE8/BDOBGIFrLlY4hEP/sc9vFY
eVpb4Ccun8ap1hcNC3uhKLAyR4lJv7GSL583h70RFYKbnkKJG1P1WdkAZ6e/tZ1z
AyJi40QLgeMQFngSxqSsBkNVOV3iulvksQgw4lilsh3MAMRwQKQwgSaTrWvxeik7
wU5l78tFbkPlzUeq367U01wPRB+l3+Ff5KK4m7ZRlLZrs5TJz1YTJCzcoTyyRpCe
5sHc8WC55HMSeU3LmrVnGh1rW3F2kKMe9wqiD1Wrl8GUfkRP4w2GElHLvXSC/Gor
rsiLWSJU4y4XTenMixfcs3IWGdI2iRxq0nT+YV5ySIIEvwNXXUOyRALoTalI5m/m
wZAwNEskhabcoUDfFCPXOrXGMsS4TXu7/M1D/oeaNiGcE7GhizJefyXXB4nGMQPG
Vj70z+lVqXHm7Zgag4kqMok34UX6UO0d6BknxEXwAQC/RfAon2M8XZb87oQbvoaT
C+/g62XeeJqpCmgzo/My9wU3l/qdEC2Oid20BSD+ZbsJv5K2rc5M+TXH2Bqp2Twa
KFC8Ob1P3SIMI1zGkBRng6EMS0TbXdKgMhoBta7O8PZZAM3HI0ksan9wjkZFsZr1
OuBO5HFcvIOexxe34jcYZ68gyZVdxrdV1Wj6uLMMsL0W6GOGNxcGJq78FR0JsVLa
lUtclYBHnqWWirXh8gfnzxL9D+v+P8lb4SETEf8DJqHZEG6NvDdETPJfqdCbgnRv
uf6YTk9jZDqq6jTgUqvW0NP3fA35/bS0pL4MEllMtMY6bnhB/hGYJfM1N2+SHjmX
XzdwVGsMHTUmgCY0rC7yhdqxeNCCi8usOixkwIc6or1ARZ1pL0/sdsCI3XSicPbn
dFcXqozZCSMK4P36//GfEt3uZ2kc1xKR7VZq87KBOa7jEYVgOmL3wlEcef+lM+Bm
dy5IfsUTJm8dd37Raq7RxxVr4xbGx15Avrx2Zy/kWrLV0IIwqnb0LlVsxBI1RCgQ
inZqX16PJlF5NmN7Z36ssvaBLMxF79lfoAbFz1pIMlNNW4XE+PewKvqLu6XIMY0l
HpBBCfOMJgCWACKRECWfWW8RDC3WUc+LawVCRxpAayur5sg/lTS9KTaQ4Vuh38py
3D8kdl5BCy14T3zE/TK72A5s9JYXqDpiAQa2qbK/xx44zns9hWM6+/OQSBZsIVu7
SX18dvvuLUqkIc7Z0TAmHXhdyhF5Z85kQ88crscbLZmasgbPlMH2szmbiR5yRb/B
daapiyTo22/mq51ln6i/bHDsQV6sbt2lAzAKZqRoyXOD/Hi4s9fuVIRCfiIItUQm
0JWewFuBV5XOh7fboZp0sATainieAJmuRjFXDbjSkc1Gxwf+tIrSy5S00x3G7MoT
V0ILN1YE6lYKcvi+GOtUYtzmMx9Sd2/JfZJMbQ77HSerl0depKB7WN0lU+Qf1kpF
BNGDY8NTB7OYdF+bkDZ4jJiBje4J3Eh/t28YgOCJ2p/J+YiddZryzm4Fqc7lNY3t
GsIAGkLU7XBXulRU/KcXTejdOHfiMFBOWHMbFzhy4HHr/EqwVVRhS66+E+QZH3Gr
fhkH0cLeH5gauObHfNC6Z11egRC8Z0m0TxA3rM15ebqZM6oIH1HxIphrLxC9TG11
uxdGraEkh0cemy6xwTOq2hQ7BJ1WnHV6RD7Rf3NZ1Ztn8uvAjad+h8+OWWxbypi/
AkZ1QGCCabro0vfpLc+6RMCP++/T4LRcXJ1W3DKqBwCy2cnyBPz+K6Df4H8pa6ry
KlV/X3b75pbF3ISsgLHrqkPThKTayzikuBzttsbqLmQ+Fxe7yocI7itABtuyaTjf
jmZJeRbJWX7lY/MDexTUuCQEIeD1X6a9MJG1XksjmTP77/qC7xu6Kg2wbmYnEH6/
xyW7iIHcT169mpmiODMOECkm1QhMACpruRwYxHbBlXqRRbUhDidssQ6yGSNv/BEP
QvePfH+2+q/cDEqYkmIjJDI7u1zd6EGEMItk9uEkSWKpA5gMTWcYBZVyu1r9K562
vJV9XmhOo8LrL5nMm/RTylYSTKNyRCjhptCbD2JrTsMNt72WC8+J1Tb7MyGIC8bv
XOz7JspTuu8BdLXNsYCqrdBsF0XgYBjtb3fVEZ4PgPtNzNLNuWEr7miSILJFUjG6
114Y52ZDT0xnmevM4ZA0YdCI8fdHYnIgWJ4BmwEWm5XjOE1LXlLc46VnoZT6lWzx
jkfiRxBk3WVoBuWcJMoxE05/5yz16oYxNhxX71UzmdKjZKmMX5JUfK04YbKYPbmr
EUuIp8UM2ZH+RKj5z0NC+GOiAIy7lH5QDoFqqpgSnD5tiy/wIXszO+xlLiyj+qrJ
TJwuC1AbfbtzgbsGkMciXmiCDvkOfaK5foNIYWxgd8kqQNSLXqCmjcV32gk96fJH
4uk3boYuhpwmzKUBx5Cl1P9d9ABu8epm+iFFyLxrF4glzn/c1hDupZocgvdhjtXR
S3BroI3NlVTKyHT82UZxKN/xW4rS2j98Qr+MCOsgi55WE3a/eyxUXagOk3uPLlW3
qmUOOhC5RUMqklY9/ZUT+3i0cQGx0aHji+sx6Wug3HfLm32I9e4r+6vcqrs97DVO
eHgyMe/c7mrcL3PPMU0UlsDYn2TgLCeM+TymxuJ2JEZdCxpi+ojyQ91s7W7ilqJw
GwHpEE8lahJiaR1gjxzwoU6G9biSbwPm9G8jEHXaw7H7x3LUYExLtE55VAe8vrDn
j2zn60Tf7ncf0I0Z9MkONyjubg93BB/LEQ7Yhl+MnKF2LjA3Hn0G6LUzQaw98LV4
yH2vjtvJTiY3GBaRup7epc+S3xpFo8o+AetQzixxDpdlF+WSzE5Yi3Ex1KLxUJJ5
utnY8dP4oHY2e9xsW4+yt+F/ebSpMVN5W9unKra+4ziXE5d1xPfDlwdOQeNjbjdv
D0QFVhVmdTmNeRhdUHnTsiqCk9Blcc2KMsuw7pCgucWlFZ04bYVI3aXYXF3aLont
ek2uGkN//ZnAjzsOTQ3d6Z4Dhp+aKKds3eGBHLUJZXLJ4wbPGKDp4JS2EV2ztzWl
xH1WskMZg48T/HLyBzo4kMdhVq/t+rJoI0p7owyLdUEq4v3PfEW5IAD7yt+tJYWl
6to9yX3M+9EeGji4ULfnuD17Iq2amM9tMSBxCXdc3yslpY1orDK6OpJPZD4x9G9q
zj9Ch2AE4Oawnj5Yazsj6ubtZBNWv1OC2kPAAZdB49xcC4hPIf3W8EElSDx3RYXS
SS+nYovtoWqutK/8bTL0nHxguf2d4/9ih7zBFYJ5DEnQTi8kEKf17gpmCNMxz0GH
rOdEB+IYa6PVKjppvtGxJjlQ3eMdTUnB3cXt1BkLfXGBm1ItJMehRGblVTJX4y09
s5FBPoCHxEGvnKDVB4WdrnQOMI17ccm5ERa+GB4CL89SUP1jRWKJKewdcdPn3QiV
o2AtE4IhKHJqDBwf6ZHMW3YQtyKvwPv8vKFlpTpAkuUsLi5XnPTPZIud+hAoavRJ
LnId5waC0MDljSmIxFbVCPAa+KrNLB9aqI+FWhmmVE0jRZnwAmJDVibVPMkkT8QL
EJTWfU340Gdn1OtbKYp3qy3Ck2iDRE3HsnJ4ZvdjSKJAP/jGtdCs0ullVhocBsI/
NxrYXdAT8yErL76EdGuBWNtQLMmk2kTQLaj6xgqEUXlUa3uzZpR8nLZvJR7Zqh8n
JV8ofnEAAADkhUbk/8yUHbfv6aIfg6cpFFjRMWX+ekQE0IvybkBD3l42w02i+ypQ
CVPH1XLjDbxZXfpDwZ+r0rF7XsZAD3BL62nUcCyiGeieBlkQzX7no6VQwmL3lkJM
nxAwfhYaCvIHvZT+WHieIL82hJiuDtINF3nfq69nLOusGcHxYMNjtEK1R60BhihV
T7Z2+dl7p3PeXFdauS437rBy8l/d//ZlKoHUzomY+Rqm6YkATfx+d9Qepe26ksrR
0L9e7W0crlzv+8U0qPOnIY2UZcwGB6UOmedzBxyxWL75h9njUESGw2u83k+/UqZA
M9BAt5piAKB3XLBx0JEXMYmpDTLoh7p0dMBnoPYjKOudx23uf9iiekODwcA5qE4X
ordW90UgzPpVMgovZRO09dlciwimBBzhWQVogau4EDolRVN37OkRcSk/ntEVKDWA
RGdwzou+eifEYYli6pbJ65+bNQhDXu49A95d8tad1q8pUlu7htHImck0p4pgvp1Y
sxwoeWnDE0FaU0lsogE4IrYV398XxfwsJjt3JKF75OHI9MDhq5g+P3Yv5IJ9AcHw
0DpgBg+2eeO02O/VE47v2WWf+knRssiWIBLLXiu3b73e/Gsm7cyxHcgNA9mDNjyv
eD88U+S7VoQ8NBTwqqfkxF9rh2FWfgzi9rLRu28oWMO6r46sguQHrynrl6JsfO2K
cXzvKZ1RgKFvxe4aZ36dFImXBwABaUZ1UBt9RA/r1uIiLdm3UBhqTprE74l/9Uk8
lXjF4R9DwUB4+C0HySE5KP87pc8T/FSXLru8VEyIWOCDZqiimoICC0RUnlAzCwBc
qxAdrPLpxU79Orsh/t9Km6NJ3AW3mQAxBqbc4svoXfT1ACiMUkN5g+aIHkMKYSJA
+0qQK3HSRjWdft4wqidaDXQJ3TjQ6TovSPg25rDUHU8i5nbG+WxvC0upCLEuquY/
Dd/6bVaA2ynSwBSDO1OnYcHuqT1UU6XXkekBO8bw7ktKPzCmfnM1xTxlpAEPLQ58
jjfsVtKmENkWKavfrG1xzi8CMz6cJZuvceJrnooMLU3jTzFRFtaEchoO5WwgYsY6
rq8UI5tL2NMETYas1CzS6VKlvKqGrufOHo29o3qf5pGRBu+g5UGJv155/jWm42JY
sbitnpKNXc2a7BryopA2k9+TTN4xKQ99B5DDwk/QQsjZk0OQ1IB6PNNBI07xDDNo
RXsGpeBkUQwpXuzSO+ikGQ9/DTwbuF9x7UCumueLf2LW1RO0PRMdVncGYjyT+J0y
/wIGNmukgINymPfyUHgag8byH9l7tqDDrubnxJAfkyAjB6Z3wNzimWRaA6CQEhIi
kqtNWLCbO2b08l7JpoOmlKasye53WiSavScVNGMed6fI22gFLu1//TaSJAhxh3Pn
qYW/a9s5hE9vK1wCeewIPJ7VKr2XieRbQ3HATccFya2TzNUHSmZKstqtUOmFH4wf
r7ATqmxzzplyughWsOuI7UvCSUKW6L6vjirruqWQQeU47abdrqp4WNXPCvKlJQnX
Oi/6TQwEJdhE+ChsQjC3X3KkfadpluINBDFRFZ5MERSRWoxxMidnUL8fDz2Xa/pb
XJg6wdB9KdgwmFPEqjq8Dx3V6KaQ368WSUHLgHUT+wa+HsqORAxhdB8emSpknIQq
JcnEm5wKcTOVmijySVFyAODQPR4u17a0IFLGwF2zvpPPmqV52wigqPzgIvfxCz4Y
vYffzgimgzw/DyY6P16H2swziRkwbYvoyE8XG6xhOCaWwRIkvkfmWlLex+e7sDFR
n0lkQyF4E3aYA841MOucfQ3Ai2v+9uTY61nNdak37OdXHDHHUrKgCie6kflI/3ZI
wtEVXL64EMHqM8Z56R1F8p7MRFEIhLsr2rIN4HidpMK9YpWVdNa5HabHF6te50zy
hbki8HAY/3HgOpZRqx3iZl5p3F/oyUq2SJ5bWUrZQ3cNgD74z6Iu8BMqn1LUnmX8
Pyb7LZmDwsUNz0hTRvmt2C7cVXeGJJg3uC616ZCPgGOSVb7HmAZ/yrA2HrAvwxrU
eSMI8xqVFGCwUlEib2OFgQxKUcLCIISVewccgQXnkuFFKW3hLkCXLMoZQy4RXHLl
u7Ue/ybAE49joVS2GyMbWJdgGArjwpCAdwTzIrtlMmd0fEPUAWmjAfVlWD5xcdiT
yC9H8ZJ1D/GBXEKeanBZILxH10EkhRfTZ7pHp3NwCVqN0uxfRiqLAjmO0Y3x7pdQ
lyD2Wg0fLAS+/uiuzh73H5VpPO6z3+WCoVITz7xRyx8GfQcSJNXEPG+MbbdbnC1E
Xk9JiKu5CUM4malM8Co+ln4rFAmcKDmu2GE9/WYRNiSyyBbtfc18PeDETzluXcAj
PYUzNTfS6YhUdUu49n2Gjr6rIgN6ru5SatLKm0e6U24HGZfYBBZWv0OIZphkhgI8
RzyZNYSZtXNEpHVOM5fumYcqTH7wzrOGrCnxUK0WEedeRRAmiXorf+n2KbeVXVqW
zqsNGhkx0urvQ42RIixV3zdhMdMUc5sF7Fxze37FlPzr4RDZo82+PWj3NDtvdLyh
SUPnUoFNFMI/3wdcTUSZTRVpybv+zTJsL1tjektkGPHm6fvFKMMzncQYHxom4V4C
u6Uc/KgUaQHEaUVTrtpoL6fsfKTHxNvmruWeKJBAmP9EY3LtQpsKuPJdmqUVSUuu
6uh3QXwUlBUSmdj2GJyyWXnVoqj7jJ8vDZZUvgoMMk1bZvzCJ8WPkKXyrvSwYeGf
FBQNMxFn4VTeyBeMGTcgHwrejfPoYAEBUZoTOpKDdLFAhOHjuq+l5Pm/lQIJSO67
6QNQN6/xN1H0wzqHV2r8qgTdIW1Tq+oxvLvRb5dB3u5AtY7lDPfT1fmcB4bK+7Ci
HE1cMpZZN+ctHe7dvriS8LhH2AciLsjwgCjkfjP7PqLxDYbFYHpqsf6YXSSUzINl
wss8/m6vQV5I3/Jm+qL/2iqQTWxNK+XEuhdSPTGrfqSk0726dUhCmxJpDVnPVI3C
/ukqGh8Ht98gFIwsfcLVKCP7BwHZ4M+9WNhsGukuD51Fnz91QqMApY3UN12KfMe2
SpQmENdK9qsBvyq7eX4GeiWUUQVWzjO4vPvH64VVVj9bY4gscHiGadndsfV0k4YI
sJs2soS2nb9/D1trThVP+MixvLKBRtfBvzrzYIuMfVQzMQB6yxw81U6EB9U334gQ
lVF4NcuTJM1azBXmld9hUk62uPI/OsKniAWUAwjxIYUvIsnW5xAw4/gCFuQ48YGZ
osV2Ey0W5tjgLbp3lf1Yf4BZ5Xq8uIWwkMcTTj0p8zNCpuGCafaRZL4R2M4Gy9Yq
OQudigqYS8UVs1/j4itdnolzabks5cGTUJh4uSMLWJYUapzeMu3tL99TJB9RAwT+
CyL96/qgCrC2gXmIO+bCUTrBLo+5XRUzXc/4MzqOdru3qZQAbolOXS6AYhkJ4dqr
ikcEKWAzlWJkxA63Ege2NLu2Yk17/Dunzmjm4opHkTJZsfWvRlftAuXqMIUfgIFx
kIesOIz4sTVCsF/kTKoDK5BbM/S4ElfNOUj8sfumPWbqHa0aEeBciUDBCeu6/5j8
sJoS11zs++R/+po7xEAhCRc9fihy+IuQuwXU5PcjQyzz6GmnIZD4jZjTqKmYY2vn
cJRvnCWlCaHsUO1lNvhNRCw6CvzXwtq0+5Ob+HJuCCbejfsUCkHl+Dq+1rpM7KyG
s/6wNOODOnXOY2HCfNM1lw9npUmcrKZcEiynHobTpql8c+nOPDZQrh841gdz3elN
r50b5/CBUUQasor+PgLkgNO0XBUf5sLazgM+EKMZxfYDLsT8A54X1VrvbIBF1XNp
Mb9OhhrVaVWOrqgJfcG8t3Sq+pvdTgKZX2ua+vEjM8+IXHKIyfarKbxxHcWPbt9Q
YYPmf2GBYfLgy67gW7Fsdh070ahEXKanRChCkuG47DQtnbDwQ5CM/Qt66E287P28
cxSzQfCTOBpAcB9pkeXP7JBJ5LeKzHqE44K/g7pGFKM6JaUINsQ4Y0zv22wBD/um
ovJipNLX1kB/6MtvZ5XK5ceoGpfO3WbiW/ZyS5XMKo2u4ZYKSE96dCMzZMmPD7tt
y8/NbPnz0+O8AkYRVYetCANC0WIS7HAGPkZlH/gHYgretrLGwGCdYAhK1iqQ9vVq
gRjA5SkmyQVNAuLyS7RcNf6YwwVz8cbh6yHeQf3xh+Tv4bc5bAxbyf2u2ktHYRD6
wkYXON6qsV8Zlp3LwS03Xji0SCsvq+wWp506KMgwtpnXqHYAwKLu6TpNccWu6uLx
Jg66PEVRJsXIhNoK/CTW7PUT28ioFG7sgomxKrKROJ0D4MiKRkgzeLAv9KKDpDb3
lpvBDsFukGPKC/aP5vSGqr8hjKSUV7zw3DPBygnX0FOvCbRBu0ylKaUDIJ1ltFsb
YQEJUlcO/kbqiUaPAZdGczysakJ2yuVc/cLCnVebgbI+NWaIR9ftuF6tJLhFs29C
5bvw0qDOQQoGPlNbZxVu5mIvEFOLywO8xDl3MCw/TQwEdskAf1jGHHaxDvCKHwBn
sCD5NGwYhVwSbl86y7LVJkATH4U14jF9VuNq/3nSvrpezUh1T/XYkiYb7zXOXxh0
yfqXPk+uCxDcO68mfWXDDFAF7EUySmMfpBrC5wRAB5e7IKr0V4gaUz/5NyKJ0Ff2
21jJdoLVfG/iH/Z4w/YL9uI7EuyyHm1cEZuQ6A1Z/NfOawYAnSp74qV+ITjHv5GP
WYaFPjnHPw4KUkKJa4SeGkvIJ3w4Nv/EsDt7YqeVJe0v0U6/bvCISjRVQiLbqUnF
OlI1iiVIIyLqbhGXhJF+VrKPJbuLHtCktKS92A7mkJexJYoFp1BdwVnNgxk/rgbx
fuEhUveP0s+8ROIlB39RqbpInAIJsYTx4eeyYvlw3pxpjYsQpZbS0jxgFk1nkaQS
V8sLTnP5maJFm4xqgunb8Ta6ZDHxRXKtckPnUNFvwT1MUMrnUF1Q+mgTB/U5bqnh
sTACbFpQpx4p4/zKcG+nkJBlDwKQ7rIMohKGtHZ0stuGUxr5p8BUObOkGakxAzWI
HTGgg6cmc2s4eceIm2YUhyJ9myF4J7AMdb+VVF3q/5bOD2ScOKXUOtv1jdwfjhCf
5A11aNA7v2I4QR2tkK0oqCwYk66U7KFYWNYfzJYZbe80N6Qtekr+yHISnKDmW1l6
xbPcLJIwvsRltPxTkmNfPFvEBfEi+FfWrI3cvkN9Yc/nTKp4cgl0E5p8iBrVhC0x
Sk/uaI3m9BuZazpmZEPy+XGwHCbkGnNLaVuzUKYRm9zUbepn7qNApq9Tv9EP+1he
P5kIGsoLrjqYIF/4rPMOVBp30RkJPWajmZDS9yzNkPBJyKIWh7MXWerHn+Wpno9D
mOrcVc73arFwWmRsxtn+KCvNhOeGdNqlJBJ3XNjcOUKcbhcSigDMapdYGnBWBj4m
j+Dd54elQDKrTqyh9gopiYcHKPbCH/Ja3jd2erPts8aTHMTHaHsjcZZNYBCM22SD
YjbpVG6QrquZS85S4ttNXkxui98e33WhX9OTQ69HuCvdL+oPD/DNRwVz30UHU+CF
wXOZCYnL7lkgd0OQsNcs6u4UrJdavoqJXi5qqdIxlTVk6fkZbLc9w3F77DkFsAJZ
b8UQCtOuWf9V7fvjDE/2BgbTZdQH/z+PPrGU/ifAaVRzR2sJYPoyFANkOX8WKgYg
FYDBKv/5UrK9ZOPPJMtTiew+oSaX2Yb2F6N+YpalxgI5zO8aavW4CZkj26p1FkHs
/qJJzkryVOjYIOwVD5SEQo/3MwhlXaImncH7kAY3Sj05sQKukWPV7fYjIHhIUP56
ZbeQZRDgFyLjG+EOfNWw/+N2KfM9TYOg2Bh52DBh/9GWKbemrehNLNokVz//BruR
KvVngVTWfXQjInSu5GMY0JvBr/mBrWjXoa0xHM82g7Jt0fHfeGiRbc98TCP5GOCS
7g7c5gYLg5Rz1EqBLM/p/VdKNlQhMplRprYtHaU8KulBYceo74IT6SDVSsw235M3
AslxAkrGdeRjMomn7pXDT/sMu5zRfF9CJup8GJEoXAEd0SqImNIyse+BiQIPec20
Lg+gngGsUpcM8ZLQmmHms9tAX1bxLN+qJAVTrzPuApP8lVNLpmpD+6c3ie4qWPku
zY9tVY0fjxDZ/V/cUmigLSIC0HAj7RsQyjiiBkElOkd3PP2t6u5C381QfqMjh8q6
cj1FhHAIFmHPxx635jBcWLrqJVnO4ovWLuZ8EBIbDYiA94AP+nKkxEBStw/hsbfL
FFAbuWHKvPurbT3F41Q7QF9i/qgF5m6PufRgKBZW/rc1Ji0ukvgBQmFco4RgBNOu
NzATzUY5iEwdvKKE5z28xJN2xivyJEbBlDlrX9o11GZgXSHwVhVSuF8FSBpmRhQd
m9i1crvKR1U/aVLqqk/hJiekHuIPRJL5c01Cl/0brAH2PZVr10pz9osBmFuSftVm
UJyzf2KHcN7Yp0yycG4RKWrgQs/gESer9v+BUAQdcZsPPjfXrwaDMjWceZoZQgVm
nNEv3yLvg57om0gGz7oNKS4dEzGQi1MLoGkdSjal1u2zvmwKZ9j0DNT4XIC5oxWg
XlkkfKdJXkKSWaWzcTAFImZ8s64H/ICCVI3dKyNVg67F3JwV2LUg6fgkz4Q6aM4Q
28xDps48dtbaR8lpvRF589+PA8MdGemdDe19mxOAQ4UAU9/jwpcci5TSikvnTh2c
aXGmLavttXQLgYzrL3lgop0AhHC0fyA+XfHmDnEfIeIOAZyAj4xokFOTngcJERX1
EYRjcfNsUXpY9ORuU0j/It4RiKaHIO3cWPSD162TpW/7Y/5JYmgi4/e7apJpsu+4
1dHroVhZ8K6eNj9wYcw+r2mWgx1yw8PdIH5Te23cfegTz5hZnb2G1es35W8sVUi1
4E4u6sAo21XYzJf7vzGbLl1m6VQEAiZEwEq0DH+QAYLBOWbstsq0TFF0PfxCNPrj
O7uhvKpfThCDaXlwTiEXhTH5qo2k8zCWSJtRfvBCHZKOunc3vBzhf4uMzoDUOnbQ
cJycdSZ4Yywl6GWUS8+skjxvc/6spFjr9NGHqyCQeqsXt6zaJjC7z1dhOnFK1G95
GxYtVyHfBPRC/b5N312I2VE4pZrstyfcBnaxFXirr8dSnTWwZHi7u7EZe/nBOsYM
lBo/LMNu4XstDdLIDekaVAGvKq74YSAE+f1lDUcckXJxNEItIJtp9a0cyc9E7Ms5
xLb5XHqlNT2Sl61Dnz/ca5k5F13dF1vVfVx9IU01a1J8xb/ZNz7ALvqh9Sc9vJMW
ApCrucQSqWMxAWh5cdX1ZQzz7uLVxus9r/9BWGTgLoN2pJqMgUTvDgCFlxyw12eV
SxO8LLx8C6H/di/WGcaSDIZR9CuWIKflzmLlFgnJcBNnjZ0XK8S82IHSmbLqTPhS
ZJ0NRzMO/GE99AmrRlMBxNKixKPA8LrvDDRzm1brgO92342Ck/olrmND9vGBdTYt
LpWFiywdD4qUTPdymZ8aEmRsg1zH9B5qHp8Bq4NzZ/9WPGWqEhtrGo9323y9KnDi
mkH+zLIJTWaTr/Itz+GPeUara/1O/QvaWeNhzA73oQZLV4UOJGURJhDH/SlqeK4y
/9L++RNKBAkG1pDmgDsJHJlq1BtzsRqhW+83jOzE/68UPVfPGojYdx4yWD2+B99F
5ggi8MDQq66JDrtinWmoQiaQ0MyHWk7TFozDbikL8kCuhzsxZdQqqh4GIgM9P/+o
AW3r0sLr7ot+4H4sW4Zz7dE/LoR2ROjo2DtypHVItB/IXr1OkExndzMPkDqpUiuT
fkQ9cgBfRVvoro8Jc5lTN+cH8HiJE6rO9x34cYxTwZ4ue7jY+WsarImyrA+F5rne
mWUSPl3rpsjcuAVeFYHGymTUlXsu3+nbCZpX9OJXwyeAYAyrSGRmbGMKfID5zqtn
Qj7ciiycQWfXxVuvUEn4p616ksgKqs0MVpxHrX1Zm8j3Gt/8TODYysUYnG/7C8GQ
M7/BIQM8B48fHSzW5CS7qI6ZHuUB+N/NoC1d6PK5bWRzognqNR8KvzGNH8pRgH1Q
goYwFTLQpwV/uebKTXqEL3a3qICPgq6sZqasVK5oRS9sjW03CaKErTYANLKdGWF1
M4kN8CD+c3t0wy+hGNdnYh8RI1MWxn7941os24cHyuyVwgi7ToyckIgkdqk9jFtD
qspzXXjlMmgwxuCpxAo+manct/72rsGOYW5XdCtUjgQkcCcqmd9rHsesPqrHOcGh
qmxtFkUWgws2okF5ldb2mgtpKQBnN1Al3BsouX5ydn8qMdX2GttfK7W3spxBFwYR
JPHRrcSK7vyJ6jpEdnhlrkl6yxULlsRw+cczA7PYdSPHbb1zh7q+LJo1pOBk4Hfx
/sNiyuVr6vsdXx9u2Usnd2gdovVv/TtABP7AtdWJyNRTG42TLhybnx+hkPM1cCAK
hgHXCbToGE5H26yTf1Q0PwuSCFVUlmn6zl2DnQ0pj3hvIci1AKTTDSeTOZyl/HuA
0SqRC4XXgpu8XX99OjwACx06KXLAp2GWRVtlI7JByLLKgRHOdsjLrB0v0KivqC4N
a7uh1H2lWrKg4A7LX9Rqo1v4/0dZw+akAsZhryrwmt4B7rNMOldTQGDcuhW6jD8s
dngqbaYwacNEqOV+AkMYJYyC8piYD9Xw3V6JFkKhpHAhG1xWlT1wmyNZN7U4G/TA
c9QwGezMKyC7BEL227EQ54JGjjmsUHLpUZEhfd7jufv7GqN+PRmQhvXOr9pxcfVp
U4FyUPp84OHtPUIkgf4+4skPQWUtl3Hf6b230E5dv2lcfosmTl96rKT0gU1W8zSf
EcbKPRISK8fHk/Nk/q4Xf+Odq8JoIIQxXnqm92s718bcyUjFRmB2oca4Rxk+dLOD
GY68T2dT63jbbb+L7CEXLPpaqJ7GrE72HFtyPTHYAs9dBFDHLfGXCF1ERlY2ViMl
6Ewn0HWOw8iAlAfhlGdnP8uhf+ZYkU8z04r0zsrvkAiJrE11oxzNoCUUFPb1qE3k
G44Yhowy3J7S18RKI9KxBk21XYSd5J882I2M+9dERVAAt8g6fNtKuosDF6H33YKb
JawQOsBWk5fP/eDA3VKsZ9zDAN0sAIXkBDf554J/MGEhmqq6m5NlZCnMG0ZcVdFm
mAGimIQIXOEUuAsCbKkFcVHDojFDk/ozUjOFZw8pD9IYho6Nt9z3kOKyEEcwXDBB
Wu8bpVCzfABjxpa6FnrNmTwu+sP4lznKsgyO100nL1nLvkIqkEGdiiLt45fI+Cr9
NEP2OwnDG/wsG8ogENl23NYisQvMPFcXYbT53EPiPRgqqeQHtZW2+O1JxaqsiFgz
1vtt+pCZ+PYoliOel2sEEMpWVMSn0L0T7TkueJ1r+D3fAOj5qb1fA3WwDWYHfSC3
yW3vTaD9j4Jv4YIr0Y4MrQyKzIi9CehMqwVWJMc0hKr32FpSwMcIrxalr9sUZgSl
Jbk9yQFTrU2TNFN6Q7nYeb4q/LLNLFuwdDi2MCC35wbu8sYqCxlEHOnITz5cPoL8
s0LH6pJlrjmw85OLCR3LEO14RnNbPLGgoOT6eIM0NM1Kz5fc4YfJKG+31diJ4/j4
teImhdi2ih/MAE1651D6HKe6QGdsSPngF0JT1bGthEyaQbREkxsptKEOQm25qr2I
1Z2hyqASNjrYR0MRWTZLLM2Z1FsUd34hY8yqOO5XtsiT+8Ozzc2Wyh0jAW/Mx/V1
We23T40fkyGjnEOybW0Mlz7DHvpkqkCMaNmXmmOncmjtTh4VgCuqpW8feSGq1f1+
O5V2Su8uUb0274Bjfrp/NsY7Q3ben4JnpEmJCg+mAq3G4GyKa4ukSgHqVE3qnHwo
Fn029q5zmhchz+exztnF0HCUzrn0MbMQ1tARhTwE5AiIARy2g8sLC6JNEQG+qrEO
wS4K/02HUL/lbDxuk1xznKpgs51dPdki2/+ydJmuuLeprOn2w7Yo4gGJA7HZQ4oy
BiExlkU2Mur6e26Xvcc+H08FLricpcC1Wt1GE+ft9IUch/fxnkLLgU5bqNPkE0q6
MJDshij+lATk6CsCWaRvTd9w51ESF5UclPDtfQgA242aZpEnkkwb6SMB2blkZQPw
LNiM9J+3EuG8T/mmkvoT1CTq0Fq+soLSx4lfqH3Gqcvtg9sBylin49hDpuANXds1
Ff4DWEvxx8iMCf6J+61iNj3qkVWhpVl1dS2qmA36JQI9yJ505ydaerYh6RD1pm71
lVdzB8n+2+g3sHTaUqJcVHWiY95MbfNhLTugJz48AzMCxCtA4jm2DfMnFs7gkh9f
6aree3bdkbdx5qfJLUvkUiE1QKvndTeMql8E3tfU9edtaWTGBYsJTciknP7MP5wr
CQ5bzk0mLRwrNtbLaoKmY5v1+q6P/+K6qVMHlHHJvgYNA+YlLDP/WoBkTlWDNVv1
wwfDm8REjp9CWXAKYTt3LyH4ftxo+MtTq0JuzM/iyxiupod/fDzkI/DKqKLHdWB1
pVjztlIyl0kg4v0RAc8wFF6jbWnB9FZo/bKm+LWIYSZq2itDRwQ94NAcDT647Fmb
ymTHWg0ClaFxf12EjOGmyh70eMqrVEgftfKoR3m+9i2cUiw964jWht9INKwZKuR6
SPTlpx5jRxddpQqGMtyXJNaOlSBTgsJUqVGa5uMiyFEq6USnvcz0RyJ0xESlCWhZ
xMoVV0n125wzsJShDkfQ0DsC8wArqYmY1kTWOUhoNzCYWd1Rr7UIy7vNMZqoy2LH
Fjt+HMztyt+AM708L37tuQ+24dB6l1cMe70w9TEtOTL2AE8W98X/zisO9oDtNS18
4BMilfytYNRGE0WGAAAv9LfWh1FMCO/P8Day0rsaiZbwB8u7vWBxRJUSFuLjwfqw
MFV0eD/R0Ly529Oaw2znWxLwo3Gwq/5QyKjgoGYOwH+R2P41XCYi26anlHLXi/27
5KXH0V3svrdshgHrplPOgAMvs3HaKR9oRf+yoWME3LMHmFL43B8IJnOW5jikmDSI
TbQOlW9BLaa6NEx6nv+6UwYpTjjVO/eqquJAjSvTUC+dPJ8z57qgeOBCByAqG6lS
HovMCdqC7Gik/cJ4WOj0u4LxOqHqXpQNnflJKn7c3JdhrUw0cdK4hwt11Caq5XOM
5AgbLyw+/FF4DyIEtbrf+w8mvDbJnso856ECfq/RnzufxtDmyAaxevT/ghTcb9Hz
vOvqO+GaKxepsd/TD4XUl8mHdJoEQCN6/HTgElAFxR6tfmGsz3KD7dElIx6Oemt6
wYt08T9x2nRm/yd6QoHWXtv+dAXjkfBOJXUNhBaVptm8tcFS5q4Y6PF8HAInUFoA
VrMOgFwUGsEavdBFHehPTLxx4WS5eBxC4/1nbimxh9Cd8e8J5Ld/gm8oX4Tw6wSR
CDyXfg7Zay3uGNMFvFTqCEa436KhCiY7LBwz4k0BChXAl9gmaE5JMeFFoJklLoyq
1u7RfNwutRk23nhx3N9Ciw0ycqq+vXyNRvUXRCcnvRMISZGcrjfkg4YetKCVh/Nb
GsH/lQRmbiF0029KvQ3i89Gf7QRB5QcsdZibD7YcZLxjZ6fV1S3jz6YSsCJPnEkl
nRx3A3WRrpdP+EUAqUeMn8XtHBONn2X+jftftrNXnSciTJgfw0TyJm8+l7U1BUk1
y6jCX1r9g5TJCwWlb2KhLNcf/376pXBZyBwU8b+sAu+R8Gx6t7yHOhJQecwWx3Cm
0LGE/l8LmPGBU0LEDeGgI64SyaQ9gGTYDDQ1nG3Z1PV8HmJ8L86iwZ6PQbfwR2wl
W849jhtX0nm7yEcgVUR4kKPjTw1EvILXmvdHzSZZd9blVJCcbpeoiDeW+6VZoaGi
fd/ecDm1pRNMw5LuESlut6k8/EyhdrJmrGFCHUYQ79oApkOMWQD/H63qYVyTpqjV
p6PpK7DTJrW/dJI9+BlhzixmabJnMzmgK58ZMPbAxNkUcDvb47eFcCPZ4b2LjoVI
aDzQgyFTPS+jfn2+PX7KBSyU811XBZkfFm6S3Ya+wJSS9d8GKi41B37zkqpHTO0t
UIG22GmFknfOgNTxntYZwFYYZ+w3091gC7xf4htj/jG0BYec1jh19OEoEy1IrI8d
0xsOENeHCztCPpDDCM+tw0nJAECuBilDEw2Auk/raXJWwiA7/ELBM+5ZMpoewT5I
/TLcnPl8q/921LEjKeuOdQAU6d09Jicm2XL+alx4/6nBFMLxeBRj4Wjoogt31ioO
gtbqFR4GqTHvG6kw7Fafk+PCzyxERuBPbIzH7MiAxUx73tJbrD5FGCWVYtVCZI0u
F8sEc+F/zKN2cH8xLJx1T2U4MpPHV75K4FGPSzgep4I2V6ecaZlw3vSH5nUOmUcc
W9GaUndg9udw46reZVm6OXKBuwhRvBoQvJrSap292/zDzCyphQbZotmjUs93ooEP
6gayacCe60gBgsk7dhFSLKW7gsduMIo/vR5eUxG4NIIqnX1mLwL1LPIawPinNsAe
c9cyKM9qGNqbnpLa3y4BQ5dgmWt/wRMjTj3Diz3BON1YbNVuZT0BkEvY2Fp0HhUs
ZPcvFPbYqvknb/c/og6XS168IzzG6DkFRQKd0ma4VPjPZ/49+aeJy7Iq4+hsv7HH
dM+grXSfR0DsyHc8HisyH2GVyVr1VJSfegqGnn7AKD6iCB8Q0wDMGnBWGi3dtw/z
4uKBNZ2kLTWJEN9Si3+Yc9GhEuiMEGDi91cMeCMUpj4aJGCvbm3AhsDFg/xkvNLy
hapczb/gXs/47wkjiNyg/Sw8MMoUd9UmvqQ5Q02MvqyBH49doUl/MV6Wxq5TWTiK
GWV1hn9LZdmB3n2RMmfFZ6qud6sJoLILTG/A4KFRCbJI7BKMyFG85wbd9oY7MjAv
jy++fXdom2B0a2aEjc7FyWudm37xQyVPlTq7WtMHZ5KNcHWZS9WTNEG+rk3Gv5Ho
JcAFVETgOxgkiWJwdReWT7SLrWNDiDHwf11LCXGjs42yXLIwW5PYEP0g1plcOjjq
rZXMdRKFAhpM1Qnt8IGQvz9gOrUUfXY21Hsi73rCm3s815xcs6//bNRZoYuWDmDz
4a+AtDwUaEknE+rfDrsfZYCjkep/dYLffpGrOuVinbgutaBjhOljvIe78ncUMBus
6nB5DfnnKGderDWjQIvnVe1nl18kTN4JZmhLU3jbOAWL5xcSI4FDaMNE0TH3sO+A
cISvyjQdA/IzqSFqDZPXAX4+nkHjYAbj3KtvMrGEwprCSRhzeXfNDxt831YIwvEW
mjrdbxtiYYy7MXdfX9uxIkUa20mE3MqNIMVEJI8VImgw7THygkFYxOry+mWFFIN1
9479m61+2AAILmJVyb52nef2xbxs1Rj8lS/5zKDTIcWRyHUkeN61xa77hi3pWU3n
YXg/hDr4nh0LacjmZu8YDtxdu+Bz75sF1lGhUKW4K5OcN45wVhy3+pP8hlYuSlCl
iVWrKiy1bQsBO9vk0sFJunrst3HIfEtTYAwUCeD+t8j7b4zLNR0CCvYEyKLMAECp
iZLbLbtUUvlak2TglGu/oy9n52Vm3u3r/NHhlNjnDGyideaOymHBTIck8UjVlLtB
5ou9wipg4L90pQeoh9vv9DOwm7zs+G9TNRlfT6A5CXDNLfiRqYnTBw2XNhm4D6n7
89vUrDfVhpLCZW08QQUZP1uUN30sSFVeWaMTIygtP6YNKV7K2+ehrfdEzXTZhIf3
pmFdlQMYhnJa23UsPR4lPr0VHaeaZffk73raGwlMWrZYqYBnRoJEaltFdnOg6/qR
JaHabe1QlprZuqBn8iSDcFjduAfEOcZYfIoUDpKUqCMrIjRIiVb0xaJkUL9JgWKu
i0tNiyyzZKrjjzptHWo60JUNINsK2x8rPktD9nxx8dB9ooXeJMAvLtXO+y3QkhG1
SHxTOvYREozTcsqO8T4cO6H0HzX6XNA83jkeuHPAVKwGOAiR+MN6h6F8yi+dTDNU
eYyb1T5xZSGQRA1tWbPGyH8nYxbzSAY17br9+C7rABEz8lIGDhqGh/X3kTxV3lug
jig25FDSxTLn6QIkyNZwrd6hq8cMRd6pyL/540tQ8thE2HSJ6YZnNfHHIyseIxkh
mg6xLxjUklpxJa9d9xIU+cheSRJUCF4JOG+VNViBIFUAUDoo1WW567qTeh9UIqH5
RmLsdduJwdblqb9MbSPxZS+p3iFR9mr+z+SeoUXyVRFM67oOmKQqcCYNugaSKq5z
lj7rNivAgqwUh9je56Y9wA2D9vYb7K/NCfg+idBREdLZBe4DlyykTIwYMaOVXNWJ
ubDFgN3zdCBoYPbMCNdQ1kDYorizXkedLIQ4MmCsbuE/W8AH4tmLdlSwvs4A5Q+k
E++hkEcHdOfZ/2ldIcBfSCxlRxgskc/scsVmLSpVNPI/6SElzqIVX7M6HuP5X32y
c1sEKTYidnDIo1IFF3TsKG884L97/NtEVEXGkDVI+37S06dXR4dq1bmwklMLxGm4
HwY6Latuf08r12ZmSXuXQLV6qNflqX3aDzcn0h2/8mRs2pJpnCkxIP8b6EADOv1L
xX1Npk9c2uQk6GZCFRmo0H28bFfRINuaCeJZRqA89KW3b3lEZG3fK6CIrS2Y645f
N3PrxrTJDZhFnfa8wscUbMoE+CcQ/00QOFzMdBKt8+Z5b9abLDpIyUeSOajTDfER
IqwBhOqQgDwEPVY5/LvpFb/PuveD4iz9N/In7VHVyMbZiDVvLa/7vO1DOhHy2eFP
ehGF5zH4Cq/vqzhN14RvzYcdp2qzdZb5g0gjuysCfjTQ2Bvc0LhbYW6IKPr1xhSD
3Iv+l6sVd3OVMDXdxBO6IKVUW/zN4k1zD8KWeNF9OTfefXp2IYLKQQtLPgJ6/c/v
yaXt5tHjqcBS4T3mcu/KPZFZUyWIoVT/lEmCB5ei4e3VB3wc0LTaGUNrEo3aLkw5
1fk5ewPMVKLKFG9IeJHP90D3I0Zd23irxne/JyvTx5Y6kKegSeXdpe0LICLhG2gp
f2/DDcoNKI4VrDOPjMgOnXi2O+28cHKctbuqWfx4R7t+GRU6MuXxiABjLwCvkNPI
ViBwiMfcZIvW8ILxwL3zZSmq0Qu+jl3s+4/SdG6/1X08MBZTR0wmtcL3uvlizpvD
8p/AZa7N9JtVrxnu3jZF66KJ4ytzKIv0kGvwoAuyrWXy2qvTWh14CfPfjvsZHtEl
UgiIN7gI2tGT4t6Mhgar7celvxLB2AbM684vYnPYxCvKaDyK/QSqs3fGDTx6MlEA
EGetQtAiUhfgp8gDH+fk5ndsG8yu6+EyRCDywKx7UzRYcouWMdv8dHqbsHv3JmWC
GtMVHnAvvy+VIozwDc38Vmjv0F6C/VEsuaCQlckBCUskReWhpBvHWiYA9gv8kOzd
YvjEeqgtXIeX7WRsCQYxCZyDCz0hkxF5gQRa5hk4u+43w08LhNuDaxbQLcyqtC9n
P6mBE+KWvs7EdS/7PEjSAX620LtFi1VNvXqfQtaDWe7iNiUANXyXDiZXYmPPXk+S
4bCyCR1yqrnwC2ExISUJxOQ/fVBsf8i4z+Z0uIjbFV9RR6Hv5xR6DUGe7HRQmlHm
4R3mvlRl8KgnFcF1qKeZvwfL5yynCP5n7WmP0hcHAtEoOrHwphIHZ1FY1PscIpks
McrE04l6sbliM9XBQo9AFHo2mhcynIW2L+ceH17baGUB3LuZalDnTnL3Uq9UhXyt
CWjJRnympnRtHFf7rBuIIWoh7XZ1LQqRTECseJxqWV+e8A4R29/gxquM8lKUnX0j
5LytDrllUxp1bjZE7OAh9SIwXyH4fpYthfYx7I8k2IjBmxgcrJ4/q6e72mpvnBDk
Db4ulQL7HYKMTamBjWSYBijSyJVJNUVkevTTFW+J1BF/8DccDiFqo8xAUF6VfUus
s8+UVTuSbU1ntE9A+7LHseW7d3PJ3VAyj1yy9KyE3QbTdQFMcAi3M+6SoJVTnofk
JhEwJV/2ZGlKjlo47uJ/Ge8ARjhQkLdoIkktj8kx1JBop12fNUqopoFzQwP5Vy2J
YBiv+GJtUR0OZRQ8HH9kYW9BGaEnaSgIShh9u8luk5beiUCV2HhD07ZNLLT1/Ju7
TYlMVYbnCG3tqjwReNC35UXkBF/ETAiiY6yIT5+rwIba36S1tYfAQf4m2KgdWSoX
SirZtBsr0zu6vJULVXwDI6XLhGtftANIyP4LYLKLoAvBVD92qTfFwfxORyYhDvuq
l3elM+vGqp3adzF4AJV/Xh/lpdpD3Iwo9XqDJ75gC0iFf09GBTAbqQ4UTo+FyPRQ
f9w52l9wyqpgrMOmGQNkwT3v4YyCtRchzIhQLlHTxE4IiEjamAvCX6KU9W8ZPyxe
PQw8vHEqY1OZ/5QY2ir/vuNTkDEnoRvGV89w1Oh8gh0IFlGJ39yQ2J+C09LRO4et
V0K5ryVg6FQXv/FDl7ixgOCISFLoNHbYGlP6sipYbd3mqNyyhw55SvzfZh53cWrd
awWU0eGbHopiTQaxhNpiT7nSCXVLghrJhFeBwO/M2iGa+hnt49JfZ0DMaUV2NMUc
X6SpgXfXO87oVv+7AlQXA7zktXtdS/2bKJhLb8M9sSMdpNNr6AyZzjKMwWBCqppB
tszwb9A2+AhbFOOggaSW9pLyB/D/3cBUv6h4eqLVwOzj6dm+vM0jefADfqVhWym/
ddsbkFqKmOUmz+pegtMWx/uvRQiopZ/bbYc0H0aSFEBDuHG9vXfqYl9OHbc/APOD
B1CyznDEq4lnpvLuXf+8f4dJjV9Lao6czgPEnLD3VWjzAhLXtTAE51G16F+GxPRB
0jV7Nh4pEIAHrb+1OI8Q5qNH4zYrTuUiJJVhfqwdZLyUS1ooLQg8YRKG0LHhyFyh
+7iMVpp/tLmJCSrAl1oZsJiN51xF8v5iMajJrdiCBFvsAjxbI5T0aVSSOa0A77To
2E4Wk2+/fpUPieAOv/PpW1GaLDCyDFTPgf8JUQYY7uX60F0/7fBhYKxIYtLI/0iG
0gWjytmnjMKdyC0/ruAbdtqj93B9DWflPZtn7zemQZ1aYzm3uev+i46W/wPLsYjy
UdVS0B95VCrT2XYrFoPynV8nXBpd+ozpO76W2ckk3JryZAmay0fw5pqdNccT2SDg
GHwaeh9TCnvrF2QZS1S8TRwK3fn0pQx1Rmrt+9a5MgNlB/5CuTG6t7u3RiEWB7WL
JFCBStd242NdC3+RggTC505HFO2r81qyzqhtcG3huddeI7zK0RKsdkG5i+kAvVaE
ONwLnGb7bAXfMACnrSXbOBA7IkZT6uvFuM/1/4ctNBJRVYLT9B8NE0AURYP8Aogq
qnSIONWBiSIBrKxgHo3mRUDRFaynypt4XH2xtm6aVZO1h4PWpTSFtqLJ5FFHnHL0
tZd+VyA5Uz2DSHKi7MpGosNxCOahEV8MrLg5rvIRoEaMzXQYVHMdCbD3WulsNUlo
/AbQmoLkmVBOcQvy8JHUQCe5f6V5nICib2E/ma2/9DamZX8K58xzSXwe9d0MVT7y
b/jNWMWvIkD7BjTTkkUtuROxwgsFClHTOX3gxBwB7PHp8/eXDj5hM/Rjq/pKkVKZ
ob/HVQghW0djj/IhNJH1PlFHmthU5ChS8JDKEQW4CXza/f+Fgf2rBa0T6ELZnl3n
fP38YqXuQ/9s1CItfQHGNcKjiw8KAnkd1+Ogw/qtVre3gb78RkK61dZB0L/hjsG4
ATC0oMUjeytbl26M5eeLAiACRp0XD9y/8SKDlCNyhfz9FtjrpNtIFuG26Cou0uxG
P8YSruzzxLJUjkgXmqqE/sRXo6t3S2cPTria8YEgpOny1IqNj0/91/oYQ3qBSeiW
Ra+Bhd33MnRg20TeikUuFN6ClTGjxmH/HNzOnATZxJYPuVBVlV4IsJnYENIN5MyU
H5A4Hw6sRCTRol9qdXk9TINp/UaGGLsT8QYJu+yPOGhpiNi8ypVFCyZ5i7gRpVgw
frXwAe3d28dahe8qPJit66Dgv7ythzhNTQsHDB+2tYc/ZrrLErBCACFtYa2uyAyB
1xEQLOXoP60FJfbGhQDfIc4xym1E8aWlGyfHD+6/OtlcrE925toIFYPGWrjV3T3m
TNV+fqQ7x/ICUWgr4XOkNMGwrmH7rWbkrZMLlVnzgOZP00Pf8gQNqxWFt80/LMRU
0MIHjVRGOdbncp3MxbBUVyNBRUe9YY8nOH8SONuxh2EPfHoN0V82FBY2E9BQmbrb
5eOl+QjN2Z+02ywy+Sr4o9eHtWpgNE7AEpP2dzVusaH4pa96qWcNp9o4u6IiAV5c
OcOkG6lZvlLFTX8B4MjaOxXxiuLP8T4Jckcr5stZjlW8wm9NIqdX3BDiOcBSDYok
W83c7R7JyjCPokvxt/3MM3G/kxSmqupMOHlnDWTJVi774mbmVGqWO0iNqyyLzHd4
+Lv5KCA4nTgTklY72tAOHSr+D96s8YypxYskJXBPC21SbQlK4q/1KixIFV76v8Ic
dEjaWH4OoMTgTpZnZW3eB8mUVhyENi0tHzejwVSC7TGscZs73xe/EQyk4py7dW8f
M1C19FsqTas2RYPJFHqVuY7cgvaJz/c6mvLWDA+pkCa0TJxfnOb42H2/XpUat8KH
5UtJOsOOiVxYf8ClFdoU575K5XGVOxTrhfErkWWLDmB9QIosUJeTlmmuAZBXYvPR
tz6nJsZGNDDrYXr+4r+ONX4G8ooXQczltwfrY6xoYuWSNaI0rWj/TVqEkGMa0wAC
RYD4ITP+7KnnAWi31BgkP42HUy9CtfT5NvTK33XOSSHf8VOFUmeShtzhb3gJDAtt
HvbEGolRAQONbuEM2/CqhugxskwYBAMZO8e4tOblu5JGi4tox7YaRdn4IvZygG8k
8myJlU9nERfFysdEmXDFZk+MU+L7/KA367pRJFY2oCz6ateR//OOa2I5BhMqIsI8
13DysCn77YWW3rb9tiK1lGBi0Ge51yjlzVkleE1HPOas+CBDc5FdztpHq8NEMUMX
rvb4uuss0CgxA2ct+uKRyVVatSdG+1ZqGB9Gw9Rc/d73YwAAyl3SMJsuvbaWh7rC
wiXMMe2Q79IVTWLRC+E57h5uhU70nhIVCaoZc6FKSusjVmuoXE8UO3oGQ2K50DHx
zLYruUgzsMpvhAg3cg7WPZPDGlJ8DdNb+uILyWPSmXxKVzkNju/1AvQ17DsiBMzH
hV1ETn8yG/SRXnwE9xA7pYRvC3aHff23wqkDsm8twDtkSVFjDdyFxckm01UpSxb0
SaILSFuORFLlhK9b6KpHenNhhf4K5FBJOml6oWGXE9W9Htu+DHHUZZUiMS6rJeOk
TjU+2o63aRQpCzwS2NjHxsFwpnnk7v9S5FM9TPcC5yZa7BvmW2vUd1uHmcPBqvXk
S+U8qG5M1Hi/c/agl5L4fxeZgFOABhZsgscziBKSvQDCalt7+GLKrpKijaMR74ev
YdMFYe4yN/G9/cKzn1+zabVyKv2KW4slgF4LRsT5mlKItKzGBiMeD8Xl8XNF60Ll
bA69ONMBzdNjRf1wa6qTiLpBNle6NzqUWkcdSgR+Ylgpg4rKV1FTMyusCbIfyPMm
iIlB3IgJM2CuZ8j4pDmFBDV5iSDl4vrqv+qDZ4bj7JCk1uADtQSqNGnOBpNi3rcN
6eSu77pj8oK1gG5RyDwl6f3iw6bEWoqcklUgQGvAzz1XLf1hDYYVskwH9rl/i8k+
O2mr7xH0moRLMf2IXIZK0wJKFWvafOO1OERgumcFd955ztQSHFXNGpomOH35tbV5
XlJiCwHwYTS4OeVdAzjYa3ljzhhhJ+k9xr6gMdtaIRe45aezXieUI+nZYN6shJMG
C2MDFog+38tSmhuluXM7X6zKPkAmizofLv/55AAvwNlNCfEOgn7NIPPC+HN/NNNt
++6PMLxBf+JIQa9BiYgnL6wBDByO0sGxUAX9IrDDqkLecfvdLiCnZopeHQsG3uuR
5T0MkT7noPJk0ZkjWXWUYydCbUBOz7o3gnQnw4vfOTIv33oCx6v48v/SxYQmKi67
A8AaBVINBX7jocQBgptKTq9T2NWheXkFNMxJVuz4V2Eo1V4QqOyJZBQZiwcjLwa6
kjUrb4W/5XSOwtHZz+j8Md9B8pLvhNWqxDV+lyZygCVw4DgzaMDrEN3/6nKQu5X1
NoJkUU0iRUGzzMSD7IaNjOftNHEVj7xtCAaQuiGTqIG+bCSZyxpPJt2bsmU0XWt4
VKHYvUB5eUReustHgCIkScrAELeEW0gsD0e/58hdmbHjhp1mLWg7LTDTI2YD/YkS
qjVJoVvu3HD2BjfVSwlYQwDPqEerolCliixPmcqhIMWUA6X71OpxSEJRRX2nAwR0
ONPZcYv600CoYd3VQI8JxP1FgVJugNDVsxGhLsnncxZpE2ofz0ahVKRknOdZAbm6
N86tzUxTBpn+RrsHvUWW1k1emHR07ylzzMXamWqba/jfm06zwwB5ivltgGRFRnA4
XMHj4SsGG0BGCZP0GlUvjzL6DQdmIL/CPIjCVBCuYL/4l0jQaaIalCoqtl7wY84F
RM/CKRYI56XvX5m2hjf5WQBErWXVdm6vVPb2B49T4/upxI+9YikIPmNyI6eH+k60
Viizjg9lLotrqlSP2T5xdT5GCOctkRwA450wh1jgz4dIvtCRbAiy89NNjCVbp1+A
HkLXkXQdSQ0sStV6D62r9ucMLIZyTkTk6l0aVk/rWJS6ITXmhlW9RoEBz/5cxS7D
EscElSkE/HNL6yIRgZJyO80w9Ui1tq2bhsOqm2bpcZNL1RTcyoeQ6EfPKAw5jvRX
bUKb6CNOFM7mgH2HGQtXyZqivUYGxNSPFc3jaoNpa0TBNXcM7rQXni400XTM+Vi7
9n9GJOtUpUP8vLCsUhERYoAx4Q3+kcec9tdVcYBvx9cZomepN2yAh3X39EfdG3Od
nmsEiqHUTkYpaIlmGwOJkdzpIKHoOAeJCAVAJ38qYSpaBqlr8lMiHwGDgyxkNzCK
Y5ea8gHNThWklwRz+U1aN2ks1zBTtPVhExJtsYMH2KhyiTdPyocsLv0Nb14c3Yzk
PetYxfqRYwpZFXDnIkugDFu1eDYjZzKUY7pZBz7aiF/Dn1wueS8X1/+D71u7ewDp
O5vABoLp98J3Fzv2I/bJQjCWAQr+90qN+oNwovett5eKK+EZkI9CaZRYe3odgevW
gytm/sNpmH+dLxhjaIVz6qbWN5SM9MvwBGhVBEASzQL9dr1v9Nl3gv4JHq3xnlhw
Fst69e+Q6Ez/OSKL4cKCzrIKwbOjsvh4S1OuqAKDAqrDW2unZDC2XZeU7hf0VQNx
KpobqKr4EtQlwkzinPnPnRIfiEZiSaZh7QrujNWOxK+qUC+HJS49KCDpF2kbdSPr
/Hx9cMoKAqJfkwmzYnVF1Am1hT3ZGkbPWMGG5XNltyJYi7G+W4g9JL6IbtEnv11E
5iKPuJpYxUZau7a5xrZyANSiDxxpBf8VGcd3H+RLU5pAX1RnIGOm8T6f3tYgqE/J
haKtHha46KZAAwLQxrbmSLZd82YmTkpEmt0T6U81XK+GDRGJjW/x4xRv0jFt7ZP8
e6Ha+qpQz+xuAQBP1d1XP8nO2aRBaGwi5EvIcvfWxmCV9OOr6phpCDXCfvgUNLZP
tHw5Vn009Ults9WmLR69aI4K2d5bDLD4rB24uociIyV8x6MZ4/Zxr53M1pTW5eK2
ppJGCgW7ZPA41tMERSevI2BPFSMkYwxYLNeUkvlWQsKzLTMMBeZI8H5oB9Yo4DMb
fbZn/KjLPivob1aWrmRQZYVrpTnX9MjDrz+unbYgy2EteWh3M/JzkwPc3FjsIyx0
G3857cZzE/e4sTNCl7+Tuz9nJRQ4j83I2/QiAkO/NKx07S0kuIi6PPaP7oNXoI5O
ghyvWRF+oAP7dEhyOhVsLV+qjjtApjxdijQ9+bHeBNHpoaiu7TMsqb9vau/GSYSt
yu0s1BP9/vmMTykkT9BlGsQDL7JjUm+EeXBhH/Epbm6erTADrYY0bm682NvP7nl0
Zfes841LYjAGHADbAq1sFEOwDjECPsXMWpWvO4e84kBKJhaDBX9Po5OAvGumbIQw
faHIMQGDD+k5ZEVH4zdvJTdJ2yu69nQEN1N12dx8fcb12wGYcoDZIhi9ZY6V3PVL
SLsCAEni2OCDIv+RNCPQy4GKAvTT36eNbwdrGzM64PmcU7YNkBDlx1GfSrYwY67a
/EO108zRsXAQEa+b4dJweMTPUfjts7oetTBeNIfJdNvFHRgFwB21FYeh5tH4Ycw0
MB0YINvor4Lk6JPPkDP2a4sy7jvO+L92DrMqMCxvrWHFAPPPZTpTmA9NKqVHtqTY
ujk/0cPyewqN6GAIiUre3DRkxPPmGyx8oErqJXLpnmODJvvdMBhvp00R2BCAobC9
3Re4L0OiogJB9t0R0q+3qnv5RRxklldP19rtRrvjFoXzCthzJWZ2Iygg8zmUYiAF
hNl3khNiGi7VRVtFXZ2uxQXyZtHlecLXNtpAhfRn5oJtdvwhRK3IjNE+NOAc+j7P
YIEW5q7kHb0qoVrwIy9SjgS5kdxSZrvXC1qPmxoiasywo0wue86GzpyKF6l7Z7Qa
PdKIhk324vwmcwzGRZ2anHSYzozPADKCH+PkUCbzIE3V3xdZDS5MwIhW8Chv/1Wn
wCY8i/2T1AkMeUBQd0gPaAQQFUxcQx8vX2SOlmIYJw14OniCIZODMSYkUWvlNkFx
nKk3V8ogqvd9jWg/TrTtHX+u13C8+gth/MZtamlEU7GoRmMBFkSREaE+dxoZF2ZC
2li5IORrU3vlTrQS/RuE1vllBVfrsb0QUCTeU/j2ZFdJPZOPSAut2tZ37OqXCeSL
PCQdUd1SApHC3ix0CMLsCHhX8y2ipF9rHEe5rn0Fdf8aHQPYxGuz6ghElcOcI2k6
51N064DH0FtkeWW/OICko1LgrYHf3NQAQSvgZc+OWYhvcJupF/w+MpxQinQFva6+
dg8MXbuyFnfRiRBrK1Er10PFmshDNfwmQem7UeYWK0FqLA8xEkVd/jx0mKBio7ca
ufj3avi5LOsE98G3CJqDwHIcXKwMMJsxLHpLj5IGkuoAWbeUHzajVT/oDENYAmNZ
RO3Zs+A2WJIOtAGI2t5YUXN5nOJLS/QfvZNDWJJtmHuVjMoWsYHrwpnpcycoUA7N
nuJg+I0X+SJgxKSTzxwDLzIird9FTzvM1d7F1WhFR7WFiQD8aoyJfSCKMR4cOYMY
kVg4bDe+xDf3uhCKr2+Kyx1Mn5E4+eyAzRO0R/795YU7UM0AlOM++0sTlko+S5lp
6z6sh+gJM4R71GPV+JHNGLqh8bewH/Uldsp4BMe55ncEfAx+/5CWAEIb07FsNuAF
gn1f1wXmEeZr1Zcj/SwsNAziE2PTnmqW9IS+rmuaki0FXuhiE8NAgn/9rLL1CQFB
4NAg2gnKJgLbkNedJdXd/BvlTYGAk0cjaWE/INJwLpU2MmJi7s03Jin3wjwjUBM/
hZl3VulIbit2zsZo1W91bspmPvVX9Y9JT2K6qCNdQTdToBQxwMpMv3le7GsJ048c
tQE/nMBU7Xu7fJlduP1U8N62KOOmKWR+8UBASroZjeM8TF/nb5UmBJkCnyyDuWSM
TPOMTwQVd98NzEI3VSnR6pcoLGOjR7XIubr1Vj1iaOZuk4kssxsKGY8N8oKCBEc2
Lvt5yWIem5nG3WXc6udmAnK7S5ZlYhAw8Uf5HDlVJuA+UvakL0Fg1oETdjvCF88l
elhzUQgSQmIeJOkdNfLcaCh1+3X/TlY3hrOErJdip9njfblJLN1sy3or3HGdm3bt
YMcz7/TeQ3MlIVNfGvdMfapXlHZ4zA8dhNOrg7K2lB/Tv9WIjkOY1YYtQR0I3f7J
enMybIPObY1CKXfiJQqNTLMijFOUNIpCMwkX5tP5BWqyvwRn6b4oT7QKhGoAabLl
LeKWorw3bIjR34j/JUhXkZh06ZmJAmsm8yLMiRsfg5Y4FBWUEMQ2n7TsFhKrs0Q5
ulamdwZky6HXLyD0ycQ7AV9Qgg5cnjlf9oOyBd8/IosAWq1B+GyZ325SEAsEN9LL
P5EvOo/m1H5VEEvz4o3tzfPLpvCazgfHpXvT6WicLSRGYr9pFmlPbhCll9wkqyMS
30PkZjNGzGLFvFs6nzxXh01m20eP0/5BRbFqB+e/65KozvI/6WCxgm7SG+GAXLTL
mx3qxUhoB2Zo2xEXtbU7oxta5j8M2q8mXz666lVBd1eqAjVEUAZGBNOy++RDbph5
FZ48J+8TlR2p2ed7BJCs+S3hb291ZLbfWO131K9cHgFDIQ2avRmz1NoaGh6cL0Sh
daBKSh55B1Op5Tpso3H7mC2reCYKmEw++q3zlyiliKjBW8Kh5UQXNFXsdNsQw0WG
Ftv72YEtpJMIv3S9e6Aj0bwQtsGKHAtCUp93AXf2872ZCQV90UryiwWQcFjDInQm
9JUnT28hmaHJFEQwE3RF0Vq50MCC4/SunPSvdBx4ffrpooRNfo9UKu9uaEoqXb4U
nWciN6mCR2BvlaA2IRD3m6j6RhWiF+6s8z00s3Tp+dOR35o6fgCvB292eL40gfoX
82Mktv0w54SzXqjj33gPJXOKG2fHGO9z7KfNae35y9XLsowR6XSuTzKeKG6C3m+B
8Prt8QtTdgtEj3VUCmK6uNiegLL+LbwN6mCCF6FteNyRo5xlLhY4ivBNdmYn5q3i
/aIghYtpDqUxscRwFGJrwNIJKfHAn51gagmw0JZt0xlwjWn3go1oOuyBCtyENlv7
rHjR6J0vUrA+7SYv4uasVEXLWN7tahf3snuPpGHKcQ7BHhlNyyfG0t+7CKrQtKZx
pT0H05T0bgfdRz/W9uQAAP/Upth3R+wzgU3JHyP+FbBTBBrte1YXW1fC9Nl1F1+K
6SKaWxEE58dbBOQcf4sN6Qs2fmvbHYFKoXkA3itozayn6glo+PeJfJnn+gcsWxeT
bgWGl/vY0AprHOuKNhnMQL+VVVBb7FuQZyln/4M2lgUMQZZAWjbcNhNHAVe6QWrY
ME7UJYa/c4/IimFd7oOQrj/ZMqNrVKZVl4vY5CqGcAHN68HZHd1xGqADQQ1YfOKn
yXs1dca2O7A1LVhsTa/AAWJiNAp3bQlaIofLwKXM/frV+XO14wbMHQkkbjMiQJoo
tuOkBOKyVPP6AXdQAEU0kJWE4vgkKRtW0DaEzZAOGKbV6bYv+X0PFJgKz74RxBE+
hVZ9K9IsJQLlxU68iHzkjyH3YCzkQF29KLFYWHEH9e1+w69IgAXMSMPJvYYJMKr8
alFKpiePVVWXa6ZgWOMdAqBaQV+Qky2i7VVQqboJ/e3L8AHucuEH34NSwzuvRCyQ
MgStI3JxETFvJvroov+juSObUpiECd97RpRL59XO2VhiE05v6ZRptDdolYC3sRHT
ngQxI4rY8cqJBQjA4oIwWxeaIkIhpjwCX7/FfHwy4Vkx/WiOjXnZ2mic2zImF/P/
6JYUwpMI4RQ5t7mtjvHo0+/wGjzOAxuxzA6ha4gY8UWAhtsYmyF8LbS1JLon9+Y4
Asmjpg95s1VJyzSobjU/dq4eErkyCb6JMyM0nBYby8ni6nm8tlGsV20Yon9eUWGy
MZhYskIc1itp6mHalsbGlg+ctDhlWWgcZw5IIWdpyMrSYByo3xQd32fDG+lplsf6
qvPKCjEAnjO7EsctW+9SBoVvowt9tIBov0YZYs5XU0rHdXE1JP3awO6EaHPunZmv
MSyRRq9nNPwo/8vgYq+cW8Ve7WToB7HylfuBztxdu+L3eACAI6O75/XxkDa+8q3F
WPdzLeJEfsuuNxP+m6c/qNW2yzqAps4XaWzLxyN4fOI9AHzGjHieB2spMQkiUZX7
AmRnGB8tJE7VEcPBwKwsFD3Dy3ilURMKPuzNOJZjOLRdJS93P4Yq5OQpHg2WdhY5
6piSsgvck+PRl4Jwqdn2s4oAY8Lw962orAFW0HFNa0ee7Go7CiAm5lfuI34R+0iV
2bNOBBsoH1RskSeXgw7ElAGYsukY6LjMBDLBYQF0fyjSAeiKVcQSaac38iUhQo/6
mTUNRN5hjh+UTA9V+x92GnnnHHynv0XiKfOxaZ3wLw82dDvlUFQ/l1UImQ3UxeQ2
U5VGeC8rZZEATiXSj/28hLafuOHbXa9XWO7GDu5UZ/cb4E5Js2L3IXUDv+RyTCw+
yYLdLbbnGTUE11eO0FgltEHcZNhsJIbjgX+DeRm2Wjplh4rhIZvSXWU6OaasLfpA
sKM6QGwYAKWsjw9otR8eli7IF/LNZZsxaQpegABQGfyeMl4fYOOkjo124pw7vntR
XWNouFQvQX9vnTIGTePFOtFRH3twuBjDttj0EGlyrReuQpFnHl0ygZ4gE7DHVBXp
A95nPE26K8GK81xwYBTl71DRJ0jkGjDqfnZ6acQDNHFfzBzccaCwr+6c2XyqxBSu
jindIVuMJUpNuM+L9/AMPP/YtsANki9IsMFZnorAbd0EHkDlHp4/C9lf2Yrv0K3r
NLH9t2kzaARVP/dS4CrGtmq4o5IV0PiibhPCyC2yAuRwBBgHwgg0RTbgk6ET2hjd
NBIJEBVbKk/jvd7U6yGSQuh9CL+9VV90kUV7OjcJz7iC6PW/d5ZAWNmTLy96Sj5E
e5VElGAUv/avP/JMi59Kv2gLKJ1xEaJeXVGBpw9OCdahydHqOY7j4MMilpyVWs6d
8XWAzbtYOn8krVGwrB2szRQUMaV2aNLs96iy48gk6Pf6oSaBXQqgyqiS5hOhJRvQ
XLeuwNhpKLRzICMHGeKzWECX6bNc/RU6CRZTgelQ+Y1SVH0qqhOzwJabEwDZfBl4
7n4QmOsaVBRfdUWs9AYs334HdGcl6h0+UYaIxGOhuBkD23c5euA4Ov/GXpOWDIBK
VLK4dyiCzWG6EVxZ93YjEZx+tPSdVenl0CFrDgA3OJ+SJqF2qmXHTH4Gj1czJVPq
Zl1DwnrE/ODGHXF6fyMbqclEYJ/iCQDphxx4y7m4SRT2LS+28wcXiNeSEvULScTI
Pqq3X63i74aYIM9+RHl3qWX+7ckaR7O5X/WXIIh2gkHqlBhMYpTz/w2L3x+sSaJo
UbKQTJH+Fz2yo7jaPo4vHUiK0pJBJ5HWZy7YaTVoMRqIGg7KgNbiYTtE2amycvm/
/7pMP8QLxSAm9T88I2Xt9Zoz7YPzu/jSukSZZf92VTRrWaiYBQYzcJHX97g8gvuG
2u/vBHx6H7fZBsghuKmlNRRrGR+L22p4ysX2V0McYGNFqeAvjXbvPTYmDob/w80T
pKIEzVmaSavvFpq7+sGUk2UPTaWZJD7NQJhL8wfmEAEYZpfAoLPWyyLo73LJ9yJD
GLyTL3xoYZSla0uRE0wGgZhcPPcPEP2h+Ih64TNN69OMgTVT2ZIhKa9wtePuBcob
CMZyueORfeuxBadvVpEzxUR4i3u+Fv8Xl7yi7myhXfzwFlVVIDw/aH0Y+xmvRlGn
aEorX/kvTvkjUhgxbJxO0JvF2M8PfXcgxqYTRHJVvq3rujrueQEpgYzh7N1QmpHn
0cxhgaxngwLRiCFZe0dKwip807LanWm/LCkinhU1adQ2vv2D6maf1c56rOAxAbHt
lBdKDzLtDIs/QRl1b/pRFdoCHK6ynOsC1znI09ye9NYwIrDB+0uemfbAscTdjYGA
WJCq6bEl+Dss7SUywgjxOEWWmPdrojv6c6hASIa7qCXifcAKHQr3UKkfRHVvkFf2
N3U/UHqFpJQzBRjor5npUWnKLFvK/rxnEgtUosoSKjNrKv5IB/GlZMEm55/w2dmp
ELlOz8StMNudPJ23jtRzOp/FuIwS++O9p4r6GuShaS67931YPlXcmEFGNG1qleGo
/QhZCyhfx8N4IESzzkgSYPtHlKBKCRgh3P6JxnxdYkOttA8FzuNZkDunOCSZ5OeA
+NFIGv4aaVOLoPYa+EcnQyJK4olyr6m0Ww5sLROXxB6+LBKG14axxPf8xBh2z9g4
qAbUldJo/004/XH6bKxvT3mfx7z6OrlvQnR7cXLFxu9YsUND2mXHaiyM3LTKtzqQ
TYmHRMVHNSeAxESDzkrQxd2755bMX4HuisAi4MVE39uekwhUrCNltMcHCsPNvruo
Ao+DXBZ0IDwfk/RH3/PpTFbe1vx+nKY7hbmlOWb9ocqhTiMYAptyBsSqShkFGsJ6
a6BmWzcRFImM19g9ZJ5gVjRaZV5hMM3T/H0XA4boH69P38A3ZfD+IvIdKZLA2IWl
CTxKFMZIMEcsMbKsnIPnD1BiablZ5pwdBqMrfIcEXz6QCy1GZ3M5R1DSmIrZF1Eo
I2gLqvYJJTnZbQ+tja3YcmajSf5DNBJ80D6g4SmalfRD030S5IkoyYLh4ZjTLeDE
HdpR0r9rGjvzccg7rSnMUDaRCBRT5L/XPqznugEjVL3CWiPI7A3sso1b3rCHRPFA
0Sx7YPubJrmMHi7t/5ANAi7+ZFxT/db1dLF0RETbdPf1AxgU+6bwQMoa1taSZifu
KIbQPgK47OVEdDyLNg7EYSDrNUg2U+FoWc1N9lvGZQpP5LQHYH93LOgr48TYVsEz
00MAIFcmjUIh0gi8SznyICOA6kH+XDAFK9wEEPGkT5wd2TRH5qaatU8pQIWLMGR5
4VCoWMM3X0iG1dttkcde88ikCAZS2btcrJYWao4bepA9l0KVCXfVwxqwsoVjQYf+
BiuVq4MnCufHj3DPK85LQEMGcGGKcJqASY8mp0yFveklEQjPe+/ftmVMu1L21B1N
qFVSZDcpOnbBvCzUQjzYPw0coBH/YB7nll4pOI6Lk/pozwGHJi3+yBgiLXBsBl0R
r+qGakYT4bXjybjfkbl9/MMFgzicOsH2v3egu3CoRR/kR1be/+VdUU+JFM1pG8Se
DnaqC3fOI6FoUlpXFl6AoDxIo9jeR8QTiy+TZ9zEyi/EEmZYczQtHbiyR3f51AJf
arIum9bqP+2XWC4CabomOORQq53fG2lGJZmluyV0hON2Ombvpr2bOFkmw3F0mwMc
2ZHBBG/GS17pDYeN2q6cba751c6GX/GKM8UolblF5c715QiAKoHIy3Y7EzXinh60
IvOaeyzpoXLOVveiTRj8BxkuF1K1qydBi8C04wO2M67li5d6qKszgn55LQV768Xo
GHGlWWOJaoZv1soaCeyrt8OVbiZ18kJVLkpVfiqXFFn3wU5s57dInLEo7QTTuUTI
4VuY4cV+sZmu/xDWgonw77opERMKf9o6q53gDJy+g5BQKwyEA/EfzK/zj8eBrT1F
B1F/N3aZWD/L9VT3Oc+kGPdv0WF3fq3L+fHd/jktxZ+y3ah+KycPiM4ntRxNWuZ+
o9OGZvHMECUoM0WT97yu7BtvVeFJSZHtzMxtJTSrOXSofNSTLhRFVidVMfEIYmLd
QKJz3JJUe4XjbIDWDanWgsUVKYF1TAtwnZD7M+g8jHly1cLMyh8LeWyCTL6JyAtI
kKr1EAZD1PC3F5dv/Bz7yWac1rdVCbuEdWKKRs5iZcRC5+Tl2SuLjNcDjvVUFy63
dKEie0Ntjy9pDRtzqpWSKyv+407gjJQQEMrwo4TMock+4LL8oZAncTK5U2H5T3GJ
y6DNdWWBqrlVBRpsIpvYubRgnGKWSnNkdDN452cDvIdJtAVfy86JslRQXhGAdvMg
lHp0J7Mw8EEpgU5ADdSGrorGwGlXAsfqArAoI/M1eseVnK2rJwjk4gJqxDJdfttU
hagKbaHXCdEJXb+rnf3mJRSltG6s4XOxLGaYibP071biHIf/1v49SE+btx7GTm63
oQKDtn6tmKjNq2LhULAuYFLsfyro9AImsPxK9UYXAKL5RaQ2Iq1w+OJGTm3+EsmQ
L2FZth3zH09hjAbJEVf+lxjRUPaqQ8BBJd10OUxLbSKYWCfuIwHNHia9UAprg1Va
UuTCmYuxKp0xZB2+g8T3tchLnpTuD1VcUpLkuNcHpLdQtw1+KI4UZDzSDrat9aKi
XPVELVuOk6NgUN8/BP47epx7A4/iRxYjJw/VIHc5TAEk5RtypA/ddObE5//p/52c
GNVFV3bch9eUgsMFg1n07s1raXWLueBLs4FUpRk60kUwjmb6XIX7b2fA5jge/xYW
XvSoLO0lVzXgC8/Lxm/oWl05f+5qIEuBzvYHdCUS6GmgFZyz9yeikAdGVhqUshmK
5bn0Hvhx/z78c5ZH48oZ1IlsHj5Nxj8Dlz9fNw3oUzYIbODu6/h++L96x8wEHVIv
OUHe1qvzxge/siz+ZTff801EP/jiTYM1hwfbxG/jX1VlQtAo1hBc1+OuCiHdtitf
6q4kN8P1ISwnZZjGDUNiAeJ9CgNdZNVs7v31grW2wovKBRXdJ5swUO+qfND8hsrS
UJgpe7g/qSvJOMtThzRZvjPapnsS+kF+NhhD6Qo4/MHMun9iLXO+AoZBRFL4wnLn
+W+yXkvmTO5LYju5noPuBdT0NiZ5EnFGOYHqPSgiCMAvzLTgZtOy5gzHxFejdOs0
k9GFkki/FwH8jfZVHzqIsPQzH1m7eIOv9FDnt+zmKbYFHR7cbq603WoLIeCRw6Rn
43uygIPmUfDobF+9EYZ4Pyj2FS4MH6ZOrk6r4rCbZ42ap4tx9YpE05RXMk84wlEk
0VWBbFtD9E/xkfVGTWI6UvPFfNO3PwsT0AzWznKT5cxKYM2R7Wo2QiSwuM5WfvW4
+phfnXg4EqYyFqCYElnBhALB8zuJ1AXt7uylLLMzTlClVS/SVTqyXwEIkNLMcaVS
NrS43pJ+1c/UJce/3WXIp11X4VV9gSmdXkAnQJAygJTAaBRmihWnDsh6eQGIU5dy
Rl3RNAAUHlflhKmT6fLFYd3YlzXgjiQwTTXkhPCmzfE/Q5SHD1T4y4AzNqhf6xWU
dq69PWb0zKaKJFikH4bE6aam6wploKmZLujSPS7zKWbuxYD44BOR35GH20+FUsVY
HFJ56Tv2juwlz668kbb4fVy+ZJNOQg6lmxFi87gKmAUvzO2bcqOM6MY+VLj1jvfK
EzdSHpLpxhSgfknkNYZFg8NGwJBzlbnolRU7MYwKbyxInwnL+U5aYUzpuoAhhQAn
rNl/XJyQYzBMBAN08Ua1LFslhcPgsUl+k6rYGMZm9niQoLUMrKIO+RMLUf8t7KpQ
HTsZSbOSI6vnjHry6dPcVPPGRj8dSKvR/H8fR+poTZmOKTnKEIMUToombkct3LpI
HMmDG6ZwIfLN+jL69pNUJUTzxGuUDUUOIPFJx6Xc75EZ5Jz/eOfJvxY4lUVPlUE5
af8Hg7WvxsmrDEFyGQ/2ukeTuXuPtyj4Wz1dEx4zPz05vvv6ExIr4rKdvvSXdEJz
vvvB59TUzptMWRkJhXb2TWn7xR34zYA57TcRtKKD8KxZIWCp7IA4U9OMl/s1eGW7
H1+n5EWpUWEwYv/LLYK5vRxRhQ9Kqy4jKehB5KewwyHIzSUNIxfK228BK0aDmytH
Q8xJne2eUmXVTz4ETMkCuWYOJMJ8w2rf3j3l6bYaJYeDHX4izKtq9zUhxQPFn1+I
R8hh7H/1nGI3qtRuRmbm9fw31OJhoUooKIzPhLoFnZo/3AOKwy/2OMvSh2lXPfdf
Zlq1JTEWffCfizz3ci69e/1Ioe0eB/m3mRe4yCDFoYhKRrZsuh7ShfhXwZQnaEe0
drJ3l2uBKF/2nRg1BnrA8QR5xuIvroPsqWnpPmR/GfFPTGVmx2SR0jRw4vbbuhyP
a4TI3jsKgbWMHxratJXDdmXfCrovY1A8CXvDmrTmaYX6f5ESkyuiHZfpyTuGAiby
/K1DzJCVrUYIuPmQ9Sp+ympSbGyTbwDi992w+E7CRBgZ48Uy0s2y0Eityt12N3JN
oXY3Jmew9rYMFrzVruv72XdlcLW82i45amLnQmCIvzR011p2LbhAgXc0fJ54IZ97
lR6Aweiuitq8DKLGZ34GlZSU1qZWnPkD6qcYVxQoSUNQKeBTyvV3lMcsJ0C1ijIM
yCE+aE9e8ChKgqjFVC+2ZfWw7MYTMnHeJDy3d4VE2Hh7YTaOVaVQj9znv0P6Ibsf
pLj9rkUSVwbxT8NIeyTSiVMyL039b5fznfrd4Ow0CQ3bRA2Ijx4Fwvt/MaM8cqtx
MLRdt2glfjlpvq2B0CjjNz1LUfKa2/qmM2yvzRfWgam/hhpVVghzPQ42ay3nKujh
suraWKW7cx7l/HtwX4I7qBHAxTAvroXHJ3UsuAc5EXe9gWbO8fMfS/Apow5IeOds
srjwt0gQCzCrh3TlKw0y6I0RamWfNliTAiVf6HD4/vIKCZKb7S9MerjMgoSMwbKY
eZm4dSVXnDH7uaMhbo0GFTECAvhmnzojS7ZxNNe93oPoM2ApPvC/723jeKeep9q5
uPfUHddfu3T2eYF67o26EQesNeLwGCpkTaD79MpAwof6R5N1vMdEZFzWluGbrcSC
2ToGpc31ft1yGtuKcsSkNl35aRmzCBM4ljipHAH9PqDIWcKYxaHDZhZH4Q9IIgmu
OZAmm1EDLfdrnMJvI7MpJDHaltrYHD8TgFfRlN11G+f3/jRkYp8BXRx22MKkiY+M
T/+dN2EoDzaEyLX7579FKm/P3cTa/aE/3FHtzHp/q/oE4DBVtnQCYSRL++D4H+dY
277Rx+tqjrogNlQs2U5+hU3Td5IOuw1zQawy13Z/Twr9jV6FSFaqLmq1q7Ki0ogY
0h3f015P/3lQVTlh5xidP7nLHhLIWc9MufQJMCIiPGdFUg+NM+heV8Jop6mTmRA0
g9MQYlz+ExB/XU3ggCwbhhlK+F/W0psCHAxz/RcclyduBlIBIHKnuC6ISLDae0r6
GdBEwYe2zpHPtIftSe8AFI8zb8+T8PindEI5YNAZzmrxyZvgklhCcP/40EppUk/M
SRTBfIb+/PMtolhrw2x8TSzEYbWS//uKk3RFlwxeZX+U/ZH3WOAECyXkjpqwg0/d
s4aw9psyzuDd9EcdMMk33S+oyji2PGonCrXYVqyck4YAkTNqqzl8yi82UI9wOGhJ
0uopYQWUxUb7fic6sZodn+defQjV1eyGwr5stnqM16gIHXfu5kYtYVD/OPAtqkLy
HdgIq5Z2M6RI0vcBC0jq3NucLKcim7eLsOqt8MRoj4oqWhgTNhWx2rifavlYI1Cy
DbfVoJAh9/3fgDBnJPsbYQdS3O3DA2yveyqgY1dc6IWGWb4yyPATPVTrzwSFOmiB
iI8k5YDVODoJgej3MuhD/yLt3N42kVr2y/3a/6ZVvHv5zKlzYWDKqQq7nqmnbUQ2
eE/Ow5z5f6sjuYbrTy/tqxjqnUVjsY5aAILRBRy3ayyv2V01JPwCkKqo0n+9q7jb
vIjWYLqSpdKo5SW9KxA4slC0nfaCSjyjYw/qWNBQUycMaU7FU4jHawLBqXBKXjbM
sMMBkuTOMfyarpdWh023TfItQ4FsPONUHA1k2X3IxIoCor7tUH1SyjhO509niqKQ
fyaf0jIXpTwUvOs+9nYCsyLJ2+aT0P7WQa/VZgRKvTmw6nzi/37QUGJPTvuSx5EL
LkYcgzsJEz40rWN55kGpTLnzG5lwjJ8TjcsD5Gs2qyq2lgBUcw35lwsUFfMQIVHs
BtKdFcB/0E7/fJd/PjgKhSsqEI7zcvNQv+m6DHIsY4yGtbMRU7dMbIncghoCc6cL
OgucKqbfuC9BCt6F0XPIjI2rRXcj8f6w35ZXN8P4nv9BAz/o6HGVkD3HqgrHUO/U
26EzL6P6R7PgbFwMgxVwhgaNZmbBIKkL51CUGMmqDflR5pcnxuKNM50Wu5jxD4RY
2IaLcTK0bTB8/TDp1gZwNoKhwNq/5r3UhagnJS2tDaLZIQyjOO3i1iOi0I71+X03
RBJVaH4ew8bT9C9rTeF8isYzrjcjO4m0gw8AdZxbgsu1NMPLfIGzXIxqQLOdaEKR
xjG9hwGpOraOZz52R6pxVVQ4l5tvbVLZZz9ntO41y51SHeUP2bEBzhrdoVF0iQBe
NUhTLdXhhJYGqLsK6MJHp/utFkBYXIRumxtEidGUC1/rXF3ZBKxKVyMWzARBxStR
ElANlHqNVYJ4v5LKD8bvgtcp0n/DaXVfFCdpYRafAArrzL+oN8Qtw9rzQ0S3Jqm2
esHIv0VDNbQedTztPyqD1bT3hBYkQfKP3/1cBSI2mGllFTfn3LxBKvBnq1QVCC3V
BHVWud/WdmJIMkFcheGXgUnXDxjSbg2ibCaUz9ZO2OHK+dVRpgxD3bamA6R3+myL
29A6CIiy/joCTx68RSNM0jNxbtKWeObRTldRQCQIUGsGV+IMMVRWD8XI+vhKBlvD
53bu/0KI4JDAXF6/DezOMi6obLjETGtSM2SaeQ0YAfPVrivOEyH9XWjC/TvreRsm
jtAru5XqA+5tdOTXJ12A6TkESzhDRO9hnnhnthKMiMSzcdf/eMsssUSU7TgXYlsq
ROl2HQmf9kWS7Rm0MI174+nlI8doL6lJdoVX/LPUXPU+Q9nK4d7bOS7R1Ryk7R8Z
kg9WPh/vw+7HkkLRDh+g0xWlEFrTDMhDK+MuqB0N8RxkkRkNkCDyYGceVVctE5DG
GWiETKxt3rOtynF0T7wrxpRp1CQoL4rCan+S4KZ+RDUg0j27IMGaS9KeX62qGQrd
BViXQOiiX9rxQRTBi9GA96uLk5efQVyGEKJCafWeV3BdTnzDGH7kzaF1jCsrhhrr
ZeCpyhOV9mk8+q8ZY07FT6sCvE1Sp0Ur0nr1RgmdujsCHPIs2l1C4NXbjoXjIE9O
9EW5tr3YrCLnXwVFfXu3nDJZqGR194UOjxZepsAZiCn5/LBmZufq8hNWnSRirLfs
0wxZ9D70HuDZFQcLq8/l82MwDETzOV90H1LmC6heUCLfvDmRyAmOwUgL2UwYZOxs
MPl+S559OZOHQiDpD2F1KO1dYmQ65ExqTz1Hdc/abQ427XHc+ZEwUUiylutNdEYK
m8vr0DUjXNK08smK/IocF3SKnlM2aToDvxqS9LQyLi/8kDb6Uk5zmaFBXOPwnej3
L0hpsteqnaf1UjVPu4lLTA3bGQTECwDK+Dw6CdKhfwHAPxfHhNcBfu6261Dg7n4D
4MGaT2ibZqIsrTnQtrdJfsagpf+lHg5O57ExSL2dKeJKpQs3bzL3V23C3NC60s6t
CZ+u+99H8QUxPoDUwj/xXa701BMrbjlXWL8o3yB+wtQusbD5xPcpO5tEk2ycERLF
+icvUANjTerqmC50V/oXM+pDWYJuDEGBc3lrh+EW/hthakPW/Jx5YK3QK4UkQ7GQ
UfxmNAYUiCnsBc7RltYH0xkObZ9GKnV/HMUpM2sgK1qP6GSTouVe47O+dfq/rn7v
MENDoYDSk6KOWH4Ln5CcqsrJSu2y+btsYR3KaTDQrlJFwNa8DAM3N52eTELMBG3l
cLWCgxT17q7YXMrqW8LzfRQoCp8b+4BPXfL5SYo5Vs7fLsbINuDN6X3kmj3qT3EM
5Q7pm0Qc3JqkEKjNzKf3PLdpF8yAsi9BOhhhsU9wSyFU3NKpw/ePf8Z62IeJBdQi
/jlhitgKGahGnVIuSJagbyNVXC4g6r3D/oZP6ZZS4oyt9bZk9KK748whCQscxzqr
DrFudVSqOrEypf081JzWUw7IZzbfgjIy0DvsLBTk4oer+u70rN8pOYqLKYTydjCQ
6ORifcbgwQQzBgFsQ6BGJyGREaXg22w0UW9GdPJHBFKXQKbXOy+IQsurhr0KoKkI
6QZveN4Ro6vrGshq1R8sBRv90C23m6em5fOr2weN/0sTR92SXUw3qOhM12XeaL/r
2P9E6TkAx3GE2xEyYoCiGRoXeiuPAMMB7LJSkXaKkEN2EOxM80R9G7k64cUcl1w3
0Nt5DqIKUxk8/18V2fzITiCFYgd7DsMKeZXxpzYukP9ZvHYEoDfEAH+bxhEhTLqk
954AjN/TZA/aYThfH8om3GF3rMfIFjL5OJqoHY9qh+pJn1KpH5BzDckaCuwfI6RI
prs7QEiRwOKpLwHBdrdeMaQtYgGYzLeWpOdIgXaxtBMi1ag+IyS53ib22b3RVGZt
5EQEMUFer3WV/hCKEtdvCqXncfARj9H+75PquxD//m/KGf+kV9qN+071EgifABPd
UkaqQP5AIzH4xbml1LvluUH7aPqG4Lx0d5AQiYJXCRBddakfTkTNtqrUFTB8Zyhl
4Ngv3bCAxOACk+GbF8uI01oc7a85tkW7hafV7FOAEWRg5PNaOZfGoTE7B5X+OlRI
1+Nlh4WipWhgKThPvY4EQasZqetzvKrN10gB1pVyZI3GU+RfHD7kxbgDk4Uh+Cq+
ufb1sCizDWG7Ge8Q09GS3xC8GNKWCvvcorH9Hfo8n8T+SmKwv44ZOItbfPrMiHPx
xxu9ted0mTQlDJDJHn6V2nmYZyVKEjOrFVGJhjwtmOODPSuM+lh9AZkDwdbgpxSv
dKX1UNjst9LV/YTKqsTklPO58E2gfJxXmFAhIsn0Rbz/A7ycRPYR6ae1wjqYZ+Sh
DCQUTlgHFsxo8r5lvjwTfWPydEfcDmgfXu4ZK+xvMJJcevLJjgH01PSt1deuGY0c
wM7s6Y6W3qwXgAl+TvELeFioK5HppbaA2Y/JzgHJ48CgkCf/+ad7s1SehMc7fPdi
uQBSOy+Uj3hpNNW9mJjDXRILzQ2Bwr2/5EaZ0UZeSTI3Gz8CUZ2tNtRH8MCv83Hm
jXHi2bq9zAeewRFEL2j/3OCctjgRJ0k0Yz5NF5olKxON/QxH9aZ6A/nbg77VUiIx
gZ0N9tVX8slUjjo+Qr3oug7mccDOSFcO8+4m1mHHWQYhWXu4RYUTWWr2Ih5Mt6oz
rVTBVUQ9ahihxZwky8ftHKr4eqMqTG5AuueKYz1KkWnCYIYSAnCIL0hVhMxIM3L/
udDYlKuNDXjCllAt3cBZL7djrv7gSLH3IM2lelmGw4hIox/C0F3VsIQU5/Nf3AyI
5qhATV+R6s+9VpwSkf4/h3eMai12kFto1Z76CNk3A92hAgeBPlSPhRcoRVmQnhmV
ex+CtLTUsi9+cwIBr/6xgBjfXRy66g5mjKJ3Z/WlDfH5iQ1rCuimH/fg5UZ89KBv
XyCd70Czu1mLUM+elKPj/MwjcO2V047wcPFV36p5FFQ5t89rej8y0JgR8RHG7Oas
dZb6nbR/bkyShMiVWuxMqNydf8pp5bI61AuKy5UnOHr8D+nfg95sM5ZpTU1z9F+s
O6D3JzmPcUCKYXfrWYvbCisyBUW8L9Wd/CzIWqrfO7AO2Z/ElIQQmJ3QZsL6ljAs
KFDtiRD0HbgLbxryarS5md33HzIklfcEgJniqZQq9se99g68Hk8C3yYPqDm5qPNr
9Hr0SXEEWYVBImKSkrNiBHlvVTAhWT4Q1pZpmavCMNjBcuu7X/s0+TBhZTjIGqKq
iyV+UBXZFc/OP+1OI0G3okqet0xvm3Ibvte2hbvgD6wTdSdyGPoypmoB6EHBJRzm
mBNYlt/ZM0gZBHxLUmskx0InHXEpccrDGQf/hmwOTXss9aa1J7s9pAy2v4zNHcq9
h0bInlKe3Y38t5AWrahmI1uSws0fghkbIyVkAsIn9BHLfrzbHrseA/K2oR9e2bPy
TauwmYwqquuLUQ4KMaWeTHBYXbSyo6kxdrRCGZXCv7V5b4Td2zxQUgYAihlkQIIU
oi+yBXHTSt/qzhmpMO4wA6ULiRa5CgX00qEOsnGPvEy8gwHjlyvAVaXIwk0Y1utg
kzfeK+fKWrOdHKuwwGNpBsqZ9gB+yB0Y4xoU827J15iTFUYa7BSfEln4+Jg0uVXq
i8xfCrrEuxt14dbqBw8seFjeEuOvNOyfRoFKwA2hIl/WP2UapJ1cfwuZAIh16RW2
CZZK5bk85IwcQQvmDwdSvHsBq0ULETu8zANeaULdr9254PjRzoX6qgWDgkyYW1Gg
82H88VIEVleI3MaIY4izRhKhdGN9WXAGRz34VMUTsFsisHfoch5ff10f+wZFRVjL
MIwnjFLXt/l9RimKWRQixQd6U2mV3lB2via77a0wtCY/safEYUFpFiTSaZ5NICxf
XcpIJIg1dXSjS0SR0O507o9uRas0p6ckFdSN9s81eBQXU6G2HZpZ7CPCp5YchY4Y
OWgT3G4HHH7UbYNIYpu0KCs8H9vNGMDAN6fwPT6MKZMg2KYTGi3iUpkq4De8YQJZ
FF2mCMoMPLu0abxESd6dxItxk2BXTCE/cgJumRXBNspkrkQgKNsLmhaMOVk66wAv
b+jcJwij/GqNkEEITSZMQebDWow/MCKiWbv/8yKXPWJy1t8KKupkLRh5EE9P/TKE
6l0Sqna/iEqP9Wp+hcoxP1n6L2SKYEE9MZXxuaj190tLZEYZy0gkWa0bnqAlsD/8
LUx8Xkb6btjCGnUlaB/9PUIovhptPJqJsk9F9kk2VpZGCmqfyjNNNWE43vMbo+t7
qoOfU7RS4U/eQRGVYinXT60ar6J8WYiUVU1e2mhMbXlRL4046XGNYnqAreQ6tBQ+
2cxw2VOf6DP6tFy8kVPHLtkpKefqd48U3DcF8oJqGXwFZIq5xkIZuoorWgt5QZsp
wf7sZ5v2aSMwbOgMI3HVcHfitXfMLbLFRAPPl0OdTTBCMaWFV8EQoSro4vezEYTx
GGqjA3H0ZiEmwBGWrp6mThzJwieOFG9fYajELWokr2XGOxxvm6GIX5/zpsFZ/9Cp
AX1SovcKSUJPTrN2XtYOKJiVTrX+GqkHhdgi2/6ExQlS0rSGHx7RbgTFWW55JLCW
zuiVNNXvxyWXyqs6piL1aLXVbKJsdmMzWFetIV/oP7fpDRtxMqjS2SF8G/HUTFm5
tbwUahmIpmERH+CofsWpxvBz1RhZ7UqrN5zQao++7akHSDwHrfl+L7CZBJNBGxZJ
DWOc7ZFNV2Bw/7BX88NYMYooE26SnZU37PaFd3PHSFKUUQO1OMLJqMsj1QRym73Y
eECwy9KJ4W06JnfD0i7uas5pLelGWMX0sa4ei81FMZ4PTCSMvvNFj8/8sEW/oyiI
so1j03wGqarb/NJEV2oJh3i9CxvRRvzn7qDSLDXV7AwCFqQESe5omtaQ6vmodEuP
doBJwojM2WOKsf9AR61GNAhp9AqppRAGpKLyyWTsedRIvN7i1gYF9/pUD2711coL
EaZEyobgweEtj7g2fryEpINAJpOJm121c+zFLaaF+KJYjpX9EWTrGXTyEsYQ+2bM
shZl93P34ZVIWACJ3JDWVW9OL5BTJnDg6xh7j1aDrt/fxpI06M3QyTd6jmF870rE
oEWZkRdXyVlPzEsqtkh/cU3Z4lOoBeytZZRin0Mb+RnePR1ztAbyN06Ue/kXVNqd
uZXrTiWuog2lk2aB8SC/HM9oMCtcfJDO+yiD4XxyRuxsfQuQ/X6NghplNXVLazZg
yD7D2a+T/21Iv42kLL0Y9VUEBZOdioMHbo1woNALjgZKZbWPdsRi6G/45TUXDRZE
Bxz80GreULEmQA+X15dcnxREZqq9MVaaxUO0+JB+J5nuMXiI8WD5bTIhyc9ShEGY
/xhADXKXzog+Ne41U3eO5Ndx2ZMjpWZdAdeh/cxxVts2E0CIqI5h4XibMp/u69CY
HomylInnsS7ivyKltnwJFyC21bPaW3nbgSxXtJdpaMQ8P8PaJp8CKX3wIZsZY3W4
FZbZWWYh3KTTkzYjWYb/mlBI252xxkLqPaY4o9m4Ov15TOVFwpcpQYoitCpxOMYO
OsPTTrGI1KpvVlFhwlLvy5P4ydgDFm1EY6TvYv7jtLc+R/FA6FESLMmZY7In288H
mTlAowdtABJLpTU5JJiyAPMmGN1dt+oHcPEirUUTX8eBtMMprxA5z0vP42bGfGAv
lXoDtXJiBMJMaC+uZ5XEKdWAJLjcBBlZQdP4Pd2su6UfKWn24qDNUsfj7OUX6xOw
AT9pDcrXHvQL/Elpe9FlBH6/wOqlnufJcLMOYWiCQAxYM52T8R1axrYjvC8fMIKh
9IrwKRpyJFvC4occKsYJbttpglEyHyr1UyMzj39XpsioPUDHq+FUNDrfyT8Gsfzb
qLk9HPUiNggTcDfk2wVERuu9BGSYT8anpk4Tuj0+oWITja6d7fTm3p7SR+TBX7iv
nPZv958PjtRI3skUIMQga+ASeGWUtktKV1o7YuPqaQlRyqjao/NYKJtElia4wMnf
0HsdMKJGyLOUMpGXzY9MslskNhEAuVYdxFhVJXktiM2KSMO1wLHnCyMT+7O4RSxL
Q7xnYi+7a8MHX6yayD7C/qQ654ZJqLcrjhLAWq9fFNk+0UjKhUDpneWPeUvoAosQ
F5U1ksw1vtSFonXObcJSACyosDosP4HxY9jCkDXJcISyNlXoHvqMXExS5GJ3OGuz
eLlBzvxDSlCXslhmU4tmYC2XHkhAWTDiuU5PH0AnCj8uk//kSgabVl1/q22Atlc1
NvZzpB7Lyj3WTSr4ypR4aDIPscYimR8CBWoQin0OZrn67Rp85hAAsFlbEvNQ3+O2
w2ekf89VNn1GBgoCen4UG8VBcgwJg+LJbcFEAEEvELXHriD6RqHDrE7pSNAc8EuW
qiE6SmHA+j2uyNNEeFI83ukz5LLs3zBh58qvxsQhev6wFKbYLMvMnGa3sp7fRC1I
h4ivfgWY6oLgLWyvFmJ+ziiuZ182wPw2UoruvCwtnbMLKr6dfDW1LOeiOZKdt1zV
zGOLAgEv/16/pjBM5kQADwfiCJVM1CuzmfEql+nSbymnAm7hgmYl28VI0JBNT3eY
7+XIZTK0TNlhC7X6lK155Gmn5drTYaQh6wT087bbd9LD+/xKMBkJeXzB8L3BFdMM
SZV19Z6iGCfCmBevfCfZzgVo02OdkcD+eDEiFDOAN/UwDSjvbv9V4mGFfO3K2CXC
kkGmeycDeTRySBdXkE8LjTT6hRIuH0yi1XEkDIP3STjhqN3X7xGgKGuNF177ooMn
umVZzFQqRCNtlCzl+T4ukBJPZvcGCpoaS3TaAjAO9TG74Pz61kUZYNcDUKcKv6Qm
YSzB9tkyvz83vFetMZub08VilCFCljz4p6uWl3YwqVtcC+LmNN3Fwaelub7z/fSa
xp4oNKdMwmtq1Z0b6lPoTPbEtl9+Re1n4yVv9qLpKJ7DoayKFyL+wLneA42hoZnX
rSBT1miIXwhJhuFoK6ZSvV2PlmMfuh3lXm6EK7od4QiKaeR6knDdJ2PHQ3O0Yakv
01w01XqO8rUdpckIrjIzRuA5s1SMFZYr2AoSeWgoqOYCnobm28WTLpSUlj46iTgU
M+CcU6J1TT9sE3BvrwdRkMTvdT/6CnFD16mMnw00Rl9NFFam1fjMTLBEFRal/S8z
hO7WKl8ahXoaWknb+49j9bIbExhENvjuRc0h7A22fkSomieUlLOd8spD9DKgFfSn
Og5md1Reo7gpCwMCQQ9dB3/kB6+i+PkgMl1t8wl876EPDS+rqWYjvJCeEx+hKyaw
ckwrPn5SEDd464R9dozkBaQXNA89R6gl760AfZsC7+9KcW1lMbKzDdZVf2soO8x8
HzGCNMpMh+LjbbDnV6iFy1P7ClXmMGL6jieCwkwaC0I9JP2VI71OuP7wDIXiK/u9
HAnZ7/ExspEM08GROab3W0LJ8V1PYEk8PN5h96C1wi9SG+5aTAz6VdKcifIYArgW
3Vi2h8n2wN9OujaohSreyPX8QYNjLxrhPCMditUqLgWsHAtfJKL9Hc5b1Hb3xjy+
WyjdMV8EOMqQJWwSOwIhjCmsDXEtp49PuoJn7LOq0qQxovIFA+VIF9Wbj+SNslyK
gKHrQCMgtiRyG8nppCWZD8zh4uo3S7/745spO+5wchSbe+Mt8TMSIaG0WdJMrR8s
2n9Na9BznPDlAJL9tfxD0sNoCcABr7ewX1set16lclgIeGRZtkzoUIWlJ4ZUC06R
1zcCWiu3Kib2T+kT3hfd0otedk3/vA1njY/be2Gdyuj+Sdh/cJuoxNXlYwmGrZab
DrARtMx2gf2f/INIdr81b3mxYvzgEbypFwTKMX/hWgJf07Jz3/r3MNl4RKLmC+Vy
3KJI0m7wTG2uUPojLMHvED55WbGQYrTvkFAzZq4msQqAqTGBPx12fLfnIL4+MG8q
OfAitno8AACv5DLsh5vUR+svH9lVAZr1lNHlBhZ3/kg6FRH5ZrhVDmQ9QQ3jnqAH
LfWp38uUtpZOSVbyX9eRo5GZiYVj+LN7fGWcWxFh9kcpd3f9tHfUeENahFv2q9LI
imhO1BXuc5r9mV5zocctXbI5+By7Q2ss98apqyqmGzQ+5ct+J5TwqQpIg0LErI90
9p1HogYLm8LYNxlgTRFQTEMoCEDvIMmn64Hdk62jccyAepPIQSKa2i07Ym+WM0tk
RGrWr61pHKXjYAjUWuHlBO5Vr4ycdpgX/uwu+lgrtcr4hnyjzlHfNGFzTP9Ym6va
k/4oPwle/0GRE9yTRy5cuE6t5PQO6zBsZ9ShJ24+udvwxxzbztO5iyDQNAmv/d4s
8SKtsbZ6AZN5HGhW5uhdQWG6MCb2dcmMgvdlhobh8IDACB7nVGsjPzPaIx9kMQ6D
AIlxPgTp667m+0g340B+Qhj56JS4Y93MLCKRFK26/C+krUW7tXRUtsIn4q+XNbgi
HoMcH3nNZ29G6VAFQ+Ou+/zWLOXrXlh0AiEc117tWmz0U5cZnMYfqAJ6RdpPFaNf
dAPiK5E9h8Esq+vEaFbg2iyg/Bezfx1vZ8QxeSIXDost70RlqBwD+ZWbHgmqGzi7
ieu9w4s5AleIFXPdw0XpsNs2mnZtrqbqmk6oqW+iA1lgA6DnSAdKjhyL8yjc3zND
vD9/qZYILa9XXCJJv9RyEgkVsRJMsqp2ILA1R4vkL5XEACjGmnsdwGAAAXkNA3v4
WMDo8+OAROdL4CHFyUeaBMxC8ARjtES/P7YYXprJthC7mooFHt9rgzycEWWS9tMa
8t34uDZOtSRNFjT8Buy8mCb6puw/0zytLY1fvIPiK6Ur4qnZUGkGipAEm+1QA/jT
yWEcDSzcOr7z6msRzkOH0DoSfk47w4TySQQ1HtPWHgcht1I28gwsOGe/u20U3CKt
EThu70OO25E4uiei28fAb9vRJwJ77NegaS9cLUeD63lLFMTN8XcGsBIaiCkMnzKs
91hzY0MB0tC3fujlAD0++KfevG7V9qMPEVK3yCaFBmaM9857WugH4qI9StCtSWau
TU9Wj+f57/KDt3X0DmTkWQjZIhad2idmQdLyaIPXrAyS9vtTW65ZUITnKj7ybFBe
GfDiiSnjw9VwLBLZYueCxGT4Hb+c1w2X2GrfxUnMtrUwlegD5R9QFxvT57vPSrZG
Ykpnne79RwFKaihxoYagxQ9Jz2lJoNdWO5FM5UoZoc/8os5Awog3/pgnA7E+JO1k
lBC1TNQmoGtrciizXq6DOBe8GgmkWpJ+Gmlvwoq35eqXY8IkUjC2XcT+65xBa1nF
zsS4eRsilHQZNMTz/5pGwYxfteVAyJ7RVhD7/NGxOKkjcYtaXV5wMBCd3/6lyqwW
3yI3izEGs266bQMT0dEsBNgndBYNtBgVVvTf2fYl1y6Nb4CRkNaLhbA4nFeF78qz
Prv5EFT9pozITnBmh/FHYgx99U06pZNoG2mHXqgDfQztBvP4lPRut0fnOAbAs+gm
dMt8aTuqddGR9d+vSBzEQD9N0aXvfTO1609G8FTBNbVmD0g6ilVWvfXrtIAPR4VL
LLkBSUhdBvWf5MEVsOMWWfPn3upvx+LZPtOMb99EklkQz1FYfx0LuZ3Zx0kqI284
cNyUViiCwEbT8uJsYYGtmO6hx5qaF/criQdTBFYNu/mOHa36C3ZlsrgrgqF4Jupw
/IFeDaz1ZrCMsfkceCVSJK+C0tyRhXP2VeVZEiDbBic7blNju8aawJ0yHJj6fl/o
e8Kk9Cm1aLNnnzsvSSH4j+Wa5xI1sTVN4F7vcy0d2PittQFgycpR/htV+lZB1QLR
Hafw7Gg2R26y3yI4p3/FnlKnt1aftqkh7hmdJd+lzzbNFFQ1AKOys8yB6qRltwLP
KUqVRhhz7dldlwCjcGgWU47eDwDTThPcHWVLdSya8/HcWfIkCDuNkU+VImzvkIDX
sNHjBdkQf2s+QBPFieUaTseO1FFiM74AmylwVbPGWVseEHTRt/cI8LsO2bWYYS38
jNgw9ZD3J7QlwJp2Kq01Ys6AG1fbleMjRu/3PXUGBx1Gj+gYvfN45yoyYGyrl37s
Es361SKhuH01vmSU9dmnLHS/VvnU4VVadrCf245XzEKN2agqoJfrntDuQdnWwxB7
5WNs28DyIUs/O7fjjSJfXQYQ/4rZ4wfLt9PVR3B2s9lFRFSOuun1gNLW5ZSodTAM
NnhSPDB91OiBP29+E7ZyIGF1VPuyKNnvd698qYGSjt3wKX1IAYWWO/8zY8bMbgfM
BJtCP3K6R03t8lDnxp1xpYsmsAJXBoBDYDZZZ1bWcMfSHmDszPlQHnLTR146XXdi
em8j1W2z2xp2PQWVZC/w1022EZzm0jydYR1jhdvwtIefAg4hLAvgVl2OQhJUEERf
TKVfRvVZ0QsPXWTnxTincSc6pSxqgOSSyrRiJJwQIUyTW6p/fVLeY3pI67ioYzIv
rLiY/+nsTUQahTeI+D7TQOilgTJHgqjQ1iYKY8viK0hV+F82WqGcSkvgDEzPz1nv
hLJLy+POWUCJ4+1LWO8AsRdmciMXoVkOaOhq8tBz24pTpiOCUFBEyZGX2HpmLmi3
+xr0DY3qr7vAmHqzUTxsl5CY7YMc7zChYlhoKkyKQp2YN5sglkiBtcP24ZJhE8k3
SFc/QOooiq49jUA+ndJNtRx2QGWIEvidZ0zAs2EJgjeOXqQxYg4CuU9RKG8ZHEeY
9ALrckRxoigm1zckTMtrB7laoAKn2kZXgVxiW+djfh3KnxW4s3+35qv0ecN+j0xD
5f1OVHCJsPboY7e78RYANqQ0yVUe28CxJlc4ly/x05daQm6Kx8hM+VUpZRHAYe0I
wWzWE4n+IknMODE+uF2Z2YbS8y7feebxRKEEX/jEkjf5dXZ77ZVUK0E4s8+CggXB
lnFIVK75an9ZsaDL+HkJSRzLuyhGO2DEiyio6t+Kl0r7uZJj7CEJ3HwoMfojf2Jg
vGmjQZD0flyFEAKUauaQoOwbkIRaHv/MSAf8/TB7kP/MHJaHD/h5lJShtPkiMhL/
CMuVMBLtPVnTCghaeddLMTPHlZRLOu0Kcvk2xhPd2/pGSBORqHf+B4alErjls2CO
6TLdMx23rk4DdqGDC5Dv65IxlNLI2hV/FRIsS28oGIMHBg+EesdncqPnfp3Dt1u0
uZbwo/XiSEnE5MmceHZe43YobPKRXO9NFpkBuhQyciMxhGXmD6BwZZejyfVddaTl
0TDaZhWwuinqvTxaRrpKRZx9mb2/2H3O2vWgK6HLN/30YXKLEzQ1Pgp9LagMrYoM
77cjwsrJ9p8FEvBI/UzKXKBTui49mt4K5YfevH8obkp8rqoMKusjizssjz35LoVC
NULHPqVAXft298caEGxOe6+PjS+IZkEGLdPGS/bbsYChGjnTSA18qttJyD1S2Hed
Ip3Z3To3JuLuCh1inkyGftDw2oeL1bVDFJwszoiXIFzchll4PaS+2BGxQr6lwDlv
gw0/ByhcGzQklgAND1AiIxBson90XErJ0pJutJB7DDkzCtamTxHaoaBLs0YB73w7
mk+zM9ktkmW4eFULjEr2cMtwTch5Afy0wsLKwf5A6Nj/nPRoLB03AT7u5O3dlUHl
v+tJMG3q8v/IX6XlS9MFzFa8onG5Y5D1PM5AzM7NuBd+Vi2yo2LmeylR/BBhd9rv
iIib+zkHY6S93eONGqPAAfQYyfV6XMUqK3M7uTvpfbVSQFchcRCbDxaEacu6xGa3
SXErEuImuwA8Ycql3Wo4vkiEpSSATrWLxFcRST39KDGnOW2eBG7bnBdI7KnmPf7p
bHHR2FW5KYp8yZVtR9aDX2XvLIoSxlhQnnzUHRQ/ORvyAozjb6szGFbI8WIGz6A/
78cGn4rMItanLj2L5pO4wyuNca0XSS5QD4S3XoU84UMGCrUBBMtfu4FAbglz9LQT
LoPSJA5AHYxijsFE7fbXJcH9TgU1xYlyErent9J96sRZJLXG2AZZrJN8mOW3Q/za
RaAxVcB+/QG4urXS5raL85lAAT9s7gf+gT9/NEDzTb5aENxnGEVSYnWDNVy6ZArC
RzP9reGqVwXFGa5eZ7epUx+JmJUAtq9TubstRFhhF2Asg6mE1vaCHNvT4fzZkkGs
ks/1/w3lzmSDmoxuTLCYdwGjeQgDUIunbib+3wSsBHPtFtrVUH4hS1mfE0s/OCde
dah7XYTypQDbc8mVik2q9hHHNTOn7Z6LhuNsMlM5+6FipnNSTyu9KbU29SCxiREJ
yXvAtrh9RB1VYb+WqOiKbHTX28cX6n4a12YgNcqDmaJEbVkFqgXmQ3Ks3WssC161
9UXufwSIz6EN06fg9TG6SImU0rvfRRP+/ZLdHh8ejhzSzmQtMvHY1qpIUrb3G2Q1
0JHsYaJs22zuH77ooRAWTox4Ur8Ek68MlCMduevQj2tJtbxS+J40F2+eXWyprh/8
HKxFbJs3p2dKTSdRvPxIYDgSQauv/BdyZ68Jm7CJnRqpJueKd3sx1uphLOmg2Lhq
wga2ViHrahzS2FejZV1quEB1gYyGoxWB1G+M6e6RT25WMhjNdcjT4kz6swyJzEDZ
fDL9TO8BdKZVSlVCxcOrOfppCW9qlXiMhSPrwmYOOHcrUMXTCa9kElF07eEixry9
/b0yRKUg5ZQsXVQkkgtwnL5W9Q1tligkryaXDq65gPUrCGP1gd2TE4pM1qXG86t+
6R/Ids1f6eFb/j1GmQTPphcEslrGTlPtoHhTo+7XUJDNbIuG7R/RCBWw/LxI5VnG
OjRh1uPF5yZzatCOklvxj2qDQHmyVQoMdxaBlTkS5iHifEpKLKsD98ap0AHscdof
TygHISgz7blgF33nJSeFodcWBGiDQIvEScqB70Yu6+WZAwgixAPuqSD+JkSQMtIJ
s4rcTlCh5HJaEsuc4q8rJ4URZJsLNnBWmEBjGs8Yr68vlmJxALMjiaZPNaWPQYmC
Bp4q+aSZjrDE6p5D0IWI8tm/35lAJRwZ9zCV/95vRZWThcJ3d53iQ7vecNiOc53q
9VnMkAqG1MGmC/nL50AaQk4GAhLaSaCq0X3sWug6bIlFtss6Xy4DHYmNmjB22Ki+
86HqHoK3QOwzSZj9NTaELGzwuf+d7s5k3yvnCWyXV2mjidrI9X/VyE0xUgHYtdPi
Rfj4w4yhiPJTVg1ar5R6S0+DReUrnScq4j7ajuiKFBM1fqkhpj4cI8R7O13U0vzj
AGaSCOt4PjOj+i/DqR++ClyfWZbpsB0SiyeGRzTMUNiFAODdmV+8ZHOzABpjcwJa
n3olma+ntT+/7ogpo4YT8xfklhpb+wf6nS45/XKTdNP33TrMZJZVPiSey73tCNNl
ag88xMZ0fiBs1HxMVoxVwc2RmggUjkJdqLttuE+V16slqnhT5VnMZRGTcYD4h4He
T18rZehnHLda5UHHDqvmlZgdYW0O7Sw77d7LGXcyeUyB+obluYgxrhEVBiP4MJXL
jhuNDvo4L6fMz6IUEs0rDibTesFDwG6sW22s1hCq2rO3cdZOvWFqIZsgN3ZeSPjX
GwLuyROMeVir9CLrUxwt2gG73FgvU+KydaONgmnY3xmPEA/P+K5/8S1qjn2ewKMs
fTZ/yZ7AiOLq095eld9PBgemi1kfpXt4sZ2fsIJWiq/bXES6An+p7KrgtUzP2xWx
dmyudpL9oXP2fr5QHMcMsk/IgibIUDQLPjB642mucZr3P/8wJjKbsR8U2046InkA
ga3wY/qxQLYEQ5X5dOKMjgq0jXrDKco23uSrnQoU1wsxborBhAqypqlq2QbBlVbZ
H5l8aWdGGLVDQwt1E99ZKp/M8AI2D9KxcbSTyfADZ5wz6KoY4DN3nBSGfkPaXNcU
66bqiMDBEECUjoyCPXTzSc31Hctcg3CDHuaagRhIxDqnLsniFWJLFixorcJ0m+2i
jB5H4EtwqY2SJxbEI2Fcif7XLZgImGd3w7eG82lU36A5zUkA5/iUUtLKVKtvWrYO
dYZ5LIlpngwEsZE4MNdEiz5X+p3UasI9Tjhxv4tFG4MdtxuFQMTdET1io9XwPHJI
0FkvQ6Sr+n+diPn4QPnE3pkOeSlgHdtUNuOYP//7tLVy34D3JxaqoM3BuxO7PR2Y
Tet3YGeRpDrKiVsWg9Cnhnio7gSfUppgjpEDzJX6dxuVRIZF7gsxOWtCHQZ32lnn
x5LdVG/jTnFW1ZgfonhCPjJp+Bu8/2kzh1y5w++71Bo7LUM3R6zC+/xZbIVPlD7F
cEUvMWZqC7AK3CelTyvVU/wWzd4NJ0faqFj/jOk7/Oho5cGhCW5tCa2jAe0F2AK4
dhQe/iIB1b/HxKqoMVt+8SpgJ95KSMaXwS103FjtM2XPMhWfin5Xn9sFonlGxvT8
s13U2mHbTwMpK8B1Ba13gSRLGJaw5Y35RFKKZsvfbLvQTDoWC9hZ+MyKUmHtENmq
jb4DQMmhTDAva/4CG/uqd0hpfUEzzV5WcdZesr/O4K6vklqkqzaoL+yjcf9yVk0V
5nCeCPQ5rE+SjdKfZli6/k9LvoND4VBEs/eKluANIAmYbdxo4db4w/VL+uDfXowO
Gz42a3flC0adkMPNSvTedg/8Mk/2rp6DWrUiQ6P9xfFn1AcnIgpH6qlk0vgw12i7
uFbHlng1eYnBx64qrxdhxW85W4whdofzZNu+xA5H0qlVueXiiTlaok3fklh5v/6x
Bkk2up3Ngry9RCxn/J//kKq9OYIbdYSx2Y+Np/sZat9FNbQDd+gjLuTkU5VDnDQv
aXyXbAHyxceXYhOnWpbnkhtrD2evux1I9+rob8HSSvmcF1HUsC1P3s+yj5obwUlB
hbegjn4PVYvBw8C7USVJZYHokyM7jaltbo50v5l56ZsT35bbJooUlA1ZsqdciDVI
bulorPO6zmAjl4bkw0ls2LHBBsxQOYMngRT9vF0lfKR+Z3NthSsT9WPyG0q9lsOi
plSZqLZwtsTWwtbgsUBopx13nDViW45CA/BpQwim5MFb0mIbJlceRi2NEj208R0B
9/5kLjgTulCETdmGqTPutHiZhKfNweYsYkzQFJe59E6SSBdzy93eQHZSTVshtNjn
o2YkaecViR+mO8xbFbMIgwCbu+tBR2DLZT9bGeMeZ1o0vIne4fD221DcKsTAQbOX
7eMc2rV/IOnzzzGhnVbXeUV548BXI7RcRpz7Rr2ZXqHe6p5SFpNg0TraxvAbDl7k
8ha9SVrMrvwLIkcuEBSsFceoq8WZJGyzsn7diisaHmZTINJJjxC1RYU9II3ofRrC
83nQOVS73V94FoKSyokAPq1oEdTNtaSmxUqnMKKssHmVdX47LHnXT0cjyE4MTNwG
DTi7uDKYAcYdAmFHuwlaBUkBdIjVHepJYVVa7yMB7nmmcWR+dOJkzbbsWZGRF9fK
qkyr1C2QYs62lKu/4FxOi7vXXDQy0eOEMcNAySredIRmRW0w3NQw/KobCi+hjCxB
5rwr5HsK6P2IFnTo2m1CEXry2EKqlU2PwrWxBOsLW/aoy5OQEOiqxWe9R3d0dD3y
ZSuhO2aw/XSIFQzwGfPUzCwNZShSGJuRjBgzAv51ZDeV9x80LMGKDvqDyRmxyzgn
zxroRPBB4o1jNBWHotAsP60lj5ttz71QaMLKhQ0Vxfk6tnwskWWf0pe2jw3yUubC
2YMcmk3/eW85FUj5DfbZ8qLv9p6VJWw7jMfBTxjz6DSB5NeUt9G2qaT1d3La9RC6
0Ar3AUBUTNdc70T+sniE3xBTvwesS9nn6LLkuKZviViKIPba3VPiQ8A3kYbFGvdi
o34x9x/QZ6fj2Gz7OvagdoF5rHyAMBxSuLLQxikB2UcRQmK5OC9Z+gz4CvhZc/27
6cG+fNr7fqSbz5ZDgsjO2WNxvA578yBADNF389zK5VZOVP5PsIHAVq+VCDRlrZ7l
GP/dMgUqyjfCZfS6nZKEk9v2PZykvg6PF/kqyI6A1s22eMI6UqQdzEiLVXp/Fq2F
qt7ZlZvdHm6VqbMAJOruQaGbcXRavPDcQx6PxoLBPqUigAmQ2b9q0yokuQLJxRpw
zL1j6lKVjXxGKDbkjAjPE2OuWCIosile7Qcx/VWXR3Lusl87n8aIFICr8FPI0fhn
Ky2UCmXaF2wtD3mZXpKk8LFsz9qaDx0l5xCf4XuDp+/klHm4eOWrW+U0wO5pgVSI
dzAX+B+Z9RmsAZ3zsX5w7ZhM23QNQ873XJl8zvl34M3Af2dbUJElF3yqkXoo6C8l
hbIpmfMNa1IWnMokMkroy8czsNY59UCAhdoBHc1SN1Z/+ERudx5qzzwWXfIyAL92
1+nDwfog2Hw85gwV8/sbmw0YSZhR414B3MWFR4anSiTf8SRUGEIlOeEBkPJnJ2Cs
0kSggtTU80UCCztE+PMzTcWvTynMwPfK2T+JgI5fE3lm9EEphtR1f2XZbgOrQ9jI
bvSo+I+Vro53z2SZCBiNA9f4OpclRdUdPqAbwdCvYXvalmdKMG4bQFOOHqEPYLj8
8+P5BC3AnPBxNtTAZ2WRhBvkyZg2N8RyNA8WfPuliVlS2bVZfxiDm+f5a2DTGXUf
GNvQOs7LqgaQ/UIun2e/JFXXR2hu77n8paWjM8wQp2onelppTXqG10QBh8Fa8sdb
P0W25I1DS4a+4RUxgSQWH5SMiiHhzAppaRwovM996KtVLsjCoCgJSIify4DBXQ5V
scMDQAnuw1fK9eXatA+LVAtdjgMMhkTXGCzXPfof0NqzFzodSrBFUrPA7FOmb4x5
cjcuaUeY0yteizjr55pjTalzUGqKMdnZT31HG1RN+skOqvlpdMeZQ/18szpmfqe3
08bNSkNLTCuzSOsUdBQ2N4HMNn35GFuAIvQFjj7YmfalXjlIC93JsWhdPTeHF9dH
93IHupveJusD7MW3zIkdCK4a/FPBlLVmPZgGPd7E4NISt9Ad/GaYmTfnjabupEIS
xjWQ2IMXVHgXnWZd5DhnIoLiM6FFddZTTAk0oprPNKVR2qO0+oNNFUX376TxUSx7
t3smJS3TsbHjp2nfcI7XXxyneb/HoK8kgJO1bqRqhJvoya6PPkFNiZdDuii7rcV5
dfof16CE+Y0DdeiTGFz8M5PzugYJOTjah7XfPYK16WXXfxRb9Nq2UKxL6lHHrjix
3aORafsgWsYDn1miIl+WYv9r5KHYlb8x2lQVQ8R9JYYZ+9bVVq+Q6nqf1sU96nba
m3rUN13E9DtMdv2zC9noZIVFGp8Qrzfqzg9c2yB8Mg8whfO2zCSTbq4HdSb/GoJs
rD9JWGiPkpE7NOFFpXpv7gAvy4nm17a4N1GP1UklrNDlwFzc+LLAH+dskA/TcSMs
ZMgBSZ+WZFvi1TkyPPG7V1Ww0bMZdWXKXFP59AzamqcAteKSUKYRH6IpkZNdB77m
UXjmgZA0xQamxxY0ANWmDWmFVL0NP74f+Vt9JUjfHdJK3iKW7eBcxGHhGuGL5hNb
gM5VCgg4ar6IevE/jf0BhuszU0TJWK3YIi7ZiB3b1yV3ZnPxEBW0eV1w0QF5SbMl
+VEzHWpJ2/SDRvgbZ4yFOimbwfPiLRCLSRLGNRp/z/KSX11mUeUIYhN0GFw4PYCx
dDnZHDsxLpUYKT4yg1mjPrsP9hnQ215JHz2y2qrjg6CHoD7+o732y2G2oZWyw8ln
mJt4Z7VoHxHqtGSHV5RK/gRAC3XISIayDiG2LlNh0wFMOBH1FAYfuo5oL95HEFwD
OThdn38uyu/olmdYBM89bpks3MzKcnSa32xib4FD+IE4XcTfOxi2RmcMgL/Q78VD
AnLgv2t1uUbRVigcVmC3Jl7CcRrzeXDxwwPOTkwEzOIUWzjWqoiHWbgzvQPisNQD
z2xtEGdyJyG0aYZgSk6a7v907YZDF0LYv2XiJz0YfAGMidj4ufSS5hWnuk4yPu6N
m2CXbbBWKi3O7DjCqg4r5m9jbDeAMqzQpTJt/q33b7TK8DVyYzxa0JVKT7mIvMu5
p9FiK2ijbp0Hmt1021Vb1ANzn7HYYtNMJr2kAg/dZkWOZrJitmRQdxrdVsDTmOOK
eahwbBA163nTaRhJpjNZZ67fItemPktmFsR/cKN9Gfi5ZASwbujSLIDkVws0Sy3x
D3QQ1KXV8BIQWPXJQ/hCc1ZNwm+mw5I8Q+0fs9K/LfyTJ7jGNaXkzhIHSsqTHcDv
Y0krBXIrbeHgqI9mimDDOWDoBeS+42HY5GgjhIfe35MPd++KJmJCVeod+8ABs94H
0w5GH8cTFP7NiXDCL94m598H7i9sgjTCA029opRnebXFiXYDUixnOCqDbahJkJod
deQRcKhPFiNwf9SJpdCOpZHafrY+frMNhd9D/ZtCrOG1xTn/V0ruonqci1Z7mh38
LnrlkuYCsUrn9Ppct9nf4pYp8g00z3oUiMMnOEoGJdOp3iGP+EFZZH4GBHceW7r4
XT1sE4Mt9nxnjRM+7rB4j3CbgyBJvFfYbsJ2qVMnVH/qd8roTaPsd6thomc7dnrt
KM6AcwZR+ClBuiIgGtj0he/GSTwagFsIsF5SjSrISg5kYjdQLK+C4ZV2em0jfxUz
04aBI5CVBMA1E4/Bbt5gDJs+Msx4jDWU6VZWgfwGHL1V8QNR9KWVBBqeq/yUO3I4
FIJ4HfrJwXOhbfcH3MdCj6dzzrnXZIXjFIOTywoNHEvbZY/+ocIv1AbJrjLcQqK9
6YBI6ktPjmy8CZ5u6Ix/B1g0zU0gtdvNeID66BJaJsl5yyeA6X2tzLNeC6g5E8M0
PVtkK7MIUWees/aOQxC1KLEhwWLoYXJCwI+6/3ubqbabAZG5TP3ul7gboptoBJTi
idYzkJEItrhAmPgdGryTwJcMKIEvOtEAawtEbNxVCO0z28xYymNW58FvfiV3guKt
AHDKUvvKr5B5HEt1Kal8qsaCFO2/uzax+vN1veC5NuqMEh+QnDQY4SXd+seYsaOd
F9GXG94k7yrhxymyP+4AV54ofCjta8duPsJL7kBmBtz3JuRmDZeIpDHMcNBKlT3+
0ECCLDyn6WHDMFmO6I+pt8DILTHgxOMyQMeUWvCyZvB6REsX5Aq9nByR9Q4NO65y
3FKHou/8boDjj7hkZvGS3qpfIQAbi4r48FckFAwXD38u1faQltTOhdSr95+t4pRL
rfXlXYMztRoOGhtFcYAeT1xjPhqAcIUvbYFP35oH5jnR6SHS3c4W6imirLtzV5P7
Wcufn/2cutI1UiErPD92mz7U26maGJtUpDmcr8pPpZaVZOdJbVXnhXzKm5WcrS2Z
WO/+yZb6bcDjnXNNOo6NRKK12XAUrvUKxTk72D6D5pxhS8v3h9r7mC0wnLi7MJxt
dmkLO+/6qXfbvqveI3ejp+suQv7SKBiniQnOg+Bfkfnz/PQViRFsiwBHcaZyCeQg
AEptXF0S7qpmjB0Z03NUBf9vRObEqajtsJCiLoPS91DMif/fEODhMcOyconw8s/T
wf4VFYWbodyBuTgnZ4RkfoqDeksiqgGG/87flao0MUUd42pOIjBvuhhnx+wN+wBH
5Bzw23htDyI5lc+xw18NdyXn0xw2CwKk2A+HUuPEV7cjwND/w7GZzFaAnBKQ1v2j
CA1ky8+byzagbCIO2V4lKQiBfbrpFGaR/5x9SRUkrTK/sc5/zISb25hlXOQy0n+a
xPR7yoJM9UcekaesBMm9DZE9fK8wp3OmukM/9u/sY67mrKFBy1Tr+ZzkGRk5SVVI
/0zZdXZnGusKpS71kXBVgn4IJpcLdtde/7sWtc7e0oO0KyQY1In3GQR1hnTOck5u
H2TfnyKdGMePpKFtq/BaGFAjf2rR9iEPIjWwghSlgyKBt8FGU6JxBxLLRpyJk9p4
Rnk/DPwNp8zEAKOwluUfWrqQvFf4j+NRdTnoZM4LOUTZ9XJcINWuALQ0++8aDdlA
btAIA1vgPvBPEUnEafWWDFy4cpuj7eTtjoCnQ4+qmjNXwXt1GSHJ+MJ/ry2NdG0Q
Mbuhv5Oi4RrMzbNt83MKmTYmHa7LO0slWFDx228tQDDSoSEojVuTpY7FIsM/yQ/x
S/LaW+tK/FFMbc4jGh8ZQh4ThgZ/YDuFcuSUvJvLvcwQ+Fx6Vu8ZgJ0hC197Kp5E
NkhoJAEZ6KeA+NbP9wUKcvD+rnRLaRkTFA2rKRIVUdy+Se2TA2xZQjwqnnKaKyxL
Ga0bqwfcaf5nj2KM9TEdNAObJD1UqcMLVmWzQ28TVokygBn9YQZBy9gHGRYmbZ3+
9wccRq5UyMnmKPaBoC2jFsbYgL9ce+jvqCQ9w+5XSgPHq1NlE7estdKWT/NAsarA
IGirmBWi5QCvrpHRyAwYCWq2OJ9uz0mMNqDqgewLg5c+FNaK1hWUdlSczJeNsHr+
8zjDE8BRAqGe+j69weOF/n4fvLZRWrahywQWHFRzTFRHBT667uumtp4ONs0PzRV9
NOxWv2mIXfiXDcTEFSkVP6cxj/ZmLgUqkqxXDa9etrM+i/feQV1Sw9bY2Lec96qF
/p00wKgBDKXDj/mptKkiltsAKF8c4eCyywoKsByeuUOo9hs1ZE+BMmISjdDPfRvJ
6NV27Zks9amfM2vDOPkyq/KHwf59zIsRPVNXaMiVKn6JEQRg/bwg43snH2Eph3Fp
vR6rhynvKmnFZVlNAIOaPDvrA9o/EmGZJlcTacDj4IEnVTda8PzDLyT/J35L8wqb
GN+qyiSmcYai4cDQbDtpYWLTTmz2YgsVXidCPWvNNv3Z1+0GQlXFvdbFRj2YtkbI
ydOie9vP75v8s+27Rrr/gWZafk1B2jkrq+wG3kralCK/NNYaKVeWuFXjvtMMdV0M
S5aPbhlhYGTKmin8tW4KH6WluC9SiAab/TXQdnazh5vdde+N4/KTB6+2l1kDEgHu
8itazeW28nbDxg4nl9UY8zg7TbDWpKYAutTw+kqlmDUQjKBwKupRaK1Eg7+HdD9A
aFAQ6QS9HH108B3GT6dLoy+Gq/fOOBVFPYY5yF39dlT5VuIOlCRtOKd4qEGltTzz
P8V6/g9IjV8q3ggaenQ2nKULuBTnhbn+odG48Xh4YR83VKBVZCs2xbosoNfvrA7R
5khN2pndPZkKMFXpJhA4VvmNZobqtCph8M+R8qevj213/+Cao6k+lis636WpQYxt
rS4elY4oRAdTFimdy5gdAQogL+/hnFS/5u9UfJvAZR2aFUojIjgv2A5/N9EnDrgI
DLlLRSbKnyCXqoz1VwRfEyBgc26WDgMMmmWKF7X/kFLayOM82T0EPIevZa5d0aY7
g9PLj0pVU1V8TRpT8yFdHITdIz1rK2wXZfTcV6Kfl1n4eRXK3rbQRi5DJshhqbgg
dRzeYG7rkarqQAi8AvZ1oVn7TygckcWokYPW2bkDf0PItIqx4QiJLYRnR6yavQGD
xWuYKhpYLS1FtmPqGQtIjU8RDUUW0U4dz5zOOdqSwiC6rpjdeDTKjTKJox9+jDTX
uk32LczKsPhzB4Q3vPU044i13u49mAtO92Rje+xWxTEJDsSA85WzRQAUC+Kw8rcY
yIH6wUdOZzKc4qaNo4xzfiL0Zl4mxbuJAaxg7SkKF1ynumwFquJh5SX909zmdGKu
PtHYUIYToLDMEc4fmSXd1GdqBzYsUBgS6QsunIjeXGB5W3bdiHdbsTYqOUDT0ZoT
GwVn6dofjVlChJCZ4PlG9FDVuAm8V9p69vOx1hSrd+k8ElU3obe2bWMigwRgB4a/
0GvxAYkZJwfNTdRwjG8x0nlqE3R4Y2js9Y1Zbuhxt9I/8mbML4FcdXxGfJzwVH0n
6/6/Abd0YBpp9KjeBLeBSGH8OXThWcEoGGrXlEajN+wVytzXtLBmWHWkOGshM4xc
OMGwmd3ARnrvnF7xIDEDpeHzO5h5WGsUoLs92XkGoVTMPnPw+KXv7hQkP+Q8YLHJ
J89j9ZtFi4xP26tarXK0ZhX2DIP3+cILVb35BQ9vUuqpfTE8C9/bDIXFdLN12Cql
WA3uQreul7TBf8SKPe3fRKLKAgJj4H5JFHNOdZTZsJM/zkfOxUkHHfpzErwuYWdM
z8wuG75oqhE30hVwpHyEKLgMaVtb8F3uF4HNxSjgtW7kvMzaQMQYWNxwiEhyZ9ze
IgYCF6HEGdMJMLGpQYtAWjAxY1phh+J2l4d4L0gJGrhGEyIVKqzBPUTrQjitGW1r
Rs1vW19cSDUQMnzwJfxpz4vi/fOGIcsGgqSBtyTvQHOeoiECL9bim9nM6gQU0fVL
S76YC4UoIWJJZxVQBcjvg5Q0IF4afyV6KIyDlgwT5ZHaLB/QVHRbR5UFicEFb1X3
hZFmYhj5I21a6MgTSv1k2X0lNkpJGSI5jXZJ9zKXXedG6PVrDoxBFkqKAQwwzvU8
dnyxuv5HUN3FbHHsE8vZlpdZzK/t7SgzEGq3o31w3KDgL+72W8OorV2X0YPCcqhA
DtFt3Axt4J3TlRDOUUvOaZpGl8pMEogJN1EvZs+BnzXjvXxlrxH4ZGw3tjd32NFx
2J4UOnx3p0vfXQ396epb8/P2SGSPGm9AlrgJjA5iINk7KZfMn0IXbyrzug4jtBVt
bkknOrxWjJNty+z0hpdLsJH0F/Lrff3K6JdP2XMomsVqQbYRVp1DLxZvLcMdQCDI
aJAmXKXIM0P3n3qU2XnrCo9J2YFQmvSFz8JBo6qOYPqHcChmnQtLu2uXQrv3bwMO
kD1ZTfs9M/h/tdfZZTlwga2NGfffxQCozvdacq+9JDCMGLw6NR0lFAI0jQdlvqDK
7GW51nIs6Iz1onCV/6G7yAZ2EPUwjx4EYEydbzcGeDnMIZrcA4HlOLDw224diZxt
v01vRY9CV6ejwYzUXC68xR8lemK4dvKesfsMoJBqpt4d83rp3D8SrJ6YubhcnB+Z
eW9cN7LXWS6vOjfo/zXqu5S9KfbVL2JWtbCfqj9eRNqGxGcgNi1PUINcovMcEkp0
JtSnlYJb5oWiY7ENEoFn6AbtzftlehOfXmJxikZZGfx0IJbNyx128yJzTuayFiif
caTR3bvQuyAwNRxf65rKXitEkgUJfmN3FQ16IDY/x4NZ2Q/AUlI/bf7MaXcNith1
pxr74Z9OQvjVrgoPZuyx+xPmXY44Jsu84yVN7V+TCxNsw4gqq/8Pj86f6bxPH16d
Y5+kcoFE2+PQpEGnB6RJykFxb42HY3VtoDqFgKiwzwcHFPujUDrLjxwU/dhYHO/w
SoqbRaVWe1eb9qJ24efEY4P29ZiZqstuGNY3/U4O2lsLFTSNkNtCVrmOEejimLDW
J0LEWR7oGjtx3MpoZWZoM/3H1ip78532ktSD0+6IIv1mEgeVcHz2xF8aZCEAyXIM
4w70yf9U5njcFZfXbbNlVZ9sTl+WnltnHigNDxRCOAXl3TTHikSwl7miIn2wwxTx
R5+cA8bZ+fppq7wUwoMrxVINL6MtUNuuPcTc80NXZ+v4B34WCZqGwgp1LThAiuDv
m6QzAChrVG+/B/3xvSvVx440wo2UpM3XGT8L/3DIizocY1yQBeXWRpY9Yvc8rRw0
vWZAPYpLZpy0rbX1rA/AQbsK2Eo3w90cL4rxBilr/CTUWvs5gp0UIh/p/pRmESOA
eegM+4AqbrV7ihZwL5w2BqQkVPE6ucR5FRsoFkSfoI+RZU+cKgSW5nyCSScy4Q0i
vzFE/OwGZ/xcJx+F5JEasFyutCboBh5GmTSrrKxSrLgUPRygR8F8t57HKFUA7ifP
xF/ysUnVHNq5MN3An+e3330lfpsHk6YC84f/FIOUZ6zXl79BAdksz7kgJ7FnugFK
wq9Nfgt5G16V1uHnRO2PX2O6AHBA8CU9BdQX0vdRguRcMuDPwEK7dIkzs5lHyn6N
fRNlFvsHsExd6whDe+bAEg7Wt4/RsY3Wr/zsAuj7IpayiFRdVkEBFFvczdePyw+J
+KwiYDyvr1r1niJnClq4G2E0uZMUDskCsoyIM88nk30Fwjxi6NIAQgo97AoOJcGJ
VQeJD16vCZtIBTTNpCU/KXkMPW5AzF+SUjMP178TUxORASrPrQMFbkECn93DHw9C
7Xyz5jFouJkq4vFx/I6tlT+FY/0iH6ZKnRB4AJbMMpLww0KmVRLaBMkgAL3mL0CW
dKpcZ3n2nG6VEHzorlOs0zaCBaSKhVgQzbpb/OTf31KWyfvAJCtsLnqdna90U+Ml
WqDaK0ih4LW6RJcgprGR96EEGAZC+Wv6Ipucwfl2gQUGxkFyv0a4kHMB7WJuLuNx
OIbyM7WWb5w1rw8ty5vgJwOJuT/CGBCDmlIueyPODRObsk/HwF6ewmx65ShF5PUE
FqwkgaVg4x88DjCy8wRTXp8JexPiYr9P3J1t53YSpW4q/5sm/eW+fSWuBYVFnhRj
bHNpsSF/LbxmwKEYkgVwAsvccg7UWZfQvYoDW3z4zxERW0oPzf9Ea8HDYs58DZnn
z2oZcRte+ofnwy0rKaL4bUvnjiFgEBcafcD6uK7qVU/plOTUA42Vv5CgCU5lwREV
O6sVe+WlAyjc+d6Ribtr3jo+JakU9C6DKGut9E0ofLsBXIxz31V+7Vtc++kOlenw
WqmtVRjEFPWtQgBynkKaVzGidPX/fz0frP5vL/FfX1FYeAmg9/U2iMkrOyf8NYra
bE39fBm/d/Y8Shxflb/9NnyOq1leEE7prYojRVkC5RU2+rcgo3tP4/1lENdnl2Lh
aGGE1ADmi0DS++Vd5P5SHXmxc23Cc0DowXO33Iw2B+rBGOWupmc5SXQJ8J41qnIT
W/pAl13A6oJ2XBTHu4LbAF9Dx1FloOKzfU/75NZNfJOEuUKGQ3g9qg3w0JS3ucs9
hptse1ljc6sdp0VEd3wz6A/QJyHgM81yEGtrw/bgwsIyyPqpCA7WkPOeIKGsELf6
1cnSwRHTnVqfdT70yFWy57hqPYrsBnkdFVSgQA1c0yVDC4BnP+Pb3EI+7iAsovLs
6QiG3p2c/jv2YcvtvkqgjjF7EwPe5CYX+8g/fBVv+k7dxUxGzJzsqsEU1jZLsugU
Y8vlKFCazoWvig6jxOYF2s2sf8bdlqhX/mXNhbUlU/P9D6emZted9HeNJEmupXJB
7lHl7Qp8jxL9J+2xjF6ojAewvlJIxtORSXD105y1gCcyfh6PabZVhcXCPTsfHEZc
b+sEt0wANGsNG2cJFz6GFzQ9NggX6fhRtVSrv2ZPK1ajla9s3xSHukyHPGpTZt3Q
8VLo2BG7oHPrnlSq7XWrlJ5Smt+4nrkB2xAZqjpBbaLKaM2vaqqhYCaR+t3WAEYU
z1dQGbGk4o4/qkDdkqpUc8eaH4xFfoSbotoXJohwYYnKqTshr8KLRXHNw6viC1R2
QTRxTlCS8TJxbI23BcKGbiSfWc+RqU+f9MUOC4L2pjTM3EDTx2La7UFUDa3P6dQp
yTsa2O6cXLR/OQRvQXzDDB2mlKxf+rhLdP1KI360TuSulG1qUtdzTHK+FhDpDtts
ME1yAiyvhSqee7KJtLKxYF8nGk4GSoqckym0oQpNCA2uI+ni/przjzAPRKDM9jih
O7q2+8RfkGecIqPZWJtXDcIXRRmQgByn+xbjfc7bidJJqAjrlp8fwnP7NtKd5Dzb
QrvI3wNGQv1AT1vaEXihugC3rHTq1FkbkVsxR3p03IcHz51Umwzc/JNuZnpQtfyp
1gWvQ6yjfG+vddW+6CWx26ixnufP+eGzZamuGsFynJ5p5ORBt7QlEbCqKBobgj4Y
eyKtNT7Y9x6P+tU6wFrvGS0pRMQ0UXdj43SqNzp5fjkgj2Q2Vpv1ZPI81LlBWo75
gmEXP0lwO5grCwKH8JGMOxRCtxpgd7XBSX23g43DvjSvipJdNQwyL37FQC1Yzmn2
S5RCORP93kPvdOdC5CD7ddx/1ATqNEpr87Zhfg2Uw9ziscFk5D9D1fXJi8hXMH3C
FwDxcidk9cuUylQFLQM/2YUgpmpygnujmO0abVOKb8obXVxB9QL8I7sekelst5jk
7f9r7PUCxwzHXxtGuKEd5W8hultIsGpBq5YJ3UjNv5BxNokAlUQHcw+qTVMcSY2Q
4ku+W9WL13GPjB88ie/kYttm55I2Dy7IgM9UKcDv1K2Q6TSjVe93bp+VMfgBE2TR
j0RsQufOOAV8i8stS6W8btSJVvTdNtYSwCrbLyg5m8Gl24XHGs58nHJV+cNoxQih
9k7kjPi8j4RC4naXaXPW7lGlVDCeczYrOopuyQgLxbHTorgvk7ewwRlOsqN6e0Wg
Xc5zg1CVfJE+URkl6w+Mzvprfi9sdSIw54epO8jvU/U3nTCFo6nUZGG9OpFhmAS2
geQge4n3MRbPm0FkRM2hYEUBfDo9z5FSEVM4rHIwW6BdIkOhJ5E3LaKpW9ASVtJw
+xQaUuKblkvc8sIOmGbnpW8mAsz2mD6V0ix8GaFoWcKWOBa1Ais1qk+vfzh6LEqN
W5gXU1mEi2d8EYfaluPsEwkmkfKYwQytPvZNFhx1CDLmziftVJkX35rfhogxnyjR
mi+OT6q9IaDWoAVO34f3teTbJOUtBSA2K5Q8KDJNo7EL2W061QGZUWpmpGniSWsW
GUTagqLvEbU1RpBWLU6lGXLOLu698ebnF0ozWVl0I7COCCwgVktlX2FYbBFbdBN9
nypoUmGm2/GDG9cntE5xovpm7RxMOhBAKpix/vhYHwAWF7zPaYtKCzgl5k6pv4cu
fpPFb0QjjWrAihZ3pzEBmjc59wB2HZ1NL0g+COOAeM/rZp47ZyFHM0yKIo+oUZMC
GFRxL7iaooGmHWlYJVsAFMVlKOzMthKtsTkRKclLGJRp7SH/LiykzMvF9KyimbNX
BBEGL3ne+nBUt9Kkckhhd4CCAoy9oNAbLjIMN+cuBG7q8cCB/XClfqWzgaWrh6iV
LFHEIgEejeG6yiguEmtIJV1IQC9/b8KIJb6X5SRqhHhUVKLcU/GDBtx/elgkEYoO
NuN2eUI9yKuma81lpxRqNC4Q4ZeMTpmaNs60NGP3O88BiA/n8enbtaRNSkj9wp35
ne79qQGrMuGTtyYHdhys2fIRwwlfygkbRbEfQGbYRfV35a3dAhfvzM4olieBkOMx
epHLZ0teQrKjC7rgWsrw6dYT0p23dsXn6/12rikCyIyCumBxXoD75OouCXam5l0x
SwzU7l2zC5CCmnSGk36DNslroL/fsFz38EQwEDDQBJBKoKnu0s/He1//Pak65+53
ZjKyevghReoMOS6KZoOUHrKwNfNh8J/DOUKH1EorNzO99b3sUAYn68QWYZkD7roQ
fTdNK16uth2yqMcTZtBSl9mny59Vluy1gOqs+/QvznoUxAAKJv8px/8C6cKTvhII
nrrIRvzFIzmiuNnkKxtDYSedB4pM+5SGl8Y54EXcKe0XfE8WNrc5idPRPjghviF0
MTyNkn8DBowJtAaCMVQTHz2WBWyJJwYHcZjmvtQtNsyucsvVpQrIOdg3d4Yp5+F9
IOYgXsD+Wwcdf4eLblUryw3t416AL+AFGkJOmmNTxpGJQelkjt1oemhA3x5tyqmQ
nS7H8W2N7IjjzRGd+sjdAtbZOytjeE8S/hFXZTdNDR0bOy72pnsZysQ+JNfaK9NW
/9kFlwfa6xQFUYcgsWdkokCrdc5Wtp9R6c2DxA8usDB9iYboRtVh7es0sc0UX9AJ
qt+sApB9BklArYRgZcjRAheEt0+tdibD5hSEFFoRIPqgVk2meo661cS5UVivCjXa
Cr7UhAye9DO8MKERRzdpJJJShS9FYBfKHzgmyJICsbPPk4ZDqj5oQ4sD5VPSYoaP
WGcYcd3Q3Iq73GZuevvunqxVEEqfPqOI7m15iRcs9hTvqWOP/fbVTlTV95Xavzrh
HX3PEIS5ZDORJXm2q6blfHwsdxn2ilfIosqeDxuUGKsXu8Hz1UE4vicU8d6d4Lqo
nI/xny1NSIipYvv6bq9OIbLYZ1oYXXiYfcUFZjo18VpVezsDmJYeuth3mElfKiiY
k3LX/vo1GcTyPmYiM+aseRHu0WD8V0C4juTf26nTijlF8glWormFvoeIg6Thk01O
C6bVbLKJ9EPLPIZEfrYgAPvYc5/zEJ0vYlIjpP+VbEjLTnHHTyuL64F3mgE3KTxZ
ashXe1g+HalOrqbmM2JpkTc1zLsVIp2cKFaeBNei+ZIi+WkOuw/ujHRCde/ybMhj
5YLv2e9PTrlsk8aZGQPIVSRTkNgReApuulJJ5md10DIlvMYtZm5DDy074lHeINbE
CyBHn5BdG2D80AO4b1yGYeJ+iyTM7n4pWApOzTRq0prKwx0kj1wTnvEi4duU+bKJ
AxeGeHIbQF64Horj2KJfpAf05BBUCuGcD3fsFjNM2F6J9e4Fe3Ai0fs9T6OVth+H
35kJ06c41kIDwnAJk5FQh4kNv11Tie/qAdWdyePC35dimF6csk8FCuvx2VJnG7uq
zk6S2Zpz9TZP+VT3ZsVAmjuTpQJMVq3PTwc1eRBLvVB4S3YJWjU34ALprXUERcGq
UKOBCpB5V5wa31PEJoNmXrd1M/l5buhEtzwyoJfy/BqzAKIGS9Rcc+2orjXInmaN
XxxyZVhsNpYdBIpCzaG1uyPneaHKhutTkaicPH9LLBJAzSOO0XQXXb2CIimU5/9G
UWAHmjGP8CNfxxhbmU6PAMnjqJkrV4BKsFitGdsCoCGeahIcZ1l+Etji/n2bZ6Mf
Y4Z1sMYqqGx/abhtyJvr3d9f4CK5EbtboelXqIBhCZidFFdEyw3NT5adczkbHcKW
rYEyo0vyGNrwwfJQ8h5uNhMlkCMY04WfD4Ow0wAv4qNnbnXe9cPVnCKNaNe7AZJs
k7lm8EpXOoY/HpiozhVf6djtQDTN9YjWYvGQ80+H55v92J8mW1+V32r/vVKIVqPq
Lva+SjjEAMImDrYTxGrolWUO2V9TJxKlTzCSb8/B+LR0eOGxehdr6eNDAFRcvEsY
p8VQxsY2Aa9lqvmBYRwlUYkzWsphKL3iCIc/2+tVjZpziBjzudNBnITDC2Cz1Pqc
Emdwm6gGUlip2XbH8TlNQFZHJ2YShx4kBJfOG7iSbThRsUb2v3gZPtMWZzqOcB6F
4BQFNF4pJMvx9JhLOZBhrA0Je+CfB8PFh0qqgLgIkDhu9biXHJW+7oycDQJ53jz1
hoGkwEAGQOetEOOVFshsXvDAeXqx+oUI2r9maegqmKMGAX+xQYGHMn/t0kgh9U7G
177h/tpajrgpbeil72276eYxs+zU+nKpuTmjAW7GNaKExbNWcmVSFSc4aVuzuHC2
NpKIqfPyFIkDUyAoZ1U56kLVjJAz+SmB6TNwwOYmxAbgHWtstrjGg6hKAc9u4Wee
v7YVUMZG65DwEboZFTeFsquo2fJtVU2hrZmIW7r6MWMTf8H/+agKJaa4Nz6IlE1E
CSrNWJhT2wmAktePRhxcFwd2HcCr26eVZNuB9PeVhCMkpeNAf36oxu7UQqK2Gij6
1L5CYvR01uO1sMoUFKqWAQsiUJqf1t2KWWyxU3Bxs8CVDte7ElZQAZDNB8p6R+lF
l66dSXeBFIK+H07M1fGoNsQwFC9M0vhE6hwMygrO7PzqDEb1A0E+NiZyNOtKDQBW
zhRZPmlD9qUv0a8ESWeej2efDGgE7riFf6hpDYb/woG2R01X08CVbooYvlGJjgXr
Z0TbwFoA12v25H02lAGjFIQ6Z7iACmTh1fFTpoyZQX8d5n3lXwiuNg5WJjXcFBM5
PrFZJyOrubg4HH+9Bite1FZ8Nd525hd1in9PLGJkKr+wzq0uhncy7kYhao0s07hn
D9I7/L8xayM7abKxZ/qTSj8KgyA2M/vEKGrJqCLiWQy53XKksn5TNgvyhZnwEZnu
8AUr5YZ7Qt7nRFdnVDAoUsKAW9wSk28GecsW7Gx49zOmUBAnGb3qZP0A0YafX8Tb
DCqCNvzE/38FeqSzPdY1yEciw5185NZCPBvXFtVypVOcg637GhdrKBGUDJszMu0u
g8sznq2sBk2hvO/8zOJC7FaSzw/KrNfWmzKxrn5+PvCaKEiqKxu3WUXAZtkyBdmQ
K4Mv4eHan2uDwYjXOsLeIpT4rdnqtlBQct7pZhY/jjg6wOxc2SVKWIhgeScb/KiR
EbB37/v1RiEjyDQ1vej0V6dDe50nl4hY/XAULKOqt+l6JBacdsd9daoSjnrxlYkk
0jcjEAfDtA1o303Zml+6bc9SFdchvYCmNKjWd1WMVPUMdAnKURHGAd4F1g/ZdGqJ
ekasxz6tIKK1hDSIUyb6UXTpKxB+5oxLr/gR5GBhmijEltE0+RU8zXpfMqXVKlbt
ghntCUymFTZWNu5jRHcOBPK58yRIsy/PT9nnEf2xSWjYGIYMMxI1AMwuXLzB6DL/
FhiuUxVGsf1pWHTfSy7n7bT3jcQnMyoEARH27nIZ0P60EGVaosBMewgfdvGFAKkE
y4LnmlAPnhB5Dz6CgoXP/sQyqZRbDEQ5ClUJ6p38rdj1xYSparuylS5rRWcpd/Jj
el4YJF87dFt/ZZ2g5pTmTMEy6PlQICQbyVM90O0vkijI6OwLqOIyiXBWcxZjZ+5o
giUdYh999tSru+CqHLLp0LB7k6us4/2V/ZHPVqTs1mlPV/mtRUgbMojy+JGHyugb
5w/qIgHTBC4Q6Ab3f5oq4p51pKPg1DOSiIBkekkvpGP8amGo1r47AEloRJq+xi5H
kvwGa2HXf/n3k/LcEEtYxBfQN+6cso46RW++SWvUXU6dXQAAnLwXBwpxYN484VNY
k1dV4Am8/uMLQFnQK31Z8/SO8Rz/2oAJh/xs8xiMPFOZjFuS4R7h2jxd2rbyOYBZ
TV7sSM6xsVp8xPVWKMLJd5wO5taFNm+fytcSy27svb1KENUIUO5PgxqVVw/9/yXi
1UIuNWrEkXWjVrL0/c1DEyInw0wY3hmxUt+lFBtQsbA5/vS5Tdg1q+FgWVKF0jqZ
eMboTY1XWWAP2rXH82VlY7TJLeqiTSA8iYF3wHSNq6s+Ibz1cM7R2itLvpBMp7xp
NwVfuKT4oIgknoJ7j8bkUXR7XCcRc0BJiEqefzFS5Gripah867w+rwVbw1VAFId9
BaGMZG+vqQvZV2z6OiSbStqRh8Zh54Ytmk6YE7Y6R5UB3y0oxvECk5nU8ZBnL4fs
5CGLDyom2FDa6YlQO3aecD4DVnePP264GNnKSizkRCQzq0GXNJrhzXxukQHJQWm0
cEEU9bRMtoaVbRkVC3dJWTu4UJ/P3dksfE2KW9zWDbalPY09ZFHhpTpw0+L1lakR
8mkh5mquBzQQY5mUtLxAs7OFotjAY4cC/1nzUr0ew15LIQG+9O0pK1nPb0Jx6HEZ
H/9pAdnH/gO7cN1REd73ix0nFUlGBTXfwSKRE3eCU2TqKkKnJNmtC1wzKD2BcWpH
YCnAw+xUxzE8mLfIXbkYgVc57u8RPC0jR9DN0h4ZyMj6KVZudiMFwL9UZIJITZdB
rJH4sHraBCnrR/WydKWNuojwAOY/U8LK6RDnJiMcm2QcP0JAiNesHmqCrc8rOlgX
KQCeazA7kntmjdh+fdcIbvttllc8wAdPI6O6qEwX+/PWtbHIfQ1vAFXmv9sEg4I1
QAr2kvMB3PAteqiwmmBtYePsWhnT3zSETViOII7Ml+lWxAd1ukL55L/zCN8YyzVq
bOtVNbRmUKvZF9/LivJX151JEEdEGH8khmt2XDL6dbcYWa/souBP9AgWwBFCCIws
EjJ5l0Reunu0Rrmqo8gX9+MmfbPTPQagMqOTbdMx1LhYhE4oug8EFbP1NNMw+x9E
hdvtMi5tIlj1WqwTDq8mZO87fMklwy/xYvbra86hMbqq+a36OX3oFYGva8SjFK/J
a157MQEZf/6uJDTZqA8SuSlyuOMwdqPBNfuVWHZURUIhSYWgMt0qlLqlVxkTP6E0
S8M7e+HHSs0b4HFd6Bed0cWgbx2RQCLteaHYhCQ6/RXcurudmGxF2iarkZ5sgVkS
BoikdHqZb3QeACmoylDSdvz8JeWLwX2DNZ0tNC0UuXnCJ/WX3SLDO7KbgtlIbJ+R
jW3YIEfKc/7LAy9xwQbBi1GYOO97TzF+vPiEnHvjUNSrmRJvWCMFlABksWvTKoZQ
m5hLlSnDZpi3RYrD1R2tKyv2hiqPw9fDjyz28PlT7jwVohk/F4dNpsqmVdrybpQM
IIMKrBOMnrMYFnyB+UCeuf3PLh41mjLMR/gE9lsltgHQ2vhHsC9cwsrQPYzUb7A6
I83lIAcyJRjJABBmlkdZZlGqpNuzI/dbgkRSDxNvfs38ykCdr3GG9jmY9H3WKCpe
0V1hcZmvM1CIgbPuIIG2qVRRFLcydVQT7qcIPKVuU6YoZ96gxk35U+mruBUO21bE
7pB2IOtmGivbbsFnO/qQSIldQSeYkICs7A6vjWegv3r8jOHd6mCTZHYGM8Z+vvD7
K7XHoPO+Ld/DMvdbcl6vttHTrVm0AbP1QgbA4WozQ7zxMnZ7TbQPxhnKgIsbRDKj
bttYxjxyHw0qfp976LJVIVkjnrW/zoAnbpv+BZdMAtWRslOFdRHoX5dZ5t1OP7sg
6rIYw97PjLJaIVf0FH3EGmaMEIzaCuNc3nTJAODHDQfhX4UpZ2pf74LtW5ekQTku
4Uq4BwczsLAN5XMKLxKdeAzpVlQF2b9pBwCbLkdl5bqbuGJ6C5Bmn3TFGvY3JxDc
Rv9NGvsQjW9Zyss3CQnc9KDeI6ToVXlNjI28Rn8mhXNOW4Id/BSbEWt1PpXYXwFI
xg55ZyO9koDV/tyFasG6K7GICs02gz2//O8TI3cseToW3uOFoGqFALtwG3H7qhXl
ul/lyPtYFmRtnTf58cWvib3tFgf0BiPAJIf7R9dtCtdvDl3edDuY/mJGjKZwxvyd
H83LZqAjHgkM4Yb6KiVmOKGO0d1noC9X4FHVhzkvvMIaMvJdRe+sMhONcWDABQb/
rVVF+hGiZqbxmj9loiCBkwaDsGjh5ytf3uQdtvIfvFHMzS0IN8+T6NlnRMq1irPe
tddhwesXdxNaaaSP8ZcUoDGHKixW7IIjStPvqw4Q436XMppbQ2FeGEbqngOv1JCx
y5L/hN7RfUyVqr0iBQ9LNO3kZhcU9zEx20QsHBoJt+311GiD/ZRlYOXhwC+IVneJ
lkzlRC3p+6XW+G53dB25jdWVAEJzASRUaLB0ymEx61mGAwfnHux9obMlxTFLc4Iz
RiORyBms6QaHWTzp9BnKUF7N6c7uAh0GVTtyGHGyZmBf0BbdFNg8rWAtsPL8LC1F
otFvyxsQAz7bMjLuBn99+6uKMenEXbOE5qZUlgNKt0WyGRNF0CuG3dPy59/8UQXz
JO7kRJ5NFrN9s6Y/GQjI5iJPb0mwJq/2gwjVLI+3meGnki6cpvUym+0vP3wPZrZR
X6woUiTvwc48siDJl8ngJYGD8rfDaUyoHFmoMGdcobGy/SbY/fZOd1enNStIQOCG
KQssb0lHmrfKqvCMjJO54inOSMuZDtYzpO8nlvb3MyPBpA4tB8RJ06yVZLgIJ3d7
NB4sMHsi6TO0H8s8wr1KQa/X98UuYbmBm84BryDNd0RAVyvvH5la/P/D77bkLJh6
TuxEC8X9jCGSvv504ndipRr2pxCfM9RIrWc4rMK2i5hY4nBgL5i9nZiRe7NHDdhQ
Dp0WcvMxKtN3fXP3Wpu6V6Ym5PEE7NkmK/OuHdP6RXCxOgUI6rcE1mxevYDTCfb6
tNClTLPybeZAMfLOLCrugc4vMvG49DhdNKxRNm34rduSAkzYV9EP8KxYNXTxHdLB
ybwy+dc0BeAs3Jl84qgvyuy6t76d17l5QThjndg4p6xxBtgPz1oAlhNpP9ofzzXy
3/n9l+aMPQyfi6fHiaYputZhYmJcRe21hGuU6cWPHv9Z6OVbOGICUEw/+wb7+ylp
duItMAhJSS4Wv+eavQ/iG2Dtiiri7yOSp6rg0Jop8JMwUcViKchqwooLNGSKG60R
CzSLKsNs9ChQSBUHWcYWHJFsLbrZ1DaJ3QHwfhJ48/HkzAwOfUgMvWOtZKGYN9As
/bv7V6WoiMzX0Hsfpe9H0ggrPOu6UMx9HiKSnIVchiLakNx0JldZOA3L1Zn0BnAW
T9mT/SO7RDb03czgB5M/DeLh1UQxPhL/lk9iyz5I06UM2VnX5xWY0M5F0rmlOj6Y
OXoacHqpLQFg47kUnjD21E66Ra/v9J9vclDvTG/HEwlgun3Lu6OTNaXVfZqhwLe/
JL4G5XWd0EI48sR0VRpxIT88VPkH0698RHuVMXH4j5YrGOPldLiapHBwjDMqYKxo
zB/Xt7socsgoK3QaTQXqFcdAID7WLpdYMHYCa9wmCCf9p2+XKa8Tq3v+1lvxv3KK
gEZeeLQovpZFdTZFhwCH1ehdvcL2Wx2V2tlfScDW5HkdzVKJOI1hwWBkh6YzgQYx
HsCjPR0GGILTBLK0BTC1336UMXsjFb1w/CX5ewp2jf21OvDZv6d5yroHhnWtFGwg
zhC/ZAJrl0JX5bU9dBbFtiWQOV7TpTXEkDzAVoeROFQP004SJFCE1VCGYLP9iqMo
bYubHyIAPZDJUuQ05rLNk2TYxorWAH/blsL2HvcQPVCBl+vp0FXWBFUrOuwdGsos
v0gZS7NteI6BmoCLnzfx8KowiYRSq7NCRTHv3JvxKouf2PmtBwIhMgZeD2y/SY2y
l/znPGd0oXPUYoTe0/PZqYWV1HFAMMYjwDTpDXCCPob3nDhHUt58C8eWzt5hhnS9
nqpvthFBvpg9HT+bYVIR4T30x20hEgT14qxfXwv3Pkre9S4KPKD4gBWA8VAqDfLy
Fxuy9f4ELGPa8KXlWD8Adwd+WcxfgLZ2UjztX78whcOWnNUPjHWNjOYPn/q70u5w
1mgSX6USHTB3vTsjCXntUO8FYTE++hkkYdO4xCqwN7l88t24dickR1QqhR1vBZ6w
GxVqppPU8B/tQ2kwB3WmQw3WlQS7g86KKr3tiMzVY9EANHhUFP4ukc7GFQijgEhF
6Qu9Ld2hEuIBsT3TTLMmTnqpSiTLcaNCVFGs24fSU4o749p6e7osnziu84W9Mr8Y
zZdXp67Sdv0XIUjq1fXZ6/vAduZCkOJxfE9gLzejNFZZ0X1QyswkqS7+51EbBlb5
Jn3Jke+2pqAPFFxCVdpmI6kmaxULgq5jd9XNAoOIXmxzz8UPln0lQKoKuECLa9TQ
SMQtqsTZ5zLdQZUX8tTTC98Q3e1aPV5P42nnSSA3Z/6L+XDVOsBahA3Dd/PrSCz0
7Uc4DImO8I83kTvSTfAjMjb0YKN4ZJv8E9opYUzX2ZdkjvDK78T/CSyi6c6rfqkY
A0yF0i8iQ0FNUnUy44FgbBFrDBi7Pq8mjcXsxx1pl7YD35xWdBqp2sYe7Qjd9DhV
MLH/4/L77osFGANiAVsQ+ST5ZcAt/T3muTzoZivAHVcvfxI2jahIr92VirI3BISC
CeGd/9esOi/fK80nbLkzDi3nRMQLTep18OUro/q2WZbA4TtRK6MfNDjNe2FfBxC9
qgkVpT7WYdnR3XqbZt9qwYHbUPkrVJ2eJpH6yMArBQ4p7WstBu7El9KE+YaHveTq
TpK7XF6NCkVQrfQx5UCLwyFTTAVKq10erB/FzERRHyRofXWxUJ62KRnZEM9IB3Db
r96AfxEHpqC5zpLo3vznlRu4/Js6020Jph0FuG2tx0rR70wL49kI/pRfUD+BeeMf
GlhNGbDaZncTa++ZRG6I/74OphytYI+BcbumGsZ5/AAqgVUMQcVOeXuBGPemgMmN
2vq3dhgVS4NBn4fYWMSxRL4cNNMXsNfk/54C2l+v2UBuj2GZpzLnOUm+ceJ6DquO
jEBKW//rtjHbKC6txFjUKnJ8mJkRag/zhRKUxv39oJkHUaisvFCkj6+1IR9sBgXd
yVR+9CQe5jMJb4VIGLLd1FPau/nxzQP3QIppzMkCoexSSYLVavXbpyRUMZ1Qa/kc
mQVOw5C6KpfELY5tWGWSpw7EHw68jh3eOxqSSYaWXYny965Pp2D04OS/NqDsJTYS
LhWNDbWCZ/4sRCG0PbKdrovOlpkFBqCjctHCshy7NIA/tw6IGVP20sxET8zTNL7a
0QXHQjMmFbDkHCaMXpjcXIKb3DnJPWgwIlX1sgXzHMSPJSyDbcy/qGC5inN08r2H
ghnsUIWVHrWksdLj6M9KAjxaU7JnZWQ2rsvdCwZHTjhEKfLBvMdPx4lpsrh22i0O
1aIZKM9aqwMcOi0WEwU/hjoyXez9/DriP2gYacmOiGbsFkcgWreycNVGiDYxDlC6
DvKcwGvJqRhGld2AzeTFdLumcAfqOYzl3f+5fZu/eNTbg3T1U7I2XYe/+Ph1S0/R
SgGGP2SV3Bm6Sq6i/IE1X0+0aHxwUa2Art11rhtQZwhAjnM0fdKD/895ZmzqS65E
TmpCdijD7nAQ23Cvx+NrFlZzr0IvkQVjIQdzvtuxJ0hJw902SztzfI/PiR12VFZr
9JA/3+yH2lmLtjcZk34xoZX3tzorEDxn8LXH9x3cYOz+XxkIoxOXcf7jykIPyKFB
8t2B8GbFC9eQsDJ3Z42Z8c4PWZcCGZnJqnSBwvQI86wMDZuZ96hJlSWH2le/CSly
r8JCX0GXR7843V8oKum5xqFtSCSoJhA73Nx0Fak+dbHvuubuxADpFY97oQEEnlHU
3QqF53j7eR6ZMt5BJrSja6u+ZOrOkdVuekwqxBV50gONkleHGdBo3NvmaFmBsZKN
ICYwPtbrtyTRGjXjt5XzLYtqqgl8icp271q1oM1dafz8BFSFSdd9A5hl5oSYnx+d
LE3iN50qH9E0gfPtLQn3rBQit2VA1U5MAH53Dh3FnqOxC94/Nh1O4KD+3xMUJ7Zf
+f6stMuvRXPTpitPIakzQeasmi66Rs+nZGmvoMqfkbkA2bDLJEn63Mt51poh0BFB
X/zVB6tM6ijTlDhNLAfp+VStwTKlmhRDHEc1lbC+UWAAWqrrUouutDNgDYKk08sP
Wv6+KiFQ8JapCwfgPz3Fikby2wYvs/l1aykZC1IQ/4pziaoynJ91YXwjv3Y9pAF9
Du7qLhqQRGFDz4hIWb9eUDa1JLxqPSdx5aW/V43RWB3sK7ARb5VmBjinUZ8JSmxW
u5MwJuBBAKW9IU4T8s6M1uj8jp20AL9a+f6rFVTYQ3AxHiZTyLWfawewLn9rkY5Q
vnGm4ygABKWYOYfz0P84OB3+Qc2iRXBvdAKEjRDungq8h/dsg4WTh6Q5qgcWvqbq
C7GFuHYn1jSSbXKnGN+Zei1lXOmrvuohNxBm0Jf6rYYSXzjHSJ+NCTU00vC5IWE4
MfuQe0CiFH5Q683JpJIeiEFpY+9EaZwDQDoZPtelgd9TRWBo97NDtFjvgUlpUDPu
0QX8u9W/C+qMRHmBlSMxlSJ60rZjvha7paKJOHbsIGn0acjI4n1Nbo2mn+L0xLDA
4rDAINtJ9AMXiAyhcvK17/1ExiEKm3WOGX9cwCnX6hCk3e+BbzEDunRZ2CRNnJ+W
AFtjJZS0d9IzxI7pVPqartxwSME5NUqV3EyWJ27hlNFc0sOgW7sMcm9qCg6fjy9B
SntvzGDImolz0ShBP8QZScbSLVCor54MjXLQkL3hsGt+MSokMrXUQeLVOGZQNmU4
+Kc4DPi88IzV4+w8Taeby79oPmgAh/llSUTL+BPhQl6atNBoYF6/80iezYHQ42Yn
wzQHFfbkLFSnv4keEz8/5NdQj0gATVlOWCQCvYfn4C8FKcj4V8HAZAmDsvbrFmG/
R4EvCF96XdsoBNMA/yz6QKQ5Veri2bm7azAXiV5VjeW526rcHY4/WxsQks0kGQ4L
29bdCGWuAwModlNYYtWCREbezWI7fQHrBojl6r31TbAAU8EQHTISftlrB2EAF54d
Xmzz7wkpK4PrQa+zLExf8iQlVGOLG20By10ylsWfXPOd4J1G1kPXLrOg/o5hrxh1
W0kTqMnvRS0/Nj/VJITPQIpTxT1d9Dc7AOSE95luUjMkf0aG2XV8wmrGylFCQ+St
CPQ7RWjoYTnZytBq2bebzvGcAN2i3tNCg7nKcRWwaqRFrs2wyZZ7cisjA4tUSNdx
sPdAbI0N0mOEJtOGrMbqBp1W8C7kVA4DKuVOI6+rWtz5EHhqanxMv5O102GgVpQV
NEEIDj6mzDBmQJqZwzZoRdPza0tNGJFTtDKtiAId6IOcjY6vxgiY7KR7AC8h2OI4
P7lhrxUpI6task4Uwa3NS3XdyRt0HW15KYy+61//3/LmNkSzAKnJ2r+WS2LNh1Ew
1n5dC+zDzFCqnnypdHOUkcdyPsM8pX2Vkk7eqvm6LGgl7BEhTdKnigrpg8m4POtC
BjKCRw4w20kM3D6bKCWrZxTpbZa0ryQUZfhWtMRQd0JKlSYmc9QU5ae/KXnD4Vp5
EOnuffNFrqqYqeBnw/57Pm6766xm2/CIGLyFzNOodoTNP18SNj3iHVx/q5xbtw6z
FZ8UYRsl9MXNv4b7+TTCMKCwY9aJVHDgo/AWQD4SuVhg63J9Kk88t7ZZzc66b29Q
VK9IXqO9vfIEXKmTgqgLKdw3CwDHb/nx3DValAdu4B5MuFy43CKn54ySeIAstvPo
5Lzc5qglt8tUTHSzxdeqCAqTNOQ4zw02mNAI/CheNCYgM4BeTotfzWHdIfh/cVKl
BDF9/2/GggFTY9V8as5nsNICzwa9/rgsPg012xgs7+SmYJJjyXY6+CtaVpJVS/e1
sVQbxLHdQoJ5cTgXChYKLaNU6AXJQC842+NA+nDariz3z3FczGvm76IKqM/80FJv
IoZ7e3lwVPAxJEkojqbVEJbgqdRvW+QhnR7L6qtV76rKsevtuHE6U9r8TJSjJVQY
zW3tWZ4eH0VUkoar2xIuLFrTnOnkyo0vTJpCxL3PMU5N7iP8YOGX4GMAco3TJPXH
Ji7YicnzZcDwnv7su7kVz+9fN+W9bc3NlRaCgivAbWzi/K3v6PwlQnb2XfUQjtBN
GBfqC//KEkJLAUyUV7it0m77qTvJoru3khCPNeLrigciNuPK+LS3FzMSMlvtxvnh
A8H4OWA1I9iP/uQNB1RSw1IWtlgamZrlcoAJ2ydZe9NTHrjJyrM201nH8NWwKMio
/765TGY4lHU6P2I15xEmkAw0pNryCIxoesP9sbg/sG8CtgUUxdmXKKAxJ+kgH0R9
NJRl0lWjjEzg0uyI6GA759zgiBK9EgcX2nT6NXLFZ7Z3961k2eeIBMrtpS7VWboq
yPgxeUeShM+pmNrtI3MerEY8p/0LT9JeFcNNcJ27vJb6QBnBVGOOqNz0FhmDN1wq
oqX6FRXFcV3jj72B10QMIX8XnFhKs6JMILjmi+8iTMiVaAkGiI3QuGfSz0pHhhTK
KToV2FYQ2/T5lzppElV+o/pT0RX6QrbOb/cuZJOs4OY2id++6J1sB2UY7UBOVcSp
yuPYmoeK+CLQu+gMKq1mn8jhyO3aubsmdTUvE6rdlCAJA97qakMlPpAVJoW/8XvM
YmbnlGQ7zVgRaTUYI7cm5pdX/M0nCwniG8Wrm62547XYYajdfi96R9xXVP5UBaSA
B3hlu9kpPAyPSut/FrKCeL1YXDj3GGBXyd2vNMVDWhrPw+uhtVqhv7+S1G4SoKlw
PAjH3WsM4Qhbsfb0iTnKo/0dJEizqOpyQ0iV10SdrvAY8wZsAG4UKxpFjZMH0as/
1pUgjB3/OEbRQwvrcymFO3dHABZqIOqdhCMMQOAzEwqNIZBP1no9ks050EBQkjwu
6eiVY39X/itLBSElgqGTTKdnUQIshYsMVyAT0i85NwT5XRYWr3+n73FtmiI6p8An
hJy4gwb62qKcJj82b4aUM8gsoAXFmGh1hQxtxZYihnt2zLNd3S3M4mIVi8cWb07n
16DNca+otwHTc/0CFB3bkf/hHVjytW0VpqSesToTSBGjFVroSHDgBgnfP6p+ghqB
1NtJfiFnew6sgkY0wcdPfIemx1hPNQBlt2KYBOQImAo8O74LTCWTyRSVWEnuR1hz
eJz1647V3U5KCJfxcwm6Piu1iYPZFofiUJOoNQ5EyObCI2WXma1Z977mpQAMCs9J
41K4sG4ke+ZymaWu5a/xLkeMaserrrMMGgSbHebCJMLAm09TD0ics/E2dDb4Hx+Z
pM1xqsgrtPyHNX2amM/v8b2mnfITUPJq+qcSRM+3RtK1M5kf9OxihmNQifj1llWR
OlTZx3vEdR7cqXzZ4NHQKcKcuDvfhJt3pj/7c6fQyATA2dnmuj/CycMmJ0H1vQrl
ZaUhF1hdMTUxSNdv3D6YaBuxYrjBkQea9ieo5Nju4XTtZlRUzaXrM51GHHzP3J/S
ft+1f8fdte480rzuksInDbBkOrDylliu2M/R0B5oxn59nw+u8/JS/k3yC+mnnGro
tIt0ranZIfxTKnrU0769jB/P3B/wA7ewUzk54eaxRO6PY0EpTSy0g5g9Pk6SAGbP
2rYmptjmMxLW/0YO8AUXnxsRxxTgaNf0D8L6awvJvHu2aDLIyKIvdVOSJCgpibn8
+vMU4iu/0Qz4f5Dvdgl9BsaOhLIg7eQTFM+xX3WQDr2QvbLAJvdv4t4j3SzmmFj6
ow7nSARE5KNDJXl0AKJhFTDCh8beCsGN9yg4ItAp6qT7zOhW+Q0L7xh6G3MRXDsK
Ynktctj89rYRFyUZSvSdlbCGhCQUZDUSoqPhVu8hrXvi6A+cchfRJj/iq4qLTN1R
sODO4bb6/XcVlT6KkL5FcAlb9dwp/KfrHGIRhQxoau9/yskOZSnOP8UkcdnRwEPY
BI9JmeyFcuLY65Z5bMf/c5hzjouxtYfdRx8L8zWF3T4qMZFIZCwKDhd1TXqySGEH
5kf4/PAxd4bGIPOPUA2YikzmX5N1ARV9w3iitvwOM+bRjgu7zJcj1JZdL3SCU+B6
T5QRHnEW0ng7JRUh9FFJLObL/1LLOOpfX3hXCEKVFmZm3e1i288rBb/u4qwwW6E4
fnaQKY9gVFumQN/P7fKiXvQcgnabxPY03r+UMZKgrk0QGxd6TByjvl6X3+mqhe83
iNKhQSMc91I0heZbRf/OL6PnTrnPQmLSNEPSW/p/y5SCglL/a7C0F4qdrjWi20FX
51S2mNeUeN3dQTRovV45RoutatqhFyOyFGPSYPXS0J1B6OjnR0KEN3nW9hT4KdfM
7yEql2ORGhgI/qhiswqq9eh0aW7OlmoI5hyzuECyG1PdXcIYw62RA2hj2+G8PJ1m
nMlENxyRFnXqhlWVg14N569+vKb0YNhtqkATW6/xKBAqpxVOO+1cAa+Kz89GbB6p
nRbBzIrRixXgEg2vCnUX82yGxZsawifwNZF4uawNXbpO4AZk5y8IjDKlZaLaGfro
3U0F6aAL2qclypOk/hXjtuY3pna2Siomt5yb194T6MGerKtY+TrFXJmZ1Jq8DBag
Fw9P2DTk9ioO+9wm/gJYsnf2iWjUMlTH9AyXAveqrw7V0JQvGSQ1ig57qOHTIMRt
3QqGl0kZE3DSlnPfuRN84pdvRaQJyERWISIFkHqF25f6HtcFCQ2212UMZVzQoKYi
Ej9uJbFf7nab/07IgWx1ELPBSv0HtscfRq0DL4yP3zFNSzPXw7RT678vLwLSb27m
rwvxrJIw+Ctcc2vx3K/dqp4+klEm3JOwC9QNck1KkpvTCdT2ZIKr08YyfJVWyGR/
C9EVzdratPM5PgHHKZewn0q/1sgAAqlErUL4XX9+ys7bQHQFtK2rgvmkFWmaxRlz
wKBcP5TTq5DMpUx/wswGDkr2Ezia9HKg9IV8WNFFz8Ui7nB3DAXnGTspeWuik2YG
uLEoqXNoDCwfFMnjgCKOBrHmUIF7iKpMWYrx3Guf8oUaZil7NB2t/5pGEnYJ+k+f
+nyQMn/EuwjVGokpRGOsfCllwtP0JV91fgZqG1gMPiXVMah6RCijeKcve83YPD9W
CCrRqTdNWW5iLuMOYIA6ZpAJMmkLKBYNlFuY/tGcuavMWlqyc8TPoWHvu6+nrDLz
SKeLhZFpPEBvwaR32U6cH3oKsAF7HMOBGb60nYp91NUqAhwQBIb0Skbs3uzuIZ4q
PDPKP2k8u732FuGTCz5x3I3gpflEu4xnGvPSfDFw5T6HDUBoqXtKMa2QL4tEJ59p
vEDXZXVxX4b8iLgCieDI1aAJqMZR0t4UUFOl8by44OWICpvtaWTInkljD0hcc43q
Ld4wurMyax2PlrksEd+ODKPfr2b+1App+z9uWyH13+KrbTGzAxFU5QrHUnvDY2ja
Xa5hCcyZGqjILRTEKNUWXu6VuwdykjHfSsq8fZOEFIBJ2T3d8K+cqTVr7K/UZgM0
mpYq6+GxzkJMXU2d2oonXgO0LrVkaRd3SPWlPUxmZ+Mqp9S18cjaKhjT5nBzufKD
gUBodzVqzEOlxNrOAvOVdFg71NbA1jZ9fxNLOrJgzpJVjMyHAjIpVlk+YrRfU6D1
HCvBjrSbG9uW0iLjWb8ZR8z/7+AV+iVSaaxL0/fdIBCqC4jR8H9A/2OMzuDn9Eqm
062pZUjy3ygHjKXEPtgDyyEwCYe0Xt2rZWR8i8jOf1FK0ZiPJ4pjAGkN9OpHQ5fh
wyWKDCUbjOVtDiGxNOdY6CIK88uuyhnP2t3XFwQwb51BlBhWhyykcVmTKzQwf96p
gmyG+cikRLFXWmNdPdOdrOkJPR5shIhk21I/IdtGE7epC9ARx+77ib6GV7/QkSzt
tgPnsQqyuxyg/b8dzhGqTJbr0xdCM2rjDTkKmHZQ0Z9jF9gHDzaBsgDj4C+ZDstI
Kwz7RfBM4UDyZZHs+cl1FTPrQG3HzTTFfb6E6nH0aEfr3JRrZSFMqHQt8FMYreD+
z44lD5DjWAHkKZPdgTNnmxffvrtpqNmpv0uFqCscGOHf9dPKnalJHbpQfy7L0i34
Erdq3JylYHZR4ASKB4/RbWclstGyoJwBINq3jgYGaMbhMppilwRYd1tTVHmqiWz4
VaNjSE8CbA1WU3z75hSqDxQ9NgVUgzSUZPzI/26LJyRroRQN44FLpiVNMsuEuMRa
pBn30vEkADEpy0+ldf3QiMoYs2Q/GJ0GAkURhgiPLGN/fzfCr6pCW+BkZVzMo9BX
+dlP7J7l57fqUwhI66sZ7OiTFd87mtiLF3tle8BjXx1uzt6BxtmT5v/XE5CCoQFt
xRWZVnFfNxrVUB+VH8cybHCtAVj3+g4Wymnb2jeSFuFOhElzIZRBk0Q30P6pL0Fw
RAJFx20Yw0XFSR44QgotDv+DigoOuL7WYAqqoUscSRjvxWlcZmvhcW6mEtGNysw8
16uG4cdBBDxs7bKNARwucIUuDgH5QtLcNqgXZZwMhNLgGIuYGixFCXXEgoyz8KZR
YJTNdEh82TqL8xSfCAL4iEJkA5JSFOGvO7lVv+NYsT1bVMfOi4Y/r7VQh5O9VbGh
uOMPorWHh72C53ovo+Dn1ZfkTvhMrEf/NiyNxVYngYVC4Kb0XzQcQv6OCQXxjZ02
xJ1gwg1upL8tfqlaVJ1v25gZEi6QEUHDPFcVhZUH2lm9HVMGOpUUia8Hr3eWpMkK
5LZxxOeN1OYq8H7A1rSd+7k4SiMV/QFIdceX0dtNBqccFxcAmG/zIhmeOie1aDST
Xw93A0FmY5E+U6Ik7oPDqmG3I2mI6/FqSZjQxnQx2ZMeay1NCyZKA8JffN2aEYIU
LJeDhXrm2dn4ejFjnYKXOZN5UJgaTIXdBxSTKHx7P/+dNGwuVHrQkMDTTpKrAwt/
M0oYwcjfwysHN/Wh8vv7AXMLR2JSOW+D5uHkB3FHx4l2dbwcEt7f++PH0Ot567fN
3FHdUf7t+coPXKzFAuX4iLn3E6y/om6fBfJXS/TFeQ5NpWoFy37s9/vlGTMbDVHF
1QwVTs4trLpnRO7/h72sCPw58xcOqVOIQzd2YK1TrgQSaJJGPI3DjyyNs63Zt8Hm
rUZMIk0Ed1aBgi0w6TBdCx8g27ZjtMkAQh/81fOuVZmC6MX/qpA//S6cqIMmLowb
NJpN1+CZEDHEYMvhFkeejjcbXAMKflpcPzZKmleI8P5pg10ejRUYWvY8FSn6GVVl
+Nx3CE8Rx25OOKXQlQdKqwr8V00WgQeWCqXye7buyKgmpP970zdoR6GApmR+fk1m
NnZeWDGq3kfi9BwGmQLjczvMJWFbd22PwDnoaBrK+Z9s3dwaYCgbCy5VDmq1dxEe
kuB8PCTpngWUbSCnU9HuLAZq8EGWq2IqL8QVxy6an4mi1SYv1EQTv91V0v5fIegB
6FtGrxdT4ewxQEaffrnb33DXFd5s05wQkbRLqimqjjMLk6LGC1rRUfhGMPTMpzHk
e6DLpe2nz2yTu3OjCBng9skrWq6jz3I53JMGxF3qZo/LyfS2MnjO9Jfy0/vwMWk1
y2pkFICYJ5vRQceGMDwOGF3ALIHmTvY0izXSmbJ69Hn8KmLnDPpeqG69hEAgUNHl
eXMP2Z0ROm8eFCdb0haJYmXn3F/ovYYlL4ePVU2xd3DEZf5U7eFQ5RnVbDUlQomX
OtS9reRv5aPy3oPpwvq/xJcNmcz+u8f6UQ3KFEiAdH+ZCUWA4sJ4jLitiCdLEa8E
KreC4pdYvlHitrUUesjjOfj/wDCm0u3VyeZi+Le6NRcKdUAkDG142GKcKz12tkE9
9t3T6nTxAC5NcKPD8J3hjKJXdDdSUtTu45Jr2z255yLmH4DInJAb6NDex8jxkDYQ
Ngdf6bwlObz0c+9saCyuo+PyilYh7AD3tdeJ5KOuG2vr1L3ZLgQ7VJzFNxBux8FJ
rddLZ68tPrLFoVqF31V8dCnFcF0hB5u7LexJx5DiFzkZZFyN4WI0nMLdeRwZYgXj
sQCDt3NPM3t4mbwEikS7SU6wGz0khVyLhxZ6wtNdXgVSBJz/4ZnUL3SxNoxjVIvE
YhW+ENgp1JCxItneB0r7GjUaIGukMOWG4GBRmWu37d3Hh7dx1qo1clYrwzdjsVi0
i7aOg42klGsbq69EP8vQBKevqeQDalc2WRPCsNUQspQXZlCHxED1U+gY5WMDMQE9
3zT3Oygo5jaWRQuZkhvDO+8myCmVr9EcQIRnrLSm0aFzwN7U1MSl6kTM/cg/A9pX
mOxCUihec0UBYZNF20ZIAW4+mpACiUTpY96kcmGYoJiz6vwy3HPRp8c9v+MaOc+Z
QVr60Brkt8n4PqxF5TbXGe5mA7hNcDnvbHx0GTEE2etk8DG3fWvMQQNJzWNyPpz1
lqI5JEIVxeF+VzQcxi1LualtwX/GB/m3bILHnLlbgaw1whVCv7X7MnJR8i+PoM6b
AvKFN95thvd1o7PEZkQv0fkb7/7vBmplBBLkya5xw7CcW7/Ew3l2G6mVlY9glf0V
gC3brUn1d0r3L2wCBERDVdvjAhOBPbr/4iozY2IHthPHq+H5uzXjMvypuedDwWYr
0sM+Gy7tfF7z6DLH8koTgsKOExJjSTWKKln+pllE5IUi7T1FM/bxUXlCLwBe2btp
aVFfyiFHgnT4CaAFhpKaOlAVOAVu/vo4rmPC0eFcLVdHaCGUV6B15etPQXRl7Vhi
hYIjmBmW/zs+FfZQjssQk83vLVfMe1Ool5VFLaanrL+V7wWGbDjdHoSOi3QtlpSd
rFWV4q9fEqSapB8YLPxpTEwfNSCqT/mW6fm+uAQ3CVlKeowBE2CRABh2B9Ba4oH+
BSL5vHo3KM5hxD6ViAj8oAkFD35Zkv0kgzz9RrJ16ki+91WSsHioofclsj0Bgcxx
H7gVQydld57WfyQd0SEASvTWZxLHBJ4DnvOAS7LU4IUOWFzd5WqeBjRKTxFcWrm3
++G3r8fJ3/hetcdxgD15XBa4HrsAM5QE4fVVcmmIDzyKjdI52Arf1Kck5ivLlVHA
rrWJ1WrZOSNg05oyWqVVzQUcm39ZFyaihIO8HZdM0LoNFiuV8XWFpWazJJP+t+y0
/Y9E5UG0Bo+18Ex+9FqjYsFCpK0nyQBgOZ3V0uoZPAvma9PMc+D9OpLFivD5t3Jo
OCniRtLS6YKZLUjktCus/q7UKNC851Z0IWWjZpWbGw1gubnIOwWLZPdNeeFkbXvF
uPkktDcx9l3kJ4UHbJgdDDq5E1Rc45Bbr6UvFoptqlzK9xnf5x+KIHvypEwgzfwR
D0dhBMNLKRVs3iUHltgaOQWfrWzdNvHnBoqFLvx+Vl9bXQgCqI3tGfulR3wtp5TL
1pisPDKlvfFeU87TNpjh8/zC5bz1QMCFg24r0MH2umJ2a4ishSWYjBIqNmewUxSk
UXpXm3Bk4IkhytTEV/ofvvxBIq5igO0e/YlrnjYECziupoLzRGhba/zzC3NeHp2L
aC6fNjQZuI9O5osogqjCphE+NviBWxN06gz73NWpMyi6iQoWvCcEnzRycigXlQBr
TsymXyavs0xN21hLRO8AqxVluX6tuC3jEg5q03lc4bVnblU2RQ1GsyiA3j7MlQAd
TJcze7l3oWhZcvsFxBtCkYOce2CXzywgBqJNEJxzxQ3sB6OE8WQ72WCs8ZsTXeYW
WksKBJw0qnFN0otCvAmvo894UZCS+K+Voa8ICewQAVtffXU7qg6mOpDDxv7J+Z4G
b4pcherb7Km2sjHswmJipqwO+GalJWyU5XahUKGkKfaE5gp7GdMWhdOc0TcDHpOH
97kI68k7wxPketYbsg2i9ln4l3qaUibTqfyggkdwvJZMyYgG5Ignhryujd7s7Rhe
ZGFF/GbhWVD7dNMHtPJbz5rjmh80253qOOH5NU+Y9xCFO99cBr1eVjWNiBkmana+
Y2KnsYJYM9gwtCdmuK8IymRrPod/GNGOcg2TjHq9vkAGQDcZaYMPLSQmgsu2V3Ad
xNg9DUt+7f5xlgeDXnTj6bn9eEMF3s1Veeb3GkP62Cw5oTPX7Atu2xYAsCe+/N++
Omj2/pzZ6RdWuAxSso4KPcOz26wLfUENvY01NOav0buP6na2KRvdQByGTzjW98wh
ewmyVS3RE+IvowA3h7OKiUGP1u1BMtgpRP9iU/onzpuSW3FywBt5/t8KaMyKmD86
yWGBVqCuForjs5+N5UbsPXLGL7u7MqqMdgDdQmLVOUpc9LvIH4JhZCkntasHBTuD
dOouklzD7HSKXBkCu9TQebWrX1yaFxDF5Zy/McVhH64/mEh1qS3fK18nFeV2PtmQ
Q8oErGaPogd9M2jktjlP3WZq7uy812QrDoGW/2wuZC6Ou2t01SU/54NyHVm0ppjo
daUbm7kwAJK9vStOn/K1eNJUDRgUkTnaP4kHtOukf1YjlYGfJFuDny7qWLY3lvPA
KIbcpfwkOuAmm/1C1j3QWnU5YQQDE9K1W171HfzaWaHSJAX56ADeEIjRoUINg8QR
ykblOAeF6wIJQcUqF+rXVR1waTwJe1S+jPbuux7nPKFsG9wN4VHXsTOAxTPt4xqp
IMrH5rZsoXkjwnaK2BQSEQv74MVYES7AZ6gU4kExv4tCXZZpPJlZ+wjeGuX4/x5g
TAOfXqFNlIRRVqwVSWFGp+w36DrmT/66OMIyg0VNEuTlWV+qHpNSGkRLY7B1HIGB
1H7VfjucL0VuPHVxVUNmHrWQ5Ocy+lnmJnotNusn//wCpTYW8K5xdbta07z3TrEM
1j6gz5EE1CYLfvJT+A+IYE4gU2KqfeMFDsKfMT1Q6css7QWLvtOSn1ecDQcEPze/
1FPGV4KRTYjfqF0KuJeOWJhubXtLgiKSEaMUImgMpmTjMKhjl0R1D1sPkg65vkDy
xBl+/UjKBsgFhoBim3NSoU9VTQP05g+TABu6NT1MbQQx675t9nj5cet9BKw2phIV
pJr6MR61zQPr3u7zqohsWykIbOCFbLCIi3qYL+Uo36fQYXUNTdh+VyGb0+8CNeQ7
qWbKn8PbAOVOvETR8n/CkqRFMY7TKtT1Vee+l+aw/80xBYYdkFFcll4++cFbzcEo
vHVo22d/vWBoRAF/NaEWzS/DTalFQgKjSHI4FLEM6Jlg6B0lwpQXkEhsEDG6rOsF
i0V66/94M7aD8aGivma5VbGiB8pdWZArWRmrBkgUXDY1Dg1KcCi4ytCNYNYLLN+c
dbegpes7M39+fxBMRyjxlVwaC1CN/tIH2MtSi9YXqa8QEPv7tYUdDdyVK/6ni2oT
R9NMp0+2e3HQHo4rwgHVokhO2DPY5fF/iTWZY9TaLElK+Jhsz0vlu50kCx/LYwMI
aV+XYkD7VXiY3xskQ3anr9c/TZlaOtezv55Ua50Da+YXzYkIASDKmZHuORrEY4vp
CtGvauQUhEc/6tiuCDOlPhGkx+tR2fZ39yl0p6IsR3tgOALGIfxgB8fUWb+69Yhj
CaTGHsIPG+96HbfisGEFDry7pfEO9hVePvkriwh675Gy6S5BmyDmNKDVaJqgZOQS
yeqCt0JRLnHANdtkOToagpPL0ACMtUd2UN6tuyU0mA0G2/8hJ3A8x+CoGCrLu1xc
X+fuqi3tkkS7sGxGXM9cWFJ9DLGB4l0ygMpkWi84qihEtPXPup1YG37iWaAM+ApF
IVQH8tF2o3PbuVIbcZi++crNBJpOpf6Z6mJvslx23JTmSMlu1DRrxT2ArwXVfxaz
d9hJgBYkPt/R2r+L0YWsZOQCIj26yOsyIY3vBVRDSMQqEWXSsDMR5ezXskJi6Nwo
1ZxfXpC5Z/3g4PlGY83WYajYpDUpP+faOfZLg+TSHbC2J5Kp13pbqCJtlQk/OVaZ
Vuh/IoDE8ia5wLhG+7XviMgF0aGoDubd5+VY/HLaq2ehRUY44rT7u8NYtxhCCQsP
SwbHTOFhEASCu4Gy01BsRpqCmekVjQ7/1gOM3YubI/bBG9vOCgvpF8scP1H+YzQP
zbyMeT+HbNlp9eswmIntgrxf2DU3vkZDtrTGPi9pWciXL6Ke3jfYw3qrFrL8qnzH
JymeROF3hJYO47sM9wXJl5Ug94NqGq/R1t/P9hemgJ+pDQfovZ6KXCyJ230btZQN
q7oF0iLLXdKjUcPN/9O/i1Fx2blUEi0U4X+mKF3WnaVPCXkMpC7t75WYRw696omp
oLR1dqomkVu07Z6tA88i9z1KPAWQHonTvtI/oc4Qp7c9/U2ksrFM+O5JbSrvSica
yf8RKNQ908n028VMn2FHimzTr93T76dBjqK1Z5AmV1n8Pj71u9YcstgYx1ZZgx1i
kprh61MrQU0Fy6kOjLbya4+0jIUTTiJxxxNckZrC+S2DS3RcpC26rEEJTVZJqA9H
137X9Dfw6uBzV43FF+xzo2b/k9W8kAeLKJuLTfsXB4qg2ZuDx/f1sTN+7qiCwy9I
pf1nm9UpH8GbL/OlOpyw0Ab5Bz+2AnlYRhl9GsAfdgCK4RbIDokkqSxwmbi8YsIN
GgtXM89J/L2Rn3fbnYppNnb6N9EJMFQykYwJXKR+6qBWvch6QmnT7YqgxBOudF+4
/o7XOzO9DaRchospN2IvZyOvrI6w/LQzmmPLflviFCK9fCkWkRXux/JgEx6OTlP5
ZZHVr8xbUJGQCVRTde1JAoGSufUiP/SVVyYOSvGSm32r5Vx2od8zetQQFZz2ALQE
mvKEgdUlMlYQthXOd5zxGTiWGaT6Q+hoDC6guDMMkPSAFKhXg4ewomqDDglwwR0d
sZGnrzjVeVThyC/22Qq6hmpu7bKGGfxc60x4+DacWsu40gLxXxqA152P1IZ10kTm
5E335h/WzAv34X875ZzYo2S/3tIqZxWMUQTindTZgCujXUYPoyHxZdfcGE9ApGNJ
3evrHbk5GNyzVB9vUY17J0BfSyrBj63FY2g3IAN6jITISl6/cXW4oql1khZD/DTX
x3RuLtTqU+F9AJpoNQF7QTFEn4GTvmz9aYtS+nxAPoiDtZKQ8wco843f//AWuRjH
egmyjKJ63kHljHXZzGU3DgA0fCd44hElEpK4B6aATmf5pbyGAm8nclvblBs0b8Sr
g6OiysfW/urDQTrqRqfOqCfnCLyYTpyiEUMlKQPo9Rd0IJgoXLhNHCgaTO18evG0
AFNX1qWn6f/YMj6gAUjGfRPus/sxVSSXSfNo34u7ejM6kHjCTnC2ijNHC2DdCY1p
p7YpQuALnNx08YiCtw5zcYURrdLKTUWleaxsMg0ri7pX9yNl3YjXWrsTlMnnlckQ
ONeyHMKPij1hh9/ylmmuYLC/WBFDPafe/I7aZEQeHBKn4tOak1vnnAZXQ9slDNRC
L38uznvoZWlQXXAt/1EXAbyiJ1RuQzsekq4eK9SsV9F0gf7YKIGWGmRj3qe9kCeD
7803HIVcxbo++9Ux0g/273ArDy70lZMQBTwv7F5ML2BcsoZswvzloqNaX+f9iwfa
UylxfBMjfOlZzTvepYfpO3fdyzqVJRTcFH0C//PqPXWLLgNu868MNXd2JZlKeh42
4o/E5Ut3c7fj/U3zU2axMNAQ9BnDnXg+OIltN/VNrH9moosrvTrdVKGRC2KVWY/h
CGUsAzXLzDIMS3nOyS56TjaO/kONZQvhRMmcVEcGtPKbyJKXwlrVnDd2QeRbBerM
1q0kiz7cMCIXbbXmXyg8IDbxOcYe4UM5jCWaKI8f8dhG3NLauwtUElajSniL5Q+U
QoOLSwapKg5+fpFP/a0whvDSrD/V/nG/S7jyfQbYFx0zBFd9b01EZT4WN034Pc2A
U5yNRgGreXQI8K2e5AgRmO9q7sLjznGrKwzfgPYR7SqNabvxjCTZOgnoJ5S/LDVg
xedqzNgdwLrNZ9qndnymhhDo1+7bHwm+NL+dRphUYCTh3CJ003359QKZHUtDvQvG
utZRR+h2+ycM0m7ZV4CeAJQvzFdVlPSwJtI0kqPWhwZfq+2G/tB/n6ENjKf2VcfR
QC9cBqU8q3NkR8BPCtgNPp4bj+Y2ebqAA2SdklQtjnxxcfJAT/u/wOA6Urn99Q7A
CYyvsemCB7AFRI3nZ0sgMhX1KWJ0k/1tajQ8StYcNB8mXR2XpaH3eZ2XxHkA5oKj
uWNDhqnl0VmgnbZesg2b7O8cJ2qMS/4fKK5nHZSPavxsN/5BIFYR71ovvVjivzUg
FV6Bk3gq2pae/5IctxbttE9ugTsV2pFLlcGj37qmlJUf2hYwn3R7QTe5ouUX9sXb
jNoeL9kujA+W5zXy73YNfkZDLRjODWtoN7hQwbXlxoZnYMJOqyG5LH6DLNUbAy2C
aG7O1UCf9sRSTKZQgxmXRmHqCOVaxfXq5dZGST9keaMmQ4UT9sPc0LdWJm2F9Uic
3+wywoY6QpIIq5E9WT2eFWLpJDL4wJhLIeTz/2WuMywC8I1lq5hcU3Imi7HI7Oba
HPCAuggJ40f+YhW2oHFcb1xcGUnfq4ENg1p4P1qXyGkfzWPvV/BfUt6rkZEtHrwF
GcGnYEWo8gcdWqLSHLaeBzI1Qg21M6wjtxlHfuLVuZfzVwI+erDvhGFpNd9WfwZT
5BoJ5RglSS6CoNotqNC7V3grBqNFvu4FKQkNFH/17DTup+IVNALb6E1mXnVDcXPL
CJb3En2bG05vAtZ5q/x/cfwK+MCmrkrtLSdfXhe7YeSz/x43hSMUx2GJqTipo3+d
h6mh/sKXQltylX5jVWqZB70r8QCeTQrjK8Cb4oUaRvp4I5YR5mBcE43LSfLxHcwa
r4KEhT5Cuwjee3ikH2yVgV87QdbmuVP+qOUvjm24oV6SF0CYtGPIZgzZMGcW1TJm
zDYYeDKGbyRv+ATjjGKuSwD8N73cU8it2YnoD8PtSeN1qBierLOZYi2Nm0SYnFkl
+O5tGZh0xrA252iW9BqL42de20LdTS5SAlhLpSFowZPFbu+hljKqRWQcbyOFS3qG
d1XO4pPE71OqRZ+sSdyfsYZVUAm9MjOzdNw/9OL1dtOHmw6+S6QzaBeFRgN5fjx5
ZBooJEPCSW8OuDwTVO0OdMj6jb+SCS+KBD3Yy5lRm3JsRktpKogg3o7WmBlAXTyA
57sTFRFvdJ2Nxtkrf3T6XiUTMRjKyYI1SQbVhmydtpgfi732D5FinkcCZezz/GE7
kPkpxwnJNAxgYOeKdgYYvuRTNtxJjfbUqWQuHpVOPjzTVReiYaN2btt2PtGEx7Na
HI3zfhGdFoOWAaUrLcFB1IG4LDPW6KGzKFSKr14xRf/e9EawUsvTTE8WGZs0iMeR
E9FIePa+pFi/ZrDyTRl8NhCjWBfqUZogoQTcO0TWTrLmXZYwmCUFXlHMy8zAijM2
t6yypcpx8tYAh6aC5oKamXCcco2Be4mv4CSGKF1RnPcUaIjv6xY3GSvTGCvcjAOy
5nYfgRWBWDPZFWZ4CUb2887KDgwzMllWVlr60drEJCXxSZaWKbsifqcovBKUgVpp
WAiMLfrj7ogEaEJYugHuj2zeegPm04XPjxsLlF9U/W2W6b199sENaGs91NVw9CYT
raj0ciA+53NxCV5UvDjbzGC9s5Yn4rPT4Gi60lSe8/SbiY73IKQsxecN+dLywV9R
zQfNZ23DlNH3XeM9Z3KyFvycMNzptKqVwPCqWwBmFCniBqMoB5FmtM7lg55a6DJF
iZM3mEd03DfNjqZCJSL9tFHcggtcWcbKtjVDHWC4s5KOyyJBgSuLuPyXJz5nBK8Z
5NFPPycT7GRLk5LZuiWoTJbtr9NTWZmj5IKvfrDry8O9+jrI7sQJuncbVwg0N9v3
sUvy1GHco5J/zZeJHgh6yFBwmMwgXPyIES0w91jKoB6ZGas8PCW0t/cSnZ9iJXCf
Cucrxl5FDoXYnfVBy4+hIUUmaSThjQpTU1E/AAMJiQIMJJfVXZewc3U8A/Y1/sgU
aoUc8TUItTC0ctETNq3MoOhrmbOVy9nOWCASLELe48X2otYh2CHeuz09mM2aaMLi
E3Z8x7EMD28qs3p0isBm4MMeRIsO+8/ugjb/9xj435edwJ0PQmRGRIF9homfKzbo
06Uva2Ro/gzRH+8xLtLW7OT9bjnX+Fclr4qjhDfL4idEX/Brs8sk6wjoknnXoBso
OrRle1M+z5amVCSQn4l/ExiodGVBr6J8oU4cReRqGOfEWqzNcdCCmlbVCmGdHAJH
T99aRbijfY8DWuepy2oW4qABzmEXtFfhl54tGz1XUTfcn51G24l7DfryMWTIbTvu
rP6IUe4nlxixp2Lymf+O+LCn3A9Yl2y12XO7joxnNdTF0Y3atpZMK+6TjyG9L19B
FnnOvJxiBonFXlmhPCJm5LMItzZSKc4Es2pw3w1ad0Ku9aueqXa1EPeLT9lXGezQ
H9HRJ6mcXv6nd5BDkfwBZSkXrArTr5VF9V/E+ybnI4cLffsF7XWBcBOEAIFwcdDl
gBOLloDI868YTKpqJScymOGCpIlmjVBJjj6Anzd0W1NuOqDdlJqU5StqOIZ0SSAh
7iXXFc56ztIvKHD8VsbGvVSzEyGY0eOr74dj0tK3zaVe9dAxvEZDpczM/6EZFyaB
ii5wjlrioZivg+HTOC6sYUChKM8jTaiWokAfkMyLNtyBRDF6BOiIzEXCRdNm7m5y
nHhXDzwp1Fq+jwl5PThbfG8qt7zBbmM/mydyNqGAK6Uumf8GL8C0avesMA0x97y7
g76ehj8O5KOmRn7/CM0mc6ZDU0uy9fWVdTEPNQE/F0eWjWCaxvwCx3F2pYChgzs7
PAnZB9lMYHhHC2WGsDpNy6CRGe1oHXEQy6ldoX/lBOW5GCA2DQbYgEmCYIqHF5yf
S0uA1GfHscN8V+LtacdLsBr3aqfrfSHCIUAvp9S5+BPUuMPxsq9fpxh+kp3LMW49
NTJoJFWdlFDGW2/QSbM742Tx6ROKAOxZtZI6UlkD5xwvDUHs+2rrGLAKKbvUR4/K
Ftso3FOB9Ytc+mHtsSwvBcdshK+0d6xN4mC1iYZrKt4zP7g8oeMzrprMi6tFmgPZ
0hq8YFeekvztd9s3gjDFTZeM0dFtrc5l2owK6hIDLQcvfCghbcBg/tp2vhU8eySO
j/+wL0G3OZGLIwpl2LBqyQ/8rsWXx+K1HJCPLcnEpHuxTTSzMJeqiBoiOY9wArPD
M6h32MnXp69glQ+r2RUTyu2gSv/hir7qzJVuLwUxnMrRe1W1/5sNyC2/A1YOmzfF
96ts0FApt1LIYSzIFaBzuJv7MwcDQmhQnF3QLeF9tA1G/iHL8uJGC9vX2I1VWpu5
V3DIH0dr3bLC2bA8DIKCJsTafHgCyUGBhkVJCnFHS86/oo8izUkilYgqz4vdU7IL
AMgA27lpeerZsbR6809dgJvlHb2kvHdEiKlMIqFf6xOcdq2+iehBPQGH5EIrXbl7
/mAAgxbb62+TICi5f6p13Szr1bb5OyhCCs4oYWN/BF1KRwq9QpPO1UnBr4UA60L2
bVht3biCHdIXoUq7z11zTaJ5ka8clQHZW6mnqk1hq/ePbhhlbRyQZ2aB6MHV9i9y
cjeY4mX4PCfe1iAFDc43edeOENm+CAsEKuOl52Q9KYxKoEPozQRWKcqJFrFHsvuv
IzrvAB+hMzUtMYM5N/w8iSlFBY9xbP3j1E3j3OzmNYgRzhtOw0Gs8MGjWwNTu0fk
ebk115DSSsyjYgmu8apAMUloejdT0j7lfhQ3ViWzxEMrv2fF6Q85SmOWku7fBk5H
+Vl8O2KWno92AeAGzbOi5d3xe+sRoMwQuxVCAUaEdxftbRv8BdUy8qrGYm7BvBoJ
wsKhiOmiXNRVTnVzz0lmsiD1mzEnxdukrYayASshc27Qje1Czc2ZLv5+UryQcIKC
Q/kvAqScUBDUsI+1iniqVqIYX170XomWVydwM2Q+av133/DPaxx7xgh3ivKDXMiW
uGCiPjo/QSS97x09TlZmoFMoP9ObyEvkeN7lupeunG2OPXPpgfbhCqabwJAkGO9v
YC9oE42deB3Y8gj+R9Mj9U8E4pm4j0nofpNooWzye2Mi55WEwwAMAEi/R3Uaiw0M
IF3neFQafsQgj3uL1Wo3ZCbzt4wmTN24Fwbu5lYr3i5Dd42Dx/56mN3U3djVbPQT
luyWzcPXb6NzfAShclODokMdIFB4zMgRWMLg1wdZp8HB3Llenf5zk+ZvAeyPvwMz
clRqWmvtIbfcq9oa4LK0gg5y00kHHg4PQ3ttKN+1nNHSXjJ0YXQKJkOIYikqWych
T1c3kbW6xwSr/Q693fuYD6nPPDoqIrMes98PCJveSC9AzYnMP6VxlRa+6Bnwq2Lf
/vNpOXXQENQ6Jzbn28XpRZBr1y1aVOcZ97mkkWTwPq8mJvv0vo7ggH6+M+FID2e/
XnxLOo7utHxAMTAT46pfm35YmniuQs3XHwIzYrqXrxccupVBspq7bA+QwGP64xcl
eKwpRXY2pQxY8xZmDghS7PPEShftTHhvRNpDLvaxLY0KIatHHVdqtBBXn15ZKrdx
fjU7sdd8HfIpA6ligwDIwy766sHMH4TXN4tX9Xva0PM88EomMCsJIPyQEWCkQpUv
kRxFKBz/pV2FMgIXa8NYmzP7Dl7FRhe468a9AbPK+iStSZyyjyW3jhpkn8BSA6s1
HWMlxVVkEeaUCFghSx8Hy3nTlz+aTuma7e2IObfJdL82VcmOgk/lCk2nMo5cqMyZ
VaZF+HEvXMQHpP2jB+GEp6c547zXFcQsT8Lcz8EBGr4tzAzrsf0S+IxB0jbg3nFI
7X5Sd8682HGwGVF3enWIst7MYIX4HjRjBMpQzb20di+8XEaQOEcl7ixlSrIts74w
iJGUl8/A4wI0bMrJ+fvG2h+27e18E9QI5cu2auzjPhyVcBdCA0Wwo8EIYltbYz33
vMDzH9mJ49wrTaIurLiMqpmf9P+ervA7vNcaGybp/WIAA5bfBOvv2Q3Nt37E1194
zUfpClt2D6rRBZhvaAP+dOZ1IvIs63fMcktBl/39OK16GXokz/edMnw6Bm7hBPMK
T3ylY8OCR0IoBYTr3ZK9y1Lh+kP8zgeM6tyD2+xAZUzqJsMnYLphbsRXUH907sam
7VG45IqI+aVw0vbmJDSmdJo8deIzges6CDxu5oKVR1WCsQM2VV1ia3SEHYfl52Eh
0mORdXKswP7Dsd+Tc+OrLDfQWSg7wPi9AfMoEpdZUIVZTGcxYCCyqBD6svMoqoHA
GpinvabqMPfNjVvQNwaUqBWJInQ9SezVwOPb+0Uy1ay/4x6HlnIJIK+IgEGBosCE
tAKCoPqfT4gmnrCi6VO8U7lkT86wvaHR1YRO6q65ahyFUbiOoyvGKuv1bVONnbdr
4y0D1gJi0R7cUihMivynUmd8bCBMRQuHgp8jnqyyExopxDUlNPfYCQAIU3Kz8vRc
opoNShdOEvxtYT/hxtug1DemicbTSmsHkkgihvDEHLES/8qFn3qPfYIrAsJvP4c+
jOeGHsZAHPoqt//Tx6LJd0mjkafkES8yQemhqCpLTO8ogjB5+b6HaADYbnagCibC
KqXRhWqSeGsfMS1d5UAQ6/4F1uCO5GPE32H4PypCmRCd4Ew0Ii/DJk5Ai8naQfjm
AwdZCqH09Dr6J9Sk2d1oygxg2e/f0894kAsR6FDzdN26eKmVGBOaPwTGUM8G3LY8
XfNA3s6Vrc4ZmYhe07w85R7dBQCMEOX/L5at5T0krZC6QWLM/buw9TI4fBdGsz9V
S1igPiBNaU5d3/S8ZUFaj19So+Pdpgyqm1qAIxl9q6mJrhmu0vmbUDTetyV1qhtG
2uNMgJGZAl9UY6ZhWhqBBiGXQVd2ovgoilwZ68msRf41FtGhJkYgneLLSzIWirsr
zQ93Cam+vLtiiHiOIiNzP61GwoX+jyR38XCJWz5T1lsETLZ5cI9M22YLXIyyHlCp
D+e6QezG7LsJiI7gl7cBMS+lUJWIrHfWamZVRO7lu+DXr0hYbC6MV38nKqqBGjZG
kHrp8xpzoSN0VY7eqmOc0/rJkjVfqvQZDN/K3ti6qodFcLX6JAvUAI07vHOrsvsd
SXlYuabWv7E9QD5mkrNKVG8Gc+I+vVavl32jFaEpZ43ZcpZ34OU7wQ7oeIidfYGS
SJM+ylEIL788Vn3L0DAsTQ/TEP0dtqB5UVeqoRUciSBBxh7x7Z0NLlGpoOdFtV4S
JlnyMRqo1NGbXimw1TBXX0qBHNcotzB8571mnA6cZbN1h2x9RDGAT7zR4VSN82od
BOdO+UvgPuvGnb26IdbweF4Pexnih01e3bdv0VM5Miv2d+95VWrumcop2Hj6lB8s
OYq97wLD/7xMCneAqcPQZOP5XLA4eDIqyrcpYoP1tI5MzeqFl8jhLaB1OH+s/3s2
R285wnnWW3qxoJuAMNdXugBOZAnpCXGgPUogUh6PVVDYUZqxRPsvEgW0kl2wy2HX
t/lak/17kjH+WB890rtm+KrwUXVGrMGUgfZ71o850JBn9neMMBuZznvTEP/8HgTZ
aATGKkVrvPUsPGZdDSJEYzSIeAk6Ojt7LFqq51UJu1Myt5GPlp25gjEszmcHsv5m
4heijUX1LBrVB6U2Mr2hXZdmwOuZc+pFj4ZR4sO9+oNQOgUdMb0TM5VSM/7JetVy
8iRbQaXQFwtxLs+KOI4o0y+tk30oO2e7LIaS5ggXF+G0U75MwY4awgZe9Biq8XCi
kWDDDKkpTLI46GTDYkZ1QbXOzXKpIzUHeKX+P1OxRyGEwv1q15f667l2TvZgOaBk
Uc/uPpHji8PFs8M4012++FrDjeboQpL1Gx5/Z5JEh3RUa4DmE3ElbvZIBBv4mIVF
lwZRZPnNMfLSzOhClJwAbZo8OJcZWsKlzcLQmWeY9PgkYYQQfFE8iUR1gLFqZxxG
0lVFOTMwfMBax/hM8DX/DmBC1NzgZtwwsna3vtkpsLVC0uAfYw6rldWCoUw8a0I1
/68wo3KLlhBhto7wYA6w2ojbz5ia6LKcl+3wd8lDcEJ1rHsHtJJgkXPT3Bb1f5GF
2jEERe4sQgrwITsp/bf3yArwnmYFxrBGbV3JiVId77J6CO/29H/eExDygXO9hldT
zpee7SAsWuBXLOQmObpGmrX9cQqTq98jV5RdBrnahdHBnKXr7C958g4eImqzk9lC
yO11pVwXcgKDFQU6lbyOmj9QgNBgaV9mgULbdOzF+Padf5YsbnWLeCoe70UmbsUy
/SFL2fSXqecRdgz45nRKRPDfQAzAnjRyifMqY6AaKLECwnhA95/ZUTEHjqiQXPvT
J6L8AnO5NIYkuq4xF7LJ2hoeysslwbbD7R8SxIWIEP6HyX8y9jnK3IhDePxSrKLk
zoR28UEKqji9W7hsSLPyJCE92p7HQ3g4KDL5GupHOWPtuBD0O4JTe+Tt4GOyaoel
q57s6HOf9cil7DXr0QN2SYjaKfEi6Oop1pyGGv19jh4/rb9IBWqMpMNJugCN3TTZ
9uxTR7sBdzOzP+cz/uSVIA/XR7WulFukOTg1LTZnyXWB4t+E7sQJpTpmsnzqd2xc
/11cATf+6YWMd//ns3E4Ae8PeUm7u9YCksuq/1t+w8swCWnszlFx1KPwFIZyPT7F
9PBjBLlGkiqLtx9Cz1xtwLiyAUudWJ7hbqHntSM7/57uQ1G1nT0/EHKNd6UK67vT
HVb+r0UGjaxsUlAFHbN+PycKVqFybTlAKRcSSWe1VGmLd29G5pVyPWS1riCHBTPO
yTxVU4/Ww0GW0mwitnucmaJ1DxtUqacFYE8pSp5XqNLGLXitQUlz3A6ylV3l5VPI
O+tVn5B5dKG/rq6d39oQ1l9IKKEDAUz9Y7Tib67TqKEbVdpvizcKVAP8jqoUT0N8
Cyklc104CCUMdOOpHDPDZI9B1c63uCvx8iAQqrnUhJlrGlRTg/pMNjMNydGoyhBM
uUEcb2Qv8rKyDCPZTwnVVPYVGl3BnVB93qwbH9P23WW8QpldSXQgbUCKb/eOJ19r
w/9VS8me2D2nPTsjm6Zm8+MTstV19+sS98i7Idka4190AIIFNt4wFaGoPVr7k6kF
q/THOAsYGwIWUfBZlhb+QXmzfCEZ42FKQUYUkbsEH8EgnmG6rnuI3H9oQsED1li/
IA7isU1Pb6EQrG82OLTjNtC0IbA9ccRnTOhXHXHogVLl0vFjL5nE9Q6HTbpYLhbC
aHSM+c8xkOB/ngMVsavkz/Nx+ygwW2PxM9xiEo53xde67enkti+cRWQDNzHVZeRZ
D18F+e91EmOoaf7D7nQWqQD3t+OspNSUrG3Nc5i8mYrCIcuATrqzFBcm8ekfZ7Ek
npbArRFue843Ryk/O4/EobRPULodSlLoMmHZHJUiZYMDELfFKH7T2BAe3x/SOSkE
ZnkrunYq87YFmtdDjzFtMAI2PSPXieldp2YJOg/q7czM5GdQrzY9oN51LV3khps7
xvvWIgHuBKQDueBIYX0Cvq5oFHaRzwj+ApAwApSJpvB031iDCTq7pOctpp8bl64A
paxKbAX1HB8aja3qldJPVVKcLNc6yTJsU05kBJFItvm/Vbkfd1tOTZGgMBQ/dlDs
c9v3c1e9DwqBxFJ4HTGxtSmTzW3oWqFE+FkN05+7F1h0S9szezDRAsjFWrZ+0Ftu
TR7wiSnQEH4jypcfkeLRdWdmgC4HOwcoBgYF858ZJWQblzq4cgnYfRWtngJvfrPK
hCm9tTTSaMZam94AarDjojp085hh5DtpbH1QvVV8cWRJQwx2OFG7Sg92eKEqBavL
wmmlkJs4hK7v220wH8E2/6Eh/eLvpGVgaNcmnav8cr3iBs1iKbTh+zhZRIWGOINr
NFCEJB7NG5/e1dMeaZLC/9zHS0xF7d70Pw9Y4ohsx3t+oJJ2MYxv6vwRrRbmhKuN
JyfRELtcbkU9rlU2JpZMu2gy0ic3xSWPUj6dJ7Kub+FyLwAsi4+ywznF5qGxPG8K
bPWHYjdJZRnKBE55MzEIyd0Ar3zqFM607cPSnWL0YC0AwJ3NKRH9IXDxSsc8q+ac
aJO7nfBKENlDZctKEI5+YnDNABLTCWJb4UkcRIhBsKj2Ac8uuN1rlLf1TYL3w2WH
TzjVx8DXCMsQ1Vsh9cCdL3gl7y0Am718tMO6l2o2RjKynMSY0fjuU2EnL/NkXNaw
/d7riQd1eOmAiB5rGAPY2/t7cOHES9XCDfPzZLwBzgBp6hfIdfuSh1jM57f4lUOx
KPR7oGRG4n2lxsa0nXWAKStupnn1L2LvWf9/qBdlRYm27zvVxmasqjr9M+YtcAs1
bFA4dgejmcC/1l7c9X7dilN9Sds1Oswj9uTkljnlrBYWEISdw0f4ZpmoIprS1U7K
2SfAXe04rxt1c9c+gKFlL3yIPt4pLckE8soQbX84THw1MnHsPmIc79Lrl/5YuwSl
ojgvDlCGCsW9hDac9kaR6b96OB5fmbFJNLyX99aeN1YRxh1dhrbmdmLUSfX5ARRg
OyxsXqWBGhu43T6cKTgCmkAcLNvQM86dHKuil5MuNyL1juqtK2o8fGgtcoPx03j4
hOROJjNEeXF/VO/S7HMb9VEBysMI0zmhr7z4fwnlsrElPic+F+I06ssBnJdfyFIz
HyQdexFoLFZkBtTvCA6gQonVxcU/4B8TfkIXzwnxbAE=
`protect END_PROTECTED
