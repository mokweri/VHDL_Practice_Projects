`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBjEiXv+LwIeh8Jh0mNxFzy8PE9UaVhkF2lYJIG6C5iVN3P+I50zcqdg5GC/D72O
aveE5NhT3noy8E71fMt6QuZedWwhw7FqQAhKGLEAgwQOvR/LnWEWlvx/N77V+fK5
rdT2kdr/GJkNErbxIEyMr9D1bHCCXKju9SnbL3ZCHE2aH/S9F6+GZvOPTee05q6a
xyT0lzi4TqsjPU6vLd3UIKppVozXiVhK9E4ACcXbGsyQKggDOB5PILqwKcWHEdmJ
IkLmUa6Y+MOjJ/ifNl3GZ67Ojpi3CDeEpQiNnAxoEudhEnw/nIhCi4dUMdz4Z7en
uY1o0DY6kZVpQf25wGnR2OWl1D93Zr8XnzvUZhDB/2bOwP/rQiLGqadcVDuAsw2B
gT2wKZFPQhuyaDaF2MGhleAXAQ5F73iOubkTsbLj01aP821lIf9VeKOw3IfbI6lj
huSL4vE7UfDCxxYg5yDt3GKgobwylRStWF8uSsX+ighDb8S+oFSbX/KFWmIQvOuP
Vsf57GnKX4UnA7ekyUFKKhtgtn9wrX+N+CNplSXnrthBQFuWT40uPLDs1kexiCam
3I5K4N88ZOrBIPlX4pj2vTDCDOZFUAVTWt1ffHeM37CpdCrrMLQ8rFHNw+V4UUvH
lBIy8Mtxndw2X+MQCUXU6UYTxE4hMfTe9FIGntIB73xTYXys9ITlI9I7skmPz9DZ
+LgF15Bg9K0vMKk5dg913KkwOBiOok3Eepw/VYIVC/i2LkpWp2XNfILg3oc++Zvo
dr4RaTzy9Epv/bNxoxpJ7/9LquWBiHZVu/xDENY2tfEOAcFUTMMRRwFLn4/I6q2n
qoYMulq/ZpBgqmS4PQsIuo5N3587iBoV509aZ6aN5Au706QtzzE0IYfFnema8qVb
KqxDD90wGw3jgQFQGRi3Rr8ksaN1d5iaUnzvd12JfKE=
`protect END_PROTECTED
