`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iz5Vf0pRJrKixWcdHJB/1J23pZwlHbdwmjoVsMgUwCwwBFs4HO/2/c5DHSU2k871
r1lmAHBZPIbebNBRDZg/lMdOGc2/GWzVWpdnQSqbFtcl/DL5eyS0RvNWFjLiiSvG
sptzMPt+WWeei3Fa4rePeFNpPCR/PmTHOwW5LVv/H9kxTt2b2NU35Z8VMK4k9U8Q
pPjzzYuP1ypwDqoNCikZeZClSKOXl8Z2lJGzAzSqUUMD5mSxUhNU7gOf7cqG74vn
sjlwnVCWStgp81Kl+aEb4k0gxnyz5tWZFmpTZAWcZ1MhY9NCTi2RC5L1QTDu1oPx
7LVqe6fVLCOyshs1Hv48e0FwcVtO6uKuOuiQFMKqAVkAY92F0dcURyNEm8luXskC
Rv7pkSiJ26Zodq6aHlE8nD/S19fkfsKZZYp2kOL8kQ6NiwJbluDsKfnpGCEbJ7w/
k/G9vb6nBoQ9pC9Cn5/UeXTXDfzoLsUD+/PlURADQ+9jGZgUpAtK90bzzHSZ2ech
wA1e+R9OTx3GZk4HC5M9F0iQqYnQiH0sTF0CixHEMUXODsmQCLEMpUqVUj01U17R
9fgArSTBrvKFEmeUTQJnuYjNqkpCuPzBKDkxEQqtXa6Smi0jS5mcDZwJmW6GCZ1m
OfSr719RJPMdxCJnECJCkcKSKSmumx9uBkZqR5K3Ow7zBfhiuEGe1w1a1qa6a13b
CgtVEgfRkGexiUvhk6so5Uu5hV65BjNvDVUb1vl+OM9miVELJIFqCLOXjktU+zwZ
uyc1HL9cVCoCz96NypTXek9P58cAfayze+eFF1D0UzOuvg5+dT6avn0FIdZd8C9H
/qmOp1GJmZ+khxfSd1IOfmM1USzWL/5rSe7UPPz86tNZQwUHtEt9YgZzJju0H6ja
yLMjK09KvroWNZGjShr7CyGmbN4M02Mpo1547UIeCD2ZPMX+NYk9mEJTOxJuQpKb
mbbUp0D/b/iF4EpQDQWe/O5pu1NLuGER865EyaqQ5+W3c0c94SM3EMAULZZli+m2
61SRauYyd2nffEZfZwWJ7VHrpxQrXeeCIJhesObHJ7IVC8tf6kH++lxBO+zSNH+j
QxTSTLf6xreSO9upO0DyZVg9h0y36cCRHGYGRunha3mvp0mGbPli+dY6GurTQaGm
AgahaFD8sC8PHuABmppaHP7Kzv3c+nviZ/4xHE2vP7KC1E8IiJvQsm/R2jBfq7LD
RQU5ZwvSjEy1Dn/frUPz7CkMno+ebaqO3ndQSpT6RMARxvTiLKo0RggNL9KLglyi
`protect END_PROTECTED
