`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOROp8xamUapusVXEqctt92WDUuyxTifCihmNjzqaA9mufl1Y/YFKwvT6EjzzNSm
Pc42cORj7PwfZwyRnBuYOhRr/deGaesN9w9l4cx8uFkYHmAECgMIfXWcbQlYYzhb
67rMhbppFYwR7/GgHdrrJnlicJG+Bb9DblVZO/ZORiVrEAbYexG/F4vqu3iiEqVg
`protect END_PROTECTED
