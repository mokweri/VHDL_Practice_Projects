`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTTXaqaGPoGF/XAAoEounjdFg7CGzgIJQPgqT9uB32yYg74Rqki5dJ8J6vlijqkM
NyaDnmIzIEy681D43VLjcc6YAt+Qpf2/W7mzJospddZ1ypq3kXYUxJGdV4czkrqe
O/r0daOqoo3IrQUrlf8Nfk5mdp6/jlaFzTaX7smWD84deXhu3WrIl3A8Z+037kt/
9DM2nWb8Ys3H5NA5Wa6CfOvT6fZMCDgDyQtSduCBlchVBX4wGVuJKdxZD+vOkjUJ
MmdEcaSAbIb7gEdQ7bx+DAfAKR3gY44h7JI6x+5amWvIkK3mOD6iK0BfGHaAHPAO
sbYb1UjM+gKBdfaRS/wTgne/dQUh9oHOk2Qw8HcNXIjj5FVo983cU6dn7GAR88CP
X/gOHZ/pUujhmU5LHBZlrDCPj91gn0z89s6sAwU3b0Py8U5rv4WhMQhseyjlO1zB
lYksB8lxSKeLiW+fDeiPm1SmPVPyRGuElO568yX19hw8bsRcc1d5v96zt/QwRB4s
jwSPC5Xngb1jCAZZGJLg/yYkYN2QLsFkmX8GJEgOV32gx6clZWnK+w9IkRNS30gh
bZy/n4iZlj6V8F/pWqcnt2j5dtaJJhOjQ/dVtPHW7liZKCkAcdB3xRlC8zKjv7Be
fz+FtIxmH5MASMR8evtnfmAyUSTGDe8stXMS+44vnd6bxwsHTXsbLObz5UP+fF+C
Y9TWO7+Q/ndE9en6HJeWIaKk0QwEhSR/iiWLmI87r1ndfkmU4C4YyxToGhS0QOD1
XZPM72e39FE6mMukiSHcUhyVbcC9/EQImIjgvYNHzIZ14lTAaYhqRu+5YL2LDVrQ
3pSUshBB6CqLQWn4jzIzZ1o7x7w4KvAQd1di/Pj8gkOOcCyCFj3KruEJ/4wE7moh
R/u74sZ9I1PXQK36i2zpJX/QEqd6ZieOgPYwgfSC+L0hQgYxbxrZRBhJv3OBk5uV
Brr96LyzQts5yvAbZ5UyJkT27677I5aUHGHDfWBTVggp7BrI4Cv7ZxObIzltMLOW
vQO/YAuVw5r5P1ObOV403stc7ACGhdLfM3ceskH1BS631rf8SwmeP9LRj7QqTMy7
6VS8c2yF4fUc26Ck0LBtuWxBvagaWXrN7uNPetBpwAl4O4IhgNo/pOmyjUyxSDHc
Tfv8+fL+VsE4vLxl7pUSAWAsWSlTPdaK4GXhMmJ15WJlGTj1uCNPlDJW/TNYafLN
Q8k0dJ9ODH1utJOVhPa+E8HZbqWcUWRRuhVFLoJIkEBykE7Tx84fXgTUJ+1Yyrt3
m8wQN2jan34Ag0+72kbuYcHnPJkHR8ZeXLdrRZUC99DV94YASdvqQyKVUSel+Up0
6yl6pX9pS2U1x6kg5+s1Q8lhaA9+tIybI0bPIrIXDQrga+Gi422L2kRAiq59PPOx
A6ecKl/LVeiA0KnALFigqYRUkjo97/RzxO6gX6dPfjFJitLalgUWM1yMk8JOrwpu
D9BPvb9y3tJl4D9doG7bCA==
`protect END_PROTECTED
