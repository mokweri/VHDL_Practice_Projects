`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ypP6duWxgpWbbEmXNoRqCjXXYXE4HMOlfiujFIOBpOUPiNhLKUEY75f5Cz1EmnP
uCAfXyith2ipuujqb1ZZfHjpc2jTKk+JtBb7tYzrAjaucSBzhVtseN7YlEZ0/K/7
cbbEoI8ll5MwCV+MvjqngB78j7B9QUKWevlbPOXumdXkRLMAVbtOuMFUlfpOXiqp
3FoLSA6c+L9ViFTJIDeLYmJHNPMSAdepiy4uMxs9R/Tj1QAzQnXcKboqWa1VOocD
jBzgtIS7LjiMEEw94ZQNJDETgTuSTf+MMyP1BKuJ+J7ErU8UFfzzMWGQFBCpe663
GGcRV4lKgctPJJYOOkbjK+hNGXHkEBAE2ibgqoGq8IzpXrz/ezgYMcJF/YdbTp9M
7Ags7caL2t9IL/BDgUdVe0l+zms2iZSZbNTO1Kj3ptZPwkXhyMB0m76oqPd/tsj8
RgqX8Vor8tBqd48K4XVS2DiC1w+VjYQkSD7qwMZb0Ig8cD/WbUPfU+m8JTxpd4gu
UDqfb4jgSvB8gMRcCAgroP2FUTvsawKefUg4z59fj00AEI5eIsZOd1lF7LUVPAa9
JTiquB/+jZghEWN7x1e6ekbfMIk/XSwp8OF7LXI1F+xAVEyexXwyxAuG+AbmYyKe
B1BZ3WXkUFBA+suOjeAGRWSUbw/XEyUUvJVZiqbqyw6tXYuGo9Q9ZMOLEQetMnUX
WY6s3KHe/ygDlGCDUvfkOaDXvgSG8WRD4oI2NteAyBhbATkfM036ykv3MKLWQ8+r
ao/QRU8zA1671wxdnH+j/bORFgoI2qQXhu0m5AiawQGPiQLAZ7VSHcagAiDsoB7i
vlDGMPaE6gGw78Rg10NKihEoj3AxODFg9SNC3+uaG5W9Vi4Mm/aJ0+4vjeS0H+Uf
0htVQxS30pHFmLyiiGgyU5hf4htQOCASBqhBUAUlVb8jFq4SyDK/ALDJJtB29foC
cWbAW2sJtbhqh9Ux8S5wMxmEsHFPxWY9/NZFBysDBB1fgAiPNuUrjnSltddEWq4l
FjKWz1fnWfDR6BXmAPxvEKaXXBD28BUisqvoU3nLl47pYMQ6HqM5YxJuKtH1y1ti
ECD3oIKWaE0jupTJqyNoUi8gWUhmv5KYy5upYCSjXMyxEXbU7P67DDHiRxn2rHsm
cZwI8bzSuhrxoz/MPSLmUg==
`protect END_PROTECTED
