`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXPeNu+3sekT9N5gXHCINOfQgFFbggPnuSoTmWggMu8w1q/4rkGNamMrGF5o++7w
Y7BmOIItD0QJcyuDcqfDtR/baBFmfk2e42M9h4xburc3c5cxDbUm6IbPQVAlcAv/
jTrLB/Gx7Kt2M1dnj9vKZSq/D6X78okX2VBrUfvivALKI68WGUrHimaFuZW1Rl1z
qHX2qNw3T28dlILr+KMuiDkoFSBJhwVYTP7u2FDCe+NUw8VQJ1cIKK6lxP8CEjYb
ikU8gg9G5j6szsrQWTsJWkNcs5TZr1cvZL7ceHacjpIox0e6OVp0XB1xIQ4QeVzY
U2ymqRJby8uDHDZA9qR500mGlJzeWSqWkEjNFxehL91z1PCF6fn9ZuO3UsH+bZAJ
gxY1lmLHW59UDTvVusX9zROLjqvp4JUwnsHyHMWI/RfAT+FkuwaIVMT/5i5aEyLR
UCHXf45jAACTcN8M0vIVtsfNV46O2v1bjk5GALglWoOid44zp0OlsswIHjSPHECV
mmrDnERZKqw3M9Fy/e8hqqJnTQLtrLgTMTWkshalAEANdRmtewBac860jwCTA9iT
lhUHmzkLKke3wNZ3KX99szRy6m+qdSxe1S+j7YIYH9XQTlQRsfV7/0llhxDIaMjc
9+GpfMt0tJbnBgie3dAiJwC9GFNfrwFdSS5w1LJPIDALrNZwl2e02h+B6ftw783h
C6iiv9Xw+vWriq8bJWNSbm72VFdwY8uOfBvrwGu3zRQ=
`protect END_PROTECTED
