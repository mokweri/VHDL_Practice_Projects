`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frL74cpPZxHdzgR2yIOr/Kraiq5rjoyZ/0/qJbQW1+Or8hFIfr4RksUYNjFvFFKJ
TJn5mAlfwx4nU2vxlfB2MYKmbbuExEYsxqYltH5p0wkBqiYspqd5eGCe5lI8vqhX
lyZ0UbtqEB2v/+wQwiZZ+IcashjpW1nSUVDuYaG86jK1n/yGXnJs3SZ8m+QvZiJB
TezJxRhR5dwLXRl4n4qSiJlGcxbPlT6Rp+yHgSvIUerSAJqgNy53/vdY4TvWG11x
pmXCz6hHgvq3EkVO/4hyAyNoNskf7KQbx47BCH081O00w1YLEgpwH8BZvelOTExF
aWEz6TunCBxKZY4OHtLBmqlw9UsiqVRHsdI66DNtH+tn/3RaMBcGu6vejEI7uvrQ
EU8ib6lQSrixIa13huDAKNYZA+mgkvS+kKTfPXdf6P6DCDSJ/H3F3MiJLVFsiTSy
DNjmUE77+8sBxAuqOYE72VHrpdeEJJ5N6ZbBQUx6RcOU5QPFmYabtt8zHWZf0TII
DLoTXYC69mJ7jbRfhUF865HxC1Lf7WNoo3/2XZ9XOIyNCWd91Az8+ugb0QAeV5Kp
GDJ0pGrilUI9EnHcIgyDO7tFZEWWxU1wM5cbMUJMWlSBCKj8esXpQ/ysk44o0Glc
rL58DfaODT0pgU38qSnLNBJSemkCOKoya+6k93f5bE/ik56PHhlhYho2Xzezctb7
LJER59Y/MQ9QOKTxuIqepLULm/5NK33j+/y8+2WchbA1uZajO29HyoaNk63K0ZxP
p4Ur8SKNWE076Mf96yVDIxoW/UsZr+aQNj0oTB+R8J6xe1ttCCbyVsxJ2jf4cHU3
e67dRyB3i8Cf1/VHVp7ZWYZjCfUpI7NzEt9S+mLdGOJczTHs/PQUP36hDEX9uGQy
/yTSWOXhSJ+iQT4Dxn/n2mcHg5lrASn0+dH73aKvMplMcvHkVWPefxnZPbHR9+0l
oN+iaSQ3ybqBLTIk6SUZETy935EPiM2k/Q2Ie/HnRC8uuSljJ5n2+Lr7abVPgV9b
Li+ixNlb4so5ovb6KG5v8w==
`protect END_PROTECTED
