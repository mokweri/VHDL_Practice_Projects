`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cc1T8vw6JRBalNJD6TnqBlX8ITjyzY15rUhLado2uFjJthqEsMI0vHFrokVlpxHs
MN8GilizSdBzULpCqMrzBt+DEFNaCM6PCiCVsLRRuTLndFv+b0eILw1h+mFVCCXU
26Tz776OdThuojE9qrrktEMMbV1p1w5w95vnG7u2KaYNeet4uhCMf8ldRwP6mij3
avKxsl7j/+CQM4a/5xFHsxnfKIixzsALr3F5Dmvjc1FkoA2umP5xW+Q3TGgQxK9c
Dv3tGrPUjgPxtTR4I2m7x8vOXV0R1/qvk4uD+P4raFZvsdlnr19H9pquHG6uLL+/
H4q8Dx9GItL4uNuwztd6fbD4dacegQ2PgJM5JZ6XXFfgKIb+iPJ7lYCgURtlVXeq
hnEoeO7ciECFb7JETvQEb3j+k1VwCA2mRpUqcV3/ndDQzzSI5N3BypocUJPn6g1f
lbvk0aBJkBSHOvcOmnkJ5JRLR0tkjnEA/3svKUDBpoQrpRksHqgeX3FDu8ZRFdQa
kIaZ5ZhsUXFJi1LeLw7/2cONHK/wBB3kGMkzGA/MdDtFzZeXtIHUpAVrqln79uh1
BhWnNYyDja6snI1gFtHUZx7h5t1rHp44lUSuXRp58sgEkpDvMEbcocJj3jkq0EvP
mXE7wjUDARjktB0Z7VFgx9c9Bj0xpihmvBgglVW0gONzlzuVBQQporyrlVsf0Ieb
EJjxyPBqrQ6P82tfDpp4Hkge9bLK93R9GwYFDQqsZ6eTl4E4F4uC0gybLmQa1wPZ
9nVafXepu+xbysfp0MIgtshRFpxVHM5GQTnVYBM26rjeWWpljuq678+upAJyUaiv
5Y3MER/ophkr18jGZrSwgGD40z5k4/RYUxixezrM5Mqldqey1SU4kscX7qBjrVDE
ROADtpKbH/FQt6wf/YA4SSVOFMJxukAI9bVrZhCMDsxkea+Kc4IXs77f8P3hlplL
v1p6Zc4McsOr42Y91Nr8VCvVJmcPHeaejn7BN7zOMFBsx07wupl8IL5s3TG9mwYC
gTtrvBD/zC6l6S9e9+Q01ewXre9PnjRnVypYrOIrolCg8BY6hTMGoHzoy4AfQR6O
Xy+vAGexmr8shkEzVOxSAXce2iUQ2m2GF4yLBEDsrBHgUXHpb2AsaueBNvO0e9FW
IMuWIYRCzAltb4n1SG8iRbAukOZGuRKU4PmXz2f7ZqOWQWsR7cqXyL1DWxqVQRtl
jS9njQGClKXgLNjqDuaDbgIX/cf1M0dEOC5WzHA2ZeoWSAq4hWhp23Rf6917WJv0
Nl2/4raZXHHmtHvKSd1q3pEvSqowm5lu8slvOvXqU33Be5kgZwx2EAK4WGAPiuxd
WCJkuiwqmoVn+LooDXrB0zWdtrW4dGo27UgamauXi31p80wiCnetrByd5UMr6WyM
kXXV/D/eRoenrP9DFpBaXGWdgDG9TvLOZxOh3ESMkuDzbUxOTw1if1hJlezb0oNz
P0FcOl+6y6xI0Mlb6+NmeOHsuNtbU9bITW6GdG8EuFlCIqlSw4i7/80gojPdKq04
UiDnfhPP4zPEypQTbs8d93bXAGsXbN9X5FM+XtJh5ceA93rCRXiCEPShC8KbIk9F
ODCdeI4fDoCes5xiiNWLjdQf31uUASiqsbyAL7/NPmk=
`protect END_PROTECTED
