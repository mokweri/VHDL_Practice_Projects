`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q2e5bvzh/tVl3vl/OZ+YGiaN625HEIDV4Y/3yacVTSfSPa12FKv3PBayZ5Ra9zvW
r5Gg8RGSx5uMnxxfCYh+GhCZElPG9Q3zFzFsIFw9t+8hRxySsJTAL3hVaVTdRenX
ZKw0nBcRdQsgORdYIgVko6MC6EbC4eCV8MChF4CoGEP49ouMXt+T5aJkEkpCQjN+
`protect END_PROTECTED
