`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmCESPrch0WBrqf57IImEP+etLQknUp4tCTNGPu+Iz/m+0y57D2JhNAezhG3Hudk
CR6749spEGZWc5y+/W6iswWfu3I0yahj70bSjzLcajLxLgMohX4kGqOvvYYllz1P
JJEtOmZeSS1MJmOkCwcsm6vGTPeQBqCFOC7Jpt0AI3UGNHORbdIwU05WZdiUJvKs
lPwLqUcda2y86vqceC+N0NfeyCY+/H2xj7EMbM+JilDJ3lDLP5EVwipzcq+auNpI
BJlhT1CbousxSWMiaT6UH3b1O9vNTG9iHb8saD+wl3SM/KJdeDarh1nd90xPrwGg
EH98l1PPH9Lp6nqQBmnoOxSU2VloJPl2h5mhTW3KELVS0V1h93AqBxl6TMkbnc5s
RDhlyfnynJK7xt2GLdiedd+5QMA7J4AYCcqGwNKPs1P52wu3TKCBHlsyLaCp45sf
65zjA7mXCmiqGhYQLhmJEK/vKQ0A7NPvPpbjWfqaFa3LIMklELtGbiklGWUCkrRh
vMjyzfC+TpOFIAz65eKOXOXaBCcFOZbWMS9jcWAsXvVlaqoVK9blb8ixFjaDZVR4
DBgsgUWqao5YmHRewxd+PsyJBpUyAIy1kwvPJ3egns1ou2QCjLvyInp94Gh+W9XI
nYouBa/KYkLTbRqNjx8shNDbLxuo2X5hX4zsnpnLncXgP9/gRv967nRlNc1+HGRb
c9OnteklCPPQ4ie50vHyeHtoAVLUAmZ2ifYpjyMepD337Vnq11ws3WKkKFHTBuaX
8mGpWKwaeHB2i5gToqaQUUc/vhdMME4rNzzIR4C0zBRjpo0JffRTXlohagR6wvZZ
XzrSeAvo7VZqB1/FdcgVNGvyybpIxjI1tTxAd6o/Xq2kCJ9bXXy16pKYHyy/Ce1H
qmNMneCyH3TARNOKAJ5yKNhRBkxAezupEZ6rzZ9dN//5js81ZRqEh70A79JSSfst
cysGxqfOZUstlhsuM8vyBSadHNDrrVx0h/pEX8Ht+TJmeGVsxVp/0GMvRpD02IMR
eK5/uqrROkzYjearp1H4WJpB3VQksA9SS1Q1Wo65zL+rWUwiSLS43oMKNaCDFSLE
lWZTKr40mF5Qhv5AykV4Xi36W/Rkc3fXHQiUKrKtVixlA816eZFksQx2gr3AmeTW
DNbE1C2QK9Zbfmm8xybd/JvH+GMgDghBEbaoSwxREzoohhaccgfaJ3ncu8DTqJJ9
fSj03uubK6eEV+bJ4/C6LP00J9EETB4Fi3ow4LS28gwz/NR7j3dtmVkff+K5j4Z8
RvbwzRw1HhugmpMfUe3mpl+aZ74/s7kqOj0Uifuhd9mGMxkmZLrw2qyGf3Mq1qQx
7L/J7mQogc/gMQZa9I4em4c2H4fUZkIgMtzTzm/HDipdcoM+YpGDUrJ+Sxs9vpYm
2GR1h97Dwsjg5GAzHfbmaEA2b2PffuehL3uBa4eVfj1QwkGcm3eCADKD9BHmTDso
r0cKW8o+EV7lm3CfNg+aRg+oBJrgaNLcLYXpoqZ4mUdIxIPcq3pknWf7Ukl/pQKZ
zhLEZbmL3gUZyYHhSD3N3P+GR1Lqp+1YfqR87ig0mH2rb7hJaXfiJ6E2hzmgBWrv
hTvSreSyA3Jvl+ojXvhJjRd3vfyQHQAbM5SNs3aMsM2GiGf4EhWhrK8RwO2dAZ7u
s4pD+1yyouZKMR/gDrdsdhoAl9hP+bcITNQBhiEXwUbgCrG72Z+lRBUeEGaMYLpk
BMDwTk2UToyg8g1jXjt8ngiJ205tqYsV93SPD9P+H1mq43lEFEjb2wxhjUKWDZHa
7Bte0ljjunAenACXyJq3VZ/6+QLa6fFWXfW2ExwObCqAaXX+CE7B0r8+zN6VCK7/
ouA9WeAllKyqj1VBet3nRyrzvx+Ba+rr1q8E/yoj0TrlzvUJ3asd4o0bm4g7yOJz
vojq/ScWwj1oEPNC1QGtXdc/MY39PGMRn7hL1Cc5YD96Hx0rJhA5vTVDXOm2dEAD
uxe15Qn0iG9ot0sV+B8uZ9I0eu42qv3wDSe+vR0DiajiSYlA2bSJoVPtHsOQHluP
SGHILGfeVdTFuE9gn2K29z1flEvnGyg+p5f6v5jzxZXkPaihkFQxYCOmQTyEIgqY
1u9KQNizq5a489qP1ShjFQWByzCJcrktdt938b+I9SyZWI+nuxVersVZRNaVft79
ydSPMz45TADckjBI75jIMSqeBFsifmyiH+soIjHZnUlZqr/AJAZ0iZNxiXg8ktNS
Txk+kxwajAzqte+6fhB3kmoF1bbwJ2oXB71qfNXBhGNkZ1bvdoswOVdFUvoB+wrG
F7d7wE0+tABOerhkH6J+ffMqNv5jonTVzoNYUkk6w6tvMCGD0aEQOD1KTTUSboTI
jmvs2aL5Zu/0E44r9xHJ93ydbOoDP3RabtybDk3Zwv9Cq/FkWHwIipMa8E5F9fBw
BvGmRW7rvZEmfIxaQc7aJpwqY3ZTpBh8KlYXUnfwjqzvE3CtiLAW774YiBOjGbDR
THrmM328x1G/o08TY56IT2n/+iO1kJJVavhAFLmu4C39WfjKRHjnoA1XILmviObS
LsWkhzyTexxBY5+IXRY0diy6aFoC5SmsXC0LAHra/Tz2+iSoDqLKrISx/bCgNLRn
7RFLWyBGSKxhZys1SFOa2rIR+DDRAcwP8DCVVXQXpS8ETgcXMUm9KKyEnKHR3ApJ
w5sthEzhCF3XnjQnjRpa5jLwQdY02iscdaHxRn1hw4TbxGwFiHbCLfuiWgniU0KP
tatnzhR9heLX7z4LMc85sO6pgSEp1dCYgjCM9Uz4iVFc3smzjLzyQxmUdt8NVU8W
5W+abGEQfSK8ylx+ulAIiK9cOW8O1fRcdgCzlkqOj6hWv1O+J/u/CpEgAL+FbC5W
Wvrcme0g1PJcno4cRXc/t4HcGFbk9MC9FCcfSQMuEGnCWDlhPAo5MnyGPsvWk2dR
lfpvELywtaRkYTZgwlzwCMOS23gaIhoWDiqgSWMnpV18jBsqm/La/9mUvDauzhTJ
iAfzXSfVGCoF0yFe6e08196iSqpEuM8zRSvX4Iox1juPfgyX3hUQ2v8zZ9BMXdrL
UVRN66sYbIqMUy+v6bYs3HCxu5zJ3n8f9Lj3n0yrDQKNmuIHvJMYCz6qTA+cQBSn
k8bPDTFz2MtTAsWDcWmHgV8K0xRaqRKgDryPw1b6qkKWr3X27RMYv7hgUAPEKTzF
49F89FUL1LJMbPj2BQavyr7BzW2DeOw6KKvCMxyMUnOYkNKZcWw2lbc8sqc3DofX
QNFGoDV66KLGQOY5xVPdKx+3x8JghzwmDaV+URi3XrMsYJjBPhg2aj0khN8bACnf
hU9rC2JbFtb3Q2pYK5vSz0gBDOi71qOpE0f6CMH21tcuKZ5TPbACq9Nh+q76KahC
F2KkuJ1+m2Q3VrNKZJF6rG39S2uJvES8gxtvYu9IdG4wIHF3ZTIx9QcoRNhpS6jX
VdrETAaam8+t46CkLJQ2VtHeKCzPs5LmGYsQx1WiXTZ07FilByp6uAYah2R+0RgT
8HjMDMp361I3rpT8XfyBpkzX3Nq5jsJj0m6fm7FduxqnrsiJNFYHe8MhehSANTuM
Cyt1XArKKT+75QGsKYLLywJJ781bGxFla4bTgYsML29PWvjwetO6HPaKVcoheqDQ
9Ip8Er/FQ4rTQr6k81E7se0oENYBYtJqaRgKyITESnucSAI9tAvrmqY0T8H1pQOE
2Y0/AMonNgeemTh3rjKJQUv6kwsaMFjUBkOuad7G5A7h4xa98EHk+AJEvehsD5yL
jzaeGn+CM43Gas07+97mYj3ALWIniudbgOR3CTvTWCbHAN0QNvNvHfRc2TeHv4ej
oZXdEMPrTakLfscDcaTvwaX6QPh/fNXHQGATvZBORsc=
`protect END_PROTECTED
