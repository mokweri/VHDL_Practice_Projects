`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ISCd3toGWvVKtNTZdqYOiVtmJKobZMQOZrc1vZB7/2NPji1JMrOHFs9BT+61ij6
Yo28LiRymrpV3Fp3MrXq7+cl+8waWwBNRA5s7BBmxYNs7Xozsg9m36plUXtWVUrG
nt763HAd9YLlyZ6JGXy4fPrOI9bELCrrRKzlsj00Wv4tqkY+EQm1iJVYfAzFCjAg
Q0HVhH8ltxPOKXyPQ7RF3kEW/uL1NvRkSbaGAo9xHo1z65ui/x5lRTb8dhGopz8d
eSu0MfxYSUmPoaFjsDyoFG075aswZSm1NAoNFa/E7qxqQjuj8oUmECEPOAn1bb1e
hWT3224urjyG9+wzsq7XxU6MxGtZMsg8fSWDiutm4nJJZ6psT+Rregh4AyH999ie
xQ8n4YRgekoShE0BEVZdsmZgUgkT1dHc4jKZHcXSKqcrsZu8Sq+PzO4tOA96MP5y
m+WumsLqesbAtoYqmnUr1PB8zEgOCn+vLbjG60iFZthhtcqzhfL1TCSwdQHqvcvY
zSr0gbclXlXI5pt2/yP/MPLfmLhA/Gy8jJGiODNXN1oG9uA/EZnw5qX5EuQ/7Sjd
jAe6s0pq24S8Ek8nSr3VcbNfZtyNOAdzjCfGM4oqimmp3IEjG0YnOFDlvQ1XhRfU
RsaUlsKfabKX0aRXvNhbYpr6bIVV/+lXX5VkufEVgPxoR7nzb5RpGn2o51SMxSDp
OvBzXeNsB+UTZ41uGybaKWFsZfU3XQk3iUl83IRiBQXF2pOcRCam16vCRiAB66gz
sxyDDamiKu0LSi5+pbYkF+UFlI4fGqjfftv0ZbzYe5lReS5bJickQUjYGPqDVGLT
loYaUhkcRVTlUn5+sp5ugwPlzCZKhz0K19EYuL+zOc8DlamQx4XQTPjwxy8DQ0Oo
6TSYn0Vl6mfqVFnPUeN5j1CWW5Sabdm/yzmwcFHi/vIlFv8oLhAaidB5w4/gQgpR
ruxYPVBLNfwGd5Qv2KCKH/gZslY/z+EcjUGKQ/Ra7z0qUdqSsFlzg87t+cmQ3bzY
AnV7W7i+dlNlthQ8Tcb1P5h0kNs3hzwAp/XY7XDtqfRvLXGv2KcJzib7/cpowSEx
Mxy/EJZJBbv3lvOzb8yckWKAnD/KYPar5szib2OH9YD1utnMORNM0JGAid0PPTUN
YElA7NdCpLHZ6d5PqsqSjBruqJCLlwqS+X1VjtG7GyV1BPSlSgrDHUb8QVhO3LZ9
HQoK/dxLzeHa7splRCzFd96a9gePd72a4osgTW9cwbo=
`protect END_PROTECTED
