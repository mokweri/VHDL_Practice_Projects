`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVwnf58YJUfulEf8p5T9hHuJKqHmjvOTJli7fkd3o2iVqHgA7/uq/AAP7yXPTi5k
jSIjit+tGqHFPCgNBXX0GXbc80OJKIrNXmu9GEqCWIGteP2OfY80jAux/vqvxpQ8
9TZsU/bdjgRQpfCyS7pdZk7FcrWnyzfGKyUKrcIXL0VLudoXF1jlYF9ZX9sfvFks
ggK1D1QUvvb5203D4e5HAUu7vBjx3GVF4hvvIE7JrDdYlxUEtYi9k8kLVtfrBxfW
8uYfuUGd3/staN+nrBvv0K9yI0opUSqVEKliUnlT3J28AxbTiO1MHOVIKCsa4LGL
0kyYtXrnbdm5nmsfNhHh3qkDeST5OT7O+lnz6AZTJqEyGEhekIl5giJ+QfDdX8Bz
Ir3XcouNkw4/XG8zR6+zYv2rvfv3ia2HIbRixVz3cFQNFIFxDGdvdrR2GidypiUC
ibEsVyF+a7w+PJzwLR0CBw==
`protect END_PROTECTED
