`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
49inFmmZCtXelE28oIH6MJbaHHQXG9QNDagYeKmGGmMmNU0W8jYm8crkCe+hPsRO
NkUz7pYfjT68hBdf21xYGTvueQ3gDSt9g3XC1pNcvthUTmcdULKi5HA0OKHGj5wB
YcVqvblpygUEG/1uU9bKxhjS6xBlwgIC4LnbsRh1NtbS8J5Aft/uSyyhdVzh9hCg
otUZKaImEYCKXoRtff/cpLoENAdczHCfuC8aCG4DS6ZEfhSu6O1Hd1hc2Ge9obZ2
cC+BpYRNIy3lYCE/oGXeXbkpx0Y/QER/gvYfhWNqG/PamHhI5g2dT2qPLaAauDQj
LrkQRXadht7N+MQHglm5wL0BYxkie+zGuAfMUICnlhepVm1ZxabBjMhSzEqum+o0
NkWseM6RWYCgXutEUu0yQZpQnSVMqR+fakgpYR8CRL6DB+iJzlbFFgUDjHoaSeR1
7rfq8QsXyvIVeyTM4dlWACgIl2K4bSXGtCvzVRKO1Be5RZGDLL66EyL8zbXDZTJA
/jQMQkAtxZNAEKepVs/CLkj1K9m8oqrXI+WUFrLRxjQBWKrgRVwrXYbn8Vp+H4oe
oPaKjjS5PAcDOIwEzHyEk95YhnH0ACOV/yrTXeQjpFmdZ5VLvGbyL+s/Xf8uF1ja
suxIofmISpHFFPFbVU/RZvDEnrDO03SyeMmR2FSMAmXz/ply/JIIq1xkxVPHQ0bu
N8Vba7l7vfHGJ9V75OWvapfcPHlE0mBdOGXIElmw9zqyZNJ3UQSKwr285wxhpkZm
PWQOwEkGzgiCoE4IkC2z48s/wn9myvKPO/JisTC7ocQdmphbyyHOe6jXWhGmJ3CI
LzGUDY4Ohc6DJR2wTiqT5A==
`protect END_PROTECTED
