`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5bwe8PG0V6OMG/VbRLxoi8CfPSkL1kppuew2dck7/dYOhBzIhuzmmxdhFZVuYUM
UABq4ljbiNtZ3vSHUUgna6MulYDE/Msxh1X7zoSw5kiz+iUgNRJU9auANSo3sZTe
LG1diroJKXRfvmHE73En0NTAS0x61MiL9uqThRT3ILmhnWIHTvGX13+KJNM744y2
0hvYwIGb3GK7djv0a2wYh0DEIgYqtsJqm1b+31jlWC9aKa1a3R0WfCF2TiK1nJ6f
4RQtOI9UxQzpD4yeA32S7Leiavw0UGDSkEiO/OuT9SnCbuj7g9e5nWpGRH6olMBL
tQWIYsPEBbmPF0bx4euUzu41MyTvgqsfYsji8NcjXyU1Er7jcBDZe677h9klNg1I
zNhPOMLKt9uDO8sCKGnuJEnPyz41aechPQG1mhswoasA4WX/+XM/gtcECv/dM8ev
CT/ZYOl/m7VSwchYoWu8LlyM1EphGSdOLvtrU0xxlrxGaSNpHIZk3Pd6K0e9wvBk
v0HsLDPe/LrOaJ5BNDp+gmi9W3CmQWyLi1YROOPL5KYyK2OyNoDr5tAXCTy4nVpI
z6EJ9+fPmXkWCwp7JybzPgcnt8ybWBsU31YK8ZJ/dr9QZ7rjuey2/DWjAHzu+QC/
VlvYmCdpgNLH7tvcV4fMmIQ1qCAOpJCkSjEp8FLWvENmkzotCpsI0+kH9jPXaKGZ
iejhJXlqV05Y2FC8D07Hra+srBeNSj4qF2nfvmGdfvTFykUBDcCKoCwpyXtCmjCI
lh+3zpGDsIQzbvMXP8UiUP9OAisDSgIA4yZKfD89N2EYRUJrzFwC7NVP8WeBzmv5
LgJSrazE7wFzfMBdf8zUrVLGYidtmgOibMXM2jQtqDxqBfzywS5c5NrV6OoN6kEq
HlEvIqTZ64joIXkUtfEg/5kDzFhtscCBX9RWGaxAFciqUCJSdfnRhctFsHo0ej7C
9LAd78DNsdNfnFXwi+SB7McEa+UEipqmMPDZfUB4BKAVVJdH+304G8Vn5ODbzz3m
8NzG/byqdQ7Mx+Ygk+8xNQzwbypgULcPdDZoRZ8hJ3TGbQ2PLBqzZq8kPxLX0ahs
fOUPrsf8bBy3Bh0xHUwzqfei5oMxRAhGO3XW2r41t5KEJkM58xB66cuiX9ZuRm3e
V5U0WjFEV7yIIT6EFJux//7+z16j+4zMPeqBW66snPr4jtUu61zkR7SGX8/BW7Tf
QKXTl6z6D1pxhZNn32c6hgYA3S3Jt5Z+QXl8K/snTtsX9U3dWJt12jkFjAosbgoA
t2/kDsXSxoGGWy4bID+yW8Jdze7b/JEyRsELcbarUVwfkIj1hoP3TTjDO4VmxK48
VxBTOhpvvuW+mUxtE/kXBgbaXnhBC7Mp7h+6iJl4kam1IWTas7abKz78EFPBs7x9
/Q5Nk02AuMvcsXZrXjChhhF6eI5P3qR0/vdFQkJMjKL3aWjf5fBae5AVk2czbBSa
stuYAfbo32LKW+9rZrytptwAAKaOvCzEsTIucZEPpyntIvlOg4qFbBg4b7wecv5u
AgeAtQoqeg1USWIxYUPZvXBwLdLrt2BZn69cO++CsWnVQGiqWTnMcaDnrGXHcWYI
MEgSiD3cja/iQHPzf87C/fdbElV7iJ/DjUDwC4b8HTBWnKefRAnkZUb1UHH46YP7
1jGpemrEXg6aYehQLHkLfu7KdhpGlRwtw646pcX4XzZWf84q/tF2I6wXv1UXejM/
Mb8lhtKrGBIZJOQOrpx+e10nkef8OhwxjaxtOiPntw0jcIHW3iRVQpwArazPTOGz
tnLciUVutDkCmY/acIhTeXxAgaRvK35IXbfr+Z1ltymRZl6hB7mHJHdS1kU5/XSc
p1amoqiVdcBYZXKlr1q2bo9LbMel8rU4bgVvspHWg0IiPaYxE/759X8TJRsZL9oH
v2Fpr+Br2seVI7ycYdlhznrH9pS8Gdo9iCQoWJM2NWCATPurXLR9caCvzsLxT88W
otYb1sjE7iZC9QXcMggiwUohX42SPWRg+sZd4II+nmoYt1fvcj1QBA67M/P7zjve
y6/uHB4XIueuXEro81yd/+UNOMpAIuK/YppyYlUlYeEdx+wcOlSVWptXfgXJOhbc
vsfd4S6nP4a6JilW6LU3f4RvIVzZEmVVJle0hQGOdV0Ye3yB+yWIGwmNG4Al//9H
93tZ04RRxa6CKTxqyPN91vz5WIb61dxw95hGsmMGRT7WvkpdUOLl9tewfI25H1na
9Tm29Na+FjMANo1kPYlr3zf8LgfUFwUEe4KBjnFyXcrv3Yt7gg06Ump2N4ojV73S
ixVrv5qqxGpANI+fuLFxd0iOxjzcZz94yTUUzTseKlx1zMrO9PuHbJLs3iBZn/Xx
pIrH5vIpRDKYEBS7tHZDzSwQ6qaFam4V6pQ0AF6eMqfxD4A2jYa692Tv8iDyPWgg
9pPhXdG9kolvmTTj6zqgtm4oGeyfWIdzjzu2H8Jp95xMGVBV/KxOvOmaUzhMUBEv
AeV2VXuIfVR104l2/YpdgHjjegN72/2rlKBZK2ZENYaFv3n8Nc1n84cxk0eZO8NN
HzN0Ccn607UMNanl/bBVnFyhfHvHPZA06tb/WlrpTrW+EdSy6nRXazzcYR3Z+n0l
uzsM89EvRCIC7tlyHylaKIjHSJTCykb6WaKXEbt/UkdG6drvxCntyRe/urBego7d
wqmpQRsottAOVIlRSxCyuk/24MR+j3J5iVrrjO8qUNwwVsT2MqK0cs0oFyL0nagK
WAfL5zAvXXssSZ1y/qEroJvGr8joBkfMTN7Zel7q97bVEHeWVCDJvfqP/LytE2q5
s+x3wGG/bRFfoXUy+GT1NaO+zLSHlcr4Kq05P7eQdhH2zbrpGz9n895MrqWQcS2i
Bftgqi6+wMuDWU1ep88JFXbpd7VN1x7mh/D1/MsqtZu1HiPzh0D4FQyqJmRWIrae
C2350Nkc5y/ECva+kPaxC2G+gFRQutrDUDsEI19FTfIH9cMs6FExFu+wWyrRlZzL
6XCOMl+D2jiJgKd1j4sYxR7wxQc69szGyyJDh0WH5z21iLkZpgSUWldug+WHr5Gg
pvbEshS8m4XxFPaKIdJgJ+pBqvQaY3d6DtS1+ASCGg1FVZD+EUBGMW5/q5cTmsib
wClkprt/ImNjSWm8tKo75kOT5FQdfwOvO5/UpL7nvhX+5jaCB1vY9ALl2hoIjNHo
U3/g09pDVLXrVGwkGw/upHVXtc9I3iamKRi1hKEYuxTowJSq0u04awOEgjF7U9/m
7HN4rW9Bvbjz3HGv4wg8zfwWWBIwu/iXv0xzAmMio4+WBeNscoLAPeeuZmtApbrM
GoHlkx1Uj6JGhUnqE20aOx5MXjNfCKJ1CbX8H139Vf4lxYUb9+SS9LzH/eajtR/f
Lr4wOw3r2Tqt8OiiHJ81DYvYw0F4u/a8f8go3+Q870YebnoreCVxXzD7i9XhI36A
GaXuXVn/qsvKmNc8RYRPStmzywoW5GDK4HrXzH47iGEuEfwAS1/SRLeV0sJHGAve
i4ejtNRBvSSR1QK/j6nC+vWYN3xJijw8krK24I7jD84IpA1mlfrf0hcvsNo4mqlj
Whxj3w5CZgH7Jo9bQa+0PesCkmD5m2eb/FuGgBcKkoG9WxDrTgy6zmVKUkcB5ClP
/+REyuWkbHniCMyWHII84+6UOBiaXUjDGvmHEvK9+iaGiFANXUD45UGMV+3dmSXN
QES8q38PjndyWRBAAS5hF8m8TZng9z3NoNeaZZ8j9F6jxwHtvwjxZlgnJ1UQlXW1
kemlGmb0GeiEGyWkaJmoYCHSwadXRMisZR45uv7QfN9DC3z2RKU6+9CnlFa6xwhq
RLiaXfGHWYF7v9nrH1TwjWprYU1pMj1tJjmXaMVUmbo=
`protect END_PROTECTED
