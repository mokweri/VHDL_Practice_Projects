`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fr6Knhw/7d2kxofpeQAtI1Y7D2EU9swFcEQ3dr7BfYPrUgDMe73U/MgLsYqvez6a
p6d2Dy7ce4P6tvSEQLrKut0krDDgcpUu94Q+bl83YZ+jYoGVm1TEDZXXWBVsEtyz
g5GsMrBkmQbRFUlM3ZpU2FRVuIHsFZADOO6ogqiUMGPa0miZ0qDlYpnWsLif1KAV
VdkQ3mwgWE7HeGC3KUANQf4lKylpJFumEXonuuZd47DOQL6UMwKlLhwnQB+2PzPC
Cn8C0b773ZigZpZif87+Wm2vW/BRyGXqqyCkodZrrtC0q47R6qPgRsiKEos2yzzL
YlGUdQxmuYq7X5MtD0RyoTwFmwbdTuuLJUfzbLYsK9+GKbXTAWEBhlGBoTkSpTeW
2+HphxaCw2vLqMHl6LBva3Zy4dfcPni5WRmv6RQXWFZrSk3hesWACprIcUzm3SYC
+2YBD0Msd+q37TXVro2ajPbjW0i2Ookp2GL/BpcQBNNibSRMozN5o9MLECZJj/Fo
sVKspthD6ff2IxSJc9Csp8bubg1d7hE0vhVvHlFExjO8myOiVNTvJ2wse0HKAaeU
emtTrrM9kEnqLZ/kuT/IZvw4RHNjbsrVlpczv8JjK2kvQEBQBZMU34OIYuZRmxwY
DnCmQA1zcWSlR91Z13167A5CYyaI1uHRWMazFe/Tvul6Tng2xEV7QTSyyvKwpaaj
Z0txK7AcHtYqRaIdfk+hyoOraFCn9lm3M9R25hq53Xpwun71tiR4GPTcJ/mFloPj
VpiwfCkiB08XBDAX3VDGYeJAxXNCIAC47k6ejZanX4iJxWltMsRntHVJaVTGgYZs
QL9PtUaT1EvWwgnhb6FSL3qhER/JJ205GpnZIYb0nc1HBxX40yybGtBsOMQxhF6N
azhzAMNGz2WYFAjvYDTREvl8cvecrC6lXyD5eptCMQmNISVW33CJ3fPmzTAS7CzV
EX4VSQPzwgnz8VhbkKYqKQThcr/glMUQWc1nWKmpVuPhjVCHqPWwiMFAeIOaxzao
h7jt7mYPEA1JWrLU7KonHZNphVZs1fhkFdYYzMadflNvK5R4uci+iRcWkjY0U+y8
CubOTmhcjwGN0sPLmoEW3zcESddWCWSmZEp+LEo2N8+aV81QhsczGkqhubzBiybS
h0jJT9LxfghprCVKJzzz/y/J4CcyKez1cL8TrlnbpcRI1S+9FelDH1Lu1snhHDKg
ntlLgz6eDmIVCEBvGoykz2sDLnHuEfKsYaKcv7emy93Z8MFbijkW50wbf1r/nzXC
MGBmWiQ7bUaWt4hmZjRADS6z6lHBpJ9DUEATSj4VvmDjEvAZwdIFCnkp/LKEleVV
YIUb7Q59lhKpbH0oCwBDf8gRF692yZGtJ4bsObCRrK3jA5p2K7VaFmA//ecrbMag
TsORI7t9ho4n7XPjIn50aQPWlnWeDSryFb2EKIRrQluSXKZCRzPYam6Xsl7JDTob
Km1YuiGyZNKWsfeGgHYBBHnYYwMncVmVLz5HXe+9iHPpqEhgRYJaamOAet2WWAvD
sXMOZuUYWaOWwnU9obHyxhhOtrt+Im5eAqM6F5beyCmOP9/E51ox2dIoZpWGQ/Pr
GuWhQ8ip5bLqM20s7STbkZM3S6769d1CYXrNMZNOHPPhaOVTk/gE6757dcnsBukK
ux+x2nevt/j4Tpb5A8LldN4A3LmakBNlH7eiss4rw5nCBwcKbTCX+jeDjtLyzO5i
gNSW9YW/GTJ5MLA1OHT+fMZ4PCKDkqDCC3WXWnGmA+rW3i00Awexe5OYijVRMFui
DSdvzqKB+TAdjAUjxbkiKT3+JSZd5pjxqWjADd70tLZ+q96qDxZRExvEtk/otRjD
FdbXBFG0FPwaqfooxfEcC7oRj8gfnp+g6QUV04dtLHRrfCwOWhh/A5gmcZrdD9u2
GfZtL0bwDnw7F+wG4pWtPGeuBvhE9yrYrI0+ixAsBrHQtRbNPRB6/aN649NcV/90
ET8UYBz2zQatX6FAThDFc2nHZKtd8M8l3TFIFcxauaSWtst+GQuvGozS/u8GV2dm
f0bylVNVa5cNSL2Pif8vSFWLE+qLbj7rWuwEy0YpDAqZIse1YKZWZ07WIap8bBJp
YDeBq/KTHTmgBy8s5EZGR+p+y/HzDcUJuzoPEXyu3/mnvZ0Rt78fW9nPROTQ+eR0
c6IrQt/B863Mc5+qhEdtN1jK+infyq5X3Lh/ta581WxHlD7BlDu9zsoZcoAtO5F1
V/kzwvs9nPUey0NS7jm+JkHhAb5eANHkLG1GTEx3N17ckhAakVmI9Hi1mOxTLWd1
rgaFUzY8vSI7f9Ynj3i0u4cSNXFCC0pBMSmCIwqFDdM83F3hAGVF1YjAV6Bt/L0B
ZH2VjCaxAy34Aw9vE1RqtSdvQMQZEd5NW/Md//FsdqJS1dOPm2U0pgp0wTYeR2Eq
SqyASFk1YInN9qP5mjzeE5aGQbKEt8xUYp/oA8fZkzdlZzKGsCquFzwFxk0aPTmb
c4nwuXhFKAqVBawS8irmUsB73CLmYb4amiOTCeSfoHdDUe2zNUue1RxyxZrx2eLV
Vgx0oqinqP7iMipHQbHAzfCbfKOqUIEhDzaYIffuz739q7hErFnH4y9Nkur/Ov6D
tRsLeig0XQP/is8DhJUsbdB8IWaKtNcVmuvWI8eVXsR8OU+SPHHSJU6wdmXCt9rc
JdJb0Ec5Mmc6tWI1YoDy9Kd/cV2mlcFZaSOQfPjGiwgBinKasIZVsw/oaZlj7yyO
5m3/TzAzNJTyACvk2xmPiI4oYVWO/4B7iMBa2uANx3DrVQm4mICQwpTJzYklHdza
h1NUGxXSUmcIFwG7WJmE8J8ITVLR+QdO6BSWgzhqKp2ASl/VjZEBPwmK/rPCe2BS
ycx8qb3W6C06I2QyqKIdnAw12zovEjM/6gxvDunO9dwFQ9kSVuEbWUERNRxatAO4
eTXPCi3o23ySYhQxy+jmbF4DfI+a4Yp8J3pl7yLSTEreRIGZ16TUp91VeZdecnWd
yP56l8acDoUP6yX9rX3A/qPl/B0zLwVuRIbRXCq3S1Td8mcOi6+1mI7bVOPt2r0p
Yb1u87G+85wfpUOmG7ohFTbYP6yPmy1H71dZTNdhuypWhabKAzPjI/IBpmr+Vokt
psrNUPuh5FH0MOvpycRK0OwYU6SBmc/dFQtJLIkHt3LDLy1HbRgtLuKMlDLDFoky
V6NeK4g2+Llvkb4PNhDvSLSkIWeIB2OuGZiWZSjQZ0n47QwLBdvcyF17q1wSVG0V
1HqaoC36TYJ+xvrrYiWo8Rac/+f4vhwPx/wRIwN9qt+z+J5EU+iwwqTAZPbOGFIi
mN7rm/3/wh14XOnq30N6VebKBjK/D35zFUIhpquCnxpWvOPpdIkNPb32djzpbwuh
bgHO31mL1hUiWChP7EtZgeazWj1+tVI8ZHB4Z/cyrLiBo4v6SxM9Wv8SvS2oK2OL
ak/StkhJSbO3HvcduUMwNtjYFQIJ4S8U0Y+iraor/2Tqtz4kJKG+3ofUhT+bn5Ft
+tk7Ne7q3p5hvfORVFWp6555UrOZsJKPGH2//i7Fn215K7pHS05tFWD5w7NRO26t
fO2VjZ293VdTWolGWtlof4/2bBMzRcIB0+gBIOhehQ0AvZtE01bDoUHa2MMc6XtI
/4m0zCtVkUGufhnwqeHYX7CpQqirGdOatwPVGUC6HVxL5DH2p47+LkqXvs193FKm
3P9hWFGMtZRT5lfrHVazQ9Xag6cCwS+hpt+939weortSDfj0G1CfH0q2EcWfbRdm
sRGnrCZAkWgxhdyziDxvKjh25/i8BBpnpiPJpRB+RmoN6L6Fi49FHDKMe8BzVBwH
9/O8hEWJ+LuoxOMz7CeKzIHGemdSaUkTvZIU0hWsisbms2x61pHRuqbT/gA7PosM
b8i8y5VVNayVEz6kGQlTs9AbopFj4qt7j9CVN5RToToBTGlUKfJ+jggyqQfhoWQX
rvNavM4AqEPgwYOU5Dm37yyEyQXvpBfvC5JB9ZLgahJk/g+bu7k2oNafkh2OPzXx
Es/v7Gswd9evJJ41UWYkTUARYixESTEfgq0MgFjp+ddlmEb1RtRKaaaEDR0/cBTy
yvTbIukAoVTdIwhIqQrTPQ5ecTHLO0oezD5DzBfX3ArfgI5zt1JvdjnUl3Z2q6MZ
HcfeK/aO2aWLW1vnfc4LA3e/U5Kb7n7KrOfLseCox20IMCdkfk2ojtYjo9aVBWGM
xKx9kZcfIs1tFML6u8ASCgwYt/9Y94Q5D6lg251o8cX6yyR//8W9QVUcxqrVVlBk
5Yw67LE8rM/wvzLUocq9Q3tvj5JPAX3DHWioj7/bD+p+vP6HS8wjrXCusb7jMeMM
UdfYIOzQGP9rHc3TbzJpwO7WJ76iGsZmTlnkd5gPDGuebr24dXrPJRM6PPDsNTr5
Satrji9TnvCIBcsJiS9Rdi1z2pukJHN1CXd3zY4g4i+nFIKCIB8b4QUpyRrfmGWd
JsrcVW6nW5zoO7beFb9a7yHvchOYH+wsowTw6RzTixB0qGlzTndcrMFy6tvxIuos
a/do4sGVWHeM1Ryfag3icgF4zmPkTR5DXKpnZQP32yCcpoVc5KgKYvrHE+wcyIPP
bjeb1i9d45s+1jBF7SbDKcjp/Pn0GPVd1vTyh0SlwdAfciBpCabCJW3vtL7q+ljE
o6MlKQMeoXmt1KDjkbDBPw+ybK2TYO3DKGdKfzMgjTYv5x6sSDcFLLyL7Dt4kxsh
PhMJzeHzFG0lrMamcmWoTXR0e+GkzWy9nRXxZwHLmgU9qEE308dIH4TiZq2CvOeu
1zIsqv5XqiA6KgG3klYnrrTivLFQXYkXhWuNtt1iISwy1lAZaLvboG7NG8ZyLOwC
S/C5xNtue6Zvhbx0dUJ0JNAX9BnCpOHjzeRkLd9+aTMA4Q5zy3aMN9RPN/ZoMfCc
MGA8tfDBpi1A77UShHeBXKdTYjDj/8p1rVxA8wGqpc5x7GHbpYw+mQcGdQLlQ75U
TYN58R8bUslWNINtsAKivdgSpb1vyCn674/GyBpfhYmAVE7EO/s/Tt1xwjVG6wkg
I4qon6BSLfEIJu0O9m+xWPPF+67H2RngSyptI/NcHbX+5k29cPE4YRdpydXMAcOp
3B1jqrE/4qSOxPJnH6vO0qyYwaBYkqyVGSMAicIe943OIF2RWocQy7Aw9FyK03qd
kz0BTfw6ptGRU9lM7Sr7zXmlgyoJJd1ROztNBjZXQDtjMJjY9y8Rwdtl9Xh2L6P4
RqibNNPQiknyZbXYBA4JA1g42aTnoecJkJVng3icbX1mbC88EysnO4hFVi1Xg3Ue
bgyozWUyEuwEI5ILCQX/fKWNMh2Tpsaijkx0D2blehzgUpoBG2ZI2TD4/L4soBge
Qx3ti2gRHasllCFPUoDY9asDLX0zaZjqBrMn3HZnzq6fOkcglxmS9EGwqBWwQ3Ns
MDrMWJmBRJCas8zLSIISZJpy8Cca1oPc73JX5ZX2iiwoy56BF8YZ3RKRnWHHbihP
o6gQ22V1Z2YvuRCE2rl/D6I1Frf6/bX9yrCWWnrj5XYGNsfMCWUFPjEP+Hjv9Fwf
rCSOZ6B54Xx7DMXF4wvtPGCeva4xCv5t/YrCflziivmS57Fkeh9lSFfTIZoiQ8bA
IZ/htkEBiWnVdNM2CND/9z4JHIrcXjIHm1RSyr7HguNWVo0aZwyc4DjzowrFuy17
OSftawFu9pQgBtvgsde9N4rk1ClYaEuIYlgaOx2lZK11PYmjav5ErdFPswcux2+y
8Hn//AzKjBE6mIR0gK9uR9Jtaj5CVvpaaXdDBBuVLys0E+57O/7a4giHzYx8ArSY
hlLLlIc2F7nY2ls8ZTVT5rvl13oR2rNPWMQYdepSmQg=
`protect END_PROTECTED
