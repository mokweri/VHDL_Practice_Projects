`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FreWuVqejeEX2Ki8Kj8YtZyiL8km6PQBmqG9xp4LohLqFwELUaVXQsZKYjy9Yb43
WXxKFYjCpYUEKhrxwlr674qL5NsPy/Ivxl1S8EYAJ1T9QWb71GP8tVBGnfo2SnJ3
kJKqqjdWmc385EvlYscb6OfCPDU3f8uVnmUTePriUxlym060Rz2HhixPfhDWOjzE
OmJS9wm9OVKYDydmlP1yfNUxzfbqfIX7W1u2l4F9HOBt23obFWC/XcggusD4HRax
m1hlBdvRqM3bwJeKB+4cPwmDL8MNd+cDFlKVMe6ZLr3HNruUMXAA6vgXcd36WpKA
c7hP597GJJkSx3niB8JE3oehGMzw91z4HHlrm3Ctgcj6SXkVPcIO40mQPQSYr19C
VmvcrHVL1P6cNzK3DUOTUjPs256VQDG5Rj6/vto98GswhCJAMXb6pJTU9zF3KXhd
ng3Uilcm0YUl2agkMMXVxzYdb6av2gHh5U1cHU7DTSuhxnRkj8OeG0UM4eAgTCmu
LQy8wd6cyALEpWRQQZlmG6P/uwh8Bj53xljXaJscGMNH9VNHNdHBoLjAqEceUI1C
QagHGrNYoZ/B5oyCuKDH2YeRfzFwoIjuwkGSKehjtCm5FidsYS9hrpjfg7TK8Sh6
8NSvMg/oZihMx8QYLSA7VRxpJdSV3BRo0Fef/iWvYAqHLP4rhcDNf5+ETfXh428z
PpCgfh1XBJfcVI7oc17K0gUNzhpCKa1ecTKFUmiL+dZsH5iZFunfd2kSYQfiS/iu
4AhsRCGGNyOBLlDhFlasVX3oQQADpsLL/5WbxuhsPDDXCA3a+xZT0PsGnhC2DcMY
yt2GhbxI0vAqPT5/AoJjnYUtEkZUufavJ+uw3IQMj6+yiDd0XklicgrjPx3soc/k
gqYV4f9zBqku1vCMgWRJivdyRWLBGYqLSxGLy/C8JPJBxfpCgEgUcGZx5WOXSAJB
DL7FwV9/jNumBIdj0WcqRFjDejkJ8oxWS0BJT8bo9e5Lwq/atApFc7SuxSVvx/TT
8b/LW59WGhjFE5yZBfuQVghySAn0pZpQaOIvr6BYbsY3BYaNZJsb3uwzsN3CfaMq
C8pib4/x/5QKNt/Cfcq1PG5R8Nk9DEb1YXMc/hfzrJpI/Cfv1AtYB3P3cgSBA6cG
lt7Y0IzTBb2KPdN+PTm2E7Ae9PaxtTGYsINj6tf/bhQe65T3oZIZT2QHNqI8O8ao
t34M9TR6Z/vio9dz5fa0j9M9Nqn8+KyFVERudIzsJMcC6AvQ5NN0HUFNKacVEPLl
6jJ+kAt/fn5WOL8orQzRTXTQYUlDHW9Gun09R6l7i+/BGLmz1kG+NcoAJmFLZz/I
MX7PkTR5QQuzXIk7IKGNkX4N7pzuHN2agwPLtb9wQuWlMejuGzgoPXzqQNGE8fTk
TlHd2eYLOpuSUdnzVxDydn7qv47JVvoeoPjJbmK+gwkCbs2Rb7f7QjN5gKhoT6xq
7902lMn7ZdXY6BxbeVW+1RO3TLtHJ3tlxJ6nRH6DyuAMV7W8LHdukHDDiPhSfXnP
ph0viSHhVa+256a3HFa3Moty7QiMA3w9g4RkSbF54A7frJ37BJpU3FqXMYlNZ96U
ioDknYqRLud1wKCAlUryeJeIL/Cu5h6w+ePmbw9d/c7s+wo+J5oGIaj4PSB8eitq
U1e90/v87K3keDO6ntZXoN5U7tKGkOwCZdLt72NcfoYaioBcxvfvmg4Pi/lDCJ0/
pQ7ade5wEzbV05aaPvxA3pXyCXTlSjoW5IjARYzp1X4FIyS5a6keraD4gStJ31cH
NgCLrtHXvgUpXPq++Di4h9iJ0rYHg+CfSMoOZUzlN807DfWZ1Erbpg/qiq+tKnk8
p5Cfp6EzUG3f2PRH62vSg8fZBfNv5+jS0wqQ8ForT/oHQBCYmRo9HiMc/0kmCHnj
btC6cQ1+EMNdVkIjQZ3etENoZCgYJ4gUuxK161S1vWck+11Ref/8jiPkJKbVVzdI
/kXJJKD5QR5B2PmKGQKuXIBwC+nR+8gK1peUMb/N5XWnJbjxqi6roZP92wasvp/x
FZ2xf6IIB1KxUFpdYzEEk0sDZv4ScJRHx9ySRns8bCDi4YZ3O0I3cNF2C5wNucsd
dp9aeZoh4kZqIUGTDrwZVCSLJthmJUQcA0U42VUIGH4K/mT8h/w5/qeQH+oOVDhn
Jp707MaNQB1IVRPGThAvZu+8GXTXl7opZ/1hv66tNZjqnoRfd/DhRmUn94EG2Fly
3YgWeoFvHl4dA+prFMkRL0t2/wtX3/3pXfNjK1hCRpLzbhihvt7PKalgk8vjo3Ug
BeuT4z/jQqlaLGyGAJV45nat1My0gU5yZ7CmbtX06HDCzFZ52FDIOiAj993qyOo/
vP+uJvAk6T1W27ztfga7ajwIVrzesC1cgcDvbosIDAdh9ToNlwt5Jqeed9Wr58t7
e+oIYxTAf44+/EAgkDRDNzDT4A0VOqWQy2fGYabgPr66mtUBn49MfMKzi9h5KAHT
yG1mmBMUae0aA5Ca/hjHYbWDP8+otFXO6Oc++2Y4BRoJufgHz2IvmaTVnnZ7eCp5
HOmsy35D6HQwmuN/d3UIENaIs521zdSC7ibPYbPGYlKpeout4sX601cWS1p9acxJ
jqxwofSCvjG5lWoWuFRHbBm97SJXcTqbKYec6dKmwELS7tm2g5mic0DAIAxXFERy
wPS6uGZlwhqoMwpf75WEGksyZ2lInBu4gHhR5lQpR4xa5cyMKRSf2WhHURVhLo97
s6DsziEcXqi36nsYz7+9nsEHCmREUJJNtfgxADqvEF8NQcfxJT1cJj8uHur5Lcki
ZH3CQ8d8hfyqud2s86Qkcc2wpxEHtaNoTwuZe15uo6BXT5llAu7zPIQbfOaZ3/cW
LKppVWrXljGojbGVOHAZuQm9luoOHyY2FTkfslf3VnqjYrljrYrUvNODOZ2WfbrR
11BHADtuEipoFcQ2zzVueSWcCWvftZAWVHAKBgJf+zhyvFBpwCCKaE5RI61uq7XF
xvDabPOFyNsdMDi9j25AdCijETKOstFnbT+ZfALdMCHl2GbxhkAYIhRzEvUyLI4+
gyTvs7ZLrd6m+G6R+S4pNqnpxyJi+i9xH3F86ZPoWfheK27/dmQWDZ79uiAuDfBp
TGU2F9SOVdq1jQcdXyldrplf2qSuxSgpy8I84EVsydS19JBbAq8Qrcst8S3HtiLb
07nenpZAwTvKOeHzQqGhDbDeJoB9SBDVElDxg3riICjHPw2A9Qfv++jSZv2Z/H4E
Lj9aEcCH+jNwvmQcqg+C8rsqU+fjolgQjSm0WMgT5Z8ZFB7AIees0s0YA6olAQjt
fYnPLUh9Je5ELEUErZEDXFMGzMHVoHQea4rQdliu3XgTUJ/SqmShC98VFcf3PeAG
jQZPNMUQIw1U8tf3xS17H4hHEswqpgw9vClx5E26PyzWVhpr/7NA9FwbNtUG9h1Y
0qzw7UsylayiEJxMw4HunE+njk66TYV8dmJIf2O2xT+FsL7YnfVe2fju014bpPMM
CJC3KmrkK7Ck+x69cHvC8VXr7d0+gXr0XR+qmWxIlCqoKVaiJ3mlXkq7N8gkl1jE
tHV3SaryAbYptJig1T8JRBjfIAvVpvW1UDxlOE5qcS15FiaquNAwTMJ/WU5nY6wX
DHJQO89KSwrgdL7XqRDkH0wJZS4CL09GFP6YybkzMuQ14xcw5WuODKRYSI+4kIHO
9HpbKKcunkV2J2iBPN8nAjERDwhEErcxM3YMprleKmpeYcTXA25RojMYXFWgW/vy
+yHiiaKTP/tiiOEcovapN/y6pSfaiS7KrnYwOnsdReW7KiVqV0Vw7DvAwfyK5zXe
pmOXMog7fD0Sg3tqhvwIGpJwiBwaBeGCqK8EQnmgqlW/tV23ewkRUXce21p0iYnG
avxBtDiiYCmP6mNhCBpBRU7qf1YxbF8E7MY3R9Tw6ZTi4pm9/GaMZEUenZcqdyme
j+0aOO5FddGSrX7UUcfPeFUpnrAEgfRFSXhLrIGEsScMQ/iheiM8DBOUmEqxhcbQ
urAbHVhwTEItfmzzZuzSxruWkzgVivNE9tTfird9ywg5pTgLh0SJjh+vsT/8UgrV
Qs7wgcmoSeVKXxKvsGVjr5YYsXaL0YXj41SBZMdOmRMwjhOQAQTw1iF6FvxDPbx5
RRbzZVgy7YciGs/etLGnbM+a5ygTEXIg8/5WtqSN6US2AFGzPZb9JNwNdgW+kcUO
mgvchvE/xNbvukQWeMchzo2Iqd3eMvH89AGAMKyOpck9cv5DA+MuWh5Rr3z2PHel
MgrwoUQQnklacb0FePxDrYiuWMZp8LKNMFovDccXow4PwPaZNngG3lwLRXQ1xZ2o
Av1fGK3pOmS/Wrre14J2E4AfY/4Rb4TdEeRDL6F15TCqD6b//XchH1S+CpgvN6LR
3hdGvgcvSvrPDqxCJ9UvO4WwbQtIUjWQrHyupF1Tyl64iDpyhY5zZxMVBpP9X8GF
60Akz/nKQZRecgh5zLklcXeJs5IFbd+O8jel9/vVJWPePkV5aK62zBC/vj4lKxpl
P/KicBaecZqNAcQB8nXT3Ko1Q7J8cVlVWvCQNLg1grIRoykY6bvgRO5kxtyqrvku
eg1JPkylVZCHPJcNctbCQxza2VVKb00tn16jEexhlbUDh4NfSvl6u+s9lJefqsvD
rAxQNzWUxa6hC3Y6fZyDQ/w9/u4d0xG3AoX7HmVSbffZuOd+oZcJUQe+7nQ/vVWv
2y8w51BRwsBjqLdTAQ/sUX/0NaCjxYXvGsEW8OZ+/PdnAap/fasIvrn+H0E0cnp7
DhfPAjwHDLfBVL5sU2sOT0wtbt85lrGgHyzwovI0HcXuX+1LynDGy5OiugAbH5aA
nWZX388pPUQscj8/JeZuT+QXfAtXnRSKAszug7zqxXIBBLHCrndJ6ngqLoSHpKrq
L6QPypJM1nGcmYr9q3HXg0vJK9rdigOwzzF1H8if0o2gN7Kmy12H7eFg5TCy5sm2
CcIotB0310w78OsnX5Ti8Mdc5+3kpcPApwfcbP2dow2hq/H26OUBoTct0Gx1qfrb
sY8a8SR8PogbVdi0RcJWwsPe4RPYuUeOibevYSNVdUYZOB4zAAxkpgjNE5dLLxBu
OLseTdKLk5pKTeCSk10hvjINjNHi8rWa8KD5aZMRXeuvQ6iNlYgD+Cb2NnqWHKAT
QDI32X5XC1AnUhlQu6+K5XEjxiS4WKXul326gB7LfCEfklwtbX6wDbqGBqI8deVv
KDzzEFuW4uXyMilaYVqF9A==
`protect END_PROTECTED
