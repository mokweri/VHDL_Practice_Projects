`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XSi/oQa879qbrUIkZiBH+2E/Xb7/C+phMiXd9psII65qwj+2R16xbESHCDa+gVb
gNa/k4LJPVM6YaRG55lei7EADRvXW+b0Lol080O7cMsILz2wpXdGEEVqrRMYjpmK
QjsZbyzIdeuvY047vIESCU1y7ow0E23XYUyVPVxFJxHDch1BWj83TFn4HivXuVCN
YsuzY20CmT3VULckz2EzvVWUEBidcsrsS5uZaumL1Dw2+3d6GwJLAdChat4i0f13
LucfUZ7cf7S4RY9BjKNZ80fqWJONS8FVF2CJe0y5lxwqC0eOi5hsDbZqktnF4S3g
tLA9gTvXX15CAeN3TrTprwaJDu8ThvdfHnwz9kZyyuSam5KK8fTD6Jsvj0wZMzto
cOuE5EEm976DAvIIdNZxgWdZJU2KkOir9+0wVMPb7Ti4TrOfw72TLtJSqIuYgpaq
3rIoLeE8b9oYEBEnD/x2QirhclQFakOuDpt587L6ZpAHiRJlfj7lj3hHc2xvIwcf
N99YkvF8N2vd2tVikRlv0f00IWs2f88fn8V1yL86+GkuQgFmE3ehf01wc0EmSlFn
draAeBrPYq2mTMMdrfTm5uyjYDehmECafZSJwmZ1AI3UFsbw52UI5mcMPhZcqc+K
AxN+IuXUfE7+puehBm+1XqllbBPNXyDUH68Fwv0Bd8scSQw6BcVgabJhJQDxi8re
FbGkl1wBX+rXq8u5KrwQG1gSkMx8eGUp1KnsC1CQ/C76GGbbGDvG7+WxOW+J5s5e
JHoumngl9lCDMrycauu+eEN7dY5cvlsrkK9zPowqEilL5YwMEGGe3WuQESY4C90s
Q8HQu2zCr92Uzd8SA/nQhs6NDQ37iIKP0tyu8sL+CYaPIgkv6kWhEoQ7UeZZ3eLH
u82huingtN1KuGkMyPDhjo0mMWY5HYFGF5dXDUsokR63w7hfuqi+ojqCGn8IU0p9
t3oDNpmHScWDDnmlTpCqjXi0LOFdtiLRMQddnnInwk0D7kNpQqxRTSVyjwAp/p+l
zXBtpdhT8/bNVxuFFdzHoBC2heZs/Ji+cqsf0fTtUHlwIs3EF4kQedpeix/DJmC2
d7NWMILmRK8k9Y+ktAppYAXS+JT0wO7biPvKfkboKkVTt7r2s2MSUVVdwg/9+ggN
s9R3EDrRxm5udGmgNmnoUHuKKDGbqKtLmyUF48kSJonU/wppSZ/AE50gEuq3xXM3
o/1VUxEFjm2r6/5QxTBOa7qCdKc/tYSFyIo3gmp8jVEZ4RK558X7bKJVAC4dF6Jt
sN+oLqi0p0Js1YYqyuALVNn1Zfekb9UWJTge44DqsK/uxtW8RD1OYY2z8VdwW1vE
4CAvJ8xFd0bCmMSz/5e6Ua/aDqrhNmba0z5rfVBPE6tmxqAYnCEskwCMJ/ldNrWF
4b9egBHF3NgVX89y/btT9OQjcgWb9A09vEg7MwrG7Et3cYo1TaJ93X7vjbTxoM3W
z0oKO7rk6y0ech+vKnAMpmb+v50nj+5hLKVcIH2iI36JIGEzityZxmU0j1OVs12y
zMsOr6Lgd/V/LHgo/Vy3fD/k3I0P64DF42IR0ZTwY9lYc9fDGXaztawB8KNsKNDu
p3uE5ckwrTUIivY4B5+HgHP8jkwohztuIdV/yISn7qczQcjDmf7b1yFkk1jDUW3D
4cx0GA6Hg+Sn5Q5GQ+Fpn5dmETqiWKcLGGsHoetQvSojo25QxDmk73KYT860g9bG
A2uCjr7rsUKsbgBGF88XowiiKxPJuNLdoC8Ytjx4eBpXW+5AvqQZgf49NpqNt0Uc
UbctpB1za1si3GGZ+Y/m46ZXr2zaYbZkTtA2ybRPe7AE4zFIxnYWtPpJlMQNd0xc
MkZjF055smgBoAz9QmG8AMlNEmR1QpIJvnVba4/0rddsOmBJwtgmCHielME3mDHz
xBuvGZ6gcf3Fm8xbc9HxVD+nwn+AXhaRZ+jYfN51N4YcqUFpB+XAzH3Xim9gvlCu
w/6b9YhqhW1CVuUGlAKR8tqyP504f2wGNPKvzkL0RA/9AOG0L2vVaeZr6EQUiO5+
GQClNLqxVuR3grOGMGdh6niINrtxvj3gOcHWDsUbH+sNEXrsy/CQlq0fYqIzvbaV
2D1afAgkYmD0nWmVfYveGfFBWD1jo3Yu7/snEGLBeoy4dRVLz7CszBe8PLGLtkDY
7lN0xqJpi5aiwVmFqxQFfhVqEQ2GihagPyH68GyWWxLOiyOzlnHb5y/EB2Qg3BbC
JHSKOo1pq5qNwiGJcFcE72XfOo7uZ/A6AiJnSKrh1TmY5Y/q9Vb2a04alpa+yp7W
H8MBUNl9xFyEeYSg22tIHO2wIhyLu5i0qPEoxXkej/XcYlwXgz+WPbEfuIpRa+gV
TvSDVGCqd/x/HaFCAfw7KJ4h5yp9Mt/Xui93YBi1GDeYSmBgk40Fi5fCll77fJIg
VwBZ1z0MpNvymQjQuToQujukI4pNPefyzw/KQNvgK0/fSImbAjLBGU2DGnbuSDN1
42xHWlJ1BWwL2qWepvQBt75vneN150bsNTOW/uHW4qXGMeZz3dm8MBnCIKf5hMth
OQHfIkTxff0/kyNX8oIwR4Kbwliyn0Y519gYHrluzD48mscKiH21W3JpCVYx6Eh4
oXKBike+MUFPvu2upa8h2r7p3xKRepuceUVoxADsCzkbm8HXrvrpsthp1S4hHFxC
DtwzGj/IpTAOPXAplGhO3iy0fEVdVByKmgWOYs+L0zPfHBhWZJ0DZ4h1V1+PdtkU
KhZmd/BUqnIK0B6nbhJEhX8BYaQJfgizXMSgpvIl4dyH8Mi7WB0mNcnMnruSCvYh
7Z6uaIBaWK52W9UVvqS8EX5gRqxygwqeM48/vT79NgbMHx56GtKcIpMPFK7w3ow4
qHTK3irkZmOfDgmpQcF/bJbe8MNzBjOUcU4d/aTtCl1NV9ldNEWdr6WtYFx6irnx
6kIpq0jD/uZgFbJtRNkImvOWU+rAlvg3REVphuJ83qud/0AGaQOoNmWNRHhrPS1C
gq+eVaJhckT/B1Xo6aM+l8LVXmGaU0+5uyI+T395vJ1zBBA5Emlj6IK3kFmlHn7s
GvTd2hePZAd0RxyFS+stiCMorRufI5c78Meh8Xm0wh3cl0/i7YWI0hEGszxmSd86
OxsbY8YR9mwBP9lxG2RT9wm9hjRuAt3oOdryrmwalcs+yj4iGWC/Jyt/pSmLlXyD
tgl3xqmcPDo2m7iuK4EXqpIMnb+aQ7UTKZp4qDxXE9Ca2eHFKEsK4WyWMHfuIl00
H1e44VvOwSMe9qAedQqsXozuk1O6qlVdDSpqFfU3tTaM7w9L0fny21/g3b2ahSzc
7/dKXGQUtIt1rqgNP5fSyOp8lxWq5NnFqC1CiHBzRS1JauKP/a2gg5k0W/N1q0+y
pBX5sCoP7OuiLx/E9ITHZGgtzr7kfIW+bN9Fvp9y0cO2o8Fwiv80Oa6ap3tS2Tj3
3aU4Txx99nQLEZSztzMp3wXIDZwVZwNts4nEs0OGzGLoVI7LvYLfPkwaufW8D/4T
EfaVokgG+YtvH/ExSwVdvDDdRqkbL54jVg1w/N5Yo/h0JbKHo9mQClm+7VxIpt/x
jF9rEIyUpQCxxqf8hB1DDFaV1+kObprqVZDY8w3JOmTIUgGP7NlZOSSLOuVoPeK2
esjgLEkjGOQaieX8dOHczU3qGn2JDrwuurWmpnSVIli8mR/o6/VdJBDHnvwY0hBl
/qpw+ME1XiTQL8ZEYZ6eLCVaFWYxNKR+P/kPrWY78ApvJ7P279xVdyxcBdRyKYZM
Lv4tz3a3SERyUeeYI2n72p8P7rh+4G414/kaWecqVXtSMcZ5wUV6rFmYzVU8Bag0
10U8lBPPFp9tWFsqyise0j95u8FhDR6u/NDprOfKHijqk9/rZ02KeO4MEsPLzJ12
avNbcWgA+pG/NLkrOI/fYEp7qAKJoVXaSR1uyZ4rC3tKnoinDeaMXy9eR1FbDGf2
nJyhjTMCyR7O35Bl6r9oTJsveEQEwggWj5oZDgPXLUI1Vs8ue4GYgEMfIObzdxNS
o1fSB0NS+SFaSCBIHKvjVSpeofDVMUxlp78G+/st8L9Ebljp/lC+Azn+roXcaPHc
OSG9t/4d2oB+kk2eM5hU3S4ZFV8gnGYMZGTJtTOFkXnDOs+Xqas4Kz48NvJ5sNQx
P+fInQ8mWiesjhuGBTh9wnYz6LwjKANfRS6Xa/vH+LzUWLVSPEo2AOeIqm7nKtWe
HDqvcA2S3SKHqP9Wg+vKDVpcvcb2f4hr9Nln/ZH5V0pfYjgxYgyFeKXPQxk0p/0K
lXeSjX+I2ZPa4cTrOltDBwn1zEffRONk7mEH5F5wP21GioxJWYvHMIkbIPXRhSWL
IO8KKq5siS31gs0VrPgH1WhhUu07vpepIp/w7knH8Oe1CnRja6F2jPCq8yWGRNFk
CXZJs0SEZerwxNfkg6UaKTHSy8fjnBuaXHDduu665kH3ye7hnd2gO+q+fiQK74ko
Vej/19wO1G8gNtvC4NsWSrKYUk0fZ212SxYaUiaivgOl+VTuxna0/FiQXRRYzWIA
tXLVDlq+ASKA1V4KFtMQI0BXIA5oORp1/sOJHmjDt+/AO2+NByccIw2XXqeyQ/VH
CVoV7qYRsEIoSETVwIiO/so9ndTpX07Lohv+0vfR6LbtcLs8HTt7ibbpauCqRYU7
4nCQmFL1P2Q50NRWcQzDclsAFWmeSq7hAXRPgrGhg9TjBDr4D5iVLte5dAxW9nLh
OLg6W2Q4JHpgvOrnWFckvFm7GX1SSwy0kj/9azuXAHRkfhLql+Xm9XIgrnHO4SgR
M08nqKqdacf/JrHY2O6SiSXmnOC+7EAtjcrmrSQ/IWRVGzrdZp3pvks/C9sTHnDm
jrJ8mYq3cHT1P9iJlTnpuM/dTTGivaffsEgYKTW8onxQe70G9RUzlgcvcUX7y3h3
kLmWQfTNCZCbmcq90Y9zvnxDt7nWAR354CZ0lgQ/2zgvsor8RzZ3MbsKERa0ZtLA
E+ZoK2JAJOrDL0Ghv3a6v86RoliDms90h0wD+Oz289S/l94AYLow2PpTUEAIS6sE
Op3yebeCVDeisgtkY+iiaMvrv7lZnl6/YeUj9b9vd6GYXx4FavApAZ2M8BlYUyH7
O8Xr0cQacNlQPZCxxRL6P2RjXLEYIq6F9pCw9XKff/Ii+bjglvNK5HAZTuwZjBBb
Zkg511Laru09gnXdBd3iSPq3PE/CKWhdyjmW99MltTrVlpGkyW2qWeBpuqI0htUw
MqOt2k1GV/ZOlDou/sEjNb4CdO5Tkc7tlbl47a0ZD8+h4TnewBzFcbuYNR5VVUiB
`protect END_PROTECTED
