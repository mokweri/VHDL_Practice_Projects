`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j22aTbGlFhm628Ryz3GU0qlb8sj/P1pBOZK/OBLagIh93uBe5teCxiV9ciRMRr3B
dDLZ9KfHuqrDyu9SxT2ZkD932h6GmqjfmyrE4Qg7LMuG9CxfZMX6AdlP0BZ/DRQy
hXvT8v/Zw81R0y4bp0a/fa15xIwChPitoQ9C7ncFhzNX4FfJu6t5eCydi1ubN+s+
YdeqjWCBB7iZxw8Gzw5Sc5Khou+XKSq9EUDJ8pIVNvihznLMyEX0YEwgax5Yd1b8
HnDGT3r4+HHZx+UJ+FXNQQUOAZkuyRmFYp0nbzkkVBbZKZIM3ZwnCjZAdpwpf1A8
eRfU0oxXOLoiuOZirPDPNACg1/AnM9JUBzEkmzoDkiqAqUKmjS6KkJgbUQ4GUG4D
eRGyHqwxmD+39up15oJai7wWZW2ryKb5G3ABETqqomOE0h/Vw2O3NytOK66nj+Ap
Pe5DfdUNDy2bbmgwVHVg2/ZOFTbcmgyrAw6EyXM7etlYePCoZyJc+xk+yHYg3Jwz
JHyDnykX5i7QDGUeiDy+ae4k3R/pQlXOitsQ5LUDgdo4trs7ausHo5scNYzKPpCz
QLpMg1ctFkK254N51oo4mvwNu+W2mpih3qKauGI5j/QGDs+3JR28AUAeXH1hkGmg
54W8L429uc+zC7ZePvxPYXLpgmUwMGik7B/VW87V0wg0sh6L+op4jjVFvhCF0nqj
el8e1wSsL9oNLE4OY8/HVB7RZ2fNjmKjbd38kw5foUeyY+hw1w68Xk/aDtnVbBzW
GPMUi4SnivJIl25H7EH7oDCL78FS1Uxbk/Zon5oc66OPf8+nMzFM5AqRNGlie8FA
ivZhjARd3bUfEm/taJoWLgcwvLVs/qmPQnu/XhGi3ynV4+1cpfpj5LmiI8xBV8pj
dEQjhM0Uk+eUdVRVuw/3HLPGl0MRTRT6T9qlHTD0RfJMz/VHR9qeE1bL0wy86jYv
Hp2ycO9nmaN1nZVOxpdWMMNiTsWelYtMFJRc3zooGgCpcMfeJGFO3Qlqp2o/kW2Q
aVwTNaC8DcfLCv5LnhEmcMIsyjA2gm9X7Ff+ueH0HIfDiosw6wUxs70ks3uAK4ns
3f49d8ljJIg9r+xU4BbSgVftSEbGuoKRK8lpMUzWEkH4dnICLOaE2FLpGGqBwOq8
sHAMEqRDMZJ88INIWfiyYJJg2RBcB5AsliZnE37xCLr7rb+BRVBvFS8j1I8KuCxi
OvS9I1t6sElxWygHYyxK+FGrkK0AkJ+WqOA3i7+DwSJ2a9bbfDYA16v5ForVG1jY
d715Qkmn0z7tvzeC6G6yCM+5FeVQ/h3hPzPlerMKxxHiF8H/dwm99XIkt22GPqRJ
SsAQKcdfRvr4Waf4ItvH6tWRXd/M2ng+464urwuLWge5h6X3PhyAAnT869flgKz5
6yQtYJ4tN5OwNcQyPX50CovYNCVBC3IBDLbQUvrPxWssau+wCRD5zwJUJZABzXFq
7geH73LnMo/VqeiO3Ftqcbuf+1kSeHCOZyTiRH6OoFDrTxDjNsrFCNdh2O+3G+px
UEXidhThY3+NxglOYQOYMzkZw5FUgKBmnBUjkOvKPPv8HnXt2S/35tlweR+7/zNA
GIvpWIExhXZjvNaDCRFEVNk9eH86A+VB7KaFzeUe8YoeLW+/jzXsJhr41fqeUqbJ
ck/Dox1Vu0aMejPqSU3EjDl5F4t27cgIZJV0pn0uGGAXo77R8nN+bBr49ATo+SrE
OeKIF4YVsX0nvP9EZw80XDFRMYNj9QN7/Sb7JJm/7mf0kslgzYc5pEJgU1s7to7z
Okqmr+VDCB0PTpaXR76KtRPkQOXQ035xnULWrEjh96CVMMBd+yh4Sn9aDROn+Gdn
wBckrbnSjDMrcc8Xuh3Wj49lskEjIR61+BIZunifqQREf6j2rpJSRuP6vkKZpbJN
qwwHCq9ap+oXuPPA6kue72Y/zg9QUGtEABjWylSQFWMgcj6ZiwBAgs11xQRmgt7H
L7h7+hzw3Oi0q4e0SWmkFsHlvtCiiWFW1BZooUCD4PgaXYLagreTTGui0QVXirUI
bVgiZlY9JJxguIGpPQCE38LRRgPXBsYengrpnMHTof86AB8Ow8hxt3PogSs74ahg
C3visRK5NPvJ28WrraQo2VwPCdXB8l3Tw61n5o8i9/xYCDe9PxfnKJ2LA/EtteIJ
Q+H4H98gblCp4QFy1CksF/rbccfp8JkpRKhHIY8WKm+CBfFASgjcdPt3tFuat0Qv
QPNgh9Ne3a9VOG8bes0tWDXAk16VcYTPCfCzB4E4mec3dvA8YoWWUnItfEQ/muPz
VC0EnZ0UWB9xwmPmXWUdmWvkOinQO7lxrF2nbpF3mL4/q6YDZCKG3xwoiZKK2YUI
X98r0Hn6du2NbP4kL0IXskmNQb1+6ziV/ApIWipEi77x662dkIPiqvROHrbxWu+G
9SAct3Y0RnopqTCreKU3x45xM05KDX9AbTvgQeqNKCRGnVcHlvgAsR8hhlZ4PXML
t4JNIkhKt7CV6YEtulzjf/MNI558CsYjsItGtukY8YNzVsv0GY2fkizSMDfBN2so
er49gBklC0sHe/FM1CrDRZa3YqIeHuMKXtpdxsvwrApFsZL8zU4Xn7K5lxLzB87i
4nVmnJZ2col23tNoIzuCuPja3rfP3mNp7bzD8ZZs9HOHTBjE6UxfJ65JgdNZtIrz
zex3G0owy4S1CzDlECLG6LQFa6OD27yJklCp+NO2w8qd1gbfRE2tuStklaSrrspR
IuDy8uXQe5sLdfeVfjDofcKJ4f/LVlIHybZ1SVZhHrC0C6znySkcozoA1DKdHgLI
JFbqYXhnr0OWhxZkUUUPKlpLHMS7ywbzRmKpgHR1UJfHS/X2RBoWGG2/K1/DxKcg
0DmM192x/hGYgivD4qG4zOgaR++z3OUlliZumHdxdl9jw4MIV6mys7+r1saFUeTU
RBV0N5B5gP7A5+NZny/VSVZhjMy3PSA17u2aozC20ry2LxJ6rzj7tNo6yOCr3Y1q
`protect END_PROTECTED
