`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFmQGOSXsTeCmLe6xqy/+qrDn9u0IDFi7PQS3nBgSxT6uGgD/G4TQMQnHIDwz+rV
0+jQROV/Zpd2PkXqf0QnmJxpImN8HAzAd/G1Ns3PAWxeKvMz7rBUVeByxLFaftf/
lIiq66foFB6ju/F0HyjQ84N1dAj37z2JQqucodBaz/MvkFjywFCkKFSdyJTBit3N
LlYcL9rDOEQtGkImb065sD+3R+dMK1Z+PaYjAdWX5wQiHjx3ZZrupa6B3Udr60OP
JSrXREA6AunT7TugDDiSoMAk1pip5RBtEyRDv59vknbBuW3ZyUWh9veoFK4M59nL
LIwtAB7SEm1RiF5TVrzDP5ADJ5HoPHHv28mo7QI9+fAORuUcCpEJfyKQfDulJxZs
+riS/BLxBU6SgOcNWF7d04alFSesVTO1z+RFPfx95s51pfQp5Z6Q3rbZhk3dQrXX
/LQfX4xIcdsFC6hSoc6rcFSlBI9ltlhE8sDlpoYb5IDOCQgWxaQ1s/JcTY+CcSJ2
QTUgZRQepWHhgs5mxw2jyDHrK276aa9xPEOFQXWwZf762KgeNohNpMZuk12nC5UQ
I8gxUx9PldCNT8bLjX/+asVEU51URKX0XThXJrWlcRqjSMSLPjAww7SlwQvB8Z7l
EaK6kAyX0PBMrC6KdBnLJwvGeupfoR85ua9G1+y7BoJgYxlgHWtJF8ozrsVPibnE
cvzkwfnBVvRXpgEUwB5+jvMjDLML1Le1Ke4lomG9m0Rni3badlVh5puiZItjBk1w
MfxYDgMGU4ab2aTsTelW8yQRTd6eJYN3RooYC/RcT0GkjQjMzVnZksUhBy71iGbU
qof868+xbeJHBmJn409fHUteLyGno5x/UVZ5PGWYdolhdLKyrGrSj8GC/UhKBhMk
BcNd96I/V/lUXTBz/NbA+/A69rcEPUsy2CMS5pvD6NQ+2M0EXhlcstbOacPFvFFA
CT0WnC2GZIyvU2Fg0MD+j6gqGn9lh9nMlGwKaUyvtj8dx2cahC25Uq29QBB/x6Ey
ybtgVwLsQfCq99i8wqlhq4qMSj1jNS58AylDORjofU5r8CvlyXaOINTbLMSoGtqe
Mover2N0G/JXGyvl7CSj27Jk+FzH3ckAD62yY5N8KoHC3uGAXbUwHPckzhTvTpEB
4CzDBBEbC1bCiB7t0j8heWfcsFhiex/yiETnS9pUzWtSkhjVaoUPQgIQ8jsMDK3u
7q2ot9TMoMR33lGmy/50qD8FQD9NWKstYyTclqoxF5Cl50GTRdnZb0YWYR43q8/Q
IHYvkSripWKLszq9nY+zZ7oJMvurDib+DojL62bd5lzwhQ45UlnxiDuKakwV5NUv
Jixaudchm7tmRvxTOySbYPA04zTiDtmNDzM57SmuJzbG/IAWP9zKqoGkysrJaHPm
v4jH5bm63s2r01DBm0JUQeCIeEPH5GVeVYsZEr72Z1SFHiBdoepO0ZyZc39ZZOvy
bmBsDshZoOxij/Z+/2IqblzKy3tvvbn/dSYb6DrZUQTOF7qsKPQRR8YrWuedeGq/
p4NmXMDGFanVL1yNFkplhLwxWgY6l9apUPfHkQFutSeK6aJzOqoMESS6CkoFB/ka
TVRHEWuIgenmO4+CPtpMP1tLJQTSGjddUqcVFNgDph9oO0RGyfGmqlzuYfM6ePC3
IP6Rd+OS8a3l880bH0gvSCwOulwzj57v2imsV+6PuuPotBKf0FljJuadyEnFM3aP
GdJ/U/BkFNTSZ6lz3T7VqG8dB23jmbt8v3QywDOU0+a9jD0ceJc/SJ6iPfWpth8Q
C0wbTICK5mr/omnXe5s3HAZVBfjQoX+9MNKbfaXfScmSBuHlMvDRPsltxYF6RdPE
Gt19iSnpAhU7UmuZ6dSwycthi40+Qo/4pdzd+5a394iUTzVPM7Lmo4wBme3goUle
kNTSRKJtXeRdFgT1iHID8Qbwb17jAawH9TvWhyzh0ZSwWb/2JKXKZrnV3DQ+t4fO
T/8KIVaEfakFD74UOBsbSMlefkOKpWhu5iO34UOB3xK9XmXyuhLoBf2+xLIMHYl5
b5R2ItgjOCrgQr8AY9q1fEOdDhu/BiXLyjbfKqJZpr6EuPTL+qgkyW7W/+Jpu0vU
7PxDqCnqlu15CSvS2NlX1bf/dNwJ2FUJ6ZRKc7tqCz8UNzr79Wupa9ONNJtnbNX6
7pXYEN9dkSNHd/4rZLQFfJZPXrjd1mtfbFHdnlmb7Z15r/BMz7GKIIy6XjBJHFF8
n9iq5NMNQCBtkkstQ6Meft5M1BgsEYHWfU616PjO1c3U9X8RLce5t9+GRvSULQ15
k2dASxQWRUXIsFrPE+ujd+SS+HjDefmWUi+4TsSZ7RhMOezGpR3jT/feYtOG/cXN
+kV6jlmQfITD4fmTH4TR0PfC2i3b8DCTB4Kzk4zlfDzpUAimLWLx6uUH5wHXpRCz
JR8fFWz1ggu+/NzdlWthMLpA2miBtQeX6UirR2csGx8B/wzTt1Ddj0q3kvJG9rE4
RTnD8aGgbBrHilhrsutWNcorEiVsjs6/5HtP1yyWFmo15xznPcwiuN+IIhJwoalD
uNLz8ouKsLb1MXl7qyUpKL2bbAFCEtlLa+p9rb8xP06sDbA4d5ZL/G/8mRIgzDIW
DXCUA5ZWrvMXX/HY103HMsU+2Hw6ogR23byE58w8GwQ=
`protect END_PROTECTED
