`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wIEvy110+8mU3IibTXSqQB8NRr3AMntHQjktJ33UNi+Lo6jmnSj70MNP1H7IKbZc
Xzo399xWKNarLd3RMt8xQqfo9UNFZlRA2mIGDc0FaaYZeFs758LtPf2ntrh8vtJe
Co5e9QKIMiTlV59djvaqxHs6FomRymIRDNGxO9GU5KI+8Q3CexwlFIwh/WKzCzIt
ffgGT74YGOR668N7JiKWurEhzbmemMEBaVcNCYqzsqitFt49f7DBo0ZPjha7R62X
UhHuqfz3oX7CT0z5wzCHAIPuZc5aOlzzpEezZ0u7jhnFrH1b2QjY+DGYPZaCxHXy
aIrbZfVPhZ+87CLKxUc/yu3bIgeY8gSyQ3QVZgUn+v3B1KquI11WbRiqfNkjSSLR
hC4ciquHP/bnc3oXNSF5MZHAa77nXZD4wEo3rDcMjVWT9K9bXkHlJ5luXok64Y0A
8ArR5xWcvLMNqNDep68xKcwRqvmq+QfCKuq5JG+GmSQxRbKhKNG1En2Y81JOuSLe
C6Rr+MUdlTltgWYBZU1sn4LuGPOiu0QvwmaJWzJl3QBMnrQttVFyFwfdTxLESThA
NSW/eL7BwdmJyrITKdGNrWrQYsV99uN2pISjlbDat0mR8ti2brT8Bczapu+MLrq7
E4Qqa4UagufU4SHWEVUPwA==
`protect END_PROTECTED
