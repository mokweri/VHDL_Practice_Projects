`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxjzhlAUIlgpqscFHxPdWjpZO6Wg+xz0ASKUGDfZSV3YyA8QY2SpLjOshmZlnGqi
1+of/basAgif6Nkgga2fMJqEmzJNO9RcPoTfin78g38IL1B+NcaP5CEtYI7XgkwW
F2jcj0J/n/sKGTbXBrlHWxctfnfoxs6QDztC5yua4JnHgZuWdgr2HScMcRyfW8uI
JAzV+5vTiArwMFAwzpyY3xSl6/1EqZ8OpntBbVvCi129jUjDxNKyEav2ngZ7BEtl
EgwgcH0QTOoZlohsXq4xEqdqhzdNpPRq2hL9H19YszXOch1rER8BfmkSq0VWrPyC
u/J80AxA3pHrtUOJ1jLHXm81gMPMHwUGvMo4UeQ9ZGE3SkitKnqlqvnBOoSTcnPl
/T8z1lz6s60B6u9wj1ZJ4wVKWUWYJ5FlShPZFhHtqP6NgpUJ41N3mxdKgIh+n7+J
uV4ApIN9C6lYZdeDUQfELgIWxfkyys0xKg1aWriGN/h4cEEk1wKwIvOdQFImXsKW
jQzXNI07qlINBcuVkS4QslKH0BP/ObmiAX5BAloAlRY62QEBt6DmR8uGeGEggvXm
weJDFH2D9ql0UGuGwXZ11VG/wWcFagpnswmKHG/vVewAG6AFp6yTFwVCM1Rxkd3V
eGlCwxzZ+QEhRDsVxPcXEBvtlqjyy6hQR7CHFpx/6i/qwuh0d6gf75w/Acokty8F
KsZ+1vNy3JisVxYu6StD3s1gPNYki6IL1XRY+W47bQCrVWnMlQS7wFEIaiynnD2e
+KsJuG9tYlQvJJJyic2b9FS+JVnVzPqfEzyagdCEYYtKZF/VKDG0t7ZWWQoLJFCz
u9AuONgPbIUaA9LMh59tReAj3acmC8gcI4G1hy8bh9t6f23m0Q+Gd8nsxhZjkTxR
4BqjHMuUX/2zkidhDH0rAe3/44X4mVD6hekUKbwTp/ppFrx//CBG30CcrhIn6S+r
UJwmWUE+RZJcJjKe1OfaWqXTqmZt8BQ3KaTbcfxsQ0ltmFyyY+eAVH9pkaqTSZrs
B6QH2YQMOeo41cpn5hFMFkovjtG95e+yZUbn1FOb6dJeF0DBwUqS0feT/fKNVNMB
Z3n0lpaOA0URX8y+Ghm6Jtr3vWLBUgHnpWn1uNtdohov/TPDVk5cdL26/kw0Uxov
4sykQRgfXm4LYqCoI6X8vH3iX6ErnVA0MY+3R/c5NsaQJEeJkPU5M4dRHyEXJQRM
mu5YToSgVCc0HjOnjIdYS2lmpKRk1D1v4ar2H/LJ/N6UPtoQ44RzJTYKBjP5xlvi
ATGh3dsFcnMoE38Uyynj1cN9nhbwVnmUHjF09M3F8vVkgSZED3/jVX34B2NzhNbA
r0tp94Kl0cu/Cd077JlQbJkqUffgoh8Ag1zGz6wLXylUBprc64EJEN6iLX69kQUz
38JQom7ZMQIyKe+36BQto5AjsI2hGnrW4TkMh+tbmc283N6rBCWZZMXqgpLsulOQ
bQyPVPsaKpZs0Rkfu2kc0tkqHBpDLplC/sP5sehkxbtJWFjijGLhTSd22JzKvUEL
vlwfTiQ0d7nApT3yQ7fSmHIjBxXlOIoa9okRNo6hca2eWWrAc9obAy2h+y6/k+cq
NgwU87Z1/LLbslcIMX/1/9wMdrdN+KjjyPX5SGvENaO8fk///t+TaWo3dI4O8LEw
DMCg2GGHAOqiS0+GxNLEvbkSANaBmWkqr0XeVBk5h8SXYVHFUlFck/ochq/SYYIU
MmS8doDI5m6zifgW7f61a2V8uZOTJurZpvDOYpqI6+4RoFj3ii5HkASGGW8rLbfG
pUPnxL0BWjheXd7+flI4gjl55NnRGXdS+n/zsr5vkzDJQznkx77AMHSImvOIK1Fo
Aof4RO8GTnx6VlO9v42u4qVxdCJJcAkmYP+33fInSatYPO6r0RBizocwI908iT8O
7JloNOtf13gbwfaDNWOtBCamcxFC9niM8vhwyiexjkp31iucO5Kqvs/8lM4vGe18
BTchYKMiQ8HP3lQydXKnI8ErTMZyNpcZqdsjuYzmg5tJ7b9abjX8NW3cSujm0FTo
SGIYvYJUz3YtF317ECqYHqTnIGiGo383iTe8ZM30Y0XYbjbOvB8eQM5twOjiEyKp
Eili5cSUNsOfFqA0yxoe38BuDruQRtFTi+rmplKTzia9Dm66ou3vJ7JQgKnDUyN5
pmiKDJvwIUJN995+Qc/MIwPLIY0URuIw7W1s1xcSWYLK5Gnf191nEH5GJoo1NjCP
mQSj5gpQZcsS9Gny+vJ0yisV1sfhpMODKJzz032S48s=
`protect END_PROTECTED
