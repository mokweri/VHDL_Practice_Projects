`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eHI2EYoal5/F3FmCL+Kc/KO+ObI2c4sYpS9YGh48JbEUr2G/KIy5i7Ye5LAFAZba
tvHbmJlvgs+S3iLLOr5G+0pV9hG8p30CUmE4zMvv+tgtmUtlvLwmJyHhfPgLkgu/
5kSRl8SxLIZz4YzC3BJQMBmsjBiS17uJ1wVC+EhzqOFZAfzPkBGI7wTvMmCkgGt8
CVkDMlE/iekgtaeQDijSGWU1Rxo1miOOycvQICaPtf0N89lizzzLCjh3D9pZmEo5
OzsecgMuCxms3swZ7KLi50x8K2n1XwtFmB5iob0nRFTBTeJnNq31IWNYyhbQ9OMo
6Ntf1BS0jutQsrLcAP3tnakdnPW49/BXLuKKJV++++KTwf9RfbFCuXTnS8dF0NwX
jnuPXOYcnWHOdwgFrTSbVUihh31wDQLyndYlOFg9YQJxszF6AYZK+FzSZLgphWnY
zhZakwCNNGTT6HHG/PWurvVum3GvlKMKPL/ifc4kyldPekRc8nyEVqBhywZoqFEu
NqI+B4xxK/C7IMcx7jPScr8pR9BEZtQMV/woXNw4NKM8/XAarpAMqt+i84Nrz4nm
Mjqv7VTfvzbHm0WppxAV7Zi0OB3UDoPJ2OzTRZ1ewOeyeMTR4djoTWo7S9soKN2q
IVec0KpbkMRn9E784wdD3EB/HZH4WwV90OJyhvVS/h8xseM6FXiCEZnWHma4vuB2
ufteAKJ59dsCn5CQ4zfZ+rFMrttI20zDVUpwdSRu57KCZlrbD8O7xviAF+2bRRwR
zy+BFPnEmy/bJPUqEatbA0Kin4/3wi0LmiufFqeArF/4BRuKL76EpUw2AqRYMneT
SQL5e0TBCQKhE6RUESzMQyIYiz4jZ4ao3InRaktmVrJF1iVyi6WHN7QRyc8jbSUl
4u1grvuVvddQV3Rb19ErtT+Zh2lRQCzWypM/5SJNRM7q9D21N84/TnH1RLtJk/de
Sqdz65qQtuCBUAPQ7kkdA5Yj/zw9FeAGxkk4qzZC+twC4Xmvw3Mo0zVXqCtXmeDc
WYW4gR4WR9ltP9npfPCc73Ybxc41cK+92MmR+k4Lr59rAB59pmScp/Za+/0SyIux
+uTM7oXxkUzbBxhhrkkLD6qPA29lGUERjmKLxbLBAwvVi9XA5rM5tLVp3h7cLDYH
n+an5uaPmwsIOqUUpUHM6CgBDJOD6MfwIcqO07t+jSd3tahpwGEB2xQ9E406qY3u
21OsXprYDv+st5lCKEQqlFgaKRqHjnXbBHSykg2NBPMotDha/LKMyW/Gdqd9CHtX
0CywgZVb2b8m3+o46Su3+gLKxWurW6YkcgCDXs+21Czu22Gx0dTIOLK7mp3Ux1on
n8y9zSGhTOxx/Z7UkBs+7lDAdfmLI0+lofvR19bz4YbPtA3J/MPcfybHoJi3IjoR
5Wvjk/rnJcUpfPZs7Nm1fJkukBeF04YrADb2Zw4fvVev3wK6eGEHbyzX0ghJ/Q+k
mu10W1JYIXpLqi/eqHxuTHer/i3QoqGhRpHaJAx0V90nhlOYVUguuDqx1S/Voy4f
8CoqcvbV0WlqBEOVI14EUqH1+eQwATxgN3ym2qarHI7VhjyMfdaiGdv9bCgAjdGc
LVSOIOBZuhF0hCLrMh0DCxn6H90bwRCBnVWpU/KiSRWGJp56TUSUgsfftTPYai47
tAXH2iLYbA7O54v+1yUqmOwkAEFEOcTz03ZnDjcTiJ+UAv+IfGlDkPerpuZDIZYP
MMBxBJQeNzxLslvgY3ORkgGTguyzYcjVYPT/cmIlrNTsbximtmQehCkO2n1yqbyz
ct7hECjQd092mPePRmBCsgG06YAJTfWYp8+B/xUUvZUt/z1TzQlIw+Fks7KOjGH+
AjoPCRIFHF7O5LQm03phAo6xZyP0x5SZslB6CyDUZn3RfDj1sKXoWmVNY9ZavYSJ
Bsa7hs83V1sWSNFDqO9/MlrBO4grr/o5kMNdyluST6aAlvfmbfJ7QPMXfTk+bNsM
t4LUqs5JJt7HPECHHpgspFlmup/ZLrJCl7ySgDDyH5yb1pBTG+F+NzpKi9M88Twe
O5W1PIaJ2zVNeuWi32uqCw==
`protect END_PROTECTED
