`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eMb93D4ZZcVSXRf7gvQB8/BEHcGDm0SjMgZYWXN71qgz2rnR2XOVnWreHrlOuY9
Oipehfx7dFGmeKaBxHTOGnRuzuBg0dmDvXJobrPeTvo2jE4/0Ne243vnzn7qM0sc
ddKuvvhLi6i6WEALn/n0AOF/9aI5H/BQDGBZHnO8pHlGgoacUEwr69f//Fj/IbM1
3iOPXrwgh6mbadpPjF77Mo2XPhPl9tphr6lV/rpqEhKVAoVqH2nQiJh8JCkqxdmC
N7G82plPnpgQibX82Iy5oaec+jDSou1rrcC3o6t2mcTN7rbXWCSr5z60/ITAza+q
IRnaHdDwsLoVr00k4GxIxbFFagqs8NJDwpp5GzvxyyLcSytXmzlwnVq9lMma069R
L5KUq8i3o/lck7n3szTYK/zFfylG06lJp2zt5PssQTvqpHTPeQw4TvfOM4VEAXB3
sBGAejSW8FngGKZMBrfNz65AbJ79keIjdYHClOKSjfzp0gHH4QVmKNQr9NzN4v7n
Ljmgo8jPd+ZLKvrL7H5WOygb+nOFr7u5J0MeNxwPag7cLMNt+UeRv2RzX+9S3Wyw
d9M6Jy7GsjSm0SxPTj/b9qfweWyY4gu+xHKkH6+EcpOolz2H0ygOZQOUh7vU9xgj
1nYyRUSTypbEXczvKOTxxtCFTPjJt1oSsUM/WW7EUoJExqIQ6coQA+jpRWnf/D9x
fNgjqa02ihwBwmGvbTg+hvS7LQgqu5lPTgbxBs+jo6YFygDAhiTPhyXp1jQKW1on
atscM4ROs328xfEi5Gjud35B9fGOZvNg8V5zjwfi0393JHsUi/setB6qJ0leIiNW
VTCSJoTEqelr0agw8w0hHDPzKmm2tiE/KEvm289VIRoG0k76lXj8yoJ5Bu/kCBim
um5ISEY64bdKMShmsXB9YJ7MB2uc8gcnDATOtK9dpLVIYrFwsTMVdUFGjuaERdOl
`protect END_PROTECTED
