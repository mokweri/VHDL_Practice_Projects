`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWG7LhN9tUDSI2RjkxNEkN43stOUlcHS0rFkHH7ART6oanDwVfkmtiI1Ke5lJcjO
SWLXVzckU1IJnNc1Ihcwcy5rCJgQk6tE0MjVGx5aKwzYwl978mhTsu/28pSLZBGk
1FuynN0sDCrcmTAbz1XgRxseAcECU1FS34D3euYcapXocXvxi7eAtSWqOx3FVZWv
9tgys/yOy5u0aSMdKfZZUndZpzPHwsqz2+QnwYBDSNxiWK+yJNzQfxW7RY31uzUy
4NpUpNXPuQLU22IE5mehmxjZSLrVM9XZdiCv/Z+I5uW23XLPqNoGJfHY2EwKz/Tb
/b4ZOAtIYf1gFWa0QhZ1axWhmW9Ei50B9mQe4C1ZWaME/hAuIi/TClZWjM69q2BI
ynVypTELKzmbH0GLAGFjCo2GIwKMkv/BNfAa5f9MqZMc+G6AeAMqNURj0ZmSiuxv
xDUrznGE/5XFuKTfa+T/45Pzkauh6zlam3Wv53xLwJziQlM6nBYJD+G2S30FNqQm
au0LZxFbzzB8x/2W1b5k+i7wbhftuSyUvO8bSQSzjIfsdDvZVlW9/BKeuOTDultk
DHokrjYz3uitMtZlKiuA8uq/uclj67Erqfu0b+BTjY2bIpP20yRuEOeOZfqFF9Zf
Qfxz/JQAHi3r8k83YLfVXPYn+A5XYIBwWj8dSthNl3LjRJ2L4XWyrcsnHXOR3BVy
cLi/Cehnydy+RZUb6AB6JHwzs0rG6Hf4kOcJDPMlNjSWRkUV53QdLlc8jXanszgf
tehFtZebzcShryZu7TOkPDvQOsnRRYED6EJbZaTUv+95H7JaRi8BqBq+Vcvouxch
kcyTh5kj8TtO1qJ0zM0l+B2aFBragjWYDRNt8sEOkJ6Do9/nhU3sdsFwU8ZtkZ8U
BTIeMuy/99t/3bw3Wap/UUICAYLz6fBITzArmAD2BAhQIcsHJoJYOJChfwQIS/UK
0fDIJHu9tw855QGnRspsvASMRozQoVXFVNBo5AqA4zuIzlNQcOWTiRp+Z3K9kuGp
Tf6WLok6y+etdACAg00NiCT3QV4eNHaSaVOuSy/voshDG+cECWgKoUtMabNAcmxe
`protect END_PROTECTED
