`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUpIGtXrnK37izzuxFopURubqDbZ/kDpPkEvfjopVun5z3IEzfeP5IM04S3rtxwl
mURgPxODU3K7F8kqtdW7pnkdvj3DHzodFqqWAopqU329GCskv1612R2qYRpPo4as
03RtxkXjLDzuOrXhUc6loseQQNuHZzmKg8ixge13Jq4h0Q//BA9UYR6Xuedy+YGg
sqymRshrpQ2bV0L9P5Dnp353w1hUTVyFGVjB456KSceqqOJtIfQu4ZbGbxsY++o2
nxTZ4y4YCsWXnkGFoizoH8R9mPgSeBy1OAkj/rexAsDJnH6KqWQ+ypSbtbfa1Tv8
NQ/b5Xk3WqqEA7rEA8KTQPqwDXkK28mb7j/D+qpz2PrwOYQcAUDn8W/A1DEc6c79
T0c2TQEMlwWJw68o2bS2xikAcC0grxLhUgqWU+hinLHrWz0cl4aFGk7N20CPGAnI
EwuJiTe3AK2lWxHBXFZF6tRvbBzETDWDTZDj0eYlDlRc1EQSsxaarDaDh5c7AVzx
lD0FMLZ6qDdeSL73GRyORHPO948q7Tf2KMZMEO+u7pfcOk4drVKzwLEBfzklYDso
YIPr2z7HdB9oiKIVboMFHgNYraN2xPdJbK+kXBjzL4y9fbo2IfRjdzWaZOYlAkYJ
kDSctocV2cjHK2vqofC3HrhdSM2G2TGO+DwvkEAIp9AGNFSEZ8Bi5xMf2gE1gRZX
xRRhcuYfGZ+B26twGBcPCfthZPJ3kfGMqryk5TyJS5N4j4rESYP5crnRpECwwuhi
fMTixMGFRc4aufoyHxvO0QEbEyGdr+NZuI58XlFnl0abb9HJ34yuUdCCDb2OplAg
FZKBsGgAIkKmDhhyZllYltFpxEgTVpyje3wgHYgreXHQ2RIKEsD+3xm4KpUquoEE
9o4ujzHVIfj3fezlnrvsEfhVIHydniW3FhT+X2eRZkDfs4vxhFOQ1OFWIlawNFWi
r37itq3tVxVFZ8ngeUjXPp/xIp0Zq0GoZEvX5Lvr/n43e+0FHafiRtIyTTuZFRAK
mJrczY5tGhFEtPNp02/TiVA+fHI74kO0rj/atVZcntuc/TUwgmA4jfSMAlCleIkj
nSVlvGCVC40V0n02L4sBj2vjWDKie+FeLLL+OjGtbg4YQB8fzr9YX7W96yYxzZHH
AogOJrIX4dJMX8aNvpJYs6tTPi5NtUdzVYbJ684pDW7ZzU0icd8Olz2om+3gxNPi
qByojR/oZaINO/JywYuwdXRm5ofFGkQsDjbj8BUnvCbbcqXCMtc3TlgVbxID6u6R
57IpYmB7Slzd9Qzp82Mgah5SwrBwcMl6maJM4TT0FYwaMCun7rmVn/o91zYx1bej
7V8toq0dcbR9+ErpZdduRVsS2pY4/CmIxL1/kt3BTjsm9tDSrY27ypdqIa3oLFtm
KAJ253RLwYhzFzjSCALDBf+cjngPSjxyC2gTKqX/pGZir1lDbcHj27ZHMKnjmMvT
DWsCZx+mOuZSBjAlM1B/tlQsuE72/fKcW6elobO+oUp7uKLaWB5lLf8eT9ZOgfTH
gSAI7uJc50RK4plzJ1o9uWfsN8hEJoujBB05Bb4ks1ENrUQQg3+lzaVR2m00fusO
X1XaSgR6qwZ8q+mvzB9+KP0+EEzyWueM7+6cTm46v47CAwn5Y8W3ukzmS39PUAue
t6J8kbi3MDkc+0k5A8sjSBVXix/UV5FGjXZx/7b9XQer06WHERB14z2Jme72bhJA
BAy/QuJESGOywaRmwc5DwSPQXvK5YaSo0cNmo/SwLOd02DhnAbtIMLN8aE/mzQCZ
RIt531C3kFYsxlcFM+yTSwIf8zP8tZRxmKubJBp71hbQimuyxyORIMe4YqgCP0U+
9V1QCDONlOXnoOSHw67qcZP4DKMN2Y6+Cp/g2KxBbqSWQO4vGleJsqYPWzV5Cfg1
HETz0AoTvGtkW0wlyzBO4blRjl2Urv57nbmOXtitI1qKtoXHyTNJZxWXHAq7ZCgu
UgwbpkFQ+yPSuA5/42iupgo4wBZnitNZuBuZ6Jj7sHI+LKZFaSbvHwqFBkcaXwd3
mBUQ98K2KjW/8KemLVx9xpg+fYnLfcsRU1jdicQUWQctyZsJLOmVLoDPehKZOHw0
WZSGT80f82+dscTtElnUMx8ANm4hBrZhFz5ko76fuCXg9Zl6im8ppcyW+wQYhf1l
3TeeGR7veADOoWzqdTqxTJnAUNOZEfjAedhyDwxeBppjvawCjBQQNmwqqJqpgOrL
bWwqDh2EalGw86Gp1/gT3mY9MDz+9TaVN/Lq/RgR6wkwHEHVGGr3HfPm1lkDd/wG
0+q5+NbNb7rPOpuRWi1yczxlmpYRbHWk0xYfe6uwR/AnyWJnwzDrKWXGaplgQt3E
gLvNyP1c6lSaUAWFhHBOlYNA3i/XzazGaxlIJAcBT2MREM2JHTHDvF8c4EfymtFZ
xCeEW2PztDal4bD+BvSbW51BwAD+P4Vmvk1thziigmNqsGbX33F84kot9M0j/SrA
GV0hQ19PUSV4F2sDMchVGitA186+zIQ3YOYfa9AhfrOJcqK1MlN4k0uUA2Nrd6gc
aW+MX1PwpBCLQCPwZKMCRBVIx2noMoHXtiJ0HHwV3uUTeKKdAQlNutzdgeN99ps+
hTPU4Y9HSdKOYEPv9MuVdRbWKQblOYj1i/1FaG5MtoEPRTuQdY8lhXiQTNkkZUxo
1p3jAmqtOEBZwuvgoNnx4f3iJv+QwqIncImobq8NWCRAxAu1jRTdIJcQN2zVhpbk
SoflpuBLG7jGhseJmZ2vkm3S/oF+2/15gWYtI3nLRs4ynCX4VJ7rpG+axPpPrUNC
HVHb3plkFf59Tb8BtBgdl9hlwp5t7CYlVsJr0p3GTeqFsRcfNqbInQIatJ+Ly09g
WRerr8HRCBCIoiAksXtfpHjh/5Q5SV2LSu8I/cVBQneIVQfFDOJqbfQqoFGebcYo
7Lvqa/YZtKsoVdovSiAu0Jk9wSC5vfrkHjS30/OdefCpAqX9tvp5aFTVzTPmmFKY
CKqz9Zov6b/YcoB8Uwmx+Wi9h2ZsKRctaV1BweKOcSZpuP/K7cKVZ6oFZcogv/nt
rVPtBmnW5/aIOyHj0jgzOLEm/nDks5BKUk3Pczb2F1bJKECjsSArhr0rBr0ICAoK
zWTQQn5Dsu4lEuP7buvsIbepOHq61kbWl3FancCtrjDCwq+32wD3iiY64X/mTceP
IisvPm5plaT/4MLKpNzBqnLQ5RtwNhbWFmW+SxN82Mima3kGBfjbBgaJN22yoldz
tpBSE4Cg5UPi2xZTq8hs0RMXv3egJrmRbuvEXdPo4zh9E88UWrEuPi99b2L3Z5Yh
2Vd0l4oOwO7dLZ/vdgvvdMWGSgJDsMKyw0cb+9l1UKEf7/4U3IAFvWX40ypuOVH0
4EP1ifaAxtCVGjJ+W5+ghtbzZ3M3y5c2BKvHPkuaKsuoNRO9+QjF6zBB+NYtq1q5
l7Ji2ubHgnKQTrn5B+rBpY9Oivs87SzqLGJsiQiQ1UvFk2naqaG9h6Ts5AIRRsst
cxSovhhKYDIworyYPkVT+DkQCNAD5nr64W5vYc+zomPMAdxoeizrgfXfsOv2OGWp
6bgoMrJOdwk/U21dMQT7KKEKTulo7UjjKemB39eyzqbNZveqRxUZkhLhG6sh0Szl
EIU03NJtWAkHG0pOmRwW0yaTyCRrqVLIdx1QNQ34w4bhhvrXHMFCA/N68fpPnhXP
FExSZspgxiosfp3clEDv7w1aiDBvgqvktUVoirYIVdR3vOV4xZRacUKqcO8EWt0p
+EMW5gWEMdSbFbe6A++eqn5zaQ0DcuFyOjyFWsdOwnM1G6K1VdvPcg6k4Y05sGeY
EYEJ4Op3vdVPp/Y6pE1Bm5Rp7hovrHlK7xpgak+gBz0/1f0CjMAaNAjKjGdkaDVn
HcwCR6RFF81eW3Z+IOyEM4qmkmqNKgAZkEGPq01pPqIQb43fHaHx6+fgxNtrG7ze
/kj4rsI8mvMA+zagklnTLE0fgWWXuyCKMlIKogR0Yv8a2snbMyFxfguLgw33dGrx
qhg1PFU1aY3Dic+iiZi9k6WzeL7+Aqkm22csdrq6w22P9qlocKh1xNjxnR0NXS55
NqloeKqOZwJpA5eIV6I5ZfIFxCVtdCofzuHeW7bzbX65VCAilSTsfrTymF5aYZgC
1XerO6xXZ+yDy0W1TQ8qRIzio8wwiq8lQkiS0lu4sKfzGHvmuUV/XLUmLagg/p4v
ErzP8JXEQZJtiul7cbc3xC9GPlaMhOje6g5HgBcZkiAdBKCvcgx9bLiTADnkatRe
cSRvmGNdbIMqn1blLOo930IXxoEvBU4rAJl2/z2HGG1+z9JWjazy8f7g0wR0Tb+z
agCIAcKj1rLmZfSVQSQtmHc0VaXQtQ9yi+8VWL0tnjBQAu5qyTmkiytols3jRWDi
0AwofYF/UBde3c7et2BNYF/lRTBpg/1wnNCv8KZpFJZzedurdIKoPcmq4I3SUFR4
9KpzS/U3wX43y8BF3zQHLECSWf9o7NsKTrRX+ngzzjWNYMKrf6mnTTSE+LRxbG3j
yV9Cqk2i3pCXUWVJNbc3pPGVbwyjr4omRZ6iHPvSSggyfzRE6SphLRU4BzFJaV3y
SulWc5HffJ8VPePcgpc7Qsyi+ePjx9WKMB2PcDRnignywTxeVYS10aciQOpZt0ut
ev9kMPIhMgWhx7r9ezozbe7tRJ9BfL9v8CRqbPfgRX2aWqUvJGiseeE2VfuMmzjv
e/2pedm1Zu52igbxNEhG4nx247ohWT97PR0iDxRTNmGBL0Rxc+vrbNIqSZYQijz4
FmbIVEl8rsWdQocGT+A4p2p7cUgEBW0ALlSkCjhyghWP+YKeqRndl0Le+pavvhZ/
M+mbCJ4ql/C0+pADWdMJjI4PKGaYqdqoEXNTkLlaRPy6kjLuxXMZmWqOkiy8VOfN
GOQZQurHnX2WcS9wFAtm/YonjexRs/7Hh6uqrujJkn3lN9vE+krz2WWwlVW6c7tU
z3maUfTMsmAyFdBx450DJK3EQwxA9TXf7cN5Fwnts3FqeKQ8DiIr3pRoPlGsPPOW
GiB6AxTtssK3u/ZHVYB2t0jAezW5cG1oZ/GlRmRrkMRIJdmRtY+MbP+bwTQGVgpr
N87CBz80doyWrJWeErEuzBnK1qnVn2oPWbVYJUUAFsDJNxDoX32I7A3zLWqsdiyh
GZWQT0FFSD8E7VeHUriI3BzyAjOCHHzdik3GVaZ9+GxOUVRrc4TPcDazRatS3h93
+s6WPjMRcxPwwIBDmo38glC5pDAWI7oZoGT743j10T7bECdPJt7+NjwTWLBETsC4
3M9duNGhetfd/iHpIspdk03ZF+sVZZH8nTPOyI0GkXHf8GbFZdrp4qLSCS0WNxy9
x/MbBPjJjnO3cIGu+Ev+PLSPWX3rFSq8ZApYPnFZNsS+Ux+HtJl2I1Jb4qT5pi0f
BVxBAywVv1ikTEoIt4KCnm2vc73ujAkqY+YSTDXryQJglUlg/PvgCpcboRRR1538
CWZyESOwLfeqvn1WvMX3SPQZuPbMKkz9UdQUOWbwPXsh/15D3xI7kXzf9zyEcMdJ
AKDGGd/WVmcz+5Gs/UvilXgFg5k5Dezo3NDFB84+ICiLm50uPRaTgP2YFPbjhd2d
qq0DmXeMXMQA3WFiKlajdx216XbLHfnwbj1H4HzcQEMdMJvlWe8+hcERSZqGfSf7
r+5Rsq7qKnvProWS9tnQEuyHsg2o+n485YoYEIxyQKKaiUmubEk6lSmgYn/hdiJx
vjRept4qHrOhE3NKyjW2Uvkad9XqjV7Ex1HsmUiSUwc+hzLorpdk+6vEC6+feSvS
8nVjZODRwHAzRb+IMmyS8eroMQL1lrd9XJU7FaSRFup87ugzdn1r/VfcX6N4bA+/
5NTYjvxgyqKeBNVI9ziiB6fOx+UsKbubwfcB6KUtfHXlZ3BWcSoR45bBXJ6djVxT
yVfRlQP4FCQrzjnxqUNUcnsRQdNs/Ch44IAsLdbIyYfo2AUctwCtXG9D4S+HRiyO
n7H1FHX8ref0iTqVZJEcr1FPg87FPxfyzboeKL2bgYINDggMa/UKtcQCgAlh1/TH
gvUP8Ct50zEHQC3k8YQH39Tsj27n9j35I7r/CxAW7OatUf1BlARYjsOlwBTlBE8k
Hkd9gJUHAm/QU/kqwcf4GdWWD1PR9h0d9CJrlkMUNFhyeOy33RLRKt0oARgORUTA
BjG1R6DBrJY9fYVxhPBBmu6I8TToA1IUG/zDiyMHiYpTRDBzfxPk5isfSX355zV9
EL+FZpZrjmi9UO8/133/8M3i6UE1DbMBQnkRnO4+6lfZ4mpSI30hU4Nl4cUcqE3h
K87Tf90m3G3qR46oUdETeoVvKFrWr8/cj1KitzwdYybpWt4Mo6mAT0cjD8JRUxvV
bS0aYCpZY9ztL4QeL7CcxGAqM5dy1+yPFViq7Q7v68Gg/y5sRegmXDHSbvmG0Sxc
w/8nFGv6UfInqBQBes9lxpxHtAH03K/xtwIMzwX7q9p5tv4EkifdPmqPK5ErsdeH
pPl6kzYeADdybVFLlSHo1C6DZwcRohbKxkqi+euwfTMpKtwIcQH3sNFEBcHk4cJK
3PE09497vvdDIVqLfXsKqQ4Bvwh5pRcaj6NzeuL3JmFD2cRM051keJzSgmFBeOSM
zuazDs3lugl8ayuO/lIjyzEKL+P+iJAO6aNYDO+tP1/HyhPl6N9aVsfmdE5xUs35
3uaD3BM5Xkl53LAFxJmzI39EEv1iRXIn0BAok3DqWYg9f5LfNXF5RW58wK+jnjvf
b3BJJS4UZ9iAokPaViDEZgPGZ/QEx0RAz4VSqOtd5GguAThCHWWnP7xPrGu9ajRp
VxVYlfTN2fmV+Xz3xZaoZAgrvg+dNwHleqwhi/HL7X8PPDK4EAuOWPyVGzO1+Uuy
om3j+zpVvnVSwjGXrPSpB93wv7DwycHA+UkrG97u+sH8pdy4BHZksPCbrR9MbwDf
vUiF3WgqSuCFm8o2Q0YPkb4561PlbVMrE4HIGRmJgeytsg90emGafAwshHOgOVfZ
qA3y/4epmWkdnds7har571tY11EwU5A+R61G6CYZ3ColwNctwYB9Xkbpb0eN7fsw
BhSIXzv+JQifjOaDE6cBdyGZqukksTI9/LZ8R2GM8AyPGSzY6X3OWGSzwgLgFPk2
CSq3T6OUvuzb0JvBjbzyQtoeXq+8VofaD3ZeC6aAVgsssEAECBGBATXGxyk49u4a
TN6i9fJXbehctsXX63Z6Iiub0cO2dzqFJBOgtqtNdXjtiDD3rC6ppLzgHlDOR8Xe
fmnAUo2x2LkGommT+QRdG4pxd33CPeuto6f/hOhVOs0MdsJ6MSue+/k72TwtuMsP
459DMQJl5jteWEI4U//KgcO9n5vaZlQ+M4JFCHjXk1xH++OlKu4ZNvZAZzWMxq1V
J3CW0p/s1qYRqBX9PrCkvlZOANcySSH+/i9WLCQwUtRvMX2w2czjIgLN5RGnW4Yf
tviTBlSSln1ROsRrt4nrKU86UlHM88Qvb/zwQ9jP6fUVQgMcxCbAQLYvU3rbO+LQ
c+dsyaaUxUAE0ZrBa96TlNGvQEGJrVyXCbHC8DddXHuw6B+XhN9HSEdLR/ppg5W3
o+4bg/7imJ3W2fJ+aVucnIUwgo4Bw9uQNxRTO2YNiakPEkTk6K8YhNdeR/1sFEib
xwwPy0uKJG3Gu+dVZ8qwYi1cfhwGzc9rjOyurv07EV2mSQn0lMrtImR03+tKaHAr
Es5hysfZ2me+BZfXqgPBuG7ZPkNbh6MRi2PQK/WLHIo2H+xFCipsW5IPjMSbwGAO
JbH0JwXay9lu5AKUsf4OkcD+xvo2bTvHzAWKZkDVa82q8fuaE+PX18/PWaeHlA4K
CtfY3YEmvNGBu4qezDR3062Ha6vtDvCEHP9Lr7UCNFNLmDhcj/RN+UUM0rOUxrJr
pimEgi2j2Umgq0XxYhgc2xnH9l1tSVf/+nMPie5xT25ZseELTbJojMfHf+eR7eaj
TIWjuivyOrj4Zh4B5NJcdyCis7l0wkVEkcr8tytAjE8HqiKED8EaV5EXWkuBnSwB
Dl9xXfstkPz2YbEhbtZE1lQMPaoDXFnsVQNRuy6H1bruC6rnNsRNrCh9vHF27qtf
ctXQ3b0JEZ5tba56biHpgIwnku6yHJwEPmEGkGvb9zuAXWKq2FdqxITxPUFrLgIW
I72f5WHCVwTLk9htK5cEpwepVZSQzARn76Mf7T/jjLGklbvWQ6of6I4Q7BfRjV9C
JBdudCnCTyCcvyiKjWLW2XFuZS/L4E1940dGBl0Kmn7pKTTjj7/CcAWSm5hd5rrq
XOGpXgXsCnXXBJiSjwCzF5vb6CPCT5CBNcHzPF9UOG2w+R3uy/LkFSjIMYzZYC7J
EvCFf20yBxxl8rJb9mWa1NmHYH8Q1O70AiTXk4NfCCpL832s8Bi0Wd4UJykulArz
L9No4iNjN0JjbLptKNogMM1uNvtfivJI2ANAmb8Okbn8tSfox1yQoz61wbAqYvQI
Rhu16dxUMnhqRl1mFLITQBjcmcKe424W7zx1dbJ1cPG/7JxOXheSGAWR9bAhZ1ql
Zl0LchhVdvchLULpnewVUSNAJwUmwZzfC+kcyNDoCwPNCPF3tOO7fL6K6s7Y01bY
6+aUVPZSrd8j7UkvrFW8l2EzkZ6DaGRhgmOSjKIGFjcHMHwwAVPNpD+dbpxqTPgA
R8tD46cK9UN54ErMRAd+kEl0U7GKH6K6sRO2VbP+I/uNfjmUFQnSIXPQWd6HkvaA
oLkNH/n+3Nj75EKFGneYoT7M7GaqLmWeUFE8xS5GoMOg1nyfiZFJAp1gLVVKzYXq
yHadLlayqwm448SKoUVIFaRZiyOssiCjbb6WrNsTwKvzqMedyRkSly1EErP//m33
55c6CJiqrVUelrzzl6i7EjxVTBHsXgSJnFZIG0BR93cE15+pmIHfSYFFP64GvKED
yWtC6FQkDeWif9gxEpCl/zKw/mZU3w1dKYQNqa0rGqcUsN/cLmtBbY3eOtswf1al
r7p2aOW/1qSceXbxBqxKah//gpw9G3SpZdZk1CKfIAGcJCUVvDxryEE2m3MWmDUs
bKvLKk06gBlVRR2Got8nV4fqT4FkWfPu+Rnk8BsAfg57rzOqek4IuzwB861c/Pog
evrzUcOp2eVyCYPT11DqAg2aFNsH4X9UJsxDC1LvJ+xIT/eH4+Wfy8LFklcb0knU
0dQKASyFdtqhrr+Fyst61AUVawSA/TldPZFFYknqY08/wCeBN35ow0XCS/9jgsrP
p/jK6/3wCHUXUYLlnXMfrRPaAs7nmjTWiKf5DStSfvz1ovn9g334zV/UzT/pUbpF
2FaKzS+TsZcSkaPxlx4bEiMXWgvrR57ptC9lwhmdAsXPiqE3riXlPPSRnnaPmBLj
UhcnsHuepWrxFq4dXddIA9okQEl0uh2HxY1TNweod4CA9jIx90Dpyt53kKRX4k9r
J7d5CDRX2h2IAIjzs3EXD25TgwTIhBEJ+dXH1Upa09rakQBTdzt64iLID0WT7xLk
7Yg2wKyt7pzEQ6lDHXaYJqBcAsSscJHoLVrvAmHL3GapYETWYJb9VepOIRJoBUdp
9qL1PDDZf3GpO7U7S8CnuI0AKrjD7xKVRKvfp+hk0RsZ1ri2WCyMNQvbNNw6Ya5U
0GXBGohzpAHj1GhNB3KnmqVpc4jkgjZ96sKMC/AQ2tt5YwpOG+DaT6z/2XYq1fOb
KhLpBgnCd+IbiBdPSRNn4oq3+FOsMKP7e9vblusY5H6LSRhTL2c3N63rfD6Hzllk
+DXyohWZHvPQR3ct3YQ+eKJx243dY3ie2vWM7GjJrKSRfEfbFhDN0AB0hG4O5nPm
+TNOk8wrzdDfuwpk+Y6bW1Ye8NSmvO6TyiZbE0BgwWQOMK/rAqfj4kD8Ne2p2nSL
OO8Y2IMqDb6ZaowcECSzLTXScjA8DfabgxLVBtKv60Z4cO4eG4F1CuiadIWJBnuj
MhwEOxp8R2Twoj2RTmUxHQeBzGs7Cdkpa2cjM3nLXMxzqaKl4824JtUgvJMZ57Rp
cHAaWfQsJIp1bf2fNEZp5vi91udlOOQEwKp5NCtIlQFZsE/RhT1kg/SZd/Wy6nMi
+eY0D3kQsIvjmzKqI27MlttT9vrJOWjxucM/ULNfvTBlMaQjjSQrKtRFFwaWFjET
6l0nfHbSFxSXY3dDP7QtR9RovkWtMC2YZY9283GtgjkSft+Y6fkns4j4174gMie9
zAgsIezrVrsfogwfkY6yok1rLtz1zNmcgJhttvrAVlwTqU38EdM9NI/cQWWU1Lm2
jwsfwcKqE2O/ZTMV5VW7F+I7aQlRxRRTb8l5sBMwbLWFdY6qFggGKHy6/oHifbme
dlTMP5HDyBeOcFBok58rebwG7pByYtySUe9C0dGSSwCxL75HVhVrw8+l+S7If6x3
nWQ1CnvomK4/lRhq6bhSNzyZ7Uktu27KUH7nCo+2bl6N1UcjZBiDOkTZAWr4/dvX
Jq+sSYjwFFOZnmAV0DjHYKDoAASaHZYEYR8llt+o0cyHN6HPNlHgvhio2XonZogH
wszWMzxgqM9g652Cm9+FBQIM9OUdV4CTO5UDtNawujaerr5xA2+09tOr8PS9IBeg
1oHgGlpC/TA4kKQ+Wxn4uoYNr6DtKzjzPyjdH1YJ3u4TviNpd8vVf6E1SLbxBFi4
bKueP+5FZO4Uk8PHp8KGQ+gFXxpeHBJcLIDc1mfOT3UALK5C0OsPs7YzePUdcBXr
W5bjhQsFRNfYPdZgI4LBCq5/fwn/dEOSPiAo0kZBPVWDrOF2CCyFRNZGDeplYWCe
YMjFze/cRGpEqFHZiN43R5uofuyZ3kpNPYHbM3eDJSnVixAm1J875ug/hcv1Y5Vx
zHNGZcLCRhGs5ysOG85oXRDtJtleZOXQfe+FxF8OppiAHUtETxy58oca4r2Z0d+m
ZOSyEy/iqBq/dQ7Lu5ryg+eQCyu6gbJuhv2263THhYRNoxjAHTe3s8WnEy9iO1LA
jB4wyO6+L0R1z6reWCgndymiXhte//dBZ+XALwhgu+xDJVnT3zTKDd7Pnm0xsb2G
H+PpkoXuxV+AWm1ConEqtRcCqjNL/XwWHNezN+004642Od8FaSvBal8JHFVZV9gN
EiaPrOkDEUm1Yvb/F6HTbSszSzqZ2IAzhUIPjkHllY0VgJpcJx8cx2R4AeE9B9vC
I/TYjFkgDxtvR3nVq5cdpq9vnAWXwnrUb0GOWt4oIjcJAGKIyjx6PYF/CANawsdT
5kdwCbadQTgg93QCjfCCUiYNZARfW3CLm+Oh023Zts1XSq1wupJsyhGn1RHShuXE
1fSvydZURFN3Q4ApPNIhcaRBIQwbINBBaAvltCE0agRFb34HzaDQyt1gv4WDn7Fi
SPCs2wjraiY7TO5VkLUHbKV3BQJxNQwbJRr81cQOX13QE5B2ExhfHR6sjSDvK1Gh
bJ0ffy+hFjlftaNC1CP5FhTqK5O0IsR2NXfX0zL+4iKQ263OwCyxMI4KiAXmzWVG
LBVpOGXr/lQ6usQYT/Ir5Smu4R6ImqdyNFGzzzhZigya/VAM+CAtyHPSffFoM2aV
2bzksEdjBhGW94UdQ5nHWc0vsEm1i8CkejxsZxliMR84GokTKxpYYZqj5I6N/0pN
yXe9yVqBT4/hKW6Y/IBZDp3ZyW1tsVffl7YiMUCnL8b3C2grJQnOkw8b4zoY+58c
htxuMixIKFtlebM75ARMCy95iyo0rdzfns0MutedIDwD6wjqMCD2cQPObil/WjXV
cExgpEScQmP5gs5gH834WyZ7n1o+dwn2lsgasUi9p+ccP44sJy9oRv9AiV8kf5Yc
kLb681pjUmakcFmx1dT2sQe/VnAne2ZrNWGSNy9Y8fnCRdq2KH8YfCeq9VgojxKP
IOCZBO7izTQTeTR3BMPfLyd1Gy8/gKYNOCVkWrvMXjYLKUY2yXSa/1pXRcxxdJAh
25JK3mCrCnOFdlpnGm8UFFlx4f4nU2UTNZwlfOvPDjWThqVv9LyzcuB7iK+w0juY
+7PNI8BTVyc3jeHrumjsuiVf6P3dCFSCHLuiezaFbA+RefykYC53h9tcwn2bJtvO
mIBhp0tyBIqa7adqqND+4/+siTAkg1pDK+ZMIzZY5EwKAuCj+eeDlyo3fOErm8NC
1Tn1F4+UtiqWWLO0uOKxsCWYpMzOhg4mgInQijPMvCPAaM4OV7Wu/cRhk8d8nCl6
6IEZZw0QbLgPxYgU3xH6ulBlNAIrBDbgAlb0bhIy/gcQ/ScOa1YH9QEdRZpx1133
bY8h770dT8+9TCn7/+zThOHnAUWLJGOeHkfq7gMrZ+TUCx0rHzJHlmuu9VudMUbI
9G7wVsUZDdtIpSSp0jVIVOPdohSYLODuUnM9kOLH3hqkRs4S6qn1KtqZYsqcSDSD
/z9+H211X2DS9/vG2Mo49Evos0kb9ioh+vM731WgMb6PD1XnFKlp2PV1Qj68u3XF
C4Hfyx54fm4mH7lXEV8XpQ==
`protect END_PROTECTED
