`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzpEOIviEyO9+k66zLAxRpp9+1WvnqxzZN4YBU0JZJN21eBkLqXEqTTL3ekBR4jZ
Vn3zi6kSjYtK2B/zXGwXjDfbS77n/R6pxr0cI5B7hcxfvMmi/7xz/HE3/cljS3kW
jB3i4lej9HYHc3hQBzc07GVwYUSj3W/pwc1COINQmDJe1WnOx7DPz8kbKHytfUyA
otEwJaJx0QjWjitpKOjK6LFk7xTFqC6vnDL2uYXRl02iHqHCy0y1oHLSnQw+UKD0
9FNX3MxVYyHA3fajycKaOOH8a3b0mCq55AnPaaw6X3mRS4/fRXeTf0t5KXdf19bA
wCIHzLM6kI2kPQQJZFRcveN+IlTQhe8iRNCYUvndzAobE5+OSpZ0rjsBRG1u2tyZ
Auui4jQb2A9HBf0RxHvshfhTIRPaqX8lWqdVgeYir6OQuQydzLXm0YGzKZ0F5ye4
wccs89xxHZyhA/CxvKem3FuLpe5dGswM53Ddku8ZwaoWbKIgQKH4R2RGLYEcF4Wj
hElTEe3x4qFwPOpE2ZogpHLhQXsLSsWd+WlXi0l7SgVIrJgSpNugc8KQVWDNZXvM
k65XKdWD3cId4vpHNpH7IzQPFTgvKeLN5YtyRyUc0cbT6FfcNcuZEHGGwuF6wkyX
K9OPgYwnX8GewfX1cPqheDnNs3yyqw0fauQlrfwMDtBK8fFjEK63ljlgh0AevOzz
nJ5RyT69BY2epYfU98j4BclCqOGEhlf1ZTCCQoPqJQp6kNe5qqnLPTpalKgguQBK
DWtdoqOXVzG1Xb8YAtBIUduwLIUf6GVopXyN57QCe7ePiLvEuga9Y5ns3JFj1z2e
bZ4BPXlgu08YZhCj6+OVk6rdzO9WzRPmjk3gfEO2XuJVzuerkO4MheeSvhsKaybv
1OmsoUTW3ejj9FrR1SS5G40pmsqI4pYm86p1qbRdmeRFtO/nlhsjtHDya+0HZ9Q3
rE696jrW7+bEV9g4nWZStZtyqnnZyuHIVTalzwItulLDtFwIs5T7JLu/HocJSgox
iwhFczRUlvM+V71QPmw6gV7vqFDzUF9HHIbt+d7VJCXcEQHh+IVq0KHYQKGZITP/
Vl6JSbDETM3I04UDiIUMJE8crNjDbHCFt9jVz1SI/pFSplNpU+kmKWGSLfkt2cTu
xKp5pMcl3AeKJ2e6UEtBiubFp/H3FylFW2P+DufZATRkhrQ/JW8an9baXvh5PoMh
DltTwz60UrdWSvGRpq27xySl1Z3rrSAMP4DNLchOdTexJ4wbYN8SOU1w3FBya3ab
77jJPJXCCNC6oVLEbgsjiZuagYy6QbxxnMbPTcNY0tlv9nmmOBEeuTOvkUZMhGw3
wuQcAZw06JZx80x9chYYWL9kWUdra2NXpxIZuPBmiQ6if0k9HpyvMpTVT8COkHem
HODvCKIOhTIW3HCGd75wHd4unXl16ZfmhoFqgRERk/Wj+iBmydjvrNWMgR1NT46w
M1VydgOigMLjlNAEiYW1yVBV4h/q6S5G/QIZkmozDVGU4WLNJ7ebHsL4bsUynKiU
erTKf/ZxVMjPjwQ2ZO6ZcnphSQImsElChFwdl/Ro8tRTUy0Wcp2FzbOExkoa8wyz
ZXlz9Qps2z6oo7NDum9Fk6nBOvBerDXOnJ+t17ukjfO24DiwW9yhKG+6Uu8/NAVJ
Benl5zhSg6l6MS7wek/u8q9Cy83Dils7R+EpfGyMjiidCyzVI+1MjL6fpSwOQ18c
wnCWc9vQrn/gy07348YSO8qdiJUvYXQDPQZptg3aX7MPJuXUsRqBoos5LdOa22QG
xmnY4NY8Luc9BZEO/4vxGyZpZkxo3VL9qicpQnfRSgklEQtRWyobvXtwV51GP+0v
Hp7uTCE/SM9FSxk4bo7fX1hN2YfyTu0U61YafLaGTzsnBGw5xZJTR9b1ah/St4ps
hdJiKGxPUDeID8yZMK8gu+Rs9DSPcWnlvlW4Zw0vzvr2539Gjmm5W0/CU6gpDpb3
vRCzsHLGEHlbklCZd6OCTnlK9BmuDeh5T4kG6byZUxzexQvg9yHjvZVMuDtO/HLc
8d1LkZvcuLY5apeH9ZjQQl8RjTqcdH4z54kVp2wDRW2W0L10EW3Hh+5W4pcfvNSU
EF7kdkiI7tpRyCr9+POp+WKOjREFXTN5tBsPa+x5Q3odYzSxfqqDwQ2JGkDuyVHz
g6TvawIduRIhaULZdBo+NydwYBPo8f4cwtfSGYCWRpXl/q+zEmV/6ULYkTkIvQdB
qjZ3WvUMa4WKjt2G2O2vR8iv+pslzqRHgpn1Qo+dMfn8CicuzCW0I8ppPyVCtTyJ
GPHqvYRtOSEAbx02NL8rkq5vuIhHOv+zPczismEzVM6ueT478qUjr2D0kgFsX2C6
eVPheR8eDEOS08vs4m1VZYF6lljAgOREIxPPVc4WekUoD7RHkQx8fSFwd8y89Z0l
IxFNQIlvLx22ZQf464IQC6f+yetqdh1CNxGfdCmL/WJ4SBcD8U853XTYLNk32cxj
rIcHn8lRZC2crAWPTq8KZ+xmSo7LhyYNOy6YHWmjjYAlBCSxug3BgfuiF41uPJR2
EOv3Z2K1w2bqI2hmoxAP3ygsZHJqjQr1TwQqY2KfvV0V2bD+Kl60PaAvw2AKVF0w
4Pk0j6O3vGi38n1uNjiAUJG23OeMo9xC2ap2aNViilHX7vtmn/5F3yA1IcVuQP9v
whP2pveGeLfjVv79pSyZK1Qxfhkof0G9NByMMDe1OuKOeakJvdrTM6eMgGUKOHRv
Ao9kgqY/Xthvbljsy7OY56xG+Xr5cJaJNxm9l+Sg7jJuLQl2ixkPaOEC0/E2gqLi
wUPosCJZ27VYvvLSnh0nNrq8Lke4eDMyncliEr1yJIZhMtDu60BHRAGLq9wxwq55
wa0kAhMtLDqk7WP4PFl108aAQe74ApER1aS6MF276aW60ZmOf30ZWgl4gQQ6cpg1
T9NQcHy6egHl9nvDQaXOeixA1wrLgBO3MgBELgo0UAburkQsnz9/ZLg/as5uVod9
ZFpG1NXVikCLcO04JMNfM/MSBVQzKtHfethvWT3rgYKaCh/gBN8s9LtmenOqnHiL
aoJnhx3naVtbtk+3AXUCzELi1flMc4yVYNpBydtSXke/tet2lVog+KnCiuvpXB6E
8aP91ns4Cx7EXnPi2lzXpqUdPfomkVTzhaSlnMlHgh27Un8om9pSuT8scDdYX0//
ixDL1dF5lpkParbzZDbgZwn9m5Ozz0wZIIUZHO97PJMzC/2ZABB/+sP3uVbybC/a
P119WOVoAmnLeNDaiiDaZZuIdkuxn3ke5co3vQdUMTb7ddzULOQGKvvEWqWma5aW
3umnTeo9/9KfDAqnUKtIRq7B4XXizVFcgOEcN62jVm7UKIB0vGqhMBi4tnw9Y25L
LHl0Ha9b/QOUHOgkQlZ/Y9bVBdS8AfwqlJ3ufHtd3UHD5T8Jt7/fKeFFZEAmb1Tr
TLrWdJkrxjTjkN6ZevNbBXVUc7rcaQbqq82nFiJIFH7NiCRxoFDlIHY4Y6dWU13u
4roH4EWrRSDWZjqoNOmJWi+uzzrEYcSlXuaQ0Faik5fxrlnnUVH0tbt5kPLY2zgR
HWJZpsKMWuaZ2Y7wSelskvrUee9PVegMWekKMtKKa9KtuaDg8q5/iBAq0PnmXokX
znFSAgKfg3YnqUWgGqQlLEJEXNneSMI4D26/f81UJNBlNUNI72g3oYyE9+YNoy0s
KPtUgI3d0EKcw83Abfy0J3wZPwarGJv43Tc6gh+MZJm0PmhjlSqDoYXMq4MeTLkO
Ju+i+DziGw/0I7Bbq0cb9YqoWzDiPWF62uw3KTVYbe/Rowhqf1Q/kD9HL5U/nMPe
TViiJQ/5mTQuti0sCNL6Ww==
`protect END_PROTECTED
