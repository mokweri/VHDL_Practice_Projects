`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Auvjj6wey+otjAk5wWqOYDR9tnvdbBbsAfSOuhy7xIdGYM1MjQUwX6Glhqz/lKli
Ybi2cr4+xpgb+RqVB6TI1fG9YfdCdSyimpDPgq9qBaIUec1151hSVOBZZh2yc0Ql
8t2KPLG/x4btzXl6kWmdsCseEgC5AWXHR/Gpyd8j3cPqSs89smzXma/fHo7N0OfT
txf5U07coy0OULbFswcRD0XYSBZIw7wfVsvBLN65BuIaVMzQtJ3lDxSanPjX8uDG
QU6L8kfvXuQnf3IH6IyxNVz/0dvZP112tGvyTCBfLbW30y5jRZ/+zMg9ZJF6A07W
8otiRBd11pAD/v1c62IF6m88nfnbRGoIMYtCbdf0J7Rke85K6WsqDwivgHUAIiQZ
UD9bCGhVX40ZNkV6wEo/vCdPyi9CPdXnKWGRTlQ7fK7vW3az+veMJ9YGz/6ahnWe
7tAMsyJlvA7q9LwZLzjHGWJd+lEd+tzqpRBwLd5jsTuK+zZflr5UjBcgBsA8fQIN
MBwGhVQPWSqrGd8iYD85RCnt/zgq9q1cjoFTYIaN1xQnst867JJ0k41MqT1o/3zc
Vd/y+YfYc/zpOH9DlJtUYMSbmTIJ+agZ8byFrRtimA2rckSeM216LdUpjOAWy8yJ
i+a8RnIMkBb25L9sSycCzE6438WAgGMa+pGzGeSKbobXzrEVqA9mRLZGR0soaCmG
DP0I+qdL7fl+4p5dPhUkFRdhfFP8jG4lRAZ4iRE5kCWQRuWuHekWq2gtNRoqGfvz
EhL65IYLMg+nvuZ5yLMh+dA2Q4FCe0/66pRckp4Q+ZlETkfvHliSf5t0evrH4pXu
HB+VAsdt/X5rtYBifnRheQcvJfiHm/E8qDPD1v9fnEAJTeYF1UK+esVGw/lJs7fq
ya9vmbSbaxrI7VbqYlnY7SzM+DEEC7I+/Sj68IUolopw5j9em1paq8XCe+5t6R5E
VKwjidSwi7pVYysrAQwQTVri3Af3UDpdBih/1Rmm64xMdM1Q8Oug4+xjFwx6U8HA
K0dt/nmK2e2EXK3SFFPaoLWDAWHTMGR4X94p7zjj/CBidSvjJQ1xCUd/hp0HDqM+
mAckQ3ZOvB08bxti7fx7sn8ZJ4QuFxgrtbDvVOEx+0xiRb7ro9I0gGf48OwLpaPJ
W3ywYqFj20gNLBnyEnG2+hEqY1GPuokWw4XAxO4vKqaVJzQaOszNAQ19N21t4WLq
NXl8ucrBnAtP1fXIbIFcrxGHlpwn2Jqz2n9nvqNeyq5lZBi1J0IIb1GbYKR+S0oN
2+4OitKUUYOsZK8JHwKyciVq6GD8HhzBePcuieslmsVFqcI+RIS46JSd1YBO453s
/jyPzrIN1HElsAoZbOVH5kXk9El64uoRGNX5bHndVuy1g9tzbzziFmrDLC74g5fP
2/S/vvXb+7JYDVDeCmI+akinGLXxcHA80lcBZvapmCpGYqYoFbkaeEy/lYyyTK3D
QoCQiy1JDOX1uT1HCyEObWlLvOzwHjCUpPVYjmiT7Gu4SfUCAzclqpIut/jaNW+R
uVKD1xK6SULiPXQDNa4EpAYZLRjYd53AHpi9SALbw1Bz9jsELMLKyIiGb0xBv8kK
oJUIhNeiLG7ubNJ3FmctNnVdlz2AmwTq98jDbUWskah3Xcvw4I7l76fVrog/snRD
tusjmTUNH9JoOls7FRuuMsX2HswA/Md99axhZk5zlxM8qSFFXzOzAEZHHD6NuItA
AwpbBg09xuDfghsAeOa37phod7eDbPY2Ke4tJoubnIfRwFR3A9TQojUuEQwZ/tGv
jPed8Y7mIVmqntLX6S/UwL/agemsoKseJaqbBYd+Urg6NET6FwwC/PtKe/YxsqiF
DEmw8fSNGTFEEzRy1qpq20kFVyMZgHfS1bsZ8N975jnSPhsps41hz8thUdmMicZo
7z+YUgLliT1MIq38G7UgiZ1rozLiJ08WRFnF4s8UWWpwsCZ0YrpyZZqNrM5m7n8F
6oGhOce9BVOZvvKJQpej/zsGkhD+paopT75cNutYl090L+LuZfEad6QjtdaTHsT6
vaghiAqpcJc9bRGriVlaWVzY1VWTfI8cgR2XshUZMUKO0MrGaw/LJiGt8WBCWxix
c0bw4UHT8QocvLy6JM72mUfNNvbrJ2GLLCI0r8p55qbDRdWnZO0TrpcT3R0d72Jp
1rLPM5YEMt1igjnUo4SX9YSRZP73tnRlInBjQ1xUSGolT6mhKxlKYLfPNuvhrs+5
69QdFlgAbXJ4WbEz1Y9epd08wUSpUIINwmTG1UiwtqMcuLDo3IxoAcII3Pf6RgAt
NaWozfMNSPRc01bi3H6y2Pz/SwXY8GCRh/CME1HQeoGWqO0yUr6BuH+xCUWcYupW
rYRjKY6bx68Cngudq06QrvU9AeqhCJ4dlghcqgbdllCzHZPwkewXGm5ACK3QfbiP
Bz1usBgr+KyVBIkw/5wmXDq5VdWLZ8bIgGX3xi6TUv8/cke5nKGPCoISSPLl7Zp7
HuhE492SgGaxcxhSxM4I2qpX7ecmS0/tHpWA3T/KaH/67wTvqamH1Awl0ML+kibd
AVvvNhgrhmD8G6tEsGicNo2ZH4KlnZEfyxIvKBTdc7AL4hEbCRkDobd2GR0DxvmD
m15G5h1IogBBTUFQ7tG/edr6kcpSsdLJGeLslQoQoPsc5R4Z1AY/0xkt+a/we60r
juLDjLokk/+JECPI9oBKHFs3K2NxlxHWDwiHrO/5dB9EtEHp3wbyvLfUYEtkxLDC
Iw4YWANzwb6Zs+QHA2HCq6/xyBGNC+GHQ2MLA+HecT8+zUukenLqkhGRvYJSbO3m
b/kYrgCBXtz+D0tyrWcg4iJ8CfE9edaHNo/Mu72SzRJGAv4QWjTWU2ccTfOH2xmo
gAam39vWAlcFrtAcmo7Fynj8wDj8rZtn8nAycyUbexRyfSJbZ1LZ3uW/Sp2n26DF
wZy1J2e+Z4LvGlqlsnCs+QkZIkV7jQI/dZJ/FiXgKSd8asTCTlddlgjXPEv9WxcG
mwIVa/t/0ec9Q3TzF0ek0o3AizfUOE34ooXgZc/orWJgQ/g6t/+kGHcmagcPFTiq
UuwUaLlnUsQRZguk23za37PfgDSjsrNXD7k4Sms4wf9EgsNMrdW+JY1r4I+AfwNV
h/HbAagc6PjEY9DR8xUAuwfofkJ/cidV+tsB/MtdlW8ZSLBEs4FxUoop3Ku/GwcS
zG09WdSl6U22pa9rQL3JSMn36r9qU0nbn+ovDTGDP5R/w96XaJWte+/r+vshF+jw
FPRSxRF8D8kTvAWqusuP6ustrxoswZuAv3sB7G2WCdkmQ3teTRgncJEvb7RPEGY+
dh4Tco3/+0L7OjiP8Ys5SbSwTxYeHEeXC+6tuy5IP6CQRryDHY6k1KfuAHtlZZ7z
LLbC1VPHwE/5aBiy1f+gPhBantgqR6uRAfYWB/Hleaj5oFPukSg2STliLS+p91ld
6h35yRWXuowvswDuGlG95+VSbonSGTV2BxBiO/u+u/EQ7C40YS8O8JlRlmFWYYLM
chOkHB59tjPiVyDmbLR/neo+Qnap8+tVuv1pPniT+bW6vG140te9t3LwP9aPSpw9
HzXTI6Nhk+IktKEtPTHoo3/mfKLTR5KbM2rHl8UVfyZEKhmAd3WOEVP9JXIpG/ue
dx5lql6UhxSaANhb+MiEeijUdYFpy3Xxalr50oGd6gE/z5RhXa6mfHxAPESt4LO5
BjhYVrZGScZQ3FrEU05aYIFCkOlVq5I4wfjsF/U5rlG/zuyQ01kngwh0M0CzT8YT
l+WDAnyweJDN17c6KakuHOypophdcbmtB3wTDL3d9ifQykH5c0zme4UWS71zjGHI
+QFVXMIypqoMSVkfIwDCY5puEnOdJ1KeFa5xtiIcHXTdDArWot6woHIB09lTkogH
FW8Sj5wq7pRhcj+7+DnKpv/KAV4ePBvdf013gAaVtCpxywc4R6CAS0lvdloe97CA
zGPQTwfMDi4F2AX1tWgaeougOaG60rGPawbIkDCUs4dtVZ/sh9kkKC1IdxZnfW+H
yAUEAsUg4aE4L0/vzmHZ/zmRqZbFzyHxGud+awaEB/GLDwk/sxu1x8ERDyLRF0lZ
+zkL962yYTByBDaOzQ1H3K4qiCr5oDK3mFOc/eVsJQV8dF+xwbI9+uItj5HtM1Xa
JoGZWqhylLjCBEe0y0wk/i/seaEuBtsNNNaItNGz4UXybhiC1bi8G1OD5pEoHaQi
Z4cdpE9qY9Ix124SyhD1Mpa2s7afeA9uO4oY7QcJjSpmjmjJY/PaaIXsYH6MYIrN
zh9vcCz3c9h+aeGYCfuOXyxtLV6w6VTFngT1INAM9nPS2SdHhfvNDIAE4lXCjlMA
+cFo3QjU70Ki3+0g9NnZRh/pUBcWgYZFncBM8WBbQlEUYF2SmCup8i3l1MU7eZRI
G043qWtZRO1DVus1HYbAmeOPCsjJ+z69iQqH2jOVobRW47QKNujTZ6+N3NP6sfML
9+LE3Drud5bPiOjItN4jyTNkLNQ3PscmkYpN4b6q4IDxDCYmMP66alFRKnZfovrF
BKkpDLJDdblyFy3oZ0B7Ad530o2/ZuSq2r2Tu2nT5uGPBJhlqdGJPd4F5isLks4a
JwmHUtO2NonIes2vYEimxCmD42Fuxrd8mtKIf4sSNm/1k7sBqNA3IMQZuzxOQoza
oOtcmiH3xLc4JUU152LO4ijxebD+IdYxfvtK5tiHZd41oW+rBFHaWltD6kefhjk4
JMYmaGraKE4PLnMGCSWVMUhRGK5ZTXffE2SFGHgHrYjJe+Nc3kItD8mtw3hpNEw1
vUAjRGzjmb5+YMd0f5oYqXtQpCbNCmk3OqaqJmtDzXn2FshkAyTW7gbQ+S1nPutx
siUgxMIqaurhJZNppSPnTaU0YBVxhkPmjvZ/CzDRBOn7cFuiaPEEmsS86hmsICdo
RXepCP28ETr397CXEF1bL8hzDbI3vqOl1gPrVaJ7lUzgYKgjIl9C8+jsqPk1Mvk5
4wXgHYKRL/WbB7QVqrQMn0g1F4zzJzFdm0F/amElBVDpLWYMq3j/zSpM6xazwfSb
E7rX0UvdVivEpo0HjnLu1MVEqJmONiXG+eNQ4z462RSGJgyrynZn7MFPKltZYzQd
Jh1yqqxgcvCT+ZXm64yxe904ck7TV/QqZI6Bq7FB/RiDEDVDkPl7XEYbQjd+ZT4P
Cysb01yaMINWc4OeXHCIlKafMNNoNvWkeTEo4Pc0B4boSiKDCPwhlf9FcBY57Dkl
pmVUVMrK3Vmb0fKbQmY9n2YpzMpXKodpv4oq2zcsdOoaRj8ZExXWGkihw9dSLA48
MzArohogr9NWdoypBHJvJWH99dxaX/iYzsfvclmp6epAP+BGn/ZE0sn16SfzA64n
G9ceejbnCqco68NCt9pU53TOYDnNmN4Qd1RVhMy/D7k4TIWxPkXCyVg1zGzhvSkY
j4GX8oUwDpfEEkADCCoSQQKxRlscYERZ6j/N3RrKFLoCNfSuLOA7/AzRuOj8nOHv
YLBpG5AaWJvj/llxt1iklZRdbArly6zozPgDKxioT3+Irn83EvaSuz1tGQNkLBKL
VPKSiASqFvNxT7k/J9r+33RVrrNhfN+j4VnlOvVu7pTIPqZIh9dK10pPG6de3i5r
WS72l0/yZU7R9kJFBJEzY68POu0lDxELzrd7mOXD6uWWNQD4ifKCJESINJzaRHc+
KKd7zPQfvCI/TB/cQVPOLrxbcOHkintOViFdgKpkQmdc5Wwr3b7Ta02JgOSrmRSb
N/jtN+FIUQSeQlexkKr/6obYtLR1quCJInNtELUzb+saq/I9sbddvHkNtdXVdcwc
hpWXDEP+KIrEKmoSASR5IXO57pq1CGG7XXQuG9GE3Ym7rWoURMcmysNY6MtykHwh
J0v18t7XjB5qnQXHLre6obMSt60aJPTfECJbNJSC/mPjMNcp9MFqurrvoTdlyimd
gWeRu8y0GFNFnoY57k2XwAvaSILW2bfu3YOikYXqPOHr4iqhD6G0kxm5Quv8Jxqi
1O0eqkls0y5cRK/bJySDWdaAhlJiYwFIPNsc689c0uueZ3Auvl02G9a/TArYBUwJ
4/QXMTGdxbZNTsZhSIOdSWXbMJPbHv4fqgnq+bZc6oDnbuINaUQczAZ20CkGGS+3
/8UrDEr1J1g2TKVMjwohcQxGb8HMXfWNmFcqyL6gHCmMMGSW/2zw4EiD482YZ7vl
c1R/edK930chxI5Ek2CxBie0iULTAAOlNz3eRtQLs8v8mmT1ytk0RhYPSAbHg0Zm
nBGYGCa0ToKPKkM61xe6TJHWjPmorwEJopcDo6EFfIkwQEOFLfIUYHH2Jzmj8ZAz
yTAi1I18CXj+64lM6QVLDpbptXfBUJesAFjhQqutH0g52nXpWvkF/y9cz2H42WTB
2dFXbRQhGW145FgPFXng/mdbGD3DHHZGXibLQ160D4+RrrfQZSxM05ZOpjXpYC0r
MfPY75XLegxqyONCulFDzkmki9kby0n5HuzRwDBhA6BN8LR7lCtENxv+QdDbKQDg
dAUlqwu2ENZQRAA4akqIzBIk6vcp+dEcVd/QR63LsVOKtBRgFrOHKgSQNO7CF1+I
akD2hE53ri/JIgH/CXMr27CIpRIDw0FVt4itf75PrW4t8jaVsUbhzMdeBAIdxWZA
`protect END_PROTECTED
