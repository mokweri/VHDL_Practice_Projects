`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sTMDV4XHvuMc5kXwHPPzRsmhMNPIxxZQ0BVl6ELZZh7q4vYtfEewVuM6OHKhzxgv
rjrk8uLcc98ucioCCTmIvMXst29ThNSNGjWUhEz3915tOQtuUpY6an0fRacp79Gc
HuMNHwtfIi3LaczuGpWMag9KFv7mr896f1jH4MYGJbcyN0ISRjtK3RDFOSKaTLBC
DanDT8HZJW/x52ITeX65e2x94R6YwJk//5T2QaOV2p9mv8E92dnwkPolsaWV4fvy
4T9pEDJTF7OnBjcVZiby4zAQio0s8RG68DP8uF+Y5vx/wlngLjCdUFE4nloRa25R
4Lh//iFBbF8mFgh6hrQQaAnMFK+nI+EgV596CInx+deGveP5sx8vrBjWd/6Uhka+
/Q0M2RTt0XngPc6FFLs6WivAsr9AZTogZgT/fhOXagDdssmWUpddrqeIfHRygicN
N0lDFtmUUKQytMHBG/0UkfS1SPJOo0wfANDcp8HCcH8fF3RN7KtNZFPmcMsqogt1
rpVlYipU5GpTECKZbf62n0x6FIpi4lJOLfr3BxsHagleuHJOn0LRWONYR/WgcQn4
ol6r0X6NVgUdd+7C8S9QfVhjC5WDkH9N9zXwaIeWrFDc/yPGcGs8De3NM6tWuiO5
kyLFK2wZQAtHdp9Ud+G184nD/QZm7NR543vfrZA4OqDAQ1tUZa6a6rB/F447vyaW
1Fh7OgIEgM3l6cIxs4eZg3S8NH3KPVKfqVVsnQtKZ2nYU7+Z2NTVayoKIulkJhG9
+CKT3YOg7WQnwUaYk+0Nf82A7LoPVarQsHIFr6OOqTXrIpf/X2lKRotKu0xURDXo
IsSCA0HdTTctpShThCY5/51T9ljjqmtyUhpBjskj5Yhoeoj+nWHXhqwlI/q6sXzp
xSazBUyGO43pFQgIVrCmxxx7DJbO69rqFwGm97YesYh4STJJ9dccaRyV/nw4fh8o
Ba0xHlsNf5HeUvZZmJEEs/M/pNUjLQZHNQva4sdEqDa9xn/8RIG6WyOfiT2c6ce3
LgNTyeclvaGmWqP+jZRRVjNRLWLZdb5l2cvm9FXngqYiQFacJg5dITtwx/yHNtzC
GJbX0WcXVZhtbiO8nbQy14OfinRQPkyzkr3FcZQwJCmSV4w+R0KH8A7iFLoIy9aw
ir6j27/78iXSvHfKvWwCyXnTfWbmLeoCgfgUIEAxKkHUNFqu16cdiepL4YACxJe7
22giA6t+FSRP8ekSHzvwffBNsXTyKK7ke4hIaJlsug0dVp6s1dr1Clh8rw1h/Ee5
oGdGNYJ+efLouh4a9eVbmYUMhE0rNECRAqX9+LNyas6BHxruN/NyrcBGclrB8stl
WJUqw+S71R8lw5SOW8tAshmIVfR9gpC5wgHKePPFauvrKqOohhv1fXF3jBSthKDY
Ziai89fbVHVoCpSn0MQqt9axxVCcGmQIafYmMznP5Lpk8KhyDSuoU/RFHVkSC8ct
`protect END_PROTECTED
