`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlZHubNQKYEG+CnTW6+5lgUry9KawO1yVSCeyXihA03N2qcq6/dRfRZezppB44RW
JRqoTrk3agv4BxRqAeb7ak/n3zrMJn3CxBpTaIE5hrCaCgq/z040JJQxhH52wT1D
LBZlsUwtg4SgvSJppfeGiZ8epys+j7hCdPo+hmX7HFQA6pwuQTvQfJbFWxTCFlwC
KnQ35ylKVH/DhW8bkoG03sJdUpJhrB610IpADw5gWjdqXXe88fLJyT5BTslk8IY4
DntymJXcejwAvYglJ64pwbak41VreNphKnCoRoP++Jw3+uHSFiS2V8s1W+qsTKNq
5tvwN4xaq3SUuELgtvvTEm9qNH9o7HcapqL2CefGbfmcSIRUC/hE/Q/begAnWW/G
gvFrCBuw8+9DnVGxUn2Ufnsvg+HjU0iJMGOarn8+BNaaxhlwB3L6aH4uIuKKhR1V
ntI9S0x2HrH39v7oXkWcVPNs1kvTKibIH1+DCNwYpmEFsbKmfswAaFM42nARd8TH
ZMVnciNQ5asIJEnbZjbP7MKy5OOZ/4X7FMN+Oa3s92+S7K/rpvASifwq1nccxOj6
EfBXV4vvuXp5kImLcyfPrhhY17udX+RCbqIVXlqFZwavZp78ENmEFRqtjkL201Ni
tg8ktOIQi5bmi8WOnCcTNTAZGY4EVBuQug5SsP5BuhxUYBtzmT7zfE1vPapjCd9R
ih1glzREMnTsB0T7CnbBlWhRCt9ZcHABsmNAn7mb6doN2hcaoF7WWpNK1Q9EANaF
wjYxdNGWb5zs2WRv7gQQ48bOcG3juLt8IBwiHncJbQIoCgc/yjCSFA/I+zi4cDht
ZH823SuvQusQV0d6dpb7X4gZgnDGn9szKGS7vMUAQ11td5BsCENytWLZKKLrtNes
0JPFCKKcec84Rh41BHFfVKfuf95ysEW1b21zgAZ2IM98eWMjjL1hqUqkYmziTB/G
hH2TkixyCYzEBfEOKNcZL6SyAnPutK7pBu3Enz4cDNRDxXiuNDzSia73m4AIGUKH
O5O31Hr4WQZYDjSV8AWb4JmQNjBXvrRGoFRa1+8R9RTdTiKc5snohBxSwFh3mttK
Bb6D/oGcm7RJjvFo3yE9J4O6XVHfHFAYABLak8andL75LcdpXzma4iTAEHQAPpXg
08iqD4IPLzaJ2b8i5lnIxt+NVLFhugj6d7d4PrKE4o/0Qgr3i+CdaVAdUOOntJsp
jmV3OWZMA9ebdzsPK+me1xSHbYXKDGuil8oXphONcBiXYlKjjktbBh0cqM/24Reu
f8q2ItknVOYGq4UWTHqc94BIFnYaGrEqoUZwLkVmFxzwwhXgqr2A1WGSfPMZyxVp
SK803B2501XL3X3oXZeHfKc8SPcJWXJJK3UmZaKV9ZEjwrd1tpQkueXfDg0F3vMk
QY3I2xrXkOcRDvVpbVFdSLozw9Bi23mDI7vreaVkqleCpOKfHC9wJTu2xD7EmnYR
gAReXkZoiz/0EEhoaJYoJGcPy3PwWoc6ut5qhkBP1Qpp/Hu7Hy/rOb48BACNm/5V
glvKVFeuhc65y9hmDPe1eXCe+I7RuxyW4Q6mjIlQXKz8Ma1DYVzagER1zqTg2lzb
cc2XnUzYsKag9IL5c8ynoZszG3iXh9ze3nX58v5N3Mpbb5p7KBG/K8Vj6KM+JxtE
D2F2VMlq5zJOPCYlczTMAo2ZWeqCHRweo6WJBMNWv3vbrau7gCVTj4CPZKkPPjL8
oaCYEQFHlnGUcwqPTmU+R7Spgm3BScv0zFy2ljZfSwODetSW2kqeHwyrKVPpDM6g
6HL0wLi/zo3lVHIUaZqq37foH+uZ6MqQ2Ts8slsaKoJiUQ70mzGHCLxSc0PKhltQ
S55fRf8DjiR3GEYMVQ+OWTKFoSoFQBZ80/jHEsw786zlkrLbxq0KS8CvJl8p8Rqy
F3u5eoEKpz+Y+5L91GepL9qC8UV3/y68vzaV1GowXj4dscM2kJJqSCFYQ6ycqoky
kGkeo42zeW6Ja6PBlMtVzzqiqKpUi/R7uTu37/XLKXN7y7UD6D9GhUXmYYhLpogI
tH0nS55oNYo4C7PBbWChqdoj7d25ZqHLnpg50GLXreF7FPaZ4IFp3ThtgANpYAiq
b5VCRszaU/18nhpVBYH9h+7XGlf3G+M2SHRNtYAnabW7K/z0q8jeDY/HXHljRZiO
V3vlUI3bAHF+63Vbv7ArE7KuXxybXzaruc57x7pYev7O062AdO+iCa1/SUPSXg4A
y4H1+cNfyDRYzMPxtAcHuQtcIhfL3boUDuDqFVmUWbiMb5Iwic9ts/TPzUJfMwNQ
9rX8hT7k8ANnNV0zRqGzge5qGX9VT81ovwSMU8VNhTvn1/6Db+kBw+CE4mMXN0oB
mYXzh5Ll9rqHTgi54wwGqyEkoLbZEcc/MPiYhuPP2/7vlg1Ew3cXcnjJMQYd9EgI
WR1eF6SqqWuwKCDcKjKORGvnqQp9Rk2S+1ETb6FZkTLwaqX2a20bfyfCMGSr7bGy
18VT4tI94LuwBO1HPpMecQC7lhTr2hwpW8gEpXhpP3kGu1LphWGynWunUpn/9kiA
Zp/GN1rEyWuAaY5U2e59sv8po0LULBE0IUyarUQV0an6esuZLmau3YZoSSWjh6lN
tZzjcg2nzOsF9rtfavTzgpk4hDftPeDw2FtVJeqY3DoGXIZ7hKJFG8bmyhUptOJc
pL1OsVDcpOFnESX4n6AWRLwr6m3ZJb8IMY7t/xHNQby3lQ2LLq7tbsFH4KP7YB+R
EU2bhJccOq7dVtWMwkjW4yFNsPNkdLvd2FmJvf+/hQebvONg4MPpF7ixJ0q+B4bz
F0+neYjblh9Vn232aCbh8Uwgr40bzFVAhDv5enZL1rafv0pKL1jlC0d0mt8n0Ks0
`protect END_PROTECTED
