`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2nQAYRpLfRN5RKmlJxn0OyoWHRZI4M2WazLPKB3VUVwsLfWtytmOcBuVQIHxGojX
JLTmSYJnACdW5iBK3Ge7AZ+9Wm6iSAWztrNxJJQCGeq/o371IM3SerHeA3TWFIdt
+gbBD9W+0mxgfSWvaPk7FSMe5WSgI1VuLQP1jn0lmY2soSRNjuh3TrsENMsD0lmc
YceGiDse2TUaI+lv+pTkGZb+1t7Vfz/j6QKTD/IhnjyuMbCiO+5NgAyRZrsqWOFq
evt3F2h6BTH7fisBmLCeqNlkvFU8C8xdCPM9x+E2Mo1wC0KGAQ4xSDnlFq2HoLm2
Qa/hI8FwXmK1M0bQBm95lYynbFW8RBG+eNpJompauIkX/cz2FIMKJCbnRbynM2bc
iwX6CLchxow9ZfT5eWhccA==
`protect END_PROTECTED
