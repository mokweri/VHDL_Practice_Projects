`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+swJ3QbdwdSzGNJdM3rqLmLGaWRdttZQsmjgiRe4GZDa4FUH3OJ/5n1eocpqKCb9
TKABrLOmFUMwdIuRMzraRaopR3eMcaXXBzqRAp3bqADDF06oj2IKiwkIKr5vjlYV
NYysSWknsK+AZv4iFFbjKCDvt4+HMfqQeKSPa4y2EnyVgjlzo/4J9d+JITzAJiXn
AUn8toCt9HSHnPX1yQOV9XwREyH4Ii8NsKuIjtZRu09HE4vdIUrfS0k4z23fpmG8
P7xR65Sf8cD4ILrN6eTn3Yu5iY3YxjPDrzLbUyOckjYkaP8VyZkPBP7PyWHM5c+F
Z9w0YXFovE7/A1f+qBzwMgkXfS6f3sqJKvKW1/dbvptdiCSS+X1a8YORBBUJzJ5P
OuWo0RAjIU6JlR8HGLYIk8u3ZrIbNmw+mIDJp1skfZUCyYS7qTaC+K/LY77FQNp4
pM6hjjUHbu8mpbtp16hk5nxbmcwSRGg9aQLuZSM6JXXrqRhStNLKyAap4gxoyGow
Vwj7cQWaSs1VCbHGUA3htwYI7bjaomkADnbeuYL/9q79HOxfwB7ul1NJPXfGQqZA
ytVAUBd78G1l3AmC2HNzWjOVGQUetO7bmbixhG7tLLAnHUgn6FFTtrZx/qI5eeSS
giHkeUDoGpdenb0DeL9/KZ7mlRe4XrG2KwxZZ0C1oY3j3N5Yl1UcV00PhhXgvAbT
knIX7mX34e64/YZ7JV8Bnh7/fxqS6IvcWBsEb4ZCuCa+2vzFU9xtVErZ3gHR40li
YrqOO4+w+Nei8FqqKj0h8BGoKvYTcK1LuFvsXNwuja80JU4kp//3bKsVFiBPj69v
nRZZ9/Z6evkbQI5WqfNXtJBLkJ0ht2bVgGeqXeDlOq7cDflULQj/T2WdnkQoYA8L
C12A3BaqB1Bw5+hZ0SbAe60kVI7Bn6mZkWNBcaQ1Jat874TbzP5o47ElmBG5i2oL
5E4kvlL5eYo70XYBLe+7499/usjo1//QUOn4mkZh1S+ij8LQNMFZMGddhs+f1C1F
rVVPH+stUxyZ+LB4qJx18t2GUZQVZnzdaYYinkn4I/FFcq4IFT0/vWIQ4IzZQIqw
dKaACg1LgqT5BSbTXW5KYRYTbCu6cOeIkCJaafWP5IX24EejJD+nmi42KCxqbA5E
xzz03QK6mKE1nUKXw9JjSnqVrz8D4ZhxBiaqkS9LRwGz/rKNNH6hvswzjewiYdIF
93Eox5ZBPBf/MYhvHF5TqJb+gIlLgK64CMbCrwG9p/N1TAKtainsR+XJ9k6rAYIs
s2pzsEVLvhGtdUHx2bRW7AdmNfHTOv9B4G5rifJ0Pnc/9LcASbOHxdi6yXwyKyCQ
lFioJ49/ePbPd2FTcTMrqprDB153BTnc4yIjN11uCHA0JEI1rfYSmH0XLpQmWA6w
QVtvo1TIv7iNEj1t0OXzDWX8r0TFceWBTYOCs0IdwTmIYZ7/lwNyODP59Ar+DtFv
FO4U8V9iucz3MvsFxMrY15rk5/ZRuCBp9tYaHHMKpil0MX2hTFE5S3fgGFT9S1yk
qu7n6RHhJzIhasfK65GdZSxdpTVoLEu7J1r0dmEyDe1u06tkk3dx2DI0QxEcrZxm
qOErtnyKhZ4msbt4j7c5u6c24c+wRewwZ2N0kSB0N72ztku28j0E4LLlLVcO2bV6
8/jry05eC6gg4ppfyYcwEAxJ0gEExW54UJKDWVsLWXahkU6u11+jhY5SrTKUzuA2
M5S4mw3MQWYq4hRp2CXDO3HFfSt7pfC+kTOp5XAAuzJqF9zD59/lW4zvnMdHm5Mt
jyF8rxsvL0az+ZcV1W4cZaVA4n2sZxUJbCs9gjVuiGSEPAGDupKx5HKm/q8Uomua
f7GxUTvrN5Qpg5SkmlNabOnkXN9oM5bTV49eE5ltyrOhrfVojuxxwxwYQztGxk4q
0eAGwoshhRkojjCdNNG/diUKPTcjUfwoRZvwgy8GlfifCOzT9eD8c0b4Xi3kOo8l
dNaaEXx+qMfwgLEdGnFl4PSq0WuoXTb4xuZIMYo3udinu71S6aZM0uy4iM+zp57d
uRyedCjHwysN5RQcUBa7/M//pbG/CtBv0MiXdUKe3JoUoL9Ql63f9WbF3LWByNiU
JIt7azlNw9dHYfKjVC+BV+COZtw8ZKbdhMK3PNeXSPm6VtUFcVgw9a8kuvt0xbo2
qExX81LEklhJJYnB3uUyMxXiLvPis6hH6BuuuPNwffXnH4MjJRepcZ+hRWDMtT+V
gKv/L44eq9LK2frx6qvyyDSaddwVpNfkx94orSllD3acZPQ7/ZnQielKqcexyhHB
d01PBglzhLSxvoNo6ANN9Ffl2lHEIeGBXy3eNmz9BAtlti5ioOITWabvvWNMTjda
Kq01/5XWEzljomFGpkU78fYChuMURbaXsw4tr/XRcnuIewE2zUc7F9IqZYse/vkb
flASQmgCYWeq0vbQZofnIf8VnfxfT0nBG+0VlilTIlD9cni+96jwN6m/sNCXNn8M
LmNighPTvkNKu/wGQc3gFE+nUC6r7IPWkkz5lRUiGK64qQZjwJDyh8L0IcQk6iAn
eWPFS0FoVhRqjj+ZqQug5EGeDqAomnHpxRjz9zKRCuWAfO8xWVUm9YWFF3/LsYpj
lZ2xpsas5EC3NWO4FbWT9/t1GJ3jJRlKaJiviszWzDTfWFyaB7gnGwJfexg9efoE
KiCv+Es9/cyT0lUZ38QHtRUJWDR8fiNLw86xHPiFoNHbWW6kqnkqXSM3RgqsBRm9
FvXVkv8NDJqRR4b1ZX7uH7Hl6My2eQa6NZ5Xi3fspdhFecSyyYuwxQn5qlba9wUk
v4i1xXzArINwpBksggUf0bAynhqqHQViCCYkyij73K3PiAy92x1VV7eMAHdI/I68
eOG24uFM+bPMekecHkSurfbfAs48U6zfENymMTgCPkYtpQqISreDY8CjOwRLPEib
Z9j6MqxLLMCqlVC2z5gatgtuY54hYEBKBlp4gUyVRnD39JB0vl2M/fd6CwBlPzHS
oX9/q5ZUD0RmLZkfDIjMFCaovQk2wQRNXFV0ewjmLbidLUhcGiqEzUTbOow+awwi
JjADfuabNJRY4OK/wLX2wnOzqm6+2mifZKE3eEVs9t7aBZ4UjuWIDvmDPNTkAJA8
tvEckRtM5NpEfoaa88dHG5tZ5my8C8vzrIS/OaDEo8YkiJk8BwC9X0WKyM46brwp
WDh4vrMPz0sqBhilqOVfMu1cjYKejaBj0rWuR+WoARTc1lltYENd8soPtJXzXj0e
5aPJeAsC3SY1wrhaknLh4GUwTR9Lv2Z90ySB3sqDX4yYVHiRgkpMRj3VeV5bZQkG
PrAIFRh/7qzhjdpo4yvzBo40gr5PeGUKrpo/6EaCmADHzlQZPS1k/qKIVB62MXXy
C7T+lrhRj9bLJDwd4iw3TB13da4Qm+PJItsVuQ7PaU6FOZ9p1X0hLKw7FCP9NNKy
oyN51ZHcZ4bN/OUkDYTV+2VS5Qf464T3o/jdHAs1dU2xRBE6sT/EwhAiDtwRfoPo
i1rEKo9BABs9YxOKRJpLDQmEIxJh7guMWB3YcvzjSFYdAsMNz/ddAVqIdyc/hnrz
4XKojq9yEFMVgorxCNAvGERdGcwc895up+TXPn4FJh/L1IdMT50zdQidcmHsMRqP
bTMWKv0We6yP1yr6yHv9gKkVAdFr5c/pYQe+uiFieBKIOxHlUgTd0lS9p0+gemp+
T9s//R7O76DHNGHB+0kFiyYmpgqKakh2sU2cs29ylxgYMJPDcsDSJDBO7U02iqWg
UZJWPgkKbr7y3KT65TBYKTRCyFchNcGdPMUsSsQzJlLjnkL3TSKEAqhYyNgWpPTL
wqP4h08hDA37P6tJ6XJoUg==
`protect END_PROTECTED
