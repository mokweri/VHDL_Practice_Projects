`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SUQs8qsPL9FNDYfInoGgSX3gD27yWAbMvCGrs65tx7IM1dMwGIAhkMe82ROY17Jr
qXq6eMQham/1ITvBBe7qPvU3CqzhUOi7yDABhploNZkHLnsfsELQK+736397rOSb
J03PyZRrAEzVywJvE+DXOV+7xkOQFLg6TIB5ebdVLbwH15hiBVsXwuGD7cuwTNS4
O6Ro5BxhP5shCB387yILvSbVUS4adaNdVbtL03b3tPkmwevezhBWY+OQu7R7R/N+
cZclXuhkkIl/FCoppCGBa3HAUbtbXhev/JVwGJQ1JU79qfHHtjrO9FjPbjROBlAL
8JXLKkCIzlw5ceKbHCGjnTn1ZNhVevkWtHxAae2CscIyjbP4fUO9xUxSjjqteZNU
ufL3z5EqGkhLwuo2D6j/IZQbZoRPa0BYyg/j9s2ePmbkDSLut2YLMMD4AJya5Tjc
5BJMcKc9jK1xVGe6WCKboAqWjqitPvq9Djw5ynjirTh3/LeD9+GAXvILPiiDE1NE
f9PxJ7wxZ+9Md0aRipUItf/q400tecRtktAam3cxspI1qjGUaZitrwfBHSp722Pd
VE8uMywI7ssAhnYlWaMpKplGT3Bf92y1LE/siTSi0oWg8ExQB7wR+E0JtK1xeKRJ
2rx7m/psHvy8Jw+lauttSaiQKNyTBfQS9JOgI9XtXnLTQBXhY3cY/iABlIq4j6JQ
nNh7UrQLWpu92NqD68VE7LGjroJaMytiVm4F1kR03gnTiuKTRdB2gePlu0ymRReE
yZRVlofYvtamqQWghw9ydP1HGuYYjan6nXg9Lgjp0R447T2WX3cXcq+H+h0P9Cxm
hKitVSDQFP0etnpSAkSsJpscJCyHDsvhmrmR0TjL1eOpI3cmY8DSblkfkVP42rcQ
p1/okDNyJUg109DKApWNTk9Vj+HXEAgHU2MsVS4acjp7KWX2MhzYW2GYI9gOOcsv
KfQm9iffOwwDpXl5r0AiM4KOLrP2POSBeTV0FO9w2S+Xsz4fqifGlL95YEAc1tNU
gsw/IKppVGJ7KiF8nG0O+jD4Db/XIqV5OAEbzA4y9uwR8WrBdbjdNqd87H/QrgWk
ikZtjM4TfqYk0ImNb8lgzGBfTCv4ks7Uc4j/ZcLD5vP8LBcwKfRH9PBBwOFTMBkR
8oKzgdXrUQ5HL3Oy8Up5Tzdo2RNmz5gWcLupbN/87J/fKXG/f2pbPjp1BSRIamO0
F560UVq4kREGuDgRltUBpBmgcxK70xXcy4RiUMAxdyp3pzFx33sislfhSP9XNRaW
T+43Xss3DPoqCdwi2A9WwIaownBLm4Zv1Oplb1Trac7udi7qqoDbrj537Ss2TSUZ
WfLoWd3HnZv7AQIsIf4D+bvUlLIz5UYf2aWfh36e6UZ8h7yEQHf14SSSLVLTmUWM
lI6tivsVFbKGGVByxOn7/sS5cdZEGgx+KCtx406imn1q7aW4g8Fs+it7B0jiv+Dv
kfsxwkYgbESKAw4AgEkp7UIUsqB3ssmgpQXOmwXJR41gnOz6AvOshQF23xfBOBWd
+mTvoFMmxBP3vlodxPoCa8ISXLssOxFGnfHE/IBL9cbkj1jfGZbHAu5PUxMBbSZX
V9M89+/ksYL0ScTkkm3V18fBZBcoZY8rUprgOpvbxdXuKyCDgHYdAo/TBa9x7Syx
A21KLgxKY0jVJiaQ0LJl3hyuDkgUQKPRz6yePkiBB0Nxc4X/6zGRVMxvNrTMzgZo
lc+edUcOuutO/aTY8uF19Rdze+xyMVhy68XjZ+nMI3Xk04ekgyplZN4MsUFRswiu
yRvWveN1kZiqdySD53vwpv8ikR6jCZbrPQoGWI3EDakPz81FqQqfNeATiSLNsrsH
oH1QiU4YY0Eu2tavfX+dSlGX74pcLmS79ebNDxra5l0kMzTxqdR1vzL0NeYjnZOe
rxewoD6DrhfK6R9DalTMXswKYWOZ3aPSVzAq3xc5ZZYwm68S7JSGcrJLwgJBbqjV
YNhDI7yMNm2ws0vgBW6sJnKXIzqIJ5Y/RS/g2x7ATBLMFgoSWDQ4ZHyQCPQvAg5w
uArJoFI33X94FCv78gpUCAziVsrrswCj68mKTdsGhXy3NxwASRCpe3dF78EHo1Uh
W0LIWH98ltnGjFApwNtF6crUbzr/6FnOIJ4WEZ8qPBac31u33cBfC/64KfSZUIYo
Rv9PN7wgKj3nU5QfhbGumQN/1OyDHCl04lTgcKb8QZno39UO2Cb5nfsNUozfYp33
qKf9w+5xgTSYSRva9I42WLCkDJR6nLLPO9qAOsILAzSUvLIodrC6xDkfhCMF9r9q
/HsbOYA7pOlxg9ZtiwE5Flc5NIfLEjVhafn6RD6aEEmfamdCYv/YK9WEw1NH4ZU6
kIw54sxo/Q0YiMWOO1dCXvHm1L2duZHu6Gc4DVWz6qpOIu73mtKa3ZyvqaEw0zFQ
fVZLddbv4KvPoA531r98lsaF+7erzsnq5f28e7yCuT7pQa6iuAuZ4LzVX/AqkuNS
soerCKf6Lmw5BSqDx+C70oSSP2qZnF9OJjSqPmIlpTsOw169S2eSJgmFO0vW99MZ
pvon3uaZRRjTFJ2jg2MdhltTbs6fiezSZJ+MgM/jKvPMiIomS2MYj6i08LUbssTA
fFxJUKjGkyEAfvwX1TAYTu995K0x4EOPYVIEUWDmFgwKiKfHfm0iK0YyRUmH6K+i
807afP44D4wTEaxZcqfC41Ksg6yc+XxnqFyA39vRNl8/z78ceOzLsEYxtZv/GQp0
IE+U7DvY/2sL9F4y2rdfAVMnzUjjWUYxLBOueXG02Uc6RwxVj2RaZBRad+PaQq8A
S/zSYhfUhaLdGO1Uarw1CbbjN4ZVzBW9Ei6HejejQq5S/HkpZKgE4TvRc3aJkY+K
68iYWFqJXQBuRFIWVs2PnkSyneFOF4UKs0kePKgKsJYWsb/kQw1cg81rGNe4e4bI
GWKqrSZnE0b9H+PlTNS834dk1MwNOphA4i/ESIxghgOgYoPGG1Ftb0im4eya7sBZ
2TllJBQR08PMjOWbB3CeqydN9Tpgq0aCN4Z7s47ojUiH0KeBiGH0RuXXFyFPnKvs
PmG5zeeG3ivf3yiIvZW2j1lvDvj4/aXQz3PSx76lTIoiSZJQhZvFPdGUVgQF/NM4
esd3UUOdPpQEZmMFuHcHU/CCcCjcBK6TYWQsQO6LJEi7iUQG0vPrpwmcsvH8OKa9
NpnQWb/FIfTDT0uFyf+2KxbUpLFIWEB/cIMWFB4PEM22e2liGWMc9mfkBS1i4icl
F2SBWm8SpcC4nPodlMfV69fBsLKosrx4dcRcKHgWX054FqhFtvKrhSgY/cBb2VNK
4cCondaxydVoauFu22Y0wc073xr1OTDT3KN78GCCB31CF8xcvzDMj8neuBxsStxf
+9mX1JKQ4T3gaZuOxjKnkei3vgTA6Db2/5ZMaRpf1zVfKs1UtBRTn/q/qJTYyxCn
QmEsS/561dyV1hAo83TdIFQOVpK+RRMifFI04vlaleGiqji6DV7IrNWIT6OkPzEs
vl5CDTOZ6VyaboFC5ROH+Ixz81opuASe30HHaT/VRXCkESVKDxgH135bgO/g/Kv1
o3e6HSp4XZb4EzuxV4ghLAbrEIsuZ/yrYHuotO47TndJ7vu1MzktIqpwVVn+BE/x
AjkHIQRt7vBdtxa8adoOlgFS1MlzxX0BOS+erH0lj70H+n2XpQcl2LauRBojn90F
Xb3zyJAHqT+n2RfY/8eoJGb83jyoRzaSxcptu0SaF6KxLWwxM7vqgOhN/pzE3Ba2
hDj7CjP5ydeKay/jLaaZOngj2HZCaxbT7q9WyaeqF8c4Zm/+7xcqkKYlvAR3NUwZ
yKHL0OBv1mxs96FJEMHnDvrob4/K8BLKqdc/cTbgH9OpsZITBosUSdDtn7pa4bHO
7uwTjqIwFB5n7UNsmmZu/u5aFSnQYrCI1p1/fuYBhjBT7DIdYTWpOEpn9U0gBc6c
cKAI/tps9P3PBDU5XFvP+gLdmW9YRchBpXWdhuVIV8thdkrtfGKLkUgnbYzx6HEH
JfN0io21QYW5b23M5Ib2b+CPHsjKWv8feFewtSjutU+ovI7pAAG+cwoDp46HJfPm
OTs79FqDEfosPCMhJFcrdCQfY/+VKL45jWbo02XklrRYIgtUIRyhvLDxsU3kaUWR
G/q04qbJSpA2kH/BNIf+XPAkgKCcAR5h4E9kNC8pDdVfWNK+Qo1NC2J32c5QmfDJ
YIXhgW6elOKAMDwSqT5OnuVLC95rXjO5VNYCnEbYijJQM3QLMy6ZmkFqjMDFhKjv
gz/6tFwy+VGG8pRIAAx57s/f5uyN8dqz4XddDavVsDKNjGGMsh0ZhYktrflYKHMR
p0d5eCuVW7iLHJNPgNmEOjr7ij5VuSN4Mf7M472OnQgPeH2vYE7v4RaBeJDYRSn3
m/I0g5k1juRAqOS6tjnNQs1xipcoOqmwHCSWbvwv/CUN7+NVPyqvas1o0e1B07Md
jj2EeNX37JnA+sEN5pjJJHPANexBrpIv6RuDkITKb/CL4wRw/bb5wU7WtYrE4xe8
BatWo3E6WTokVXirStkPzOnmjOisf1esYIf8CAlbKlEeIrrGI/uoE7QIbVYNRcIH
De9OJEt6+0sRERdyoelfcS9tP95Z+MIrvZLQ6vejE5h1eo6khjS7cV01b/2isOKo
ed0+NkX80XfcsxyCw25Y02B39V/AdWiSVisqj5UVg+JrAJcVwB+8O/4FpONbhAGS
lj97eR+Dc0gecgoGfAnpbI3Yj550IKLxgyQJvEY36EFIO0iLe47d9xTDe8cq+pSF
ifa6xN3dBPcGsf1s76YdPn2o12Tv+CGTFil0AOwJWSQMYl0aWpmyrPY1l9/FjFLZ
Dr3xGyMMYqP4Ym7yTIKeanqiGHpntILv1xFejPuCHb+ruiGMGw4ZNTGy4MKn71yx
0zblf+PQw8ozgTUOQIipjVUUBe/cIrVDPeXb3KklCVGPGjUU0MUlCwz+EbMZcxpj
ZiWsbKWVXEy84hU74tYKM2kk0jq4adp97ex7Orbk4tUHWcskrhcgWVWkf06AMfPP
ol5dMBUazkbid80vi770pKWrNWOgIMuthH+AMTQbvSTUHkbTXpS8KA2jkb7DmDyU
O/OkFNHZo+97mEGu56gSwMnrZ+t8O08bFs+D/to/DFXSaOoFymZkVr1XHyC64VAi
6GFCOMs6AjOdg/GhNLUjitW78BKTeIcNdR53b9MBsnYoozt5sKSOt7oZfMv+Ger6
+nqncEZ/4axTlHh9VzUK4hx2RgwShSisxv8OGgI3qIPcObikcrhjjXIoOfjxPcxN
tlntmdvIv3JvxYonutApfMCI2iKEEbVdLSxhGHE1cmhMXW3m4ixqrj0CqOrzu2Kw
jL6czU3qHHH/bIOktPRcoVIHVu1leOPZQRrdcUekwiU3U8VA4Z/3Onx4a4ZFaBIo
XeW0RzLL9q76scYAp8rV8THQE0p2tyIR5DI90ngaUYrh15/AViMzINQMpv8cfSIP
pNS9WVju/PunbC7r8kpy+r2ElwOmETB9IZmm59lqVFYR/6jVU+SrfMLCwAPjm0uP
L1ahkvf0DycQqPnsFWuU6+pVGr18ePJl3IaubwsZy62Snn/17MM6h4JDookFUs39
eW2g2RmE35WJS/D+WDMZgroceVYPhRsvue8hf0BqOJBA1hwSuTT9E7EhI3vn6h7A
CN/fBXIlia9w+jdWx/y3DYAuKNI4qAL4xh71CcncGYQaG6NYtMb4edYYu0OHEXvY
tEgul2XoNCPQGPaMEKQ+aAh9xtqs64C9Ufbc93b6DD6+PgSILJa4tDelLbh6q+Vn
zjmoIV2Ad8PjnKTA2UJOPijSrGJgdqiryuEJxawVE0NZT4GOI8V5qBt21KUKHS+i
oTc3lTy2CoAUnznRcNDL1tJlTJTrOlUEufCRMZzpZOoMxsZf27B6etr+rUlcb6Ns
5aYBaKsYhzHlgup8IJVd/NPQr6/35S/FE+mH/DJpiRAEC0tybYX5gZ/iEU1PIOac
9RIMePZ4hOCnLcYPRmH0J/D5Q3xcSf+Tw/lxESWc1rvrbiYeWJGuZ/Whsh6GUNoF
B9V++Mbm7szQs5jnmrlqLnhk2eXcjZiXbGgcdrMScQw0p7nktPFcMe3NieXFXA3R
4KhZYJnhVWhlyFE3WEd5STutWOPk42LNYw9oNMGsrADe+QB0pcXnXejHfANSAnq/
eB3LNW7/7D6WN31wcBh/1Xte38XpOAzR4/b72wiU26OhWgN5p7ANcI3oPqHzDPoQ
+49QT4jzcDfHJGL14VlQLLUXTsxhD1l4fMQHqyJM6IN0AIcSEf8ABIj5sgrbhXjl
22SKZGh9mQ9qvnf4CEY8yWGsG33ROLrMlzXs+YC0yJUa4Syuxs4lA2X2Pl6JOpFB
Z6WyiEA53bsx5vyRy2FXjb9AIzdxb4t8yw2Y1F+GuosoJBHjFxPFPIdWNgZAFgHm
Igstn/qRip3qYKZnMMltGvaEVbWmLc7JTM7azR6RUe3ejNyAU4lIXVjNZxlhjb+9
VXnAoYClnVeQBucoBwt0YLTX9JM/RXQHVl8+xJAfl5kVH8i7NBEHB28GsB++Vsbt
DpYhTZ42C0Bx4Qe83abHCdwEYpVkx7iXsMt7kWhnWHkA2GM9rqoQG4R7XZPuZFkt
kevH8m93BJQWL96hLdquPqThFIU1zi+7CyCehcGA6wx8g1bkgEExxOxwU+qcRsM8
aB7O4DFeDHu3LuiKc5y3PowqXgKeNnO1qvSj4Dbx4e7BZTDNgPzsfSB7Pfg/kkt/
5Ggj2Ykis7yJ7bzshgE4rWDbbr3iJ1mJThVI27zrnpBdOZkSTgJ+EpZTCNPTkcqq
yQvWahzRCK06m/FOJQ1C2y6wjUwFy00eFNhscGz/KXyOdbP8eiiENDKWhZdjr6lt
4AY/cnt8NbTqGpLyodxt3nyQW3UpiGtWC4sf5GJTkU8+GH7CUh0Vog+fRR/dT0h5
aUhSJCHyqyxavqCBjsbE/sV4PxpEmFUCfvYRkTCCY6+Po3j3K5Xp8x9MO7i0xSx3
ZYxNOmslzikR/ZZBimzr2L7NBod3VjT7+qK7hcDMoGoYl2gtyCJnEt6CQtLFfwqi
adcKTmq5TWbNoAI20pU8ThZ2HZ4b3tVAe+cXNLVfBjkt2mgFQt30XvBwfKeDjH07
T7myZIUHMGg8FSGskHTAXvpQxxjg5Zi5wzLqqDmHk7QCUvtkCEkgZk9mlRto+iLn
+1uzaGY8zClRQEgKBszkO8IDL7DFM8D+AVJmcmNgh+zB/q5GJIYzM+p/5B+IqLW5
xSFRvRwfVTA8TSq1siKTS5A0rx4JFDqhiofcu3MJjRURNAh2a1aXKJqNqUKxUTab
d711DaqW7W5oN+l30OYAM/phWPug8PHXP5jSu6F9pNOwmhinDV+B1qyB4/WQlsh2
AoHiW3S+buka1F9LKKJ96uUSfpwqsFDPDUEcOgP/ee9eoTjERj5yI+HsHIGNaIHU
o7AoQ++IS62BUyRJP4PdDosykK+JLGZsfZEbuIFJMap2sIFMOnlccdBGnvsNXLcK
lUrU4vSE+lZDfz+RgFKJggpa8nW5sQeQA5JW80c8RKQgapTWr54mTcXIJ+HC1D9O
5Qmgac0cA+zP0NmoRizjKe38hFmW6E9FSnhbpk3uAtogik0D2vNEUCLj6IysjS2X
JQw8vKoB6ZMf8a6fvGAoVMxRqzLMAs6ng3bcg7z3L8fvDbEJuPwxPOa2EOXgUoGM
fEuVh4lM2zulnoO0phd1VAG7i4ZkBTZBJwSOxASB88ez/2X4QHaQvB+81V6BGC8D
vP+23nElszPI/NHz6E62cj0CEAjOXpa6075E+goswM33Y6p9ZQWrLLUfS2AA9VYc
FMum+AfVVoEgUeap/CC16u/CuvRG7sUczuHrLnJHl/Rs3wPGm8rPKYfsGbE4OPvB
rerWrhoxqTOZWukjqCC58c8cmFzFFKjOKrnveeU+NgTmPoikLpIF59+Mh6jnaJ6z
j502RqF+vYCcCLyBBND/+zIaUxi5rZoIyNgMXc2olnvYQTTZfUO1Yt6Bqx+kVf3g
O2UnylyiPMJu2Lx7sNqris245k2mPe+Cc47YTNBHk4SpGHw8iQC7sSzed1tm7Vss
vK5DtZd1XNGIozcfHOAsEcVISuWFTH/DX9kzSbeUl1BoCcq4OBTCggJ8cbe7vZM/
1xOzQnH3TbvQJslFdWuh3XvwkTrnnvwE3bn05uSm/D4A1F5ZaE8X6TTJBWTD+ePW
BHOT6pcKRAgzlRzOoemCOAKN7t3O/siivV62U5OgYvRfBXfDzJPl/5IoWHxL7qE2
tq09RQazxI5OZi5k8rD8xkEwpXWOoZEj6E+D3NP8rMCHz4XeLw9SXteTy9p4avaA
StHLQDgoFQ28WPbS+Uw580PsJ5NC6dArK2S184cndvPlhUcK1+TL7pv9XhK4H6Wt
6fu8teW6GygrIcOW2Ep4rEaZGTdXT/d1B1pKqVWgfbp9/JM3dwX1PKU+9XZzdO1B
dz+Aif4stG86zJvcJKnUkbnnWsl9f+hTyNOzEm7Y4fNshV3Q1D71BdeNOf+ecgiI
b8tXKnW6+3DFJ6sCGHgg06SWgIdcg7dnFRFmDg22X3U2gwvTWIbUI2hb1bKPtqpz
ftJcQHM9AmjLf2W1fUFSx5QLTFxxTX2dYwOErrmjNIktKxGHWoCUV6LtEleNzmOr
2WSRx4l2g40Fhy4WPiD9yujN9i2ZDf5OxLjUinhY8LfGaevdRIrJEzhfNFeiHNo4
jcRgyN32HjMKBKH+O3iJS+CldAb9m8ti3xhmbAAvmCRKpK2mK2HGoyROy5v4c/cx
2qEYnHlhQ4YJbzvv4tz/Q94MYbJrCgS8HmdqVJSFepCuHOUJ+sENVqS9gRS6CrTS
KAF4j8yOn9M1fv58Bej9oUQnpRQ12O/drGQ53cG2cDSoQzrvE4+DGLrW9TVbNmX3
0UW3v2/VRysRSNRDu5DPCbgYdQN0CZw5rzqyWXDfVGkKr2RLfJTEyG3WVg364KZR
QC7N2rEZz/7i8sdPdug7gfFSwjFswjhgvcad6LBUqkbB8/UsPk3KMegy4/xOEEm9
5nEnKbfzwnjmFMRRMYEaSeiYkfcRCmE38iYJeCwV5Z9a//3HDYPiNbdO11ceIl9q
byRe7MuxWo+hGleRym1pfUnWUzwnoax9aZiXMHBfRJ6wVwBnKYYj67oKxXpsPu+h
bzoOWuRRDrK9vinFUqDNg3tsSFtSWZxhUT54dnsdxyr6RXOThat8/M6lfjTn9j3l
U0EiRR06cVSK1WrfCi2JDR6mcEjhtRaP85TYLxYaoU374W6/dV7TIQP1MQ6taf+u
RlXWtNUhPcChxYD/ZgfkpROsDPCSjWyl4A+FsBY+04hHZ1u+z2kI5Bwyoq9MZBaJ
jXwID3HZByYmwTdbWcOW2KwRyumC9j6f7rS4NHyr+e9Bq1hlJFdtEF3F9/v+k7JM
AMznFY+dmL6zARJXKsKj4Qurf0rIQjbywq1EU+xt3JFihxalyzLasTZmfbaIPKeq
25JPSrBlnZAS7a0bghB2tMQZ072kWZhuDyqikExvLgmmcQiXLepoiQwhkwozcL8I
EUjoIHNLc6czAg5Kf0YPnXS4+hsGG8tbDVhLFRCeY5GEIiVSr6Tft8xs46BWTF0n
yrDcfxFC5n+XFuvwZ91+ly+CsUAjTtP2+fTCkkVBtuzQDmrymAbItt5yQLZeA0ud
EBx12sBescgVHM5aNTWzLQ3cFzZ47Bxip5BPZWU0D4KpJP1q3G5/UbSowAygg9tb
+mJVpKUbXqiMa4omd6A6ENvCtxldahfOUsDOgvn5Fg5DjDmZsZvM5TpENh5kiJT1
1EVgtCYrKORwil36l0/HlrRE9GeD58F/exRiuI13VTLdldiQAoMsxr2kttWAfpaz
tPKWSrFy8Gr2WY0CpyE5bWNENm0f9vUrp8SO0pI/jTliho9UO1BGXmE18DoS6niU
aRsK19I5TXWo2S8H0EqI9O5Sni61ngR7XUBo5ng6mwu0ebol3YT+fkF+PNtWMgiP
5vED4eigYe1TRqp9SRwtN4ND0wQu42/HjiGf7KsAzt1E0kvqNKtpKsBp6aoM6QDp
JVd1KVWqUz+IctCwNK/WRpXJD/OqjBvJ2CDpk99C/loHLYP21vpaaUH8vATrD7Sw
qHr7qWmp/0nN5xIpOMlWUnawlxmBjM5ex+rRhVkPy+uxYImCWQvDcrVpD+E/d3WK
EduPSSv4E7WYVS29KTYQDHjbM+7wnPV6ibWFA6UdOvtVbPdJ8RvcjV0BM3FEiHFZ
XK/u+bHfqA6X5v6wQj09Eve9baC3S2wHzxayVn2uEoUzRRfHZSJDJ4TxaLOz76xI
8z1NYBnRnJnoC8kwsPUyp47w97+O42r6StXRGtGwJVGFOnGBaTLHPzUxjg37cAv9
YU8iLWiGwS3A0JfCEAoSiKj7g/ohAWqV2q4lE8bzXbNDVvUw0/yX5QjyLsImkDFd
pBXSEM0+hMYgpbIUKRVB/DeCGQkLHLWixTqisuYt97B6Ugtn//XW79voVLVZyCpL
r5HVnUAFmdZP4t2bj44mAqdObuAIPyRzGm0gxlyYhlGrKDTjEo68wqiey2COiu6o
Emn7zZCaW3ZfJofBb6qH+CNHt2xC/91SfgRaD+SgMAVxxTvicAbolX6NoMOLPk7Y
ShqeYC5cNjCnPEmOWObTsFJZEUwxfVCv+BXcv/QSe7eVP2FBzUYTVskLiBoYD3lp
jxai+4ya+2qEYaLPy1Uzp6ShT2felGrsxgEYotse7yGdHvHp4Dk5r6jXxSaOCY62
Znx7ue1amAZq1TdxC27bWTc2PVkyZQZeYCe8m/7U8+z1uBMWIuIo8b/pc5rvpk8R
iXWjtnVX9VDtEBdXzFwk8C2Bmj++GmyS8iDWNohi6yWP7c40/EHA+wzW3wSZR9iv
1YQx4NXlZgZu2SJLd4WM0AUD9Lq84ESESC714Bf0yCTwRfH+CMB4kV2/lfjXPyTM
IH1MBvBguHMcPmtNQU+NQlUTWWHaExh4B7UmJeOmRAr0f2PDNABpw40ufzUqMQbz
O6Ssm+IrvuuN2mCDa4zfmMgQaWhV34mLXp7cRTZwd75RMj/CirHsdtKC2goynAaQ
4azRZ2PazA1vLjKZ8O2rZpu0+Xtoc9cn/eGdO08fc/LT/y04acp9C//Tr0U860jo
148A5ZNUPxEJ8o4VMmXvLE/g2VHsk9ngo21fgH7Lqcuu2pvujj7fwefCL0e4kmum
CQ82RX+DOvELbATTeWpLQgzy3mjoiMCbgUvZTCU/TbpyXe/MVywdT2ICZYDtplXI
Nq/Ly5yErge2JV1iQrD34Arb1XDM3YEF50R9aZaU8mguNQxMQL+tGEd/oP1MCFcE
uEpm2eUREIjA/OhBQhC4l8GIDvxxHUYMKA/4K/z1ThMoWT6logIwzsgLvwcmdFkU
TZjLDgdmdAzUyXkog3her1DgwgvJAD5RQynuVWZZUk+Xzgc7xAtr9l2WunJ+dqCd
rGbO6thYGBoY7rwHoHxqMu9V4c+ek+Hylu6XLuWKsW6/vcHa8LtiOj4Rn+fuelmL
zzV7ClJpEDGhZq970CKFTC3gs2anj8Um8fhte7rOAoVqr2n68FX+pnnsXtV6ygyP
uHK3atoh3kjclMThT3OIoQ0NdxkoZEFqv+4eldWt77w8KKndx3tsgKDzguevFN3r
zON4J4LHS0NDGiKs+x3QBqWJKaMqiGCakdQoBtIvx1LQp5NArV2zKFuh+sJWDo+z
Jv/Af2Gar4nspwpEv9kqodM3y951Ghb5Fzmofu3SyXgbqIEMZTageIOVkE1sL0Im
PqkyQt6MnIVK1yCBvndehXbFEeqyImnG5+awakkFki99jNoE884kYfx2qdc6bOZ8
Xa3pbsq3Mn+VD950rXEMSlz+TMDL6k2wahZwKptMRpZMCBQIxvjy1jNhHoTf6f5O
n1HhOm9LNTvJacFJNOxhnNFwCBYYg+i8eS+inDiNXYU4ry/EjHc/kNxibsmud8DL
9WEXYSNQq1jIp/T84akhcvjan4ZFJ0MRwLy9IMDpnO9IED5HsKET0ZBs+X+rXgc+
WxVq5xve+DIjPDTNW3OqCI0xre2yM22KoOtNSRRqDAVKBFo+NzraqcacSF+dadhS
6mquf9f8HEoy/vSH7ZI6E+GI0W/8cEk+IiLnlnwSeVad7HtD1c/3lBNVt59RSeuA
U4DpnSk4hKsgimHLKLmou5zKbw0mYrTJDNAeSzsaZpiWnvJsqW0TIebQwDslbYCB
1k7Ht0UTylZgVo6lDIbkVAjzgnOXwSbSz2wzPBuBvPQiI8K+f5tsigdCwkSvQdMc
Op5R2t9SAmrs5uFQkL4ABGRrfWEcGh3H2/QZs0s87I6/jgCBNsfQ7jP/GTLv6nwz
LaH3IFbT6Ghsv1af5Ej01VmWg2JN2En+P7I578sq+eQjlSZLBtDg6pvOYXOjM8iX
AUhXYpMzCorj/RQkSgwzTi28ypl0EnoC7ARd64YIm5uhH6EJbk4Ke7VxZ+QPV5US
HvHPgXU1+3ix9hZXOS2ip9dKEEe8WENdIywhKqafk8AREPVUFVTtxre4m8fXEyXf
4OvHIyIz4aarTXD7YS/o+m9SaeiR/tFcnDdbgtde/5Ukdei7KlwWswgol7iHAup2
dicCt2wTZnFS5/dcs/mCZPrU3dRVjqiYLtdPASZcYj7rgHMzbNjLbqzqrqj0FhB9
FNda0wTa0IGJhv9pYzb+h7ey/8mXPdNVxuk6PH2crN/ZKN9fS5KdsnyFnKS5upSy
kkfxNv5Qy7ZvViXzvMWdQ9xnx3t1iiSh+fsupf88GoVtP49FLXyN2svOI3Eh7v+o
wGV9ndXr0Ihk9I52pmdtuALG7Yz2wnOLR51Pv7KNkxSQ9QWw1W4ieFTQyJJnWYlo
xBVDK52Px5il6TAGQnqG+adxoR1gHzG5FEO1vh5pK/8LkJc4lNSX/yunYeJjZy69
C/i8P9ZWnZVW5C+1xCWX6QI/c3/8NbL3ATmSivN68/+V/Xev0B7v9tI6AENEhtxd
atXBJBOCfTT14xvkqQMdBe/B/o+Ge2uWxdPDIHlf2iKhoe7YQbPVHpdnwUE0+4IL
AHkp/kGzVzdvHErrfFWMmmDUsQEIN2TNXHZtzvMADZsQ/KlkBSLX+Djrd3aZQAYA
`protect END_PROTECTED
