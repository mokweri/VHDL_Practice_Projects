`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
womsHNBdVbdkUnKVxVL1wcf/q2W46a0+iRtKsO7bDon12tArOPlv8u/w1KSaUxbb
HarLdbPKoBDfNphcBIDePhbBIsHKQx/n2ixKHUy2yhPmWXn8LUy/tCgKGanccDFw
ocje1kXQd0M8tJy7pzTZ14VOh2gsjcKjBJ2E/kxAGOXm6i3SCJ/AIHbcNSxvyZWi
AmAhqFIeKnZn+XESHRWGy9J41NiWnjLhSVPzrhJ/ls0K4zRZUVPijy++3FRf972f
sxjD85pq1tKkB+5CZ0i2RhACKfNexAgyB4XhD+Vpd3CRPyj60A4eE3HLboFw3XP5
v9qvZWXAaJbejSDS1Q9+kn+CkCwilf1ZcY5s3HPtbqsk0ziyh/qDZDrTfKkogk/e
kS2KhsLlbavsTGL9Ie6eK8c4hlnO6ySCOnz1j4ryPLdWxRtyD4rEN0Uwv8GvvKxD
/DX1VLJW1MW8LzRCt5vbb6l0LJclZRTLXGdVZ26yEQPREE3HWsl9LrhGdJSDHk69
hPYsVyZOnDhphChxGDLCfU0J8XnwjgQOdXNUnpSqGr8tDmuLSJ8L063xTyxRZrFX
UEOqa+98jk6mPkCU7xHIo/wQk83Dc4rXqRkMcX4r8PwJKMIGv3wlGY5U7wie6p0O
wAFP6EuuVmKhhv2etwgQVdK46/PHVNk0YGloVYhtUdb7I+oPvXZdAeHW8T0tdLvM
SA9arCBEbInKZrtzCRpos5ubtOgTkRD2Z89gAxg1upjpIBcVSbUZdfZjXaH0iP94
yr9sMkC56HeziXIqpZ9Gz4elS1ywsBtGhYNg7GdfRC9GvkpZfkjXZv3d4wNnXQSZ
uUre7GgyAg8/vWqguMXHKITxILM0l/5vc03vo8k08rAIwodSPy5VKyxf0qnThXIj
W6OnukO/EUbZOzD5tftEitvOD7Q/eGHCV+yiqI5lMHr0Nm4zzvyMjDxpFgrbxZhJ
K1T8XHGS/enprS27J4eo8uqXxXHsw89pjQW+7kIleNHUmJWd+UTp0CGhzrXgYhP0
OCjfBGLWN8pTpGe/fUjtTCMRF+2eZd/Pd1yk9QZr2/1ruY4YMXNkqMkz6TSN7g65
/5VM+uAlzmW3M9Xx2l7gdaYPtPK1uW3Ma8m7jrExqSszm3qrVV9SzDZ8YXnOJnqp
/NVyeh1fsgHC8XfgHJ9upxMltV6eZ1m5isqp5HoeFI0rcq96hOMrRHK/6HlED3P9
ityVtitLtYINfM+c2m2Hy+cIukYBJ/OyUgyWlCJCQ6w00bkX7oCjVrIXsqiTYxWU
MfZPWldCLRkZfcn4CEJwEn7Crv/apvx1cl7ATwHyrctCKhy1/rTUeUL8ohMh+8YK
BI0J/H9/7bqtrgpWGoxa9ZL3UmE0CZWtpTl414wu1uuEs2/Q8xMkjp0nLCuSvN22
wJ1+at7kRwcd0J5tJNxcETgBDpdVFXVUD1G5ui7iyNadas7D+LKOg0FyWZ/GOyZf
KHDF03ed/+k5kzGs3QKEDXSJEtz+X4myuormLuXNoE9TtQBrVdsvxIcP+1l3s5md
BLD0OIM7oz8rrBg85DRpxGBQUbQzO35pxOHPvYszkVqtqhYlaQ1oH98UccWq+RCE
x7qe6HOtJjsnHRTSpQEq5t/EMaQM+9B5L6uyCIvyQ+yj2aiSoRnh2TDjqUY1PY9d
gLEQE7tj6KGAtDajvAkKp/ped0cGY5FIM1Yqm0QR17BLwQJyAVjhP1/DcZ8Hr85b
RfChpmrS0X3vzw9bch0BKJT6KxHoUCRoCtIPnRFXWFwEc5GOxCCjbN59VlnUV+dz
13z0EETKrF4cDJRDL2z8messIdwMvIrr4m6S5paXCPlaic/hMDyLNEvCN6QXnxwf
O5STxEgvDeJGlWuW3SA+BLfxESHrsbr1nAbNbl2brTsJUzoYY+j1r2BVuNiGmNHG
5zP6Ad/lMJiMq7YTc/Sw8bD1oQ3L6c0rqyhyV/5Jtm1Q7iCO4bs+fGHLICKZxEH/
WrunTvcC3gCTC62W3IjUKQc/DUfq5S85DNkhCnbkqLjdi6DTZQC+wlE+gMlUJblv
KUGMkXJiwZKoboMUzGtRP5x2qhNs3MDduGxnnRghyl611DQwRD+UIRHEtZzX6Ghw
iWfWQbsvXkeC/WCXTrrymEGXz+4owqica20qYSZDskqhsS91ls4f8/XdYGTKra/g
baOKuyEExxNOhC9854vNevjoh/nw/GnWK/jXzxStqzcA2N5HYl2hH9/qbqrxQx9p
/4fR9Kpbdez2+G5MXwFhyLSWvcT7xfOXLFPRA50INeWjG7Xw+ztajBM2CrT0H+Nx
AwLYITJHXdrtteax7fUe9x74ZSNnVLpyikMQKjSW5voRan5m3aD59iDCJlJPfeQd
gO7HcL3PRtJ98xIDRNnv3S6anaBcYvEMrJPhpgNZItvvSnUMciyNjYKS1nQdzyae
TxQYdS5VDFU/QaS492RUrA0nNy+h+WjyP3r48ujkyMCKo/hwnFh7ta+trZfOg+0S
Cl9xDqkvP8QqH6moboGxgrTKqQae/VSZ4DuJwtYEs1QkO6ggYRkq8xPa5MxJW1c1
4zBWqlN9DZLluPOd4maDLVVUt/vIDWeLwbbkIZS0NCHSx15D1avsUc7s9X57PXm/
toF2eRAIhj7fHlY4qr2DrashQE9lqW8qECn4n3GZ0m3e2kS+RQE0xA/fjxTJwPjP
1UqjlfF789Rc9ZtnJvJP7Qx1vEekohuWGLEg50T6v4fYqf4ZJ4LFwWAfRcMh/XM+
ZSZHOWVALXwKzfiDvq7UPJM4cbHJMz7mwxsDNXieMe0zbX+cyAQR0PRKR84Jqh8o
+ajZ1FXQbXwec25jEMG45pKGRJdVkUhLX6DIhKIO263flYLjHrBWwpxpKs4OFD2M
Ngsz3sXWuh8hTsUbjdm+jRvQx7iPud93cxgeDwR9kLNUDSX8DYr2yzm14/t1HFjj
1xZliCaoJ2eWA5NQ/Aoxb+0k/jTp//+ZjWTF3cerWxNT1gVdD1rHncZxmWfVO8+5
dV/B4msdF8PTDlRmkM3S9+t2vGskPlJFCCdFd+q2AX9WKBuN/uCMoASh/66GxMwy
BnJLstPOq2aBnTn1R/LNCHNfz/btoO2BEfbOJt1wfnK7y4Tkyj22k9XG5EGtsV9Y
GvTUr/BYfMBJPgFkGDgd6oX2uoFYFanYlZl8WR+sir8I/zruHcw1cDl2es1wRmV9
MqN/Zz6CvYZr3xxJWUiA9Xq8+4s4UAR4tqAJuus6Hr/kaFNqp/yR5HaDpdJD6jxx
Nmxy2DQsVouRFeTQiXpbt1yMJblNuYSWlzUyJWTG6ni8ML+gqz7d6wDXJ63nuZzm
oc80NmxwudztJCA23kWbltD6M+pv1Vn6MQdxUMkyNZNtO8e7IMw24Y+XxkKhcpR2
SIDKnAoq5Z/82IG9YS8YkZzi0ajcBGDb4imzOewd7AFb+UP/YcymJ0VnL9qNJdRj
Ucmg2+QDodJTeKGyzYxahpVihJG659tyY9VoI8p9HI6Ow4eLKnhcpOfTiUolHdeS
`protect END_PROTECTED
