`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E+muMdCvNP9GhB2G58/W6+yfgIVAUC7G0vQrweGYhj3GwanDWv6aTJEqZzLwfeGR
USxb5HCdDhszCnwCXLVoykzeQd83XsltQyTID0N+4DeDi4ZUs0HdBvlkAv+QFnf2
CKHEbVs+phFMNpM5TrcUq3eXQsxMy5Dy2SCMJGLoyfp3SHo2m427pQxaYAV/DpLm
sITQdVlbeFGkbCG0DZXzWE+ul0Gmfn0TPmTVsTJq1QI5/DqcHKgPYB5ABU0pVA/W
i8BDLtAQfPSvWTVUId+OksA1XTLfkGz28X57LVcuCiCjvhmEgndF374/pp+ySqeg
EybysAz9L7z70bogfoma1RZsqZYUkWk3Re4mbKFixcej3FEUbZVGtSQwFyn/rcBM
2XidwnXzOjbr3clNN4qnlljGgj4xffIxn1p/m5111FmiFXHPmnK8sRTXtS3TakIN
Ty3LQc85iczhvwZgiZv/1emi6IrfuhQ8wqE5o5hIcfYaPdKFWkXzLgK+IIPuytP9
YcUvPHTKWRqVuCfmVZuCFEQkF9nrXVxr9lMweYH2eJ+cRQ7KIKwLEUMeWHIiS+LH
G2T6TnNTWIAKiHN1ADLCvL5ljexydllNitCAZDmlHNbQBPs9+2tKVey5/Wer/0j7
cMzHTUrTI5gJTMgdPFthgonDsQu0EC709h9cqrrynQRzf17IolZzAmnHUQwHoy6m
cJXUEvvkKNq+T5zP/YjOMdw7MXTdxeDsAjJP1G9aKCFF2MkhWrBKjhjUE1ijHjQa
5UHh3q64aDpuRuddnmPzp6E/nCpLoEk2ch13JaOz/bq/jY51FattldgwYrnabfDt
MDsOcmdJD8rC8v/igDpBaHbRcwxRO8VU0LfJcRRhtmkA0GUkBpcOdaKEk/k/CU5L
wtFxWvrOQl8E7bb3eiXLJ3i9mWIxRDFjG5nEyUNk1fQVYpaGGxlnrUv5BLpnthyZ
HioCh/sbkjx2QFOvqcYVu8cWUvg5wSewGiP4AQkcAtYKJfY3xQ5POXJKKB505aFf
Lk9fQIct3TQfzkS735VXIOmlx5eD8xFGb/DsP4LJ7bKSPT6+8OW7TTPdzMx0JgpR
4H6eGzSvfF/T2ktUMkzgyw70S6efrtNTnFLlSYzLh9CawGKFAM93iMxY+bE+G8di
+slJb94hr+Y5W7XyLXDpvsWMQp1oI+vrj4Hx9auZZ+7qyQ83Ju6EXpBiulvxZsU5
zx3fnvvft3CBgzvRgdwTCcvXzlGLyMiy94s070LazURfMy2An7Kf+EeryKlOSvpf
ienDw/TMXo8wHStH4cF7E8tciWevgRoqcG/aD2LT1TjWjZ1q2ylZIgCuoxYCYqSx
C9UsyAmAs7LhelzZdJWf7X6u3utQ3x+rGYIDU3E8XZ6iOKYd91t7sGmYRrDzZVaC
xWQh1C+IYnf5oG+fGjjHxxxUK+k1ZBVUj5hLvMqDBo7isYloVvivokIH9HoMvCP2
pgO41Vjbpk6OEPSnqev/7xtfJzeeF/kY0mYpnQQXm+qhm6jnapWSFdfFdmfaHYWz
+olxaQ4FayV33F26k1ZawFWjLN/9H53jh6pCTolfBHXlslazX0iJRDv9vipvQktW
dwVQdjNgQwI36rk52lDN6ESpV+PL888kEsd3O4h2cYmg7u0kFqkbmNVjm4oiSx1b
`protect END_PROTECTED
