`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrOyNNgqHv2SgoDVo5U/k0e+3WmUxnzmHC9djCaWO/TCfPPQ/4Mh7zFgPCnVu/yM
ZiSQde08/i4fH9IgB8zhtdf9+iimxD4Zjb1udoBjMj0QLGXb091XzimWQqzIEE3k
DN2kveUgF7nTjKFZoT7ACiKkPs+otM+c4HNVin4mXad5zKJjfcjIJK62tvZ7ReiM
DGHwR4pl7kEwSXcGxIJO0LjFDi1q937x9gfFvkUb4Jyesr+PLnGGhtRg/V/ULPEs
CxZli6zkSpqL/zBiwzuqORIxgYm+fQPccVewWnkthRzCU2t4MlYC07qCRyJiXIvK
2/+aE1JTKnpDQjzVhsn7kkFaInGlSDW0uednXpHfzg7EUgOK7pNMLmNqOz7AdGYk
/8ttDGUmfzcLBDiZtvyIST4IQZ9+AW64n2KFB30C7LKhBkB01ah107DZV1QDX1as
805Iqm9TEOS50L/Ud2Jpzyi5thdq5mVKokRKitTG8TagaTRtxEOf0Sxew71J3vqO
pNzVVpYOS08rHO2IK0y+NrvEUg7azxGtAEi1sX18ycriPiECtUk9NJ9whz5pE1vQ
NGFuby0ncrSL+eWTFUYCVJaJC/Rd8JRPf5/n/6v/yHSfQCoi5eCplHjQkV1c61EO
ILEMv0CwGVtwgkhjCcU/TMviL41kgI0NfGmVI8h1rFnSPCXQbFJufS6l/IYmeZJK
JDPDRm2cluvy5Vq5uPiA7cDr5dLCMhVN5wvzd4WRvYa7Rhp1lqWCT5niiVzvX8Ju
bLkJlAjvJkIPiL3G8eTaJBaIlkjs0fyQ5LzyZLGfbcjQu4oTWMAIUePWpXQuEh9F
sYm3bBAAWpMo0BYCUDvncw3DgNhLZCtpKiVnHfGh+SZTW+yym5BchMNFRiJ9f5KA
o75orxdQg0Ti4vCmffFpVUOKBU8FTv00h1DZYDdGLAqxlQrIUwyc73fglEurLtAU
oBT/w9luVct+C0qriRbzNvXLZsM0qjMFh/My34T6Dh6BjkvbNB18KhvTwgeVEOED
/nTLNm4IdJhKjYmkg8QtZm+LJbkvZenkcw2QfBhNXMOy8Q1UDG0UkXHzJM2Jvaxm
C3nxvB1bNSGtgAPoSPO/Ij3ZJUHWGCIGkixJXY/bs9wseOA/4d+y1gxa6wQa5KjU
aoiQDtysfb+/8LDv4gBIW38LBILPDCO/eTT1Ys5dLsXWuCaGBespMn2C54AhQ248
9B0HCjgNBANlsgBeGCNRSOVH6zZzxME3uOQOD47rAtSt4m4W0i5BAtuJK0IX7ge1
0S2VReOeWBweT863u+DbSiqY9qNI0UMJjgRVoVGppIAwLCLTBZYlCavXtJ0UrYZx
JLSgegrOMkTAjIwE7YJmSwX08cxCtSdPEOPoYgu1krH6DDdBZVlkrw4bgTY8GklH
kj6IsPI59Y1o8cyKMv6q6WuQHKimoCI5Z375yVno9e9S1RxHb1zrxFB2kanA/2bU
QQsK7WVTa+97RvfInd2Rl7FTGMhC34qR7ndwTLitE+LImKwjmhvs7EZjpwyG/dpW
9i99EnCDCcysL8tX05XQugGJEX0iaUVZMj7P1z5sW2lDj2ormhAoJoFVWPabj1LD
9tudkk1+wOQyaPYglXI6wk/X6uBGtTKh6jPcr038uwW+UTD7qGJt0PfdHsVaZ5tT
1rhmmpn7qZoPjmksV8vY4IIwZr5Hsku91BXH5Z0cU1+ybwDaUv0If6jFuzeTm6qq
6XNomPke1Ytm2kJqRCZZb74IQBCtGxnQ21QMSVojm8HBTgNJjtBPnZLlOlmQafaT
QH6qc96IWpd9JPNwsfKLjS837tNWC5Xj772p9I/6GeGztEmbAgS2VeONtFSS/Yev
rI3JuTwQ+m7Ydg+17mQnnb+IgCIYkkrbi/odVfjD2QcgAATpR38oLuSgBwqW58Rx
uqOAgRMLMFFhVevusukvlYyCnTBpQ1wxDUoBXHqVUV5MJsQXwUl29+wG9/b3ISTl
9UY+5GmiHmZn7AqcWStGUs95vdhp09Qmd8Smf0CnkTMLbmKjTl9FGAM5qYC3vpt0
ASUBtZjNhaU+3qElXyir7L4QE/5zWLCE0VvOT/edZcdeG8s2QGLADGA1/S/xzRoa
G485OPRa6l0WL23MQBd6OWjiNGKV+Rw1rMH20U372ZnzPp8hIHm8QogV7bUa+tQL
Op9CXkRc786O0jHyey1uH6whyozPIsdu1ro2B3+CE+DZFzTeyerdTGqJIFYa0COj
ogaAKUMW2iG9MsT8l6h9ykRF36uzAq1+R+78oNK1rsPBZ5OIO9cmLo7GdXb4cS2u
HzY1hdTV8tszQb+OpyekhacgjOJGXaqzUYitgYGsSbr5HAaFCbdHLau1PVDsFDqa
KJWmqchGEpAxux8hF1Ti2RSKK0JdJbuKGByjQYg+FsUrrHZlWcqi8F9OuH42sFhV
lKVIKVmLA1DTcoMefd9jka4LNK334UbvUGiHydHLQjGmYLgm9zUqTYOKaSB7hvbO
sVWFm07IYGkLM24smplI6U0H+K3vRU07VLZP0G5qDvpQa6DZtAS6quWWid4of/eH
J9qxD0bAxUw0RS5MxV+RZ0UjloMGEPSNcIhmL8D13hPT+fiHuy1oviXtKz8GuWCq
TZe8Q7iOo5lm1GD5Xuqa2b9uNybPhDSy039nv+Ra4ynfVn3/yM7iWFLCQHr/i1NS
AEzQdPQ6NrTMV6x/t4zcUDUdzHoeBjC8/y7Zg7qN9iyE9c0HHbQXHU9TQNZojjgN
QSPTBHeYVbxylOuR1EJV4fJWgZjlL1Nr0HU5flNgehdSnD1Empokz0+AE8LcK3Up
AGFmYCm2SyQpGZ2uUCMLW5W3Wev47Urue2eQkyjJoG4KtpiKUyoSO0pAf0k+s6Rb
0OjlSsyWeXfDmHkEFyECd47EkXU4YwS1ex7w6Ja8dGM37eJDN5a0gBvjd0z72fLI
37FN7XHAhpnrSscUG7ZCdlcvXE01704E1vlwYp4omRsgFgeLUU1OTu2iUrSg01v1
TQDQzB4S9lEr4ShmsbiIw5keeq60PnF8DsYHl5CYrS+wETsz8Qu/1SPIXojPFGyj
IBARDrwPK9apBhNvkg7AgQNqWqkb+kUAdeXUUDmhiAyv715lND+Q4T1E2ONZZ3Jm
FqH03NAeGM1bIPOweg6dnjG2KXY9u5ca63dPV6vcGAAye6qhYxKK5vkMWsDLY9wL
d4DDs37+l29mApiiHmUCPWYjo/VHSLLPIP1WRCqgsK51UIg3FQC9EDQdEC1XeU3L
9wVLC2Xw1CaHsG2+rpAd0EMn8GLgAQSK6YWLbrCtP9wNGOaD+uRCz96tfuCHFVQ9
8GTbDESlXf9R4wtJVT/g6Cds1k6g7BXDMpTPs2ft4jrVhF+CjScBkOB2yKMrLeKp
sXNTKCumtbeSUKpHlrL5sUwStFFNx+sbbqRM7t6aZRD0oGv5pl8QmbCrpvf4o72E
KgBXesvXADbSNGWiDcv47Ihr202p4xcRtmnIF67pjXrin6jIVgwMt5RQ/7Gd6enC
DkzmplT1yoxb/udOldZxi+0EfRmrsSJ1xD7c2XyKKmkAlz+o+oTaepIua1X9VZ3O
gNz52zvG8YmOXeaA6ciO57be8L4ozLNkYRK7pD4uK1YTDj4hAbiPOCsr/e9ovY07
uyUF2QnB5Km3QO0nu+9K2iIg18MATcCALNTHBGfuAH7oABHlvdgxOajoMa6An1xP
FV/AqG239r9WDlqIVrWI2WZfnL69GAVGFmui9iQBuxRUZ+eznyHKY/3IL9n0qMdn
abKRexMJSSW+q5iHu/RC63aFC6bmuMcZfGPI8+fy8q3/RItYHtftoYW+EvUxXXMA
2EMqi1PqBhrrzhKY03nFU8cBSOGcFYTthFbPiF0Zoyg5i8gxkVjG+Rdk/Foqa8Vt
IQGmvOtfrsva52ssJdmz/hw1goaGJvAvOEBMYcIpq6BPuH/rLXbjy1gQ3mIlg9aU
J0pfqQcKD4R3FC/xP6hzPz2UgDy7dBaFUlB21a6SToayw4lHDsW7bplGbeaOcrNX
lkwY/s734Sqm5q2TXRLkjyALnibRwxYG+n7yNUKcYiUKJ7LcL1jUKZO1a/fmHT37
ncVez/q/k3n68OID+gfzYx+bFc4LvjPBwVQgn2R9Yreblgb+qkEZ+uf0OKXXPNhU
kD3aydVwTO2tlTihiAL4lIfhIqZNqYPGNc2Gbh/Jmp9VxZR0XkArutlVKzqljhMB
Xh/FrPByNZIu8HXkw1/AdEUy4WQwf90bHrFn7xlvRAVFI5IYWQtiLgbz+/0xKj/W
llMA6u4cd7TDTHA+ThIMeon4/JG3XxvnQIyMaj9o1ys6Qmg0DVJg0JWj+EyTvpvh
mPxs6YXaBmtPrimdJn/1hEFC6xzNMKtwtAlYQca3E1rZ4gDLt8VbHzILmh7+1IlO
IGqndD8WWfWF7dYFzH+dktA5JRLzBRy1N0rBqvZBNlygBmIEaACfcNvyYKrTWlCw
`protect END_PROTECTED
