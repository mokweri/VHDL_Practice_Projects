`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rVCQ+640P0RZRTMqkoJFwS9uLc0KILxb7IFYt9Qf38qe/ayIg+n3P35GhZ5U0QE+
llXM3KlNILZ/379/zYuPMH7G+DYirk3pscodE9lnettoI8u5xj6QEjrrpm76lobU
MWu2QnqTMnKSK6Lk9HVTBImgwsP0CvT1e6629oJ5jG4OiH2aTk1YwlzFqpK75ux7
SbS99hp5iCGHO20N+ChCnZmGAnym1rIaxjIBpRDZCdq4yHnWuuKMReWTRLBjev/M
c+Uk4/X7FPqfjb/8F6cSwLXLEElHTULeJhe1fp1s+vasGs2+Bq3fQtYlJZfnNpz9
7Rusxx68gp6/dWxtesLRMGHMMRyj+4HJxu1ozqBiRGsOVQ8cYM/WTzquXkUdMB8E
nY5P0xq9dEMPrC6mekqhMhHURhFEtqB6CWa8Nn2sie86ZKHYYZWkDEBU7/JimFDd
8RkCnvtMVd2s9kFswomwCSxz+S8bLrUzruQ653cviWDh4Vy/TSBFQKXhR9OKYolV
r9MOWqIe15jy9WA3pcvGFf8j3ifabtgtaIjx7d/75P8tSONwV7OPVGYEIQiGxGss
jsENXh2aJWjl501NuBSBtVH44CO6AXQRW7AU/1aL145TOyAWJdLgAy3xWC7dKflC
2Z/dni5gKl2T7zkFOYom8oAuLSdc5MiKHdB1bBldXCO5/leWNhY/52eSCzl7ns4e
MzGefhLslDU4/lflKIh9PG4E/2V8Qh8bl11F2EUOOAyOGe6j6tZSOeoSDgNtWRvy
AP1I73e+1RoLts2ePswPV1yZr7ijEgJSUCHDLB3Vfl2yywY/5PoPjRaU78O5zKHz
IqqUwIbXG5xepssa1EBuuk25qvrQStL285CuWc8xxlE=
`protect END_PROTECTED
