`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCeSxE6oxScwg0pIRMqvtN1vl8h65VR/+7RmvvOhFlwatwMysjPWk3Ohg66teQsd
+hUjZCaHor8ATom6OYI43sg68hsRXMxuFm9muYeLMFqaABnCAN13/Y1pzU72nEgG
oJzpJZHyaW3EWYxzCvvjFXx8lHhse4N3lJHMna8+AaACL0dLdPSs2TUZk0LxTIDT
Xz1wOJ6wIedtkVuIRilfgmoZoS//aTVq4GVD+A3HRcP+o85dFKdDzzhywzjWBhUO
yWP9vLXGk6KdE3t9dPSh1vBiveT73/ngdfUm6Cp1B6qCsAwMCQ/9sbv9OVOqG3UV
Q3V3chmkT4t6uA0T4YUnMddyu0nqaCGZhR8L0OCQiK7f2OttSMkjaQ/EClYKAaBL
SZRUsJ639BNYD1nWLX2KDHBQRat0YXFGQzUDhRvgWqShAqLyfio6MvKBcxEeJS4Q
uCqAUQMgRMpMkhjFvf8QaHEyu1GWO7o6IOyqcwyKgZmiK7Om/rWnzhHcmMOcDyA0
pQC6TNJMEs0+WRznlhyX8J4liHntX2egn0agIirBPCvqlboJyPGNVUGyUcSylcxX
dgsQTsNI+urhojze0fQ5jeCYIr/PaG4NrcE5Azi1ANGapO12Z9bzyraxQMfqNnBY
Wv/4hsBmTC8Bhqzvk58nE1VRMjNoWgnkwlL8f8mNlaQPL/1uXd4rM8cGs3Bw6rLc
aZAl2KnK37ujxytoVDnTEMve+Xz3Ebq/ISCoZDBECVF77mPeblMbAyH54paatDCU
CkECeP8iP6IHfHrOqiWHUmFDJjae6bYEgUoKZybsQx4Cblqij5nB0J790Ltd4x+5
Kl/Met9SDi1AO8fRiWoPgyeTPxlyk1uqEP+p7+GNKgne8MihcsUuJGM7vIK9LIRu
YuAO0QVf4/M7oUK3zbpDZ//JVUmHA7qwJ1OI+6DPVFJ2JBRFsK3OU5GqD2yxkDyd
dnDByAJ/5lLXYKP9ShRGllhBO/EZn3rEJbxBUWMzFeMRy+7bvQ+jnLjO7uzI0Yhz
8u3GN5yXXkIttlBvYXvcUQAbn8xG9OQp6jlsPtA4HI8jEiD0fcsYeFvLxZKu63eN
a9vJPJ6a3Y+DoehGIkrjjXtRUg71LSl2D7d+n9b9IvZdNtms5Lds0kaCr7lo+KJ1
+GtWUfhn2G6ldPaFge/R6GPlX5FANctdPSfTF8AuD1gg0dIPTHAwV7FQ/rvCDNq+
Q0C9MV215JAb0AXJMnGPGmpA/A4kHpPqEINV33kJw0aRMocSW5/pxgL+qce9oUdu
M6WmiSFxVQrfhberb6MHD9aWkAyol7Ap6nq+MR3VTRUWsrP89B5iS5tgGU2WcJye
+Lwt0l8rUJ+ZtaNazq7kR4LHDEgNWdxp+cTQ+ezE786QVdg2cx/gZsORHmvB3Oiq
1YjifE1WCAVKxOxmxc2UQrt1RzrxYTs76XG8typ10XLMsnNzBCfG/OQbvuyzgYeA
KcJ9N7WkTwUKHL8iys4Nk2Z60xspyzJyE/28ZhAfaFAFBTvelVDGkHx1wRxMIYzE
f9/MysSYFukvQywVTyB/+4jErqp/Pys3V8A8Lk5FXyyH18m0yCh6cGdLl0SuKqYB
Ls3ZN5dBwB8gVRe/oBfrGgzN0s5rLdhNqR/m8OALzZQg7lJzk7h54Y8a9UCj+eTF
rwCyTJ9xO8HmiEjgXwOXB77FABkDj6IZXhzquBjhKki4p+XvDf9nvtimDXafEgGS
ixgkhh0GDA3IiZJ1OYCGR376nzDX7ziojUNIlLmqCOI=
`protect END_PROTECTED
