`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxcFNC+R8u2MzQx4dhH91r65jlClwrytNTjtRzH6YtjHeXue7dxr/vEEgpSk0AuR
RWG0vQXIZGPThkVXv0XU3EVBmJXmzmt9fJ9S9RZMTagAX9mPPloczA/uDNs23aM0
wNJ553R6h6cOLiV1cbWMqFARo+I7iUmwapE4Fj+DTg/XltfW4Kai6izMtOq23gSu
AuaFI1nVZtiMOyYImTOf4pfyo+0r398oUxzIjt4dHRUV+dbWyZQy6673L2+hsYSS
cZfgTwHTVHqNnP6V/Kslr7rP5KjA2mRlddeucxXn5K9f4fuzvGGzK0B8EHsBUhbH
lDc5UBk/6Xb4r0ggD3xmT1GbpgTvqKOWyWQ8FAZiTHh+tm3186OusNDyT2ykHRFE
BKdDM1zPv5uBbWHQf0ilGoyhOYeqCgynV7lYVWlkG9svX2zR//iFyzHpb16c61zC
jDjdQIT4UbfUlX9S80l7/LTT6A2FF6zcnc10PeppwaQCuq1wh5MydLXrWcC0pLKf
G83qWIdfQUeYZTc8CT3FEoAwrjpMgeGyd+yu8KXOezZ0WO9XVNxY1fxHYzpZFxEQ
1k3csyJjfUWLdLQwpRvewALwucsohbRWav8gYl8dKjJwdmLRIx9OLD7yaiLUD3dK
Mhd8lHGh4aYO+P9/qri7jbtb0iR+pzOalxfvyTTdu75xD1tAVkFgb/ykxkeog9bI
ITVEP/xxqHViplNfFGgZHpGvZJnmUNDPOSiNhlM9f+L4G91pDopX/VMaeiaUQWQr
h2LGcCfEJXEo9/n4ybeSobFft8E99tqWNg2XlKGNzERsylBWfafrVZMQsW4mwmv/
0yOBSYotJomnBVUqAJSE2WETtZ7FuxLZorr44+wYljt0UDFrqecE5hPHNz20fzBz
793a96yNZ1AJW5vZVGGpL3SxarfDPtejrOPF+YAFr8UuDlvvgNTDFda3XJl+KRFI
x3obSVqSJDHuDyl5WIB0PuBZo3u0/KjehYiQEfSZkXfrzMU3qpVhmh3ArvpI1j2p
4Ky40hOR/X75ikQnc74LcAa18epgqicEUoFGRQ+lcAugAdN7uImvKfKa1OjKq8lM
WGvU0TNDpwXNigHSCFzLRsttPgGrOs11DzosLE6w70vwYn6eo1awNXrS/T6SrpOW
zJIZ3TrIU6ohgU5tECEMskYfheODqEML8KMB6fGiHEVbiUYrSYFZAIb8J67VX4HH
RvbaeRREXgKpbTD5NZyQhI9u7jgKHHTvIFYhwF9qV81vixBCz79i73toeFWanWHW
CbfM7xJ5AI4irkVponOVOItAFW9sUrhNbQycUutAL+G2nAPlNlZI/4RA2fwEcmLx
xev8mGZfFdWqnRtDHYncwfqYwOTIM3EoytSF5tC0tfSHEJ/FBEW+rY9VH71TfT8B
GNbvqMP+8rsGxDcsKXDxOf69Kuwi30aANpCoZWxOA/w93Oh+/hIkvYZxBd/gYqJI
YrwetZAnG1EMQT+H0bf93pH6QUy+q6eG6dG2qe0gEvZU1bZy8bDco6l/CMjHOVSC
Vt/uoi7jbMTPY1IuZjUKcFrpGn0RcAMn+HoqDV/KxdkV9Yh+3R3tZ1omrvVWgdGG
y3tvHIfVkKw+jF7pbGseBf/l8XDwnwQhuDF0kUwL5z3OAaEImyvAdXLWjstUO2hF
DBgVN5ZsLdaPmbkxI+NWS1SnMXYQcD0HWhZlTy4aEPCKzX7D34bfUlop1NkT4Uds
ooiFbKY5tT+ffCOvsud6Ew==
`protect END_PROTECTED
