`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gn2AKmqOZfI3m+GFIVY/4x9BA0uXq2a02pEqO++FQlU9thUdjJLwT+48I9yqedL2
C5G+wYfKj3fAC2NgSpFqywetq7PqebGcFMrlU2LaW7gsWRwlEbMrnRthjN75/YEC
uwUw1PUfOLDadIR8t10MFQIWl7epLRqKgVq5+D8o2znBssrFV2y2lc10uJIrDM4j
YOo8qeMB9x9rsPKx+ope8a0ZoGCEq2BlhF6onfVtvBnz8GXGsMIexEH7xnqW/XKk
rvjeeISPrTTtVMpKuCLJzfaKOLjfdhZFfG5NLPhIHacj5rlvKncBhsma7wxNJXl8
nh+7DIKAq0SkqRehbnHDcjbZS1ilotETB2rkxzx2sMK8Z7lSTWYcOIfVwiDt304V
8KTxH7WuAilpGuis/zHH5LB4qT2jH6XZqwlbSP3tZUr34yhpdBq7Uj9MeNsnI5sP
QateTRSkcTsZrXgZOu4BOqDJhs2Mt9aUCvgQ09vR8xh5VyuIxywnvKUrPbUgVUd8
TUnMtgEe0WaMZrVG4Y0In0RXo9JeRNLB3BxpBKJQUSdSEM5lFiikCTk3aRZ1EzT1
YHDpxQEw8IpeLcyJdR+zNUwBKquWDD5XA36JK4ucb7T2wH0O0qEzdr+HVPwj10iy
gHodnJvD2jlF+jvcK1CezYY9AoLyUMUqViZVq2l5UtqY5Fsv9WzH5EShxGhbqkdZ
P7H+Qc2wUGMKokgowrjREQ6E/Q/4bIYlKlUeerss0xie+3dUmDLIKAd/GiYZjFcb
rj6TiQWcS3++jzAt0wrb1+rqa9WekZvQO5pEf3UzNDXNMWF5gxumM0XNCYLh7gVA
mcErEw8sVmlmJdRvAFJmssZ04cixBq0u5qX7fGWNKnOs4fnKzscEhbljPqb4WZLZ
JwrBFxmGai0uDcsyuNBdTogokvv9RIp82NrwhD9tJoI+R97BofSky3mNi/Ok7lH7
bHr6mPXTeFKbukLOAeVlx7me63ZlHwS9lHxa7ORpWIgAD5W/d8m93c6XPm4Uz4XZ
XyvNwrXppYVeVLrfIaQlIQ5okcirVcV1PSofkfsamkFniQK7wEJ0UF6pZg4YM2/K
O4nfCwhYSGYNeZpCXBpXjBSESILzbLO38cj5Jg1YXy2YuU+TDqPJjgEjMVdtNutH
8forzGD5MWmZVd5IzZaMfkO64K6PfDW0M0VIItz3ILZh+0NuQIozQkQN6b7ueXsw
hT7YdZAFV4DYQXXAVPNdKCz7Lg4bKJTTQfJ0e+MtQZYiKJcnU0rso8Nt84UTBpYM
i+au/YyWCLwwFf7t7SbnngruOj737CzYpsIVAzUYTZ2LCoK7snUBFjNDvqnZBDXc
BSH9Bfg6oMDZ5bidyfsl54SbHPHTVF9GqlOQ0W06hZ04L3bUfb6x3P8XUXoAK8y9
Zz9FAWP5symgTnOxCMij6s4FVpeCztTNkkvQqAj/thB6RFi/EXc0XAyu9tMBGvst
LSYV4E5Y2/BOgeC9uhRIvO2Qz2XJRZzsfvdBE2+s9epUljER2DESc0CyY/h11dBK
GVmitGOlByZAR1t1b+/oBTNlRbw/0OWiJAcaclkCvSrbVqibnT5LDqzmFlssPHH+
1GqzAzBoCx2BOLewlhEhVM9O7ZLiFpvE4SUZAZRQ4xLfqSrrZ7VnG56xUsRuPUjt
vm3r/xCJLrkdiGmiIiAmgR1BXilhhegXi/1hm/Lj7+y9u2rY5bczsOVHk8NCrdy6
V5isWh18w25E5wCLSt387aRwegoy2LATI9/gZllXAVFzsHCY9MSjbi2haxMeqcNn
Uz59qA6kxqzRMOOAhwd0ERMDVRbcxQYEamY99mHqBc0C04qk/Mtf2WxsWghmgqmB
Ie3noK+NHgx7vmAEO4zPiXsPAQh6HPyLrnYCqk4VpGW69ufthK/xn4ysgMzrRkKd
Q04aEn6cu39RS/g0RPYia06Y6itizecCWp1r1O+4RTpXcmBkoEf+94D4Py3qrai6
idGWZFkOhRYspTUKlP6kGsbGHkziN8lGNBRioZZHRBgP3fqNX4Z3a1LTu+5fYI3c
ccCKqnZYhJP5iSyjPZWQDzEYOGcRk/4Q62jWspY8RPvn5BkxdREKi5tOPaihmXbX
O0NXKAIhk0s0Ow4CHy7oP/1SBF2aL6jgrfBNB9qLx85dfbrBHHXZI5CTKgTHn7JA
UHCxLMgRn+y+3bZUu6biHSqW258W7qliq5G6Dosr1k9TE2utAPsNrkrtjW2dzMze
X+NE7EzfRB49IjbSeGLEXZQu67StI8tRdrzbGTD9V/rIjE/kXUQWeo3p8BQV5bvs
5CK4CeFfW87hl/+bQ7exrVXnrHKijugpl+9GtgjHLszsbhDMgCle2UOZvT3TZDs8
Y8UKOkY3P52eTTagmEmd1BLC6MOEoJ83vcodL088bSRDlhab7rTsCbd0+hm3yXfP
i8mfbC1TR3p6lLBsoJWvGnDsWaBpieV2jdmMHUlegDU3V1/YUGLZtQw7xTjmQ0Rt
IRa0JEJLsoo8swKUbDbTQbX0ljlUzl9udlrVgrPNSLd7fUhSV2m43z6yLEVqxul5
sL2sxaa+j0qIRn/vMK6GeWcRb8GQSmo3x1KIj5QDnYvcDa64zQ689vcRYrxckkIY
FIilalG4sXeOJvzsgzD8u1MvqoLXTfs/GhfSBQhW9Jt7hAWaZD8DIFlXgDcka83B
56V6LUTnbSUmmsjsvK2Bf6XkMQPRqidHHOYEmYAtgiFZAsWdTsJBDcAA28+uK6SO
aDt1Cfv5LDvK3vDkhPaHqGZb80EZH03WVo/AxCUJ3HhR/IrB+wPL7lnh3Kkh4C5u
Jeq1/3xZSZFsodM2ZlQn45xMjkMAk8gdt2v9Ls6C3KB82Q0twVo2SgLEd4FRR0db
HxzKoBUESzzM8avYHUTG85kGW+6d7vXTXuOrIfN4Nu7ZlDq9QwuekWvVKufgqEgk
JlgwGElI7A7i2Pi+Y9QstooxYjvdMt/fZKTg/pMzDgntp3qAHu4aq5O5aY+n5AxM
P3EixAvRkAb5C4voU0vQbBwe/cukwSIlsYCRDSlNidVdyNaMLJ+Wau+UJQVaCFfD
aBiNBlrmqLEjDRVkBVrjx1Colnc2jVfBaV8Lo4XEywj3/IbOjVCDiFML2b8rc40+
yI4+PmBWpHVJUrijCPh3GmE7RI8vkG2L3y7xVoxgU0Yc6rhbMcSngyE6ehxsfVLk
NSM2wbzF0xBFSPS4Rw6owTpGJezFoMzyyBOTlSVwKKlssRW8nXna69CLtSlxR4nl
b2bzl31keHaIFigXuzrRS3cWCwcc3vCUoxeZt8Dr9Hhd+YSRCpItJ3spihVJJoYt
9q+r5wWO1S2DtVcwgdSixefgdPbu/EeicldL6RIGbQ9QBWFKcTfDGMd+mVIDi/dS
FCcXwNYn3fDrd0IlDnVdTKwttjz0BMEcvfRCagXCeFCPkQIIQtJ66EinVMY39DJ5
lvn6qN0DjrK6/gjmnkEMHXzUYPPCvQOMCdlGSiOx4o/RdchTWqecFyuiulr57cSM
M9vBuH2am4CVzCveLnIFiMmtQCz8oFwWOf/NcYXPtIaB34xKrD8dzh5Ny/QNgKm2
IuKs8k8n94h8yYPRyvXrFHMrSxwVWKAAuN2YJODKOyYLL4d9mmfULXvk7eHWeLkl
qdimEQMg2x7ogc4/xGgZ7iXVhBb9aH7zsDdMqONas9r07aDNwq4jb+5PdVWyzYRZ
xuBHiR8nywTPfNaF8VreuDC1q9JAulh9AC5NWlYSr+BY+OBgj1C1bUjI9oF6+MN7
9O6+vpWpvq6En9XQde3qkGfHi0nwhcZ8pdZ+TXzflS5KoDzZDDPCHjgM+f92ilCJ
/zWfGg7049KLW//M3/AIoQpPM1DAaqcLX/q5URFGQLjurxFq6s1lvNK13+NTPeIn
5udD0x9xfVu2shwY8vnm1KOH/VtA13nyIQKYjyo8jR/H9UGhkfDFmw+aejBJ8jmF
ppXgwqJ8zpLSlTMAV7JCuHb1uOoJyKUEvq9ekcPbooPxXjUNGShHC9Ui80DrqE9s
hSCPeoyXdmLxpG0Ylv5zpaqehXaOrA8H/2Ak8/dIYCfj0YlkomuYPWXV9MZCQQGc
Hqsk7Ul/X57Ng8oZ3diqubEV8pLn4NV2UfhnVfTPzSqsJEb9M4GVMiMSQAe/d167
P6yb6aP2wJhZZqxhRJAy5aTS+grDw+ggAcMYo3Yhx9LZGXJfuKbRJyI5yUHKk5ty
W/WK6fWU++zPIUVJrrtNx8tNikRZxZaTyIDKM9wKN4K+9PmL0oBgZbrVBmFIzuKi
DlRQaZNgL1w614S4Z6VPR7VlfW45A73iZlrK/kfFF+omzrxkmxP/Bp6bphEBSAEH
MN3FSXDm5gYRGV2SEOR6qlIJpPXy6nZOYEIsE9Q9C8RjQTG11w7BAff3WYZfJTHO
lTpbmg5nLc23HXkzIffUwExhRJuxV4bf0hnGvYFPf97KV92TJrc9vfDMsfZ4/zUG
1KDIxb1maqLKPuBL10jxWT8Y0Vz5HEZHyDU+HFlXa0eVqLqnczJ5xltdh3P0MAbw
xWRaevM0y/8F+SW7RJdhuI3P94oE4gX0y76lDkuvz/pWoxJ6kWemmTtkmUJY5rF+
cV4KkW0m6Dv/8MHTe8S6FGOwF8Z/SveJucXREMWxZO4niMucJ3+rR1L2k6QE9xsa
hneRHyOB4VMj7n1X2840QGrQJZHYKGZkqOsjl85ezzIxvjjDuAhn20OMs8VCKM93
3tNPlsyI+aWThgyBpAo8LMujR0auMuIuHvlLhoVSU4gul3mVdYlO3ifwrZHdmVm3
dMBTslg4dO6jf2wExy/r+kzk1yTbbP4GnRft3SYHelMzffR0vl/m9cDQHyduddI5
q7rI6XaFV2EU8EtalA8WVBKL6pBpRq3xSJI39pxr/sPDa0x2o4K8uM4gC0jQ72q0
FgIpHp8gEwYYJECOztNEuzXuthxJgwHEixoKDy5uIQkkkfhwS2qK9B8DaZmojgsL
czWXrp+OhfEC8WwypHXpJJXCiF+7g/XUqzMuBmpL1Uu/yxt6Xh1WlzDTKMGHu694
Cz+HTmvgzpAy3X82pa6b8YVGbPncrOunFW3YzqGWf7joBLCtONnfSk19C0/EKSzQ
0uqJOKxOSXGqJmQaXQ7VFLeI+hQuqZ6LngUuLPLo0YmkcdS+E2jG2/UatleKJOJo
+O8NGI5F188amYKZsU38/uL+KNwu32iLPNyRrKDhMOOAKkVxJIiZLb4J6DepfGK2
p8C7r8RBy30JaJzWjMnd+3tCG7XiASpuaFQ10RyWnFS/aT98xQ7IO13SuS2kdtDl
iIgGSEwrh4GR7HJyTGBmaq7e+c5+k7Znsbl/y1C1L5RcgJhLlxjcquh4NjPyb24L
Ge/VnWgpZe6re57RRV2mdY3P97UEzHdXHsQsur+MbdRpjRsGfVoup+3bJZuBDyaA
ArbdqjstNaMAcxxdAh7fkA==
`protect END_PROTECTED
