`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDqO1ALcNXBqTyUcP+yLvFJOMpwI6N3exBftD/+6ccUeMGQyz2ee1FDGxBp3VvLi
JggfZM8JbtIYrRYPZGtz636Jgc0r1nehTNoYbM+P1qPJuI6kjEPpud4eE/CZ90aO
NEFqWf5AQ3pVms7E90I41SPx3PkwXMf6LLMWWt24GZyH6tfsUsXap5Wd+gACk5dV
WRNmQUgH5PnA5PKRUyx9Kq2yzV6zJBkAG3SeLE/FBaUaLKug8prLwabTp+TJY6GD
5yBuZxEuQdH2Ea55i9P3RhoZVwReyOUB2yZO4iWeh/GjTI/qcaikLEPLSel9XE65
xRfKKav9bPcJibDEQ0Er21fwo6ZrR7WRvKqXenYLMUY/rL6mLkrWpFSpJJolsYlD
JasAmqVPhmyZwVLXjw3hiByztHvOcO5WvhUmNgLMs1njLjEuWRK8mmDQDkRKirFf
kx/x52dX3VRjzVPM0TdLGI37jbZxkJ4klWqCXkXua1a0wU5IRiK/c2QgXXsCKZ/v
nEa+Mwuon0ns47sYCFQUyXDSyab5fXDS83NKUnuTbAjJeAmIbHOxb38479ONVAM5
+2stnuOzkEKPd43Gob+sFq/bWbM5NIYENjQAuEo55kzkBbgDlEV/TLTr07LeYpVU
ladde7/nnnA+jYxOR13NcHxgFc8Yxo+xzj1ioiPv09G4DfR7AXiZSZizxo11Wvso
Du6Sq39un6FJW8L7lbLpQ3DrxlCq6FAaEvie9+bKkDEBLPDRvcBv/uPz6aqECQXu
crJ5rOMFRhfKhrbfJeF5qOizKuAN7k1jvLgsuMdfuZ5ZCdEN7DNDPcnzjVAojE5j
SbEuPxiHKNGekr3dH5q0bSjBYiwEYrilqXvbUXUcDTijcIQZvxV1Mb+IainhUT4w
GsSlKz1ouoCF8wmO+PMJNKjTZ5O/Z1TJXYgcHbAAQrKQ9qnD4ECd5w9k+lOyi5F+
XIvoMKnIJbowzae/XKgsLkKicJKTFTcXDvISjGdckXDJqtR2MvXkRIKQKTvsnBam
NhZEPwjhF7MC+AtWpqUy9nNdXBUjcyztl/MsZMPDzWIVHVA+GpvvUHlXoyswvXPY
1Fo3N3maQwHu5We1rjvvqA1vB0INA9i2geN4ZtaFHYMgJC3xHRrDGFC3w90bqQnd
Gy9+IY+FJO545h7GdQelwN9a//etGDgCbuW42D+rZj+JBuy581F1Rb5wecFDdzze
yqlm7331QYDcyrv9WH/SOqibUGxNtJBuPFlv42rnhFMG9Bbg/92hL83QM1HEw2m7
+dAZV3qVSu4OShf0inesA20BrHIYqnIYl+Hqfq5aGVbgI5QzWpyXyLUHadbZprRP
f25BpPsoriqqh3ZvrC2ZmzwplrHs6bZB3W9c0UjFyT2f8ZeSa+WAE5srA70Dsitz
3+nFktSAgGA6HFajhtXq2f8eC28iM6sGG+tXOwJDoSyJ71rBYo1zqLvpsZ3xhR+U
Gfdcq0oh7KNYwxHZGxKKv+7G8aREh3EC1j6OKHdiN7w8XSGZEanaLiuzsE4rCtOv
bs+l9+aJ56kSufBQwXe79S+4l+gj78RmZ3osB1YpYc6kYmL7DHQUPdBfg3My7++3
/pC5YMKSGjSbYseJtqbmf4JvVI89a87E9zi48MTGtZJ1d/v0E0eV7evokda5w866
crKEq4HGTMqNTksgFgVyx8L6WljiTDv4KVMPI5r2dtLgpsagLvJuPbc9lVPcPTlq
+do1Uni6qi1l6297rC51pIX5g2U29hgQSyFeOhw4Qh+k28be7iUwGhlt+It4K5TG
RnEKeal86583YzmR76ZdpyGBL9zf8JPy/mWB2d0sX7e7k5cDzy++SOTBalgmV592
XK14OOe3ofYca3T0G4ZOR7DU7OUs0Q+46z6K/b4LCS8FiCVz6+e6+7XGg8BA6o8r
8ZLPp789bKDWeVg8dOPkrSXxygcuDtLINdRExqe61SrV9A0aboxGFcwV8kcQdCN4
honTLVuCVm1a6BPLLnki7LdBoEYvoW0khXqaGHhf5QdhIT4aAAT/NJuTw4VpzMr3
BC1jAYxPSDu/zSrNkguJu5zgIT+rjrEkuQT+60Mkn62CmBsETKy8E4o7CoWBHUTF
Yt/al826EC0g3nSqG+1rBb0hhh6TzazjFmhne2cnmfuRXOCFQM5kqoCc1+hi6tEB
DNZDXecNibz7CYQtNLhYNrASg0/Wu2aqIs9LA6qz8dzpH3qmC7c5s9Hw+RoKjJMF
Z3j0NVGNIFzM9w/wMkW5+9nkB8sC3BDfJhXdvNhi8jV/rpCchSKj0M1T9ASJcH6V
2NmzJluGtsj0ctoaLk31L9vEImWWnuTaaAj5dry+0Owntpk/wKP9YyN6Z0aGA5c2
Is8PL8DvTOwNxIpLj47UigjnTKaZ2gGrWjhEVHPPll1IB+CGpLV58ERvBmyCoZvn
1cWXf26UBTguKvfXGBDRD04la2B2D/hEl5c+DXr6ohFNYvLsDmh5JW2QlsLu8dEz
GHOi4/ISDfcYgr7yqPSRwCUbchhr3ysRTfIRbZmYNLrl61GOh/dZO5xvi7IA6lMo
9IA7G3YB3PGS4COp4su9unMdgqszs2fOr1KGNsl908UnOAuukTnF9fRPBT7nVXyN
ScY080Xm2oPs0AjO18R8kHWHLXVCsW2cGvstvbEefRB7Z2/2ntQNuyLqXQvUBWN/
VnSyl1g8lcgD8VFUsN/Wo1T1cd7wKCeiWAbLlmD8Gc/P7kezuKSRanPEIbPCd0zQ
kmNCKWx1lzpm3UDu3V2nsoVKzEkrDGnBgJkkniXISJOkJChr19f2ET7uZimTOc4m
s/fZbLffQ62KEtbEH+1rAKeQ+5nl24RTzTFEqkHD0Pbll7p4KS/G5CRTyUGtlqG2
GpcXK09KIHASSz3CepB0xZTeTYIKWHxr/bRmoB4vVweFrL1M5QY3zqZLP45HJiLg
ocJDMWS0JAGMZvdJkldYOFXJdc0N8Wvf6fJRfvlYQD7Mnh7+l6N3j1lH4bxfaFn1
flQgSMKXrI2WjGYETlrFVCuvpqoVOwpS8Kfh60wWLXuptTxiGVkzW8BfDUSL8E5i
FZqjPOiQ8WIs7Vw8jshXvN8muTnS2UhsCjWGz7EiFm3xsU/uzRmZyT+bAwTJVO/r
q+EetsNkTLg/xJUiASrtczHxwRpkPN8kfHdvYyRAdeL4q4p6tfiU3R7POK/EhgP6
Gl5yIcZIQC4SOXawsyqb4PZM0z+cAUXdiCNstbIBnjC8drIpqwkemPN3SiPjiRZY
Gpqdx8Lmj/QzUkd6cXT6jc0/KVB9AryC8rEwS/e13Iz9FeqKSq7i4qsOG2FdfmOF
9jNmfz4Sa9Rtbdy22Lz65lUex3VqajFQFDqsKaKzkv/YRhVX1IRM3ghjo3YseXyv
3/WVQSrO2170Il0+r8ZJi0lMi62atdr1GZ3+gIPidsn3gTYuBRhy9O0ud1xugJTO
h7Tp0tLI2IfbRYdtg6SuZq2fyHoghZ+tSBx4L0OMGoKCGDHwBMOg5FnelcdKMzZy
nj7BcO9SFYdrAgeFA47dw9/L5I/4Po1Em8Lu29tm1IekAQW4w/y3cNSO/5dppbEn
oS2/FxdM5lqkUkWUiUx60pyObjFuDuXVHN/CxKORepyQykCSVhxEw9DeNxTtFKdM
QUNFh+BFa2agMVoROHy7lxg7o9CV4hIgS2eYqEu5N0HZ1lgoQChFgrc3fFMq35ky
yJxYRQZvePNnoKwrviyclTqBM64F8qOtlZMaxTagqd2BK8Mo96jZYjCDDZyT0exy
EtQ5/Vpf7HU7pvQ/z+iJOQD2HJKzBZelgwBD55gFiZYLWzPl06orw839Xd3G71LC
+YICupVawIeD3SGRb2PZ0XoVL6xX8OcGoyqCt3+C+SxZG3+L1cgPWG5NIWZaIc/v
SDaRG26vS3G3mKrK3FhVyemKmrsjBCy96090jxrBT7h0T7dYDN5QkltcrXOoTZRi
gP/quKAzwMQ31/pOq1HGG5500gng47vS6+567NDBQfBZhTBBju/L7bwvpmz8cPmX
SwAXnk+dtfLynaItxGT8rysv/B8j+muWVbfpONraOj4zMd9YU1zn15cfNeAG8UCJ
1D/Des7sjvjJqTr8UZp06UpyBAxuBExpwK/CWwtLO2+shHB4Bmk42HtSfq8Z9/AA
GFe6n2iqnl34IIZasY+Z2lu/nI3EqrFw5IEOcQAyeeIb9JYZTWXPGU7E78ftHSZc
bkaYssE4n/101jMRREvApr1ZGitkcs/CNqrPTAOsfVzkJCg/BIPzEDpJxGSd53N0
CJKKCbFurGTKNZCg5VTADyByQbt6T36oQXMxKHAAE1hKVFXNUM2kckNCsZkEr79X
n87nJyp6ADEsOwcq56biYaaD5ePXkXwe3JE+IepiTbOrMQgTqSBi1CE6nG0o7Rq4
GmvY+87/ej8GdJzCsQqCh4n2ynrIEEexVi2oO4Uj7jXOOPiB/etSy/eSisW49KWB
2ROCWwex4I2T6rtiMarpmFOuzpOiAn/wifGFpSbaEzAHkVHEFsZ9oXt8WmYeAl4I
AKNyCIXX2Kejn5DT9VDhdnqnawO4XjRVqL5FqLHOtCpxJkwdcFdrKtu1jXnW3/ZQ
PzAyq2z0Gdug+aGAXa5kGl9TCKIhCg2gqtoGLf9DIhIL3ZYLtiYukRoitwcoAXCV
pkz1366xTSR2gaUzf+IhmSkR+mMdz8KZnMZ8bweyUKqF6apdZ/FrDZ6DtvHlq+Zy
nUdit2Gc3V94RdVedWTIRKPu9HoKPHngjDryDQQokkJYBFyNIq4NhsIPPK2bA31d
lRC+h9Xq/8zuKD/JVKt0wSc5MyTVhN+trLRs1j92sjG7srMsspXy4o8Qq2bdhGBv
E24e6WvNC2CAbxdcYp6IJH0/MqniVBiZdypTEoj7DtTOpl+GZfmBb8BFn1/gcdbl
ArZTQ5a/Fhs2MpNHoH/v2CjRPDs8SlKJcOV8jykqxoDifP6fZVLWojxEuVxwJ9is
Bg61rt13VBFT9DmHexvk6zQ/lrkY1Xi3xHA8mIKbWfgFFcwGvXxMlCLU9OWAfOba
Orx9z6s5WdTcKidXc4rxv7xNkO0BADUp4Jxao7/HFNMEKdIxxEYuybAMGbF2sYC1
9FXawxMKcKo8B2yHDOrXHmGqyDEoFsny9h+qqiCM/CEcJgqzNmpFepGUVgY771bS
E4rK9j0NfmSuvkpT+mp8jInm1kVYLAPM2DraELIzQxbQ8IZKKsGsa1vL5yN+XLdD
gJLphqopOJKc9JE5ExeHk3LiebYfri2U1OHGcAip0s2cpBSlcs63mC4w+n/+ZeVe
/PEERPO4MRDGxCcRmnzq0Ez+xhEdavVoAraawl11Ar9TPoJOgLyL0d2p2Hxd/unw
gW4F84QHHzjca5MxvKG0ki0xktbuDvaPo63HI97+n5g+BA1yWJpsejl4+pQGGzku
M8WoDsxwd0cQ07wOAa6/80QWa6yO2/TS8Kb/HttSOUVrWXexEkLmq5esPQMJDPw+
n+R9k80SQ0dV1VirSi2PaXPqk0nJVfcMjO3AmKjV72vBv9mnJvOMm9VAr24LCoBQ
ZNg4XSQeQJN3rBRxELLTLE5D+S7nV8Ew6I+VvDVQQv7BK39y8qv6wgvOiJ5MyKXb
a6JFnvYHW2RoTCU/gG5Yaf4c96n/XA8q8Yc/17daVl+kZB83YdU4MmIO+9aqa9SP
EjAtex0U5O33rijMJoJoDTAabQcMXQ9bxzCWfTSNTnImh2BjkPho0JiqNQ+qZxXq
6N2ic2hyAZAIjfbdcu9RZdYPltbva99CS/itsjatdIki2wGcxcEVF+JwB/k7B5qC
2nsCM4qPqysQIRxP0peVeiaC/2FablJKS752e3fpf6ZaSTeZlyvj6MUYpqkycPU7
fCHSD/Lh6gKOyjxXH8mvGctXzJ0CeLnwVHitnszMPADqBpDiqoylcjDVeb2USgH+
z3EEkRlP5ZdPJ6AY9PjRcQR/HAPy5xXC7nVoj9tmMOdG4q8LM9+xuWc1byg80WK8
9IizLuLVhfV1l7YcVXjDi2FnmM+/xb0une5Bvk6Xo8dE2Cwc63gTzhHfl0N3IjTl
+M4RXIfm+ZS9zr9AsB+FjxjRSx3RIADVhsrWQoOC7EiXshr4hskRfBt577IL//GY
KdGmFoFLQ++O6icg0xxE7N02zm0rfNdtQ38MJSaklnLj/ZUok5Y8q1UyvB3+KQ/6
af4Ozw36Xtj3ZMtU5xwOJ1vj7LkbW37e3x38Ez7kT24bvD3h/p8Lad6JkSdxz6Vt
sJPlvJx6A39cleH8GJ2ybdZTessV/ZhO/ShLzxfwumfextAUy9NMvmzUKwQyjZAE
kQ8lWJzLETTcMWQYQxZ2tCxaVG+IPiurRVh//SI41p9R5yyQY9VMCO6aGoDcSXxX
wEh8xS+vU5zXAxTEKIVRKVgFiw9D2m4+T6QIX6wQzd94zqNAw4GMDRgeQEtTqD0t
XR05lYptay0dgrm2pOjXQjhMPdCtW+0r8XUrHXVikpPcPs2bTu50kz4UU9NBpOlv
kx5jbQq6ia2tt/sYi0tA+vY9QmhBNhiKW1+AX6yMJgm1iH0du4BDuo1PAYqJZFZ6
Agumz2SqBJvGxgQqs8UutQmSu2X0JE7Om2CtstXn99w2bTms3j2WiNg4X8cyFkx8
DIwQfLnqueTS3dHW4M0HfZhmz1PUElv+8nh89BYeTeIb6LZZKxLGHhpNuzbhKXxo
w/nC1/Y6ydCGh89RXM8P+Gp0HGe4Y6JRGRoEigtFCdtYjugEF9ut7ipDRJ+tKTRb
+lV0aIzq8ulOvi4YZ+POpqSwijhY4jONRf8P3kGSCCswMDqjdSQassR/LpfLSOLf
qRPU3W6iDbxhBVYupr8SLAnQb0csuKQLmar1xp9dn0I7QQ4Mii5N/8bF9G7MgABz
AnhvpfZ4DoBW5xnbVqAnUh827tN0gEYybjv8kqppgqIQI6JkO2xus+/cPPWt+QVH
wQK4tQdr+GKb+IQxAIBv1QQoZ0Aw17GDa5C04ZonkwwX+PrjsR8Ty1PYtYTyNMDb
AiZEUBBD15uj+G8hPyIlnBXpbznSFFnibJnE75g6T0coPNCi0lOXEhIjR7ZaKoDg
feOLhHNdMGCHuqv90TuDoH105fmhEg6dVm7wsrBWN5oFpulRMLcj7TtWf/Fel+3T
Db9JaH3n4pveY0jQHG4MRPsLEXIyk7yV5Ldv5/XlQ/tGcyyZdysjPwMOWbQsdxQ3
EtQdbDiCeMgrxXuH0AjNUlluzV0LuM2k7uFe2dJM/xPd/nPV7rvdEfz3Oz2eum3F
YtDvzsuBUDI5hH7CpmP/U/r99OLARpPT8cLDK5meQAf335+BzQow8tDHNEceo1dt
NtVQm50/2Xvu30aRC24A1U3oUIqXbPRQazHV/viRAR3l/VrK45LYCR9nE085AA65
XDMsGMiie7Z5DDo0Axp7+UP8N9gltkMtMmDnTpveGAor+esjfn+o6xF4uU05Wz+v
BihhDr5quTD/IqjlNa2Y+y4NWsfKOzUQY/QutmkCt2YYTwlymASGxLmzA8wHtPsH
eZKV8izDH+jC5OO58bkcQ81Z/iZN5jQSPqD58thki/KkD57Ru30ppq30lRwQyJg0
dhu82Ty3FRgS6YoxBEo59uMQoM74xIYT+xT+ySQkeugwnycLV11XctyzmVZbcfEb
DWL7c9nuZHGrRoLmJF7/+OlGkU3xv2T+uGA23kuoZVjwu9GpzKMhp65qMUQcMo4D
bBHdJpK0QezxXBFRbGFMPncUMSJ/yx+ROTDxNsIaYjhDr1gPORBNuomLuNP92+m7
E7ZHM/+bsIOTgy5mJGegC99QaEQ2n3ba+SDTAfCXOtuwEd68IvS0yonHtyyYXoFC
7JdOOgAAOi40LF8/I3aBzmyRzAjf1IvhsVCzqsxgb+w8xutxHTuYCY7AUwBd5Z28
rDEe1bCcUDXDlHfvl5uXh8lYxwjjqxM/+44Ai31XhUzIT+buJ3QpTPvPnUJSjEOC
KIeSahxSt1RQg/Ho8a/21QMF+CWcYL9HrBs0LxP6wDX4fTmM23MPoD9i/ZkiEOQK
bGDh5iDPdxwD/hb/8nUARsYwlDYZK+ffNrEUrBa1VUJilp41WkutnXOI4u/Zncbd
i57HIYxxUchSt9dhCB5ewdXxDP2/lWLN+esk0vuWz8IHAwOH3I0TuWHL93Tdp8Yc
cseiJkNV2nu+IwmdjzaWxVVqZ8VCWIlMJNToZjJvv5x49QVVC7IcN/4r+mELs6z1
jTvL5NeTc6QUyG+JlxQeg0lXC9UM3Va5gaQein+icQX7+wcanXbQCqtv2SxEpCYo
sgJA1aMgOVDFBMn2LMAycVwFu7JYJ3y+p0tvr1KbLBNS0dzBsgkOQYkXvpMqMWm4
RDP3/ZSFP2gae51acdcCVINSf6vbXfn/fxuGLvSEeeXTlDgNRPoqAkC8BPrM3w28
Gf4oTf4B8RibMrbf7LPrt/3Rtv9r3KkXEdLfxW1uGCTM6tQrip3L4eyWzPZOrWwZ
T5ZtAPYzs/LsphdyIVDh81/IOCVlKq0LgVyP/ZnUrhbQQJWWwiJXuF/CfintYxLu
JpMAVu0feX1fZSkLbNV6NsubWpfd3NopkpT+At/bXxzIOHw8e0RQQjMiDIvXWwQJ
RQkiWkRGZb52aDzj/KtHXGstJixmPbIROsHYFIW2y3Or1RzB9N4RZShcdrxMHdwS
8PQH64dExPbCUSK0X+prwXWmBTtFf705ZMEz9vAjvhtYF64xpKTQvBiJeu0NL9dI
KPa1v+0tRSyCv9Bhqnx+UN2LIlC7XzKbYb/o55qcSZfSwWtinYlkL3uobZCwYPY9
4kdufE8xpCz7zJcEMSCkhLdaC8YYMD5WDiHypFJm9tYghsQ2KVI/LAJZElV7g4nA
7i0x6BqBhXHXtwGrG/C/2vNb8Wcjw4KinGgU1m5XFVDnHI0We2fumcBkVTstseR9
eIca2/aYerVP9wmyOIC0CLivFgCIOGNnAdRlqPSSAqDpot3gVRbWSeIeZ6yxOQw/
TzKV5LAvmuFCWvAWFWcdom24IYBjTXeIEjngrWEVmLGzDNN6shIk5Kd1bZipyjF5
jIxu07VHapfdOCi6MySJYrqDk7D5ebTOB+jVFugp9lwI6raRPCdRt3Kv+r6G2Lh5
52avTqPnmebdDc78VRjp/Dz/Y9dRh8nldY18tRGsKJUxgFTmd+5zUsh1ZGfEaEVd
/+HIP34mv28e8Sz18PbrP5F/X9AdxIsMrYd3LwRahWv3kWgIRXLbHopVBfg2pD5W
Rd/KjlVjE/UdsIAQ8lMrNDaJHb8d/ZxdbhHaRTMTik25BnqpWacriJWeiPUqgm8C
2ZU3fBVw27Ivj5Trdo7yL297ajkEfmjtloIYAKGIMP/R9paLxBXeGmMD8q00t/VR
JELkuqrfJLV9TPzT486+h3wck3GMQ70lenLO6ovexgINa/h2SlyMI/IwZhDbSbPd
vIbchA1KzTjeKEFM09cFIQ==
`protect END_PROTECTED
