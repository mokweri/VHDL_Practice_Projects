`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrDq+Fv4lWyKx9izvg6LENwaV0099bgIaMRTPTk2qIHZK31WbXL9zYJhpmZU5ZkQ
ZMv7/baKlpqTLCqFGCT17h63o9i9Hl3GsLTi3kou51v8r8rzk3HR6LWi1yf7WquU
qYSVPFgmmHzD9DKnzFQGqOdQD8qOKWXcTyv6OXw2IiFuPZRK/q97Af9tV72EuYO1
0u77ZGpfhCEDW7MbrIYYmAB5fxOQfHG3RuhiEiTjXURJ4xDNbuzbQ3jG7UePY23L
S5XB/o/1o80Uvv2/Pp4C+rqPUSxUo/+tL4zRJ/+4yV+fiQuU44mgJYrK5hLS/6lQ
Ity62tDkDCaThQWhDfOh1Y3HxTWEPzi1ZeIZrfdPdNjEgJEAgwZhc+5XYTcjjBMw
fQDAo6sek990HZLTwo6Xm+tC90V7H1IrN+95iswGHyS1vcEn/qF9e74lvwUn+bq/
kPHts2mRdTL87dFFTPtFVMFahJeKVpLkO6wGo1JjKHd9fub3yvrCiNWX5Y9CeRQc
qeyLdoaJyPuN93Gu7y+FlEfL8G0EQ3qzjvvDma2sqvdz0RkhL18jPJh25+tBc/f0
4wt6Xkte7IApDG9vl797mop1wFObRuEQwl2UXp1i3Z/w/B0AjYZ+jrZsoTVobmwz
nx7qiH5VErH2VAah8pPfBGZxoFEZvENlHbIgqt/ZgEK9A20YdsFysYANZpxB5/I8
OzZpsMbe5vq/iYqhE4mkdy1kSkFTL//Oy0MsU68OY1BRlXl7XB7lBypi+/CsFXze
yL60dLHyJkOnvO/1ec4TAipmc5gq/IEFKiT3NfvhtqMRkn2o22c0UiDpOcaJ8oSX
Ejn9UhU+oPWSmMCrmu7rSNdn9ruZV1gLWuhXixcm9MnX/oyEGKqGUNqaV+b0SD99
M+UUaY1g0LlFV7SZvz6Mi8xErbWZIBeQWISkLaGnilGEJlPGucvaBYdctrc3jq0R
kT1Q9xpF2HEMBB4MOfib4uFtRM2Zyo3j4fwzY2z1bO1ZNIGl1kEhzfI2VO6VYvny
aFy9RnaHPLldqCcMuE7cDm8AbXqxrTd7xUf3UjVUcDzQldR910K1b7wdcewnhckj
wXZSWA8wsK7QJBIWbceXzwYHqhY4MQz+5GOgL8n3Q/YvRTUGPhKLcoqTjse+M4ug
Y41q6kbfIhUDJjrYRWj9YY0Z0gnoUCHHD/HxLsFRiotx5bNYc3DXao7+EK72CjtD
sut9WPvuA7l8BOeT9izKeqbiFBOIFYNC8CpbbUOJLlrnrtgC7ZdeiItBlPHvrimp
WoKu8fwWa2ca8w6zWEMO4725uHXz6T7s7bQWSr3X7fSXQKVs3Qg+t3Ibm1Q5+hqb
QV+9XNaWr/Rqcyf3BLoAF6QVerKiuN4GFiMQSO4P46gsKJBwuLMIGdLnHo+YmHR8
HNIryBc6kv8da71XGvjkq+Ee2HoDHbda42WPpc4KIoFQmParU9/1fTVktroQ4kWy
NkQAh6kp162uGpvIKGmtx7zM3Oi3nd82kIChtEZQG1kxA0eHPZY0FXBHT6+q7KRB
wqDPX/W9Ac1xG5OmmusRfke0+I2EOVX2YDCu/3W32h6ZIu/dTS2xV/ac/v9k96+4
L6LMNmR5esX2tVYH+BefO7Y2HBRKN7g32nF8kQmllmcX9nDxeqYqdx3r8wEsCx6o
kEeRrKR63JkD2xzTZqoLdO+LeSbhI+0vTz9eyPsueigDSg20BpcNf9TYzwK2twGk
lyLY46yJawOrtKUF6cChhQn2tU73M3WeN3YYb13y6oNeULkYdIt5D8u8PFXE9or9
MGkKjRoPN6I9SXUqIgsgu6bSyOQY17GqhtPLpIzX+Q3lGL7bHi3eBDYtx8XErgpO
No5Exh0SgH+L9gUs232Q7+I/EJJw7snDdFG2b7WUR5nq0E83+r5XDKIvzJoWVctw
1am+D1hQXJXdbnbjq/lpJyBDA6K59B2io72Aoc1lYFkQXpxIkEouzcU/0R5et/mT
CFSMmXyTUA1JsjZ+FkZbUg==
`protect END_PROTECTED
