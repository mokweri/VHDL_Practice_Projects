`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/4PVfrr+NWDpULumSF4ZciIy1JA7NfpwHn49gBRvMoZd9ggA/rHsfKcJtGq9xr8
XG+bVWH3ZjRVrx8Bqy9zSuD/WSxS/a627MQmtDgezJ+T19zjGbI4smGKvOivu0Kq
UF66CCr1SzbCIlFlj6RYXcKyeJOYsuPKLOCtsnVcjMbbOulxct2J9Y8+ge1EDuE+
827A4cY0Z3kDUn+jzTNQOBFHXZomxv5l2tbDZ/kLBUAcCsDqUsb28gCyoJhs23Ix
DbnpCwxKZEQO8J/UEGzTYnsXUJHdtDPMugRqcsOFgUOZ4k2RHA5J4CDHmsyTQdHP
nQ46E9mQYDWPbDKp3JBLt0JAv33jzxDAl8M20dAkEQXM16WKLDiIV0VBmTFu8Lee
yHKtzDOy+tbc5HDBIT/Ggq0beGyAUHSvBOjwxr1VeHYhBoSkmz/81Jslm4XIMLmW
5gPH5geMr4HRABv/5qhh814M0PRF2lH0g/WFF97Qo1htZf0FeaP3MwzOgyVNq6MJ
xs/Lc0gI+gfo6MHXzVl6GI1ao9YB3ob9HTuyjJ6WukGevxUpUkzdqK/NEOoK1RoI
N3DnxZORs5T+zoMmApxVdnzNS6vmVPc0vg6LwF8Pc5+LCx4lp7RieUhkUm+QmjZy
bAsvoMa3ZMypJk8JCv58vFCrpUw1dQ8yV1FFezfrSEg3YlbAE+kDPtlumxqqxeo2
CClzU2jlcfxerheZdJgTy4Jv3r73GRXI7FWkAbrPPdb+sp/A5yc9j3GRm14F/4I2
Kvr1kutpxHkDZxbhP6apHDzf6tqsRtgW6bCcVSgR/EuJrAFflE+8R14xNzBKh3Ly
`protect END_PROTECTED
