`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czWQT2fsfVXE6X5dVUmLmwj9TSbFlKc0hdYNkxSaoaUJzCpt58PjC2AhYoJyyfuN
eGKKK2gR7mHREszY/gj7ltbcl1jhlQLe4GDw9Ps/rekXpZ4A8DlySQs1++x3FyTa
nRoq5hZUqBYrAuAVkZlvpN+M21utp7zoFzMoCy9QtTuDwOrsEHlnWbmGqlcH3hZg
QOVekwleu0AbsmI5uuOVl+/XnJVoEDdDGl6R2TkYmdfLAER2xz+c1UOWqLlKBK7X
8oEkQt1QM91/0I1ajZ8dfC9heWPpInDflBepi9c9gXKsOhImDeDU6kAKAsz2sGEE
i38rStTEoYpyIxc+z52jMTlxCTCPZjtSn9QMdQdoUkTVg6t6NDUgdJP331bxyAdA
h09hDjNlYSSnEkqFNu04zZfONDAfernDuto91gBGHaqBkA50QaIhWkwo3Tvnbrzz
vvtRiRp9WU0NKbszpdjHdNS1g3VhzRpbjXF4j3s5fMVWXrXkeZweGOTPwRD3NjfK
t5YU+GqBR6E+z/5pBmRR90wbQX5D7ibC3VX/f4g9bCiABVVDS0j4nfunYqP9XuTu
8Rx7uZXFlCcHYIvngOxp4FxBW0KQL2jorWxlkgIrQtxUBASi26fw7QSd6g4MPpLS
FC2uqPcd0m6dMn6t3G/z4OR7c9YSOCYT+OD2YZJNSaonykRLxzsYum4xUMA79zys
uSrebgfCOwwNzwLzJuQoA6NwpK+Y4CYT92u5TnqJSjg5LmT+WTFxDAhh7nhCHzQo
CgqbBMlfzWQaaqh1t+xX6sEvrrk91JQtnePtwQ9Uwu8fRaEJYU3yOy4e4YK8EpSF
dWC/Ggh9x22iA+gNJmc2rUiQlw75sLU6efbw0kXy6W9HYoMRybgc6nlTKy1cjC5W
8c5/0NrXIRQanAI9qp1QUgA/wKNpyafUWyeOmpYxQ27uxXlSAFA/VTWnHTsqXnor
K7X6qeKr+cjljGrqH6DoOnwsJgRb8VxZyxNdEoJXk12ONaLQjBCOMlI31K+nJ9fY
bngz1PagHFHXNUsrZWxv4Y5qOrhmaotvzGsFcsFVAQdeN3okoQ+dkSi/p4TIX4rH
F/2mV6j54oCFWO0EYf6PpbbMQ7NFO/DGao6V36M75/8fpn+HTzE0rAeO2CR+tsgS
myIYGKFLKTiMWmDOTMWeWuonGXevoyYi90A0xZp3TAjLlrb57kZD+D3XVAywAQDn
ZvGf3Qp/yVevyOSgsFFul1QRAvlFLeENikXofIZFpOS4M18u8vGHRH+RUImRxPSS
17U2RiTHTov2e4DNh9UPWiXzGipv1xvdtkmhEau5Y8lo6ODviXkDsvNTk3iN1pgW
Cfhn+38L7G7ZC8Xum66mhr+jjEnf47wplUxfrCV2p0+NE1PgnpYuIEhxFCMMXj93
ehVH3kpaLAi5wpCpcMLKZW5fpFp+mjIw9DqZ30I5jCGwLAGMiAgcfu8kYALBJfto
m6OmsVu2kgEgTks8zRsCfTDJ4Fc670wnx3HbqOFOeOKnYz3mfL9W5tUq0RM4yJDF
MVqH9MAqFS3p3OJaz8w+pXyr88kn6VjSWpbKFUdLNJ5Bfn/4xpdvoxmVLHxygFch
eYh+embApYEo6R0YnvaGywv45jZh2If1YP1YzlIN7sCREo4SgqEn6p04qfuplQYo
HYz/pXKUnNBmG3TFFwPfioYOqHA57mIrw+8C6lskzdisLrQQtZ0qVVQlNY7OMxcg
CvXytHJQIsoChMeoBYUVO9/I39V3Ldb7PRHrGlEHRth4xzBi2CJcZ1HvAVVUpWmw
JbO4pQdALPwQeLbC0cM68ISTsmBKJd3mYDROcbM8eh44lRR2jKUXVfXyzcpM2+Ub
0+/UTXa1P//VcNGAgvqoN/uLURjkv8ecteAQBgdd/qpA8C5mImp51Rz6sUOFcDMB
T1A10naUodXkoXyQjBG29uSQy2Qm1evUT0qck7V+QMfj7m6mdF3dBE+cpSSdvAw6
gkAqWz9NvfvyBKumZ4EEhczqbmdRpFn7z7KaIHvQOCRO2Pe50ufmKKZCpunDskaF
ybK6pHYDLSBCVkYD1wErbByq2+PVDVfjTxTmzhqgZ/YqYUjvj1cTDdRmOKQnkqRZ
Bo5jYdfUa1g/r0MftDj6iAauBwclaIfSxa+mDRkFlGVdcYJGUzENPAtekhlPFkls
Me4Z2pa36gr/UnPIbWypc6s8Zsroaijvg27ruPE5/VC6f13ZvjeEQASP8gTBH5S+
JHCKByiMLpHCgsbVzgcAriM8iKrJaHMHE94hjBD2h8zKCdqqoet8Skbmd+egvjdA
q1AjPlyLhXk0AaeyAG1PAcDFX/yfpyovuFUwa+8Ziv4V9XpLqIjJmkNQNtGgNYXh
EmnNM3gLdzmvPgGuAxPs+CUerohYTBj3fyeibzLS94Nm5+FK+dbEM/nQGcpLRUTA
WgDhd78hzAB0hvBIu9TXuQGLoW5ieS4y/JW90/HsusMt5sG9IUIpfURUFSA25JsL
W8wIpSksW6t63EguGRslt7YA2Hl0gEkqqfHhOJUb9DOulAb/4FeT/RG+ubwpFoF/
b4rZ0RORVNKs5MGl4nai5VfGOPLyHBp+psD5gpB2hsoXJD7G2eLFZcA//YxDN+gK
iLw089YKu1eWAx16KQGwUGM/e+GsNjTDsIjlnYvPyhGtXhfYWGvz5sRgbmU60DM+
h2Q2mwVRYGGz/6dFegU2NO5L8zKTYHiEqdKmPIEzSzAwBaRb+GT4H89K2W+n21aS
kJ+DkcuWccY2ghvgW5ejWjUojF2Lti3MKYD5AW/cx1SZv7+vhj0AK4ARaUPEG4bd
oLCiryBQaxlZF5fJYkEt39xP7j2Pw5hqnIef+yN4aEOi2mKtHr0bxWXQ34scVTAA
RxxJ2WaS9hfG8T4wjInvKzkoDCEeM1Buj2m5d3O2UB1KVtFDk7ID+wzeDoKuGAI0
KASYh48mYz7Z4Ik7QVPi1tLLmRAOB38YoPPiR9FwIaQw8owihrSXyT/k9O0rp7mY
2LN3qfe0bPOAnos55dlkklN85HBBh67ZIz925B5swpZY9M2SvgLudladVgsw8xof
jz0Ys4mlzbAwpNtkVp1tqc3wchvYdaNnSqdGmgnAlctuUinisdDvBX3PVLkm+FJN
xAuU++qVPCe+fLuZ7FN6eJ8TKWhbgc9WPSsoatdfiAhs42WFNzolWBH+ilzRdVXt
qpgEUGq+Q1uMpgExcHQQ+5Sh/T4A6JXtuGRYcbyeFG1nXx6JVgu3bsi6p9hDifNU
4lc6blOYTHXeH3gUkGjGCcbeQ5VrxxGsKFFKNoc9Ekg1ZNR8kANYHV2OdD2ocMuC
SOrU6KXYnlyNtU8Huy5FCMP4G86/sIP7l1oU9bbh1F+rpwnSMAkTIgcNmMK5TdXq
XAyKDwyXtXKB/ZM0ljeBXgix6yiStzQKpduwLJTOjDWt9TMNyl8y1ajcvVRwwGOy
zNS6wTgU3mzqUmXFI8Wl+oh6jeTfj3kWl9hQ9CjstlHqc2vET3aqbFFqtxbG8/+E
1QL8ZQJhTiHE4QDlpxSnSsL1/J3ycmwCCPYvp1aU8lCI+LIO72R6m/+iIeAtQ4A1
BPzSMHpu3H6v2hleRT1meNj+1b24nIh3ScP5J+diTvTPypqbpQV6Jy3DkcmlRR9B
fpYne4OlG1pp01yg3K7eejcBLb/ciAfWhoMK1j9660Az2OiM4On4fFOyoedsNmIW
jSiiAYFSTXiI2yO4/N5N9fukK0Nty2cvBtu1V8j0F6NcmLBKwiV2tTALx4Dwjbh2
RjGKr8OZ0m0iwx0Z1gQXecOeBGnu9i+sDOCgwNs00inz7H2c8PhDAIXToVILHBgo
+tSgsO7vNim/gvbJ8HBqp8wVpCKsCa6b6MnJRIGNPwd4FS9jYAgtmU+a+5n89LM6
xftPWGEUx9v590raFVryXsuQqTtZMAPkQc0hECTtjUI3YSdLMBekWhiHIODaVvCu
pRbvyzD+6rZWHb7ht7qetfjEB2hvqd4g9vLXBSItqiO/pnHWPBYW4RUEHS+lQwEI
cNTRuGmK59I4cZkvBgNoxIWwe0C2HLeUS2RIq0C6Aw6NHBv1wFQRVYAgVjAWfHE1
uI/GQ1TtsaJLYhiQijAiWFL0HKvZCXep8f3Ciq1wLmyuSFf8eb3/RxjeRpE3iTcL
dOZv0GuoswmlovsWZEba6urntbVh9vOvc3RzMmMZSf0qNw3vNTuqZmYsf0SOXc9q
JkmATriHEh4YlHGYX+ZDenqp+rSsdCEOuAyYMl9BGnN//ovOThBS9cLyj7ONb6ju
iM6NXgIwWqJhXF+tZesgCF/W+iHCN4IuTDuEfxNo+UpRT19DSc6WmUHgJ8qDXPK5
oGZQDHBN3+skdE7tiL+c4PoHHKRCW6MOJU6x0Fuo9mfcKXBGJbjGKBZDj99XrUxP
prYyveDvGbjis7ktnRMpWXDqHcBJVMnITqC/6PhoUlExOeLkJudpqVYNnyKox//e
BPvxOeqhJA6uzSjv7GTbdKIxaDvsbdUyPN7qJrokFA6MV4A43UNzos8o66duci22
LrW61/QW+PI5LcoK2RqMs/BdJZ9hzwUoQQ5bkj+UY/wYGpcSRf1amR4ygH9Q6PSU
sQk3jp3FY6nwAByh9OETLHITRpo0A7jzSts7F4Nd3KYU/sd7Svc077xQM28SmH8X
ZjjCJchZUQMhdYpabQzaIlqUOSKTXUP8A2Y//GI3n1wjMmDeHRQ1dMnkvG4h2cjk
Gcizyduq8p+LjzI8ZwrZNXcMzUCE0gnnAwRpEbHVlNGEUcwVE4SmRb59JpbIBvGp
W2rsJRxjYllMD/nei3oyR46Xgy7DKeyQUMsD0exzn6qMCy3MeTdm0KAKiM0P0KIt
Jal5NaxuJt7AltJVep+TLk6+lohS+ecHmYi2xqmMPr4ETn27gqt9OhZZ4BHNiiPV
5W4RseU8kI7PFRs0LIFaInznAaYQ5QG5p2hZ6frgZ65UDFBgfo/qmYq9IpPjRbGS
lDooVBCiAzzod60rIJ33v6Gg3lwNxrfZpM/yJotGtT2tBTBBskEYlgd+fjGde2Hh
2sACi+jyL/gQwNEbhEgUDhlNYBU1L+cH+tki45WgAZfVhnBXz+j1MIQT0JEhy1Qm
c58CR3bRuHroacsy2PRatgm61ox0FyuCQaaIst0n6DMBnKXNG3VNpqDPsO5x/Rad
0l3SN1qQ5sc/8JR1YN7p4yoMT/Aj7xvpuTtoAXoVuZZEdOtbyy73xy1mLIcRFYIH
DFoFwtLFSb0fLyyGIyzWJDXYXq5sRJKptbHxzCBEb4exy7r6LTuHxAYsWGJniL65
Bq5TCOdUQ+VRjanVCozeFJf7AwGvysU5HLbBZ10oR8AvQSbSm5223qh/FcPa8mmh
HuI+esFhzx0Z/n3rgOYMUQhszhuGPFQOFceGJR+mcpucMWFb4bldXSTb76AtTEYl
vOZvOF1EpHubowo0GY2I6NA7DOdgTy/wWtPLazT0crfNqBnl9/veW6g96ka6RS74
SRXrMzcn4R+cvjHS4UKp/ZzEBToJrhmOP6gZVZAxeNjwKNkRoYVsTTvBMDVQRgPD
F2clUctMhIWE2IbLOtDXXuhqI2oS8Cz3/soqgJnWb/SIFb/+Aewn/DAZdZt5tt+8
TZcp+fweIf3WcyzpQ5hu8C8lfI/x6gbzhFpJ3aXitvbVMeEaJrDwSld93hPOla4l
VkPg23ezLxb/JQpVRhOAgMvL6xWBi9fztMzILZxbwsrrpO+su92UafVsCBW1Ca7W
uQEWjE+9r90K3U1X16WQQy1Nry02we7tBLHp1CVLFKps9HPgGas3UA2RqNYSqkU1
vxhNLEUiZKTSQf4ak1kEAauYq5p0ClMDEc1zn0ztWBwGzTsFrOhx4fxgcerg/M0p
Ubf9es5lVMyvNHoRtxmH6M9WEjDeRgy/uFf3vWZ07B3qCa65HswhBXIWwLggjGHc
GT4ZyEnD+AQ53l5t/qOFgmgtkyi1i00QI0gPoyye0skmROh2LJ8ZVIfVi+Bz1+2v
1pUhq2tqRw6mRj6w17hdTa6rpORBUXYerQLpQQwosKuITT5Xudhr+fRV8H5jl/Nc
ggbGXfMx064XpRUCU5nxy9AH2sTVCj0W1RGp5MaQra++kDFJ3u1zSpthFhJUwBS4
e2k2sNvydEwGLrjLU/FBi0d+VvSkRVtfjNkaGXT6gsGqrCbgsu+LAIkRzAmhDwvQ
RmKhFRoI7Eaf2vQiwdoFERTIeUeoqQT3Zrwa5NbcRmF0Zy/O2CmHzFAOk/DU74m0
owP7RXvHRj+IUrtplWFOe9gYwdhZK71MZ8/Kq6RSt6r6V/LIeOfvjYYwyvCr+M/M
5Dcgq+KxXWn/w2BDYXIdoWttMJzDc52Tp/LCd7TfGc/zZn2V26kk3FGIPL8ovsdw
JSs1gTafw4oZN7voAqYioOtKrioNBZxyhF1lV9oCdv7n1NIZeTLw37nqra9xV8RV
krR7pD7weKT2pbLskzEnrCb+096lW3NONNLCId0vYwzaBdaDkff8QXumIFo02CI5
i1himr5uhSqU6aR1fAjmzfDl+dpxB7h5kP2sVkAz+SA2crz6G4riOEDyq1oSS6hN
uGuhUVG1M1qJ3gmt98FWZaRn+VjpfceL+TTbt8aHwvdrGS1HNn/q58q96VzXV/tn
hl6Ir4i0od8Mc9Feule18TaE0OeiVK9eGet96o/nTIvuepjJ3cxg8NSzaJO92Yny
ymA3DFl0QyLiS+hHLx4QBpUxJ7BYwn/XhT+0bAt851SkTTWxRKxXZNprdy1Re52B
OK7RgLPSYSeMav0aYkf81etKxe5wKhBTMSSQZMOF67Nbu3a/7zSxq4p76gQ3GbDr
3nmGjBciT4pWqpu3pf5WKatwwOn/TChlx+BJgz7jRsnmNrnaAPsmvUuQl4lZWFuu
na2KUsV6hbl6o7gJGNNuPAg16xuryLppUsHGlIuJScJXhlf7wI4N+vOs4jGXRA/T
rjz31VnKoU+sPdDTATYoMo9VtYXgshofbaC0On3nv1kVOIpf5t5qnDB01FYCMMxa
4FGd6+pbIWeDxwNxNOJrBafOBzScaIy1B4Hfz/jZMHjB1HsZtljBzi8ZWXVZrwJT
SxMFy04T/4MYw2w/nISZQYdCqzmmVbINrAzGVMZxmNYHXpRoSZkSCUbTMR9CYd9C
eSeY+Ms8lkEOqDaVXhVNWxIXLA1d/LMQncXT574jfSIvxSz/NOpGTOkRAe91Fbve
8NfdYA6m0B00bY8cRCW5XSFGzMLJXQX/rdaea1Wmm6fKewKBa5g9YX5H8uouyIs0
DSjJ32QZ9T/sg6RuH5n4q1o3Z97n6Gx+rAWdfqUyyi3s8wIGuCoAYglA5VzKSQTS
rzI+R2afW88FHS8K5IdGgZ5pnF+/I99vNP+Uaw8zsjTERw0KRXkZC16kkCN4Gsvz
aecA3349PfYTaynGuTmSHtCxOp46uKU0ziu+suUC8NySQ/+pZ/ghVweSaKS3s0Lg
6jlOLTCk7zWjUWX8+M7HuP6TS99pONakRfJ29W0Fu73nGEZjGJergC6mkF/NzJSG
cuBIZDpBcoGOq2XmoGnsZxyOWXIoil2kQfk6OJdBjSUlbeYBbSE/hgE8i2g9ppwh
bru+ECthi8HWGzZ3pdTqL/k/Vem41SpFovwruHpISAHm2k+6hG/czebj5E1Nf7j3
KQcqUPFiBJNGhZu7VSR+8rIxRwYwc3fll56js+sxoKJobsIBg3gTfHG9xtCQPhYf
FREUkClq+LUZ5QscoghUhQ==
`protect END_PROTECTED
