`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QRK/MEQuI9zEGgtW1SHyu5KNYPbjPTA3P/GX6s8tqwMPFQDgr0IduO/s+1VYSGlq
GxaLJuaae5W5OcOywmduJGYn0iQ7EeuFybI7eXXTAlYSOsrFeiklBMcg9CsDSKui
Mq5O2PLgmjX1NdiN6wCt+Hnywog4HHlgF6wpc4OnT000WWDePJCQ8Ge8QRpOY/I4
18+Uy06XR72C6nC3XK7+D2fmhV6JDGc31zgnvN/iXoIPCAwYpnV8Xer5Thwkdv6F
MLpCcEEBEICno+pL1R1nwKy+fco2rH/ZE3egf2Z/1LCnwPlIVhUDWGIBYebyH90W
C8kz9FJ3/3xeMYD+0r+7pnYT3Hdew5EkX9zWuJPwkgGNG/zdBObtMStxQpJ7XdDq
bKrVlAzUAFlncwOskFn7wNSjxRafUWzRiKbyPe54qMWMcnvpPW34fBtCT6mZr0bw
KtZPiPVmh4kCuqnBKnPFfisOMM41DkjFRT6nyoPDcKgeKyM4Oy/17Rm5NjJb2na+
0l2lDcdlbguHmCwxFUEPgMmPoS9vNCkrZ6+tLH2vBZ5h+NsGNexojEIlAnpFl27X
ui8iO419zwylljlTcHdav5d7jHbgN9eQPwDtACbnXBLmWTI4WJa94ra0jeFewPRl
hgSOyuQNP0WGkqPWz+kPa1CIRXzMghiX2GWlgt5kG+HcZzV4E8uFnHn5rtAfKFze
J/hdUNOTGX4PIL3GB+1CVasvs0+Oz5It5nBQvmTx/TS5UQ82gxSo7viK8HOMHBoR
vvKaXjeV38P5wGP/6Gk/VDzZ3W/RNU69JRHlxUJz6nJPuGnhk5Rj+xjcHIK3n2W7
j8l9IGvVc5kbyUkr0yj/7WdJYcwdUIYrBzz2+R8d/W+2mcQ/1MOls6ufFBmhNDMs
eTK/UGpOlVpX4GKyYkBmJnaqd7Ncd4Fd0GMplnQmBKCJsiHsjw3PHVSNutD8NiB1
xDQ0t12oR06vW+wZHMFDUpXw8BtsEzBPnZhdzjNmQCJODMyoO0q4FdsRIOCvLEY2
`protect END_PROTECTED
