`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ltHJgm7yDbeyHmvMyXS9sE+rcJcZh2tP7WEjF0l+EF47wJO1L3iXiBuIWcrA1d2u
3m9z342l3EESBLdKS5e99VrVpAPiSAEgRjIkGviRq+rf7yMqz8VHz0K3oExQP5N9
zpL/o4Qbed0Tj5/D9cdD1aP0m4MEaWh/xSfnmDixpuWvRSD/Lfrsh9EzV6lXJhjj
vKJVxDUA0rfo3wZTZOIHE1zVvZkZgQHw0jd/XieOWO56Vxk62E4UhvCYYrnj4sRE
Acz9/jn4OurFxV6z1ajxc7c6faoClttP6kltZXs9bieLIUx/VZsDxjpvCzckLcN3
GnGoWsztIPanJOezNcssRH92utHBXyX8EeL7ZrXA/vxr9c9fxl8daSEJ9n107Zv2
ebfGw7OwkEtJcPuE0m0NcLwxGDeT97loagOSOCCC74vvmIObD0Sf25j8w7h517XP
dCw6AfTx5cpfj5iuupHI16BJ+EMW77Y0X17ceq3Dss6xp2/jXYZUR/VGJ+1Ltz3w
2FEFb6iqQ3Q+sWKIbI8pP8LNQDrbaAt8ZZ36PvS570JI/+fFOBYgBUqeAFFKC2sl
NXI0KJrNPRKiM4PlnOY4cU5uhiMg4XuUUgfvEJW/e/U5Ke3fzqvEOZBHcZ6/uIvC
puIAvK++3htPkp03QIxi/RT8uPQiQObSxHHttB3MB/2feCKGF5Y1bozoZJ7zYv9p
O5wF26y6nq1/kcy9sG3xGXMv4N/pYH4S94fIRWwJUrDD+MflCvaEfa/278hq+AGm
WvAYzByVVfgnPZO7637iFYnzJrh3WuLBfvlkWgTl39UZhxaD6G+8Jj8H9C8eql0P
b9CvOgM8cV9mSOt+LTPHv8ALZ0RSzCpfilc0Gfx1j5UTiAYcWZtb0efakgsNxbO8
Ioic6UPuE/NrrH3Acavw7F2JzgP6qhCtosJF1SspLmZlUrQXshCbeqbtwGJFo9RM
C5qOFEVXzJUJY16eeIUQC+QvHJDC9oIxoKbmaUCnfCiKXdCd+MDO+NTKzafx9ejT
7stplPkb8iJ6akatHEhf+Xv3QUfyb7JZoLfvCwQPLdHBR1Egg+eCKaFRQ0jyHLJk
S+zG8ImqvOPVLrUPsjTV1baoJcvu0XTY2FlZ0uRNO5eBLCO6W1RkTGQ5XuzKbfCc
j1l9vlNa3TDpGKrqYNdA3iqeX0uqbjetVRdqzP/PGCYOAjE/gdzOgp1qEUEWzVTa
EcuUGMQkDBLe8l6iEpN5UE5IaFuCvDpcefHwLKHh/uMRxrPN7qz71V2XaXFleWco
hx68L8hs15AsCe5piMRQYzzKfSWXitYroET9cQDxBsQ9S+TaadRqW48BzZxkmO47
gfEKfkzyzzVkmnCUcCvl7fTe4qOmdiJEU2pzPc3KxN9fG45YnqjOc0jVACaXH9qT
sMTA8ScrWEW1LtIdlw5taiMgNU5FChrr5CX1c1jbG9QwP2Edclxf+MXEMDu7dsQB
3YF/U69jrFZL5Iy/F3jJT7uatuvh1bLwQTGMzQbm+D/osUeIy/LKgAHlX4XkvyiQ
QLbts5z4S9YpogZRKEivUQg0riWmHaOvnrVwibJ0IbQHSpsydhr2rLruUqdhMB4+
8yn6xbZPyHVYr4z3kcDIqHFU9Ku6MukIRDvzq0NSKG+tNhWEao+GiaSsHR5hOIwG
AeCEJscl9tVPV+PulvqaV1yjCOl8UPZOYSQXzq4HxNpdP1ft5+JooyktzysAdsUh
JdRcc1f/B7ssuaUlqz1lo6xLRTxu/QKGun0BGJcBaj6hgmmZU8DxEeHBDhvmjcU6
hEMD//jaSLffV8bqfMgcuB/OTvK5RjT3TZA5xLxKzs52GFprTHYTayfc2G/1ZpAO
pUo7p9XfY3VTvCK6tvwLX6PDCKeIXs9/mN2bWqVSJ+g2Bsg3R5cDocmw1QSTKDK1
80gImiALvwWoNDbmd63uO0x1RJ5KmJwhRSbWP66xW7K3zkJ2WglSKVLxvCnp8uIb
SlMT6W3CBThcuD1BEF4jLG6dcsgcyY4NYg/mI3aT6MCZxlj0kotD2c+hHxdU7Q8k
n/O3++CKYutgF5lyblRa4+hgOuM/I84jdj5qsYOhPfW6npJmWhsIiE7OLU7JRexS
1pQrTu8j8wKEFVlE7yMWREKAefJmD7nqjZwZuaryhEoyCesiD8qQxnYeu/hAUiXU
alOL4dRy5y/SCjgXTau01dnmIGbJMSm5JRzfP+E0/P4Ssu4bqfiRsDfpooysZ41V
DmN4s8sVr6vBkYaz4dj9P/qhP7aQoc79dlFP/Wx/jmkEKrA0EbIGMvKMS0tzMKlP
KABalAOJwxoxdzXkUjNjlGUhjL4xj4NLGNeH6bUWDqaxjxWILmdH99RZFTRGvi6L
etNKI3TmIL0VWGj3U2JZWUgDasaoo+CLwp2Kj1l7H1KAmhryDve5XPF+U1OaTKjJ
1r9MbT3MsN5/T4aGVh2bVVw47CMcMrMQuWfsWn7xCCPyNBj5mEqne/r//DcIvKsi
fmfgZa129xqrw5rFWZ9/EYSTgIw1/5/HPqDaY6gMUH9GSrLMWZTbPPBv6BeoSGAw
Pa4YG3/pcJvEEqiUOKS0BuN7Azep6m2cUV3Vx9g/mc5q1Ux/ZssSDr9T8hJ5hNrA
/oqVdo5NxoACLfF5i9M+I8Ze0j+pbyw8Gt9tbfdJOj7/PIZCbH8MLBWnGZ0clMTh
5atfA5Ti6IJQie2hcNYbM/5rSwylz2U8ZMkeu7ForVESrOfPKsTPqdo0ZEqtEvL1
zWVTWPY2HEOlhAuFcxatGhtNGkV27vE9yk+lW2EiaPbpMDm6zm29gvlotQfAJCCR
fuF3totQHA/LgR5qqVFoKbpHy2Rwkh5zGKZZtG5436rgCEum8x5tASs75y4dVry4
gDvBAjINVjgALowEnRLBC5yKDpYqpRq0VzAOwHTRxIozxrDnaYzFu09XOjPXgU4m
iDQoUdtSKfzdTt0HEGtKKXMOk0LWKOO712iETBd1T6dRr7H3ZOulfsmFY1du6ly5
sn4QKCgUMGZs0tofP7LNWRKWyHC0jbLx3NILbI1W/rp/UDClLFQmxFJUtDkAyd3C
XKx7fKt896j4ZG8a4pV8laoFNdZ+qpBncx3DPDja5GGR7FjLQQ51y61GaCMPDxJA
HT85t4Vzd6tXfaiWLNEozrL9SoapVPg7uE+Wh3gTrTwriZFCNi6ZZC99pjxu74lH
4C2/IJn6PEhqkC+OyjHa8wiwu1kYcaVxWiqzfVMDZEXlRrWksBZ2ELdOc3Sldrdn
EbasOFvrU4kjuWGoRjtUyqWhI/AMbcziXVaM9v1gdyLOnj0T5f5CC//q0KrXfB6X
Hu1x1832WKtj1SWu0cxFERepjp3PZHhmSxEe+hhjbFcSXfba6+TPgSRqphep/h6+
SrNpP99ucOcu4wHLFFNzUPX6cmtsdjyUI8kOcblyKoz5Hvng3B6EJUtoxzHIZlQq
at6kFfdmsbMNmQ74/ztkVKwMD4t+AdxyTKDDpeySRuSN7GpW9alksjTuMbSiW4Ue
e4fFIQG5uGEqDINqrcEm8F92sDC8Ng9C/EwiI4pDzubIiFTQcfPHTAN8x4Hqlq6k
dhkkkT6hakymD9pD4Eel7f6m1zCR5L4E/WNrNCVfRDRFUmUdrDMRXW7lD7TkiDbv
RwYZYP7FqspxfgivuU9uKYb0LBL291I5+ClMKUseJqz1Mq3kjqsPA1YnHSps9nYu
RepvK6iT8SM60C9pOg6XwcLg5Em/4hW1hEpDlenTvNvSONFgilHULIIflldhszkB
jbqAeMCrDPh4fmLDqCWqGvet0NFoLrjZjIQL8DAbRgzpsc8AA+IcrHdsD7ugOrum
88G2uf1TYqKD6ixXvCSoaYLwNv7xdlg3PoZbVJCQXX+2Eucg7s8TkI1Bc0zSZu27
Ly0VaePX3C2+Omy5pmzMccrFeDSXeaLx30qOCRQ44ynxxEe/evziLbhh1eti5+n+
oSjaLszAP2pKEYQdLx6D1pCmkKahKw51KboNakq/5L5AVcLQZs7QV3Gr/98i7Y5V
uDT6nlIFFm1fBhBQXdTomLVHHZWZQo40UstyezJ+OXKzTZ2Eu3udASuDQuJWO4Et
rUlbo9msejnjf1qlNHsOCaIJJ2QxEUkuyCK9SuOD5EVZpbe5vMOiiXEDISwqgYOB
B12Sebz9LdFHN4vxW8VlamVL7bDgIWaodm6NudsmrCnpClV3WfIcukd/QfFZoW6Y
lVpLpDzm11+FoLcSAHIq2b+sTyEjhIr5tbfkzA8mxcQtJyUY8GTQ3Kgw4xhTiYAS
skSvkEkVv5Gr/vW4kqS0wUzckNFgaTbl00FHQtk7tH/XmO//AgBlNR7dsj0Ac5SK
IlfPJjvK1Pvo+OuIgABiz/pBGejY9LkpQjWgl7aiAEC6eN8/j79oqOIgJGJycou+
oVDc9CXsk5JUHfD6dkPc3uCYlEcDQiFLtcxvg9SfldA4eKUegRFvSh0a1Mmeo8kW
1IgPW6oD5t2Sc0Rq1s0MgzjcnoWTZShA9kDT7FYc4VIoDLucsfSxMujFG+BNqzFD
oUMJhsY/7kcQKDTok+Db8b5bNk+gbd3QMeYzl6GSqx6wz5bxvBFcvoDjP3nS0xkx
JPZ10iCjkFJ4P27p9DhEu+JtQekr69uiSzQGzfH5C7JpePmISC1kNhh4OYG3Gevf
2BpHRbUpZZNDUBvl0wWqeIAp6FtFhXHny9xkl1dZ0fmvhK1Y6GmIu1I0FgF+Hags
iWVOUED92TFLltOc/dEQxDfLnge1/VCZlRdkZDJr7Meq1XvZvrnHYreD5aMhzcFO
Tuu99lWFKpy4hISkFHPPYGSH0e4bP5dmAs66yvxydkSY4zlt8JDRBxQGk2OXZAmb
Di1JtA0HHr+n7xqsNFMuHWh7GNArCyE7pPzvM7vUsL85nZj8M/P8BxkS1XuRs0XB
JVqO5hTmB6xbevA4r/S2FHE1vr+Y33PjtOiQW7QBnsSdsqUEyGpyLlzpDrrDv1he
vHXxs8qavRfuvmy5TRk4pam4ZYE9BZZCUrBLUC/wwUbb3EEJhD0x2R49r4OgLZ8h
BU1NEkRxJ1k+BewTueTnatYdmO7WWB2OaW/Z32ZT8Mrj8+PFmguMUFJ0AjTe/RFJ
NBRBiz9TV2cSUKtM6YpOqvq23kKv1AF3NSQcBDJ6LYrN5iEJ45UtvYBhxRUMlRtm
BWp7YKbQr5jFvK3hVFMBzWBmTJZD0D6l4OkfImnV4kYtI2Lf2Zwbx2j0bpGmWlmH
HEGeYRtIT8s2RIEJE655RSgcB3A5rQqphTsN+LnDGOYI9XZW3vk2FpFVP0RJ7y2S
Y8AEZpA0y/RhS8i3mv6+A/qrTaRsj+ZFc0LUhfbDvDGjME0LBpFIPIndZgho4x/G
Zs2NpeZIUa7/zreBCGmC+dEdBqN1EEitti7yN70omKnDZUelgEJpIF+rOvbN++/y
w7RrRhXtGgBb+P+mtZ7A+MzjW6Ah9pnd2TZIYeJA5x8bEvEZUgyto9Ii99I013th
ZQKHiRZ/5q4pgD4J5huaJWoe0yT5d9HK9sJDnsImQENPxkhDTtAXJjMHXUCfk320
/6eNzjbvAZ4Hg+79jQZSsxfHPTheFKdfu7D3hXIlXMesprULUpz2obc/+WzWV4hE
UeFdndVGtCJePRRXYBDAmRmO0YOzAYl5dk8uvjjPlvM2j3WH3a73icuHKo7wre8j
EbPLPBClbGX8Pht6kaqjLx2AkjHxr52CpzeopngsIP1LvrQ+4rPx4AMpRtG5NN2C
cXMhio1ergyILB5vGxeXgIqLPjzuW8HdtQ/grAywZXm3aJ24wH5wqaGndE+QKI4C
T8yG/BSOO5NPXn+n04zFssSHi//ryeTqIgXqprx/O6y/LGcMHfvudxn5U8V5nY3x
IY1HXUL/mdAGN6q/R67rUwcpWvjv4FD1Bhp9YFpyR6B63DAabpMkeFK6jWfELalv
ZMyq/edKGsgvzdzpnrDm9+nhv/BcouPqqWQBMh0H21a6K8KPVXPB21CtujayG/Wz
gobm+oxg8RhUyqmDxLn5hAivxwS3m3BcX9wWLvi0lmTios6b/rgDc+mO38MeQDT7
lDGPOkwogAeaE+GYW2zn4w6P2pbchDqNy6+VuLPo3YHRm97w5pSdc8RkXLhPCXOX
uPiRuwvWxee+a3XXoDbhADMbZ6rxjoIhrJVUJhkmhMaOvDs+5J1h2CgBdB2YzlnB
CTaTbkVIcY5c3ZoLAcQl10+1Cv1so4roaj93sX/Q/A5HYX0JLx6KaLL/NE0sq49b
tAgAf8AwYZ1qJ3EGaO2XsWaW4zpS0XICZEwWF4GleHfe2uSlAOo4mpLO2fJvr0DA
tMXadbHfUQK+y8lycTdHDjuaQRGiwPWQhEZg1W3YLcyLgi6AwH5zDdz/YmHgQWpu
jG1Uuh675V1KGTOJSekYloTlzCYDtBMO0OeW0k3LdF9CgOcC7oACGzHXh4uknoHE
5Xfrwm0W9pVwIC3c0IjzggJBh6cPF7CFqwmVKFKW0Ycv53NZ5W65+FM5FnuZsp3U
QVSpMTHgtuKtImf0MXsONf66OT9QntHicscx6cpAMKobdiuBdQ7p9rk+zAO9xFZb
wwsRf/xplYaiSvQ51qPf5dzha//FtKa0j4lpJU3SBaqvD8i7BOUwxs5fkZH5KAtW
24+6/GxuBQ18LOBFjn87/CJmGxL0utCPQjYFT0oLLZkvHPSQOAkCfSvK0B5khxCS
v5H7rLdPH4EFWW3oA6gPMFuMb5EJrZ9ImPL0ZuyMbbROJANYLHOXbzlEEkHPL+Ni
MN+NGkDUIfZDKqNhhbge6o5SNuWGqLaPc2v9N9i/a5w/ejVls3k+JfUu8zaGmnfS
jDdDwcRdmoPGvZf54eLO09Ne38ITnw5voFJOOENfGoFk1VZpGHITEpxPZpYt20l9
iBGDf5Ka0wF4nD1UQJKuxq8tb+uKYhK0KMpj72j0jqYIDiyZghBSI69gVlOe9BMy
hNfUW530iBgdhhdJM9nhr5mdroFOewrS4lXy94/RLAozZvjP2y5pmydieZwQkrQL
C3ENjr4+q9ksE+KaRExtdDprZT8yYJIOl600DVsrp467fEfjtEpZkR40Vk/w41p5
9c58UAQG5GbjQRBn4pY7EDfKaNhhj+XIk5dBU/NfihCtblZXaZ/O80vroOEqYNwZ
VWxThyNQkzEddiTb5U0tnjnOZrNT1Kz+IWFxVN3jvIFHRvaxMjrcVSwYnukDCf8m
gCyYdH33Oq6tgk7svMyC1Tje66lrc/ZPOAzHnF98vFxTFZom9/kYcpyWZvZL9R3i
LqxzNnf9A6B69sbkpMx7CC8yvWMEpdB0ZpE1xwKBLstpCb8Kr7hloJBxNuaLsftq
ZcrWlqu2Lkva+V8+7z0qKuCcDloxT1r75XSlu5zWUpKzqvyXXSdpOScGeTteESlL
mPM0DFGNLYfD/JnrmMNzyi6l//aUgs+vSAZBSvaHgJx5qlOyUjoZcybgCN4EO8c8
lqIFhwbqlnEtGxqGn/jlzbdt8pIl0FPwy3fd9vOzr9RCwYUL+EWP8KtRFe+ygJ4l
2wjYXooxYmR7XiJaIKwkJycOIL2HIV8E9j1uPGIctKCNe/5+kmkqxrFgXkHpomX5
2qdRylebdII2UTi2E6xHQxNkICFdGGRf3rl7voLisAmk3oIejKo8W7vGPw0DN25X
SDD5AI6OCLIkSSxUveTgS9m0oUbLjme9SJUCRJEXCmBS3MWxqC0VMa5IIQ6IRoYZ
URYUUNTT6A0IAwt3cXgfSu+F1Ax5P1hvokIWE0i+yePuR+QZjb+WPvRPOSR+0uQt
3roLOAyorg4vP1zAysg0bLyHXNBPbF3P2b5yVqtYQho4jFtZppzwtR89hbAehNhD
GkZTcm2vZXvZIVWIoqOgLWcmzaV1AcFNdkfWD3z1yNIp1tNEsiXwwOehexE92B8v
6hbAkOMLySDUAVB+qIVkNGPfhk2ExfrKVFPzCxLaxbo+pbs2cOAZu6F94q4YU621
tP6KkOJ8zbRY0ASsB685CLJu9UfWx9JogRZnh9nVI44zGxCCnLsFW0YF79G1EKyB
6Ql96jj6hv+T+uzFlgeJMf5JiVW+z1yG9aUFQSlzJGvZ39aitcxstV5gAtXptlbc
YF4VKGXu0OXBInKDsTeLXuUmGrqvtUpCCbtRhyx3NyHNRx5OALcNjIQ8AGYVzVWk
z+rlP5ym18MMTPgBMQq/hg3sr8R0PJig1F4Qd8goTqjamisDyqd1Fn8ML2mfoiF0
+WbZ5UPTzIJ+NclbrHruqIS/aIUP907znV1k+2999kW/DORCXgrlLhJ25Yq/vkiJ
Y8cPT0Ll6ljQ32PhlwJu82qVpuy/fUgJBJnLdivNlhv+7musXEKXgh9fc3eKGx+D
fOEfI+HDhYHnMnRzqBVKiJ3GUSP7QcaoQjPA9MNh3RZcizS7m+9s/4qx48FG8hUR
mvPt00OIwPZ81IkuzlWecsgd6EHvuGww4GP1SyvVzahU/9RrCgOWvDV3WDzmwEU/
8M/nXRZ2Cdzh094KUWiUDJGjr7hRcaQrCmYwaiFRQnQMkYVL0U4zzsbXj8XKGkZu
+Ny+dYYG/BSLfDhRUqXk7nM+G6yTL8BhGfYBcaJ/3NqVSiBTMXXAssRc614i/JEs
l+fuimeVjrk9JCWyuvkz0Tj//C5rxknTOMT3AqzABcHMnIbAKFeLYRdXAwWHjM+F
jOFbFNnxFssc4vCokxduG2mPom35YwYFsK7LIXTRfs5hj6HrjI4sax94QfbBLa0+
11sIBSKzxKwjml7gi+wIKUil+C5TQlt2oUyfTZyKzVmAPDTQg5yz2HxviOdetoZp
E2NRELwqExeoSCWgvv8r/gRdaqOhx1WHPA5HqC1QqiKOfnudx9tG1gi7BmiyAJHE
gwCVhUTQyv+WLYjsMurUggx2QMuMJHDelptcoq9MPrxaNqL4aKExk7UiBrum98pu
Zra8luYiNuRHvP23CyGltbHU1lIWdi+ff0Oyv5V7JmKRQKUA25dIDYJ2Hp4CAQ2c
IhuAEfo8NjmZefgHWtYHHHi2AMszKy1sYNiiAE2/qYCVidRJPpicNCAkth7usZwy
tHAn3sv2kzF5BRKUF/FI1a34ZItUUdjbHTQl2tiR8SdJPi8IB49YiUIipoLldjAw
++s0GykqjNrveEOP1ZgB74d08dwp6k1vmYKz2eYKC1XEEFQxUrByo6/Gmz8uuxXj
+jJ6RbcgzM2YJC2K8pU/VIfiJxCLmWa23yl8cEBzZeHD5HUgRwfsm+rNYVgadWPG
D7SZLJAd22ekQ1APv3KJN7o0d9UoGv10x6VUc+aizO63kO4AX6um44UBpIc8j4Jg
JlvPZ/Gw+ZAlMIHbK7uGhMxo/Dv9oQqApb9bYZQSUVwXmy10xOtOJd+aK0VGcTtG
W5k60gbPr9zZuZOAwYNN4QB3KxjO7N/lk1B1tgWpLVbQn8xU1nHL8QWvB6ztWd2r
6emr3LmrkW3y1mn407GZ+hpau8Gm0g/65x6RjpIUQUkMqgUQvtd03gSv2Pj1v9iq
FDTT8b8vYP8wyPuX8yN1mpV+vm/2c6zS4/WbNV1mps035Dk4uX6YYW3kGf1/Hsug
f+avpwB9K7cHSAy5DdkGugT4gLPjopkWfoS3yZ+GOCPJqgUvHTo1+lkOFjstWyzW
AdEMsHLUWy5j4zPRpFPugDS6FD8yBEodsXzkFDTH3ssNCA/3WjRqtRDGcCDmKAN9
gl6oZONnMDimOhyixpHLkiMq2SP9Z0QDRViRFn8gDPrUyyM0jwwJHHQboxzr8P8s
Hkqgwxi4QvcY1/A4KrDM8dr89dAi5ZeJg+v23UK5YOUgOsKObAKk1ZIv+vEAb8g6
L7iFkEwM+ZAIynSBiiaWqzxlOpDKcq/0qg96nVqjxZfJf61jqRUCasP8pGKUl2/G
tytWHhCGtF6qqYBUbnAoJlKbGZ7tL4fRt0GGwG4OHH8YwG59Rrba/ci3ju5cHqmg
rK1oSXcz5GNiUmklWsxqEDF4MGAOkcJ5oDfWl0rX97KRmFQvxO3/V0IkShrMZw00
hDHS1VtJ4BZJBMKbEIGhMVvyvVz8dO4hl1hVoq9JsJ89i4BChEgv4nAWQS8wEm9P
oczI1rr08w8ld/1K+jZZU+4PNVKMmX04brltG+iWOk46g2xjQiXNAnbFR+h1k8hC
DV/kszFf+xmRqZWt31RDzpoS60qR9OP6SaeiUXKS2+2mRkRt3yql3GgzzQOsX51x
+m01mU0lBjMsJhX3FwcKpDd5N20RMkg1t5iYznfSXK396xk7RxQv+/XPQ2h6ucmo
QTGbYGJMefxupYz/0id2MxVHnzeMN/j2M9QRVhlVPEV1jHmK9/GvLEpeVDzHfyWy
rfgEFH07wcc1BfVRBDkX0ldbYYD/ijCmNd7KbvQTDZklXHQG8OC0+uH7254PMTrv
CCE5XSbZdb8Zyq356xfSe1iSejVDslH+tjVr+uaUksVq2q4Tqshvnb8ZT7YWA7A7
KnzSrmmF5HfRuJEvgPdT1wxxN7um04OF/CcfZvnVSWZnMmyz2TyjX2gNy92ssqjQ
oM8UlQP511nR3rZd6pHUFhPwnVkhxoafJFilnwi7i6hHYQaR47vlkbAASJGYOww9
HpycOdnJ5DU7ygLSKd4ET+CVP4tzE3oi2jR2jYPsSrNpL4UId/LMqYkPZO/zvi/n
pmAKLdz4aFnKtZ1LKPNsntMANC2YO3/1Jz/LBw1cO/Igkg+LAfPL4V+Qdl9P+hIT
L9PalmmHvKTsuFl1C7NSxBy6M/S9nMCzhDZxZ24najYfvH5nHPz5zW46Z1MIlNpQ
9THTZrdykqp5u0v1XBezKaywWFcUwXjWdaFKIe4egzWGvgi/xHgbUNNpxXbea21U
2kE7+W30TSrRanS54cPgrX6LKc15w/K+p+NToWFqFBW5bwNhSOBnI0UyIUyoQ3ef
hzXSuY5G4/vkI6GsiITVYtHIMZ9FOkSqTNvRj/cwMeRUWdIJ+kvY7DS1yiBa8BtN
A/T8dpUZuwNK0+r9vVoJ832OsZ5AggdnyiEhQFueuNe/8o1BI/4U2K+gHzKWG0AP
C81PGdIIDvwkYzmhXahspewoS5yH+JJjAOLLWj6Q0s8WLXmy22zzPYg7ROo0tmcg
KVorZsoHbnKkCm5G+LCPakc9d7wxzXFrud9K1uVUwuaUfZIefr6FLFL4LtJw2fVM
C1fODlTb+bDpbKSM/I8EX37F4sL0gUc6ZRqVieYYsXMnbrLOAwaw9eTSRuP2ou8s
ICX9H94WY0oIkaMoAGaBVvg+KA1iOiw7FbYTK6q0897cNIvK+YMwXxZrcP4MFF8D
u6G0ZrpBgLaCMydjVC0EmiA9wgsH6jM0rr9JrBnye/aJLTKhcDns5rZwSP9VvV38
7UCU/zSrltjd5JVhz/LuAg8EyKsP4Tbyu7Wb7hf0Me3GkNvZKW0uRVL7mNaCpFOW
pZO6qwswJj65vB2xsVXu0s1cIkA+vsVbq7TN1tQPbGw3XwaSHdZ/G/yh8z0MOzXI
572ynP8zZMAqZrEcnmPXFOZL1cjDtvOB4qSavRoEtdIbqMiimo416jwh4CMUigPf
SngIj9szjCy5ujmxXDeb0GlL9zsXJDiPQvDdROX3Bg5HCwLZTEtWJ3TCqTn1P5jD
mg4nkSxc/ZrFD76NMAZVMB9LFb9QpteVpiE8JMtSpAt2V0wQx40Yc9cDbaruJyvy
q4gFiPToJMZIrK7DcZd4HhtXz60BtfCw1I4OrOJijwHmeYL2TNZxFKqquhLs1nnL
YO8Txly9GrjKhoR9fq3bYjDfvhAq0XIzgkfr43eiX8xbRhe8/rjGV1PpRvVioCX+
7uNd5yR0042YW49aKfJ2G8X85kWn1qr4irvLdLGV6+q5IPTXFdemtVDLBIXEKgei
fAaLBzJorx2j4ottCxfbWGOp7b6FVvF4s06u8/rvUA4JvK4l6Er0hcMwctI5Taa9
DhePD+aCEkAGOH/lE4BZpZ97ZGMv83BWNDsNG05gSa9PF4PIphrf2PkzI8ZgSACZ
gIL+ucq6QVVL+pwoJc4Kb/ICpUCEFFr6vx3fNGaiuhTERdpt6M5BRceh8posxeWS
6GocK+Vq2wnkiA+HrcjCHCsSyaDv7oiDJifjFzW2vqRNRnRRAPourYS2aKQQm0Ey
XCJwdotf6+2/A+CpvgqyLcqf6Gcg6Mw4QgKWo2izToxC/SMvUDueAAvs5aI2TiJV
jF3gdZSnI4lHM/wtA8Tc17cAf4xMN2AuOejGz8TRefmKiJJmMLNvw1yCf4lHfAcd
d51I7zrqStg5MXLAFN77FRp9jDrQL2l7cWCbXW/Um+ESCAuTAmdXeAtaQhyaOmnc
v1AFNgD0pGvBLaYRowAoT/naPTqagyd1H3CmAumJtzSE3gMrOcS9Lg+bZ3lYy5AJ
qm73NeslUIRlqm0rCpjcHheoPIS16j3kzsuujNWV6AvIEftq1OubxklImLTMQw6I
32Jxuwlbt+4D5nK1PTzo3Ugybh9Tx21ZELXYPTeEIXpQWpNignCELJLumXlGsU0M
9pjL9wnXQ2ovtZ2jBGMFPZQKSWRzq6Y9a4XnRkr4UvKv6ZC2uu+jpj3AWFfIPsqK
4wqVrmUD29ulDtZceCiMjzNOqYtL5UH7ARlsius30M/XvKomCSEBLl7vZ9WQxH65
5Kg9dzt6t3zPJ7t1nRsG9MMs41q/ZjFQ3VwLV7SpRqHBMbYVaMvlrgPm64lMG2AN
ln5kDag3e26CCc5f/odyPf7tgAxSdQn1lNf8IBzF3ucBnjEDNZSlDx4xIITciN9B
q66XWjgbzPVrHr+Ny5GRx2cdoJN4ySy8yuk7ULpmGeSNpuEj0aUGdWp3t7gm4nXJ
uGHa4Zdb9HlAV9DMnMAvsrqxCSneLdl0aeRaHhByWj/v4x//Tn4fte438+O+SGha
a1tMv72gxKWIujFdFsLerr2I9dXELk8jW/cmZ5gknsP4lG9mv8lEFUPJPkVnEgRH
Y4gwiUwKo0Lx5r9OEGLDGzenPbjROZAl8wBqNglaZknWYYyShOYIg+aGdSCuVbW+
fJ06rl4R7SpxENgGIsJz8gEDOilwAf/L1K+rQdBjC1+yzMRkbwtw/UeHJMmEJV7o
llfWnetpQhZTpDgo1hgAhjhJemwF0XO1ZIkOW+MBkCGwyz0CsAdtjRzTS5XnoXX1
NBLGJt+OzbrDkq7GM/2zoDHUPuAqaSVQIjQISEV/K6jOuLXHNKzWofjoqVkwE3IB
BiEVktifT5UT7iLrDxZEcmWQknEwX8SQdAVLQbw7poWJ3pU3k06Qo5JAQFsPSgBD
920LOrzNJkys1eyyiTiU94N8NoLgo4IPMnNsyrQTuuRVw9WBA7WAzHpE3v6wtd7y
ysFa9943aNdDxJWguNO2qiow+TLg85zd+alHkGU6AnpIyidSd14m4Y6bBpfwVWXJ
JPlxTa1qHa8S3MIZcPpE8NpI8Ds04jmluSuhg/fpk6tpB1aqz4C65h3JdJF09ij7
lIolnhygnxSetwYwicpNSCkI4raGmHM+tJcsB1RGYZFVpFR1J/tOddHhotFJOr30
/zIIQ191TnAmcNKYiZAmfIrcQH3MMv0jG2udR8f8LPTnZ7HIdF/3YbWymj/NwI/6
MzY40QY1sk9sSkOhhbTZtx0zTvB7slgasFouJ9x6EEY21UPm+hACNSPelSnQUCVj
Vitr8bsdKXp3cPLNNv+s7z1JRaoevdNvlFuKhN2onRrya6ap7x6OV4CP2qo9A+at
h1ipdrfe205PFxAQnEn/rgIWf2ZhTW62lRJpvfkUvEIco2zAyUcr2msGCYa7JKKr
xbosIf6vjZM2sJEUdfZCK++SIZsLlM7y/duGQv5Gmz6siHS6xEi26fHDOBtAPrEL
nOdS94QfQCRJR6Sa7IJVpUFWBsQkeHIsfSNwGDhXTwsefSxrAEVPfQqkowvxgxZ7
5UWeB0L92zV97xWh/Ov6+fa5gUbHVDAyuqXQsi/GUeVtUrcGkrV53DJOYHmZxNG7
FfW8VlT1Wd1i7Cddigu6fcikYUG15PDnG0Va7Kv61oUhuWxwZPfCGs0HMbcmm6jN
Bm5PQaXU2tVBw77nUE1tlnQ/clYwOLgE8RQETDle8Nb1SgOJyv7NzGrgx44JFnCj
G1db9i5lDsfw0v4wTqFIuK1vqx+2Q0QGUQgfLoHe2/8Bm0z9QtOEcnhdvzoXOxfC
hZYqk5ffSZzoHCPBdGKDI5LpQ+UFkJmyAZ8cY/vrtMjiLjtRGtM6ojywwy1nUMf/
cYlMbNtBZU84kxa+r+lBCwQPYdLvaZtNmHzgSqomSO22h3aRG8SX8H7GxsMRDm9X
2ZYIwN4bWnSq+qJpaDw3wJEc1sGWTyJTv4ucr7UXo5wzxHDDNBE5mk+hyPOMp0yy
rV/RFFDHzABev5JaBIUuRF95NUWQzjdGpfyJPOsK2LLtW2FHIH2Iq1EOpQFpLv3D
h4b7OksaAybE6IANzLK+mDnriqtYvJzGy6dWhU277c0w/ZrXzSuvovCQhF6xeZuO
0TdJudiqdNN0xUPkTr9VGDrejW2GvVs6RG6EInQmWhLTb1KH7n7rvOpdYLfVo1ew
TklgnYZyJhN8Xo0JX+Iiyau1l0Xn6iIkGHCX6FbwqMb9GNp+o75zxzaDNB1lPAAe
5DVH6poGxS1VdyomMDR62HQU/dFn4zGJzGM8q1NLOz4BUe0uaiyuIb+Y8rnzKa0m
/SeMGnAd8i8O57SMjZCZoJ+hhNbNhe1DaGOMsmvDHnMgFlmmuiqQa4vtuR2+sxVz
6TX+dT7mvGWi6+6KD+/SMTk4F9qT02bLv5K5RnB3xjbA1hJIxcizXsz03l9ZULF2
Bp3QL4vgM1rlRlVfpKYtcDwK6diwHVQ8FsD878QX+sd9qIaQz+iS2wNW9FyUFNwL
WuyxzqYhRI2MoHvGf0aIdWWG0uoiGOMg+LNtoHJwmQqSGJGgEAnsKxTgc7As7QIY
RFleC0zZOyp053CtUgUIqheIYl3iMR9oJyTFXDS++QWdduclZMdB+mg0vEcRktvq
j3YDbXsuDfILDrAK3+4mTiFwGEV2aE9WrtnQnulM8LyIvI3G8I4mGBYH91Sd/awU
lhHPB/LUmcWYzBoAjGp9B0DOlJLhLAec8KLxuVaguYo9z5YCSJnqDyKAbCpFSSIa
RtPSE0DZk+WhfK9d+Z8hj2K+vEbNE+yA9ODPkRQSGIzBuCk72nl5s1zC1cYIimgS
Kk5I3I5mbi10SUBBbaNPld6fUYClYuRucqhZnnou/E/jlBN/FQsnFGLfXEF00y/K
CCIDiVgEwtqaogK+8/QHMmRKRoW1fEBmQVWdW+POK7scR5Qd/Wjf7T5tIvmqGKAH
En+0C3cj5ouEK4RNk/m/TRlCR/2bv6ramI8fY1UBismGh0mKDnM31E4rRGA1n1T4
wniVnI9KjJolGlB8B19C0u6/tBSuwV5V/IVqkbPHpVrfiGkq1OB+LQoqF3DFnJbQ
M2kCUuGAGS3Mc+qPgQWaWfrchPBjS0OIqQ6vU7WV7M/8HlMslfRjIWao5lBlrL6m
L+3iVGz9kgZvX8Br4iwkJ+9F51L6jFE4aGMLY5l0bCvT4ccjGBmd6INaYatBv3NM
KhYRAvt3dmLjxYtKWsajQJG655COZefAo1SmRC8wDLlOS4LlFxP2i3xlfghDknLQ
BEwcFWJwpRkhqpWPWbBkITnvHwO1II+t0aaRwS4MdMTQcjEvfP1ZRtzPhZ080Q1T
nlKZlzlwhc3blbOWTyITDRXWzktM1czo4eDcFFEstJovxO3FAmbm/wqyMBY/cjzq
S4/KKt2npIPe/nPIkaFbhnEv3YqRJntq26w35XmxBv2wLoUTV42g5T1yJ/F5mb8b
1BWl/1BN/RSrt+B6yXoJjGdUeRww6VrwsqLsVKNiBJkVpfaivOHVmKOVqB1lKu4l
nV0k98ib77Uf6f0w0huZUIoRqBGTOaIvjTViWC6gQmrGH6SAwW7fdu8rCN/wX3tX
BIBVxrEsEAwzW5sNA+3Ae0Y43mKnAjXFapLFA3/WZsVeHN+1xkRRqb6zcXmhQQUH
cZ8HMg5JJQjWrMtC1N6ChLKKE43nxeSfD70lZONlUn0IWiIxtpPtWprLJ6vh33nG
d9qNj2qDqKjFZXxAyDs0PiyiUKRygJwV6Rwrqg02uSQOkTTmSS8mbtRWio80P/1X
JxEG6GQih9+6M8aMCnyow1NsMYLPMCIFMikEm91TMVzxAe+AUdkf8RcpkPGNWmWb
4JEOBkGnI12qcSXLKiKv+MLLFifGcjoezBbRLwKJcB3YDVodAebo9+fE3K2RFOdP
+t6TsRqEaLsFInppy/N9TvGLBqc77sqTC/jmjgF+tDhCrXu94clQOAPndl78Cutq
ATdb/zJeqbk5KKRtnsQmZ0Mdu5513eQ3fhER8wmtptCOr0I1SmEetJ8KjRwsmuqm
GnIkOuJOMqL+DuylpdUEConEbNfRZvnlQC8E0Z8SJwk1mExsSaa4TR4BwKtGuHY/
8GCmjUe3Rq8g39rjoDnetSPAYB8GcfHPU08X2Qs1sa/zNjuC1hXA0WlcRXvIsXhB
87U/k/q340kYv22Np9bYr7OXmRrEbQezPfTym07fvzf2m4gVulfHhEssgPLlssie
73sMtWaOJP0cB2x1hbz7hmud5NdiIHuQRbK4tB/MhpFWfHPZPPELoNughxW92XGh
FlDEZdcQoyDoQurZiK4MIYmUx0wSygb/HpDHGfY5MuMXPaxQ2gMxw8gIqGwAoLpr
WZJ6W+n5MeaUi1EV1gD70FM5SeFMy7eqKZ8VolfmqVN6fymnLaCu8HDChbjBLwVz
meVg+1UEdrN1nA9c15tpOSb4NCREhSWkO4bgL6xQnV+GuTa6neSP6XtiJr+SWM9E
9BsDY6eq1NHFzZK24NRRRsazjSnLTBg/amMjNipU9A22BYpYlQzbsDNEfruS7Svm
j76wnFavT3vlLnXUarAvM5x7MXhn5b+SR/I9D2H2icKIMzBfRm7A4AyTg9/kq/EI
K2LhuB28YYwM3LNIFAK97iECWMKrNq2rtTZnMDKVdQ9YzqSEEi8BmHwP9zX0mc+O
dVSRkWGbF/HfPDzcS0JGoFWNrNixd7FIy1+J9OAcKmO1iv5/8h8qaXnVsjH90yQM
d0osFHgb55hLOWEskR9Bfrq/rC/990F6bU4IPI5cR6eBXABrPOIntp3N8tgxFoKn
jsPFSwYowWXOS41ZWEbudTl8q7YNxPXMn8ztccznNyyeZhXNSzhsEM0oiWu8KKVB
E/fl8koXDlYHHPQ4JxyxewYHoahJRJ3JKpmhHtoztXTbmIvDJnYqf39iZOxpEwht
tAUqWFnup1J7f0CO1wKqU9C2e/c9JWWidv9tS7pwy+8TjjUAgIlFO3HbI5epfQO6
Zw/tMo0nYTG20WHdvjcGwLhxokXlppur62qJLL1WO7BAgadwm+8EBOL/v300dhZG
wbVUs4tp4NojQLJu8Qc2O8Ic6HuURMKgTSy4rMRg8oRbux7X9OE5ig4ycTfSXXix
Nfug6PoWoWBGIdFQwzTJzwiN/2LIAr/Hia08NaARikKYo9Tcs5WPTRFf+f4Y3moG
grgip6/EaNiSlCsFh5uSlE94Wh+5AZNpFoEZTKaFgelohVI6BLJXbtVbqmV3SZCC
JlXdgwpcY/xI3Mfldhy0c1kfVwCpPVNZa4K63e3KG9S1rxZK6L9dyYX5VsRrZ/9s
yLqy/x62dIOdRBmmPpzfEo882AYl8L/L47in0jY1eH63AWGjKWXgCJ7/KrDYuYfG
hTRZ1Mfm5oWTbODSyTC8T6xEZYo9vAUmcIwRvXTebwHrtyMi2vitICcHYuaANX6V
fKDWVKyV7xkIIwh4lN+I0Zaz3k5jBNq6Yq2kqEqCw2wgYcuVwOPYBRldrVuuT2ki
P0iPlEScx8SI3TZxYTsEaX3gF+YhKmQxjo5vySjK0QzKo0ZDdi/qMNFYSB2w3TEK
0qw4jq4TJf5xOiAQiww1fs3gVOiv+bQ3HFN5/X955KEcQpVf8kEroMmFe1MzKgr6
iwtwb3A2b4KtqeeJaAFju29XUqjFOX3+vD1YnMssRcMHrHSpQ8XlaD5mXRrFrFGk
Dx/nEBTRoQRN1tdkZ+Ghs+WWgvPB6Tj08kjNQ/nQ/14m28rUzVk7bq3NPhhnUzm/
TtgJFKEMYs5IrGsTvfFnqr9kU/YBIjOG/b5l126NHENgf+OEHTfX1MK6umqLH5J+
2ITJgpLeatEoha4XGtcRwQ5TYqHBJjvlYxKUj1NSB8nEDlA2vTR/++Nx6Y5SZT+4
fI/F/oqNm7y5R9XT4vgA57cf0gcQxCgi+TlpsIWEQMcgyCAZlOPXzAoQltPhziXv
9bQr7MrU71YWi/DwaVVILgCp8d+IoAgIv2eqTBRldZwTleB0tzBBOtYbFcuGOCFW
txdVamLyRYuJsabyzsSkMmN3AGpfDGDvS/zAKeirBc7OnCCjkCqjR5dtC7v9mFxO
1RueoaVFTBn4NLcEr53r6Qpob+KwT0+zg2DmuR1+rOA18S/WmdhmwOgSM/mnSNNb
ceQKOfodcYQyfFTdUbFOi98+PnJfhJZOnHtMPmUamo6LK55T/hbG4cHz02JmIcxx
m6RShT1+g1GWs7+2M3wA/MgyQiC6QWsp+OdnsNbp3EsvoqYYFmZCR/GNXYllnziL
EjaSvidhlGYiLG62+1L1iAZNbapewclsGAd1UcOj4iOo7upOPx+3s2th/2yfcKz8
ZH3Qqt6Ziay1nyO1KgYSTHrjG2aW8RFjTrdvmAFjLsUN4Le7YuxK4/3PXqlOhjxg
ETRBiap9DBW53Rcn3V16kxDKcHUCriQjAMo5Whz2UQrEDXhWqycLMLSH+wBqSCac
kanZb/6xQapANCME8tA8VF63+UJvWAJf9HRK7c1aSJjMAc1fOXyppxSqyVhwVZ0j
wjOLKtTtKNusf4rzoBJSvyV45GclIu6WE4ajuJP9r3F69TXmC/tVZd385veSZMZg
IQEcT4e4/rQAflsSibvvkVSctoY1vMHmgT2LX70xAmwdwTZM4uV9ID8/CvlllIE/
mYwvUE2GGRpwA1W/KGUWJYrAhtDruYzUQGLVYkmP7sQS2qsSRuhCbsJDg9sc3Ylz
ofB224xijx9fNVgEcotSKy8RREn+E/cpzajaSqYmxMHj09hVRjtHfGdYa7nTQSD7
E27uqWChjaVZBAYtlkF9MIx8mcmZIAY9Y003UYbTsFpOIoxYAHRz/xhkTq63wXn1
tq9YVH10ek/UbMfs74+xqVfMh9LIvXweRDYKG+VdMhzNchNmOWNCwKoVgQWc37q7
mOEq60dXKCIk2rixpixLKSDtQ6T+FWTIOIyO15eVboXXm21eR2dKMtnGckMBf/k2
Q77Wr3kKfvZQwnZCDq6f7Kwdn1Veg5pBkCFthunJHbH1VI9tG2nxW9qG0tp6pYtK
kG4TdP/aheJf/+4YUH3gc1w49I/VCha7QCm5tmJfGBfllmBTUCDd+s9G8a8cjUOE
KdwRCRd14PzG9gt71R0EvoLs7QjuE99+BmP0LrvdHmpXn5NUb31tL8h9NgZNB/Pr
BalIu4Rv8nIE+5ARmYWeP1eLo4IacHvmvjjsVdLuGZNeYBxwVzRm0dvFEnulmxZI
41GhHj5RnwgJ+BxOKP2l5g0mvcDhviF4E2JWVuVhFl4+IEWunNBy8LNMzeRXU5rd
EyUyK8EPeD4KNImB1L7OLQRmnh7tYRil9uGqL1xiFOYAvG2sqPfe1PvuxppQVkW/
07br65HDYyQ1QvJleujZauPSk/BxlHcseMxmPhFjEG6aoqA0g1ES6ikLoMiAiSfU
RJec8r2mxs4FLTnWnBciTxGNhimBK8IJorKh3g/FfLc8tDWoLcIjcdarHgXUgS/b
FmWZQyO5CuZwH6QYa1MC6o4scODtKqERqpmqFK7dvaoaemuutfGzGwHhCbx6S1J9
02IuwmecsifiY14r/ExyEiUqOpuScnjV7dXhyExERETNiQ0nL5Nf/uqHr3eq78u1
t85E3KhNplfM/97xdt90cXsjQGJknQuzNB79S9pM+KNnYYJ+wb29khMD5Zo2hJAX
byYyWBF4Kol43JIdhlipJ8GIspcXh03Smm8FzHChc4Ks20n/u9p5dNhAyFw9XjRP
aaVuR6u781IrulPGR55P7I+Z+aFuIAUIsQAkp/2atjWy8YQKclwLerL8+RnvhOLB
qzECMtY0iRaaf8hUZRKhSCDRPcPxEX1hIvhC2aVnpZiZjcpj3+xLwSzOj+ULysbN
lCN6cKc/kx3FhMqOTBjYMSNoBsDwalVFsXOMUMAr5Cwo1zuz7t0kt7vpHMPjU7eZ
Z9mHVUtyED+wodX1u9ZqZXAQxbBn1a3bEhHuQpbguJ9OA73itujEdb361fo72voJ
NZZjQPuM0GVB/wGVOPxblQXZKP9l43wsd1w6+zj5Zve2/7G7IgvEoU6dyhwUe1Ow
99JRAcc8nfz3hPIJxgd0WWt6zx3Xd2WqG4uL3aiHbSq27ZSAJKqnzEtRao9SqzFL
mTqN3wiZVUW3Nw5Dk64zxc0CCuPpwNOFFKWUIByIfVA5uvgX3D6ka8XawNEdEQrI
Sk/9IZdDRt3dcIA7uIxL1BZGg3ssBMH4vMtTnXa1q8JuuOAGadJl+Mbr0EzmNSUd
GCDOG3T2/VgnOBgzR5Mfs+Ey5Wd8rW8OjmE36HvUB8oBJpGQ3luUHXSkKnMlrkqc
9RVEzipU8O6OjkL4YMOt0bdp3JH1qgB6YeA6npmLW/a3PLa5bColHqgjZt46Wx5H
pj6G0JOfMfsT0GGc0/r0+qBoihW40NhfUIZnbOAA8d7sev1xPuK8qjjp/G9tFcgI
/Pja7//XvDE9O0s19G4sX75tLoVHfRQgmRFpQ2V2e5ovywZQxBznictzLfQwaZ7+
ClPjWLl0ihqfcZfZbmOGKBGO2Qj7fXwJBc6ZZ7ibYTpqL6vtB3Ti2hbhD2eTK3F1
u3sxjbRtSbd0ae4WCJsHb2hhiYgcoO+RQE9skfhoPSxsjSn6IKt28U3I6avlh3hI
Fkn/eNreV8Sif2l6Frf/R6BLhtmc0t2yN5ob99m16SyUmOxIs+ZWxRHoOI7MAoqq
9V2dZfE/MUHywUHJScLXIBhHYS4lyGwwAdviimg0/a8MZVsmCfgGX1cOOQ0dNXiU
Xdf/HkhZaHUsfGUZvxhb90wYGnZsEQKMz6BtjpP/carzrhSxHZWipu1mvoN2B8Ai
GKH9fCWUTfSwjTsdv0pMWZVVvyp7vpoWAMa3bg8TZ5HhpXFwghsfNoF5ymhYhs4A
nS9FLdVWEIMh2jIbKnIK+ecW+okhcnVhW3Bvui3gCrd0yYFv1LW7ZWooR1q1QehD
pqJVHKei9EmnGG3xzFRpnx5Ulv+sCZ1/ELtLEcxsudUpoKA/ykEepgcdZldAwH1F
5tQa0YSCA4DHGu0Xgjb1IEuCQcgxWZHsCM5pl4EDlDB+hNLcIT11WQQNXoPXzh+n
3rBRVNSS4UmDa/FphgDE0xUhXKrrVdIA+AN5uwy9w2iNQucZkosksjpEOVn5q8aT
v1iUgWB311r9VpHGkMqLzlxQr/hA5J213U3v/vI6mXpbHBwrZy3wf+dOxxN+xWIx
IuFFTQqx2QnE9W9w9nx8WlLEjNPkiXWkb2d0kPAu/aHIYLvtLkvE4bPsbz2hrBxy
QkHHAl/st9XlmCaWg48571KKIooRGICugA55Vvl7vdbsWRY/fU5FYiWtaVx6FRVd
e5wh28dPOdyFpgjRNy6BdOF5uXA0kxAYGdOn4jfVaAFW0swS8/g+4QqbqYejMHPp
fqCMbeP9s4L+fJDx2g5cX/utpUD6wA+mZgDPrVbsqy+6wID7mCW3txZdzy3GCCkW
daSb42zA9PVWLoMgOAvKYbPfjerpGEhX/1h5djG7gDdY/vbk6Y4GwzpdjSRm3Ma3
nvu73O5yOIjfXiRMPVOGaRjoGjaDZtgwybsKwQw+/KcgB/QTKgnhdRgn1kLfF7CB
mtjhbjl6KuMaxpjL2jwLvoGXHuPvJNf58FYXG5/RAO3rprnVO8GxKHy+0I0AQlTV
cNYbit0z7PsU1tkFhBF7vfvatw8OiKZCA8wtHhehZJO54ka3iLSNnJjhJ44wBiz4
A/5DXNCWesQDtVt5zPpZYlNotlwKWqcSqo5NSwAWNFf2t8weGjZYggsU5pJZFQf4
lNcO8tQCpcv/z6SEKrj+kdT3K9KBz8gUygG4UlML1D3xPxVOI9I6QSZ8/8W/fu/P
XRux9NdzTUCXaZjUPcOWrgxHZXjwk3GOs33KCL1hN+ymnTyRJDtSDt9nMtOzF1be
b3COMSS597kMI1CRNKqxnqy5MqVMMmY5Dm6uU6cRmuoYD+NfXVEIIXNn8444NIvI
ncdCnJOmUfoW4A4B8RnuWmE0VXKsUZqO+3Zusv2lfd81ckkdh7v7xG4BwlHtV9GV
yAg6gTzMRBwY58SNvAa1SjP+NWGll8UK7iYo0NeY4/oEUnpfVM3nmkx1nQ30fnmU
KPGWQXZhg7VFkKkJJrD+fh3AS6MD3LP7N7Pq2anw3VUj/gw5KUJJ87wXIR7rF1Z7
1SVmtGMPbbG9HW0r9j/+uC77O9h0pImreIgOoFC17ctibOCXkL5BRxLxy6aEGj8P
IFAwiJ7r4O/R6VqnT58xgT5BsFJcwObOdUL3JSTrPVbiPHlBZXV+rMy+JJezqd2R
Jnpmgd0fsCKkdYb0OHi98VM1Hlqbb+vF4fh8DrWLy2pQn403aNQN4J2LsyXLEWY1
LolfjG9X6bq3+opN52KcbByqOt1J7bUStbnHN8FqTTFcWBmJmB4uoGcNaSwszXe2
HZ2lwyjCmszholur/7ArIF0Zyx6g/NblL3r/T/a3JVwRuqc3ZgmxSilHTYYISayF
KcxP4SvOLZXaOq3PdLS9uX89h25oQYjkCE1T0or6rml/RlAS8uBtyGNJ6kDLJvRD
GY1dEvL9aJa4RX2O2Z66AZOXLgVswitF46fTGTe1HDcU1DSwGQgqKDw+tMREWKMx
yMfJe4gVoVP8A5BmS9xf3GOe0HWwhOnu7pMKAstnbBST3hoa5jLBiwu+diYfIHd/
wJQDUSHV6nQWRqK9tq/Sq+quGIiLBD4c+MUh4nvDTjlwA8aFRuTo7lpbD1CIcMr4
sg0Pv8pBVI9NQ2wMeZ828B6nNHMsqB1n6C1Ah3UOZE+cfTU0g1XlTn0qmOJuWkee
9PMVUGXlgWXlF38aaOZdW8DOvuaSe9aVIPiqRZKf/qNkRrMmM1GGa7h/HJh42kce
vKxKZ6u7805Jp4oZbQQrSnzeJ8Yg4KoO8CkhirnSlKw5tiUayS8cROzmJxW21kOw
UwiakZ+fGPbMTSdhIHlqhdnOCbo4cdH5gS72HpkRPMdnPEBkP6ZfBmTNhWSRjF0s
zP47ZJQSYIcRNQID1T1oBZ299oePGiWv6RFmdgCA6HswrLoFIpiziwAJByEbMK+v
X9At3NV66QdcjFqxOpfypwcRf7qaOLoYiRgB1gexO+qAD/oxzP9mHgX7J6yinqND
nxyTccbmWiPrLYjw0gwB3aZFeX+Aijy1h6hsHL9oLdsoX8ZKtY1QIdCZMbHmipeu
BPs5iSbm3RxpylVMI0XOmzHnhjnqBJepBnTqHv4+BHirpY4VdW+OEfWCfelEnmvi
IoI0P5XMK2j5PdvWD2L7km0WK2i45tk23mMOEFRp3+frfPBOkMZbG4zhC7LKBYAW
V1fFzOAZa5wolPk6zvTEOwH931lw+9gwr+s0jiQEqp5jzkLdePKk9+jrGupi08k+
mgzJxoK2MjB4PJRGvXcDORIWoUmEdqO8GulA8yqmKuKEZ3etgSwcxPNow1TuY1MH
fiAMs9HlQ2fNlPaJRyacTDztWXQ3xlB9zAbbjOzEUAR5MXDYgjgVmTo5r4DkOWfD
O9+WN22HO4apkzGhAN23+gorf+9WE/bCz5pybN+bIXqM10MHfxWKRYuf50oXoCJG
qhxvMExOGGp5AzLO7/toOzzb4VsPYdJMS2sH54ThF1l3bj+o0Vc7xjUaqbvn1QhA
Cs4ekJkr5Vo6HM2PxA8szlerU+oEXMMtxdFG+Lqqds6iKgdy/CT4GDARqvJgLFwL
C8a1KRpVGsXdvXNUu+XqHVk8SqeYuyPjkOPht7oI2R7K1xh+rXVoVVHTSkp7yQoR
VHMTX0sYSLudE2g+PTpVqqKgfEBlw1POOP0zm7DdDWxF9T4MAMIGGch41VTsKGs+
GXG+sR2iokJ/U1V/7E94MRWcKY1XuGk95aQ1jWRqIAS/KnfHu6DgXO9+6VL9Mpze
Lto+HpUDPlDkHF8MzJSMoF9USnKiDcJeRr6LV/O4z88lzgq1UFP5v3pHbKvy9Cx6
FQoMYREu/meHiZtish/E1jiMS+0t2yI0knwjrW4cqnDbu7fiTi1p7ADg8I3bY6Iz
EtMfSkamXcKdCQ4sm8qEtDxDLLRN2Tvl7k2z8FdodbcZcJN9QwHN67RULZFoy8ak
awkKGyf2AM8yZqwDnwML/CIQ0JEX46G6BifP7XnYXx0=
`protect END_PROTECTED
