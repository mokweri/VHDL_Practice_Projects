`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U569pk0Bzt8/j6ADxe28gMSkj/OTvO8yQVaEszAHz9jIVEIEhhAJl+zlvtd2sZtr
eoybF1/D/Wr0j+42nTeHUJrp6vOk6fEm+mYAtXpgc4ovNRknWxQnO8GDYwArLaWb
W3zikxee4jX3VLCoLYnRfPWnShkv4XWkC/qgS98oQBFrE9suRxnWlsSEwetyhBvj
NEXqL16xWtqyOSY1cNqa+PoO5UX+rGyOvbBRDqJXDysDeU87PCJEaDcgC22bg3Pg
6gdzRP8gakXQ+Icr/qq/uSkWDKw8aFD9IIkG7swjkinMGMEmbP0lOM6Jy9yLi+3B
afYN4QSB94fJAbqoG0u8XdPWz0WJ9PF0d+o+dYvcIGafxqTymIuqBgYONOg9ImP+
tCZffh1Iga9uaZgF9I3ao/c6eW9LuSyt89jiaTDjNNoZbLhg9C1mUkxiYc/Gl8OB
t/fMQrjzUxPjJq6n58Esy4+77hwOugV5r4cfvQ5hZZnA6F+UJD5z+GEY/SlWIzDE
19Q5WF5FwEwiLgt0AWkrGkPtGRPHUg7AwXOEIAHbipFfhnf/spLgKob6AFI1wFae
aFX4kOn+D9HGby5NdYD8j9YWE3F6yFHs/prk59xyMV6zNSlQf2Q38Xw9RJ3M8x8U
4bsNlOXcVYsxJuiATzR8RpvsCxHL1gobgNd7di1PxRn+LtfC+3U7qlf2k4tgNN6W
NxruiqGML+w+a179CR3xhT5B6IVWdPflwJOF6MGLmZcDtDdlgn8DPy7/HapWp3WG
b5aWBS8dkG2znQcmsvew29dHNzgbeXZeE6noUJEHvjqdpgD040PWwnttJjhYwUMK
7XlYH1jgaSxxhbePsvvgelZ/HSn2vZ8OCYkj8KYt2/SJCtm/Cevjxz5fELoLOsg7
kcV6dVyB0y2QMs6IXy60r/rCDfkJ3sjWe+9kEQscFVAVgrQAy+Eu5U3jKPcSmwaH
gqWZ7g1x60D2TbO8B69I/CGHtujtrASPtSFsPF9oHK7XrsdSmt4roOr2ZlyfBmho
VSmMN0P4XE59z3iVy3/j/PDZcNE1ZdGUXR8ofXu/bC9qC0VxjPx0Tbas290owxTk
DLcYE/oxZ/jd1sC6zvAXjZ/OUMmxBFWwLC8vt/7W7tiMu1qwixkW5276LXIVqXyT
fx/qnRBVLlT5aWwpGajOLduMCaxm+HscM+MqgPFIOgapgBDJe2vU8EJ6JI6uDxHF
3Tb1l7dz3rSh9C73GUfdTZBFtt+B6JUyGL8JbXZReSm3Rvfo8afy6p9eK4QTH7oc
rZAF2xox+PvrG8iQQHUfgTvl2RSNq4ZEU/p3o604ONWqtHvD9Hm0UfgV0eNdIXap
/5o9xuTnW6lc2EHXByymMOSlVXiJ85010Wfd0l3Gp/T0yBCCjt6R6/A67YF5LATl
em9ePQwJI0hiayFJM2AwCmjOBBlePGTcueR/7SZbj+onl9qDc2ua3a5dNmBhKJFt
WZ9bJUao1sWYu9Zy2ZH0BSVpj4lTx2ASYpjTdySwFWlWWXB421QqcC3ccH3NUh6P
TqL44zSlDqgyFpLtPf9wxtTf+O9BazGWyGZO5I+GhfX/0PGg8SpKm+r3kBia4hAJ
aikuGcthu+o4exDM0byBB+XB/6AXzFrHzMxfhFfMEDZ88bJnsIc9KGaGzR6/KUSw
oI9dpS4xoHYu2adAiM/uoyQUkAZ+XyXULXpyhs2Mr6CyIg79yIi4UWvK/JJMfAGM
Pylp3TIq+ZL2Pv0fiZW4zH2ctqPkpPHwxYuItdbqfFQtQJLmbo/SCMZNDR5LC9wx
sVmprGfBfAghnqfdaKdrPn71QZMlg9+Q0jZC1O6Ru70B/PTfLa2xuIh0knOnkHIi
h12RIerPhjoXF+nGXd6NSL0NTQM7SI5UktAOcHR/JPE/QX5DCzBZEcjMRX+a60TU
6TjYYZlw2E+Uh6Xv6+9S2grAolbE6HDzayrtWAVoURADwKvJ5w9pfJlVmnHQaABj
Fi9upsXWko0aYXUxhY6rfRLU7SUd5b6NIzHyXaqKdjEeTXNE6ZVvw6P4qs4tnI3h
RUIyNamt+Kj4jBtNrt6oJyv6jqehAoMHPiX+2VflroZjd0JP8A6Z/MTAnUdnYNuG
MjsGMli9Itoi78qzSeA+0sYUr4tNGwghl5zWYAhvW22nFYWIxV4ZFWjvgBc7HWnI
ZqibjIeXx0IBCjzD7WfWbUfmuQpseTTm5JWB1Omm0Iml3qJzmfOLftGFVcpxLj8b
lUeobAGT/oLSeWTRgkgdmytBDauc5fAKweTHzLQFOyMVtERbVP3EyWfCuFiCmPEA
ITZ+CBt/CQ304SjzjYVVkuW2nPCrkGufP0oDkzltftNzPkP/vrQbRg6mxbaLVFt3
eQUfu1T7nLK/2VOjNacs/26DtgFLnhqFhiCLbfjit+ey6ohaWzrOBmFfb5XKZshF
74qefav2hp/XBX6HdzZvL8tK2qlldZV5oo6oaru9NbwiS95oVbGKQTe2lgBGyCmO
yHqitqh5CIKepxn13qCdthwtsREtJJh+UN8JN2pIkOsiDycKjSxY0NZPwV/2ZhDB
DjiZyHKIVI+XOpNLs/lHKP9e3nrBieM7YJ0uWWY8hRChdGJjKzHbTanBOtVKJIY1
pK15oHbcnya01iLMy9sV0Ck8A0pc/n1cXKsEyBK9h43YZkoRryam9oxl6hnbYLdX
JOcuxjXAh7+e23u2FZfYlIlo0FhrRTbOERNNnljzV8ueoWBq8fl3m1oZq00lt7Oc
MgJuFKFdPBjKo3yQUh0o4BKlB4F/8tQjZItNOLo9AQcG1gSMpdwSZyzFSSAO+Ogf
d9I3mJ8wxPK0ntw9oLGcQJ61iubguL3Y3tSy8ezO01P20A8CplYyPpzpk8/RqaKq
az1/bc/Xx2B6SSfgSef07oHbMtCwh9ZEu33VM13BhpyYaUKr9kb0DmsXFEzTjF1O
ISK/b5Ss5f/0z0RBQCuk1hO0oFhptMdVI0Yd0ZX4+U7CEnfxhd/jzHl/r3AZnLBa
GCrt+M5vnTrD/vu4XYLrNjBjRGalC8CAud4vO2SdVX0+nyVray0kVsI970Op3LIY
8c1zvGs/qFca8D3eQe7t465kQJmtm+uo9jlHY2XT3Dvy3ISRJPq/0hl2Ea4xRwSt
lYpA081xxOcaKzL33dgY1DKZ+NGpYkw1+u7vCkBzdH7ibjmTuDO1cnz76rymEtR6
ngVx6qGVHJ9ciqrvUwl9AtoVsxHFGxsrFYA02f9DxNB4nRHfRNusFOvh3RcLo5Au
RqW9x+kPkd8X3dl/eKsaLpI1633njiJephPnHczEe20KJekyuFoA+h8rfcz5tKL0
TR+zznHwCYM45+QJCuiNFqznkljyeQhJOky057Vdv2Is/wrtWzvf5ksxPlDGf2xo
w/Daoz+nlQ2muIFEUx85SDY229UfhoG7qGdiNWd/+CVRXJwDoRpp5JPdTkgEvFHw
yDMq42Z1aGWaYkHZCGCd198XrLY5zyEVdOpFMM/gM1gDf8sTYE7Gbsg1PKUedOoQ
BV8bCnnyAQzAMNkSUrnTAJ+2dcyVh0MwxkWbVJEzq+EZIXbSZAYtdbf7BscGlfWP
YYvTmaqVY0wamjBILrLvCQ2iSDwVDIHR+7R9Lo6Qqwqpbk9/1hbosYTYR54wxjhO
pIYxXUeVniN4sYyLIMJi0MEs4wp9AvTpeetp4/kFjwNcY2GINJbEvIrFaAZFYi9j
julinnSUkYn+umj7pZjBglOFiT3+yHzRBP29unMAczs2JlCJtX06bpApOYkzAIc4
mP1Za6dPCNSdIb80nHxkd6LTrTFjJmV+GK9yGJH99rS7hi5xp0cwj5cmPO4bEerq
4J7e6V8V/ylgl5FG0X6sK/4ag9UnaYW7eO6hH2TZgSkySaHK5xaMLVzE7S+znBel
lSKHLRykj/acv3XSXlV8LsRG9lRg2DW4N2MQyJ+lK14D+uJvDqo1iU3XYw4vtPIx
EYGvixmn2oQXjdceyaS8r3d53fIDQQVzYZkNP3SIp2Yd7Yte7JSomEVk5MLGWw7A
TpQpzSYwo21jav148J38YIMe1t2VFjslI3HXRFLDrgYN4/F2Ik7JEVltTFlqlBqI
/cDpI+l3qLM3TJ9EEa4TejfxZTCyb2IhxFSh5b07qRtOjKMHFjfhBWK/nfLW6Rjg
0GFO+zkCJcJi3V4eJYmJkj9r/zfgLhf05T4m8+V8mhx19kFnHzwycGB1nL3/FjeD
amrfc7WkpMfdBU1+3rSUPpDWhEoViimT/kV2wTMPSlmv89+M34L49738tallpg/N
r+A+EWSUfAKdHt7J6lDsCS5D8vHCcLLkoCQxr5QzenHTaJP3IrQZf9GmSBlD6XBy
ELOmpd9ldG8lLtDxJlfb48uTBtym1yXv8pwLHKmQQDKHXiyLPR3Us3RlmOZ2X5ai
Dz16rRUpYUNO6KviFsCy1wK+HuTIlaL/fECSLnQNQBS2WToM3YOAKyRoqabmkCLF
+f1Px44h2tZKFc382d2iZ3l0AG3hmuJ8vIphT28VW49o2RGgAxAsZQx2qBJIOCrC
Ms6mCk+QR4C2scg4IwP6dniY/LNqYonjY7A1muDbenZoi5RAkG1Fr/6M9JVrTZeG
fFA0gEU7Iji2glmejf0KihC89KBZpkee3+3HmMJBV68kLmh7yjOP9ITtqphmK9rf
4h9EvMKTTO80Vg/fNFRAEFWHJFBmms2WrzPSpM8rTavSPgwHZHnBcql72Vy0D1P+
SHAJLSlappcS0TfylsgE5shFUXensEgXlhX9G09unG9hVOpIYzECumdLH3t7YzBP
AfIiNaQdVdMin+uL6p/EywBrQYYA89K77ILv9FERlK8hRmwB2BsKH0c3Uv7tcXaV
OvJcouKvfrlw2hTYipPloKMkiJGfUH7JBDkD0mBx8gceUJ5MXJNnN2w/5Aq6iJUB
6rDPNT/nlc11zfe3mnTUBe2JYbIkMpHEN7tct9H3nrDZppUjcK1BTDiXAOlZomEF
iYAYND3V6ff+skO7YEdrT5swPIHO7/DKTHSmH8TpoUYNzoHNQeSvl59d0x5w/4MO
F0FmD6rAjJhgACmfizvGKDg9QnL5Lkk4b4MuXZapE8b9q8IidM0rN7KAAbd1SMiL
rhLEUlOqGJNPC5Uedu3cIUTF82PM1wMyRAp+WxwtIXjF7P8FhdTqIV0hPsrAq48r
VKl888TTj27O0doRB++xoKXSEw/Dl2nm2exB2mMFkJgOVGD56s/H/D9JUd+l2s6m
pk5/p4DFCq/Uu0ESbr5f/8bIsof3zqcllKKHSzFjwBCPKbM07OZG4PUN6FmLMLYt
5xajdXK0uaXkjw0K/JT5AcExxHdsWs/frgQ+bn8Ti3xOoeIjEgq9SNQBHRE0AtVi
jBvGUbNTkjBucjUz+a+x4VasuMYRvgEnvLmTrgyuxbUM3L4x2a1bdcqPjxXz/NJh
+Sh30pCB/mJk2fx5tiPVV4bntLIFFRhjmuDQuiu1ZGs8k6+cc/MIedYq7iEjdOb0
y9lkzU+KVYAUtO21tKVTKiq9LQgPRMwfoJUDRQwSHxfoTU53Vs92J5nVKgnvlK+b
5uqBYr8OmHNopcBgqD/SjNd6chJokj6kt0vn/8u2sxbnZ3mXrkdgsUyWzqDhS4r7
3Ask87ujiagzuq1y0l3X4mhDTHVO/7vpUqNc9hy2PLvEq0X6x7KAznhDQCMJzweX
NukwjCEMcN6VKY5RWoBdlU13GakAslgQsy0cAvqUsJVCNijU8/43JaqKHukfm+Dk
5XrASWGZ1Tq3xoN2jOZYkE9hPA0VieUiSvo18m44C8VW4lG7ct9UtdewSk5XFYmi
5uAYxCA6hsG0HR/Lp3zvCbLIdULL2HoKVLWJ6XVjr9W2xaj5G3Wwvg3Q9Y5IqKJp
7Kl1V2aZVxIKqYn4wdOZMVQX5cgwRNVWihvm3LtSw/nfTZ48SYwBcJhy1NCVdQz2
ZCoRJxwDL6Nxa4vXVlhEiM6w5FzxtQ7GnaVmfJY+Jl5Mcj1ogwhyaCre6fReh5g7
RPhUupF2pWjZHbsBPcHOAMJTaFmFmflKmPhES3MBtrgDknQy2yx5lNrEOf1GYv+w
geHllhwmHz+4F11EkEjm7WmhwjLRlUFigZrWmqCHmtHWc8XXlgoyUO5p+7PMuQ9w
cwPr35/LVFJ3UMslrMDloZPHGUUAOohz/98LqvAyUZ626DI+BpZvDrRq7tGlAIfF
A81MmhG76VZJKW7PK7oXQEQqrefkro2693O9+GuCoqDMIoCoHw/t2v3TTvfvQveY
VaM8wNPpziXAAuL7tF8q2aeVj78IzgEhLbIzx45KATbKXmN3t2R+E/9TdGExQGa8
JoNdUaHEwrOlIaLPYV/tUdCph+TG1Ta5pNPtOeLIljTevayAUv4plMmVQ9BD9ipu
4zB1X23V69vanL9OcS6iVtFN1Lr9berS1CLl/MTzvxxg5hDdq4VZfg17rpQT9wuL
d+GKYiJVfdgHbyo5hs7FbEMjhYgesobqwwN6Tl97StvVsVVLBOrNLd+iwsTV25qF
Oq3a/zvrcz/jfeh8iEJH5Tvj9jQsV7uUP3uKFf3RtHpJtlssg+94jO5841B15ZaF
RiAGikgN3vDn6O+dXhIo5VC1XJqy4KWzKxz7VpCm0XjVjMB5w0L41qVcRqezlR6D
GZT2hoGsc0bki9LGCL4dBzJ5dbHbzen4xMtclZD3M93Ip5SlZ/zFmVN4LMqeru0B
HYpb1BmGnNZe/FEXI52wMvlT1/SIJGhnpMZoV9vHJH8WwDkwhEBEFHzhqhJVeZY2
6QC2AFirCYN/pOrwyPegsrYAtavI05bsQZAu9f6pK4ZLeMbzpvlQzuJuyAswcrAY
GCsMpOmje4mEhDRrzZPyUTcu03qyDck0+k6rz5OvbynZbKkgS9LXYCSvgpqmVfAr
fI/z+r7IIphBpDFPDK902mSJ3lU1Uo5mWDXKzPxdwKdihCyTpLeUfYKSpf+tnupQ
LqpIpIIJVCMHCUuF8qex4g3KnHYGomO72KQ1DDOkQa6W7cfMdgtPDvvNE5PSTLZ1
nV7HxUlLCIDgClrqtHsvvq5qCnhMeCSFQTE40JAJloQ3tqSwgpqoh+9sLote0FLj
wpX6ikSz4QojUZlnCwJiSHXBgJM4cEqGtp2/KjiP0UpFPhgdnZ/kNn5sGTjhcRrH
7WKAzG9/LTy2HOwkUgL1BSMJCjf7tGvwe6O3936TWUgKO1LdrD6FUoX9RWHjUbHT
EQpLfXJkMigQIM89cTJDdkKKm3sY5KzGpMzHhTY8prf2s0MXwgMLfx3UUtORmiNt
E+7tiNKYkiOQ3BoQYJntiq/0LR3DzzZct2Lh9c5t4+WRCHhC0ad9Av8m4x7qS7Mj
+EOumek4nMlVrejlz//P4cc27euqo5QHcA+gBgnNe5owOv/ldKMezikhkJsdvzMl
eNU4JSfpHmr71OYQzYlN+QH0arP3sebtceAu/1DS8k+YHQ4CeaGOzy6yY0coJYae
HwpNjb/uNDrBW+Nt8yPEO57lwAbxhjCKEOTdS+zAP7UgU4Un0kFvyMABT8eeG5vM
dbIVA/d003LVeF6NaXzC5WCB2xZ9uvE1DdbeG6/053B+6c7qvOyM45ZDr/vy8SGD
cmcJ6/wDEUCdcY75cGivQcICjq3aKgeINijKhaDPWHnaRd4ZCMR91UJeonzVeCI+
FikklpRcUs/kzG2LMxdtN/3COkQNQBZaF2mSj3WbCI7Sw1TBqRi/Isam0d9oV8Ip
KZElL3sNhMYhUeQmj79unGrX2ThCaWnY7cjFFdv6Wdb2iI7QpYDOfNlN3ukYwWE4
qwmjInZJfVOqLOZXVUl4ZkUU8Fn8YRO3KAKC+OMwDxwEBeUYI6WJ4OVVs7jGXdt/
NfL/sjfFc1StmI1l7oVhc/o+5gFBdMenXTCc5vQI+Gjy8a9W0B5y7pt3Xgfb7t0k
V3FlhG3HqgBPVPbZ9iVcykTYpauurUdtn6xwi4CzRcfvgYJDgzJdIh37F8C3JM5X
ZHaQfI7wE8LSoUYAywGPl54/d5gw4GgGaTJoDIuLin5lYis3TxWAPtT/u5GCNw9p
ZAUeNsXxcd3jwPnp7uM5pl5RtIG85lwEB+5ccsdqo8nbCqcdaJmlXjSIsyF4lVcj
PLeLi5nGefivP3bVwx15K4xBkoElr1p6FY4ieEgpemQslAqWp31THWpzn5raA71j
DwEbEdZ7OqzsBncXAvDQPbHIp11IvwMyRlgh9pnkQ53YcafAGTZ+wHqhSWfkn+Z8
h4CtkjOQ3ffaQC6ZPgZB0vg9Yba9O3DJlzi79KM4NB7HbMcsnILZ9DtbSHqOPhhH
3WgWBKVw+nCveih7/RG4b/Rv5EyiB0md2Fa59GxSn9UuQag0fxv/6LKnpcVaRGe0
Un0EBubf9MfiNn0Bvw6QxNoLfutKvRBnx7/o/qrKdOhCTLUrMfyk20GsgF6ZJVEX
A7SUKcf43w8sQszqE/NyyMXbVFmywd9WUXhhh+gnqG59t+Qk7GzQAYwc9v1HQ+xz
nL+rBBxd9InYRzNt12/bYYcg/54ZniC4b4UwzztCJc1EDSHdX7P/gUzV9OQ1ILI+
56k6o6dja2H5pm9S/XavycvUcy+jWlmys92lyUVvqQd2bttQb2gGKqkJSx81N7UJ
hlhFZ4VtzRC39jWaSrNVGcD/iaRp+xVJv75kCEpXH05GDXzwU2z1Us5ZZ4BbUVEx
OH2aGpX/7wwuNClQyf4reWeIjO27PBQwDqAy9iWpAgGWzhVZxIWJUSXWHbl8stHa
AcsMBLupHuVJx0bBN/huBb+fZ/8vzighkZXroCF/Ly/q8eyHr77x/fWoXyXx1xsR
zs7neLr+35e3Q2eeLJTwRRBkA1hhSqKKkghHiasqeCtKTLlVvTmvqWrqEOl4UbjQ
AVfxwreHth51YQUJK1eKYPj6WDapYnFGxDNJfNt4E/icuhbdIs/hJU4LPETf+mCj
kJ2eMd/Dxb5pKq3OgDFff4MAzI1IWkdKMoSIut5o40Qidg6tTGUG0lw4EODWhFA2
0K/60MinpDOSzpYc8YT8xaXTi4bi5vzaKuApcJ+TaxoQpHjCvq33quLYj+IqQl0u
52FeaVFYEJMGOthgofqpRY/YE0WGPbHlprWHXEFJjUprPR+u1QJmweoj40nCYsow
tKxZQLYSPwSrSXjrLKOy7chDmxN7ghkbngjVjeCdVGYW8CwDy+rEz2d1P6lzx2yn
TAjGNrSFqplZ/uYXJ3W2JMaioDD8aDOEjF2ebMgIRzROnTRahCdbx5gbfF8t/olL
ePFMBbzccjeyo2fyVizdKzXT4SqiIQWw3NAvk0YC9yLcXpVmcN9qnTilmOaQzt7B
jVmZiOm68BjaaFIyRyxNMNqmvAiT4mMEB60m1aqHVVN0HGFVOQi4qs8sEoBblIGm
NAN1pCwsdbC+9HNn4clYkcUyJPZsRIRbVKgFH8NzTsMNStmX6fVViO5fufZQWbxL
NeLE1ENwML7r/ilJPhGgqQ7TVESAGZSiPgc6jeuKnE3mWB3uEgLZUbMvVAe56brC
EN0pBxcBYVubfnjxPnKeshJB0aTsYAANQ6XMybKUclNDwzlsXHXwkeJ9m/0MoDpT
l6p+XIdS2baFtDuTTU/IkbnadH3FYpvArlHn197fnyK8AkTfqDNk3KGs5pCq3OHL
oZhrB6U/u4V68qUTJ+AFQz0W7oiLMvFhyTe7zSNvXLwozRd4EliNcfkkQUxgxxtm
sielyAU2iQ2xKh+b2xDVoqKw2RlLKVuodYfhrO0StebhfFQdPaf2TeFptYdpewPA
0HgQSCEOEH15IaurzKS+8eFx89fKmTbGUK2gLX6B2iWAgiaLfhOEFim+7mVAUHiM
mzWnShz6/M1Y/UN4Tqtfo7Br6kXmN2yIQD+Kb7nBFF2nV90ks5d9+n3og9CVUmZF
8xmtn5qzWCKRcSx/5FrHFSIF3KhhNww43wJ7WE/fhWugGY2gxK4ZOYdcfjYOYR0w
oghVrJtTWuLaTs6UlxamSf7g8b+d5nCeCdvvLWu/IBGPmTY9EHpsio32G/hpTgON
yeuDFSl1oh9i9QbgPhzRxMUEUsCGdrB7cZUMFnGTAlvSvmvs7Yd4RUr+t7YWyR4g
0sRBAnjG3heqmZ+tznE/hIBSE7Hbii4Vwp3Rsl223elKp38MqlgRbJ0u7hbw/0d1
lz4ucZ7uAuk+WeVUpykPnI4myF7RC8vysOwUKkN+mv2iShtMe3HWe45ixxmMgvt4
31GKFWwJzC5uAdbd9ozMz4d4m7gj4risc8iTERXDEixJFGZzFioDzTuKdXBOG31N
BOIDZ3YECqUlMEdBXxLaIpmuWs6YHI3tsaN0+3eS5TayXXwWfsSJYpP5e4TvtNow
KQL/uHjSfVbB/Yyl943NGdLrjBWWjjf2/PPdMJqxPLZTwRL5LlOAoWrxv/qDA+08
VS01hsmO6+T/547Dbtbh4JMHxvE0HqqtgwnKPkcjUL9ra4C5ct0WfsNyTWiI3XEW
6fo5JUQfy7aOiF5NLDbVIDFRcYjjHOukgMN7ovtOGLr8tSmCVd2cFd9VFukx9PC6
CI0X0u+ezx84ruhaN/ArFpua9khXdHoAFV6h5JkIw3iDhfDpE1JiMoG5jzxBMfYn
/cSVq2e2qosb2J3Pi6Mmj2E0sx49tJg4bAcYudzB6uRD0UaVwLlH4AVvKwSuEurV
AZJ6dTyHXhW6UIcvitc5DXFnd3OcXjofFemU5qtEKN3SBgu9169Z/3ZI30A6gj1b
yrpYM1dPzO8kfqfwFwYxNigJXvJPCQfjV2+aEdNejT6Qat5ElsbuCa2/mNaInDIa
wBfuSL7iZLdoejV4papMYmuhz8Bc2dJDBbSJQtOJG71WlbfxmV5pW4DIbuZ6S/B5
uWQShD0yNy+CYR7TYysGRYBfOxWfPShBpghzspo61z0=
`protect END_PROTECTED
