`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvQerzyXtmtTqGtk6uzrSgREKpio3ygI44LdvLK9MNB9dOVAaNgFGJ00+XtzCfOP
TfS6qLzSypXvnO9EUq0CVbXrDFyrNrYu7NFH7O0QPrnjOYJNaL69GWgmW7qei4Kr
pZmaECZbMfpBNPfVZSX//0H6Z3Poa+ut21oSmSQKibKoJ1kczO/rfUV5z/49nhnh
iuyivwRVMzw+JYpTA7U3JVgmcrEcmQ8mk2jcfMf3QxMYyhUzaMuorKybHVmRP9qX
ifHyB+pP57/gRgl5j/uX0H6jEo+kcl6PoyBeaEHU7YxulenMLFueThaiLo10jDWc
PYHzNCf/Md4GIbVhtKJKkIZq/Wy249MwEPx+kzTa/yQ51H4PnGBExcC+ZnSstnYL
fT6qPD3XY5NpiJ7XfFz7CVbEhFPoUnoPoATwU9OA0tsqztRdKag8xk5kOlYBC5ZB
wAPcoYZ8sjT7hAJ6ElXlNW2yhlvTBVtGfN1r/ZHPrj2rwu47fJ483ADbbnulXF6j
IIWaLj6s2/JEUv44Qe7pEG4K/QaRtAAdO8atN5Y/VZhkJC9wjYGYxOnKJkvrw/RJ
5rtEStKJ8dC8qicTgr91UjOdXI7ze5NG0HhmiR5T2C0AJuCcuSOHBN2KVAagPeg7
ZNfljYcUaNJHVoMidZ1AEygCt6adS0AmikRiRAvM0NNm+z+cm1RlXZ2mL6p51W1+
muMfUbOA1sz08S3wQD83MTqopkGip9Kia3iAGolft43PKOIOO867dTgH5K7ClUTK
6F1SWn3NWU17OpbDqusz0SUJBBSNcdLexPia1+kZ0ZN8rIfJvItTkUEqrxAy+mX3
d7raXc1Sqzbnvyn+KBFVQKb2Zhj6MC/DXsH5ocGCuJitTJBrbc6H+GZAGYNCeZ5/
6NbLG1RWpR+bi54S3Ow9QWhKqY40NGIJE8VARYCi52dK9Nd6vU1hjpI/MpSTQlzm
NIE7obdbfl3QmWnEhzeA7Nh1UMA9BO+3GA1xKjXlaolXiVIFLOSTutGzQGhEv4wc
71cIi3L3+SWP7XFDgDftA5mhyQqQbWWZkOdPdCDEaRG4GnNZXE/3wGItQbUxaQDC
STio15KJZ8EVgILQeWPRj8K32D/eEEjAQZu/ix7N0Cur5+UNdbcN3zlHYrPvqHKt
Rp5VxBOvhOGblbkhOC18FsAzFoZSgNKS2KHhUFJ17Q+m27BOG7xydQTS7HjHfyPk
GpM0NHzOcD2oZAc9tZMNW85DreclhFsL49TTJgkeJVHtOJDr/kXVkoTZEc+JbggX
YZsT6UKTzpAy2fIPMJtwd3kdyya+FgCKe+IEu136cq6/KJ2VJ2iuGTBedwXlPi1+
BY3AcKtko++7WY6KtFjXj6XySoT0WUo1f7v8a3g6wEVX0zyfVSBFg0/ftfTfxU4y
SfWuuSW74bFgUkdSrHCSqxpSnItSxVhYNZf+MFQf7uaHMYP6B8XZv3yAdc6uz947
2cUESzZt2gOF/52uDxoYXN2pdbS1sf+pi8xVTNE4LAEsamChOqmh1t6/cR46vP7S
`protect END_PROTECTED
