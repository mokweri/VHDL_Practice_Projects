`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7TAjmtc2zPdEQqghRWzs8plB7PZg4xnoOdulJiEu/hvX7GLoJHKgGIf/nwZ5SSKz
dLvxQIcx7IA56OQ9hNIe0x/ovoYSOlYM27szcX2pPxdK9NQcRHZfbuqty2B9Lc/y
B516moYhvJRxNNL2F+UuxD+vPhX7JtqjdI0yBJSsE4w1wD9SL6b9VoOOg0JpkkwK
OYERRQ+6z/luGmnQ3yeMI/lr+qQmdy5rP81+PRrUJIdnXMTad6Vw3002IzspTRQk
qknrl7aboTHDwcXjfIF1tI3XiymbRanW1akDFq0is91i7ZbBj3xsudUbzOt+cTYP
YRCWmqFyQUlFVPVV0XhiwVfu9fywyrplPEO7quJey+XrZK+jKHcVB1GfkwALEYk1
PRIKUV/UMx4XHs0rqMQqjmlJ67gZSXTn4eEoiQYBG9YrmhTQPIodMNCSgg8PPqFg
gqVRyue2EaoU9TnQnoLXw3vQYNW2qV11duZI11XOyE3rgMSBJ+Jb5Afk+l63erO7
uaHbVALeU8nikwT1/ckCTll3ZE/XapS1Yq0saXCrKCCdwG0k4/1IXEwzcl9zYqNY
MaMJFsGtXHVdugiOzbnAa6fpTiteelcF3C5/2NWyiz7GNj1dikoEDTKEE43w3vu0
IerUqtYGSPjVe8j6aA1kxEfX1nADEeguQMpbeVDm9ET5htCqBhsJhE3gBT9QUvri
uM7zgSie7oLCJBOwXfi8zahmV+5txmMUlAH/EeCEj9bn0imY3XFLTjlbwQbm3A2F
26ocZe1H9A1NysdTMm2JystSrcfpbnt0MxKdMriRhNvvMpO3o9vL+u+JqpKqLsqL
7ySeCR8Ere0mYfCHVLXoAA==
`protect END_PROTECTED
