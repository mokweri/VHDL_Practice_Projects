`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0Ala2kYFqzxKs/9eQzKvNR1NObUBHRLAqQP0zyG2FGDNpdi1Zje8bDKc5hD8vlq
NaXNhSCw5VczLeWbj4EsjayiLN2XDECsXgo51W2KY8ZPep24b+6h32RjCFmanGJN
v87Fq0EdAwtJr5Q9OBiYIYBNnFE97ZR8fa8KcHqag7RaRKk5AShGx4buNehjFP+0
a2TqpmUfb8JjLThMl+iTvVC1+/6Xqrt5L8PW7lhbjmPYNXEzyKRIJPG2Iivv7bNX
iEC5ormbnzD+/BqOV3xfuwNmyZz9iQVyHddXZUeGoes90dwfQKJrWFNzENeUCQ23
WqEUOHZALUJoxZGPOQMi/XXP0wmEsmRHc/tB11ntSEaJNAABkgMMQGjVbYdOqNB/
XMUsb+KgRx5iiogEKiyCrS65uLd7nmuqy/xSC8BbW8xI5xe5gGCcAWdlcQH9cMLo
sA4xyi/OobQuAMqF8SXJitM1++pGGzx1/B2OZjBOk0800GG7F/FOtZ+wPBmtB4rL
Viss5JaqhOPN51GAPw4fiwpmuSZ2VeIBIdSpGoHL+G7mMj9zqlYXeT4pedg5VQSc
g6kVCffTGedl7YKF4acFDvMyeC+7HqbYTSDDUtsBeUFHGoK7OdXPInmTz5ySXyxD
8elTKqMTWNz2ff9Ho3mq1SwFPPVK90uFWs2feYUHn0N7lrUa9oIXPSWCGVn743Pt
GyF30il2Uyss5UU+ud1CUJeLVErb/tG4H1aH+dpyswRN2HembXgBBIdHxpgISx03
z+0vJTNl2o65Sof+8IYyB1F1C66zUdxdhjr3DpB62j5gmzyCwSaIayKOjlk7a837
afto2qgOS/zMrYQvPwu6BblA63Eba/x0Wg5SityaFYu0RjhOATOQBQ5ePNYflh9o
WqTw9YStXhJhfD3XEVj4lV8LYZcIgWBhi50z6bE7I25iZHiRuhNLmCHKEPUXIABM
hualKbi3Vv1Gasju3sLosylpfvEPfdGd9TdHLGG5mRxXWMdTXHQgfhegIMHalzsP
4H1KHLYDyTp9LGTrmclFfQyVt4Qawu6D2FDPWAay0QJMbPBIbZSO7TbKkYTUk30A
Tq9tWNIUiU7oq4D58WOhdQ==
`protect END_PROTECTED
