`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWtwZTQoaqb+ohFcTNzf1Od3eWxTBBmI8Rg+dlvHSppe5rL36ooMaIkh6/6Anim4
o4/pGEMEUwEyrPJL5kUL+vmABTEBZrZj7N9EeH8OnQZdZL6mnuvKaO+TBiS6mPLK
xhdDZtuTTia2PzPOoAbfTjJskiuzALTlMoB2KwhpLsu73ALWYui4T2+PER2blAEm
X24DzVuoR/C6ezlJiYU0LuiUTfI6NjlEscROF9UXquZ+xpuIV80oH/xpjd67MSrb
Ex/uY1BXJ3Ly/PYmx3Bc7HEdDfVB3yRjLoYB6U+ERg9R5bIBZKFD/H5D9sROyeS4
eTyfpwPJvk1O+7AC7DcwBf1ackemPCyrd1JYqev5D7oPCbzoPxhvnu3DCRA/IdMW
XbxFB/U7U65feUMpefFPHnW3mSWW6RORHWsmIu6G0P3lHurFFHLW46JXPPe6ALTA
XM1F3OlJZIDPcoO/xeoA9Hx8FQyV21bAt3U/Q7QE1YcQ4pt0KomVtNdLmT3SR3O4
rK8XWSk8UUzeBvqn57Zk00CCgVn/fQ64QRIrvuaZchMpuyp/Qz9LhEWDiOrrAWsV
MsSUdEuYFwQIMMXwiKChhQE2iXjf9LzFPOnznwUOZbByrEyeMA+sJm+g1BypMPiB
rW3/M/GJdESw3eN0F4M/R66DxY3sVDKKSQc1fN+eQ2d+QowAtV0mGujfYd8ccuC8
816A1C92BkpdbsFsMHLVXcAvbMvImFJJDBHQ4d6DGM+qmszCWKBsJXbv0JvoporM
7uf8vEodc7v7EKYanswkttxWDRnBw1RlHeUpZK851yTMTIccURZeGt705dwdOHbY
Cha6sDd4on4D7JEbdWKAOFmB+Aak+aDygKR4lLw5dqlq0mqFNUzHmpqSbFAGwn/3
DOpwp6+4m2oCY8xNbkGkusP2HwOfYyy/5C1KETAdXgh/wwaObhYCP7R51JtiK6XC
smINHwZTH3z3sShJSz6M9GSpzJsc8gcgioCSw4rj71Dttt9XZEUkEzyTaUCqH8Hd
53jdc0tCUBsYK6Qn7UkJFYV05IvigQ4AO92Sh8zb3F4AU7wuZ9MfBaydQKDVsR/I
/IqpGFBa5qXeoFXRceOOLhQUH3OfIl86nfptb4Xv/L3Dr2HXmIOtcLuMjDX5z6GB
7kxHJgZMdQGwlQ0AwCImc8EMps/mhR8t/ZznfIdeIFM5GhhaSXBbGhQ+S63lx4lr
j3o4iaWWEkunrMk2BWJk/VnCMuWTtZ3yPAPLTcYWX6ta7hkshWP+kGYbms+fUlNy
48QzU8MhImp+cuUoFoWGHrGroDSNISskX5FQy3tuqfFXsHXOdY/DUQpqLtKglBlB
K8kdlpVe4FQjgGwjXoFLVyDDf/kyTUZQIqeqVjSSJ0ywSTjMipAsG0Zi+rDOzsup
QRciCL1TZb28uYFvTtLahkEFe//Qzrl7Mu1j997kEKipsIA7IOZfRy7/qcQyBISh
+Km/UiUXlJuW84fMUWeWmEaZNLEVGF5M/0Yy+svS4Z4QoNnVmkLxvzEQeGzHs+LM
zS+IahaMoET4InaMEnCGhxiw1yZinfigguRE0F2SRt+7ezr7CBKx2Nb90R7u/Opv
kHBDIMuhwmPRPzFR1RxFXhMyOUudrxCYUj9TQciggnaarUoLNPv8U26BFzsrrXc7
AsOAnbWWofigwrEjFuq9dJjaYdYBB1ARrOpspkdOk0kcy92fsz11Btv1icglVLPD
AbC7IwJnxNjNaztWnniSgFRWdFbunC8vq+XUrM6H7Am9d/HQQom1L8hp9RUj2VJI
8qPCh6iXhDSR25FDBIFTTtwBdAuVQHvQxgJHhQq3t1vaFvuluMUEE51LZwxu6UCI
4khFBzhvsw5hEJKjvKqnuHAiWX5FlsFDl28avDu9ZOmxZ5sQij+SAvdewrQ//NSz
GueP62t22L5KM6QnNlAuhjejZCTNjD2dvhSE9XMHYZMXEPUxaJ+5ZcVu/Y3VmAiY
69Isf7+reKJe8HbyiG0bndC1OqU4dsRhx6B5wjB77K/ZtmiA9J6Xxudl19XQXvDG
aLUqavgD9XJSRZzvDjIe7ClO4f1bcbgKjMlo3qGgXFhshK3Z8EU7pU6WFDH0Rupq
sVfOmfnseFj3sGjMwMIxFjUJVxq+ntcsNxjszoHaMepblseeYC5dRTe9evZIypoH
YLDt/vVfYZ5SCWrHYTumWhtHbMcayPP4wMSwt3CK+EyS1FmixdDx902zy2R0WyRS
y+zjKXROh4lV+7wFVYzej6lFbYYcTg9uYsHeWY+GeH1XT9hyKSd2uChq41ZkvlSh
ZnCats3LJQF783vytWUnfbfvoggiOnor0lcZ2M3BLJbIjLDCSttCkveyJQvPFcNZ
4QzRQjlVDQ6qBSqKtFUh73QXBCsnTE0BfU8mGldvKVtyMNW/BGKdHVIPAebZL2nL
Vh4/05ijwzTFtE8IgZgKVPo3ttotl9JQH/5iaa/g6Kv8NPicMGQa1Fl8H7uOW/ds
An4TwZfO5jq2xv2NyYaDgrl0mrqmGvlqiDUdX3xP2Nwv5wxsoVNkNWeehowCNV5v
32JUR8vVN3xDmQDtVPJja1UPIE8tJIQT9rwDQmOl9I+Fk7YLSKL4jx4eT1/On9r0
EkqWeG3o3mar1lJDU+Wp5dVId6anSevZsezahoMOVct6Cb5bm0rf79FKXPHx6Rqs
N3Q/zRWIOzj5b8CoVPGpjNXOYqLTbf8N/eEdud+46evA1TgKZp8OO9n74BztOfYE
7ya0L+sUwyFk+2rprvLg3xZA3zcQELSVHYXAzahK14319nW7RipwzOII4XeagiSU
5N8bFIfTrFshco4ioORW6NReN3DLOiGMZ/CkGvrcN9FEyseIFIEHXoUEqbY/IUkC
Hy09giTiFr0jyyvC5Pv50yidPWqAj5NVjbRuKtABF63vjghtW9kyHPFSq2X8JzMc
AdIDl3Tnh+gNIaDS1/U+aYoOB6CsbrHHFzHIildRuSoMqzCDhhGBJtbD0zh9nTER
c3aI0kDoKI0lIAa+KsXSOL1itcSzBa/Uq7KvHLDGHE4xgmjeFlyKSaHL2LFUoJBh
8Y81GuaYgMNxDWoLPViW2+ZMGQCx+H1/8mWIQ97zfCvz7UkQOQQleVg2wq1P+uDI
d+UUi2oVW8rT/3MUuXNiJGB8xAoT2q8GEs5R0AaYfKiA15zl1HDEqjvCZm7S1jUv
VJ3KejthPmfuirpH1JFXczlrEMFsMym+3ZPBRQDfMGebDQqQbUwPONJr6524SXkJ
m0yFupWxQhuPZwaxmllBiy6clUIzhqA4n7Z4EAYHEQrtEobST//1KRionjlxZDAH
BmiSc3fhvNKQqKb2yuqjQRcUhlGyoOOREvoX7w2VIlYCG5U6J2G35cqB1hLJkUbw
3RY0HNyYIfgp4g/jTZO2GXd9x2SiqW0T6yjukA0pQIkcFyGJfMRnNHknLFVe7O9j
oZotnaGkeXeuuR4EA2KruDn1wZpDGq+C8qhszAWj+vIpgCYYVeETv/xDGQVcbK6M
HN/88mFMbo4h7RcOebfq1WosD/VmjlO3fN+4n3aTjfIle+LwJxNMxzrdnJhKTZ5Y
nVubKZjNvTteQLr0N/TrYmhEu14v0crYGOfsPqXJDEoOhydN2peWl8syX2uaC4U4
BoFecHoGhY12XWuUmer0eg+smxXBhUAwgzYS2iVWL/wtY25sMkr/DD7luPNOJtSu
RbyfIEIDvKeqJWbdnHXIzeTr3U/K7sQfsu11MCXiHD9YDvLsJGMLzaWciS2x45QU
Wq5ZRenJhx3p3sLFZ+b09PoBGEtdHPWPuocx6H1lmMsLEvg3XvvL3KPdgIzNEaD4
eUaocQkviexcoHY3OxpTCKx79U1FZlBLunDyt3SywlFBZOuEibuF5MVUsssgW9qB
IsohbFEpSLGfanfLAYatVDT2NsyWMomMl5xXE0s0xSfTfkfQVEKCWxMOXS8jBdJv
VF2AvKFTq4Zl/r3m1U55G7o9K/RUb6bUoelQONgf4rXjyrrkTsOfxMqGUgkObCAI
/JnRnA5FSymH35wZndH8K5GA7A45REzgEXInwrQKOt0QlUM6RCZE+Is3pULerllg
VFFj6fDLmD3FRv4cuBnxX1wgDyEkIvAsGRPFH2rZEsNetREuSVR83Flx78UwUJW0
`protect END_PROTECTED
