`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h6/h/sv4Lup8NlyUBpkMiMg9boWs9T0c0XrQYuEftEZ29E/W30tM0sLnfckqggND
Ni4K94XsiO1LSD7vKTAungl+RI6hCIcFl54li6+iDIY71IqInHnAFwGT1/Eivdmo
PTXokZ0cVQB8ldrcqYkSQdUd7lWmSJ/Rp6am0hkEZXNfathdYwcP/73OuxMR1l8E
rP5tI4eIJX9k/aj2GEc+aZzGq/EpAs3fKdfl3KD59dXezgp41K2mE4CMjfuhNDUc
Z6nECflhopRVY4JULvXrD7G4FtDJsSbr3wkdqVdbehp/iY+wOW21MIGe1rXaklIR
i90zfgb1Hxsc7EXkXLP5VrJ1iTnF9i+N37N0oDyNnDdPldqdywJeSWBULLrXoJC3
5zLc9Ifa9fuyPa8+AAOyVamz8Y9ccP5R5MuzpkK6d69a396aAG81mpMDK8hkhPPy
sNqCGVtEWh26bJW/MKeZkl2W7FTRtOWT+FCoo6NzFZHPMUsl6gs7Wn/COu+jejlT
Vt13ZreZohD9KSLDU6acbkEypKDBjxMXtydsSPp75YDys7TopHBuxXQGFr95skN1
pDriE1hTLw872A0kWGeMrEGDDBH746kdjo9ZJ75Bt9mecWYFsm5s2RH8RpPiVddg
ybP9I7MdA7UGb0oiJ6DExXLAVDbN4N9xYOWiQZG0+nm4UV7k4jFdXd33ZyFsE7YW
UsLJ6p7g5hKMVeXOG4r0R+qLwQ92Eu2JTA/O+Q1xQNn4ed9hAsDpCmTWEcSrUBZ9
itWGqtYRlG5HR2yjGv2LBM/Y98XAgCtI3yH9vXyIKK3HG8QcYC/KTQGEIJLaBEN/
D2BmWkm2W4qr1A+BNumCGOfVPKPxOZgmnnqnPbcjd6aWEKVc51UkkFBZsJHlJbJb
MDjo8gkash7IopTzjt+yPL9obGtE2g/bbD9ipD15Cf1NqiphFMIO/UaxOUZa/UmM
VauepJ2i3925cjyA8kYKFho2Y+EasMbYU4tdCsZUZOgp+xfV8sM9Z2J4iclK6/hX
Sy50xz9UMVjT/Fk1Ga5GAaA93tPkVxnX9cuYVQ2I++Uy69vDFFwcSqPj59Pvc6Vq
a/tyNZseT6a0t/27P8l3J2PgA9MhaQrTeQ+VA0pWYx3mIyi8rTU1iPRrk/A2r8ME
TzBMT/LH/fvjKobfOZG2bXpygk7JeH6H8M9PhKLZ6M7UM59PKDR76s1/TTpSPUqW
2A2oZZ44EHqzwJNua0eRmwv+2auNC9tZpr+SgEnlqPf6jsyjxrJqcRnLS8fVJw7y
1R0/bFRGIDlf5uRd2nFyK/GuddGKC+N3pUOef4Kq1Qs69WMzEMd4C9P5VIpWW3o5
rZjPbGA2kiW1rbMHQGMoWAkWHXR6g7up77kDJP5rfFTZ4fCIUC/PvNe1WgUfBCcC
bXLb8H6+7vH6KpBajv2NyKy2mfwFPwJUH4Z64C4kHpJI+awZovtnlc9Zd7iJ99ZI
wDZg85Vi1TwC3RzE5wkXjXTU3ss1Gchi+6Ipsb9Oyc/W2ttR47zsJml9oZ3C+Lls
kQu7a+rX3RHLJ2AaHm1l50tv5LlbEiGBbkHMq4H98YNcrLrq9NdyUt7rQSRGFvtx
cInheXbF9/RKDPZgKlk2xKZxe6xQ9v1fWaWfwkL6SgYEm+lptnw2+T6VtxVylNrO
igj3vV3qTs96fp7KnWJUPpjkRmuHbza5X8xGlknnO/fqAtMb0PWMkQOtnMf1jvMr
MvPVp63LPYHlxpIztTyejHagPdqO1lsKh9Y6lclhktLPVPgXsnsJYp3rg5be+7p/
AxyhxQeCT7lUJkiOjq6MwRf8I5QVN5F6Zrk11sWFtHFatydsYPLTw4Px7i6UfylM
mWhNPpY5IVCJ7lj+dXL/qg==
`protect END_PROTECTED
