`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9TvvbuOWyahSTI2S99n+oCsggnh8U9gqLMXmR9uKSVQGv4ur0PyezxouLUaI2U5
G31vxtZgDcumLs764gCX5dbtDvvT5gsWuuadXq8EtcRUAFU59wy2WsdxYUs3fxeV
ZHmSaI05/StfIiRB3H3SOd1OBicYZrqvo6zIz8NjStOYBYdmZmqMOYR8h99D7BQq
9k9IOyFHCMixqB1QBLcpMcjpiGtHZNA8rgA/JZPPcB3RCJmkEe/j8f5bFGgyP7iN
yv4k9Fk88TD2nyynvxxBtleTChQT75wiS2Qfib9gkkFl/F/MCF+8LQBd9POlk7ij
b8Al5PTeqnEeibzAriK6JUmn8RmhjiMjE/CrBb/cstoXb8ZeKJbLOzgdVNN21C5C
LK/tmOdr7YuvHysP/VgdFuW2yiseMXvYvRQHXaYxfQ6xsfxGTIufl2jpsulMiWtu
2kbQuYv7h1h1Xx4e2trHWOIs3B5LUsBJMRoiXHkmyqpS/eU/WU5XIj6Cm/HpLIg6
C/P7z8FYRcfExiVLEAkaF7yFTMSHHRaG/MtPvrsf8uavPz0oO/0Uu5PI6tVEv+R3
FwOMrOO37G1ceUSc5frfqW3DOZ746KiEAWgDKr8pmiypg/8pGiAwP2eA7jMZ0Y+L
92v9V6M5Z+nfDivixw4gAm4hDQE9kaX5Qkn7Al5EDJRiMoNPuxRYFJcIj2DpmlIx
NXigA4SbwZUBVeqO6dCgRa1M1B/OahCx87c2t0zH6aHqrrNYW+nPS3VAgCiNNT+u
Hcy/NlCxuVeDjbmg8vKYAJDhLz1R1IJjpwNxbkBzX/lMxY2NJbolOpxNKGxGCAZW
IC7fUf7UKUvqfic90kzttQ==
`protect END_PROTECTED
