`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KfFDSm/nU/SOc65Ylo7H4/x0zOysen50CIsRqU61Wociopd16Wj2jzm+gnZhCXst
c43uD9TqtCPEcgKnUY1t0MmUR/bCV/UWkD9j3TUrvlEDDHXIpv9HyF75gXZr5dBQ
Ga/4egS7L3vOKFcscgFqHON+PXAZ8asO0s+G2IzPtSP/iJlaS+kdAmwXOprG4/Z9
91PTb7hidi6lenSk7QCfGFB8e3sOj6e5vT8A3adB9LHT15+B5j+9laAJv4YLP2VB
em1gE/nM8JhT52SAemAcpiW2o81+bV+9q1EJkEc1crJBag684/4x+VXdDthBi0WY
F8C+Fltubld6nfIltKdqMrci4DuYVygEakyDvn53zcsg/KDh+awcZol4dVWxnsuk
mVz6XHHhZgFJIJyDQU54o8536FQoNadeAFg6diLJ3kN76Sp2PxmHrVgQhrhHsn7W
cppcRXrR/t+JKItURpwnqcugS4wL05r6iBtMcBTY/66UNe+Fee+9Gv0mfXBFgBq7
95GuVNuQc/nKpzPZL2gKV4YAGrM5Z4X48q13cQQiGXYkz1/9XVPcQi82fJpIfDXd
3+84ittb0psDX5iwrOvFyviPKjWqsGrh7jTcavecKR+DDXJvSfA8IQVIVbcAGKPZ
mqqXOaCeUtR0X91XU2sM1FsD0Y9RQvLnH5bJKRa871skF0RjPjIGV7/clKP1WTt2
dd1LOAbGjsN/znBoZ5SWypuUpdddtC6EoG7282/2eZIKNeJNTzGZTIVz4Qw648q/
4cGHfpqPLNk+03eqsnpjHA4MDniw8+RHbnbuqiotLzmKEUTGoTH4U1OeviXQyq1S
McFiJfYdTrYYCuV6rk0ETg==
`protect END_PROTECTED
