`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GA/FAsgFGPxAvrspCx6fn2QAQEYmZu4cR4tjjMkmUS72UWE/ElkavtnjSKNeuBQJ
fPp5jO7Tx247Qjdq8C8Yxa9ZngT0e7GEtulSAwrt0FbKUdzNJoHSRYyEMXfSjNRA
LMYGceInaAiGpOxyeWTXO4kZw6C/QzQy0FYUajVx2eSpI8AwCq4i1RvKm/nkArRr
VMb/IggyvYFd2H8ysHXx6gNz5mTpMN1oluc0ZYNUlpzOFj0rbaTuHP/5vTM/9cKW
WMSkiswV9rurd9Z793OjY5DLcimYqSIjx/iYEz3HUbEYkYgOILUprnzc8HMOWRSe
kzzxfltjqshFmw145Raw3uxxMyrFpnUd+DG/AkGWvdpzCTqY7Ag5ubZFRZRt3Cy4
Cc9bKqG9PaMXkqCD4gwCkIWVwZzI9fyQO6O96/VXr89N9w/wMgKyVywS3CPTFAGh
iKKcWxcrxgfEEO5OgZ4J1ee3puLJllUNNjiqTtPQy/KiIKsbO+GMEMc5fIOlUZ8Z
uLfA8u87p9y/16Di4r1FY7OgvXhp7YsPXM2xggqt4xr2BshMXRGDHe5wXUCP5DVQ
NB1hHtC9Ct6mHrxViC4VSK+e7622YcIZdq8l994M7VyzusTH/4KYSMxqXSePtMk/
FfsxOyt8hoNSRpaf76KvDNBS2AWPsNZ2Tmf/fFBkYo7qz8dKI8Ogk21pJeBcdlNM
ax7fZOC38HWU4k45grD512nWKfjS4fWsOrSYcxd3vjPCO8LK2H8kvrvYzN/59/+7
UBN4WPZedMYtg6iZl7TGnE6tp8qpqBVnTWnBC8DjjqPDxTlJ3956RALCxiQxEmDq
PDFJRchbOj28DLyjSgtmhnOmRTyMK9UumeqfyhCZrAkjlWM429753kuXEU3HbNvc
Y5EpVboM7G4Du5TVp+MzuPdIzPINKuiEFZozSohC9J64MgCW6+LESHgNKixxzBtn
rAcnn+R10E+cddP3NnW3njNBPASDnu6S4eLhhSSqc6kj9jS7MV2gkBGdZEvEpHRs
lvJSCzisQaAe/iHov+92boF6tppY5YoxrrEbF0kYNRodfxchKEsl953yiPG9ww4i
rfYcqQBCTRlLkgl+xRbdWjTNTesy3crKenap+2QVxNDPyLnpkMy6jn7JL4fAAicH
y/oIQdA9AIY/HiQW4biIiuxJqieMBmUbkByfeV05roAEaSmyrrSonekZBW9Ymb8y
mnOi6onsQVg/lrfSfyJrRtWu9CvMtiaylrzsZl31lE26Ez9Ej6tMlzfw6s03079L
34XR7EwZZlyUW1XzH3QAwjkSZdf+OfTdawCEkbJM+P1cizg2AU4meP/+xSZEri12
TJnFnAeiN5YHGndtjPz7PjEXUD+5xHlUGhow+WcEloQg1gVfyFZfjx366iyBso5k
+UbWbOn1sFtJzqe7auAj64+S/cbFjI9vdJEzGVWunCZj+VRC0ucbESCpK8DYltTE
C8HecRK5js8y38sp4L8+vcn528kQizAV7cn9vkNPWwuEmwTAxygp54mEi5i5QAQ8
1O5f+XAVgVVstSF8yO5aybyNeR5TkfstyzPlZ2OsbmTEnPo4Pd3wQdOaiZs50+CX
xvKiQXFREoQUw1Ye/BIAJjkIha5YwFYug4i/HFvBzcUPMfHYnLqFIo/IsRA/ADBC
xe4swvEJShQjku4hNALnA/4ZPoIO+5M5gUTr3q4ZGJe4JpNriv3653cf3tU4WNv5
DqGmb6H7cewUeXmaSc5tFq0d/RdFOndeRAsnHvpTi1CptAMq9ujidOhxICmJH9ar
lkp/gbbc2/AEXueerCRXO3cuNyt7m5trlPWuZ4N1PKSrFSXbghNtJ+UT+9IJvy80
UNCA1FFbhG3RZyfGZJnkHbpbdxMvWxkvLQ52iTcD3TRYr0kojIgP2V1PY9qK81Xh
LZ3n/IFVfNb9N4HmpuG+zZ1bGo87kb4Bv+TftfjysSR2eN5MBwjIrnuVadxEta1m
aj4m3Yv+o7heoLEME3DzLP4YizIEyBwzUUItG7rkT7Lq8u28oH36FyRSMvWDqjwy
r0Pb8Bl3BrZ0hf1++ubDFlmdRLFw2KnplmCUUYaHFNwMYuyBWys5RWyDUokzL9r9
XftjsTn5QbXftqA5cC0Mc6v/5DF0aQcE6cw0K/evcHS7weeYL1hiX+XkRydBOvi3
DXfNczyvLJdu8BBbYnR25mrgYivkIP5aao2oVyWKdQEoaEU1NleHNIn4ScAW+DvX
xwesJFJtMwnxJczmmktvKcYl+CDaSTrbhdWieAGRgWvbw5JAf5FxpLeh3WbpIwAq
2aaBdshpEqOBJTjri9kkcWTDDVIBuQDQG4xNox4BZ8k4Dwtw2Ey+sG28kpmAgalA
nY5X094lo+x3778+sVOcmuDWZpthd5X3mTC99libDMbqqKYK2gIryj/wVcbeFaQ6
xOjs3dGk+R1ZV9rwN4uD1lkS9JxfTmhNIinWMb/ipLFkve7kle7cZYwQXfW7r3ng
iJoyuZXLsZ0935JLAaqisDMuvqnd/qNV0qKMuPcYKFsbzU+oVYOF9tzapImP7oi6
IhsmsubWeY0us/iEoprsCX9rOAbEga9Iji89FaxgdGBXYFUIFj4IBg2VvNEvkA0K
dSYxM7RWYzrGgFsnqV8fmjeKNmICGOME7nDz3CiXaVkJRDZwPOg7ecFlEq5QECbY
XiWqCsTdHKMkarAECxDnXJyJ4UNPZIprKwJwlTh6/08vd2pXY/HCv/x2cyk9ySuA
MRNpMcUMS0Ra3qKEgp7nGKA7nFYkrBn0ayqN9ao0fVOk/WocGNhBCUwTv6qNxs0y
Xh6wpMNhHiClADnFC24qj4/kr8ae30/hSf/YA2Yd0XAOWlP9qaG7r6aicu93Uyu0
G1NA1U9ycvFHBQijC9HokrQuwpAPqP6LZVQlYXus9o2YWeVWRC0QSXN/5IQW4xWG
oFhyiH3qTOn71Zvab5JkK3RoQpnVQhgJGS2DHkFBsMj8EqpSPheiPmEJomFKyc9v
W9UjE0hjaR3bOn+ZH4hdpP2HDkZICMGpVSQ1Oa0/ZLaPBbDbIzRV7Bjbz/fe2bxv
dDjPvbvJ7Z0qCQJMEa0/WbxGxGJG1sh79f5sKQHmXGXgc2IOtjGo3LSpdovyCQHD
Jnk2zfyN+e9uLQ6QCHBBGKc4bl2GrWaEUdKdI+5iMhLfVaeargxDeXNGe7/nsYJq
8dCKebxpP+s7Pdi1CGkqA5qGUivbieanUNQdu+VBE7O6B2IbSbncB/36/fTo3PRH
VDrVLwcvUKZ27olSi8f/a+dJaaWJ7P9XpVr/7JCq9OS+IdsA4baKr7e0bzJV1gHS
iIOZGf9dcdMackr8nUiVKXyduni5Xvt0WfPZy6Q7KM7v861ditaEggjomea5wwPg
Zc7J1DCbxxP2kf7yZsN8lgScF7Guy2w1LWhT7Ixl6B8B1J6L8adVEzSXReS07/I6
h7pi9yw4hyYnpEOcIWuS0j5kM+BDyRhsUKSPOJLn5eaLW4RohGgM3cSjY4Exhx2q
/Y5VNXhjwzMzub3EP28EliKAQzVLqjzqJupu3CauM+C/1v3mKu8/gGD+dbXYlg/w
9TRPmwg65BLVTRWLFS11zeak85787wziryNDGSk0xOULuLIOenInlV3POhq8p6xI
5AdNEu2YLuyDrK12OVwiia+r+kDfjkdcxlB99klAovBjD+7EuyUSLl9zEyHhsMOi
ShnYAaWRW5/k+T8PrXAXNG8QZlNTJzQkxNG7UQp9bACJJJOMU0VuQXD32V7cmJa0
bawBaNeFij0RO9EwKeT44MqLPU4VX+eqN5Wz2mu3BPCg9m/pSESuz3K+tI2s9DCB
0z/8WKyjPERNWomxMYt/yw==
`protect END_PROTECTED
