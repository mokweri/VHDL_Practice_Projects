`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dimu2BL7mXZIXmhqdx6xlnWHWSLT0ZFrgGud5r5bkPYDcwPFSj3aC7tetty8jLpZ
xROmpRbofNTv8MNROsaYYns3bbbK0MN+SoTA9WnrD7ELW2fHJ44F3OUaIfAOJM1r
UCr1OQr9FWTyBX6QvWcVWKZrMOyRLenlKGi2Qzd1KNAp+ORsMR4cjPF6RQA7cZwP
Xh86okgU9Wc8AcL/5ye40INQSo1/UeKdCOVUKE1W9QO9OspBgMjgeRTJBUsWSjAB
YcVyFJ5b4h95CNaoElIO9F5kIW/N3VYb+H9QJQ1WamNYmNuqhp4OK2tkjumdIVfn
UpgU0ILc2tTO2ix2IxscnDM1PwA5AUW6MFyuctAzPRHLL0Elm9oJ7gCaOLpcBo+U
WHHKI77KNgpbtvn02kI8iDhPioH3j5BU4fEu0FbvcHxT31TH2ac9c7onaUIdKlWV
Y7XWmjHbSymMIJvhdlXUgaU0ZNJ4k0VaHW31RTVtR/+22+F1BI6xVnuuM3NQltXD
7dp4VXGTKXYJwtyWeyd2j0WhnEbBLRo+DA+s5oYrcv3m3tB+A757zsqesLT0CyuM
rfkvHqwF5TMp1UkRgKdOiwWZqpJdWOg9tlrybkomhDwGJnkE9KjROZjwH79Lx+dh
YYRgOeClfeXSmPCNrBus/9+m2IEwwdRv23RHL36UxhNgtOVCj7xkIt7RRlTKf5VZ
KiRUjhRPRl+SCM3bwdBfZCnivHIYTpAWznaksBOzul5EcuvbnaJ2PP43PF9DJZMW
pcjzCeNEzQDZxz+brtEJf79MMJ/57wEvPfFWDS91kN8JBj6Yknw5NSNBIevDmzAZ
wWMX2q6HK60Ti9XKbWgYflF5BZTNH3RmcltO+vvq5rGeaJ+dztt+/NjV/658YEI9
eDwvbJADuYl4fNCZ2nlnd9r8ij5RUz1hho6BB+oCdm+oz5mmZL2E9DJ9X2x5Q0xa
YTSyN3TK7xcZdjmt5Ix5tjNnQOoR31EaytcyGu69zVGrOH3G3xUjuULA5EpD9RRG
PZUPVmTIDLJzkoF6Zvj8VbwC41IURxgxl3ouISIwvJMmdI4Ltl8Tr9cfdkp8mWxt
8TkZl1Zv8qTUnelQrtXUrunK4yEwP8G1ByB+YooDiWy8vYiKDFoX7bwJTeQ8/7Ba
87pzUZJWeSwJv7OQq3vFCEOBz94YNxdVXv4APWN5VdrbCBqsk6o5yT0jy1x0l788
Mpax5lzGAoZeJdwMta+oVY8PbBcBK/fumeRAtbEoLOk2btxFuIUrJWNnE8tg1j8+
g3ERKTmN85asdARK6mkUmnRF4i1HcQ8+/py0AaO1SMukNSk3Z7y/xoTUW7L0qptK
gbQX1wZ9MumRP36T51wJ0E9CsN8Fzd+NGK54bZ26kxZJQJbjxfcBix9QbYsZIzK3
3c+MPVs6z3WBPC1yzcfco04i5UGcDlKObrQ75zJTd+hkvQcwJufKlTCCNly6Wgog
r4uObPa/40PErHKdhG71v99YOLX2PeFBKBWOiHYm0T+IrMmZDj2AUp8da2jZcorg
7nOVfHV4UL2XiSB+mr7T2J2URkWaJrLK0GbBiPmQdyOJIsrYOrAU/S7O9M6MH8yl
K0E6cC8s/p0rsFai6HD3Ab2HY+mohtJVcRGctrE/R3itZickh4D4O3V1nVdrrMcT
EUuwPrLRL7FXrSzcYNrRDAWzH4vQj9VT04s+WJruSfYhC9V9unNcxG7FjN+fQ03K
ORmM5d8PYuTCpqCuyuUZBOJ40D9r5AIEikPK4OzvaMs=
`protect END_PROTECTED
