`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwbGWrcyzSOMXHQVeoNNckdsit5cO92H4BRTkn7lHSr6DGTlgN734YYLOdZ3oXFA
kKpZRQ2JbeeM412vhp375cL7zicBWinmkq5nagWyqVxdRfaQB1yjpSVKdTYjR8Of
9tZDosEqdZj1T0mMxhLde2DvCsljkLbfDHU7O1iQO07iH13JKf7cjZ6f9RfQLlNS
u5tQLByHFO7ttXpCz0mwZauR8KRQY66zKfIvK3sRyyzXQFdHiFoSNlfK2Yy2Ygbh
REvP8ra7BjadF2NErAvaqQpz1CxiQnSIc8gSrUwRu/dkviDMvPGJ5HiHqO6+KsFu
IIXIwCVzhKUCHR6GThf2+FiCXkVNJkirhmbLYU/2HIJ2v9FMJv3EsBQ6Jz3YQBEf
NFHbYksQYomjDAzwJABdZEdktObLq/Nmh7CmNdY4FZqd/9cEggMN+33YgP6VCnlD
gXZdKn+XI8wzxKMBLK8jytW7tFTZfM1DVu2vdacV6R/v7sjd8KcIU1uI0ToRgJyC
segEjtyPir0YgZfmakJIQGTujTHYj1UJCMf48JeNuHZfSv2OUUJHsqrWzI9bglmJ
z2GHZqUuI3eC/k6DTFA9USvsSaB7Bc8eFS7XWG1d0v2F+/g0wDlYZlNlowTDOxTe
IobQQS3fDNlR7Ol12qToBxZmKQk/YB+naSmWeZOtQNj0/wG5GYHnKCZg7j6XoErl
rychAfHCEirKUDVGySiAuHY68W4eEqIrGXHtd8bhUvb8qZth1A2ukFXNO3ZACPp6
Z2dgX2ntKkKG9kwoERrVjdWZcyCr+FXVVydQmJLsc3tcA9Dq52SXWqDRJZJBW9M+
l8niM6AZ5ZtBB2ObFljtfM1S/QBvMKI6Womd0ttNt6dHpSg8snyR2vdfI2YP3uYz
GF/KIebq11dAtz3Kvz20JEYizO8BK6kQidHk1LVPumTFByGUoHHnn6zlagkURIeV
b4n931Z+NswokabBW3uphccBHnuwQgbzE+mYoCbSO4YySNCVKAUz63XnoXk9HIwD
h8ED9Jc0MidXEQJ1gYJJFgRkpOd67Lt8JW/yJJMrTL2dhPe0BfAKzV7SXjdcEgBs
AMzFhHSXb9Jv/5KvK+a/BXsFopi8R6fJqc3xGqbhxDTd852oDPybQIUJ01hjVnl2
Qxny8ueLhB5JATxDqnU7YfHxgNMeGDQl1B4Wef/4dLJJ79w5FXgpWIjNudxw4W6s
rcgP7n3RLMQMxsAG2A/fA23klveFj7ZQ7a2/wTLKfJHH0/ZHwAh+ZjBXj9NY0T3C
KRH60HL+O6TK0Vsb2c7ZUKgexSYi2Erz/7FFqIcp094IGAEX0MBO2qVr4DWqGg8a
6pz5MH08AZ05DNiGUFLRjjdsr5dcKNwurvIBmsKab9uKKF6B67q9A5x0rsMdjT6F
wlE6RSOXrOaLlNCB3yTg5VV4YUoXJGUfQO/yo1dTO1+ik5HT/FTYDpmAJ/GuAwr4
fgiIkeGjuS/YXOLUK9htFpeZWJfxgtr72a9Vpiczhu6l5B19sDZ9c1Eh2DoCnCIk
3U1gEVPGPyFgCQ4R8a8Q3kIe73cqOUiD0lokl+KK3q/tao2ELk2Ykxb8MYHDJIg0
4W2rJtqCtEH0xcJX44r52m4YDYZYa9CobbY5UxkN0oxRShBAaMqHBYdze4ojxkkn
dnQYEWP3/5k8VBRhWy3An/7YpLD2HBamxD0ZTDLUq6x6FsDJSiOvZuvp4ZWrjD6v
0DRAPVLzD1qBz9GCzX+xr6lQtsgQ06n8mAJ3smHgW3Dal68bua/bUAAW2YRB2Fhd
ht4BGa8hFEDlUqAcjaUB03furEJhwz154jtj802j70KCR3hx5Eaad7609NI5SW0P
0sM4SKnk9Ldb3fURAUggAsFCvD2yBxkQPQcvk1ogwaZ7oBU7WTgVde7Tcz3Oo1x4
P17rfjFT7geEToYYn9wY2F/RQgp7YbvD6pxNQZFkXFGNZCTl2v2cDnoC9spDlEXA
U9FVRRQTPUThPDb8B1j1cr9P+1Ncz9Z3UTyqmqK2f8Xvfnepbx7z5dR+IrXC04HD
UChctPCFKxW9S9zNEMplpK325nhx+vwIBlbCGgc0+xEOsvisUFDtSarTbnxIGs5+
4z8EkWdcpKR8LoXrqgjGaQkl/OO1RvVzxN4qrfVR3Og8SKcp3Z9YQfqGVLPXIPVA
Yjcre8Si6Cg7A4AJvMRRdjtjtIyg6PVT3jpMXeXpoHU4vbYvBARb5ELSbB6Sm//T
d0ORJ3kDbrM4PDFYIuZu63VFW4VPPcFg9mh2i+tMx6+iup6bMPsrTx4NpD8u8aaN
EfPmIOUFJJBo+0scfSV638GDjdjqYkiU7b5EQhb/6EKlnoBpOwlBJXRx94u5yEaY
bvvAKiij4Iix7tyTbSn+/0+hx01YRHfBY0OgDlXCcRDLRcu/HBm68LDEDV7HITZE
iqUqBGPtkcIAfKkjM2/NYsyEad4sFImsR4ID9eymMNhhjW0Vy3Y0eTPD6MJWcvQQ
eMwm9nfpkJVJqKkW1S1rNBOEuNMeCoiD1Q8v/q61Hdf2dFZl/Vs7d+4HWeWGWRAD
g0CHLBgvfgYf4F6aPJj//baqCIKO+t0yATdw2aPkSX/3rPIAxIeVDg+wEkyawuaQ
kzEXQOLlCxPKmN9oVXGdIAF/6Pi4SQc+0DO9DljTuiutTmDc1EBW1fORz2yUr9ow
cA7tb7w4mz7cCwCOCWYcViJOAcIYkfpLG3cH6NMWUFu3KQ5mSLL4JQGIyeYZuSoa
7i2y2JwRoVio35pDN0J5lM3a4T8W1yDFHCzNQlH0HPLFZvozeygf0QCEoNZRfZaA
12gWqAzTiN76FGKfcLU03t6+lcVlgAxAt/kQ7qHkAYuDCDJc17N5jvGX5k1oam3h
cMqylPpx5r9Eow+vY2ICUbCd4kGIiL2LdyV4OSivkNCXnR7AZydStghXYU6gI8zz
jPeaqQTFCl7n0eW1OURBv3zt2ZoxeNv5x4Y7EPZ5Js0dfQpRFiVwZT4+TcAZrYYG
2wIWV5lwvs4sd+XMaeUDmLuGd87swjW4S35krr/YocrPE1ZW/6U/SQt9QH/aq/9H
ptXGEk4lVc7DPfPq43nlQO48U8mBu8kiCHmWU4SwNF3QfsOMcyMVhD65UR/LvhLV
sg9n2cLKkQp0BQM9S+Di00AcVvshW4XVb7eoYETYxPwstB4Jg6QuwpEUi+fik7hU
g38x+8gcIl4JK8YX6I1c4UNzX+cRyMZ3K2cm1qOBUT1cjHb3Fj/xWRxzamu1u33E
c88VLvL0yulKVxWns2d4HcZcyu1QDmnDz+dZclRfnRJPqNn3H+9zHJjBgXJ3inVh
I+vVyi/wXUYZXDElW14SP0MWujghH6cfDpj7Se2x6SSIXhQ3J5fWHu/ywWkTcRmE
NQgj96hxMsQc5zuTax2WmKqWwfjYsFYTGA4h0j7/5OqhHGE5EFdrwLQwHdAktpVC
V3sZ1+2lfOLwbtw7ohyGWv58mhc9UoooHruMg1cMXVwUMfKz83M0Me2JyOIO4ab3
tIK3LQVOxwdFCMGVGP112nXBoV8QB4OnJLmB6oh41zpWh3y9ig0IBOM4hOgz1Kua
4/bYXPWq3sVySYHaUcB3b5CZidHK4DkUiGp0nZ/9+/u02r/M64Fc1Rg1a3CmJ83B
QAT015LaRYdfqtQoRfa1s2hHvzzLhLWvIzTimwJCIHMDOz7K1CqQZT/vvDxRGNZv
CNzYsN1UH4paqb6e9WqPDKNjv4uGfhKe18rVSuVJtwmtkbfoXc6c2NLx/bQPfnAO
B38BsenA6wJ2TSZ+ZEanQJu9alZvSHHR7Tt+H6KjQRGxDJhStkBKeN3jqmiTLBHa
MSHJc03huEasir1Ngvw6ug==
`protect END_PROTECTED
