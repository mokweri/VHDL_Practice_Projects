`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nrjv1hQ7MReUYQYhzaPkFBnO2+qPKTYg/tgp5Rar1a3KyLz/gPNZFgR/aE7Vdpo
XGZ9dWW+hfmCMM5iWoiOgBaQhee4Dw7ozvZ0q0nme6+gUNnRjLeN06UoE2GijU54
1+wOggSJbgpc9TGRhaQfexbwznpJ1k9KR6Z4xHh9Fjjhazz2HfYGJUwh6FJZkdBS
WZi1yFq7RH9k8SR07GbUIsICE+wtZ+jt09WGHeb82Rtp2xWvSROaulUu+l79MpMN
Br21OUcy/pdfLtzFXB1FLPbfwh/32LtUcy1fPIw65OUGME1DPnikhcQG8hbqzoqq
SJZGqM8gfjElJRuoOwrgKvT59FixNlwkMnzhI+8uKd4YA16NOC1y2k06mC0QMxNT
31FqmIk3+UkKGRJkZXmO0SQoItTSHbeiUSyNDfSvzQt73Uwuk+XASvb47KXWY6pR
umvBJwR4aLPQCpRy+oXusip+r4vXp5Md3t5+OpaBjgGZSNMqwpTVVVJ6XRFUsFrp
dLervujVrhbAOMc9yByCU/zk5vRglbpHD6G6b3602QDXVnqifEXCIaWCWgA9mmQx
8h6vQRk/g3aYqI4QeJIOEv51g5f9qkVavgrl8FjBC2kUsGQMLDV5oL0x1yQy7+g/
8M7Hz9z1iwAUo1nTCRMQh36P31ikicC1CxqQSQUYGCDWVhGzriIdy6BgGcmOGKHD
SKiDoAaJA5IY6ejQAwL3YhN3fPtrWQ9YXLv7Yf3qBCYxWIXW48KhSt47CNdrOyky
Sb61QHm88t002JdYJEVwcq3ippl43ZV3Oj3GKXqcUHL03GujtjUoN9CAK1IBInJS
mv/vUS3f0d8hIOfULuNBjqDh35ZWP6EcCI5vhorabG9ocjA0B8kWsUQ1LdWP128a
0943U8w51JnxsoR8E0Yg8EgB1KgFWh4cMtPqPHldbbHVhgLT3yXag4RBhJSvcbl1
brYoKiae/iZVjHotdzbzR0xrZ9txBkppLJoguwf6b+cQHRYSp6JxSL039RY7twOC
fp+RC0udfW14uck1M56bz4fG/s0P7hgk0Z32/wx663T1ZMcmmBWRdZuujQsS0N+j
47xcXg7TGxQmWkS90DevT8jO1CEh36ZMD515ignMqAIM1X0up7ZLB3fimk3p4q6a
/l3ZDAEIXlXBPCyLrP6DRcuXdZww2TRO2+tR97oqdjgoFPwSuNlSW/pPIYu5RaCB
/RUB6cKlKYK0hZmuaxOb/EXeFVvkgcZAUfKdkOZ5ssOPK3WYgPr+uMdFzpQXnzW0
0uf6O0sghKQnJTXffBbz5g==
`protect END_PROTECTED
