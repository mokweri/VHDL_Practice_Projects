`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9BVeTk15s4t5343yDHQ78e5AerOnzjMf08Ndpjhdvp3gizleh5CoT5qqp2BySQJm
lss8G8yUOJz2r2HevOik4BDLiL7cyEQrsweo4xKFIcpr16EUXqp7sKKjkkSYqOYE
J0WH7yderH0xTF2xnGr1i/6SHkjbNHZh2MQcQO/i+LkmTgDQFxutnxBnOwk4VvuE
5r0FLd8pdb0pWgKgg1/WFGF+wTZsfY2Zy1qA/cuL5nioUfdGW0JAW1pOnagcDzPE
2mwtOtZ8Kk9jzUY3EgCvPVh24ayqSmk0Dv4QcaDDEVgspe2Jbw7bsi6yD8KRTsYX
Nac+WwMWqYsNjJjivoBpVlKJDqbK2YqTWgauRYVH5ss8WPPi1e92GxaoD2SkIuJu
xgKHwcFHB+rCmwc1djTjm5czxznfSZAtDLqAFshIiGaUfPu575BRgiS7oPUWC/kk
8mzkBqs64xGNpbilWAQF8NOXwGhQqdmZUjgsV0H+4NlpE7+v3KTpRnb5psHxyRDv
WYeofzWub//AJ5Y2d2GrpM8XJdNmy2+tIIB8xR3Gdqz9/Xd3D9dc3ntRpTx6hm3c
BRhy0KjodzJOwY6/KA3ZLpKo8AbqSvBTWVHlamV63xeUctMOxDCniWmG4/9KQFyu
LTFONvIkEI+srnTJCzY1SVNXUl/V1t0a1Xm1b8qzJy+TW2JjKLDODCU+uzg6yK2Z
kdVS7k8dzGY1V318j4fUf7jGmPIe1UbKpP1JuhaqxhYRyS8mz63g3s2KZDRI0mr7
vwxCXPCNk4/wKDueO8qIdu3KvJw8UsiMaX5WnaL0o1/1QTeFkNTsWlGfSUukyZMc
m5GLsRzvq4hPUx9shX9CZh+0LzZAbEeV33IDmOcZowfckElbc6Ozo6DxZkSF94uL
OmsQgtahWhI+fLFrehxZM4xCHPXIjd99N6ncj5VvSvxgnxkq54Ikn4RJ0SQEtr92
Knrh0g64hoM1B7biK2Zfo/pcBy+CuwJIKPa6SERYRBH2LPPssvEFHF5RzuzeDRaS
o4lHdJmYeDQC4fR7h4oIEojN3RpYRwwEkh2+UHTDVNcU2NoPJDJWXtBhLnETxKFJ
d+r/EM5d1Ki+lUnYUXFzt7zXg+SOPHKzgjCBTiluP7k5JxBz/rB/DV/Wjvv7ebfO
DeQZdlN6GY9cPJWNbBM/xA==
`protect END_PROTECTED
