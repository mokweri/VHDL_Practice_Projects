`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cC7cDjgBGFesvVIjkEqqjBL2qn3ikk362j8KUC/nsXmbHsu6mtiXUTr87V/d7/mV
uyRWNeMWGmE9Z6iYUuYBBIGwtDBNbtrcTHpvV9/IZZGwAp7dD1fkBxSbbdNJhobG
YygSpBtp+OUkTpk4sIZ9Nna8GuELUJVXf/xTJL4IJqscLSt7Yq3yPk0ovKRInrNp
5zoFdn9KIa4CWZfLJxxQmPhwZokOLFnkIMdFDtV7ZqDC0mVofcPVa4wve+UU8kKX
vPKextKf0Goy+goDIHxbvdcj98QlA8WMCR6NBjfkOa23/jRm0UgElyFTuNakzMtm
bJBu6VpHzYNzB/v3GroyD51srODvYN8YUEjJoPGdjaj0qpXT09upQZpAeGgkduoJ
5NjQT2Gm2NvrRux3quA/mpXKwDMqqqFgmeEo2KWveiqcEuVPQBFpYFXXT/T9Lyfx
nxVecqdHu1o0DHmGKeWX7g/OhnBKA/MHAZiAtairphgxcpi9iXGhqBgDM16TIzFZ
pHAop9bHaJ4hF77EFba5rvBellTu37tfrStjSya20wc3zbjB0+jjqlch/Ue31EqB
kGI8v9cPJHEBcPQtF2HSqVwOdUESOWvixFkJ/dB1QLFqoF9e5wWALhvUuXwclNQj
98tfMYr5K1cZcIJCm2c1Klx8xjkvRaByEEJSNkWWt52zjsW9WNQFT6QsloVemoS0
FHAsInGUMvwf1PtxDrkQ4+h5H77wVmDUg1uQICzepeLelqxhPUJosfPSSI6vq308
gll4s7mVyNw2uXybMIGx13GPjx/9hGLCjefXxlwpt6hkVlo2gH1sZWeewcMZABZE
4hNTGWbj/zdxH0TNayEGbI0NMkf14Atxac2EvVHpvPD3vuj093DfcJi8P32et9dN
c2WBB5mx2tKWGarxZIaIUQNI7RF2SnRza2ZQgwtiF1WpaQ/o27mBiSK1RJGNSeEu
9yPK5kiGs1cOe234YVwZG3MsJOi/GOzwVKLcGbvQMvsWQV1H1Nt+3wAZ38esZzDQ
k85IluZbbS9H4T58VyExDKXrGcZdBLGqImB/k8zwUoq5Lvw+FN9JA5uGzyQr1jE7
6cUeVp0TR0M2o4vmeXWr0bvBbFxERMwzODRg4SgCr5uC1AZiWm466hqLfPPLr+rV
KjTWne1Zn11QImUfggInHSpjwG52IlACxp20LE5/W+EELh/howG37Z7OkffbRrmB
ntw8Yg4EO4KKmt0MB6NpvILP+T/UFvGBjdpV9cpjQzHwc3Wsngcn0SpwHVT5B0Np
`protect END_PROTECTED
