`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eIkvlCe7zbQiJVeQ7lQ9LuF4m0MDLJYhG4/NVz9WHQ68/IzJfu17qoRpWgURcCmc
7MBf8hIT3RN6iHPZIwCStxoD1Fw57FpsFOjHySHSP/y/WYYDtKMgY1cXChJvBpQh
nGLLP+BFCoowyR8AGtkdOStWZITLGkTvDY247lyyt4g4XWj2F3Qf+Bx9CXn5Jrkg
rhbakfoW/MOJ4buxAc1E7Uti3CxbRzSmQGimW+qN0p7Xk3OImpuTgE3qqqyJ33Md
G5GYrhup48vmOPyW2bcX+g4UyA6cprS6vqr/bavRwMRowv3/lYCjWU2+CsQ3TxAp
1xhsnj4kn2cDwtCzaUN7ookMUtkNhw9zdRhhbYCHcHk=
`protect END_PROTECTED
