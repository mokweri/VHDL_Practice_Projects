`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Po6JoqVQ8EljTXc+iPbAgWpLNk/LUFhg269O2HolN7DPE9HrhLOe3Av+fINgwl4
W2Jo3kI3VIN87Qglo2GSvENTzHwZCEmiCZl0iOkhOgHOPP/6teC/JINDX/OvghjA
E2yTIoBveQ78kuBHAfOVi8cRPUJBwwTaFqmR85SBJJpQHU1RrpUsiVZ34o8QrQri
5Z9M0KknfsRl61g2TPsyNl0hXtLNTi5RLnu9Kc9V9JhZSyXLpQIvmNTgzt+eRg0d
5IZeDnaFD9zsGuBILBahssAAJQiEGBIiGM5PCr2JwV1XuVQjfjTQmiww5ey3ZDPY
82pN4BWrVcdDZB3u0YtgCWf0yJ/U5SjtB6Jod2KRnJSye264dzXTNqmmQhQwa9U2
TG4l2l3jrT4Irra6i/RxH6RREpDIdftqxWxIdVungnskBt+QSS0eetuANEtJypAU
`protect END_PROTECTED
