`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISnPY/Flb9hF1Ns9sCdR+kxdh0+2DhFFJt2EdZ/4H6jKtVCgJWzjOW706yullr1I
1/c2ZALFBorFv+fWKgIt4B4NxwbsUaquxt3bO/ZQsOMyEtlHPsbmysfU3/ZF+Tmj
EKiB1jdMMhY9uvV/+Sgn/fNcD0GSe44ISl8cIeHk9qx/hSWRWm3sdn6pqTu/fMGh
RLBry3DgB8zATI/NMTKPIiXtxtjh+GFKcfiLLvvBhGO3AUoyX49cd6OmpcR4yYBM
hkflOjJzRfX+0T8XU1qJltnm46rkrt7NE+XHYpbCgNTvsVZbXY33x0WmC13ut7xT
HdH+Nr7gXMwWH2SDov7Rj/B+gzozL4uQ/YPQHZiUQLn09O5lTeGtCNuDaWmFJzSC
2DPuWuGkLPsClh6bfBE1otYCZgC28KOrvkSw/pLYc/uBjpPiD5nf/noQJAPHEie1
ywLMNMg0IaKvuQfiUzLjxfMa55IduCaX4fwSaIsrwZuELedbBpajVeKzoLB3N/NX
YleJQ3lPfU3p/T+uay6eMzWHwSjCdKfwEMFEk7KPyElUxQvv3at39V1nULzNBL3l
rEg9SY0OshIDoUx0xYpST8lHj6SLjfuXQmQmB0Af7CYXD5HRho7O//xgMQWaNCYI
t/mGrbfijvJBauVo8eh14PH8EkawLrtoG6RyMmaiaT625Q1WKHdTpMFFIswwk64Y
MjU9LImvVVmSISTwLb9ACpGUwj/wozYidDoeWO7vMcg=
`protect END_PROTECTED
