`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9510dbg5eeMBaY09V8TjtvDDgZDhu1gMrrFSOHqRwY/2dRu7haeLpAWUDIXQp9h
6c8843xyvL3WLdMFrISO3bbXuJZoVY/3mTrB/E/1OPRA+l61/9Ifp6Chl7afNoo1
hNagt4iJXnruDjW2WAtBTNH3FEHcWQUiISZHGq27VWw8eqhSQ7UAh75hm4AtqoYV
JtnaIAPnKWl8DpdoaklTRTLhmYlcDpwMOA0jh/ad+5SklPuZE78w5rkAUqe02lGF
MS4jsv+mu5xpa2Kgq0hUBldEAx95tA6Z4rv+ZZJPmM2eQ38DfS4mb0tyG0w2+lJR
bR2vZ+3n4+MMCZ4jE7irk8+cvCVuIrCkQPy7oJA1yfJzls+5cpWMaP/rtBcFUQqs
5+8E0xv0qbb0w1wft8KMb2HkkhxNbrPI5msa12HbiBGIPJPE62zH1/YJd9Kj3nu0
qxKZfOdfpn7DaURSlHRLRot2RBIefC6XuZj4QwZ3LKK9m/Q7QvGittDMN3t1D1WY
n5jlu7vv8elGJszFTEZ0Xk48wfMaR0DJORvR3rxtmHTIOZNfBU4qRjC0ZNKjXhfn
SRtHY6NgVjCCYdZQ4RB1MovtZTKg3XcAb8dIJFbW9AE5r9Ov6MflUo1e6qifH6+3
FXaDLKvAB9KgCXa4s5TilBi07w2VAqyWpLvdCua79zOyCwpEMy3ZSLPXXV3qgltk
rO/y9BsRIV3EKqfvavSUGwhnBjs/7Zna/Y71o+iQLRozbyh4jhZIuIx6ZJyYQNTh
z5HDG3lhZRXND+UGW68+qpare/ckzkDQfF0Fs2cz/qdyxiFv8dE9q7pWFt8DNc7B
6V8aoi6orvQn67MZdKX1Vf4JxCGW0XqiB1O/7pA+RFVfrK2hhGZ948/KVJH3hEpl
sL+xbmhK966Sa3CSvufk9+u8XetP2Kkic5+TqVhTKju4gLTUKYATK64k1sZbICBc
jkv0pd1FM6iPmNAlDjmze3mJsqU9wwR2YQNdRoRCcNsl4x7M7dW0MuJeeIPSC89P
zUKbGWtGzmhWgbS4LJRURnUgDqsjsUvKFaYXcstqYf+UUIfVy3DpDv/Y7kD7I13W
9yNOBufPy+pkhO6yhabCLFFXAXUEfbD2RCuwDtm/7RHWU3yVTImBauN3Cb8zzL+K
oJCaYKcepPAGyk3aPS8+V7KkrcDTrWcwtbRwS5o6+HLvl4uV3a1DsoLALG3o/7Td
j4Y5YLQbGnxcYfqxlp1oVCC89emENO3AC8R6h0ixLFohIo4Lb48+1Xgz1a6dNU/J
XWIr2iPVKcBDOsEdpvLu7F74l8UC2JrEOc1ap6YoY6fDY9mP81I3J5Yct6Dspb4j
Z96/yFi5iIfEYFf9sokVdB8t1LaO6Ks8QNV+Db7gLerp74bWZ8Zz+uwRA9kK9y/h
8YJT1mqcZPmOq7cs6ArLCPVRxOVDHUQuiWRRGfaT7Xmrptn1sba7kEvTuY/R6PCg
sO0xK8N6o+Nx/MjDl29sTRaTI3Kbq38WITiIXx6pW2EhOcnkGmLT9AgtWDWF7T7k
7DhLBZhhpkJj5+R3pGBid6dbdyiI5Bf4gY3F8U2ZywvHjlcnU/GHMBFjOsLEcCC3
/urSQlY6y4WLN9CJuHhFmun2nACOlxh47TU2dYNJqfC/YQUt/BVcsZeIpynNYbtE
2gZabRfYl5WAw8g+LXY/Sni7UYvUDf0ObKu7MbLfehuXzZs5kN4N2trBjgkwJrTG
hFBdH+tEE3D6cmhMeQSPsrEO5QQ3oG5ePF5SRoQbH08=
`protect END_PROTECTED
