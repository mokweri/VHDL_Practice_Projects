`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
owZg3CWVPFms+QHXrFEUOVGdN0evmFYFrg9fb7NgphBvosqaNGhETxDHjeazebuF
al4GaJe1ghygp80Fmy3tpZV5zvsSIXv53Yy999s2CfFxhi6ob0KwXny6PbdUP2ke
BpHUYvx6I07zORmCS+wMU02m0WOcM6+aIWxHJ2Rgbn0hduIfugPjTi3i9tv9mYfp
zrFtnuxW39I7qN2apVtOkprnf56fLO5/yewqOmFPLMd3aSQ4/RWWlvw5erpP0zZ/
OEfoHZbt2A0+XQ7hqpxfpQ9+IkR1ZcNPLo9DYZ1XoyIV6GPco/EvHqFLcIMRBiIs
kso7Q3GnuA5Q9NO71OnKd91DtP7aEdiefhj2vfKkJ2d/RlNpw8HjwgudZ6nxY2EU
AiQl9eVv4hkzceM/gazw87dgES181ZU8jcaOaBwuDq2yYxGf2sTbFtXf5KO58VUe
nabullzWmDavBoXIOowgwbqvUl7ztRAfJ/10XvvoWpoZFP7NM4pEgX1HXz/FdCke
zxZbQ+j5gji/GKyRstk16ombooaVGIQXA/xscdObxQTbLhA5T4yOOgF3Oo4Rk+/4
cddHWMs8E4rmq2UdBn2EECAGNpZ8cMzWo1BrkzijZaXiVKgZwUvAaTioQ0hiBepd
7bW8t3u1d9uNoLsPtzy99M2y0MwPDSJoZKnjw5/e8nM97UzdxJVIYviYZXXmZmgF
rL5xQ95JbLipntn419JN553GYnU19xoUF19pB8x8xmBgCJb+D1hMKGLtMkFGnl3f
lL/lAtg7t/kAJ8zJVJGLUsiyjlQQ8wvnCwyt6YxuF4P+TWc5t+P84t/Cb6k3hJ7H
ROgAMD0zqcdvzx14nmvm1mWpIiCdXzLaVJ5C7DEWuXtCkWfc+/prlFJK8xyUnOZt
tFqggHKJvbaGipKmT3/0N0+mTnmGpfbCg7xfNGpWe9o36y4/DZMmL30wMs2jCiHw
JOK3k4ep07UlZ++hZHF28fL0j4kmpbhKb9njHVAeab0T7tQfojfLrJ/iF2HcM/qC
viyezmG3hkmpyLIEeREVYItFDCfGxbWzF2PgvIRTaZt4J2f9RI+jaHM6z5iKj4FC
/Ho5AegKfIFCFUY9H/1oKN5Uw9f9h/u+YOa8aPsQZ5AD8IpmmM68GJ7eZzCUhPwI
khIDf2yTbL9E14AFL0Ris5snrsA9ubOpNS9+gPVq+/4U74WJiQdNHCuJH/9snEcE
mB/0KXWP8WOIPbNtNmWH+OUR0lCKCHHa3lXA+R5V8lpkn53D0zK5uaGndIV6bptY
E7z0N7US1hGlwCLqJJX0vdlSVMUklTMXj29iOc/kPoH6S82cV4RMSOB1cYnavdXh
ekaNHpz1/4vJlhuVU7k3qNujlBT1+hM2vTtQjNLWCO5OyKHUIgvofdhTvnU9+Z4E
xDxLwhdN57AdRj/sgF/GQaMrIUH36yNFGiuAQ251nTyjTa5BTe7/EHU+a7h/AW5v
o+2XfAvQsts9VP12NbRrPkQHtYSdxdT/PgFm0784AG+CMjD/OIFxsFbu/4+1Sl7B
acW0+GdMlYU9cWQgbanLRZSvRhvN8puTCg9/l2kM1qj2QVTGK0lwfC9kflJKrkLI
D+G1/dlydyRMGlEnQ5vmjLwfYFcwJI3eKneIld9HHbmPTH0jedHSilyC+q/LkW1D
33u6QSt88sZIBLDAfxtVz/JmMiTDquyWm7TctL6gU0uDfbx/vpAn2vaPmvMuiM11
20droeLyek1x4kU62shbdGmD2eUzU9AV4s/SBToCg24O48JSp1yGY13OG111SpsK
JISZZEOOLuxZ2lzr/KxLFPMzGXe5wfJKCTAT6BkF8omXM3KvyJ6RrpX3jOmxQ1YD
k3iVX+Z++jwNYONL/GJeO7Pes2MdA7W+168C+nseTx1+5arj7JKxc+pnHZrJ78v+
sclgy7Vbr4cNOqmEFUglV/0QCuvWQLxkc5QKAeZUt0BeWYlNJPZje/MtZzxfFA/V
5ZDtnvGgpDdisalsC3NknkHoGoGGGgNFHj4f+KiI64WHaSYI1UFdLYNqJYRiS5oI
nYS95UyjN/hfs/lBb0HrfjMeQa5nKeUhPvOa4fme/JUokt84oulaD8rWl4dC9GTA
+EzMQ3sWvQ4mlVJccprn8lxj/VjD2qv4pRXscNIZVjVS+bUKcQN2MOh4aBMcbzeR
sfUivWRRrKsD2r111T77d9dwRPOiI1FqEthvMiEmMD79UQpgSC37kdwmhlC9ss0X
JncCITv0uQ7RwWJWUhOXykj2seu/Hw8F7fqeKG/VupJjecZU4QgV3tKZL4TclaVe
7QfeC6DrUNHAQSM/IrkHDl+N+9OmGzq/zL3z6qcSLL6iSeyof3SbvxEyaQEAzboH
/ColYy3a1pBIkbKvVGLxfPdLyG/fmUst2vfWyR7DzeNv3iHdivo/vH+rO8XDhMv5
lwf/0SNaYdeCKDmERnpjqa261XEslGpzIT6YWgS5g2h2oRP8DPX+UVoU/seaB7EK
XPHRDpT3yEGR4d5qwMejv7tDQDwjR4xLYxbfv6NKK0FGBbePWbVeg3UeqcZCYKG1
6Eo+sw7fiwYXU5qTyDV1RyxImUbewkj6N1V1+2Tv19R3vJvBXV8H42wH4q5osFcA
vIoqGU7SRrecrQBQ+WohVUg+o4r/vVqEurhrLA3uZSBZa2V3l7YEsMtCacPWWcdR
FhBcqHn8jvHB1hLn5UOwWSAuT5IJMygHeV46bvwXTvs8zN8zzyrN6EukiXVfxcT0
Kr9ArRGE4BF0QRlPG9XvhnJut1hRe8gi7aFrl/4hpOv5llhxeDrDGMCZORUaogwz
fbXkXBzYkIkdEaaSIJnr3LWZ79wMhnUhdQpQ8/vpV/wuAwQuq7J32MQRpJx+2U3S
zOeMWuFzR/cwwtRSN5bfhz3hJvPQ7Lg87L9IO70pZv6xHD16Si27GAZZ+qvArJ+1
qmRAuq0e/l1sRCZ1G732wJOp6GG2pLat3gdZcnX+j41kzWuT3+QriXP4o78tB96e
n8JZUsqXJ7FO+yGPP8MBYoAA6ivwafeo7ygi3bx9Vw+IkCorCQeBhTiBDNA6MkZ1
gwKDQNur7hgaR/FMwkrSESMZwwkItjX3NstLtT9ZTmUwWReP2HqC7NGCp+pBb/1K
3bxHXDfDQrdhJimXj+Laxxn+pzaTsJbtx9aammt0JNFxDW6HkT8HLJIYdbqyloGS
3HmcUQN2TbNFwaULMLgeX8ac48TweGzGZZmGYouthSaoKL8i314JLeqK85+WYuWU
E9vtNFeOzeAM322Ff+VYr2LOERJUI54ZgDVwzVqU0kVrY1bEIuSYyXWyzgbOngIU
9mTu2PbVps3UhQnz4RekKKDdrinB7j0OiwjMchYW2ldc9Jwr9oPtLBmT842IXD/5
x54DyLyOVMBsYYH3uKwn+H6UUqXbPT7P4/i/SBbOM9NJdO1+wrh83LPU+EsgYZ5t
UAjyXxUEVosvD5yZvwQxvBpbezLkc4YwWDhfcdLEkNNQreUspE8ULoZJtOA5M630
MqW56U+SDMfmyy8tmCyTQ+ZtgNLboLh88FKA2AgmIyxYEvpKIPLr1EybutrxT9oL
5Ufu7FFR/v3HqkTBo1uXCRvo8BWD9y7GR6xIyr0hRMBs1kD5MD4W9Yna5Pm5BXF5
GQnPNqLVQyniUO4HrrMYEb79ZkcHrtS1Y3RaVwOgnG1MbKqSFhCTCGt9AyH/L8t2
ckrOBFTNPKO5CXK7UlwQV5nG4zjMOc3WlT3A28UJrtZBrlEpSsoQiuwnEp3DioQ0
PB7yDABV82+weZhALB7PJINkd03xWRbutyUSNdEzLMByl5N3voHiDllRbzQ8kckF
8L2ltRsHMdQ1oTMcNnmPCboRhFtRUuWWoXrGXdIWb+O1s/Xgbjc9OFewpnpEwuWt
ojOE+72f/uQd2rl0ccRRV7Apm9CGtF5MOeuqQTAgvA8LJTeY99odQ++78gHHHntB
GRfqYtzxrC1u1GH/awTqRpgqt9U3aCVuMnqTqIW6Ie5HTIhT6U7hKrQbzJoe0ZTP
As6hXlua/mDadK1qx208xwRI2i4iKj3l8bdzXH5QBvtDg1I/SNOg+AhTERKlkA5Z
Cxr2DJ88mpb/18Ei7X0Vcpg7/FXgiShqZoiG4dtT1tPAfGCEU5uLDJy76SeI7bqb
6FQFxXJrDM1LKAk/8VBuTxyH/Q1hZdakdB4n9N9lI2lFBCAJct48Qbl6k7yNomQi
AQcWcISVOUhwUD2pWr8JOWy2BzS5QiJCQ+P2LLAY4iWS+EWQZKhc+ksCfTYsqZFu
eW/pMk2r/F3S1kirbMm/S4AlpSbUgRZ06mZ82/D/NZdRfAYfZv7IJm6TZLSWVHSA
nPdtz4eoaR7bV124HtwwCuk76xQ5e9B2jD65InaIAvRtOkxzADL4NI/KsGVod7Ig
GmuwmjfV7cxk6+9PCxL0CGCvVAyS91g4HtvI6cVJO51fRbKV9dx0T2o2xdzyP8VG
SJII09NVVBS4U0rpFhgtodELrLV/bAVP9gjjVCkBY3LRkfws3WNioZig3ntLiLM0
d61puW1bWU66X7edikQAwTo5BYWehviS6VFbM16KXEwMUOmMpU5Oa2A15QhN9XoC
X9KX+QHjAstSnY9GJLOYGlFdzVH/kUGxRcqYl0qD5g//fnTrD9SDJ1BCzg89l8Wu
wXT9x5XPKbBnMsC5BobUJokzoyrkYmp+cneWD/95NYFWBsy3xYhtvFMFDjJFdCeW
Kk/Gq8J2/lno9unB+2MuzbN+9DYlzm4lGFR3Ztk1fPfAiVm+IG1UC2mOnXJyZtXZ
g8fb7TqiaHuF2hEWar2I63mxInXl6JJSGHi3zGCYjCMIZcm6fc38izOhaEcU6jom
R9v0ExU1rYWN70Bqf3N2WRYMT8/6ESb4ZF9m1GYaZer26cmdlCC5XxCz1e4hiPUX
+nmeakD7wavw1OOO+/kUkj8i9fD01CFxC58TfEpSCf8MR/OfXEjtnG9d5Pmw/rot
bxqnMDdzo7MDA9MP6lKW12itGw9yGcOXmX43hdAdCuBWdrSzbLr7Aw/pHCgeI5h2
v2QO5Ua84t5lyONrQu/MJOUmAX2VjXypn8KmzcyQqCdGZ9Kbq6bfroVcstblFPip
z9AY3QWqYSd1HvzY0ln3hPtRLcGdI7Znu9q79AuRn/pPA+yMGB/+Stwk00e5T326
3ET5oJ2fIacH+8UW5xSK9aG+EV4DJ/RxReQfmVkHLYKkqtGYkti1LumGWv11jAYv
5zM3bUI7g1yezAxwnY2WItuCZWQffqD+KCTpLapb3EUY+SyqABX7Bvvd3Dc1uqa/
bza/I2oTbovt+ONG8hpl+DyKP37jg8QTklGco4XC7+/n/KMoEqBshaYia4ekkyvL
9nqiteo3CCNa1Ldm0lsiq1cw5nv+ZLmbOn4yi3uXsahIenaPokBaKXMW8ashQpZY
rKm5j3EckSgXaKZoXtl8anokdLGzn2Yl9O5qwxk1VbXca4VqzDZaZNexZxdEWQqS
yKdmn5E+ErZWvieww/P60663eOlAKJIufvtc+NHlCFnhQHfcnKjcE6wjLKfQSMtR
n22okFwQuwbGo5639xaz5BQvolU0dEMhKFzu4JE/P/49NdmYhKjNX+v5StY71ZdR
O5lCU/270sNrXYwulcNeI5A8D853c0HJTCdHrpJvXGG2sh5meqfaU4vF/k7yglqE
aregSNM7UyrjzxG596UWnXDS6+t22g0nrBiO9bxCnXJOcPs4eAwr8POZ+Q1RwPz4
bMiXaM4zcCsnCTq7MpiZwaz6hV2xT/eVLM3ZDhAO0QINShNYLwac4tmm916jjmct
ihrComQxWfbcgLqajJQ2l1CyHQIzrhJrI8JCWw489I47lnVrPDRHsEPhW7MHFxix
MTB6hT/bjVokW1BZfmWzQtw3hFzfi8Veb1rVhnNYFSZ1QpBLWItNuhChiocEy0v4
nMnJgKQJDEPQD+N55ozHD31wzF7l+Z+e2vkFxHbXyvmddmjxGkwyFh3yFCDqcEZr
nFzhnzDpXfdKRcCEfxrH/vTziASZ3DxpbiRnwHpmabpeta/9O/KJOrtKUJq6m2FJ
Vx0BZy0ps8eX5WjaNouJPOymMG61Hf0j3xjpvI9foJvYLVJPK6vEFaF4amFh9BB4
IazMdUHH0o2ej9o3mTAk9tfF7AxQHr/G9ctdloKHQmQyiQaDZFWxbefg+dtA4gLJ
mTDegbVIDM+4yBS4fwWgbhmzhH3Tt63o/bIkXz/7M3oy5AgVFYEKk8zab+Bzshp8
rIdempVJ9Wj2QGmpCxorZ2Szl/HBTTDSmiCFJu779vKD5qx6XspuqYcjIF+z9ozT
ar5dZzWA2HMBvPp93S2iPWGAcjfnFeCLsyJTuvgG8iWHXqeAeQT5/ES2e1xqdj5p
iaoCU8cUHdYBpy4qRdLTIhaxzfi4bF9TIgnvo6qxh9fZW7I+K+fLciT+W4N1rHec
5lGF3u5rpm2O1uSDL2v6hVcSE5cHI7rprcD9PMjfkt4kUfxAydXeEjkbDhl/toJY
6WInhMIp/yjzdFrtJJyyk0tfIP4XptPZg/BQmlFjmHplbFoyDlcazdAK+35GQDl/
0GJ9L0eVVjwDqDV4wwHKI5lviWYUV+7ff21FZJ8hYweAFqPq57+bsQqJ70xInlh0
uPGDy/DFlmET/4YOZwA1LdMdvzYEP8EG+109krivIoqIMr9gBm//TxF/GatzKWM/
1rOEvzF4jaZ66+QI7Ws5aEtdMYmw1l4OUVA/1cmFAe/aGg8uop3saI8kkOSrWFAe
1B28aZo4QtWhHrPM1p+bxNN6jOAKLhNkIAOOMoELLrDAYe/qmtPCyjpSeUhfPwes
lfwasTS8rkUJrTL7ZVxQCJE7NYgM+Z2dZ5v8C4xRORSo0UihfxXc3PJ+/vxvG55a
wt2Lw8pNniGtVSlr7aksYyYmAr4YO48Qo8mGMuxJUEWFhA5/2yQOIzO2+U+LK/J8
WSmLoyp2MhW1cuKrMeegtSNpiFqXGAAKKmIYYjkL7KlwO2drrLVOIPF2J0pwfElm
WcAckCpvHRfY7ktcj89i5Dw27V27NO8NMXN/MpdTql0Ba9Pls7W32bwbr0K5Z48B
np31eD0vad2rCHRvGRMYdVykfeJBzfvQqONK+4ELustSPi+ReGCwkyDfagTnTEt6
RtUz4hRQ1/fpSFjlhAv08oSuosHcUlndE+P4v70rtCXRKC6CKUBbAUqp+SgOrAgI
Iq/bTnechvZoeiLaDS1u3pcQhHlsnZeqNvMu8ekCDyEkOF9JcF4MnX9xnGBHnDlU
QVmmtgv3u6rLDlBU9Sli7rIai9k96vljA9uf1sAYALcyZu6WJJzRb5FST3xXDI/p
UMAz531cdCBEHGB97mSF0si8NLDbofd2EPCdkEhJFh0/w2AEo+WIhctiC544owL/
DTCyGAVUidVaNzAfguaIQi2rhePKE27e/EJqsqqkz0AocQGQFqm1nNe5p6K2Lrcl
UEHs4T8W0Pb9HVNrtxSV4ibc7rzDZzz4TMabm5V/NF6ogRxo+LzRaqCRlUyKcJko
rBlQKCjpFhNEbPX/UmR/jSsqVPB30mDIv7fC1lP3gDVAHUsAiTuoK/bJWtuf1pqC
WrJuSb+RV6Toy0uujAQy5tnX2hiGAlrwwi5wNFzbIEIZdzf7V0C9ogwD4bfJUj3m
ZF75rRrlanHXeAKiwybRbjiVhItBJT3LX1/W4AwuOKVKtc4UarLjKHkTg0YV4J9e
x1Lz9UuxMr3i+y8C5qUuRkooyOuVFpqmZ1Me1Neu+rCjKQ7WLwqJP/FKzqCBOTzG
Kglqe7rJh7opCaff+G2lXCeGkCBQ47t7U58jrW4gvMJnpIfs1LJugNxbyJ3mtKL4
D7nP6dbaQLWG1u0XXDKkbNHd82jwfCGM3ytMxghhiCvBT6vw6F1K4aHl8f/k+PqN
0PdoIr51mnKAGz7Y6HZ7bgM7umypNfh6MAGvP1otWQp47my9+E1pUEOALPRF3YC9
T9JhZ2oofsBK/evlFIHoNH0hEHuywZb7H/e7tmsYFey6vxgpXQ6imYOrQgFC+rDm
s+pkNdb74EIUoeRhX1bNcyRsMiX0VNnZwjHU6sgbMaXNAmCqbBbAb0Z7Ys7b7aZT
hTkHdbFw6zotqGoBX2P762p6rY6BYC3eSRtL33sopcKXBW2xmKKhVTpEPcFfzMes
Do6VIOJ/8cBqCPmjqur5YP5XeCE2Wx3PHjmDzVVTQfCuOZm2Zh5GBde3CH+7ueck
2UZtT6zBepGE7C9D7I91pqJdqrejOnFznnyTHk2hxtYidU2ynats+nLFXJq/9Wjl
PRhhidGFFHYUk/L2dYK0SMmyTTRzi6Q2qLOYzATKdMe95px1TMte9+0K+3GXD4B/
vpYZnqF5ZkLGzNeEAU1D5Nb2w7oQyJxH7qbTAqveLgeS67LFUkJdCN7n2yOIYqD9
5xhI0t4IlfY5qVfSIgaKKfn+Us3oFeTLyKVJPMd1cPSLfJLjl+9jZZnQOHztj2s/
TOhBmVICxjovKo0eV6qUxbiD/Z8brJ18mWdVrVJ1E0FQjLY2zeWXUwcOwOS94WPs
IjhD+3fpGsj7d1+85/eQFAwSR5iJvjHydvN31i6kYOp3iuzAgKc+xe02Q+tFROC5
FF95yjW7WrNabJxw3F3V4w8XEcJk8xTa37r/OQsA4G0qgP8izaBx03E1lpGY4iY+
4PSLdEBKbD1OIf47Spsv5B0BjM4lmA3OeLlOjVh5+l270FfHbSns7wAmnXeT8fSK
c/6w476Idr1hg8Su6GEOte7QyrFQFNUyc5SA12F2oY9c74IxtwRyGqdBZkoiqzmu
ZAcob1WA7FQmE0mdeaa5rsdLDlehj1VrvncFL0EUnku6Yu4FFnr3WSsgOpL3Ct1J
oUZIv0K9rKPUMkj7QXLVhX/ub5yFERme4l6VwRyzUr9/ZtTrxok9kR1FzvDMWoqN
CiDirqQI+nNf3vU2Ya+gify/7xDS6EWkFhqvC2//HqqW/RIF684qD6NeNlxrKrGB
bM7/SBfhEKBcnDAZE9lfJJv5qMBopfD5SwYCVflDkEz6qTkS7hvjKnFwRyYjCMjl
lcRGVwUbVrfCTb2RkAD7RbpYzexbVE9dp+0nivsXms8h5tlEEWqHig6c8R9NrDxK
Dsia68Qy/9dfx+ua6UmTGs1W/kGDtnwFecFfq9HurA4FDuMDXP8DimoWySAEDxfq
wOn2TfI8EN/zwkDYCzjTgK0Lu7xhnWwTyaSUIvBQ5nAPWovQAPZe7ByfJUm1J0iP
ynOK9h9d0DC90nsuIg3JDxKsbet5Nqd9dfYaNXN+/wo6FHHn6sRALDo04w0Opz8g
ceYI9AmMeJ5uFtdShy9YOO9KyfB3KmI/rjFJ4mcMJ8BMsBxnZO4e07FdBRYqdeqy
ZVrT40eo1buRfHCgpLDCv0/UWec7ohBuiojNP8pEG+4p8h1rKHnKNLCJ/hfnWTvN
uSr3lkLmzNUcl/WtJDFImk3QX0WDyqqTolAzrPJd63JOaE/PLb/S0BjzxuCTEF08
QkJiBucY2IMbP0xN+bAIgGQXROprBR2X1EkScsV5npmsNPedYX4GXhzt2xi4el0i
mExbkf1LxfsCmk5V0Kpo2/OmrCm2xLFs8IF9ktCdh52h7JwQNBBZJujBe699nEdU
FipN6t94jWb84KN1RdKz2si/2xb8uXctz/K4XcD1JS6Lt+W2ibrn/a0F12bL6CCW
QyN4BzrKd/45VxO1h28fT6ztvraXUD63SFzB8qyIzJzVCRdofBuT1pr4x0zgGhlx
n4OQcBrbP49CYNqZUtYrZGJ1SE6+P62rosBUXmBABEYcmjza1c/vdyvTzsyz6oxz
wlT1LZCkcXJhD8Zdb8KrCi503oCpeYVwBALaaaYmTtzBnpY8vNHY/TBfB24xErjo
b2koy7fcokpcxy7nD9+9TYKa7QYgWU4pWXhjmr5y8W2sfwJ/KW9BUhXtdZ58t3Sl
BgPNZKX1mKMrTQzYx6Htr8BwIDmnseDvqXxWkd6Fhn1gh/F4vXNpTvdFzmuIbnnQ
y01cvQZEKS+wd4icwAjVe/ysUbhrtgiJnYJJ8CvkooHSDI6myNjrAIIhjXaReMk3
tiTP8CZfY0zCnrkULgHNQaGZ/BBvXhZaTjcoSBNd0DkovbsqT4o1yPukDsPik+RW
qOcC7ZAGZoLzyBZ0gckfLAe0DadYqBCATzBzwp+GUEhgd6JT0LWtwat0sWUJjTA3
eVNkgM4KMge4yyXENtwcMz0SWbz6+NB4l1KQ2FVY9sG6Z8nWYnSHi6MvAy7fjAX5
OaYhWrswDH76AkRmSLmYCSGGjewY17GA5vsd3k9MjRmXXRp1TRvRyi3/V8pHDylS
sZ1l1ug5uRSAqU3Dj9Nihfn+giEdugxdcV1MmRMddCOVXsXPBtaBEfex29vZ9Sb7
pD0bk3mhPo0neqqgGApA6dSfeM49dU8/J62nkw6nTPX45pCYhFwBXftoAhsfGqrh
IN9BbyO30p1jkTGl7HaLyz7jpKjD2SqjbUh/uuFb51rGhuCBk0dHjC5Oiu1q+qgh
TqihUHKSLX5e8Hcpfa4YAtDtJ1/1OqgHEjzDAkbcT6ygYGDh8V3BneETadvQNzWb
o+SxFNwctCpJ4/THF6Y1HXpvS9XDo8TDPKwFF4SC3wkmMQ1fW5LopCSiQVIr/eys
K4BKr9FLUY7QMKvJ3y6Fng/l4ExR9TUQcedqREN2+kbV9D6F6Ni1D5IlhXSAaR6O
PLZC+8gFPdAlQ9GYiQ+GNLmLbzb3BYqhOu7SIUGAY7ceaALPX2+dCkdtEuFxGL4M
Ps35BigO29DgX5M8/qkNPAvsMxjFR5zvbtOyE+3O+yMgRDhml2PQOCty5NlJivBk
LV7an0wu2pY4j2p24sAafrfTlg59GqT6bxDAtGNqnmKZY6zpsIk7wvU7K9JA7BBt
iaqLejV/853MBeYJpKB370OrDtu8Itj+J3F1B3I8DhkXGQH8NL1eBKlkGGitjdE8
ZRDwo67XLAVxJtOd3Dd1MXmMlLlAsBKk6VMGF+3KWRDwvAnl+1j3JLFK5Y0Qdp/T
MLVtrHNNjXeYfsHCnMHDvpowCv+z1xsRI67KyHQeDcB4908K0hZNYC5GUKWTDmHP
u8anv9t8vJWn6cVWITkNbAr4CGfzrQ933gmgqqKLluV1inpiie4EhJ9/gCBFo17A
UFEiICiYGAdzfJzrBjsY3x1+LJf+me9ZcO0x+jQhBiU9uqg44zawHypA6DYBI6L1
k6ErKSVDzVaIttF4TP7FBKOrSwMNRXmd/ToHr9nyTucuUZ60Hw/2AjfH7KFzJcJ0
SaG1TP/f4ssYRIW5hA4QifQi8XjNV7CfbKPgpHr+yw4FS0II1z8J34Cf/vUjDNFi
ULpby3x083PBzk/pBUwayDB0GuHA7vZtmY9MUaK+N7qNs6yZ0fC0rRMOEo10YNF6
dB1nHbCaIWhNuyMlwgduPpqwWlp0f5G+yG6jqf7ioOubXxMy/S4ER6CRbffrqckC
LDqcuSa7zLc50dyIwdOv1nqyG5bWsppnpmahrEksH/NwOlj1tTcUiE+kHsHrqfAA
KtiBCsNPH/6zvG0rTH4a3JD46JLInKxxLoxhvXfeysYVw8aLD++3p11xUt2AC+vr
o5QxJRXlwTPXsShyOkl3nyo5nkvVLvkLWl0w9W1S5ev++iBM/9pJsvG124T/NaDn
7VbGHLATngEfIpu/C+L6pnjVvxjXcodGHaidAclJj0ADraW71/2nduzcoQQb6FDD
1UkwGC+80Q+H1H4QChr3l2M40oomikz3yMgJlXZfqT4aLnL/cFEJmH5HJkOCKpAG
6IVYQiaBIkCB0qaMbu/zPho1BCmrm99wGGIGF9ChqOMFM79t3KvIUT69/GmIw+ff
KgLLWGP6G7rpNR7vqCFBrUCPWSUGI9zSxzdNHwxGYIjMILuvFvhi7x6Clyx7PS9Q
FdSrAI0aSpJ4YE5PX3oNN5EgyH8ckdbhE5KCLhJ6BaNwgOs5VmOYtB9XbNvwdXlo
2nid4PZQ5mCURufkA3b7CJuJiqfkwbwGnMtTVjQa5rXlntaW1Jwv0tET+GkOzEU+
itv6749YVvgJinKsJErkqQ/glrlCZ+BgTNUNAv/IuatR1cHPs37Q4WyT9RsILXiN
UL7AW1gaN+OnFXu/xS4JN7kyZk+KdXwGggZxFgkRlCk1L7xrewlghMcpybgrQOMc
NPXgZSpqd7crsVLzlTga7mcyS1t0kCWG2Rnqagq+0J6nSIL+Ig8pjdEcTmUADNsd
3+EIutbJSgVM/p2aXQl47p9xIFcTxa8Oyy/XQipszzdQ7vctEusWZwCBPJhIhxG0
3edscN7TbQ855ZYxHuLw6nLS1it9YyPPiSkNqZrCwMPfUiNEKNzzFN3iANNHqKjc
0l6J1ZMHFssbjmmxGsDFo+noFSahK8pMDEAZVg4pMKs92ua7+GD/vtQxFDiOjmUo
RvdowvINWk7ymA6zrrIvnWIDu5DFNGTUa2L/w8qqz/4M1cH4iZ3RB4zWz+D3KF9D
OViQME/7Wjl+ZjHBXcNxeQkMv4wrbK2NPtJN2kxclIBdRL6H2ndTA3F8hQpMDajU
4iLWAkAAR9Lybo/5aW5GYDrEMSV0kOlZQxEA0ttnd3mCb7Iq0eGPt7IF+Bs8jJwR
IVO9ai7BjNeQ7iLtSHiLYRTiWtlI2dPwC4c9PXuSoQs6sV+Gc0W9MyVBB+g/SsOJ
p5x69UTEwYpeoo8lXtbVZyL3wDE6WJ1TlQ7p0/ZjzzC1hqsiH4SU5//bRCShHcA5
u3cgN9EMOW+gAqVOS6LccZyA0HML+Fv7Taipg7VwDkAtLL9qTafEXUvxzosoeNDh
bn1qBD5spdcowNbtXpyrlcQ63ZQfPLKLadL35nAN4b15IySpP7zUcUozGeAuJ2nN
+EsMGDCZbGGEkqxIjvqqkJPmA+0Ju0DOgBCTPYecCVcb9m/XJKepIOVdMVZ8xFTE
tnKdC8i0RLIFijp5I1tUJ1OQZLAa/cfM/6iqRIsyf7Ac6UUNUtfQEiqppFa6ipLM
3OA3TDdR21qUT6MXZ4McOERRGdhVfazSTS9cc4vCDl80M5IzTCZRHIafinhdp6NU
luXjJctXRQeGn7VAzvY8oI2/9cJGtM5ZCam1wG2HZhfakxNr+6DjC6DXSf1Mcui/
6HKv7CkS7WLlnkfMgVGNhWI7ypxsQihQBQOeTfAe7+4bhP4wcElldiYdcAcm+ff3
tviRi3+KrMwqPTmGqxQ9TJkglU25jnIRKt5ljXBqye8TAOf93GtlBbitc+p5XOUa
mA8suxquH1iGmgeHuHsI2joO3FfR9V7hfwLvcbigUMCxiU3vQeYFCl5lICBrAuCF
fRHknYKRKUL8pPwQeVM6fznJ4u+coG8EhYigOz9J4OElzspUp950tOjWjVODlJCE
rF7dI4hIf96x6j3gjRrUTa4Axfi+gp0EplbrRDw0PYTPi927zItZejXyCtetCtc7
LrghA5UyIxEncCJNAY/RwYL5vfeLmC9H0xV4tUYZ18BiISIwIS12Ns/A0MPUZSPx
o3PSEAYdUvHbIwhqO5Lxso8z0vYHR+FJT+L+13eDq0jUNHYWS70klJX+BYZzj55M
vhLUlFXiQzQexq501K/46q6H/NAQmsIC9loyewNL1zKdsKNWIimJ4jV7K9dQ/JsV
i835x2/A71dtcZ5sX3LUJpYkffC9eTfi6qPR9W8Hos6ER656fsjZiiu4zfEyQ9v3
JW3ys8m+Q/qSbvtEzMtbOpctdjVcPJRKfSjBSP6pDCZddVL7soT4ck5+iaX4qSkV
vgRcNB+CWVroLVa9Mcw665OwlNnGQiugZ6NFDdahH7KfbseV2FEp8cRu+YAQDJk8
ojUT1LwB5f3NLOLTZdCSchbgwsBisvMbjeULZ2fBmX6INGTEZrbS0LSAeP7YwxKp
E6cLeYbRMg/Ud6RUyl2KaswNVAe4dlYoxnhOmlF9R4GeIwOC/sq1HwJPrSoi7pDN
3I1kPUU9yWk+gIdWDSuDLNfyWqQLP6aanH7zmk9GV8kT2xzn1VdYFhOo6eZIkxKO
KAcvmGEOitjm28vOmVOmQRhWDyUE/P0YGIodNreQLqhVY2llP1KPY5pBiI0ZXFM9
w+SaqXi2zrfvYeZGzekJdk6wRLiiAsZe1fztduIguWHBHzjEWGScjojuHtn9ZbQX
8Y+yWC4gb0zy7CqrQ/FIkQtw8736GPuoZFcd4yroX/PBFtsNryAdGPAH1qTGoHhD
mOAkX4qtzS+08IBDq/E/NPsYDogrBMTOunIw8qhEFqcY1QikZLubOdTM92jtq+xd
7k3t7+hiOB8PlqoGjH1a3BkcAySOEt/Mpsdz3jasbJ9taeYBBiwRMRdPn0OM1w7L
9qtUDhB/K8Ed4lzCcHH+HtUBYlQhG3TdR8FBWiKjVbXzIaasoFS6LaTUSvNrtewH
SATPz7i302uPLMnt1MbB8cyTyTuHE0tWUdSWGRICgbX8XOdX88eUktShpsXm4nKE
CMapfkqssMgC2ooptHwHV8glDbLYhkSorqLX9jrowBCB6fEghMtXs0qAN1eB6dL+
dymuRcHCNOrxzSTWC5Zkkqn/bRzvrA/s1epmqfP9hHpLTICHufrXS+MSE7+QIolZ
OhOtpAmHAWUd4aAxM36my1RZDhvHlncFdSk/DlIwszpu4UpzCbarVUFBpi4Pn+Sa
azdD6pBYihFreZFWfJH/TE3adJuDg41PMyRd+G+EEdYgxV9MQXqADSM5KhRwe9ye
v4RUdHA+o3GMqZUACthfqc/u3gqdOfNPO/l1VsZ6vGKKE7nN+QF5QWIyDzBPmF9p
yxXbT5kTFsEmHJSs3DYl7Btcm4r6l5vWpcwgaMh6g9Jh6w10mAVQ84RiQqR+MwF0
O0oHtuXIAd/VoQo8RwKVIZ9aBP0lf8qlJldKDitBQXRMF9NtD/YUJisR3DB7PTPD
frVJKjjqSF/nfVCRVsRP6KjnFB0jSFVt9k6UVUIYYD64RrydoYsN4eLcJYYrNrcw
/VqW+JgPRCUTRgG2E1HZcM7lcaE/CmLR73hDpWaaRvIjXSuXK0If3zqPMYrTsOYy
Cw4leGixqu1Q+9zh0ZpPws0E9wlsTQu5/OOUQH5WZO9Fvza+IRuh9YlBugb+MKrb
7Kp9sXYtMsqKESAJpD5/FT/ptfhF3dAscsQMLY75+3xgeR5F4uk3xnRLqRkKHaPr
2PxNNeFzqkKcFApQF5Z3tF5ixEXXajEr3XRng6rfgOg4AyN4gjYIphl52KRVwhSs
fPA2dt9smDGTs1Nb9YgtH9WHWbt03nklYMSdUk0AJxjBnsecfx1dOcCY5nF7/8wM
KSgUw7Q2czcGpwq9mRjnxyxmGVaVIWIxxCi8Ev+yBOVdEpQnJPvyr/JrNsO94aDX
80Ce45a/NSdKOxjr43Wji0JcWQTpCD0JXqi47r69YnE=
`protect END_PROTECTED
