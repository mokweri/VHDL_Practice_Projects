`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Cfl2Z9GRYEi8ryOXANyFSE1nR9qUtgEyo0WvUlu9ElT0RUqEijOgTf2ac+iSDpc
pKHRK9Igrhux9W8BHpgXncmDJcyWLueErMC/5UFB5o612EOc3e/po+VY4wt1Xhfd
zSuos/th9tPxiCPDH7nWNpXDxMusq2fax/y4f6BzvWUZffVwVAnLj9+azJEEAQQG
y4NyAW8i95jVY0gSeI5maBwfk4n2Mp7acA3ho/uG3/ykoCih9GvQYXaPbo59wKan
XW3PDMFRcD0iCZl072kc+FTylTCK1xR61Xjhf1dOeVheP6v+EkChywU94fMolLl+
Qk097gwX83ZudwDLTdymrvFFO3wIdA853Vozh41wUGKA/O8Sd/2Vvag/h/9I6GDJ
kveF4s/8k7R44AeZq1oD56foEqv1SqZgSyzk3uRn5k1j6oPbuPg/F89BiJD9yxaG
aG6aP62JRWOlWFaCGYiO6VG6wiCXMjbCiq/jPRTO/mvsTsm5qo9ryprZAFstQHV7
Yj96ZrjpYRHSdFPzvJj7ESyHpCajITbqZuvLSfM4eFpcOKTOXJfGBbG6y5i4NMNT
daPiMHxtDafuuoubpMl7G3OdR23UbOX4ZPSBjkFldiC+6zCACZzK5k4d0l3AzBmc
hBm/+C5DQHLUS1gt4Lu+O/zIyBJ3tRjMhT8Qt861+INf6+IMdWv3hduJYtE+dXlE
BJQQVOwl4lMBsSy/Pc1iUr3/z/v15V/63DJHl1j9Rb95RJ6OH1pbCDKwkRGljxjJ
gi3+2ZGf8cxbYtuVuaK7uOKkA6jcLQ14Ktkaqinp4KOxWyYRbEjHUSLSc3i6iz5q
hfVLoe2vCJ/jHG4VgAePwbBVbS2ycqCR60tYfASNTmSFXnYw1HT0DKg5q6Eyp+PR
ckvBxp3Qy03OoQIahD7dIYbWkxbX2deef+rSswz5lAXtVe+8217DYtRgPulUIgWe
/tVqTptu+J9jdCMqfHn+D8JmqVH1vPndpU0fJtCNJ/xrz+ew3ORDTAYSSi8+SFym
xExEbCyHWLHNMf8s0IPD1T49KridSaHD3PVIAydWXUTaLaMOQOQXCi2u0fLQY3J8
r56+MJN4RmNCpxeJCaJdKFzsWT9mRRgq4AFxDHZHwvfjB/Kj7hY0dkSS8+Be13W9
e00gUOFWOzh2398a8m9I2kEQ9SN0kfk87WY5hZBWAFIocyz6Vqv0jUN3xgJEB4QU
WdiWa17xoepiAXGBiVtsrX246imifirO6n2BsopFer3ISkapF8nB6SxjpHB8uATp
RZcurvagWpaS3YT5saIBS7b7xTtD6l2dOOdkmECFGy/Rc4FtWLrMkyDkn8k4wtCp
lDzX7OUaXEx+SnQKUu3cuzFY7JTG0uP2BB94X9RtxpZEggW1jgNHEsl8aym+Bkx6
hpOjqQjWKoTWKMJzlTZg+0j+3Q/it2z0hdN0o78F8M1bF53cbwdYjnh8bDpNSJHy
WCb/4JkieMRD5AW21edOc/mxSuQboAqDqXM6MMQahbJISrmtbmMc/mBhYoO58BF4
muK9hvJt7vu/hvAHPmtRk+JM522MUpXnaIXShP5aZlqgj3ZWZxXE/pN61UyEbIAd
MWyuYIFDc3DTuB5Ccy8xOYbAYIQKYLZzbd9+zu6acBw4ai8ApXVfqmpU7CBL9GtL
mRvjJ+kBOVLcdz8oBWSTigc89oirymViRgrR3rgKyY05ac/T4Tu0x1EQ0dpIPRt4
Y4mB8cC9oTKfLKDypnABQj+5tyHRKl+pp0Jjy+FJkD5RZpHtlPKHjYp8P4sh+gWJ
no/nwYgNqymMhQs+zrKdcEyPb85AwKz8j43ERKQCdlUg4jDopowoAZfLEd/2nwqX
NEat2Pke+HZvrqM6aNJSaw==
`protect END_PROTECTED
