`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycSPtqtv+7goZtPrdG0UTfi7f2h/JqyRkNHM4qD/1QV4d+uqJg7q6eaiBTOsISwa
ZedX2MQ+xPYwd4yg7jTEDm2SEUp+hX7Iv4Q1g7k+R1c806cWVCGT+Y+LafNVqhCu
6qH9wyujMNpsu0Y35bwNHmx/jJ3k0nMe33ZM95HQmtzT3hxX0mVnQ/rJSrn+t6tS
3PSlHg1NLaPAtbnNu43ey1pPLltjZjk+cpMq+okEk5K2gHkJVOJ0VB5H6qWb1otq
eKiYDHFvjOGWXVe5+voUXnFWVHv4EqJCB7+bO+pUHtsZAafkryWSIxMfRtZOQ3TI
IdJ0zpurrRbshThtc6GaDrvESzdaVK1uBhxwjac3plegAOr3PtZtA4kxh0AkcHZ0
+9Bjm95lEQ2CVj+tC/7zDzw1KxwjY2TVaX4+g2wMKRD9np+/gYn807UXnD8d98Y/
SbrUE1R+gI151+ee+HtiU9pWRFktyDKhsXOogEfgqQ3AmrKPmC4qDOK+gF77Ic4F
Nd7lm420MMSizGbnpepM/iAP7Fv4Iv4Q+Tfic8YAsk43C4jq/1+cl4q822fUFIQ9
q9ge3lVi5qb/D63WXcS7sQj9XzhJ6AAuNdtPdRHla/9yDsv3fP9FgBeSepfzzGU3
CgVWzkWupTnRppUvENjNp4S/b0hLQaqYCw/2ChS0MRjING0slNg3dsFIGoz19LRH
KA/SsIqLxFBwtPUtw5CNjDNdXXuDB4Sz0Ik/u6m/mHTyC70Q+K+UcDWyvm+Yv1A9
Vm1JJiLLlAtXY0EdaV1yILzJgwwdtFyvQK1FEZ3KC/znzxD8VxnCdE7tLi66VuPj
MIInsZPcrV1/xkrfwcqN7k2qcNG6gtdJ5iqdiW4mNMTe0EQD6wThMOb+JJ8DGg2H
KIOVDLCF5Lg0VUjbIWdfoTEDodE3OCb4nVLC1IEpo1nnSriUJCixBqyImK76ktYh
GA0Xj78iZxOMvJNNDvfEn0nKJYdr/MGbLNDvrWaL6I9jN9VR8jIIfGIn1iBYj5kg
/t+ETO7IdpK+t8HQuzFim7f1Yk/ks4jfhw3XaKWxf2ZPvMHe7nNgpCIUSeI76PvU
GdocPlIbkiv1NJNKlQ2bGesMo7Jp7/atoAdU6NktyLEGCg6o4+qEQj62sNDCSFGR
Z0cpAfTEKAcPNUxECn15rcKIOYQKuHWILwCYMgPYsG5VaXNZo2sWgohy7+6JcUY5
fBtJB/Ynb3OXn0+HBC8+5WHdt+KwPFhwFu4FCsGXyF0rKC+VtyQPQUf3dnZjBUHr
d1zAA6IHRq6XNQTAtglIwUykrYt+FlQ62nj7VX4RoqNQhrRWi0ADkhh3jACqR3b8
ZztoqDXDcojLYzXbKJhpR82SGfvq8VnEvMk9UY7vHxi4a/uxtp+wYYLML/okf8Ic
ZLRqzMzTEz//DSWsSZzeUHI2UkT8mQLQ+ajlzVN1TuiYP/3lHv9mQ6ME9/JyE6oL
njSKfTlxE0io6ywD9rfeKjPswI+ouIsSndiymaV+h3tCy3fM5yUPn+MZXd0qBmk4
skgqNvJFOWCyl8oW+Atq7jwGW4Z/4BJWBW4FLiW18kAgR1beppUF7bG7Fo3fkH+M
H2uKRTAhNAN7+jqQmDQ+r6lJdONFY2t711UdikmlRhNe7qXWLH7/H/YJ08IcO+yg
baU2KPKiKUsNAwCeyAkHOn9FWPF/72TS147d+LEN/utmwpBBraPBm7T/JoIdDt18
PjzPJyr//iENr2ik7j7fk28Uax7UERGwxYwiDhZNXZehrfYM1evJOhu42nZIQNWV
c/xnt4Q9djgAfA4kD2q/8WbeunvrNT9RTC8APYBKEDpqFPKEm1WsFzKANhnw6Xg4
KnnEra8AXpzfX+asaEzTsoRswnhko7ZapPUoTzxQWIdQpcc6h5GtwzfgEGpnRviR
H0uBvZYGTAF79/NL4czd/kSjBAMJ1bGkFVg12aruNguDzmpO1VV2tRpcflMJtwfJ
4h1000UwrDh1RCSWfgomQkkxp/nRZMRylRiQYS2wj3XdWxBn1ZSaUJBlvYG/uGUy
3xtf9Arg05ExGxYC+HMMi3Pj3rwImC5LoNk01k99z1DWlHHUt+c4VC1xG4GliWF0
/N30wf3MZG8/oxpNmRPXjvWBXpCsL5ZtMvtKvSPfoylHikLNlrgMSInfwVgvwnhp
cq7yU4D4dX7I2qgDCOQllPHI5Cp3nuGsipCgJXhD0kqF2iR/zQwUa1SKGVPlQlAe
3CnY4wWOSlVDWWED6Jny8KWBmaDGlXaZXTDLzQlFt9GVxoKZToAycsKm8nAFoRP0
82HAMK6lgeJCFda1qIj++ZRJz1NN0+K5b6Suach5PBBDRzZ+2hIfWxQglPifPoKp
y+en68NITnk70WQ5kXofV7oBACVKv6QTPMXxPrfgO5fiuBVcIDxctKowMi3eGYJK
BNxiHd4nnrONWFjZ7Q5FCTw6WJ2P6oMDRWOcpD0vVVQMtLutu0lBZL8KQ/zX9s1N
xaEMDJXxP0tQLDmikCQFCT0HtmKX6ILm5UD21fHiIfP7nmpFmyfQTQrAvLQxgHcR
Tep/a7ZceX3h2iedptGVT4a5tVPJKaQhpDV98P0DO/drYf4ZOIedeCPnZ8Gjr1Pk
DCnJAtZuOISgMT4dI4hPc5i6gWrDI6KSuEHLP5e2nLBm8y6g+oyalwoMRLTUMUiO
akcLWPbMoqg1EquuQyVc7HGoubyUHpP2xD6/z+oBkNjBu8heau14ezFPZptyCGFu
0lfv/4RvjcaLvfh3D+ms2gmS1QvO5WY2WnorWvBWZLhLov6BOPIk6B9VLASXOaEc
+kTSGVfS3D4PSmfgbx2yhO8wtfQus1aPLqVQ1cedeuXWnFTqAM3lMLiwzX/hwZ/+
QjluM1c+MSejcdV9hmdQ5ndHjiRqmakzk3K+yscwZREMo6wFLe1oO6N1h0dhdPmg
nLOTlh8Kt4uhZbEJBQCzCDCd0h+j3rAOcfGTAbjCNycz921NM5eDpB1H2CVbbay1
MEHCK8wT4/GgkduuFDEt4uKTSAKZ8BimQOKAht6Qt+Yopfk7Ph3N+hZ5Wp6yfJjD
WIsnBvMnkcQc15uuLNRvq7ef0fjvueLSdZC5rIzDkqQYdGIY5BmbA40Us4SMpvMb
VNrrkfqzqFV1HolS/u+VhdO+VyhFAs79Uy3J4NXYEgleosxqETKilMZ96UFU9C2h
aAJn2dRCpbhc4bdo9+FrK8c4Oxe9jlf6gftdWC+a1wwTeNfA85uKeBN3lrCNLcqt
+l6f528PEf1YKiig7LVfcrZotu4j/l3f1Kd6V1rNIQV1Rlj1jvmffOg8uW4TjROe
3SmPRMMTH/QutfOyZ1eoFHRil77h6ChoSZluWa6aCWzeRcT4XeK5h8LumbwNxBdj
3Nz3oW0PzL9/2dM2q6DbyUoKyMmb7ExznqeTPTiHDlDmEvmguRUwALUKOYoV3MUH
p7wavgtOiiEEQu/VQD4e/SPvf985h64G3/DhF1qNw9x0gnWL3WsD2eyM4mISxqQ/
LygY6G46CQbnIoBe+z6IS4fFvdaPp+YUyvtf7w9lBAgERrdCUeuqfEJGyAMToV3N
uvdFX7Rrltet10U/HXJBd1s6fwt0q2OnRVRRWMdT2taU7SWpaBT5v5fM13xr8oVK
KqFFjfLLVmaJ0ieqYy3Dpfn4o3JEJdjLWcyOQFMa59zdle4tbYJ7fOP7+Omfz4ol
8h7cBxC/J8fwhgiZAxEaxb6VNhbIUVWbPp7XlVK1aLVNUi922nU7s4JNRH0CD7sv
5xaXtS3mL77Wv5sDmg3qyFAgT1LLo4RKc1wE4SHSBM5iBPvZ7ohUxAtZjg5UB0HU
XH490x4CAvLQYX6U5QrbSXTiSlQnBq9q87OUbPORTIjLs8j59jT2jNhmt7SBRMBj
VdYZJOixLIeoPHc7OHAh4xmeRu1p6yxYaXQlQDjtPv/ILQJqWzhZMEkIlp+ja/gk
TBtsbnWzunf6DYLY1U7QTLNfoQPQcsfHF9ivgY8TvqF49akEupkWnOeMqugfT9nz
ZiBdW+q88emZMnHF+0keF4kfhTRXGQ6VKxyWYZ8hr96tdG5Y6SxgkH99usjuE1S+
wWHMifm2Vjez68f7m16mJozs1H6EqbTVdcumDGEk4yQPk5sY0rmc3H/2R7OAZeX8
N/VYgOpgrpFshFm1LIdJoORizBp2sijvWgvOTJ4aRuLLabMIU9xuiwPbdxd5otUo
c+uYJLBnmxAALROWL5yCPnD4IdkMiab0UaYRBgcgYpVOKVu3NW3E8a+2rDSHe1Ad
`protect END_PROTECTED
