`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqLt3Tp9788jyVjNsz9siQVZlVbLzXaKmzMTRlTYTU9tb+nOUXdrDU78OvttoP/S
35sjt1TA6bT2ttY3qHmbqln6LsxdGqoyvNC6sMAtztSV2+/CYSOBOmDbcxN0w5Bh
Zm3asLBMiCG1wTCjSbWoISpUWxrQzCJds0AF5WjhvZYaAYfRZSPa0PJI53dOHpuh
dzC1cSEg00wWX0K5p90vJqqzRyoyCv+PMie2dpJHE9/IEgMN3K8nwidqOXZqTiN2
pjLAcTpRkZDfyuZLLOuXHQIJhVptZAylA/dDaCUKBINERpHjelWYsHNtq1M+kkOt
u2J9DTzEpTsEkM7rWnAz6aeFIhUTxnn1IxMRIZAZ8ZHUoREO5YeWdu7BCgI1M9Kz
JfUdNgchMZ3Bzo5Srar/25B/GcdGDntxOH+dcXf7rhruAOrijgu4wtI8RS6CG9+2
ZaLgblA3X+4KVHByDVd4GOfTzR2teYaufgFJVfAws1lXVihJhAD49k6KANEHQkJf
UCcBC6u5k5FFFUKwP8jAKskr2vHs5j/4YtQI/YeBvaFb2QXHqNz1mG2b6tHj7UB9
fKFO+NJDqSw5cWea8ad7pr0WoM6SqhD86NT/JhbHGecUVGPFSAI1iWMvoqOV4q3d
tEUP2kMNFP9jmLCFWRYv2XuFo5AuG5kIaqnbODvUIcpjHVk1ZDUWapa+b2mYpJch
REtWHEIDwpN4WnDNbGLUkry41AcVYOK/LLydcP2CMKAwlLi0gnq+RxWqR/6fF+jJ
qLTLVkG76f7BSwacWjNs9pXBXhpVUwIn9Hjo5nEkKKiHxmd4ptw5bmRQ+7VOE1OA
8qPG10MLOToAkqw+bLNGnzJBZ3uqTl+j7ZOg9JamKZlffRRbS+qsB1lJ/3mEbTuq
S+stJhAe0d81nYfoVzRkZAgzrUIdPhwYWjg9htsyg1eT41OJ0PkDgL7Bg+0bDrlB
5HdUR8iEjhMiIti6TG3Hq4gBD3tdUMTOx+vmaEMTPD3qHYwg0GEIB4u0om27gwk1
QC6n1Y1MUEQsdCR3ADnyCafMD/56fZqLy1FH/d58UdPcRVA3qR1rthpwMIM+EIbH
s9S7NT5tA1INoO0TKiAZARw9B8+rbg0g8yVQERU2q5OWEeC7z4aq1Ncakk8RmXTj
M4wLI382iC1U1jXSng4u4ayZ2/MiolL15rnN+TsUEWE9IgDOhS0kh9i8uVnxwDYl
mrKqwxNBsdu+BbuBntvVS1pFXsrBYBG2CEyJB4q3uwS768+JooH0CfNpfRJEHkSw
KSZQDi7kbdT/xlQ/QCeOo6kio9FcPRh57Aaxsp9W4brVjHMPhWQJjxfaVqc1xOAP
gu0LkuNXCq5ByodY1Y8sf0UBDB8xgOaV8mDGfmgDMXR85X0yAEPIhrNNckMbS7TH
B3kougXGQDETtUPLCJyr0U0jfhkRwB5v5a7aTQTxSkgNLW1240D04Eb63Wb/KWd+
NsHfJTzj6PJ6wFkrs2AKFp21E1Rka3CvTJZ1hKxgiomUWdZhnFiIqpZ1KNUcLJfI
tkqXzCTBkXTVki+syfBuv/zeFfOkjwZEXn1Y6194MZohw/JIOPE1K9rrVCGlWr8D
Qm0p5vGF8VvpjMu9mRosOLLRJ3s129UOSKihWl4xVs9f7JS6iRTKUCQUA45z96Z/
qdhvD+e9FE6d4MIujxKuAUtJ+lE7WJQy+G27djIImxGTxcLyhUD79JlKbRYemVeQ
h/ZQo7I+21m1O1z/i9eBn870DilxD2x5cdFqQqJC4fxmDZG1tTRZpuXALpXJzPt/
lGVHsnWQ07eXQK3MNB/kQkRsM+XbJL7Ugmj20O/XIyLutj6DfWEWkw9eWF1bC3pA
ilwV+1opIhvaZOuot92d/gME861gxbK+GgY5EsscxWa4pBxGWA6mMUuxFZd48Uh2
gCo991JXd3gbG8ClPmMnB9rqtljgknMcV7mjpGnIKpE8pkDOwBfrGyUxr6WDeMuM
7tNkzrvq3hSXB4sIYCtT2npjDm/9Pf4lnianCVFZlOYBMUWjosNdAb3s8629FSeP
T4SpfH6odny+6EEgJsikYEnSmVBKYjDmoohoqWESEtmi2SMyZMHhEsVT6tprM9NA
rCPa0At3SywmAS9cR4Cz7GNUf2RTJCQz8vqbNB3Z5t4PbtQCuL+mkGRBbd2KGWJr
nqAMRpkFQiuT+/qVAx6LJoLoV5aJOhqdqcSdyNgccNsq1AVyMnrd5eW8Z6oi1DPn
7fvAfNkCYejKVmX25qj/u+DjvjEdiy/aW25/GsT6cGsAIPG9Bbq0G2AoUsNGHyOv
wfNPfYaTRmhPNdRP1Rn5IfDKJ5OMM9P1y9L5miLJimmYkulfQkpDcCbI5jFQHiDD
8XLRGEzO5gjVURiONR8vxjczjq01LgsxxYaWNRD9YRX3YHpCMVIHT4ZmSWNCoMWY
0oQJNAEMhkq3+Hi+WGzoww==
`protect END_PROTECTED
