`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DferJsYPS6EbWAbV81XCb57k6qw2+sDpOkj7A6E9giBeEHAxasUaNg1Q8bVDJtSI
8qbzD1oxhJVcNoJix8bMSPxTfjCf2OnlIean89TSAhF3lp+CKVLop3yaruZ3WnNc
KC8SCV7pfB/w0M5KzGzaDkKLoOgAyUfT/MWdfqmmBVbHvTQpYAsGPi+fSXQGKvXw
IRWFAWZrWlS81jMpOK7knZy1izYEW8wZuv5/mPRmPzp6saTilrxqOW32KMZWaVlq
uyorHeGQm0Bwpx8DhLg63wmdWLZD7GD/D7nUqsJMrVQcsZ/Mf3kDhHLGr7vNLSxW
fS8TXfJL++ehac5+wTjUDvspWri59FjEJ0Yidpel1OH5VlWF6zrnZSH1rL6ckCGZ
GolIZjX9E0Yfja8c76PWB9ProhO3GHETjo1XuRe8FilzUoSBG4T78ej1Tc0+Q0gQ
SgmEcZIkFVHi3WqElAhRkvlcmqkfL4CJ4O8alESxxHjlbCe9MA/3V8T+jeoTtc/B
ahnakRfjIHTPtSm0ATNtmVqalj4d0oMv82pQvrs0OW577D+atOIWLAIB8tspdA1b
pceDeeKkWSbr6bQLjmjLPhYSZiPhQsC39zE4YZRlsrjRtYLoDEjCglm///ZpJPA1
94dxXDKrQKloE5XfH1g6llcZMXAUMXog44VtCOgDBNXy6kdHRL+q1B6jGqAwmgNs
Y77L78y8rBUtnd5SbYTnzLYFa45/x2WOwwFlKi/LNoEM53UDDCJtVIhbx6ENM3j4
tYpYr0flWe1vwq3v6DdzxuMpwU8IUqMeFQTYY3cpZhM6FEpCwf54slgt33YZOF+m
q8CzOYJrSVd3zov01LfIs0W+o36KMrUaq/HyB6xgs4KjpyCUyF4kls2CRE6YocPD
OcJyT+ky3l258kEwGU74CNayCHFJYU8muIHqcHVwRJEUMCr0l1gtAbsAD6Ju+iBt
ntLvsta1K5MO35AUJYbKdFORfoVCt7XSVjP55U0fkCle0h8fDuOLJKXqKC69RgAv
nqI5r4L6Bi4rZsT4CUm3wLThiBFI1wpm5Ncq3P67GUg/JXw0iEi6qrEWMjjhEhr5
hctSENJ+z7C6xIFwZsHU/PS6VdMDcBjdkT+INyn0TQOoMKR+rbI1Z9M4BVu2zRTX
91+pA+0Y+FQzSwXt+d5d72ERz769v9yBtEZcueAY4TlQYZEkRnlZaqLIWLWYkEl0
a1qdtL/sPUMtMbhYRAaR6SMDwF5+r97qs8RHLtA0rPjxVYwoPFu/nf/GdbVCbf5e
fiyFP69kbcUuwZayPD9sqh0j/x7/bB9QxX9v6vJP+wJ2GdPQZNw3W81YR4H47NL9
msn2FkYt/kNfjnfCqw9O7eicCRc1k3vH9FyZ8YeeTlPY7RDIEwHOGZYG9YzrqtB9
lwpJwzvlzUoFKg0IT0ny8wO9s3qy+4k48Q+Cfs77o+w5Ek/1Noj53Jl/s3X9VF34
r+tViLFrzf0fVeT+xQNKStTsuErvsafDe5E0WQpe/FP9xedJscCDyR/BYcG8Jo+i
gIWvkWVoUhJ6JCnkDXws/Tx6N2ddQ3U6ci8Yi2VZZy/afkJloc+tfqZt8pcuXgDX
+3uRR3wkf12w3x/0lk/u9N1cnAP7KVal3i0Og3NOj2w/Aw4REmBxZpRIah+4cdX7
/02FyMogzGVe1BQFWFj8IajeX6NMbn9VbWy5LQxJqT5fCR7P0NPu7eZiufdVAbMQ
`protect END_PROTECTED
