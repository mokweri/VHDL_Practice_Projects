`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjssCPQnLs3kT20J1p0yqdsKe9KwRYXCXUoOK4vfVAWGifml64GlOBTmZ4ngaUYj
csEarGoFHrw220jUf4bchTte3yuG/vMADbU86SlIsUqdQP8DSFUKrmurpDVoy7dH
C0KjXqz4YIT8D9sBT2g/ieO+0Y0HkaoueXnNl/RxsJSh6xAFIcBRRgM4zvSdEQl0
3bKEWw8LlI1PsgqQ2A41rjxahneoJV1PRKcKyJlimfVaxUhFXgZK6suZX3On3nWW
9RewgEe2OZTE7vrL3jOJD8hJJgIljmGC5/z+RkLKmH/djk3TMkmIexx13Wx96HjG
15dXY/fcP3ToQFNdGJZYC/0kfethaVKHuGiK+Wy2gTSjwUr4MjRHNsXB/WJOZmQ+
O77yPiec2/P0HzQMJhgvqBK0C03kv5H6VSmk9YGvQHjeSUxlZR9kKLmm+iIDv+tR
iOnrBdak7HpI8L4dn66pP11ISNgHl++PkfKvnn9J6AqEj8L6CwoPCmp7GPwcb4NM
TdNsMC6lGtlhUoYWfdDMBe78SlqwDilod4sPI5c1AXgi+V8hFJBWqDLYnij5l17U
oLZx/3Rrkqg9kKs8/85c185VXLloyWXcfWgXsfOTUnm33l0TXWnmfjOoeGs9VsK2
nuoLbUPlG+TAIZbGsgu8lMTe+jJtlABq98/aBGMeu8KAPF4eNG2OMCTO7xpmvlQj
XDISslexmAOkBgYSkmdjHKQ7anWpDVTWq8/GJnTWou9GnarqeHAQQtTRp9sEaF3U
mIK1QthShJJLL4FYMBsU73nbNmTUL9XSQ7HL1XOKTRauqX7t3KXBusTdvE4A6s9O
QnuyoOgsQY+ExkyjvtQIVgywKPyU0geTugbCGZmtBEQhRvA+inhbNyzqkr4cIuB2
2aKOE7iUPDk/9TRr7QR19g5xQ1h3L16Xn/9fs941f806WpULspQFOBdHZwsbYadJ
pV2JVgRJh7+KkhmxOIjgRIgHBvMOxd39Zt6FVoJf76Xjt5eMVZvypcJjKpJm7Jea
2J1zxHDaT2eDWLAPCxqDRnqyRmslteqpC8lUzXZrJL78Ad/8iL2f7nTWKYypd2iq
ua3yNpPgIEUaqBUifv7BJOEkEgjIAPl27IptaEjDEYn0vbXcGbtvjSi9eOUNhlXp
wvTsPNF+Ft8mp4M5DCytjF84WICOok5su0pWJVCR2O3Se99rHneLCpLV+/laK965
ZzcVhxVq/fjkyc+icHcaOe+GZq46grquOlmP7JCj24/Sp/YqlvOZCQSdL5BCmMqK
ntUi3VPfqQsm5+j4pPD08p6pR3Fm8NPNS/gI9LQl6iDUiNxQtUtiah+FUf7LGcZF
AkuQhE1POUiIlCnnPcDi2bfFIOn91+eUnJldolrI+cQjM9++QC4089XKMUoT8eX5
AEuUWZdnAzh4FpX7nANLEOZvkNen6r+IvH4bg99xsfl+YlW46vbtSSPchvoVM/ru
LVGrkaY8AJmZcevu2athYZV795V5nialjxvmu1C5TDnv34rcGHHDWwhlG3EknBEO
vbuKUSNqiy0Nwc/jDRKQGvI8GEzGQWlBxh16UZ9rauK3JPtjB2Iu2p5pXVHrZWvp
xF3S/0TaWEKGV7JrZ0o4RodVmZF5Yjcho88C3VbjMwTr+CFlmkr7amMWAbwhWpJ6
3ANhZy80K7+p/MKJOUQwluTGtut2K2jrXZGWg4ROnFpA/YXjsKgKnQA5sNR1fEVv
Bka/+boxUAiFco9vy63ezSf4dgfab7NyjkI9C0XLbNtV02PD2lqdzEC6H4cWqPKm
AVbIhH8yQM4hudyRDNPD5aTXKR6fzsX+1n0icqL/XYwyz8NQT/nxGkeKFQ14iB4P
F6DaOwTQfYN+HimSSXPQIbBCJZZPaikZdnw6/AH2SQBgiqkl+7/XbsLT3BsPs2QQ
1u729N96GYqElmEEKY1XuoNLIGu0zX2Dr7463pzHf3VL6UqBwnKurM8ft4FKy1xp
BtxO5YtRYJB8F4Sq9ajRQe8GVtXonUy0wGCbeRD7KrG/G91RSkXp7D+06px/Wtoe
4Bg0drIGSAJeJFFOAqsppxNTB1EjsQTRoEP6/XkGd/uG4IM96j2wDbJMpV1gji2f
iaH5thsgS+w4e6RX5y//OdAtXHtqruNi2jrKLVJEi3HVB3t1SjGmIazM+77S0OeL
uoGPJB09VtmN8RL2a4A8OLLyvJzKVPvLsT94h2tG0ICSWLM5wqglUuKyhf3EaeU+
0NCg+L2uBCxyjMu27Mq2t1bfvSCj9aldYxYdZ5v//1CoyfUCUkitBBlMte4JWhBa
/gaKyjI/vmfuY1mjjfoyycf9ONAtUM/DMj52JOaQTPIsfWeKFQkNVM06JdJ7n87x
KvLvxxvJZFKaqzK9b82mFP/V55dws2fKFmSS0x5iSwALnj2V4sL31OZGy9u5EdDf
SZhfZ7IJLl2en24UsebXmpJEzO8jSuq0Heaqz3Jm396kAPojx0SDJUlP7f2tfY6B
PKPhD4cz8FyWJVF5HsB95/7A0hbZ3U69Do3VvFjdJgWLQjdMjL4InZfNq+ohxlu1
WwkzAWznPDldQVlIc3M1qR9CgnN42nTPGWswF788Gfg0ZgjICa7e0JESb1dgXUZq
H6WhrSnaWADI5qumXvjzF0Lz/w74hM+xSHXuKnQmRJEg9BscBy/h47Lz1VccrsqN
Q3U3uCP7Cfjfiyfq7gr6t02sTPlwtNHBLtCr2gExTOXldNdjA0N1o/N580RGAF2g
1wEeTQydBxQxDGzrOo5msxbj8KRxto8MuSz9B3BOG8/cT4Im6D8mjOkfEvnXORr+
TARVURPmnY6qf7mRclklTEvDAOvoFHXw0prYXzKveOt4AMaoAACXmtcrvw824hAr
Z4T/j+0/CrPotgXvFqcvJTHks/fWDL14ZFjbNAlOGWD1hpyH5Gt0PdEyERe/LdF7
J2FYVotXrm9o88hehBloDumA9I6cnpBb7109FAmI8Ag9y02xKX4BfpmnEGgb0gIh
QiYCCysBb18lsL3IU1BPfpYd+Yh3gD4tltAWroyl8ei8Mwz38jee+ferFjgSBSyx
j8anO8D+OVh7mVLntKBX0a0BAU6WXN7C2LfH7eEE3bU+JSjJOwY12KGJHoGnoLeS
zgVY1WOgp5jsmcleF46mwd+txrcAh2Zzib1ncSgh9+AdvoEg4/GbukYr6dy7iz/B
ldnNgNY6QsRbTo2qop6vSpCXcHrUwher0HDnFh7NNa15Ry6DEuVNHpIywOlObzB2
+SNLHGCGif3jw0ebHvJB8dS0qCsRa9FkHASGRxNlZxHSWB455EG1u4NxwSi/MKsO
QZGLS6FVrXoWyfpp04qYlbLolIvQhwDnP60KmzbADezcDVn7Nz4ABIkXkTSlp/vH
7pIu14Hww1DGlQb4AIHfW3h4ernohONTNqIBm+x5QLaAE7YohGpM7VYkRU1QgR0V
`protect END_PROTECTED
