`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
998KF6mb1oboA+sMpAd2Yqjmh7k7Gz3yi46lTeFHSO+K7AVZjOXYrP9NKO3jYHO7
2mQZaQfr7IIS+rYQZZXjR5eRaTlKIYYIah0DDcDUHJXMvy4aUF1/K2fp6WOOSpjD
iuR9aI52jjVKNUL65P9MaBdJNb5Cs4zp7SMYmK3rfZMzXJuhNZhbAp/lYebxO8ad
VUzPEUKcoo6g2oqMD0aD5uVAItYYja5tCBNoNpoMEzvG5Xw0PGPVsbBJYor+HNB3
FWEBoIr1aBfmeV745hp6lCNR5clARDYd4dv0SmpUJSFhlbT4YDG2sFBFi7RDpbx4
anGllDtE9BT4OtRqUqMjt1e40VwAjd55MAWy0A8/8Bb9qPKzJmz6Tp8QcWwgpYEW
52GUethZRK4m9vXRCegs+kwbmu9feU/e9QqIC8rF4nrM1QyaCvlxKSn4KZ/sVKoa
cTN/4+mm1zQueFdqgIlVoKx7z4U1Oq1KzUtCgrhqEkM=
`protect END_PROTECTED
