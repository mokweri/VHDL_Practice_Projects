`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faGPCHnuZiaGz8Z03bn4qGjjfHWYvTFzDaioVAzCz6FplYnG016vXfmzM3H/KR7+
xY4eaHjR1Jua6GCcxnvox6iTe8qA4fCLjtltr3Oz8tQLN0tNlnxuoTgVXNn3vAiy
C7PDM4TTQpM9x2IczfMyw1MmtCBPPVBmYq7ol6/WZBr8WxRjU7YCKf2p+/42FqiJ
obIHBRWDO8tfuhnH7ct0GSOlCdhzdBcvH8TyZrq+wPxPkn3KxwLGrHO0+18v/EGB
Iq2qa7LcbOe7inrxqg3C2zb7DsrtsKNYDuv935A48bMCJan+xF/kPlbS/jz2vswJ
dI7zbIyG/Y46sor31hWDrIJj3f+yW5GDRdwVY3nCDuIzaZ8a+s2qVMU2AVAtjk9R
4lLD2swQAAB4zRkTzjhFu9dOymDmftrUhFRbD70/LmF3ycMDJp43bBOVLtxrajOi
tiyWl6qo1lku3d5ePTIgjQSiep59NAWEzE0V8shUyBbF/AwBp/8GuSDuH4VDHJk1
czsZVyU9CbZPskzlZH+iGVhbtGTR2crzzkk+0ceI/qiyGXKmeAqEDUzWqY3Nwdwm
01z1N1un3rc+Cs5KhHTGJixJ3UyuNzgaD4BFEEWopeNTtcTBtlmWLGI+p3zPEHKe
R0zMraNvUFcy/dcN2ed7fbsOfJm86Qq4AnTULRDAVH5NPSvpg/PAHJltEMTk74hP
JNMYlusdTT5zWyWS1dw1ePUqknl1wcnqJLRrYhvvwbJxoR9EHBuL0HoFpxY3LR4N
YTnHU9tKp8CLiXBaVXTSe0ToArd56aCtL86HSwhkop98JSgFtbmNQKLQHKKaou8/
T9RFOo2LstDKVw6pwCekWE1plI1XFEd5dHyVz0nYwlczg0eU71T4StzS2XgM+gbK
cYwUiYGzQdffqKldCG1Bfx5+Stn3fi7dLI0T3X8EFQAhB95gXg2vZKE1pWRRDxqb
C9SGcM85Optt0UNyHEGTRx6keW+gXNW6pM7pQbSXvvfHW0VqJCQWEZvgW2aaYcPw
Za6ynqxg4yn9MjmKyXCUw3cFL8hID3aI8yZgs12QuI2cy24Q/tDl7aQv2YTAQEvV
bIjPg5eddLBHuBG8sv3WvsgmidVQbTQ81JiDmIfMr2ql0TkMpSHybCdUDsa8Rt5I
C9d9FRIjS99xmVk0EROyjV0XC71iFNG75DQP2f/SFOxkO65u2k4y4G/kdf0T/PDa
ZJdW7CbblXqYzLxNFvLSDPxWsLSX1PPvYkx+z0kCDvsA3H0k7q5cMucTnyLGUWVG
Oo9o8USpSGnHWouZeMKTsWWU1198NEhGVHA3oQYBZmsbv4YWytKyFp098rrwClIy
AKGPe9tPGHi87lMEcOu9xXsiATxMKSOy86TjZ8AHKWkdTalYiOtUYfGaEab3Hhgw
WGyNp8i2nkZnLhUrzoqcxl+FaoQKMJYyJxAtNmt8xcz9r9O1MwgaKrwNxBdAPeG/
IJOKh1pnyhK0MklSbfwgaBYTmMYNCuaCe+G9FWhpHhiv7uiJFzskK469r+//F0+B
VtrRlPwLj9KL6iU37gbTpQHAygbTXNqUM068k+3Z7LedR8QV0k+GlVpFMdkToAsz
H9owLmtRv4pNqHGyQw6sYvC89A+aazkbOnkumGYGLTWmFSxX/Jaa6I8kH+jctSWY
RN57Ol8gvMp6i6AAthIjaFTeFF7XMmzPwIHWmXEPqSZyA670QXf5uXjyKUU4n6zU
M+Jlq5vu46NCW4Q8s083lSFki1ad5zWXhdrh6lEJl6yeltEZGcSUz0HbSP/N0N+o
poEYvq/PyfSOwdGHdvpYaEb1dbGuGnwsVdwl3mcCTXFyFbXCXpwzeZzCNYszSs5e
tnxuwczFtP29Yie2nKjZXaNYLa+hTV4opNfAHBbMRIWeG6pkcERUB+6JM4MBlvDn
miJrUryUOsg6Bv6f2iyB1O3rAbdSbz3MkwuQEfFldI4tDKpeyECBPCWj8jFiNYgZ
DImcNlpkXwVjUyL1HFTVxw==
`protect END_PROTECTED
