`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8J/91WBsgSI2rwJ3WF66LUF5R0fnyim13m7ddvYXxar2KOXW9bc2U2F2a0HL/jdd
L4QXX6mMpYONkPcv4V3fv6ZleIg+7dgp7HdvkAzFPhZLDGWNT4n/8tpYjqFcr1xh
T8VbO4BcXG5pzYZTW2C28tsLYSd6sIVXQiq9C4AtyhsQXSl10VCY7o0v22P/6wBK
id80iCNU8iqqV6x6QPe10072TKXWKG5qCcl2pJkydRUci9i/ocjEWcoc9xvt8jMB
MiWsuS1O3QartKIWbLKqmDnSgsCEaCag5gQJvP1dBaq3qOXHHU8agVtetmT5xAXH
FQ0vt70PFcTygXlIC8bTYkqJrAtIcK2DeWI+jhxDHg1xmDVGv5BIQi2R/jkvTAFr
yHv3RY6V0cW8RBlj6ulmFrXn+WYuvCL7l2S94+HvUzwroUoiLj7psuI9nrKN/Tni
Bg1CCSGIV+vVBpRaR8BhUh2sKxpGA6Y/m+RaRO6tpgjMD14OUntCjHh3LljC6Q7O
3tkqzWPl648gF0/DVslvc898Oqxxt4xADb8KWX7ILJSrhzLK1CxII7gs1y/ZPvlT
g/khCbm4PAtX+6OCyxWg9XAsntZQfwq8Y0doW9rxwQaFG4/B5hjLcRHjyvBXgo4g
k6Joqwg75K5h2gVVRshhX0xoYz891RZTG+dKFs+xmIL755g5FU5vW3UdnhT9Sn3v
Xs/HzdXKWLzeYlI2HCL6vXzNRjr3qKI0cEf2e9osYIMe+g+3z3EleYQELEA5PbhS
49DXYkHT65sNJAjRFQ8B8CfoyHMW4Tcsi4c27KW2V1HSN2dQNaDKbB94P778C3Gy
0zi6jTdnDjrRLMYajXbuz8q6ynzGr0AD4dvFbscvXXTc1e0RrvbhigkLVpv0DSLy
Cr8q2/lbD2pOqKgj6MzRbLdddXEC7NwLgvFGhBOMi1hSaNZ6CvdAsOJUgpy2SkI1
Nesaq5BPmRbbfvWjm952HR8y0T75CtOZtLiX2y+F8PgEAXs6xMIsDoqkYnF8odJC
4dyKfEzU2Q5LgGonRnBXl49Z2pWcY28MMLJHbtZ+w9Y8dKJ7e/5J9+ED94BGbm4v
S5vN1G1YsTMVk8eTFFRjlV6WAukW+R/sgpqJuFC9yvx8KrZSA/xv27RIKtS/fX2I
ay2sPAf8/8BeSPzPKKVpstjjKJkuWJ/vnVeRAxeaX4bgqogKeeQ/PNiBMPR4JTXc
JCsQR39iVtVKV5pYhBxIfFz04Yao1IjcJxFO0P6BOZs0pXdFCKfHJZ0brXfjgaFD
q8GOh5n97lIkULy9mwk8M6Bfa5OxC/YzVcikBEe8F/vtL6eti2mNNd+KmgHYuBQP
zRWRUageS34qoZ6N+paaz4pY6ss40iUkbLcGkRry0/xfXMG5TUYROuf4LZksjjlN
tEk5bk7srI5t7WKQsNwAWuT6iM/aaaHvsntYQ0hHsBR1SOCv/BnO4+oJlTZG1HP6
3ftFV3iiIHZ4JmQnpSicJLtNlbrW70+I23n4auk02rJlP1G0yfqdH2H/cYcq2dkC
ao8BZtG8uQ9vTVrdksnfWA0/4GClIa2F3roD9fCGntAn8xzh/odV/tOXsNL3V3G4
4BrWCAhHTArXIyPZMagY9DBGa3B+sDC2sh8GGM91KBUxBW2THMFonsljjdlHhfdL
VACl8MWgvfq9vQQY9L5n2b9sz8OT2KiPcL6FTbI/QHDHeZrHNBuSCqq/zo2gg5D0
vRVV3jQkb7qXXSjq5E+M3Nn2nF3h3XXmoC5794tvtz81OPkFNRnJSNyfvz463/oa
+b5i5UvsUhf+8u1dENHBO2YNt8AuD1Mo6ONLvQSr2khdkcuV4Hu/hhSM/rF5Q+93
1z99hcGWg5fkbIgGrKYpDdO+7XpMZpSuo6ioxOYvzrI21Vx5OKiTb6TDLFQZpdqA
1TAshZztJciwfD9IkLKOL/BxBUcfcmfuCsigsoWw9pMvyyO2/H/X5YnDsgrTkuCS
Z1OEix8BsoKDxLUrHGjNkrvjIhBEFKNBrg36Lom7fzsl2xtd3gWtClbkZ9JGbL01
VMSZhLleBJ1aujHVOeHcUPEKiqyopztRO2q3mgc2oK+INOhY8qmDrZALyxy2oSyI
TIrQ7sjDH8746kJp0n+z85xzJn8vz80LpNs5eRXgslcgiCa9QFU/eNOoGP9q88DL
+J9n65wwyP6XHQL4cYoFUfu1DlA+KKdWqYj+FLBVU3w/QHyV8StzL58N5tNP0BaY
u5hNtjkyM1Ws6JUldvIPmU+yC4AjJ4SbivWDv4qxBBD9hjQlZ2e/EMxp8k7uKj+D
K9y3D3ndNbNdSRWu8Nqft0xIvVUaI5C7rIs3qlknl9KX+7Ql1zVsy0ZAy0V/8/nD
Zvw5wgpqwP0k4lpJhNc07WAUqsdnhu6As6vyt/U8nTKvmrwcHAtVQJanKUidIz9G
laZFfVq3GuY7hxMfDJVZ8Ca1oKiw6wGxNPslKhfH2hY1wxMMP5Dbr9VKneU7hKV9
63DcENHGTrQ0od2JGQkZ8VWZSlfB7GQyJRSHNX+gHwYA6H/RgyT5A437N5x929Va
GX3qxdeHgvnY213sfDzBLZNdccJAaZcXf1BiskFe+0N5HMs31jdhmVxgx8r0gf8T
j3tCMa5NQwQ5MwCF8loArKdk0Ni+Minsq9UaXVAIHvO3VQE+nQP7GlJis0ea1531
EgD7R+2zLiR8YR3ZHfoRBRhSuO3Fo/qrXqW3Lz9Cz4F3/U7OCUMu5gofCxTgdpxq
tshYHiskjSqyKLqq0ONp8lWoMae/sbJTfe3rJrHnheTjz6v8avwp1mL6mbNZOYif
TzC2Ab8qxXZgfBeCQ4+5Ciw7pXQ7wzcolS0NzfipypD2a5BUq3FyVeRjEwPTZS6M
/VChc/6CjTO10r3JfmuTpr2vAwbGBlb4XIL6kaIGIQFsHVC6Mmk3X/h+y15itwku
WMx7dLFSvjPQySFHaACMoTQhT5H0zY64fRkmeZSLTs9i0R6s6f0eOhvyCgIT3mmr
4I2vMB5AWWtZiSx7EDVRwB2U2kg9FUnEhYVLU2eRi0Udf2ezudpim/2zUCSHLsfe
gccJ01uvgOvwQ/UZzdIeREneOQRB9Ik+WcFvPHxThjAT3+diqgU060V0sFwYaLKm
mcKCOTinkvdegRTtNVnSGR5CXQgyMHzG5/qsk8btdenTRQzw0dUQSEstZX2Ayb7D
M4Wf2fFGpMxHno6wvSRER45LMab2FIB+KK4KYHNjwqcZxo0bb3nQZ3uCGtJiLd5h
fBfejPvhN/D2frzjv04I9OrAiLzahPThTCcBxukqpCzI1xeaegPf5by2O3xzeSLJ
R8EvSJuAKfypiOw8TQaI6SQ0ALlrn1LTObqRIt7d7xrEUK1vJa2wPh21k+RquVTX
jVYF+DBTqip6bnzqGpLTv4QuPLBdn1Podj6FnUcPl91abStZjgx8CDY+n3Qy5Oea
/smJPDDtZ4l5C4uu3SMwol7AEw9dHK95+4MpT8k5OSdbr9OlFs23ezdtmnH9TfIu
iHLAQUFH4r48FmBtxUdvWx9zXf2pqjIIN2t9vBy4KNyh01kxRp7tat0mU8RUvVV4
JBBoI2tLrHZxtslT/m9IE45a/gj6IlKEqkXDSwR8OlNTXnt/MR6Wici6jNTteYqj
vEktlDz+Y20AKk26cHjSXvAFQtzRzT1vQ9dX51smfa2ShXmY3O0CZ3ZsM3dWZ9ks
GI+IOjNyD50RguEIkqVRB8rYhzEWoc3SDJSe8kzQCr/QhWUmpWNAcH72+VikMnZ5
GGAodKQ8Qu2Br9Yh5Mfm4GyGsKdAsoFVEUs1qPCCTGvWtrfPbhUvcNw9IMouIQHV
TnB9PvUL73XW7Uzf6BhEviZZ6+9F9nnXm7ms58KykPT6zxIQr3vmKygdPwieCmFW
QmdkAxr6UePtiettrCOhd/x6fbOMT87trTNa1rEEavajJnlT3SQAPj/tewVEYcX5
ZQcR9jeSfiRN71Xja7FbvhOfFcDvNABEa4cuGWsj/Xk/Isy8RXFR+x0JVFMYx+IE
2lowUUPvmjjcVNqaAlK3KxTBNdvKh9b7bfiGKSr02CRdZbiAlINsYS355ovunR7f
V1xe2JpNU7WorIaYMsOIy4GHRjpb0M0g/d2uSrwbmbEBibzM3wkzJjzmrm970AcC
F7p4JJRkBSQoLJ+1+KmjMejm3pFSL9dbqkT1r0eCkDpRXg/Ci1ylfKPHiT23M/ul
VEr5BYIr/x2X9oOgtwhTlPhd2h+U2jk2YgTtq2GzwwBcNGnTZAPSMd5H4+Oivslg
44w/L2t1uc9JxMjv1B4yUerFpBVIOUusDx45zyqpN9ZZwIfLJbRRzd9Fr0s4/hQe
RIG1mPAOQQtW6tiCZCy5OAzIRS57aAOvphH8GVlycZsuwUNRk5j2NoU57FmArhtl
teh2UvSsAOFcKwsKjQbzlFYhiSx7Z9uBN4vh6Y9uMP+eWxY0pBMmYBBF8EoOfocp
7uqKPa6RC5lnOdKpI4PGdrBsVR4F6SiAHY4VNnYHapiPw0VXPkjZGCCk77FC2d9F
ytKcRSbaHl4mSe85nt4AjYUXhc8dIIcquondTw9NxP9t1VCiHQoERMytJ74x6taY
kR5IVmoAq+PN8MFJOO/I//uwIrwTpUXSndc1MgRayT7FBya5/bkKofu5XeDvuSU8
Ihja/AV9Lkqydw64hJZRP64vDPL8KjCW9zBS42xe3J8aqhgJi7g6cX3YoCAeATrR
60U/l52IGPyPO6fguIVb7yC5JzDJz0uJ3Fpg8wP+p+XXL8SiU2fHtoOrU4MihKUK
gWsf13uDhOS1bkcZCV96VXNo0jaHN9PlxnRPzPMWKmLB7vf48eFp/MNSIThJEkcD
Rp4wM8JedLPaoAAFGajVfwGiAkLzRSnWTyWXEP7x98TWUEwpxM9tXOXEKmw5OUVS
NPNBUjbHeGM7GRaFRzFYxphJe7UcB39OtJ3YLndUqbrruNLh7sXBoashNhMLAB1O
KT4dd5SgpoBUk6FTVX6rbruJnFdBXc0GPNqMLdG04FOVOYAqFhUg3GJHE5SwwOI7
eSPhmVjif8H2nDYup2U0SEZoUTgLpf1ccHGDgOBtWBVPC5AEip7fMtKh/wvsvpJQ
RlUJD5XEDo2Oh1IS+2uMWWEdxOyA/EosRvauWwQQrMSlYyEx/2K6EM4MM/0BqVJp
eWvrh5BgxAmzP0UgcejjoXhsqCX9yLyveDFh41JXNJ2KQNMg2X15tYBozxnxJ8mv
c/Vpx3mz/axUAJfCaVGShdgk+Iwb2GF3U4qH5JGSzjIzg6NGG1no+NkViGpVVS6S
G+EmhOps1/hWd+R1s+MLnGgpSsPI1JDedlfdAEH9RFMam8IevduzkP5+BTRiOxvA
UToz7zmUe1oOoM32v01jigs3ZudBN8uMTzaO173GnfITTEkTvcOhS5kuHGTaXAlE
MEzeGdFpHQOfFuO3EK2piRnQAJPop1OVpQk71gSFtycVry16lJgctjSWo4CZ8x2U
DzJA+H6KiqWcFnEZfQRWPWaV+XYbjXm4OZ85q/ixw8sV5TlJP/CsrBYGQy8heCmk
8jCrCOQrvkF2HmUc6ZKr42yyNMESF2ZZYSTZAz/CKsQIzajmlyhXVir6OJs8da30
tbqR+CwMqN1mtNeugIADpMJ5MZ5KOAadSy54v7gddA5ZQe9bbFR13bp8gVi0tHPs
1TEWvp5pISuj4I8LACTkBO+tQTgrGcxTWNh4hjRDPTHF1nx8zgg5Z1AXEDDTn8Jp
eGn5CDyt/Vd4fZvnG2cGh74TMruRQAydu8VeXWLSWWXjfDguCZ8ggaskPegHMM4I
ODO6PVIV8IaXeCPUN+tvmThP6F0ydlsOvnUNAJPYunS7Y+u1nu6NDu/44PnjlyFS
MIb3npn0ey5IMgIF9SsW7UtgFdkRHp2O+eimb23ioaqMwKmpkykbWnN/M18II0Rr
pTQxE+LpnsP2OGlMICwN5fEVELPtEjigsYvRO4YCP2HC1Zdy+v/5PJZjzYIQTUD3
H0HjWKwg+OCQEwOpp4cXFuhllEiVgFmaJXOV48lkJDi7P24b0PuzqY3eDWqj6sFo
Qm/2wKb1dgfEntUqXJGXeqGnkZwGG07u5ABhRxCOQqIavyKCXv0ydfZ7t6r+QHcr
7uFlaZ+NDlTeyRpFHbljvyNSm1/1vqIAeR4amAzVXvEpnDO/QMOdbLEdlYB52pOX
Y0kNvQHhNVzp/DVNN/SZcpHILh7fTreYRB4dgMnJkxajluDVAYeR2L8mylnSWPaq
cOaAu4K18fPDsDdSEZkabEXKMLib7ZeV0e6OezoqEO9cBNObVpQeadVorZRxxeTK
Q9BmbsQ3zFikR7LgJ43K1CIXiY184A+VoePkCVP7NGvICaUvxdMvxalk5AUlYUWI
yuA4KmOo1YmxgV16YLHf/R2J2ZYPHFC3zAbRhl+hE5AVYtlPc7FrEQtSlLeRAAnY
mvvvYTogYaQ107qrixMaV8iN6KwFh78Nk0OiBpFiaXyFSLTPCuu1uAXDe47FM96C
cE4GDm0WO0Oy1eVdJhnFRp9vSrPH6YaB0JQBwYGSFgSczMXYgOmUw/btR1nP8ArC
UvrAIZtCM0vq7tPcm43eglO9OhfSaqJGyR0pSU4xrB7SDCytMY8/viEO+4qwLSiU
42UoFwWmDs+j548ndTEI7065DE+AYMCzNrLa/Gdoo1kJE2c2tqtRwykWzaKDyeG7
v9Hkd1JSBjW0CdXqlNcPU0mMwPWGJPAjgbQMWtm2WXuxEd4gUZFtjoA5t8I5B7j6
ficcmLg1Pn88kjVU0VMI1Pl0Ta5YrtcO/gGx0PWjmplBBEdvT3c6eI3Lkfp9F1tO
GsRulmP+kKGnyB0QLpLHGW23W6Raqfo31M08JCOaLyLTuGZZ//9CzNkh4FXt7qsP
Vgghe3ynTW/7kwKWJh6SMCU6JIZeeGHnP0QjPc4avjfDJuEOmQ579b2GXAVUklfn
nc8/nOQKSzNnPd92GQOW5gp8RjHzfb8tOdM1z/pnO9NdpyzLjRDn62o7vDmbjCIV
SIIR9Gno4nRMqEhUnWxgTn0M/EzPEyVTJv4OUbqCqwiU7az4B/2f/fHG4pWqwo7/
i/CtzPDJqHMOhk3ZSo6oLqSt4t7dnorj13EqwvPzqJILa6OGRAFJl4lQZt5unSJO
ftPDIFPmvCj6xq00fY0Rr+NB1oQxLTlUuOTHAiDgB9SGdnddQGZEyRHb+JujvEIs
2hjoMXq+vTDDoo/hYKumfQBu2B2KIRJNfCytPM4uwXrQGvzh475bYM3V9sY1dBU9
PiAUUsWs4XNxeQxnabA/H8SBZ1+49jLPMz3J9l5aSdCdy5DSoL0Z0Z33vw0wBcB0
8h2eEzDZYaOIX/gn6bIcxvwznR3z4hE2urtihIeU8M/iYkcTVaQU+W0fsmADSO6S
36OT0BEVMriDFHYfWRBtoGXPmyXi9VgvFIkKTbw7gWVG+EnQK7PF8rktZHZ4UZzl
O94sP2GxIf/q8OeU6UhLp87taZlmyCJzsb+6Smie9iZcHH5SeFQIgCh1y6E/WhVd
5VQsIWjFXL6p6w53hza0L5e39CuBna2qLZgha7ofUBlqonAn1xIvRrrOveFupjcU
xPOJ/ZqjVD7L56Qel2M79Bx6y8+bNQ3ADVm4xoKSu0mzc2Nxt4JgPUOv0EXvaYzT
Ndb8NqC0rT/8fubyUm+UjqM+pzfrHIV+xxF/Sm6AHN2KzoIAOBUJtGRtOB3mE5af
bB8CYPIZBh2b7TulZISzE3x1oazZCfO8xgKZacCgfhSEWyeWHhruHoz9JMb4vjcS
hixBICTxGQOUr4zBIvw8s41UzNCecgYpOw/QksGYgzL4Cqfm1R3njnIgHImbxiYK
/9/UN2gIKnBkcY3YIs6hKYWzWkdd48+2aVD9QEZrKzNYcCcC7X6pZJEmO0YulZeR
fYF/yZVtoScFkq3h0Q2WoZZpxia32XwcG9D0wuInpv1zAZ4enD3iB9iKUloHFNXl
Jmu0qwJMqjBWSrt5yk31VzKFDXqmYz/UaVzpOJPq0iNkvHaXdLP/z2chBPrrwvDc
Nk1qbVxv9QgLxoz+PddSAHmdQim8A3lJgmYsWHiXbnfOKTiufFXm3pb26Zpm/QvC
Vnzgx3Cr8CNIqBVFhf7mExjNm5aswIg97gLib5jLDsbJfSxeeQxcux8Z/ao8/3KS
jD0NdvQnr/6gP/OoxMHmDpIiLfwnAdpAOU8LwejVJGMrF+GejWF/oA7M/kFG+cnp
qZrBBQC2aSIjlhY+lwqTff+9mgbwBJW5WWutF2w6oCNH9gXhALAJQjTNbXkVXDnO
phwZ1dh5Zf7PRDMVCuEG59SfHLTKnKSIe6XoHW9hTKe4d7h3tGRcVL5QUqZndpkN
LSKWYKK4YSw862AnJogw6Nz3gY24gCfs+UlzFrs8JBxziNOM6ktprzUyuFc/MUMM
eV0uKuBSeXUsbZXpm9s8TaAtSSG185dtN8WPGmJJMDgNGM/QUpdg3oGR6PNnhHsN
+QW8UKEJ3cdad7GvtPNd5D7MROBhDw1/cfpY/HrL3MC6Akf97nHrIZD8qLOBJMtG
c0D6lt6ri1W5E8318+GV0WzerDX5BxPMcMHwwWQDIO+jCFESH0LORjvhRcDc02U+
OKBzC1aCvxjw79fl/cI9D7KkaW9B+ESUp5m3oOazJQMsL4qaCxn5t4/zKwPefsjH
zozGphJQyu6/SKmbdP9dATxD2Rdef5xLbtJc5ImMvO3vonHxLYJH+XlnGR4Im1xU
Ldxm3OepWsFxdH5RWCF9nC85v7YnkcC4UHTzIa5KvgqywlbjPXxXfA5UcAygzDe/
8RAamxfevZ7BtEx+mjB1TNRZ10wKj51n4oFQ4jn+jKe4FyFh6bAI8AV0k5pNi7CW
B2eyCrCz7F6j7o1IXMra5Tq0PyHfoT3RaziIzYBPyQi4birms7czgyVCGX5+3pb4
xIB1PcmGEhXwVWl0uj0lAUHKZ1bUCEDWGOOBrfkHz4SxqIzfurUGEKP4PTQXJ/g6
gP637rjSWIPRvsXjZ30H+5N6Ue8tXrdrwT12fTzfGpqDaypvFxKzuTToVNu2Me17
UXR2hzGqvYZzkKF/QVbB6oL0HGBEN46sISAsNl0bxaHXhqQKx21LgQq9Syt0bo2y
i2vv+QtCRHNCw0dWwIBr9+qR1aobpUI3bqqFO0WcXSVgy/lR4JLlkpRG9dNqwnWB
CErwCjOmCpkth4CijlLXu3EanndtOM8MdiLQ3vaTErXmtL89O7UhI8gI6TucOfQ+
YE7FeDWPax6AkvB0DAo1drJThsZrbs7KNl8q7DQnAPipOqkdGKmbhBog6BvkPgHi
RwaIMyw9vZNDFJOzj7vsv5lGC2xlIuB+uuEgWiLSjNLKmm+PY0n4K4de1X0xP8Jb
IJ44hNOJxpFZaPOWjgbrvhNc6g5n6bts9nMDAXPtoZ3TntlQwMJsWyHpVk1kyhNB
5ghsIXKDQpilRh9LNN1j30fI+30oC/DmRMm7lanf6XzrJ+VdX18L0zun4jVkCTnX
cVhDYvc//IWC7iTA97ewJJCdZ2pYYx6ADCgN8S6LkyhSHeyM0F6r8e3GSgE5FJLl
ff6YbKIAVND/WtkPHsw1hOKRNLK0dAbUGLsaMrtcnmj93dfE2/0vgMkTFGP5p/3+
zc+Sbdhj2nv8EAT3H1Nz2YSPre90OpapSjGSzX0ly+lQWbzXywnT5G776AGrLPYO
TG7CZkn8xDjLOj+JPsl7lM6GoohLqdsVMCg98XUTpXsprthkPBUtJ+DiWni9SB7V
71ZPiMM8lCLhbaeC9sJPO1ozoJXf51r9S9qVfSUVZ1IZS93nmAmTLhOuOr/+TG98
K+gd9/QPWYFX3sDU7wuUR5TNeAkwqeylD8ttuNmfxurwV4tAYnOFJeCykO5B0RHj
jLCsOen683NpQTz3aQAtaFgJV8nQXMjvd+h8YKnPBNoRIIdedO2xpx7o4V+cWtJv
Xi3MmmV5WADNH4QJFlMDw0Qo4lbE+/eeJsbdWmdFOPDDJmTCI8moQ7bJ2+9AhUOP
89CTLYPcI/jT/WarZrbdS3rdL52PQcKnfMdOfob3krwyP5KYqXzLeZy5JZFE2lHT
fi1uuxoTTZjk+A3lec0Z4Mxm+WcxmS27XaWHn7HiSDm0+XnzFC2z84xgmEq0wS3C
UMh8fsDjmEqTwSkkLr6cc1DvWRwght0rqWIpCjRuxzYV3QytS1dF1ZgycKB6b01C
I9MX1u+r71D5Bk176s9W7PCMQTrU4Mj/XrzOuXeJaHCZyvrTNNBcNUzUF3pDU6p6
aPz4tkV8gqvJfcq5llZKAM/dqftsuCX8R/iPtFXEQ8HppuKIlbYsqbFv/xFOJot+
90uTau2+A66MZK669d5lM09qaL0Wg4WdFVWApHBzbtPKl4gEjA+nDIGLg1Gk5pGP
skjfbE74mVYRnIpgfd4M6UvMxCYrxK49P1R9YSlL8om9OM0AZv3XEbX6mXJmRRnc
pQ0mGBgNR1oNrHQWkgHO9nGZ5W9Z//ACKROhNhiVSgIHvEB2Ee4V84oxA8JleozX
p+R3V7FOudp1OO/6/ao2sP9Nolqf9mMPmHB2YBcpj4oYFiIQbRla/fbLh+BARs3g
mS4/87PX0p2iJ5tHhV11whFLlTPMc6bD05oK2oV52m8GeW5tSAlddugIcESIqynb
GtXP4LJa0GgTrggkz8ucbgtFaxk9Wi5baCYxkOrR0CV3PKq4nbRQU5tul/fsr3bI
7D54yw+w346Pxe8BorC6cFgVuN6YY64RmXF9NmMzDa5+kXznyA2gZ6MDtkska5QN
VZecP7H8q2aYYpV4aX80O+VYxjgvv6BLjSX6kGCDMCMM7wE7m9iIeZ68yxSK/7f/
8JqjI0vP7SJ6wgMIKHiH88r4eWSNMvaWTrbKHjBuHxSusSKNeh3C0MTOjxenbHgd
uivSykMDp2uOGB4d9y8KkH0TgF1mL6bMwmrkxIfA5T+XTk/y6r0r8pv6nSdRiTG9
dy7JAHKFb1KSG+hJAm07fU4knWEvkyCQC56EJgpvIbjDdQTeKsnJrNTd70zmzLLo
yFcltZEHHR+S5dTGcnAlaPRjwABNmL7SNpXmD2IeIx/VIbMnfFUXCOzkRheQQo6+
yks/Ucq81E7RQt/P96u9NsURWpnM5aZLJIKSAl9zoiLC+OLRmyGDBupEelovIkbh
FfBql28jIhJIxnNOQhRU9CJc7Kvh9EGyYfrLLy/Lnevx3Z1L+n7d02gr6Pzu1VD4
WFSivUpACN2NTujN5AQRB0aLmR/9m2Gn0TiEePRn5O2Q0qEYlNPSV2hNSR3qLc7m
/7IB+ZHh/h0FWt1i/UpuWI641JRqcde2MxzuKquJlIKYciBy50HLP1JnyHS1CN6/
VamiN6MdR/78WLoPVLmbPewBsHLbtnc/XVWF0is3g54xFvzrchbWhGN1FuaiZ4OE
woXZjYNEVARdfqbJxYBJnmxXLe3wytaR+zwfFIFElXr8Ddd1GdZLFHEOV0zEfHY1
VqFww1tdvl4UEdUIjHk/IRgSGAR+ekNMZK4QPhYkI/yTSptpqUyCaMFRLC6w8AUU
/L/RpOZqedffiGDl9sSHCi6WA/uQug2qtzWYtSVM3VzDH1I8wkO2MwbyZE7aA3Cb
HSdTi9rVgeo7LYFrQPtBg2ybPLSvlYsy6GmAu8edRxGI7oVVjnyiHslevl52GG2U
WM0F7oGo2hB2NdO8hQe5kMevYuYRwkB5NhmUFzzhFsoegxO8JYnZH5XpqV96XJHV
SwnoXiF9J7rBT2B2yEUds72Rs9jA33XtTQt+CjNa+e4TntSjfO3VtIMxMsshnBDF
3bCFvudW4a42a2vs/IYjN8ebaSIX/wlDmBJjh898jxCG5/06hv7ec+iCu+TIkfrr
oziQ+VcqyRQwi/bfimdfwutxb4qW4VrbGLAyGxVIFwYqulj24P93YPzts2V+5ltp
gv/T/fl8skLBlIACX4TA4skRmypD687pn1EOiCpqiEtTlRX5g7o9Tm0ler9JXTsy
tRKvPhm9w/SXrNzvka1YRGcKn2wZlbNgo4sAE0kiK1RyF6W31Aee6jnOgOZQ+oFu
1B4FfhAE3/gjNjE0uUtoZesuiBQ3wK7+pSX3zDH38bevJj6F/XE2heZa9JxHmtJ0
2+Szd/rwWwQwr5xIvj1DJ2A3uTJRrdi3d38Lk8xQcxcOM4jUz5BIeO3DsGXahIzj
4TK2JDUy0eppt1GOzeuMprw1pgxkSbL698VEabDdvkz7hgBMkopOwjDyhjtLFITl
9vDvdFlccNBWcfneV1RzvPiTUVC51GLetLruQmSqN/wnEZWTnxB/4wXqamF19AoM
3M1Q5hDae3Z0eOJak7LG/XYVoNI2c8nQb+taO2TJQjav8H+otkiKgjjMoE2oBQOj
sGWLO3JhROKzG8KcW3/rL/pdJGR99/5jRPMGZ72kwYqh4fu4Tdy0V4hZMNl3ij25
JZgvTMY4sq0ai/5gSfMxHx7HBNEhXjZ9wGgop9KbQCH4wwz3y7IqvVUjgcleEbJ4
Sb+xxdMSXRkNUo1hSvH6AzmM3URLLG9yytnoi99quJUZhXL4UeJAFIUCsg/TIUld
o6iMRRRuPpM1GIUxNyju5gZg1VAm8fcceqLHWJam143swLVpofQIpO01naN2BL8X
X1CwlQzB/B5IrwkyJrS+gwggs03wdNZKG0zeEMc4y+wxS0S0xCfuy1ic+GGMYVhg
e/7ub6iYzGjsm6CEHiwNsLRynxomKeJ6U4hY3QAhfrtWiEyixNGlYx8gpsBUEOkl
mFXTnJONk/mEfp7/rarR25NUHuAjTiJm+wM4h8jyLROkLElPsVLwRJ+oCs0/dRJ/
q7u9fQNwdaYz0HWnBwGB+VnaRtPrsYoEDBzh81/MDjzYkf/Ga9wOhqllZ5tBupgG
WaXRgBYfoD4rCt3qQrn0t85i1UMtZCjcR8jK0lhbRFZTVouZBs3WgTdFqnkSu+RD
AXvFk/iQ1fwZyGId+FUbYISlQLmh+Gz1f3vkMXxogqm/rSbkNSiP2WWpYg3brOi/
37lEX1byobPokX1gVT9awd1akicDBtDm9C5FFo+aGQDclJxzRTQsU+jD8/VmVql4
bPn4FmUH724m+xpSbaBb485/NPP1pHVNU1EURMMem6NaDd+jsCDK64oOUGSHUUMp
WRIowyqIFuDwrq7/HylMtNxh/9kiNUbOgdRnVyerfMVRkh377aGt96dBQHRnjxX0
F/FhONoab8e/+Iurk444+O2+7GXROwyQ+VM47guQrml2lDO/NFb8Z72IwVl6XOKr
3khbPng0BI/pv+opu/MW66ALB4V/odbHFX8JfzKCmftaJpzM2QZxVDA4q6v77u2I
MZsi5E98EwDg7j0nxu83JrMHEJcePWIFnM5s3HRJdshC6Zv6En4wdBJGNt31Soth
lx3OQygCfoI54Pj6Lc8rAVMV/ErOCd8mYTArLAKSO8RytLRqHYcGvyLe0Yf6Kl6d
WVieNaFI3Hmpaswe+ozwBEJ6zaUzh3crzcsNlpzh1jL6/n2mAjZx2SXYaNa4XRAV
lQJZal1IDN8JnSdvd+ZS4qzW9Fv3vELumOx70XJeh5ML2v+zLKeAeDiDrKMOoT7t
aofb5YmjSoGRyDrva3XLCEhPrQW+Gffi+2UUwK/JV0cqvz7b2zc0aTzxFBFZG50v
FD1Q7vcACabKS0yqJjKcRd7cRDHnjE5HmetUsQ7caJ43nUQ/kTQyPWBNaWfpX6Gt
LSY8FgIZhddXbJaco3tzat1CsHrrVFaQjfxCFAaTjg4lYgMjpwYIAQIrYQAeiW8l
Lbme8a2GcglRSQDxsk81Zxrg2hPwqbFZQdSUsEBDt8lLTkGEulYlbWiDLrvNO4P7
BWUgcJTT2SSAWxbXfkWrrfw2KidhmfTTJizdV322Mx10G5JERDZyNJLe/5i5lyDi
VyQMtW8DC6jTHcNoBxQr3e8PzSsh8Q0vnGj4U6HvVQtRfNRG18hKxvICwPqe5sjD
iwYgwBcJtvIidLVDt/xuIDNkZ0aigXc28MRB0V7sJ+uetwQOj3RJCIE91l/uyWt3
yQ3CRJEwfCEfuHw+ocVt4FKJk8S9SQ/82tMqzv7P06B8hSrbM3gp5Dx6DCFVvbhJ
u2BSNI3E3m30JgwwcrHAlMXmKT0z2IaCvL7qTyzWAszmu4t1t0gwCviufEZd9wkp
x8SSFjwMZx2C4WcXJOzbD2UNRUYvqwk5gHo6LjuqQErT7U2hp1Ot4qGIGR/1XpWn
7pVMfaQNmsCfJlyWVbxpoRGa3D2rIG146ASmWchKCj+yqb3BJAUWHDafglc9ttbB
JCnSv0ncD1ixM2227heYbn4PsPxCYHnRJ1VP4MVMtWV20+n1a4wza/15G1IY4mFv
R7JhAKnuO+wkIPjqyekN7rqiLiiXiU3BdngS8vbyAN+wc1cII2yTWns66IkkWrYQ
6rMdoDHtxEQIIBt47VNGdtVJ1OvyzZ6Dr1zVZ+vjM08oBiaCu2J+dBRj2PS38toy
IHPSFPtG/Xm/ez2CS4eqGttuFsnsJ/qHVkCcBUiI9PaX95ZPR9L6iNXu8WHoSG8O
/QrvewDELtAh8vvYj6lGKhSklAOb/PL5STvmqY0D5/CTJR0mV5ef9sof7kM/0gY4
jq9iyKYBrLSis9jj7HhZRpcE+qzoTQQ9v65tZ0XZxJXE50Axtiu3/zeVWYbl1yGC
XlK5UezOnXipPKOK7Un8EOIUwZRj4QGK7rMGKV6ZPMiMIUU920Z2MHhUKqoVOPNO
CaTu5ZZs2FRZAT83u8rm4om1IEvZZC7iQWHxU4AkVSiRPnYqzwfhenGi3JQ8kdCZ
nVJDPe5Pid5RrwByI9gbSU2oi8eL60kBReKCLiKDL8CuSh20Ot6KUE/sQTOX/wyK
bjCvshQdIgCYsdxyIpG1+GkTWDpJlKwYmUs1mdPAqEMQwR9DS2v+3PNxWEzYsdRv
uY7zSgHuBbzawC8xAmVFguxyXps8MVBDHttQ/+GmdgtVJ/G2BpKtH1UC6SCc31ge
79BqO/p+6iqZegmaBqiPsXpDrJ+LK6vOyorVMnTgRuoY/qXBEpt0kxONIGJF+8+u
/M6/ACRDyIgfapn1nkj3vOtjdHAtR93MEqTFrjaD3LVI4U1XTNRbf9JSfLlapIJb
IagaFJ8nXJLuUAU+qEkfOvnFUGGMeKjFCAWmk295Cg0VqcAqEFnzujccs5A0s+cn
8S+gN73qv9tBBe/b+w9DHm7/5QA6nKZOgCB1xKBUqH6KCxIXY2DPZGexmIk3kR10
CKToMH3FEtCeuemW0rxR7vx3/POrCjWsl7YTRRnujtPeBrUheNbzwUA3J67NFhSw
nDEiooM7GAwZCGW0Jl+aARqigUECfvzKXdIpLkLU2DAnJalIvPFFLz5udUqj+vH+
7HNgWrJ2E0ntkcYdovMlUhM36tTQC54rPuNN7HCX6J5C2wDZqg+Hlzx1u+X7v3ah
C3xy3DCETWITyjqU3KGEx9r4DNBJ22WkQeN2P7IkhtqNkWEaGd3KD53D/SelzQEc
OZ7EnSP1S/yu2NsEaVTAReqbjw94fsevw8hCH59f/mfy2yScWnoEXKGMDbez0c0u
5JojiM/E+sprTGtg8WJtA+lht7nFjvpPbVgdteFcXvu4kLLMkN83oI72ShRhDVeR
EugCXlVELeVYnnAX/PrfFI+9ARr3Rksuuobo/aksTXx53JNC8yIAojFs+rRh2Njp
NyOLd9HLViMWYsLPopmlkAYtB2A6+YQkZgnBUNL8XHOZ1KxU5IDOJi5D4zdIn0PG
WlG6g2y5ctvXXeHXA1hzfdT/rD6mKgeXsvOJte0dmh2IPqj3hQXwlH+pGrf4/cEk
vDLHp3gAemdxHVmd6bnQzGOOadl/mXzYTwwtKRxCp7ELPPUEcntE2JPTpUQkgiXR
6tTAlFUQ/CXHUH+YieG22jkkQQCvl/yAbeW2xdSc7gN3bXdyT8Z+Y473qPhAdpHt
87pr1RsT4tkJ28+dMty59xqA7Vt1/4VsAFRU4HCW4KsxiTAS4Eqq7dxXhQoPsx6t
jN6ecJJoJbHEUTzozH+eKAqNgN1WUuL6PT5yQDDPuNI4pObx1OX3eeDtljiCTcA7
rkw2BxY+3L6OFzRfN4jnPdrE2GYXhLEEnmp26wEW3zXbiMf0PvP8VyAYofXru3J7
Anh+mhjVcN3uCeiZosKjpavrRubea+kmxFudpCXzsOLCI7ejLPRd7svvtzwWfZhJ
QDWepCxhlbEn4yfje7TJNmtXe5LOQYqVZxPnCzWCV1XWj9RSsc2KTjx846IioEsd
BE7/o0X9xZ7eRPgpTj3Llr0m5UvRIbuAE2wHVIk9RfbThxAkt6hnaUdV+vbdQeAz
50b3QBNRs2fGGxnueZkmiR1Jhdw13ZPSJjeNNF4OyX6id2rVWatf1wwQpsExtpLn
Xt4+rFLYz02l+1G71rrtcCB4gfCmQwgY1jg76WFom90oek2akvmk++rSM2FsApow
emw8OWxXVhJ1wCoLhWy81thAqrZN6BlQ2ATVgkh+fdtYqY8zWMQPpnD3hu3Wn310
5kG3CcuFASNQ5NhsVtYCsDotpxQqrXPA4C40CSMiDDya/ccdk+LCxhx+x6GQaZjc
GAirmgyoATu5v09ncfdFuCEKRgNWN/YXLMZ4nWCDVuixNaNdem57IyiZ0iaw/NJ1
U9ZK+X+t0sV1ocnhELpABp5RsxeMgQqh/YNsTtsnX7WVIOSktT3kahgkCGa+Hi0a
/q3Z6QfF1ECi3l8Yj5Sa/IohCNkNkldf77tZzx8hzzjBTlj8T0uQ66cB2TMQMADU
GbAmliJUhiRbju7mFdk8bIRuPLPsr8cKK16dvrkLn9IJFAQFj1fcl5Lfh2OAB9FE
HlM9ifWkV5bSPLao/FyD5v4ZKUMcTgHcastsxtKn129pVj8J/TYvA6une2TMxAll
+35aoeRsulNL7AC+GNMAlCyc2PJsD8pFrDbVA/s/YuTFDPyI2il7tQsXmbOgNN6+
Voc15OY106B6zb+zzrt8hXgKJfrm1aI/19e0iCM7XzRsVOa2HKUwr9nepfJvZL2N
+5dGbmZminSgEUsFSPnhf4Th4cfPugoJbE5jPmwj7IqGXAgkhLfJiBrk7BOjTzSY
KA8pGTFa28tfM9LuwM2NXS/GuiCafy7/VliU/J4PP+V/FGIEHYWxk9RNCfkc9VSe
8xlTb1Tixwv8S5qhjogslWnsZF75+E5ZFYQyXZhZKcyXsBL71OTeze2+J8K5THE/
yGYdDcwuXqGD8cjg3TnZ++KJ+3Ju7ZipNpnfD0Yoqj3zw6CpLwh/CnO5dK7U0p22
9vg6kQoXDCFNkvCuSj2yPxxcLK5h0N9aiQFoyutHgFWtSXH+1lL6hAlHn7zNRxk8
5FSM3ZvUDxDysAF6+UwMVsGuIJLUZqs0uUiZ3WsopSz02CuHPgZe/rKAWnU/q2FN
N1m5EekztFU9OVJspJrxoXUwKPQhEXZqJ/egXAj88b1fIB97yzVbovXl+yBRiqJb
P5u/E7N9pM2Bb9cNM0iRbiycpTbokYpwHni0fmB7EkDMtE7S7gr57a11LbfZaYBi
vZmXZfR8rEjGPiykLl3eMWMuuWP2lWAAypueSuzkHV9JMIYigYdP9FS5wjOdrVzS
eVqmND+QBVDYbB0Mkri4GTupo8v6xfQic7RPO6JqGA8uT9jxms0jQ+BnnGRvhImA
Aa/IyOlIUzpxwurzJifbmABOKI44fyu1Vs7HRRvoE0B3uu2w4uyxqIgO2OIKWBJ7
KC7CALEmFkD9+RjWlgGLPqTxI7a7Oq6jxsROrc/aUrZftUXXS5ModmkcQMz+fMsO
EF7vjnqM5ejEtaEetrwY3CzmuzvJOIOVzmPPjqkq298cPU51RMe4iEVxTfy3DtT4
KTbt/n8iKEn8lT/rVulA89khB9g5ZI/ib5yrXK0qmMhW3dYUt22CqiQ4l18K+c1+
rOcn7uYHDaJhBXjAiCEq7+h95giMsZuHycAeWUhx7MXdyTHAbx/QNsF23FBCEK6l
FbCEAK/PdO+czI1YdHvcd8R8CJS2mYa7/pbgdQqsDtN96qIhMyBDfHKmsfgl000k
qYf89Mq/DrUBYD3N6zIC1tiUcIsUbjpBxOfp//yCzculQFm5ZjQX1G27h2JwllpP
S2iNLR0SEI91n7OzlfHBf2A3BeDh1M5Kqq0Jrxlv9z0NMMx17FAP5rrF9I52uSCn
QJ1i/MiTdeo45wcQ+Zezxk7Id/hO0zgSyEU6Ddzd4JV1EjMkryj0mavy2PXuukGR
IinexbN0IniXAafNRYjgLra1eXF0lvP64xzhE4fc5TeNnNQTVJ3Zvnaabkm6SCfC
FZrs/v+Oo+n5xb+IdTuM0nv08E+ZAuYyubHuyS+sqw60Pbh+SJDvYCaenrNVaZ8n
Vj7cx9fR/a9PtKmPmY3Qm0X1Iyq0HZpHZ8QxRdrsOYPp8SJ4KkYjyP8radmUDwcV
pp0fLcayUgwQjcwWONBOT6QmRyQ74Z4he6Voe4E4gIKbq3FrYOq//nQIdgD8FaV9
nVr1ZQFnw6PTE6Xyk3TuU76xhUbYhdpAzq8rDIyefWZ9yqFVstsnhqbsqLfxgF+i
2Qb9uWP9gIBtTXLLSJzno+vQrZ5VusrghvvTSpKgI1/Jz4Dv1O1B0YdzRAw3fD/X
MwChEHyXZ12qRtsuwvlruQUxgj2RBE4iblMBBa+/DDESYbn8ipDKoYigduBvU/aD
EXFqKwh+Hqbe6kvhfQ2ns9r4DGlbtjwUEW1Bl0Gh+XoSZIJ9qjCE99We9Q1MJorc
Zr/EEIqzCIP9Jj1vLdb9rxG0awzIR5OgByrSxo4EfW61jw662ZUUj8ubl0dH51Vl
CPhQwAvlFgtNS2Vnyb/ttSLxfEZ/GgQ3v73FqAUSb9WT4SubnOpQmy18oiuOrwqk
ntmOtweGbPAC6HFH0Tle+7R9JTCUq3nfc56xM6LF7mEMtvIgOV7AOYd2qbeGBiCd
kN/ubAcqMxLH4sdkgR6V4RsR0WgoghDsDp20gd3wF7ldllTv+BZXVZCJe31PbGjF
F0vtKl2d3UdvcNh0IZqnBA3VKjX850K1q7qIKorekwZxHUT6oJyuXbI0MTn/FbF4
Bms9qZQM68W229AWRaPQr0Cs+Jv6YLzhHqo+J6TGW0h1GO8wwN2Eg9nuj54FB3sR
DY9VLfvjUakgMxPXN/Y7ExGHsSUIdzoeAhnVa/3oKotfZ9BEEUIOSqQ6aboUGpay
QPOlBZLUq6so5dpIHZ7hZok7b0y99v2rEZcF4Zl8gYP/G3Xb4/SKQMBrCDnie0sn
oNXIs2oqqVJkjWiarbT9j+JkUdEDQP5uXz9e+yiyW2PCn142B/oEgbDc6B5pEr9G
GUGWMbsf5VaE33bco6Mh3mqyAM4WTNXp0jRapHjHFJ+wMzI6/ewb/c2UaeILg2Bu
XU2NaFqF2xeFg4YiSecflx37bvCanzGDtshWXn2DSXzJJqBho1CpykDdSKXYbwFU
R01oQIw7odeSI4ehzs+WkvxMfXglde9FpWMaWBABqNbN4x8akWaNOMdosJKbScYs
eDIuGTiEHYxkPceql+Ho20e5LT1flh4jDmHR7OYQqFZHSena8mzhXY9iq8Me6TdO
3SghvlICO7vQH6LXL+rANnwu6O0xyWMnSeMI89cPyGFCVM68Lo6Nk4GGhjp+hfRb
pCSB0awb8olKSEZGt0/MXFeFeRi6SIeep5J9Tpqh20sOMdMi336+EV0lPhMaixT3
rJHS/wTiD3r6F8TbbLsqUp/J1rrlQB7qcSG6OyqiUaKnYDWSLgq8YMcL2fUE9NHb
j6wEUdoo76DfOV+fC3LfI+iGfMSGHQ3ahZSVVoBuPvv6MqjX1w+ou6XitE910VPS
m3l+A6m1buHMbuFNssLn2ClNasbiLZrPDKZOvnOWWozGHe49L6jn2JcYJN0I6+PK
6jWD2rtlvwU6yJhFp1L6bXq+ibt1q8VMLND+Q5H5ZpMZS7ev5fTPpTJuDsHJM0f8
f40uiSxNGWui7PYktpOuwczdX5j7Z7TNMDSzTlUJYQkAMNzqkEyGtEvEU25X2SeY
XFEJb5cM4+eH7AVd18z0qCgqRIEz53aph+sZ0xnZLNsD1iUXEJ7eXencUftJLADw
w2mgQFTy8ej1Oe0wc14yRqJxdetMhGVMFtte/T9qHKFUHSKMp/t8rxQ5cxIdzeeT
inh5aR48HfaBJIYf8kUmQ1ZzBHnWWYZ3nFniZ40Jag5OD/hCST8+ADL+gTepIh/F
vpPC8I9yZ5XR/26KKYeYDaLM6Rh575RfEJXDaTulPsj15DSdwbFicvQGpZXxwPb+
gtZlh23pZIxLIDragCaUKBsmOf869s8r7DOIU8qM2n7v4iPBmhr6jTpBYgeADTv0
k0IqcMzZHujV3DwgvNNezn3V/t+7pX3JPK+TQFofcGF27941k3IUj5tYt2Uufq8q
W2yTX7MZB2PxlBYmc89HKpsCgB2UHjHawpMT84DkbUmxkZL8MXfvsZFEPxjeZXDN
iTt2jf/AFmB8Lt426nzh/aLttx2OG5R4ObxvDg2Bq/xqu3waQW9hm8vHKHbfGaFx
lw4P1Y0Kcghvu/RbybNUYJolRU0QXGRTpG25r7QXoP1iJ33yosbKctwDvgtwKRpA
DJ2PN/DRnpNJhvuRHxI7mPFWTcRqH08dL8zDPcIAe/FtQNe+vBmInqHctyrTyhAI
B79WSbhOB8GNE7ocy01wRcbk4RmK5qE9DxXrTyqhL67Vk7D/YnG8+DUFj5OteQIb
PE64rC3vVdu2tXIYEXNvtGzmpTQbdK5qb1XzOpQOeXyqNC75XcFInaKCidn+0WNq
V74XCwzXHAGzNVnjFCONd2X+GS1+UEbZb0Hrcl7R/crXu74YiOIh9drsHK02I0Oe
LAsR4w6rAkYLxRzffOI/mKuVrTtNMVXF7UQsV0A6GY/vMMN8edxJCcmERlsJdLl3
mFZVvChzRu2gEoWZqPP7ZMCRzLEz6N+0Lh8n/2p0//IQUf8Y6/qdMSU7IigCR80h
4phXL0ebY/d6vbV0RD/lIbXayI7xP3c+TOksJiGWpfoqaeaSTF3I6eONfQOn1Jtp
SyWECFzTqYVafF3XmaBtRUKMp+9kZ+QDPkfH3e7CZDvrH1GFyDHh+PyHVWmJ77UN
y0jGMvwpqk1Iw1xAk5i8XF4Ai8PO/xZuInRsCad8I9ARLjbn5/3vZLrdzrzvYB9Y
/FvzeRXGJBEugBBnmfkQT47Wdh1D9CQsdKAvchTgHGpwvhNOAoN0ejcBTcdhTUfB
SgfREScPE7x8fbPuITcO8RNBNCh8Swi4CItnm7BjSmtnbhhY6HQUXu2cilsOq9Os
A/F4rW7958D6Z/1q7nwAo9Izi4qFsoCpXG64Jcue7ORiU2oP90YOouR9AgtSzmtX
Mzp7T4/PEafGtYYpSHD7ngXS+q/wcWum9omqoIxQmyCrbYUuDSTTxQ9SNtEN9Xzr
BQ1c9Qs6YoKhATAykU/WnRFyuEQi992YhxgFwW0b/OMvR6RqQG63X/NytZuQkX6y
8R4e8UJtCXL5nDPWoL5JRV1f9OLH/CTTNgbiYNbm4xTwPHrdyT81Ps5jVtH8NqGk
G4FU1pwCbJLpw8SXjJhy/GsTpM6s/cSH36l9QGGv/wltRKez75lgEbaeC7eslHq4
1htLLzR2WhFhxwKrA5SC6VKRl3iO0tls5eALlFDmLiMyPtPJkkkmEvnifZOwxxk1
vkxn6KW/JDQlG9MvBkzv3Lvvo41eSpG6yHRMavuCV2qmntF1JYqooQMBJCdea60t
QoCq0xGW9y/AzylbiuQsQh0EnuMkcWtvZHPsTkw5qrRngshx5rPCHXmvNTtKttbL
yW5K2rtb1ROkhJgKebXhb8b1d769sr7KMYI1eENRlof2oVmJuEaMRJG3BeFy2ND9
kTvFZGXclAV0pos/Z/WHGhhMgE8ahgh9DP+ome4dZptYm4HhT1fPn6io0coYWJ20
QhILa1TpeGE2e+bnsleM7k3gN06DlkFWUa6TjYzbpQN9G3JeY+MSZLkXLcYCtEJA
th+AL5IkxbAO7V/+0EblVc5SoLQDOsUqEmnv+A9nzfOlGhAL1SCNnRwtSRst4aZc
hahluNOYPLLpyaGkgkpla63QGwbqesiBlRFS90g9tguAs8i+KwWZicwAmeG0oo/d
+k925huK8rBx2Lw4LbKpBb78zo/ydB+YQmDR0jksz7EOU6LZ+odkj7/Es8KIsDKc
vZuOuTWFW5JMhcEOfNJMxQ==
`protect END_PROTECTED
