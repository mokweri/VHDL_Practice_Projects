`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73m3K9msLXLQM88t84bCZuCjCfz969Frn2vuUXAovE/F5YmkYEc/y+Hk/ts6P/gA
HTJm4cgs39SLdLIJictGjkUTeTFSuzSfv3y3JZPIk9HIAo81/7Kc1Pu3jB2I7pna
ppnkavaBid7NLwaGqojZEufSZDj2s3XEkjGXKIzb4+3Ke7AkALO6WW9XUPfFxZIQ
Yiy4651FHCL8Po/RRVXSn943qHDp0w1++eKGr3GUbvy6sHM822FmRnykPZjbWb6e
E7LJO0ulqvgTQksP9GPdKwfC38Xgky8u+Dm5PQdnI1q7YWklcipKw1XWL0P8IgfF
L7Yf3RmHLqFsHoO9WAH9Agy3y/pori6C+GJWweOFPddIwEX7xKfZhymQW7PIjdGO
+cguI5X6qZK3IYyk91uZX1t/TeCvsKrxCPOmqVUJRmRODg6xofzxJUTRHvd5TBqV
ayT6KATYTX+8VZw7BOx3M8qFG/P/1fJTWoc5cm/IeMsIPWJJOjefYu4eBrtvBRcc
FyMNgUbExkOcHIYR0KRxv7xMR+4pXQETSjAkCVbYTVwqTl/qkAqcqX8bl8+ukLFN
OgG1G/nwK2fU37kNG9zyO0r/ilWsG96qOuX9I/7ND8GSXH5lYbjjDVZbPBb7K8i4
LV6fwILAlO2Xzm4Hp5LH25SFnEvLKKgR0FaCKp4UfWI9ZfQ3FGBAzA+ih3LaNGTy
4vBvz82HJDdih0sH7L+TifYAWGaONYEKg8TbYTkxhCl71sycV0Ztw8rgo8DoVITa
YQXDITgfproE2C4/a1IT8t9jd5WLBMb651HgmUAPawIUQ9nGbnFFXWPvdW5Vo8nJ
0WmyzTDbHiGMWtBDgjcuwc0dtZUcLb0La4F0YNWqH0xDf+OPNIxd2Ir2jiig18Hy
zE76e1MKqlk+Y7n2IaRMMlgLPvI6L9+A/ir/D1Qsm9VcdvQTrxojq0pu6Dc0ACUA
k1DFv99C+fihwPtMqTfHW07l+3cEgwnFdtlb/NustQDAco5/0oU6ZVDsKtllbJ3D
W0QUBeD/pYD3+X7NiE9nJJx7XK2CgqGp15kL/2RfMqfa1Pysi8MfZSA5kSfHullO
3lVTWrcj30q0TkpDY6cjs7Ns3ZztZ0dvUkS0Yo+CJL721c0Lk8oUOrnX4xcj46Fs
lZ162wm5mj2+5UJGioHGkk8ST+B9l/4llRcP2fl2etibGC1qTWV0FeT24riTuxGU
p495fp7cxSOBD444LHMF6zcHpLl0m2lKHIm4c7Yreqzf8fd4HHWffWO8Om3CUzA0
vIaRfEBACytIoPD1fy7RXEVy4tjS04nViN+yhy1+DiIdjn8errmOl3leSz6NLcwH
6DVWdSDhJS+UJDoAHJpt3iEQv14jc3oOeuKvE/DSVZVRmyPAhefuG+ZPdf5ShmI8
KZCg3z6dHoC2LPA5DFOX9t2C4dNoedT8jS5zd7qWEN/0eMHP17QOCoiiXaT8y8Tn
`protect END_PROTECTED
