`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DPMYnENKDxi/LPucqN4j5cIKP7pruYZ+zvscBoL4s0MLCHi/dUCqyL5Qew5TLQpq
k9hkxh/o6G9RPxlMBmSS2U69N6vGsEE64Bjx2WtanfhhG2SLPR6khrWiM00+MDDl
eLk4s6NCvYD40uPTtyBJu+1E/UOtOG1PJZ0w02GRHK5YdQamGqhCT6Cy4E8KBbT8
pAllkH92NtCRkwhMDtPyrzEGVDP6DTbBAWxRXEQUyLeJHf6P4RIGaDLWRvuGwVIg
WjboBdiz7uCKtClGueXyHz6HXsN19MXRrKUjYkn8mWI8B1C1k6DARRDPIKPnZfKv
LzrU5Jq1g4G4e6j86JCOSjZ+JOOURiwVxNqCHpJVXLevfzprmIhrYl33KUCtOEfZ
MWzJZroBQG0cyjXLTstuGTO9UjJzTxR4f/bLGiWnByk27/ZyOqf5Z1PFcxT10YtU
GSEOV2xof7n5KXxjeJwa9f647D6iPxiFdH7rZ2NRQ3qCm80+xNzXODFXpTpOW1vC
SmUxpGm8l45NY/n18FhpngWKJHH6MDwyp6E6PpT/X3qJ2OW9fKV2xd4u1NTmTXaL
q+YsfpEA3QI2CHl1L45Sfa/f+NWLqShdF1JH+LyVQvz71JhoDd0VxF9RW2v9b/9c
6w7fTgJ+L6KkuTI3wrZcynvqaPKepMEwhD1enjgULiOvqowyMvW9aa+oERQyZtDs
6co+r8w1xtP3EAPGzzGNwLoKRRsYTiPNsZy2JKa/29/M4NMsXLBv2Lx8BN++uhwQ
3LCKWPqAYPRf09EbUTUnSb+dNyvGaHu914ew6XqJTNQ2HLLOiwZXWlvlEMStXxcG
nSpE+o9B82kzIvCaOv8qdK5Lkn2wzg9TyITWBlEPHeEy9cf2n7N+dUMad8dIMea8
PuWsTl3aoGZJwqsXFQcapqvDbS+a9c+pl3wRA5qsLMc0qd6l46pj5KgSeIcia12v
cn/hH+we7Z1UvDYRqX+O5bmyRa+0jpPvfbLZN+53vMHopKNO6MZBNVZwaK3lBtGc
d0lW4QdBrlrA4MrtNCCW/yDDhFOF8X/VbzlGBF6N/GTNfkrturwHu7vRCucf+CDe
GRrtOwBmdezIdBs2ZafVIOlu+JL8dz/84ImHtlOkZ/eBg/sFddBnNeFuBKcaMPrb
EseAeZ81s9qB4+k7IqtOi4NMs+KNjJ/1A0x2aL9ZctTPDaMNr+zkQrHKea9RKldO
5cxLh/yZf9f66KbrKsjmy7kjfL1FaijjsfbRl+fEk8K971yXop78yW/GstkNCiAC
Wa4JkFT0E5Us0EAjTa70YAfThkRVS5MgHeHxe4lKgdVAAhnRmbHXUkla3E7eVuHF
hLtTQuuX82PV+O2ILGTxGM1mqsZOjYAl4hiK3iL1MB5XI3L7U8TYIDg4y1vz1Avw
uuUdAUUq/p2j+hZ/rP1mrx1+5ER7Fh+5TZ2k2O3wzyK38dUJZg6JeB29Wlrp7avf
F+ecEyQQdMBGMHAdM06txsVNoocA6eGPZ04MIhYAPNtJTW6yc9rQUXlRxzOKr/tG
rO/SWdq4PAI0P1rMWsGZzeYz1EKFlexhypBHK+5FTWw77X30tsthrb1mZsUT4djm
kI+OKJ+dQcJ4LgHe8dW+DampqLqLqxsRQtcj4x8oqhU+XM9AV8oIYBvQ5llgfhvs
3FSwEgDPuvG1W4RHEe20NDh5tglPK292fUXIJO3BXFmcaLehkaDu/z8nkHyLNV/j
oq88JmvUBloiN2gX8Usjsmgk9TrMbqSrP0PsLej79ZCmw8uCjk/G6g8R5Lu0b9H0
1LSEF5KMof55raKQlS23gD54rM+Fbuke5saU6o1N35XQ0HvABB4tN3Fyv9M47Grv
35AdfjUHFxcKUzQJY86Mh5b1xo2G23vEAWdHHB84m2rRNm7xhkoME26JPPtoNPSO
1R+H/zunrT2qogwaTCMVvVpNo/ngrq/UkLXzR6FAT+gyFJl8s1Mt6uLp6fhTGudy
jm4u4eBKgnImVT6fprIBa4OvmASSyYz5zRlBhUtbaPW3TFdU+vWAweWIHEkt/FMq
+ghlk4kHFSIXtOuqUpj6bWb3+J+yuxXzbrznTr24piltmXj1tTzdaNX6yvxIgmg5
5lJ8JZkKAc4c+ej63fqxqtld+M+tYFL/zVKafn0sp73li+1xSIMmXM5PnS2mAcDQ
JzeoRu7ENdASy5zl5p7xIk6SGA0pazcPiZOQCeXL3HasRos11ghIBmrn6wb0Wmpz
U9DXSMa6seIdzipkzYQyK+zpjehAFm4BA7UoetXnLwKQgY2vxZMvvMP+InPq9aWe
vq1ugmbtDNFN+uesCDoZ7wDGFycVtiprxJ2o+o5S5TJ9pt24pEnISVu9xFubQxRa
VTMnsFK0lGPY/qLSucAJeDmucGh8MRheIc9ckHUTNIWccsEcYGD5bzJ7h1tjhVhi
kIkq2ee/7W9yhWjbbkOWOA7D5PrysJLGqWfkx11B/btDByRw21rpEfKHDoGtQTYU
DU/RZIcXrp3Ufq4IweMzD9eZwXeHo5qJTC86PtP873Bb4ebFa8xRcs7e67lXa7g4
OdB6c0TAeUEsUU9AxE6I842o+xr+U5u98AGydb24mxZ+bQCE7WquxDthluIqCjFB
qa27XF3Dk9foiKWonDr35ef4Tyt9bnsvHX1oKjWWD1ohtNHE81Q0Fep+1s3WLulT
0uwCuUQhpqD17LCVQ2Pk6D6753lIWVdS65Hy6p0MWfXIJBYjZWQxe1j2E4uN9arf
uOsXZ29MVuG+2HfeFErXrb4ariV0YFezTy7LTKhUVo48HC0D2QoCzGubROTVdum0
/+Xc+CVMXz6LrRFJY0Qw+B8OEWsCV92CGkss2TBWyDWPMBIlgfTN0Vhy4EssvLvo
TTCHEAUozUT4zaHDaU28nEBANQI5d84CsdvGyIKNkfqBb0gyKQihU3FMOkwZN3sg
GOTKM8oqp//1us1iZQ8Zzeeph40Yu3cnv6aHBgSlr4+vyEatw0Y0r6GpsXEPwVak
4GGUSOzyajaq35lQSnKbQ2XhfqF9kfHMJ9zKCNwMfLmhETBJgHbEBwmLsiNYOzfN
5pVQ6HrTvFQH8o2wxDfAVzHyg83N7iEbHS2Gjf0vZ01NhAYIwWx3plek7QcthC/6
lxbaGECD3nJQMTGDdsW6grz4Kjopn58zSo0O7c11SBsh+h780EUz/TPn+7oEBIG4
F07B4bkP6EIoqCxGMVawjkxDFuSkxidyfKpXPnY0cUHazQOuQPYAlpNmPIudP1QC
0Xo1hhOUngwpbOxLSsghnvxbQ8FxAeRx5QMO36ZRg41Z8xLn0OCXClA3cX7aOQVi
VxVJBEPy8H1b7XoTLL236szFnFStKe/fiEx2gSIKdAtKptXY0RDFpLqXJYVmfvr+
kjF0o2bHTWUDjsDZp3gsEmWpeklEXXAxJQ4s2vqHORxdvq3JT1yEhl1/dqsBMong
GQezFgZmp3MrqgBxlX/wVow7DW8C2uvC9wC/Lf7iFuFOgH5cdQBIOIuEQECuuqca
n/kNK9F92FJBgHyS1YnWZqFoVJnZYc5/QT9vIO5PlxNCuJ3k3Yg6/jebjZfS/BLm
94rutRrQpaTPvTIE9Xgh7OVV0ahhYlaCJQ7Xu37b8Ygpl60t+LfHkpMu8G9XqYVj
8gnISZqg8VxoDdjodjJ7AiQ1AS1iz6yyiCX4H8zvpeJ21+yryyt6b6PLhUi1LVkn
IbW/HPrJVLqp7jN9QvPp+Aea6CFt1WXLAYxAJ8p3hUMOqbcscENOvE+fUpQF8pTX
wTOgujf4TIVo4U9ZKtLpI0m8WMzaTt8+1PLaxp+Y9HBTCCqgaqysC2jqM8a/hn1W
xJ05YM66wh0ZDud8DmOVEktqC+jYXiIAj51ZIjSUV1lUS8xUnkNoAImO562Gll2S
ea7j3ZpuPxOMgY+EJ/QUHYOWQlyA2ZELCuNp2eYwt28c8CaH/yJeZn/kjNROtwE/
m168nfQcT9g8sBHUQTTAp4qQqMW8PdJOiFFFCnlWXa0l8R0LovghPMaFckJkWfoh
YDfZcTajgltQFdyJt0LWI+9jf6w7otFxoKpPzpyVq1odEHIzyN03cl8hxEHbeyYI
8u5Hw95X84icKZ0iIjGDksB897RLyKmp8x2w5Y5hkPD7gDCEBpvxA3GyVD6Ka7BL
hwi2Q9bQbM2fGS/EGD6SiU36G5BGglyC+jOprZ58jwT7JVIj4mA05Icisv0LdCTl
yIFcLDe6vOk3mAw9Au1DPI0SiFkX/B9gWWEXj6zDhd+ATsNlc47w+PkYulwyZemn
2INFKYWg/zX21JKcUrf1jj6PbF2mG1EhQ18XW+9vaD0btygpDUwERF+JZlWyiXPT
7aLlTSXCTf3kv8N5FWgV7WJQ9JBsNmuh0OyvT4aK+6RezM5nphOfB/vohmHJ61TB
UCBW4mJiqsNyP+tSKKkY+GljY6LHFRAz5b4IOyVt1WUt2+Dyb+5f13JdMGviGupq
YtCPN0FOX4p0FIzhN0ii3dRlPp0wRe7lJEvgZ4LiClLDmNwA5UzpMKuMqpXoSVRS
rpDIRReFPyjd1Bob4MTWreYDN4XVD/9bdwacKIvBbtdtQG5oHKPM2lR3/CK+7B+v
+LWVM9geCR4NDTx44jQJ+7gdhSyx58FWh3SrKua31iYji+45SP5B4acX7NXbSi7S
rGlSwOULB/LFDbdujC9+WozuL8xPn+DrXMIScn9tt4r2lj8HjxshgJ0li5x43jA8
4hikk9Aqf7yNyB2gRW5b2Qa0DOELXsN/7UphzId9DFKbH9zZfbD+KO/KEw1efaWf
N9GpO2L26ZVZL7xKnhv4CwgkbXymJFCnEdwdRmE0iGQtxsOS21kFlu9kUxKQufWA
JJqlhrHCaPu8YUKlOudnwciX2vRmHMhco2/qjmMpea+UBXZ/GsddEF8Di9lOT5D8
OFiSxCShjYdgDaWHqtdj0Nz/m3u4D2fMhE6PHUetNfnsF0KJdaYaLCiA3Ss6knb2
L9yD9+ao3emKbXwnM8PAwnOSGxpWdQNERLdRXC4yk3cBaHY1u+zrrMTWEOrsmxn1
i+tj+Jpf1TOJFyq08D5Vs61ixYiq9eTUclqay3nHVwm/ENYtpo4ZYeZwyjZUWej7
H8Iz3A7FyJo4avzyZAidlLmp9oM0QoQ11V3+YFvt7ioH5JyUY8yBqQuG75qiGON4
2KfL9Mcn5d5JQ0Hcw8l85rtrvKNeTsr7ZBsqYE0fr4QufeEh4yd6AuGqTlx2yhaX
ktciS3aDLT9rSswmptTeH4GESzf6/Z4exWs/xKmrF8aVGpp4YyjAOlAzPjgSMvIM
gfjDQ9+EA7fSqusGkysQyTJAghAaOJrJL6vvi4fnZPRuOmJu5MZmjOGxQAqG5rsu
VpAacCZ5KET3r4oNq17So3rm9weNAWUfbtPO3Mat7CSW5VGE3HZOQtgJLqG3H0cC
CwY/lS+rPck/fIF7EohVbd2/wDL2ZfeC72ucyJYUUI9UYXHxZoMRdo3wXq6fYBbA
nB3RLtMJiP5EMqJchQuj9+lHujeTUjoSsEgj6fcbmb2R65RImM38NI0el5e83Dgw
BKqSFHWmK9840RPtGaYOgeZI3JfaOLLLwXbsNmbGEKt7Gi4vn01ptEmVLyETMHo5
KulilWvTEoynR1VQwdrOhSgWAJe5Ps8cibRDMWMqb5Unabhv6xnEJ74GBsCN9JSt
T/3PVWhj+WELp9GPPm9prox3g3V9V043+IxRnFhiu/6aUJH2ycEGHdTnMdjlnQzw
l31iWKwjHnqM1UsprKDpKcJNb68TqCoOLbKDEl204fzf9lGURF5bICaAIJplPNE8
iMSsqrZlbSIN1iXlJghgUdPgsZOTHVl6Qh9Ynfe8vWQZcT0QMPohOk5I9ORh4InO
aoAQ/2sVZsbp/zgvz/M/7x1mTSvOC2ho6aSU5abktN2HQqoDxk0lxv3eq3QWWqYv
YcRpXAQPlXH0oj1j/ZO+lCLqqZ9KUtfNdETfQ5N2euFkv+z/2bJfpHg8bfDXIE/j
JtJlVrSu9KmBq2VHK08lUUIHvmKH14TPcXczx9LE0hE/jfk5PUYQfuAqVgpTGjPN
VgBjcSpp8AQxJO3+tcuF7MX0vTSaLLFBPa+IhGock5m/JKR9mTLQFsPg13XwVifd
Q1UEYOS3amt48GiNad9RhV7ZDtnYOMJWO+KCz3pJkulxUZxeTKwSQgb1+ylhGm9E
uc8Vdc2fJtAnlAUjEHo51Mb24upOSDmrqQlS0Rw5+Z2RTNcQjuGVIPaZPAOxeCPy
Ll6CzemxgesBCqmK4FpksPWjfyIZwjf7ooxgCXf3VkrFjSGm6uIlIZ1gDf7CKQjx
gPfGuVM2pUcGtWDGkySusrj1rjt/UflO2XJonqXVPUi6kJJJSMbXw44/cNexE9lf
NK5fb9pkgrRseM3txB8CaYcgUfOBbqrbObmGg6GJrocJypzDy781Tne1XHJ045hc
mNcu9VpSwgGLDFK+T2dlGljv4Hm6AeMhajPvkjTML854n7qsA3UPpsNvEvhjBgZ0
7xxV7hS12T0QwWguHBhF/2tbizZH1s0FJs70AEvAF1cs1sfClh2GTPlNf6Oq71lB
sgtUhdXLWJ6miviCICKR9e6GAUcBLtDK8r2mpyrQQDKGcN8AUT2zSaThRlx7/i5z
Y3Mzht8z47/5BinSNvJN90x56ybAjcLwyNbbA+xUT08KUsoCVX3p8+nZaChGa/sa
o3iFaLItgLbUlhQAMz4BnMQdMgTqJkh/La4PrS+jjzGTzRtrNIPYAMZ/pydZK+kI
JKMwyZlYiM4wCAP+9fsEWiQsMtCk2d6WKiULnZL2WjBt8FxUIjLd5PgZYUt8uyY6
gVa2UzeLtxbJ0T1zifIpqeH3f7DlMHY1Ohp6WUkQtTimS9j+1RJxXDaZv/w1AiPC
XKcbp+SF/lY/35dxLCJoY9hiBqMChIXeo2i2s7z0/psndzDPTLpflPknZ7lEl42t
z0GIbtBH4iJEhnMf7l1BWfP2lbfv5VINJjUUMNwZRzNaGhJL4HVqxw4HXOorKn8M
qwPFRAH5vuSdyReYXmnXgoHhLeZXzwe54tfY7aei4mAhk1GBiZzRydTb9YDMPmIg
IOou9FyVU4l75D5GJPsrbX73ek8KORh1wJXNddAXGVnvZqHYg5w0CFr/qJakGQ/g
zeBX+d+wsm3IDZlgDXZhhKORZgOTNDQHEj58KZItc4zoqGxl0wC9esWn8fE80/js
DoTEYArADgvDfUNAtULgj/C5HlUOoUePu70ZPA9mKYeuNQcVqlriD0Mcq+C62FSF
uVypuwmrkxMoyu5Ss8pptwOWci6RbsUWjzPpk+l77fusVaIX3TEM5PeSJ6R38mZi
m6tTMC59+3E+N3pIsuT3B0J9aPNk3kUPhClG2TjD1c+nTVlxJtCS5WF9+hmc5v/M
T0pApx1wL4em3dTz6nxcTebi4Hp4QpTAXMxd2Vv7IqpMgSEKj9MMSTYUGpaRIgDk
3aPLtOsQKeXofrNsbrjNLybY6cmgHymqyjP+rnslk1ioD8k7aKrK1AhBUPOsDnpj
/E0SDIpj65Y4WZqZeUbz/oJcqB79BMhicn00ZS2pauScYLvgg62XqETEp89x/NpO
4Q09WMw/7K+woXWpgKFjpiKbYB2z/Zj4UAGxE94yugOsTZd1AjAaClDPIEXvCDzn
RC8h3yOCTYjn2le4uFqqrM/Ku1+Mtr9PBfwdpF1AaOq0lERCafBeGuMdcaNPUeJG
8FLkmeeJTZDAx9ebYl0LzVbM7az/hl1RQsFzAihg7kMr17R9SZV7pOsDtDwS8DpX
918714c8kIlUlMm4PekGYWr1GLvGVb9x5vv773CcZGDCBfb1TgDHKzXMcyqdooxN
C1ZQC/yA+qmkY6vigd5e2d/ZnBu1Kv3TBEbVbCJ0KWFbLdUmYzMJL0rN3LiU83Tz
+rfK91070qsJJ2LPF4jKV2JyY+JoIYRFFH/5Yiq9EA2ycOOtm3bIdeSbrKhDmp4h
nN5j2e/0Fe0Wt1NHaMUeySPkYhxFU8DY63Zf0hkkBnWyrc+o/9Bm2x7c/RgHz7IO
jefBMdzGFXR+LvdNU4bYaUCKus9peGDfUw+VdK+srI6yazXZPgqs+c/6MTjzuGMn
JBp2dOeTC0tVu5jCQoBH1E1fm3VDjX07X5ZZSSuQhKTSJu2eNuXyWJRJLTwvn+Uw
04ZMqvkcZUyLYipUoWFOk32E1xFjhHJOypktBgbHWozvgQnQiV74k2hyU3GH5nyv
RI7wZdTGfh2KsDtmLxetO00qX9NjDW8nL9ofhzFmUDOPZqGznzvxSrEot7ip5BmQ
iB56RuNfwqhP03oatmt6iNCzmU5excjm5Y4TjOsC4/k/OG2TqM36QC5lQZamZxjv
Z54Vsl+PolgnOLOnofufZM9/RJdSTx2bWWx4jZbTQChIcwFfofI5LtAyMi+APJ2Z
Tlzid1QcNv3yiLthmImDpIFcLSdi9MMUXNz6d9oTM8u8k8uF/RTf6pwRm21l49Pg
qkiUncoSbESG3K0ESr+thFaO/NkMCvHXqU9PsHkek0dcQlVd/drFm51FFwqu530e
BZi7gZRtW8UeRe6OnoL+uqr4cSEpTT8LMRQJP0y4xHuE8CtF7A+bNNrbQMqGx6nO
5wK2PtdxwoQ2O8O407If+GIXgx7jxkxfQ6KGsfK7ceaPAjz0LkS/XVTMSNfjF9B0
N9FbEcvMIqoJalvdV9n67E0pi4gu31ve704aGtj/PmVD3dF7nU5AOqhjAgE1Iw+J
Wp1oFmZPYBGmgOrlnDOE/HlQUFOce1Xu2dSCn/krVlEOqDr2VNHegL994l5duMAW
ijKrkotrrxDBLvuTsv9rW8Gbb6I/11XHq9StbDZavSoXacvO3P8vVPZkMjnM4XDX
5JuVGsqGc1eL//L40zaTLqyknU0gysCnHXAsdqliudoPxXPuf2spmoJEM0EtIvaQ
jnC6/oAo5BkbZ1SIMh4bqQ3uYF1wzXVrlHsYBrINoZK9StqqPVGZeDshVsk5XAIV
O3ofbKFqSSaT/RJOrx6HaQ==
`protect END_PROTECTED
