`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NoqmLPV1QTZhXYlM3Lr/0jO1uJv0w9nKzrqZKqFYR4zomxnrIQtXHaznOWC+obCL
G+iFv89PnFx3AT6ABmXkqaGRjiFGrjl3q3tZjYjLzV/qjNfn+jvQDOcetb9GeP7D
YQZgJO5wfz4G5B3yNpC6aUF1z7mqMqq/319L+Kms9Nx364ig3kjAxddAGtJVqwvK
nAx6FylU+T37ciu03tPwBVxlHQlAXigMqBtqR1mG5j4lRfJO+sx4Dr5TrFr8N4Nz
Tj7FnObTSLHM/OdAkAmaGfHI3US06tJUZBzOucI1C9Yj3LzsD8e8DrWR+sTzHVtI
rorLHF9jMXelUtwVthnwKsxDjwSEYdMLDwPCIR+wlNJGa3PwuV+o8XSOa+FhFYnc
LVLK740Who4b5GDek/eLpQakzJokti6r+bs38oIvG7Xx30SMhf5jIcsYBNEzc2BH
CkPsYgGTS07VQJzwSFB4+NjSCz7VSRKmaKGHsBZl1e8o/wS2Vrw49VmqVDbV6mp0
3J+1o00HdlCtn7B0YnkL/Sj9uPdJm3tzApbv0aneq7oQwlc3mPKeDvst23LQI2Zo
nWxqmy4FFTXm9EEiuYp6P77bPBYcG2VlRQgKwpXFiwC382BpZI2CPTWgQeYN6cAH
FXhs2I0lkCjyTCtwsTaVbD/BgLSxYA1u+uhYj1lpm/XZth4bEOZspRcvxa/S1eYe
jV4vwhiDWDgmJknsg0zitep9o2Jc0jtNUkv5vyjlnymGq8yNf/R+3Gm2y/QZlTfi
V4Wn8JtmqB+r3W3MrUL2Z5uTR9lJE5EmMNvGZlouXR8GxEgDQzVc/KT8fWDIhwcP
r0gASR+xXzuNYD0Skb7PzHdKkwUsNiZ9UtVThqTwH+Umtrz0SQwiO6oIdy8ZQoLk
hlLypEMyPWJSf/kzwc8WGKUwL/P1vT4b9UuhK7lmAChSFTKwZ9fJfG+cOL6UROd5
`protect END_PROTECTED
