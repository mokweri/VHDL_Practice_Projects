`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAiUdBgrp85Bhvybw9xMHKVd0uum+mO6Ew5a04F1gFkbCfo/+MngKD6KUVrakY2B
8d4CH65nKAgMaG3x5f5W0WQ1hb3/Rc9nnGOHh293eU67LCEeoIBF9k1Rr1oAAIAt
LcBRSbrjfdxNLsNfjaeodgfDxkOvjQGFesEtnCWoJWgcC04Wt2+evIdiQu1vXod0
jwnKwDfbhUcCu4BT7DHkky/EWIvL3fPJ4HZRAHyTBjhFKtu8LkjsOIUu88DQ5T2p
kA3oQaP7YzOJGjvGslc2di1S4QF78oqmJMcikult2KZY2EBAC1ubL20G7+k5XjpO
n72UBcYYMT3ebBTH0aNu6jpRJVrRkNzg3zKN88ZEULqzPKjbBdGNvuCi3ux/ovPv
2n3wmsDeGJj8jxFm+V5XkflwMDWuC6lpTvV2+5kwE3OsK4D91nl657kunyuyOXJm
LoqQwvbnwFgGzzjus5JLgL1+czZAPLlNVytwYFKDJUrTO2iHsoR9jUkJK0aPiq7w
E5LExba7iaAmJDfpcFvoOkrk3MT2gjeWgd7kS9XJIys8UH2y8dFLJDOPY0BgCszm
py6W0NyeqUp2TKSv3nWCWFexIfeh6WPGbU+K7NixzsgZo+qYoX2yML/IxwyWL1sf
e55o4f5XUvxBqeOG3facGEfHGJHxjExP8KeyD20cZEuoia6wtYTzvTtzO1tSA3LM
67PKO9Fkym4GGiaRGHXLmVJ3OecPIyI6zRiJLjoh+yaIDK2DCgq5g+dBg8TZkdRs
UJDdBrQmygEXANoulFzDN6Ec1wvF6fO8t7PO+QKh8wStbLdy8q+DnnrAEM+4ok3U
xqQJy8PZ/nm9M1xb1PDAuxqqGe0QUCM8O0VvBiXvvzbAiNCUqjQkR1y6CUm87glT
85fosepJebi7UXzGEIgav1S0DUxqMAb89GwAzhLscP6FYR3R1SDRE+H733YXyRNr
blKKHXBXYSF5uEtkMEIMbiMSNhkSBVuHApyKXQsiPN8qCyoBnLM0DbhDmZ6a+lPg
odU3I8TFtp8nmzmqQa70s1vR0Daw40+rUjKV/fkqSN/HSNjsOQOmX6VHaRL/iF71
gbpm6Hmuak1Ny4XzokSxC7HelUxWwHr16fYVKL7iXvJustaNfIYU7SZXdL7W3tgh
KCNH3QlfZQKtKR4W4dnFHyjVbI/U0QscRUCzV+CwgXiXdmUvdgbGtbMKFztylE6i
Hc/nUh1U+5zgwc2Wi5ZEsa2K1VCuu/SwRQX1fV/p89TK/fid+TlcDEYMLL3hc7Ss
wnPrCwjQB3VxRnx+ixDBAB2+WZLxD0jSM8YMRsOYn61nIulYew5FrH9oc+3wzQST
SPkWeB4X/GLhHCBRqD7fXFixSVh2UYN9ukRzRDgYNzM4ZXRKSJDtdb7J9Q5mk5N0
nOpeH9WxP/Axy8pPJu/CLJsI6Tgbsd2E+dpHrUZw1ChKnvviVLzS0QThwpJSRZQl
0VZdZ7vclMekBxiPXvj6kfc2qNyrCkRWQeHEhiQ6hczdnhIIsPqIdbUQzVlUw1LC
vOcaxZoUadjuRB2v7iK+oRVZ50UI9soFWdj80YCQeDfzhpeo2X4yptqUdlDgGOoK
/ps/JHDLa3o7czOx0Hlto/mJTyT+Wvg4r60MYrIUoXPFkyIfvXlbQfW20XqlNb49
SpDPoMCuT97dZ1J2taekMaYZJSaHn1xpukatwpXtaMOaEVTCLPDXKN+QvmH/AN3E
7Jp4uvey19lfp6XCgWHvonxFeV2sGGbiR5kPNj5gn7tN7ZvnKgOU9+//3zHJeeV0
S1UAOdqVRiCUZ4zo+YjM61p/Li2nbBCBDThsXjlFrPxyMspTsDM0FH6/EozhT7aN
ePGYqJZetpT0YvvynaDZugdchijTHrrpb45LBgH9ZLkI+B+JlsFgjYfajae61UA8
tcKZ/VwjrxhnVBtXnGc/qZUIWhAoPjqlYF2ZmvmTKYUaV34/0wQJvDYHKfQh0Tib
C78Fk4bzNJ6bMNmXpESG+NpI7+LMBP+KjdD3e+Tr8JHwBz1u4C/UzeH2d0o5Tful
+W3rOJFhV7wQH/1mukDcrwZv9O2mdO0GGJvBpJ/IQ3A0rT96Kx0DFNn9Fqbc8Vto
p5P9mg22E+6123lyRWixd2xgRBiTbOLDl05wejGY4fW5VSFaPgetIq/g0qfuQTTS
JGJ3gFS5venxYE6Cgo7nz63ebkX6Wg4FE6u0qgZ804CXvCJXgIoDU5AgsS875V/Q
U8emI1nD2OxxLabFSpMgF+SLrfHV2BdGbJDhFn26SkG0KdpwcYdEReMyZAQV70Tw
SLhpcS2KdbB36KKkcbictj2VXy9gA4RDT8sTbjGjaKeXbSnI3cG9yYL7iGoPv7Hs
I8jOWM6krqi9Gqy7PaPu1YmXq4G6q6QDTh5dWOYmsOe1NE6TVvrCD2AqrVjQHbmX
cn3B31NrsFQkIjnIYNWwUU1rkQHkOCSJlSt5JuEqIERGiBDPA0eNAdZFHhnHpmkS
2cGY9xKCPkU4JLqHvJZYZ0kxQ5IEjEGhzvTK755/mv1fra6icGQqPuXH+7kTSRQ4
QzJ67fGqNvOzllAnSslDKvv9UKWpOJOz4wppRw9U/JHbPTdsP4uMVeYFgT/ot1+L
LDD88e2gUhUHqN7BQarwsVdtdDwDEfqbc9DAWFsne9nswj6K/vG0HTKCc/zFlCBE
KrvO3Y0tUVqg/pRoS8oLy01vai1y0iDX0zdzvA+6ChQhYoYlIdTcH9oa6lfEuScX
fIsv8IIY9raEneyYb3xouCDTCbLksz0/LwGt+5swRqfZbP22YMi816/PwsuyxTmw
3BPFF++t2PP87YMrqfl9MXOHIBZZAQHk4/oIEzIW4oq5TOD35Mme36sAf/1BPMx3
piYjFpwyudaePE9wXFaOiWV1rb//jx3mHuWwccx7/IhiSyO8loUG0FHjasmA2WP5
DKj4QfHK84lVnkmxxK80Fu34xYSQI6Q3SEjE4QDtbc1jMVMHLgbkV+V7qS7qJ5wP
MCW+qcUQ8Jhcjj51miE9rcZktsv2Us9KH9JGeAr0MP/ulKi/lv4q3NJfaAfeaHLO
Vy2gZQhH+ZYYumsk+5wJNhrrYYA6kjFCWm5Amfz2GY+X1dk9eWD17LJ7WOn31jDE
+aD3Gt4USnkruZhKhuwoC/AbTZESdUFDt1anbrTPwDRoGACxOEVATj99pZXlBQnp
XszLUxncUzDetL2F/CP/qCukdZyCWEGYJujNlpN5lMnnlhQeGp6goUjhwH7C/crA
vRVcrTUlxG4ZeHCeOc8FmaQ0z0Nghd1xq/fsyNn5UZJssu4Q+nnQf0ebzZgdQhA4
Fw6YB47YKAia98TncVyznV2lLdJSf0BJDNA5lW1jt/0gR1pOMetcfizK5QWPwNLb
jnhS6JbnAdGMLAyr1xWRZDMmM6v53k615D+ZSRa6VvsPN1apn4U5ynbp0lQ46HKI
v0KC03CwSEeI+WNX73sL0Qj/ED4oVaFWw8i7BConYPPuRjqV8iYqV3+y4lS8559X
3MgDdKsq3ApxzpmLxx35pJlv2ZI1Q5YMQQRGL/LL2xtn/ZrSYdlZVkqbBHZr47tL
Sq3o3p9xY5W/5QK81hO0RuNo3p8TekeZzAyToO7DhiNV0tQ7bqmICPxvoEpRJe1D
vqwWsa9K0bC0Bp2QDsGxQvxsjk5mJIt9f8xmCnEHYKxFHfsbigYxvWiJJy+H4+SU
X9mnl/KpbN6KsKNLSWwne3Act83OqPiUdU4UH8/pRsGsMK7zbolchFD+SB9OvD7I
pomyHE+Q7x6aCZ80mebz6l6On87dYirqmPw0BXaS/q5Mr2JLaffoV4XRrGXTZwo+
M3n4hzjNlmO5saTADz+de1TV87aRSYXqp8BJaXyrrQLhwGVz+SJpPrulLT9r9Wqi
t/jFYbf85g6iY2x8xK0KPi2WP1Oi/IpRa+v9BzwUXzOViXt738r5/70mOQNqMgc3
bj4S2ZTmAWHhhyQO3y5u7s21Coy4jfrNkF1kYSPDEq+9tBMWN6JYGueq80e5Sz97
lKGvb8GhXni84FUdF2rK7jYuGVXqQTORVBlnszQ9vuj5RNcgr1EO+kdKHusoeloo
ZOzeW9gdeX3wigv/U21doxRwgLdVwB+GH/VEmCAdIoGr6DMC/gok1aZMJLQgAbJc
F6MwtfDtyp5+n7vtt8US8+l73ivVS5w9htL0H82CEISP/D2MY42AnSpd3Me42dI4
jZnbQ/RDaJUIuSjzV1KPmhPnsJfYVUEWj3l108zaqnFmkmVDpOQ0akg+YfVBguWH
FRAwLW0/qFYU0L71qwRimD7i/7xC/cgc3zdZt00N8Vi507uRoOUN2UAT7ZvvbcZV
H81z5vLdGK1bdouV1+idQMVDACixmJQKqKFZ2spQ4jCuMDvdtRq0XxKbnQEsJ+uq
GMJZ21e2rfzk6GxIlRNRK2KS3Q+nyt8sMEedlbFugI6CPhu23x3j3xwOOQBRz7eZ
RomkxaEGs1GBRcOTEwdA9z7OUKOMWbSOmNYCB4ob9toCnqOoCfJ8d4Upfp9yvgQW
d5j/HPsGtpmLmDqbQbqE5y1lcLACMKmiJyggA+Nos/utGO0EAODcTN9aKHczMDyc
lKEXyUNDu+Jpy3TQb7WhG5JfSN8v9a//6bnfBL3uvwxg1s2KAjANOKZkXRhDPPLh
wlkY2zVTH3sys1fi6ixdRTYq1SMRap5u28foeJdLiwLITcywZhssXq5mAf1RtLsw
4Fbm2QDR2YRtfZ5rM2JcLZP7+gUzw1Lqk00Mx79qs62SnTrWxKDElixbReYSm9n6
WPYPXY9kSP5OU73/2Ow1vBdLc+lW/jQd2tw5oTzO0emDDziDrnRtvvpzSOBiEOqf
AA2b3f4qJU2T19Ohzm56SdHlXYJ7y0IX4QmL7ntszHPNHsUPB+gADjGwfIBMOXj4
uagxXQ28Rwf7DIiUnbPk46Ea/YNmfRF5pMx98U+LL4wDy2jbmRcq8dgaT/tY5jJw
cFaZXdLNr8Z65dX0H6C0jeaJawvGNyu9MXdfWQytEFbrcgHC+Sy+aM+CsrM/SHiG
8Um+alw7NeVsFIZfGLMhUEkjXIotIzLoCvkyskYTajzaJCLuIMH0ixmycBosYD7q
NodCgu12P+cz7jEzYm0o6ZJpGx95khdnqd5Hp8tbP1Om0X3LX27ae4RgMdmPIl14
SZxUiRVGft5UzlUa3ZrN+X7gwhkKgVEjtKNV/rCMbL+7WlA3hUxA12E9alERG2SE
uDV2yrW4CoAjTG4C5tDEmMsGYxAOHmrAFIDDWfU1kqV0+9yKvVqmpKHyPrVFVEGm
CUwaGOXKcSpDo2MtnznzcPwEgj2c0n15ghR7JroqYgXLYIod9KWPSu9DAZvlcI7/
OPjLaISJaiwgcrb0kfaq3hSZFMv1L/uZR8f/lo2Pec7Q/RshKk9IhR7fw0fBNTMk
W3AcAAQbAKMIka+iKZxDay04JYhkgZHyHpXwwx0VhO+V/l5UTqiTcdl3gApQqCh3
rgEwixovdjuJa2Tyi6lWJgRWkbWFf45EvFLxe8ASJ1IJh2IAizC3k4GPWLPs7/fP
33bzgWA2Ju1PRYt6DwSZ5boyzGiu/StaigO2Num1pY3aKCSYQqPO2zc1aU+gOCrU
256hw/0tGwuOvzADXn1R/z1UBuSep48xholgLhayDcerJqKOxUcJQ9U+DqLD9MB3
N/rltVOZjeESSQSP4qfgrrgZPfGJFL+eT/7g4BlhdoHt/vUTTWHb28GXVG/0n9nL
K1aAH+TbRaXhgPdyjQNtfoEEQ0ncKkBfxkPL3fLYQgY3MQ/6smjhGDlbjtwxnWaG
afBuUtD2C0CjhHPUcdRFUnhk78WpOLM1TJhQ3taU8FU2mvkj3aWzSw2yTt4FqwAY
RtEpkBPXh2FFrCmUGReIpZntIf9Ganp1xkQDTFtPZT9z03mc71eFSSW9nLVuUUeK
yGl+TDHbqj/x91rfI80IYabXlSFVyLZlvOTPHH5DAg2vLQKutoiAAD/8Q6y1WXGx
XTJ9jyE279KmjKqCnbPvjQFEofD6YoIDp8CrOFi9/4opK1ZIrzoyEiJehwz4K3vj
oFFP8vn2WwgFSAG+9M5TqGaZrwGAapSQHpk2ZzaS0MOG0EeHVeOXLDbbTk2mjP+t
V3F/ojbMdaeX1ooh417JVm+SIYRFLLu7Rh9NqOo5hkGpT3C4aEgR+hnrZhy1jJp7
fOGluBeu3lNd5sI84rT4HZ5K+mcLEGHQFfdVCHc8gWHJIN8vt5DRWkWMJdbRzdyV
oXgEF/KIWEI2T9sVL2m6hAlQGTYYktuVNxw4NWyULJdd3XRT64Nvx/pfqQfkmmAt
hzkPeQlzHo/6HGfWlEAyA+YOlMrozu6Fotg6Wi7acDvkr432itWAmKElygWHdn4p
a4crpoHRugeiApe6MBuFmqqHD7ayRw3VX6QdKMlPbs0v+I95X3/0Y713fuDnkgkQ
xndNTougBHG03ENqiN2UP/01REx+8sfIzXNn/IQjHTHvmt00knDtKSlvcXmVurKR
4ZrXYvCDXneWX7d9hsH8c4HjwfcZIAnOs2am8Qz/StgvtSYgxnBp+dfb55PIaZHm
6a88SBPohYntp559NNSz3p4uvdNo6lUbehmLj9xxFHhFBN4Ren58jgptZK6zDD/P
SuNCOKXv8evA5Tmja5Xx7zuxLIiLoyuxWI92zRqmVXTD9tkn+/VoTQQqpOfmWtv/
RQyw5jC2rLi+ok+S2GMkHcHBdIMODEzEv6X3lGwng41LNKzz12QGJHYtXm0lGfJr
pyK/FWsjOTcltBtPAN0mvEbjS0TCxXGIWRkwoUHkZP6zD8maVPU/7K+RRA6tqNs9
ZeuyJ2M5IbR6QCgUkAxPDkpn+z/IL9hTUF1tKJxqtw88Ca3kgPfNZDyMFjgS+6bQ
FFCzXhT4KlKV4NK68oc+45K5m8Es4DaPh969uoDw5VWIGMldJmPK/xXyUXkGm6wj
OvQFPbmR0NjFc3jls7oSmSbZmowNJvM8ZeUlbG2yLB5GYu3BbLTJ6o9APz47CaQi
xOg4BcVBbSQFWCHsPmNzf9WrQIWdPlSglR8UTINgMCVJqL0mooBJ0HWdgkEuCFql
eP65woj1Nn50eoEzTTBbQALM0zM/j0Ds1lTmlnKu/qNqIrj0KDoOKwopQJlbcVnH
5peo5r4FLep68nb66t1ygdPj3bQ3MYyFGJKT6ZTCBcJDkvIpBdq4fgmLIlMYifqm
yAbkUPmVjCwmkFzjTt9qyRJgZI9udeLVMlA3oraRgSrHr+H0IQrSP2uZcEJEcuBt
7Ruo8fjuTXpOTsKcaCk1xiHMzJBkec/e6oIiCAMcPl2bC+Iq6DVWW40a868gwQC+
kptEhmZPFyKeEjwL0iPdHrJxP4X91JmGOrE2sUnWwhsicVPQN3JXDaP1fgDgB88H
8b7VOoYJyYloR0n5PZP6m5E0MBIXsmXlvqqtLzvmSGocZ7CBIL4iUw0UXrcAWSkI
fD42mZVeegJ8U8YLqn6sryLRG1n6bHN/mc5xqAwa2DVHgj85vmCF7nb+NK+T+Ls2
PpVAjfhjX6jpCESO7Ro6QpPWC898TC120iPZELPLBGZth1M8dcqaz64mvIrmZQZ1
Df3So5t/zQYS7+ciPg8kX2D5DXfHHiNtW4k7vzSvEKH2TR75AWjimCMOV7kBJCuy
CvUT/txI28ICTfybYFEhKkI4tbhtVUA30uKlLG3LM2nfUbAfBjQU4fB5wlVLJzfl
BFViIkC+GbWDE0HLMsnUKLzG9kNiAeYXeF0RSLDJk1eJN0A3eWxBx/uRBaXRb/2m
7buBEzCBQuRUu1P9OTUgA6ngMj9lyUoBnWU29EnfXo+yn31ZXFo215bzQJB9AaRV
g2MKxqHLAsI/gRBXwfTjA6IO1rD4b/z0cKblr6D3PF5kypE1SSohglppceg4kaY5
oKpv0q43kDC8ufC8RZUXQI/d+Jlygdk7R/XVzVrxH9xU3BxRI8ckhOqUCPFrKGyf
yY2KV5jcy+A4tzFHLUUidYA+HWM6NrtChT33zxM1Ty1d4UOEgniuQ4J75DcF4eEx
cURwOnzbax7kpVmSq30tE25ekAhVqCEzDmDCzWHy9XDr1crvtVa1MkuGiScZB5cA
fXfRpQUJD/uDIq4FRjzmjxL4TvK5n68Obk0KAugO4XmM2Uw4BlRG7vvp7q96fy33
BNLARFvRjueR1owk0MrdfOrhTLwF63MaUHCsZfabh61Ydb2xojD8zk/Ch4S7UgE/
iR/drEQM/u7yNGbvqn9L9ZgerWDNAxMdSspJjwD1ute2bU+jYnjrFTkzgu+DSFIH
CHk5YECKyITMbOTed3RtCbQ/jwPKUDmZ8RAR23R2ggLq12cD5XutBD06CuFMTSca
2b3W8MsUiY7kE80ppSqZTNerDhD5FN4zoNMrYCeWjp5TRHtRolNs3noW64HbwN90
caK5YxRJc0i9rdEsYzGyM9Jx69eE/uj9FmMjsfevYChDsc3qYqOW0//U1Ov8dwoJ
ojQSzr+L+GZiWI8YzD5SMoIWsaK2ypCmCFQZ3xkWmCNfK8HzAwQzqg94bM36ftY2
NdtDUj83ljY38leQ8f9OWXhmqtbilZumePJuIz5dSEPBoKNqf/lW1s/vjYeYZ4S6
xBYzAAwWZKH11oQ/zgXlDCNrdRC5xeqqBSUcLaOuNsJMc17O9kJWc2TFGDgdncdO
YwQ9paj8DM6ie2c/ODlMxJxItktR79Xr9WY4fTKnTdJ8LZmmFG21pmIonCohu7ue
pys3PEXjvqQUKsGaC/vWT2WnQro1EzntiyJjxwCFeU8yI6jrN519fI6f8jTwqxHN
Gl745bbb9CJYC/vez3HtRCohPUpHMV+7CS/XnWMr4Q6u/OZWLjjug0AhVomjsrhz
s3uVlKV9w5Koy7MVVUqR3F0hzLmswuLHH5q+nWaIBFDWkuID+7VSWjCFmrWKeseW
Q/bwlH3l2370ZU/WqLmBcq8Xg2y8NHTIKj4spSnspjv9SD5f+SO8Cew7H1mVUVzL
t744OxUJ/TKJHAOvGy/774cSlPmW7zjpc9b/sSBc6nRFArfnUXC5OsGmJkgqGeB9
foa2Fenpb77ENTJRn20UP1rLyWGqm19m3od39zltw7WUwGGxgZiSrUcIzohg1EZ4
b0jc5b6zvSnXqEdJVw3voS3A5VFBb6HxdljglgVhg/nhnSnuOpiOxa+GQ4268TbZ
NqgU6+NhIsPxlITYEwgWWqia73dwoIvUKJ04Zcqh+msc0z8bAcAKpsOtVWLDJbFq
3MV+V3thq+AViO3GgZakroJw6cD1537IxeVT4HGsFjrdTsyRC/ZKVwdCDhR3oPjd
2Pmcb+ntf/VVnfrPQqjW6ZaRkJLpHJWTXlxD5POrkS1AoX7JD2oJJV+hPnyi80MV
UbwQMcIjT+wEBuy5TNCEEybAzKc17Jf63hKCRzNjsGZWzRB9SJ3b5OgxXrrUUL87
0Bqfbq/lEwhzkUalVLKdcUtrprFK52fC9MbpYMwRTLs+KCxwQ8rYAyUwlz5tgncK
Xoo4FuwH0WY90pY2ijIxzEPv999xEjzNqrmVrbwt7wIKxqcnF277GkGlUtoUen52
igaI1DqFNKpKlV7+WufYmFgYevQXwHRLTxsgVJuPp/kDEWuCdNHMbly1pL4YLY5r
8c+ggoch0vQKZXwyPhzj5f9xj7SgBXz8FVnIrtpcqocAk1z5+H1cofBCZ+yHqhJ2
z4HYUy3/TQvIDZ/MxLOnTsYgW73hvQgLt+2XT0a4mKKZ//h/c0lG+6eobzlB7jrb
9Gr5s3P9wytEc4bLm/09pagUTnaz0qBBISj5LWHTTy4x2zpWbtZzGdWpKIZPRJlz
hkhziD/PDWDJBuI8jtWISJ4QGrCjcrlA/G1PKkTMgJfgR3CLmqacVHIq3DOKfqvj
XOgGAwAvX37ya8N4AXQ1A5A7zvgviQDuCLL5Em6bCd6tRyqFaj3R93vr2SRoICFX
CwrL1TasrTY9j+QXFl247o2HHf+KYN8tSGnHBH6CLOPQQyIaFRbBjSS0D/RhmNuf
H+9UXw62vTmBryrgw2crCmGjQNy9GZ92G7BJp4LZcWXxI3TU2YIjXBElYI/pVlsT
709G0X1UXJq/+SmBtVP/vtFO9cBFjra/jv/dpJS+LUWbzfEYVNq10ush+MMWh2mA
xxfaWGzvNaHMBmuMSY+lM9+gAvTUrQW4WY33HlFbppKJBQx6ngrK/Nj9K+gGO3hM
4cnMeOUkX8eOqlGWLrbf7NphLtOBxnwkCxb+Tx2epDicfVomPd9PvZvlmv1z5yN9
GnfBvt71Jn0Qb1i8J5ILazZHZRxPHvUzvaK2Ao7tMNri1TAPd2r5KR/M9evWXvMO
/PH7ZDAVKbawGbPjSxBzk7SQZyDK4TSu6iEEfKA+9dmfV/88VCQhRk+pdR7+j9tD
Kp94GhjO26NI1hQBAf96zvmuJyH041e9cPw7FdyeBh7Ia+P/2+H5hf4ekcAs5FNU
AXHh30CG9Wfm73ZZ94AQhhaIU2H73Q0q7kynVBR/zp4h4Ll4bvDlxp2NaOueiH4m
ZsL7F8izmtXTaZ2dfVavOtcDHHGT4bOYvr3KXBGDj3h1mtXZGYjPj8bZwwVK3mHI
JU9IomUvbM9lBBb8aKEksdW9XH3MEOi3DScpFKoRCDhYZ+Zlvck8KfM1JktKMtiV
fBs8m0F9SLfJqSkZcpCtnNJUoLKVW5ortnmXS/bteaWvEXFl3/BoXhkxeAU71WlK
tnkwsUOgaulyzMg/sYjmS9Cw4mZtGSwbgyTtscLlW8krOm2maDGVmKa49zYgu3kL
wSIcZTpm9J96HfIUtyt2JJ7LsXknap7tVXQyrjPMKys//wiRVpAbRmLj3KFI0mDm
tWYB2DWegUdqRvN9JTPMHJMUYVbFguh9nux7fiAk/vIpdhHq5FJU/M3aLHA00k2l
2Niugku1C43NxE8HOJUPsaCnsvkwiRzK2jfUOayozeG3eRyY5YCVm4HE+3YSJwQh
NmpQSIliSvwt8kPsyRETl0ahPDf9Dk2arFmGmuQRXfN71oDXRWxtWp5tgD5UlAtr
mFNWrh0KFHy42/89EbnU4U20bS2Dvv8wbRZ6PqKs4cKAEQj1eP05LCGL8tIiWd+r
BzYeiEOnypywBLWTpdTmMV91a8vLOzukHSku6Un7jpawpSIBw7ILVJzE4xj71dBW
LMzLxVDQVlk/r4ThLSdtCFn+KmsZKZKFbh705guch0+EwzaWINF4U5Y7zaw5EOoa
ZIBD2zfuLxklqMD4gvFXfUD/99Ae/QwY+0DTSQZIQeMVDPJSunC76m2xq2lzL7Lh
+TpajoA0hm7OKvuxGMTxFnOpitjVezCj2YIjCugW65dQJdzSBH7jVyNX73Lur5A0
DjTyhKWmcuyxj8d7LduZO971fJTnXkTYJu7NRivQHMKmHPc14mIlvJJ6hf17pqWA
Z0qB8AqavIwZw4JP+zJIWDKDzZ4S/U/G2rs/xYMcgd4bQBGAO+1JSwzm7ImBVcyC
Mh52XPWKJ6mRXHruOuT+Sak2dCQUMWyxMoxyg6GYqUJOiiY+3bo+Z0z8WOWYXzu5
pKWAADmTs39FBSmSeLLtEPTDYVYlNCw5RS4MCnT/MPZSzr7UmOiigUC98TK/2qxu
JvL3u7Ga3Y+5ygf8hN0WTUTSvzv+ZcLWpdLkYk69fRKkVYtbSC4k/UOY4ctQtHyI
Z3g4V+EmXMvJXhdgyJMm0/8eRY7n5+re+aGWNcprSHqHSmivGnDcmdgpKtAn8RVu
sKTi4KdKWKGLalYV9Qny36OZnN8jmHVL6uuh3coU7vjwtBWyFY9zU31mtXghgoZK
taB2RSkKqnKPcVyZXtVYOWy9eoUfgIsb7fEqh1pSFZc0BCBffcmJ5Z1gvVysWBf+
adrvfFdVKO4xxiez0g+pk3kU6BBnhTgVXKVtQBQNDvt5/iivM978qsDFSYzf4t35
9DJ3telCShJp+ZVgIPUIriilvj40CaOmIU2NPU6XumoApt89s+6A6aomxaSt+P2G
z3Q+SdxbXDYhjs4VV0Xq+9NufLmKXe2N7qUy9AVkyTHJN0ktBRa+PChy0aRljXYJ
RJZMQCoEGrRqbcTeSYlfCye46XwrUGB8sr+5YOg6ZAjgsNQ320DG4azBFwm4LPKB
XP8E+EP3xmBO+cNRSX/3gGM7XqTMjrbwsFOoFaug9rQbIKnH16Xhn704Dk4ds0rX
5ANBfXvG0Isl9m0m/OYeqtDer7bR17L2UFLfhf2YrQvBTmxXmalu2C+xJ6hnI3EO
MNXVkpsBw5jSy4vIohLZILe9ajPYilnwNwciO4phn+zDZShV7OFylUCMZ70k5LXE
bG7N61+bOfSiC/ZoJE72/Gb7gQeA19nTar6ev6F2/10jaV0IlrAUlG7NQPmvLY+P
Swv8Qts+Yq7HrgWCJUECI6sgylooDuylMEhaksslq7ry9Jmi2aNaZYSmbnZkDlWT
hbueDa4JsZSq4MlnXmsEKVBjxPPuohwQ6JBDJi8UzM4/xTPrIS/9yvor12751OIu
b57nFSgbZTLtIAFTAbyZP9PqdaQr0iydIyKYnsDAhqc3ngyLiQqux/9IBKn1x4KN
gymzsVkBVE/L9VyAtzYKa7QY3JyqHZsJkVCn3muPZBT/MsQ5+hfXvWVeD2d9jAlV
gHnDboy+iaMmufrAP/hFYmyVkavHyIFJ2kjEpyg1y20SYNjU9/16vROuPpnK8Rld
IACvSCNQ8INaQpSnKstVwgOXS/IYugzDn5tDLZvMHybxBmJyOCSq+QV2kZDRg9yF
EchsxtXnxL8cFtTx1NB5Tniu5ZNmhXEhOndqdPuW9BLU70IEm9Iq3XwiO2ffMdZB
IaYGfx8BlD+Agb85AFGxO6FfTgHjFZw4eINEe8XQybQtkfqsnfbNYGoTgAq1bkXs
8NOTSOswhQdOZmuzdkxLvHngaGqlynq7SuT7vh7NliViXI89V+WC5k4yhmHQlzHM
y2LlLi32+b5YlBWBwQqW1U/iZmcSebzdEbixH5jxtJTo6eLBHm0ELGhCqqLNcshu
ipmlp++yuR2pQyIUn0nUZWfokyHzIhCAmMFv2YOeL3JhT6SR2YyZ/TLC4JG1wkDt
RBq0vA7ePqP1gy05ESLdnkPJ6tvTsGXiwNbmJc+FTtYAXV/QxJQvfbc0Tcoisfam
JpKi3haTIcBWJ5fL/esGIFZeEPmN91JJWNZ96uBFbaFdD8/6TVb10KX0pu5/rrD4
a4X8f55Y459Qqm5+tHJgr/c8A4pb7tT97tesya5CpEiAIXW254o/fre0V2510WSt
2cnsrvNBsnsShv/yhuC2poWv5mi4AMEOSgM/+XLAmj0MNkJ6sNl0oWJvcXEra8w2
I++2E9qE3wHS1IQqG5tbctyTKPTCBCYWP4+bZT1m0AQiahhXOzhpxtTIwX88qdq+
nw8f6BdYByL0Qn6Gqh4jVDXseUOwjRgivNnHRKtfRhLQJcCwNVw1fDpEy2yfgrcM
PSwDafq75Y6YmcC8P2ZHYHEbnGyyYysLNZwFNv+vXYdG1pYV81eaVSvko11gN2YX
SUtD6y6xn2rlJyObt+W+ubva2pdXAwyL1EswTt7rYVzXKgElRm7KVGC0smZRKwZz
Ff3mnZQYlVoqKnOdMrUw1V0CaoV0tLn+SHNedyJTRdRc4ijx8Kt2tSou68rcbYAV
uIgEvEBTKfzEbhoaI7ReLYySRi88AzEbXIYElh3K3/QyrKVi7+zJ7+LrcdUMasTD
8h/XGLiKSPVTb2YSRZVcGkE3twOHNRi1IZof3CgHMZbQF7cAYSpzvFQdl5i0B5Zh
CuzZ9v39THjpT77LHATZwDFzK2muaYIsXEWPUNMJT4iycVcMAXsOk1uH0MwtD0rA
jHBa1H9rYyLRE/qunFhzfisrEDJmn9mf/lsdo1MHoh/FeeXtR9ZZ7dXk7asJYcKf
H8AtVDQYDFAqy7m9onsB3/BSbwW8Le4FNkD8g4mMI/znjnIqDqMRik2oqYpWnQEv
qV429nIMSxDPNfiP2uZD7roZn1UWHpknkV3ArPT1YeKBl1/i7qsZvW0CSY2TWgQ5
duqZtzDxJtwv/hBLBjF4e5ancT/iK7LlDcfdv+DzkcQntA6lGJLSXsG6vPptR+6y
tXQUW2vrce8uNXHYsLZRjaXdP9MD84XFEah+RUAMV3l2mR5P/KXVmO5HryrWFauz
7K1pW3sQ5fD1l1PA9aE/aZKaTrdFIySGzgVpB/fHrAmryPsgAfLPukEt1zoFs9Ao
9b5oUjBdW3+C6EmCr/Dhw43NGAVejVnyAaYiIHFrAU7gSeGklWFr1BtmtKp61teU
ni9o3nNm+5o/JviNINRLmXcWPufhXQ/ESV6qZ9b0Kis85/oHlQzm0vRttEBmft3r
PF2sDQglWgwsOoFL0t0Prc4rk56hJfb6PRd7mYfx6Ay5bI/xd8//8SmSw9f2C72M
ZbvIV9GbidsfaTWcrQn9USVh1j1rgyjESFN+By+7VL2cWjcadf3cG4iPyodfbQYJ
5ZdjwLK/4g+aefDwQEu4nKH7fZe4mD+Q/UDUb6f0Lc0UTLm4qj+8ehwKv1gqQb6m
RL6RefbZCeJj8wokqRXgd3dhEkD4KVXDb0vIFxqBxXdTIQlA1M58qarHoXLIRXkj
rbtB3R4mJZcniVlKxnn2Du77ErtvOGI0YdtOh2xLOdh3Jw2OMop7KAProS1Pd04/
iml949nZzoxEqd+kgohfEwqgj2exyw6Oc6ju7oAB4twsPGqETaSpt/m2dL5KwwMB
TGwj1dHW7S5zDbEOYGvciQ6lBd1VCi//MyruLZU1D9wu7iYQaqKeKRvptCNUDebh
yW8toLLPdHWt0UyTTPx2Yh3jGOf8z4BzxdBBtP8nQrNFuhr1/ky5GFBXpM47fp0l
ZofVHV71SIfrifAoXUNJSm0WM5cYFTW1C0m9vkbgLGpksQLb51bLGUPN00CV+NlD
ia2PKcMUFrFSXqDdeFA2JF2NyJsF5TSRyK/BcrwRBpXp6O1nopt9YjLcb83MPzl2
z1+IGJX97zIqvOzj6qZzHNr3+d7+RvF1V//2DhRor3dBH6lWv6bpYUhrDgk73bPu
t7aMWzzqKqkaPXmdfJlwcZgm68mio+UiWeOUn1J4hcS7Z6D11kORP3Qa58lUJI2U
bf+1xT71enU1YCQM0AnUKKfHmTXqu43YhInSuRYouK6zolxqWU53Ak7TWgOxL5VE
G3NdCL/DCyCT3nuKZTn6h9AXD08u/Ni1MxV6rAVzICTzpBjWyerKvOMrHOuHYwCA
18cXgkOGnGCcmgf42+uV757nIV8BZ06b7Un0H16pd/oeHgI1FVaYNY1fwHQ1FIW7
MrpElyXhC0DNe3h5MNOf5ns3H8kmjQtDAEf49deBItBnTjQcPfDSqLTBUC43lZJG
YnfiViZSD1Mim2kq2v3pOr0kNXQL6hx/zWaEcJyeKJhiQ0z3lXlq7XBpBOLPx4TO
qAtHU8XrZ6NiyYEO4bryvVRtq49MLaQAriCUUuBgpkpap23cXTR2Mau+/rRYPD6e
srFISOSgEq5egTrGuiC34SeUjOmJE6FA+TKnRngGn7VUky2lxBYiES589sguhX/M
IGEe0YbH4sXZDCzv2EGTXrYTrQJfsNRJ5M9huYqRU6rbb+TnsexjUU/2jR7KLCJ+
n1mfUxgIvDPhPd1kksSZM497te6jfBn3uDd/0ATeETnRUeD+GTV8eQ/oyat405rk
t7hGVuxsiikWVH01kz897MVyARDFQ2pJDfNoCpwzNEkH9S/OqQbwKDqA/2nxVCj+
rHczcWyZG+HDQ72XvjYQ+KpE5zKSp/pi2al652b8Nrk2UPCfcy4rHB0nCS9qGqWB
vADzTsUTHq1hDZggkOb9pICI0WKERiUx9SzJqfEOT5oVcdotDBtoj/cfn7H2MIZ+
tlJTgUOqZSRNJ4Ir3a8OXCNvMjWIqzCWd96x/c+rlbeW/TE+WrGhZcqBDZaiZgVG
cDIk/cCSJTa9o1x0NZUSjXYwDYT5ln1wCsn8mIvLN7hpFeBdf3vtYflyHU7FtW2S
xGD6gAYoVFWyA4QOd88vAueIV7JWmFjkTVtjv/Bi/U9mPXkqR2jyLxxTxzIL0UGw
m2A1QNsvjboZntuAWa8sxGHV+1olPS01KZQAvcaiW5uj5sLXV1EelySlbpSeaNlF
zVX32k6vfSWds9RO/QgPrkzTjzo+bloDe5NHmp3T1VGUokKL0ygFn5bkaAmkNwk3
JyxXekdaKrqW1tDAQDHmY0rugetdyqehrYtIsRb+K5+QVusfEXinFIu0vGiItgqn
HkH0RRw4q6nJf/ffxAk1qFMfeQxPfYaZAbNjL5O3YmQBiazJoakIFyV3tStZF5ib
HMSX6WsMwGiqSw9KihF3xzt2xNafRXEy7rcua4BLV3/OdiRHIHy7B8daNGFl7Lh3
PeXf3q8bh2VuQL0opY/YULfx8eqJxIYVd0X6TkW7VCHdvxCNkvwCKiB0iNSrRyFV
Pk79+YDU06GsJJWcOwANEu0otpKZxFqvDe6ymHF3JZievv7/IZJm9z+PCJvj2QtE
pTy6Vx4s1xOE0yzgWDchBqgtNZcjBtYSuly9YvhjW1GyerDQsCQRWdOOtXWM/XgC
2oWnutf+H1aGne5kV3UZDrx0Ehi6zQviP8L2XU7Fyi/Re6iquVKJXdfc3UIqnzdt
XZeq/JqdHenAhtnATTKXGWh+qaaTUOkxjg1q+uwB/21/kGdBbXPi0v7Etqpi3Xur
kjG6EpomzY49G/L1oBCj25PxEGRU9eMZmb7NCB3NT4AjDVQp2G00X9GEphQU/t0V
+KW3HtVz/h+d6/OqBlWeSZCidNITWJQLslcFWMpqCbGXLNWat6mgZcp1+7S61jiN
9KFe+6H3ChobvhaIPkDi1bd88Bk8xIvEiPSTKc9Dv8262k/iOFoOw4fu25U+7LdN
UNYKSGUPHQFZoqsbkaHiJLZ19XxY8jYUQ3Z+uW1Pcmiun6twrCByDd7A8UN7KwNb
R136ycLRWyNHj2bYjMeflpTEuB7jSTGjVvChAd/+d1A34ucPq3wwmQZy2XMVWLGk
+ZxupkLJS4e14KI/phYbJg7Z/UZfoBz+/hLgPhKtvxPhFUUCwwzHMB2zKqKJft/R
aIeHcU8HYIEl8jP//sncFUUNf8tEbZP3r0Kt7RZNIw6bpjKvHvxJUuoIh3I48aVZ
nhUsSXmskYUCmKYORG77zgV5N2F3SFpXhF5gu8HjQBOx+ElCOFBvgWtluS1zyUEy
0cr5e8zEmFVt1s7ymNnSYw2BUzjSsGbtbbB07EyfFZ8IQ9Cip5OwLqCXESYlWypm
Q2SP89m2dHF41v4z63yxjKVzGeLqctTZk8/179vPBtv+sIw8L3g/TgfGTYyGw0gM
pPa0WEbS/ZOEMd4w4WTxsUtejaTqddj+aPSVuSc+JDbATMMrgoYDnlNAp1I7qtBD
wIKpUZVtXm/6z+BukSoqToTzf/syeuzT4nhCilxyuq8hE+dQL8PsMfRDd2N/6GoE
uJ0zyq7fUJITkHZBNHn8JxePPDNwsgN5OlvOq4Mfq12swbtwzkRjicBuMBRPuDbh
i08fCMWyHEYN3sB9w5ZtwPlfF1CdoJbRK85eIbvn3bS3uw/Mrm9mInG4GveTlEIe
PAslMi4WIgPaH7iN9bJxINdnnliqR8sosCKr8lIHdWHOvgK3AY6MHU6G+9O0Huo4
fJbKE8knmblwGCA62E4AVgHwJVx0b/EFpG6tC8fh7FvEkj2FvYtelQFRLTa5qW6/
7DbGa6e7mo+F3H0O8YWfbTjfQ4HZ/h6LdJNcuhYzcImHHnGZu1fRCvJhuv1yG29O
yYTbHSUWBYkRUP8v7qxVtjRbpBy0LYo3AkwWkuaY2N7BzjkEELryGzpZr9sUD64B
HBitKw2Ch0fdIM6/dT8ybsFbTTnZBtppvrzoXq+ob5TtIlCtAhkCP38m/3wVV4z6
wy7NmbYDvDCAcxMCZhU+y277vEs/O0SqduiotJwV5bt9MCM90toon46G1McUEYoO
lDIN9oklQaXGEzz3/O2KPie+XfJrcGfeUrvji4uGEp7gNwvrjCdOfhfhpJKeTmKY
tXK465zBKK7DAnMCwIdBq+hJNflQ/mwUkqEkK4CyQWOoX8YGLBDPQrXkUFbTyX3e
fziX7dv9OJ7Hpxw52rXvxoxGhcBYXZUKP7UeqVBz+reG1cM1Q256T1Q5XXnMkeEk
5yYiwzakWVW2rEj0MEp9IDvg3+XnVOt4n7xOehCFKHxWqT8/vBiDw+mJdNbPG6mi
Wql7fCNiPoBr79M3e9ZNSsncs3NqqrisemkTWdeH2b2R9p/Opc7IDkysgLRJJ1R1
gB8orV0jCmc5F9mkiOice0+FYFUdwcBk/OPtUqL1TvnjGe+BL2XS4ZRKD14AD8mb
sh7y3Gx235NGkJ1vOD2zvBc4PKnZPoV3TZ5lh0UnSXqxrIct6JlEcv0LBv370yyJ
YPLjaZnTEtKDi9GG0gea2cCJ52h2Musc/MRtaxL+OYaRWFsRiq1oyqhGSf0wW/No
yBUgj2Xjg7UgWtezr7iIIAfds2JEwRN++OffQJk7MPXIsK63kvCBjGRYIrVw/rjk
ttF67ToI48AXmxebZ3fgoM398EdV8T82HchUL53GdznupglP4EMIHqRRpfg4b1W0
Wqn5RifnE4HTjZ0OiBFMgfDm/yvWN+DDffg7rhOLI26PAex9InubLve026Wbwt5t
hcl42KEXfKXJ9Y/4P4RxPCRTBH4nMz6Ub8h0XrQ7gf3cYJezDoYhGy4mJ8qN/3p5
qDckG4S1fXJFg4IGmWLYUmxwIACRJqN/mK3HYV3qzadNZLQUJgZullfuwgyOdWsU
ATO8c2oSaSx/7aFtB4ET+7AKBhZ6C21X9nxgOMJ1ZzPo3U1gvPQOATDf4azQl6Ch
lkyGsGmIn6/o/LJLuqCmpPsbc9yRyeCta8yzFgmUSgZ0BLEcp7g10/vtp6DI8yK4
kW0i/SZVDVyaKmFjv+nIMesLNtahf7lckFzK1iXNGn5EbqJS2kLdEAnbS+h6OZYD
b0Nj/HHRXVgBaXjN3y+I4f9eHEHOCW+ZPjR2tvjC9yGzOjOEV5fNPXjUG67/lRZD
POrr6Dzi9HtUVvS8Xa9yQfct8JG8dgBjay8JrMCurSWCcwYKes1m/cY2FtrE4JlK
ID27esVQPON0ZNOiGf+h/wweqy5IQP8TwCcuzOe577QM9P8R3zb98xOTXY55QuP3
Vlz4Wu/D6V8JranYjyuKGUb5bRWN8b/+S1roVVde0iebffWE+qLStgolRa7gnG5X
O+K6FH3Q6HkEWD0i6vbqy/lUdh3xn0oVDPQtzhkI3jlExcsCXRz1Xj7kRqf3K0XR
8rFUkKjmILtKYUDvZAno3yWjLM7wEiuJEbXOLfEMbbbrsNHCMyCuBdhQjBMi1xKS
3JDRbl0uIVcfoHf0TgSEOSOPXQBig4hrGPU2zpmKr6eXjaicBR+rYg8tJBdEbpgc
vlAQtbEKQmBrSGZ1qRzl9zK3sKrL5oyrOupwfV8GgtYJi6djxxdamvFCU0sXHHOQ
R07zYjV5HwSQ290v/cI8siZqc0vDzlOnGfG2GvdzxKlqrS8JgBqOmIGifaZoz55k
fODlIWsKF5zxBZZc4o+takmvzVeuNhBCGziIkd8RPLEV2VOXbA/h6+6hDl/e85jp
AfQI3MoT2xi1mezrnqpVejq/dkqOEAj9l8z71XeLh4vu6TyWWyrhORf+5gkYxkjI
Tx0XL1k1pKaD9PEr5eUGlnBfQzHhEz2YFZQFRXtBxOl7q8FcvOpaHY+YsUQhXj6F
s3OXLxRioJcbeNVK8/TdeJEOMRUjHgXMxI0CE1iLm4QD1/gEEW8F3vFYdISgR8Y1
ki91KO4gkaubzGkuvrGo0cO304qwca2EEXGl7SRM45wDvducp8v2+fXbPD3VEjps
JlxJpShuNoacUxLt3UYUuuUkULeyuhZp8ODsP9u281UMX+XPH6O+TpI0xVCMeCHk
5YfEt407Y6n7vMjuE0bmtepD/ZOB8Y/lsgUI/fmqOsuE9xTAuOR0UrMiOpBzCGl/
+sPaXM6sNaRzz5ufF1Ov2yJM/n2id0XYsVcdNPjq1KjDwM5cgqhC+Q4cfdQIBV9/
631wNzTA8uYHrJR5vIdiJqlJL8DgNbR4RlOJ4fC4Qa/cdbPYynA+2xQ8RdRfWF0Y
jy4EqmJARofGlmjB9IKwZkP4EfywOGvGRbFZlSn2v/If9W1/LKB05LPB62P+UGvZ
Nrk2KeICa50+ZwIU3gzrvNdNVlxSGvSc23v4YlcDQEgBl+z3ytlzD8W/IKUr/f92
4M6Z+elOVH1115DiORHHG+sl2e4KxG3Ec2Y+5c0uJ3C9nLSGAK2TBO5g18JK+HkQ
J7R7qaPq83aaCOAxbP+YA+tiOVie5YO21aOVY2EK2p6OUWoBvoL3Gf1nWTRY3PB+
25s1jDh5DewSsA5oK00t2jw5lHyovFRBzooslHlqlxuUkBuX1UCeS8E5pYb2P0bz
gtC1iWuVazeHY1RJNZzJyk6E4Q6ZulvgtpsKpViFIy8XqJj/k8TUZP7cltyzLoQu
qrAeA2AO2Uy5xTS/gikQFCMFv6GEV5bgB8K3fXnolZxmOHVodV1yeaIdJD+xYcAd
QkGzWJICNJps7hp03dsaIJLDRoXoGbq1jyYpA7qwjKoGwJQlfMd2A1ziEWIEh6UZ
lnEr6s8dltTHm1Y35Eup2q+k1i1y91fpO6ON+VH9GjQGUhGH8n8i+WtZC1OlHTQX
m2GDpzK5/cQAZVN6VO3P6Sxc7R4DWQMbp030LUZuiVvflbZWUqqUdCRC9H761S6l
in6qWdYX36pgDNz+O1PhpBOfBh+Rachoqu/EA9CcmhelvDf0rrMwZwmZ+SIM/RVK
qy+Pw8Yxj4gB2oo9dR92fh13QMnTwhLGUFK2CoW5xUXEHI2G97lErMy+LxZCML07
4Hw7varwDpD5rCcgFWmFzezkJuQoxJzxuHuMJuJh8yIf/R0Y0znlueWKAk96lLnS
z/csnHxy5Q3G+sPyHWFjs6lzXl4ACA3dAnvswqS15y2qv7WNoNw0cHACSmIWZf1u
n6cj7DY+QsWiUrN9ogL0Lzfs8uMFzZd9NJU893pvnoowvnqxDcTga98Hu+0gqCyl
Oj8QFcnrZ28t0QcKcYmJdoMokfI8XIztyNBrNHKoWX0KeTa8Qu6ZDsSjtrK1f98p
Bzk3e5lPEqqaXzTtWUMua3kYF91v075piWvDndHom3RBtDyt/0GwXGx8p+iNBn//
8B4prBSzI/MIBz3WethZ5b5fWJXzlqB3BbdFeEi70c52XXn6VY7rbVl570mKgtZd
Ia1B3LcZODX6hG8hrUAtL4gTrqCxALrJevJ0IaCScBQPUst9Z79fuIkyMgC4YgjP
kwErxlbtcWghoyYSOZR3rkGsXz+k2N6wOeX4Bf1t2lDu5qD25AxvlQkOksQWSR7W
u/iTsH6lfCB6Tx6SvEO7N3AJaA+3e3YzdZzHutdXogabLMjpnE5iCZld4p88tdO7
qVPmpaUSvD7MsRi+ANwM+eCHoSFDElN99uP0PfnJZn165YKzZilJeqGMEAkNAl4c
7J/s1HN3pM7UXj2Uhp8yc/8pHtoGs+96+aXYGIePOwm9LL2y52rIeKMkPWHSWBx2
xWiL9Zqs5HjFPGcJndRYuEPn6NKBBWlcPw6iKRLgiaaqo5uWYbU1DTgANU5D0nMh
N9pbhwB8DI3gDB8n29M8DIi6OgF+dIKvvIz3ZVa9/PckHm6vR5okFp50uXd3Xksq
yyBh5A8V5yOZWi97/xnVpftfrPEvV6+GJIFspL8S7XubOBz4NN6N5A/sZX9bXmw9
nmDNzKAFx+lA863OODPLjjMuboh8O6r6NEFGGE5jvl//sovMfoeYEDldnuXsf9SI
FvBfAKuE0MyR4kf0ykKf5wQD9BjGph2AfPworxPg3zmzmreNYGk24vk37GI4DQjk
YdflEHgeScB6+8ykIXJOsV7RiaXapza5ugvYmMyHWreVXAqQbFC8eNT5UFwtvbkC
VpHBrJFzAh42YKhAEbYdtNE9/ec/fxYaO2t76aH/4rW4X08GvZObiTRvBbEgPB6M
qde6GM4FRei5ZJ4DZ3SeG9PI4iAb4DC3ll6j5b3emrSk39yP+CMxw3lj+D1cc/3Z
OoSzvIg9fWkaFqmqshSMxhjcV9j+kX/NMOXW/ElkqED0Cxg8Q4jSmC6YVX+8t3fn
UBHMtVOjE0X2wUYwf0V9rXrDlZyCXZN8cPl2J0itzAzjqhyN0lxYtVohNXj/sLDl
SJxuhZ07k2KrRzKimgu8+MYnMJIw5gEChJtJjstCnSAW9yTROV6CRZM/1/Me0XKc
/9SATjFLKzU6JtDkKVIeesnFrauqZOAccZyqy1wi/xsfXI7xs3vvMdNhuF6AKeyK
pix53A0M3q0ILB4ZI8sAm0DHC5fDfvwf9M9RRBuszSJUanIUIgML9HClH55TsK4A
7iGJ+AFyBKrAApPb7DTc+PRbGVzHyxwWeh5IGpJVjWNSvygxQnBOWSkj6RTfTMUz
0+RfKKGP4PC4rwVJ9anLWvFpK7VOZVsriU3muBJKg/OLrPP94I8mwAoUPXg6lsCq
uNUwEvcpKP65z5dsxrTXruhuQ/tKyx0Cv8HkCqTVs9oD6ZabOQtBEciN4PnRV76Q
CZKmSt3PXpNdiZvfWXMjs+OG+7SVUAj4vZk72B8XpEgkyAQvPX7U83HsA3V9WbI/
Iycgbq0ofcw+05HaHawoHz+FoIqjvFvzCA02Iop2WakptMqs+MifhnTll9fU1zo3
b2cPWQj0mQQRmNmAd9ZCVmhZjs0IHXmL/DkcQuEfoWDhiu33HwzObzivASwrstJi
sHNCa+bKSw1iUycz3jMnUzEBm5XFOVTU1Ptq6/FfQSNFBroMrnJE7T9eAnwaZLhh
BDcK6FpR8IxI5wglm/JDuyhpB5dWZ1gos1rPTpchX6BQgmCVuKLZH1564trpYGRD
4NSdSKcwz8qlkWn/mwOLB4UoCWJW2EVE5JFeFAe2k01IsAXo89uurC7hZ+Q3BVZl
O3bvte5JrSaidwTswGhkadJ08rbNF3C1SDLIbMvjXT8t8JNrI2sKOPsGMiP9ogk6
bhxJ1Jxl17UOEhOfSJcCC08x0YWj1EjqumCpSezi5bfbGi1cwTalMNFOnrophHlV
yfhTQmrq7XFollIN4ZcZ403+M2SxRcaH2wY6cTF0F7H2DuteKkVobBi70eERwWNf
I8KDdFRVx8CHopTEi9yzTehiNjvD6ep911VsRm/yL4QfdLukffEZDQmlezLdy3ec
V0hyAr+2IJbw0MCQfF/RI6gR0CMebz9AJn52CuEDBcJ2Bv15CJdjZkQrgSvSzzLA
NN6Pn7Qv8+GAtnCfc0EfBJR/HLlSyang8k7/e2gismLRDE1AEDSO/5FQa64HxEMr
NOhkFZRmjL9g6QL6HYxYZsxf4g3qZLnaIXEhP5ulcPhJxslyJlU1WftUHLavWH+d
U985FmQRyidvf0lax5hrh9AdpERZazPNbSpJ+jMznYpDU8K2vb+THJJAggsDG+ny
SiJdEB8vt6NzcRgwD4+L0dTRlBLlCTKdJN++03erK9rdxLdboQ6ROCEFr4W2t/Xy
6QFtFx1EaHq6ze6UntvIzbwCE7R3qnP0hf06SvYzDWOdx9q7MEt274itKFiWM3P/
iYSvO96sBGI7jK5PgGqooCCQZDW7d/bAEZzN0BKPVMs2c146zuxU+tieQk4Z0SWR
XQNm4ivdKkw+Zm9JKv9LSBPVSTwkWf9wOVPXdBuNraO+OtXoSaxeRkyNAvgE3HQ7
MsfGOHLVi7tqLWcIaZM20l99gKEiZqCzUqSE5zKsoH96+aR03F+qpZW0p30oAvsM
u8oWex6A6EPjN12sb9bR4ExEVf22lEBURoqNQF/4Wj4p/mw4ibNtcUuZMHsvMVXp
7nTvmgt3WaWKP5jbdOhVSide4heFp/zy9Q3r1xFO0uXlCrD1RBBV55FOorD1VmQN
SV98yli1UMfRfzDOrcjavNOuEGRyz8LeY2zUL10gAFgo3z3uVOndMQ7Ht2K3V2VE
n0zrARqC4t4paH8MuZWmqwYmX636d2z7RYsdBB8kOuKvQr7+v1pXrsUZGGfoXAFp
ASnKQOBq4ND7EeSkwDI8Qhg41R04i5i6Dks9zLjK/VqXtq60rz334JXbVcmVsWRe
/jYGl7vhQ4xvyQ/ip7fMrsXcMeQu3uUZ/CndHjJVwhgPKvl/68Zi3FhEoYhsDi+v
9edse9Nfho3yNg/B0YxQyeEp+o+05IbfVSTvo3A86YcK/veHGoah4Nqih7QzPSvi
os1axGgnX95axVRsC0EUxhL3pdHyVSmQ12cpMdDYee0FaBmL33h7QABhUr4+ZJHO
q3PuLNMO6z6N9uwGz7xBtf04Q1i4LOrF7KqNCQiNDHpQXz+yni5Tq2VaqXtY9JEd
cTrQ1WEKItisPPenNk1GkpEFdVNiOL2tNryM9Z0XcGDE3CL8Vl0kkomjqFBjZGtV
KPD8mahs5Wm9rWz43Tcfj18+HexRHbYU4ncke68diBceEs97zXHAIv3tW+X8CG2B
jbEHlUI0goojJlXmB9DIZpTx58i8WJQRJZBzuYH1unkwdSrqXyL919njlVcsQutV
tcYrHa00RDcOydwUwpnk63tHY52+imj0UXyg1vIJTY5a36kuxTW7H0A6pJJd0lJV
4FFJf9p8YavYJJhAoemU3e0cy7ILsvcKQorJd0tNAUHdBBQeK84QMulEE//6EKbO
QPY6soRiwQiGeFeNokawIv8MJNz15iJwBzpMmIlOTe4nMjFXGHxvXOfzn4/r+66w
SdHOGvjzcAA6DML4qHNLeMHfiKbst726dk6Iux4PlmX9sQNhoC2+0wPpHfkoc8T3
Z3wUqEzJZ9ICXRtFBV5kSdVjVpOaSBTU9dyq1LrqT6oC3gI3j3ND3pKtbYStmK/2
rAYGcY3a6lQPTvar4rtlG2isEKc0Wmel+rv51ROvV3x78uRzklVESr3onEeE3efX
UOHIvRp2vo79kPsfb4ljDkpFmEC5UgoNbfM5LoKLzDJfFcs7Baz2kQQBgG8vBFIU
uWJ3tU2m+NH5Mo5cHbyePJaPX6BdTgDU/gZZ2UOx3kC2Km0wnJ5EP0kkZluRd+HV
vIJtSkf27TSaFfKMPN9G9hUu8atQ2f3YGP0iG1XEGrh0wqVazREubTG2pDiGYVFU
2mZmbX39voy5/x3ndDzcRE3DUil7nV6ajNgzq7+a2LwUce6SFGSrYYRSbBGSKN4w
JDcY9e8MC8vOXcRL9UIIZofhDJSpZ7FqRX14kKvfQ/9Vwcfy+YD0mTC7P0ouvzqN
aYqpnCiPGLM58e/LG+072TbkzsJia0+XX8Cnqr+4qQftKSFxgW0hFX7WLssX5oPI
BEwiRQmcpWwSKXfYLoFJABtJU5z3zb3ZKfq3C7DoK6SpfcFxfgh2Ey/e5DLr6YLr
ZVLCynkQ6pht/LEA/YE/Yz+9BU4VH2Qf5FcMFsvVjusRXW9I3VDKIFo4bMTouPaz
U/onM83iKTurXUP1OZ6Uas7zIxV78BMEbMuby028q3Pkz/v/9RzNEQ4OLecT07lC
rf3dDd781wkZDYUW5lAHKAR05Fq48HBDGDQvag4Sa8EF7EJc++xMuFxp3tU4BPlu
DuDW+yymHa2CdJExv0qL/Cl377B8syHY86ZAa6UVmRS4byweep/96UwYxTmwDIim
/q/M/zDoaHgkbmniy7ORqiROZoGOeVR70UmwK1aTw9Mn8TghgHztdIZRvB2S/bSd
YxvTVGFr8eZqCKRnz26UkPVDcSx63MP5CwxSesZyAF5IucnexPX9PgeAnbp2IjtO
phX7fCjmU+I2xpyA4dR806+z2kHE5Wm8wcp9atHduUDvuU3Fw0P8dnNUJFk04pjy
e6Kabvyp63gWsc9FLvzFPOzMuPB6BK+ZcS5KOSloytR4y9Jtfm5q9gYjSqUdx5RH
feg4mcPczfWqZlNnM4hxTSsorRkVK2v7vjjgzDirWt2bJ1TN2Aq/ptDZPCt+58G0
zZ1bzGeewUV8agQtsJidsllrCfms2j9AuzEFKjBu0i/wRsefsnA3nP2nT5Wu016g
EsLPoCLN3wmZTp2q1VviseAfmdT6lIJzyXtFNeBMDw9Fv2YLMtMLIKFOMINy1TBN
U1PFZ6WdkzDHTQ6iT3MnJumyQg2x0gDn8w+3/8/ZfSyqhuF14dnCBNX0ByXQpQdh
TTvAz7voHsuIpGBFCHwqpYJyQglVx6WPLXllq3gw5xlmjfrfSlkfKk6XWsuQo+QJ
onxajm09HWj4T2kYqA5W1P4oac+6uOZMhN4XmrxiuFRdzieioNpf38bcq3qx8aqL
kj+ove8NimV6F9XJwsNlHYqyxPRkOqeNziTWfjnQ0cvwjFT8FfCq2K5cGvA1xdFn
oDyzS0n3rFAoOt+MOrX9Y4sabUqowgIcwJ287aU9n4bXdgLD7EdRYKn7LQ24qFtT
RSku35k924KYRoWyJMGyZvZbuUhw9xndVexlyGzfamz2YLnxOS1Bxn4zZzFEzYKQ
U9rjjk5pcwRUquMX9P8olq2cwype/BfSOwvED75e9AY7WkaoGMWDhu1JqWEuku9C
nDW6rqXGLB8ahlMEK5hZ3OEfc4lwst21Kuuhzq5Zg/VaeKSNJPtoP5wxW0aLvT5h
5gdhiFLBIyvbDR6lBBmtP8G2jcbxolbuVgjq1LWmTmP6gWhToUGPq6fdXjzoWPAq
QvUB3WnFP2nsIUejbVzMUA4xsG3Z1aUXveSpiwIRDSJF/5BAYLbeiyVJrQ/Ih6Jr
N1I8Pwuv+5PxMYx954U54Bs1RHn2ztjmb/bezvme9CFPHzpAD7Y0z/i43QZBa5ea
a8uCxfY3zeRAiC0ShBAl1ww0D2iuS3mCCfGkWri/zi+o7kH6wLSNOGROltV1PK1o
3rgv0qryY8HDAsTiqj3W/PE723ONS20v2lIXgVmgTwkBE871A/g2aQaEKAHr9QG9
ktPlQ+PMDnMlQ2X3ugnwGjHkQauJmlLJ4E46+xzeU7YpLauNaFcGbuwIZEFWauvg
n/yk9fOaG/7469OtUOazA/5OWfNJVV8m9CXd+/HHs9flA4Jo9ZQFIOHYVtYJRGKh
4GdskwnZU+Ve2gT0PEBYebd+3lu7xVpHItppOsP49cPISRf0zGTf0S6r6wpZbiSN
YaL7r+5y+Yw4Z72BfdOFgBzT2KcGjvkn7HiEDKQ1Fti/QPzWQgW680YinBhirrYS
NIEES5NjuhZUszSBLCGJG+Jbfq//Mu9uqbXS3KbJTYVh26e4XXo4DZEu4Qj/wmX+
xB5IeQk2yNQhX5eUNOxM4qxGeNKfs7vd81RsV+jUSE+S7bonsi6CQ8r7+4iGtlGH
IUhylab+k/odW4hHQ8Kc6NzoDTo7HdncEl14gGH45EoHKkT5/SGif8+bkbVhThyY
U4g7rhjK0cfiL7oNcBKE2p56iV6ZrO+j6dL2xAEDE+xsmcajiOEQyv23sH2eZgFB
YBilvhDHOWSw+OHMaSmsYA5D6Skm9GkxqNeMYpWHVave20P1IxU5KjojO5Iw4W0W
dL5QT80novbIiRFrU79o/apdaBwz/H4PRLradWsu8XoBOEt19X0sso4Y8mrci6FW
wWfGBUHIfFALDJffAoBeV3dQVTYAdBlaY3+xim5r3CFlaRzi19JE2iE/W3FHUObA
b0+LQsTWBxPMM7XNDgDjO3KKswhBgWg/zNJqw4EA209GhtcWPafDLuEsFsVXXkAN
3n9PPEQeY/IthMIb8q3wP4RlZW95QCA2+36iaK3ip+UhcRJiOyG1sg6abHXQLJ6A
nCuDwxLUwAQ3cSsSDJoJ5P5k46c/1ZkHpmXeYer+qelI1P6D012gKIBmgIvoYFCX
CkWosbhdO/ABm3qvIsMNR6xPPgpmO2KPZYWQhiXNDzfL0esxhH2w308MdR2cZDyU
tHOfR8GW4TLiiJKe7Szb83NKkw5X4hksVrNTeFHR1bw4kse/rV7dARg8nsR39+ie
Ldriz0OZl0pyxOHVZgorDz8p37+3YUoZKbZs7F/VY8iyOYucrjdU9vM1MZm8gpSY
0lB/rDUd4zOGl3UszBJGVrKoyLiPG4Tp1JkW6VyJkhWEiRmDAo8bQbexWUl4lofO
mXWuvQu89RNXYJFG0JihBix4JyWI0QGSKn0QKBsP4oOtycInP7SEbUFO1AJZkgjH
OqVGe4RZmeK6To6gQ26IoPq/nKO0dfS2PXn2QXYz99XGt6erCWmlzx2YGNekr3Io
UUR+8gXhoVneE5ugp7Ane+EuBOCe4cG7B1Gr9Qx7I9d+8EinmT2Ctx/AeFiTwXjG
pJ2nzU7eTH1awWga9hPiOLgCmCo6/6aUM8IGSCSMnh4USDGKRZohrU902Pzto4mu
ujYcXzGhtEnONvf2nLXnmFDIUQ7Jnn7mugcWVqEw9jj9LUo+sHG2yCCi3mswYRRP
Ea3G5ntGZ56tzfD0cQinvyOyLi3xo9k3uA94To/AJ9CU0nWVzxa7Z8ecVcFZcy1I
oRJ1ewJcBzDYrhUQwPRdeY/sTjRvUGpdyy76SKV25J0yoy/J6P79/q0D3Ze13BYV
RQEgHxlqnSHvf6R1JI4vr2MoHyupaRBEpD+q9GwRIIKu0N6BlTsmDiQbopFbbxsT
dBT0zz0gbVe2whclACPyGjGkKw8ncIz4bjpL/3TifJ4LeQAaX3UNzybqOcCMD+h1
I6uyGXyp709RrNUUXjTWi66vKf+dPpmxgFFvb3LK702Lc8/VJ6Bv3uOik+/45wkk
0TdmXnWpIymUEQNZ2VlS9F25qRIVbOXEwEPSm5+Hc9hbrvtvSxszlpxahIf9aZn3
oeg6SZVCoF5U80e68DMLAXWnS644A37/I9uQGqWv6r9yChY5kd0rRPE70RoeDy9X
a5s5qHqLG9tIyY95OAeQvqCO3qNH3XBVRbsbgTS7K3yKBa3UXELmQKuHr2rfyz7E
Eb/3JnW9YkhoKN/oNjmf0KvMyaJw46mWB5ELk8SI6LSFOHESEyoHZvlEkf/RpsTY
uR7GWPln8euWHpqCpdMJte0l/h3z9gZstBCHZ1Y1J4cw7b3RHNcw13+BGqZx7yCh
KxVBu/XpU8jS4mJuFPfN79u1wGHcn2Os4q2BmbJkiwDV55KP0JJJAIjh2Utd8bBg
YYRGX100Cv9l+nXFECnqZrtg/RlsFTrK2wXygrNC8Y+ydcNTulf1vWhgxKpi9ycK
rdYe4G9LeGNimBGOOPQ7dMsdbw1mX+fUMxxDqqHcIEAmJEuEiwbpNA2zKXfffpNQ
iUSaghSNsmh8bLe3pf6DzToExWj6QxJexf1+U6dknoMb3hcv+KIzwWECxEgaM0z1
CMq1OpPvCBkNcpMkWuqQQ8Fd5F0AAQI9sEz2eCRTski+7foyO4JSnXhCQuNKYOMu
Bg7tOb4VMhT/7RdlbX12wa/16eWAKRcQqIc0aq92xvlR9cIq32JbxIRuaKMgMCNg
eLxuzmIgrIxK8hF260L2k6uQUNbqB8ZNHe/GeZzpWUrKY3oK2mk0CB+ZMgSkRyet
vws+AFA06JKS49BNJLyV9AXHF5IVou+KI7UEIFnNFwgFLbjbMhODoJeHH/Oj9IJd
Pqwx1zA4gIMre6s3bsOM1WFLOooPmE6mlvLDlHKo7LVMVJJcifKcwLekOPXAE/Ns
jkROivkDD1v42buRAxGvjXUDSst3r0jLXMZoGdef1sLtSaXPpaONnIYv2CTytFE2
9NCr3oohddkO9OFj0H54TimzgoELJ/pMUX3iBeGExMB7JvxuwogE8Y0ajibsP5TS
3LZQUVu+ca9EbNAxZPwRlmG/OaJLevQJ5TKwbX0JFea+rJFRgOP8NK/+ZPV72zW3
jHYPqnCxPXKrfWXJMTBAU73g6u3XpC6iYdFqo2BcWRtTCxjvPlKs37ev5TETcIY4
j7RiupnMbjTS7CCUFwMuJHQwU0qnqUg02TjHA+R6322RMEuPj3Lh1fOc/tXsSQmN
bDAPAI3DRiBn/cWu+ZWrybrM8dNhW30aD15qx5QZf+vgzcL2e2Yy/FnpOCiT0yXP
bFqPWGE1aIWhAfmTxKq2JWtt0Hz7tGeu48UI++VBZCV4D0AMIySsCAoIy4XPLvuy
K4fIE9TDWIa1z30oJ3TUWMlGYGha2tgUDT8fT/E2alWP8uL7pOuf2rZ82cbR8ton
z1e8cPMdv2k1oL1LUfASACK6FyQjfGkNsqvO3ybYxJb/B8ImfT/3B/55sXpJK35V
N450rzv4ErzkAiym6WAkKkp1Qhkc7DNaywKGUKwvQvIuArdXpUxAFGr+x4HBZESQ
za7EIdTCuqqFv3/lIyP0K/UGyd3KV3L/LOMIcgwpzf7bk43sUzywXVGcA6F9tnkq
ZLwUo5NRsZ1ePH2TEk8XB8ume01ZjbP8K39Jao8jS58m/l22RNiHtTdpk2vrJzUC
RshiBL8umEdllL9kJ+ZuIlXMqQN3bo+Zjpg4R6a+IsQyE0P8IhmQyOSdt4YoSWXs
xGrNqbNiUNQvDfq/2ZpvLzU7qlPh7HZXBtZEe0O+KNCgvXk59KYSLhnxiAl8lbYR
Fp3UAhkvKRQ/wQM927eSFdeLq7D9W5A8wKmd/XYY5ndtW7UG1NoOy52BdR3hjR2J
AG8sXitkc2cYJgnlg7Ur1OcLVGOr9QXuVt7M0gdawEICZRR6j0EW/wXUI7iKgm2x
Gufx5nIN3uj+m/1VDq3hpZl8JkR8AUZR3RpTe+5zkMi0gFTtzzsdOUHggU2R1Kfb
lE9Qjj0QUTlHF25G/X+FwMcLB88ChlHJMSm3PztmdnZEQwXg2XROFxtZptPX0fRv
h+8gMjr38XZRlQpHSPvtuBBrk4EfT7WDNXYDe7EgkTg7kmhBy7Adw+3AG+tnsCQy
zskVEqpg+m1rHdUOkM0wE1e91R776Hr5XWiBbVoyoXVreUzzxgLisHxZDUnchQYp
UhMvk1m5G6YdJdUGLwntzD2cmDl8nZ+lf9XGIqcTnGhpL5FzcgMuhUNCCQY184Gb
883lgJCu5ph09++S8bandAhstg+9Ix2joAoNnMpr8hl5ZVXzaGrATOu5p4Jxs13P
H7d/OC21zrjfKTW7r4PFcWY32IaYyWqotIB8EtfQQZxNVTXEktA+y3lm7CqI3hXS
Y7Nn2ylePOTeb5jVZQOIWjfBzkZUK8mVUtC0oc9vdZr9i+jaY7XpoPuzVMZdeP6v
2bqfIH6uc0H7d9XcBOQgGhF9sZyPzRK/XCJzJEDEfBjnifSUXc1CZk7DKVzNeguP
/9waFNr4agzuYcFWlMR+XwvPa36iBlwmPbuta2s7P5Kn79+O4p7rRzLrTiSaq+MG
rYjecZtOA5QYU2voi9H7De7FeZU2cax0EKGcWdA9dDEia4Do4lEfyKwl3pQaTNq9
CbcXlXGIphu3k7HJzJJL4aJZYPVF7G0qz46czqBuCUpKGquIA9TqlCB5TBPXSLlO
abfr6CbKw6uumK2W+LjSbjcUbqBP1IJ/4pPMeHlkJ5O588+2Q2nILbiCZjlED8Hc
9BWsm/IYsfHfP7/xv2Gfws3dG9Q2COou+ri7jJsjRKD4VQ6Jpo8NZ3ZU5o6KagRC
nDhSpPBmQlHWFEKb0mHTJuVfe9imSZz9i4dkB8HQWenwh72Irw/LbK61mkMhzkdC
btxLlmsbwe0HTzjD1pW/Mz5LamnjGZIUTXkwnF6vc4x5Dn9OruUWZPtWC1OcX+Q4
XzJ7VNj3UQD7v/PyY+U/NBOzyR8GKmQlWGMXpIiASQ/PSqfnJLmY3ueg+GN15iAJ
pSh4FC437oAZN0LQhTF5wSBQlOVSBZd6/Fvq+wyf/YV+547isvfXBNoSw2TDGlGY
/JGEJWdrWkcK4WjQHzIgBsLSTw3MVAo/bNdvPWMn5XRXlarcntNCn5cQRR8DuOhW
a6Q70iRVaEE6Z6972kleSuhK3lWGoylVh36a4DimG8Z/0qXCz7WPTMo3fL+nZ1vW
akDXm6Ctz/Cn1LUgCA8nvJp0DBgSn0RE95PO0jlMreVgwdKidOwv4/HZx+MVzBRb
tN9UQvLw+z1+O3o/bPRftzvLMKJvia/PJOlmhQ1+QxYwZfmQ1qwk1evWvSXgmAOr
C+3uh+jOUWD3EWPF5nqt5q8DYPwu+f4FqRfU2LRAAqsXcZZDvjqvHc42zGIRK+mI
Rat79QVgE/FVdJmVb1WCSiw8BrGedE0NqH1ZYRxWM0kBaKhXJq1I93/S3SsvoaZj
8XtgQaPOvRZVabl23xzD1H5gPCrgOEi4/CxFiItsy75qKQdSP0MemcDB3QSy+/NY
AbN0uBFFORZqgQq/XqeI5JvBcp3MuwWO/QVdLKpw07hj+W5S7jWfunsGh50cRY9F
WXAG3E0bArK/Cx8sXvW5A3rjMSn9HQOMEaFSPIQvOWhsIF4h/t+8BbiFP4Mm1Ebr
XU0jLOYUhbFLG5ZumxZUXeBXut2rtOZBhrE/z2cvlp239bsydcfgwMEMnd8zL18i
ul5YJkBNQRRMYHTWJA9YDvhfYlsLKc0oX85tYXrQ8ula/ObOIKBGTrmLmbrJdTJf
x/f097Hs1eFIdoOij2YRRusaQrbI9dwQjMQ8AlQECXzxBPN9O+wolXh/dE3sBjok
iRA+2i9DUtMjGTVkg6o5FIu4cQxAxzUcX+4O7Q2TUZgvpImsD6ahnj9QkRK+g5TL
XUO+Z+5Fq4AS6LtOqp6KvvDvqXYVltPtti0OcvQ/jpVdOmJB2fdHE/6p3TtFhJEv
9IHeQIQ+cI1h4kuKkfhdRwBjgNLqJABozw/b1bRYZ+ISai6oVrMa3EnF9JAOsyFm
ISdXF5AW3ZODpit0792cNxqu4xAw8p9q4B07eZDRG0UZh82o9sWf7yLe/juTZCM1
tQL3YGXi6GKs3bUy1h7rcD2hnTBtE4DNOOPDz0mXJgz5yLliFmAitToRdtQXYVjs
J4AWq3ieb8KM64HPZafvG6qa2c8Os1DvDojdrTaWnTJ5y7TMN2pOaeFlveT02eT9
Uy8ugyg2me0IIviUptCE6NnqC2P2KfEjitGIzYQ0mug+hCkWrHYLWHtsu/uz3Kye
PXPcwLdEWsiZzF94F5xKq6hPUN3X4L7M8jT0luEekPC/+Fq1KfgB9Gaz3A9cRsvb
QysEiDO1wYcrcamepuBi3z4bFzrhdrpCu9R623RaKK8+3og8S/pHk4R4uWpn3/HU
2ztOtpwA0HpUahZYfgc5jlHicajky7w2L2xclKiOVgu6MzhVNu9jaKCmzqe+eRbG
gsMjNiDCqRBRG+Dpt7IjlojTJeyhYEofKFhefIPSaPoG6WdzbHRSEVv8i/Sb0MJV
/htit3Hz/bR/ElW7QCKJNeI4svkSABFPK4QsuMHXBotCXk9fsbVvBJNyPEf1lvWm
D7LzYjGuK0F4WQDPbWs/8QIYj1zANcr5GlAigKNs4Z0fVYw8eRkpNEZdaMcs96s6
rNbM/IPvFCyOpqqvLHN6MOB9EfC8ANVxOjLpcntZu3yjFAofbxfUWvDTa6DNv4pW
EWmPRac1ASLmc8Kc2uiaUThCY2cPlq7r4PPiP82wCifOLUJmhXnI0WvAOuUCE5OJ
IF3dCWwREjvAaM/Ni8gMpG5555srhzPJ4zR9mxgXAYY/aUzb4xWVOqHdK8nPW459
JbXbTq6xYIn13nAALI3n+wkY0LNZE3f4QsTeTQypg2pKrUD5ukk+0n2mSt9A36VL
jA1zAMK84abp0ES/ZZRTVvfLSMVJTvlYFHCmtSj7gwqeqT8kjqslFv3bj34zHWVf
b3ERl3HpHrC99f3TjC//L5aKSM32UO0glXhl2UHoQ3ZpbWNglStdoW2QiFFebjA9
aeLoW7kx9THQnyk9talQKVSBvmAExi1o61s7+L9YLJElGgWxvGCYvBxpYRBwNzBN
jUIK+8ASPYxWjucmCORwCH8Id+1T6cdIGJsCFUpbBcbmsV1rv1d1UGudH0x9NKtM
Nec4UYFKBa2tTo1sXi/iNaqu4jWxudq80cnoxE84r1IebKnDZ7MoApBCPYaC1t/J
OJWZx7oumQvjliqr0BB8wnSi0yZ37usU0amSGczfibVMiYRWpxHkfsybQcmX/+LH
UcAg1Jc7SNN6l495/14gsK1+MFyxposiwWjFEPsvXS/bmKiiwRd3OZc4zML6IT4m
MUPvT/N1nAyZ8b1IlvS1achRo5oXdz1fqb8OZ8bH+QHkVng4pK77fDn/MFsgHnYx
tj7DuR8Lo4IvgwOyl7hGf2kcKbRiFtIVv0F8wwfEPwQmWTNppCU873tkbmlTQpR7
4bzflph2W4T2PV/f0pGS4pFqyAXXP9vV7gX1mAJmZzqVnqa9MYvcT3/B1P7JLh4W
sbRO7ttYHyDDasvxQJlOKrB7B48F39csy0JRNpgAM9rB8jySpNHo9J8U/UinFNEd
GC1rKQ+n9XvL83fKxwNZBu18qONiY63Hx3QKAXnOyq77I0Uo5KPSFTSOCYjNZhEb
U4KdYIUIABEc8cJNCkae/16lUC+AclxeUFR2JzUU1xSIT+S13V6kmfbzFqApzBj7
sVqhmPY7K67PVbeZGuB1OAbwKirnBPrzvtY9ZDZv0HbM6kxrrVKj+TVR161Aa+fj
ryXGog0Z9nOStVPvWFtSokkr65/xFNnPaZ4hIM/0fQlvRsxQrsO4VoORG+gmRJBS
b+wiR+kVRXET7xze0KMLmGinJcv0bWdx0K6vNmzBwNNDxfAPvzXab7CBoue8l5ww
Jbk3zU6jbZrjBnudAvSz0ieNrfkbZahNAf76Tk+BIif9jkb73tVQNQy00+iBacN8
iklS34fEI7wguueuT5VXKeBSvCyuDs7l3+6y1qhzDkaYHwrrwl8qmP0sJwR4jviU
Dg1v9L2hIUHK2VOewbg5QMv8jbE81ciQx+AAVAUYM7nPGJCVnibXWzq2UWgBneJE
oK3LybDcY7Td31pw+BTaBaCXk9pKgGLMKEMFxS4qpTPM30onlnIw7Ce9wkbOHDlU
3mFFvXpduPkiLOVrTk+s7S+vbNNa9Vfg26W+aN/nPgu60afuW+NLfE/dMLZLlgJG
FDzMfI/C0Q8tH8v5oinn34TNmE8R/YHK9DcmHl+rUlyd2EZJ7It4GW0geCOu07pj
Sq9IGjr3D8RDoBj0QZF92vbotc6y7ntZBij1Qj0pcuz+tNljXzeQP6abgHIYASoK
+10F3hhWSxdCKYomoLRWB+3fwkTCV68wW/2acJKA5Jlteq2PCNTG4ik40TjpKyxW
AGxcYGY6VSAIwunn6Mj7iKbb5gz2PrVJGizzdsF3jDEchI6PU7QhNVIeAen/nHfR
meb1Z6fQ+AbB2yxvof9BBntLGJ0Xb7CwJtGcsWnhJvHKEjf1kCa1hFaCkhoCrnaS
aaeICGms/bR5I8p33Sx+b6HuRKKwbDL532UqVSVq7GFgBpVUzqOZ0lCl9dWbc96F
n0YKyawl5rw30a2Op2m2oEH3enROtqLpSmnPXW6EOrDrMjkCWlJoxplZ9qNJo6C/
xG9wz9R0pBC6ud/FeOR6eVaCqODsCn+bHBVFl7umUV09toKCZfIQrrAzgD5H8LBL
Pykg9zI0AJshTXD5nLa1zmVVIlxYZkt7F+W9IuNw0Z+Z8iay9+ru7uGS2+0GU9yS
XM8niaKIMEjta5yp2hFtCaJH10NePLERR1zcqPT76ECTDU4Q2QnWQF2i0BZQzbKd
NU56Xp4EF5hlgfqZJ8yEvEOKpQg6BtcbxgE6sQ1SUxmGQ+wiMG9I4f2CzrCFNVnn
likRvP5hQugyNyp2GyN/yTTeLWhln9xD2amSfVm8mNg0fN84bv4NzArG6MY+7geu
Scm5IGzpD7igmdHN7NA1gVRc1NBTRctqmlDSbkZqgqwuEEeXloEw4s8/urBtd2/M
R2E+rzc2gPrbpazOnfaQhqxtn/H9s2QFGfadzUa9cko0CcPaY2J7RUCzb661xiX6
Zo5OE2X/4yH3gch/AAjAYnDm3IMXjNaCOCniDJ71uEH0G+v/j2w2nlJS86afo1RF
ptH0DFp8vTfeA95iuC+pGrLgFdvv/9yxQxyd4KtGA/6CNeltAse0OZ/i63mUTvrl
yBfLp03oHBsGuQ0DwTVPBI68anWNDocDLfwWJrRoVv1zBM3toXCfqQDuFkChJXQo
wjEzcoenftCbBZWgNIg2c5QtlNPY3RCvfS2KQ9Mfj7a+xWMjSueiDtz/i847lWVL
1DDyWtPEgDT6Bh1AXQU3NOG3C2wZt9DPH4P+Y1puoiCwL0p6hRT+okAiY5/mPEus
B5dqV95zGrX+i6H9QIor17HuqwWa3PY7EaXZLpPhKnEtgCrXGGouTQ5fam6fXbAs
HKaPpRoRo1Opa2XcBwT6xEBpriYtePEFCcaJUDmzMdDfu6hsOjgBYKRzvZkNSrNO
DaCoQsD4tiS6eJZI15qghXNFAHNHBrXIgDxU778MPb2mN8nu0tlmWA10goNVOLrl
6y3IEEhGnopiGieJx/xLOFn+wmWLqws1j3AhqDLeXxbwlUjDjDTI6uGxWl7wpxWq
mxPENAm+IGm6tr5GIWI/UGsSkz06CE5ejtqairslYuH1bYCaKMjisw4OfmyrYl2i
BBg0vrMa+mDpGA+p5lboLkOqBEYmxqmX8bwsqRaK0q6INR47Er9RuYb02OmjLBc/
iG6MIBE2UqJJG95ZZ5b0ZFwZAmNswV7FiAmaP7avMKyFNSUJFCSbsZNr0GlfHt54
wwOCoOceIrClVhIR8pQL0Y9PI+dgj3M1tRo+oQpFR8/RbHOGwWrinQnPmovlW+YC
3FV+9Zfbio0Hni7R9BTT/4ccXU/Xaexqtf4beo+z0KimwwrHVLCpjmHq33LyqNpS
ND0GkmiAZduP+7KWJm1p1rL0l7j8yzUus5Di25b+oqk8jMjJVyxJOk0VvZGXnaBA
Xtlg+ZICQegUqGd3EOiahA62eTc4QEKvoUpca/8vNuJk6kc2j3KGrXr5G+Zp6Juw
AHYVFVB4KX8ZhSdzC/wjWGb/PZNvKvARHWDa5a+rInVzJJl6Wcm/JMi6BWY5zwiJ
Pe5bL9vWiUqIdjV2CO8eIAZ811oPHTA37ZbtDuWcFstIGeY4+/sRpFVgbGHWYqh2
SHLu+grXnUYEbY936cy2ZiKqH7oE6UxsIIuxDWBpncg0ph/lsbp/f0F6srDgdUTo
UCxRPzRFKDnVyafupWSMaXOAi9oDCKfcMEHtvk7d9krU+b/h+C9hdh1WlIFbRpVC
/2XRvOiSqk+KiAU7nvCzd/3M+zG3cHAn6t9JryKZ57r8kIJ1OwqfVepaiDxx3gse
d+S3z0z0IQeK0VHMCXwqqomy7kWTxAV8XIYkcGMYy4qpQrwJORtIX1dupusAq4eT
60XDuiLJklpcIvvuqjgWQsTyiXQhEHWOeApEdK/MkUMa8UUUjtWtkxrB5Ckd9ifm
xzPoWosgTo234w2Rhhf4veYegfcSnH1j1IzxtLwsY3YNVP3juh4gdbO6W4PfFeSC
uNbScuqUWjcmikhV4vMw4Pn31uBjiwmarqOJpAcV9zEwDbbpQ0ZHU7OWT46iC6q1
D/3oPHO7eM6EoLldCC3FVC7OV7D6GR9n+7h951OpdNa4a2MdZlrWynqgKw4xlKhf
Hg4PXoHyb2kZed7h2SB7SMNvVtx97imIzmGZ2pbQ/hy6W6HPkfM9s4+spgf5mext
V6VOTH0vtwKxf9y7xrKck/olEhfGIgu0hq1aUYCekPOGSzqODqsfXQjL1MGaozNQ
VEOLHsBFaX4iiHbov8UPJw3tXsGhUUsjce1i+rxRVg16O8Nr7iEymEWjIRVIzRbq
eWcuKzIFPiBkp5Rh0FAHoKTm8XFTWXmFY2jPJGZM/Wi5WP0Abk2sZw76fUC6iEgb
EMCkt1lxmCoIneGz6DwDav3atNfa5Mkgy1DR1CRZ8DAI4L+Bf4GKeH5GpbaSMmOm
3/Rm4LGObDQt7Tm15bNBPilFVWRQ1oWgyWninbeNByDzqPw+QuBGCX4EKQCVm1Q5
TNiP/oX19/6atIKM5lkPkpxYk9esLXe9Asfuxgi75I2uuCqiwS8cNRIo2L8S7TcI
fMYmKti1i6N6HJnT8342vbXUDG3XwvmYLkv/xqN5sA2CAUS6uuVQnGLxe/x6uPNn
6UW5tUCo5kOfmyOMeRsE8xjHXfSLlj7WHr6QOxVFpoHtxLDywOQQFGUoSx0VHsCk
Bkqz4Tqb1VaRuv00y3MGEEf8awqKX7ZFieSRwQer1qx6+tMn41dtzLIQxFAxFZaw
+8fYYOQHummpGZNJ5ekBJVRKZN+XydSjvlvhweBQIO1+9pUBDCFrt7qRoS+1bL5d
oHV4OsYfrm/7i1Q11ysEhrSydCa/tWJOv3+IYvhJtpg0C5pj5UekFU6I3Fy1DoHG
93yom5y0QuOhqaP2y0shQbvga//tmVBjyIzPdw/4EcCw3BCEvqusllCj4MZqBap+
WtY9vwD388ns8Ciwi7mkChT+z6BRqBGWHo9Z8hnKIzrnWpKbzFn71uaHoxG8afZR
G3vqW+iq0ZB7TLEHRdCSayEoLL67pUBiOL8IJUNul4Wud5RKEojH/sIU9i6V+Syz
I/VdBSbWNaUDRj7DUpc175q3s3qSIB/75JDHYTQBJtw3oMbbKYnkC1c8YgkEMWsv
P6HfBBKVdyH6k+VUGOz+2X3F2A/GCWyMlFi2i5RD5pzjGhLTflIRymECspB4f35c
S4hx49Y5SMRpl6GjSIJ5xrj60zawIHjARtcgeqyW+18Z5/+mzdAjygpUQAmKYsDv
QTcPqM2hs/v3+045jvc1KNHvqMOgvAQsMj4WAhn1W5NZIA0jrL+enU2+hAPw5DCp
hOoxEYb4YfgFR3HjTuMscrHXpmPQAetlYQ+fd1ihmci1ADylxDiDSCtAnamAQXoY
ZdnZ3VKbGg+4jJiJ2yh6g5Yg5QHatjCtyeTrgmJb6yIXM11+JC4xrDzVNTJT01nF
EURU+/OR9wPaqWUld7NcT2NqR8yAOna5YYtLVuCUqtaMKAKnSh4fEBwDfotLbxcU
dwFCiu2hhKSGKL1PVhb+M/7WUF2YjNDtoXc0GA9dp7jrTNvmyD5+5E+5Ta/dHTkn
fpO9OBCTj+J8dU/tLoHiqGcr15BTOQEJdduOOfsCGeMLZZKlk5Xp68yVahLKzIk6
M6SoJ78bOJW5K7CdKUyx9FiCyp/4I8vmsqrbGS1KgJ6jY2GrH87oSgN6sPrd8PjS
usCKag5p53MzWelK9RCJ7kJ9UWyKXhbjmdIZYVem5AC6ylB49+E85nyZVSTqUeUa
tyh4HBsSMSMkAGC+j7jDy4IRW99dF3EebMDGLsiiTY8rA7QRRS/wvywCK2sWmjfE
wMBdSfP3+GHDKN0XxYec5hb13pHeoKB99W2bm0vMUDCjV5Yl09zy8cV7thKEVKNW
Kb13ibPv424h0iWpGHg2qDDwKV2WwD7NGNKyTxPBEMLmWvZ59X4ikjNZyxqikhRI
5mUcto560wtFKUAiEu6y+WP32KYWWTzFOOVo6U52AH3mCZctaq90QEZz9YHjrzFS
SIVQKozO7/w4VHLOm+8F5EZNu3DAVv5UuyL9CR/g2c4pvFCSF4wgQOd3S/RC37OU
8puATDay0wsm2Dui5kO79sW+rzrvgW3zShjlyJlxh3c8uYH3s1Ri2zJ4HU/+ttvt
hkmJSOdIjPJkh3vFzjE9cCjA49xiKu/8evij475juguVa7npvOgIGNFZvTRuO4Re
umTwyvOrhxEaguNcEYka8kLPC1XHDHw8WLIYTFph3oNiF+sHN3q77xNuKJH29AJ6
VZPxASJhZPhYtAShqH9tbBIzjxtFvAtKHvmIxPIwdx/Knql6vxv7ih3J7ALgcSD6
1viXEpbWxQisYwsdFRmO9v1S4sfd/uHhIR0/rBPLmcV0oWvDbmxdQSd4Oof4KqrI
jjp5hCOLD3alqEE03ytlqL/nSC0N4j1M049RR9vbmYsCUtKUpnJaIZPk8WECUSer
vlvou+3S/jO6z7rnpWQEVv7Xm/KPUwvM6RtCmkibtSAiUIYLx5jQYGmwsTC4BVN2
DlQffunCeXActhRygdAXHBIj77OKArdnvjhQtau0uJtxgsi5hg/7skzdhC7iL29T
9BnjdvKDZlO6dGt+rcb6wyLziSUwM+7V7XemY+OMG3XT82t7kDdPJOj1fzZPLmOl
QdFO8NOEr8NJ1b7ghew2BxrYSxpqJGi1kTCS9r5EAa9QNoCURS8nP/7VwFf78UXy
qNI0dAiopICRbB1pwwFi6mTE+xKuYmwIiHwL4R8fajaBMnD+ad0gGPH4m7WOH0SL
CIHJGVEwvbpU8mnlcajy2Ug8TCuCen3EllW3yqDa3gmpRPWvsT4u/2RBQT36Bggl
4ZQWcQLF9XYb/SI8PaQdpuDJNWYdKBXPaQy0ZXK/iB5VkuHCncKouQZRzksy0TZG
xyUUYAaFJb1whSusePo2OYUDqvZtrt3xaKN3ib4e9XUCiseKW6Mp0ImPBJ+L1VKu
Uewhzh5EM202Ao2IMsKP2WJCxeFByH1ZkFpAxIFaCWRA2m2kXO9PgbcLjjurbwX8
yP2LMSE1n5Dsph4z+VtYnRJ3Kya2+cM67EDcgZKeUJ+1Os89WIRhGvqR9TkESBVR
8d6/wu7uUVJZ264CBdtCXHjhtAPYvuHi0sjd99lSZpHQjuGjOem0XDaxPSpHg7YG
3AtpEpqpTAzJR9GgW/rVuk9RrCoAWenrTGP/BOHQpaoPPbYiRlFVGtJuO7TmnFdF
RBHpUmaa6xdEk7DQ3y7Cx5ZACsYi1UqsIJtCSn+F6zH4Mf+uBQTEFrfk/dE8MGgW
yOZ19WwNODeA0DE8ln4XxQq0JyRFsfiBjRsEx6HMrMB0mllm2CMubjTsZN2+TsPb
UDJu6Tc8nAghErdProz4jnfm/VDNpEhI48ZRdNW/mYDh3IyUQnlQ/Gjt+amOm9xU
j0VgA7i+oJX4wU3BfEVLxnEOCQP8lZdHt0ZCc585rLHNs4Xb+cX6+AcEm/uysZhU
Q87Wvh5fYONNCgUchGEVj/ZaejRXBBma57raz/n22+4Bln/VoExM8KINo3KI2dz0
XtHBmwt1qaM3JuK8je8Is9U2EgwdFaVAzCW6yKI5+qBMdgAR9A2UPksXyoss/ZUu
/9a5+wkLWzAzgF6PZ7zm+mAtHaBcVKVsLfrmJweksqFTuV2Aitp/x0f5yJ5mnIX7
ZPpPOYKBF+gM03wEgH1UMKPIEYKcIfni8J4qtI9AP6WCnO/nWwdPLaEULq+/Khmh
1QQ3RAix66vKH692BWGFSbQMVcvI+rKp/+u2kKWvHnoZACs9MvAgvpOk8YwRWnkJ
I6vozpk4ZYITfNydPka/Jb80hKXeMQzTKyChzEI2kWeyG186ueVIDbCPmbPdjaCP
/o05MiHjUJT/Fg8fQoHnjEdvYqSfbiKTIJU+RPVLrLNLvEHzN0C4+DkiDBGVLuoa
NsVwywJUhJ5ocwPGgZ/PuSxnom79fq3gFeun55p7am+fZFtSYS+Hwiluf72nwQUB
Adtj+pSivAAuXMNwMWQ6Y+MSFnKV2hCG7PMSDnLkDTTKUJGsJVEx3piNvfTHWWaT
WP4Rtycjwb0LcA2LwaXy200Tngu2Y4U6icdM+fsHqOhR1OsKJHxKrPBKMCz0r9Zl
0jT4TSRYeGbb+sNqalD5YS2zglcmvHdy+rNQwHreofQ587Y21iqCYEggIjyGcL9i
kbBeXkNFGP1p6/Aypy8KGqYsJQZxG23L+TWVzgOHawqFtiHtvoGV5PUVM+9iEXOw
bgqj9p5RaiwqWi7Z8V4MfFXyr7+Zj+Nmz1+/nmrs3xNkS/m9baOjyfAn9R5GL7Yw
pQeLN2TAhBKySLhGouMZd8BbW6jdzJeplMSVp6DN6fgCSZioHbaN0OKKgAkEO1p5
w1s89itepozvgNAZKBV2VmrIkxz4AkDbrFxkNQMHHBaSDBAwXnVK4Tg9OioYGh9a
G9GZz99bxG5Q3roJWkrnJZ7sIA7l3SjVLRX2UX2tqqH5qRyqWYFDIRpqUxNZqDvl
EJt23eP/N8HUDbAoT9jvKgBnZjVHLTcr7Wq/dIonrgLn+6n2TiDkH/6DDjge08+y
km+5r5QazE0IXLTN28btoF/yA9vTiMEc6uF/wSOhFUW3rodD2pAkSxUofK+gPSfb
6kajvr+CaJQtphocUV7gPwO1NrH9Hftl8NsChTOVnBlqvExx3Y8EDLqAsolXdeDe
VJVcATPgeVsdOVi0wfsu6CYcoohl+OH7bGzeJ2A224NrYsqX/Oro7IK1gAiVtMgv
XrMcZDxtZDkQeKv0FYbDmMxDnf2NNNZM0oSBPvilw1M5N7tH5iGZg7DR0FJ3jA7B
5Vj5g4PXtrpyplyX6b0BZbJQFryCEuHdZo7rvB2gijfQBp6PEmEv36yEHm2FTIZe
fK1GUMydDjgh7ntE0XDxdikuD+KntNz/lvNV0XYuJEqnjBx/SxwvVCl2/WZJO/mB
+9MZCdhY+vmpQFh4pMy60vCE2wXsIUMOFLvmKwYq9mWbFkq62oi92OCa5ZoSoU9r
PXxXUz9pDwKJwbIcRIcZoA05C1y5W3DTCPuVcFISHf6uaf27pqWh5qjC+5voUA4Q
TdMlcywoCcR8N62XhfpW2pHW1u9ATcNCCHFV8VWSwYQIxmt+6xYu2q6MHi64kqb6
IwVQ3mSxMXTdZb3oX8Oz4gDjus+YRx2FzEziDFlJCUrMPTx/ak5kDpmYc8iWOUBu
SuzYOyhxTp8r91xxpKXVqmt16heD3X2PyByzK9utvm+KBvweiQ96R7IwoLdgSGCr
Yqr1NkpHctUyJ6samdl5qwzO75u3PtkGtGqjO2OGbF+i1eMw/c8XFlNLtw4BHzuu
p906pW4gJX/xOpR0EdzUYoAsYHoFd5KmmvT3Mm4bhjXLT4/WpOelxahkvrrTmnv4
reGtuydlEgTFvTnouFx1+b/g7hkn5uesOYA/ioDci56XqwuY4fZbulVaCajP5HKm
cNNlnCY2ggHPpY3WtsEGF/ykhq2Z3q3M4HWi3sdh2k7T2uKq9AY8y9ByFU1Usfuq
4DTvnltkgFw/2Yu41XGGVqx2N2ORV4ELoBKF7zNis7Mah2E2Myh8X40zh8dh8Osl
9CKvmBFN8FugLFTKcmi2GUMOenxazXFTsa9T16REtc1nLe4taSGw0MAqZd/8DVZq
x5eangSGrYQgEsCx7j/SL69+W0B+JDos7pZtRzEMEhlxupEyx/4TUyKDhdOUfGki
AHarlgb5ML5B4ERGhlYuUKXJEHRoKsue+konyEfHane+kwAvl6qXo3CsXj7YYY5q
eWZGs0iBDdztQtCdrRyEuluzP2iJVTM1FSYpp9jAyOc4qJqSJCmSittOF573Z0Qp
5NqTDyLmWV8Wm4ld7/UvLKiY6U5SLWfSO1gYjYdZKWmr4bbWGWS9o+VXZh0bKtR0
xe0V0YIlyx+10Exr4ySBsHfuPfY+XATsMM4w1qu52uKw9N4uBjISrHIcfpMl7+XR
zmavbEEQ0CRLDIwePmihnuKU5wKieCHfcbIBD+EWmQZgRHqkaAZGBQdsv64HuCip
93lQcKEhTBfuqWFeKT0wDgIsKkQm22VWYwy0DgxWKFHTPTKGCyseIAz8iGaiavEM
RTOMxX62WVqCvbv/sqa/Ql8m47u14kBLJFJyYBB48/5nw4yeOWVuQrOwS2T4iAOM
ohW7ZbJxtnm9X7MzMOWnc/2aQxntLxq6fdZjpbyFc8KzV8Rg/b8hmkmL1TL2Bmdr
1ERn3fj+SmSTC0lEbk8loRyAQHmhioGJvTrOYyGUkyriNWXmA1UCXs14Vy1scCQv
8hlznphH8DfrHx2KNZSxLIQYJP09znJF43VtG5U7C122tuEDXabogza3gIlRCf6V
AS0volgpvlsVV8sUPpXw42kwiY4YP6Y7ZhxAmK8as+L+DqkwaDdweN6Nrs/Vp2/K
p7ncdKyYs2ZkiXWPdgMZqGsBf1IQgfbSGB68hPw2jZY8x3rFKP2N9YPZmzp0WEH7
WIeSwfF20MWf+iBplOkJGESOHiRt+mecTil/p21FQS8jA9l2eRBWj/6loaBkyNfB
44jNZ7ZUv2b5OoHu15xGzr5VdeCxWWcsGCix7ybtph6WOuJPM0NndEy6jP3sehEw
Cdw1fk/zYQsdlJAivWdoRZJYXBqH01PI8+/lK1aP+D5JcjfQ1d2QYvUKuL90tEPD
NHiD2Gtqco+PtTmZkFSPjfq3EE4HRumntKw0/+Y2OBqRKXIqq17a9WRmb/K8d8Mr
Y+LVbmw+UYnA0UPOXGwAuZpHOAoMdH0oHJLOoAyYsEbZFsqIgHac7ydq6ffTXWzX
wrD+aiM2W5CEwUj0INbO2E6QR4yvFLthlwbgOrVmDhz4nk+6+UZzVnKWaootuI9u
U9Iq+gSig7v5KsUz81oELLBpSbZ29gSzMfG8bhQOluaWvL82xrQ3AVKAubTJu1yF
HvOFWOt6ITSbxDld+lnHocWYU+s6duzqXzQLP2cOGz9QKzDB3G1OUQ+tlBwEwvjy
NpSF5DqkvWs3XWQaVo0hljVZ6PjwVc3ZF58mY++T3oFIcHlOGGEm5aE3ERGKrIIQ
0x6ZWSTYDaKGBO3Q6ZErY5lv2WNDaO4a5tC5oTILj4SaDxu9Xu8F/a2OaVc31aws
SQJglNlFdLkURNfg6wVZI1HoL5LAhjrnGW+lATvZ88Ahiov3AFVc3KeYXUnKUiTV
MqNoIKsq+GDiYgjwtXUrJdk8DwKSYrW/b95oyjDW8v+gf2fhfC1zaZ2HtymRpdE1
ssfcOxBrn98L9vc4vpd/xR95ZmLPkZGhYYBa9b5PcSgPW4jEgsGnRmaWoowfExnY
ITsbEOGKfEoPM7iQp5VSy1TZsAsk0GAgo/Nzpd7I3PIWRYtX/gkV6BnFlx19EyNp
ZgAZUSdSlnecz9pHlN32YIaNxKeGOQagWRO29ZLYk4EXzsYgHNqyGlIMRhTVvCHx
Uk6YzVQf0ReKj3OTO7/9KnN9oEkhyVcMm38MfHOAhJGPGyXAqo0xjVpe3tGX6QB0
aLMV8EQdtACMrp7ONg/jzjctcqHrsGTCfbeQ6a9y/bHBr5TB1t4zuMQk9DmiczQE
cnHT2fQloOQxy1mKli+Zk/2Pc4lTMDO+6AgMDJh/Jos3arWwHUYQsjQhqVZyjNYa
92tGNjQmaCZ681e3aoQk9pZXFFArPRZj/NbjgYoj8itMJhydMLBH5NB63UEyddXh
/JjD5uePvULPI6rIO3GyPafoDvcAh5BZfzjnGa+TA+RxYxEBLY0X93Ot3NYPvZiP
RaeR85D6Ze8HwfKDiKDdiifvaG3TAN3tLxAdmdsXhUXJsWkwz3SumRUfrPwQ6UWi
Q9Wc2WKA6UAswMV6FfQ2nkobpVRO5eR1AAPwTuEeWE6bhAoO2xyi8D5LRVrjLL/A
GuZABI3cVyKTumiMdA6AKN1CCpQMwgFQemx5i+sgsQnaOXmnuL/8DwtzuuNDtUxI
b6/7CcgdJH8m2aggwbEIiHj8HWnh/yPyJMF0zpJ5lUpyvHK+v/IYRMV5wmQKl+9R
QFaNVcSKBhbD6NJdWjQsSkPCXbvG7vDM5UerWbAe20kwe8QN7LWU6g9YXRGl4ZCG
6MrkblyF98spfeByQEhSuu3Dof+3tbv2bKzLs2ckaCpSFWF318u5KtXXkHWSkJIz
TmRJOgQXk0m6Utk0C8LRz6F6L+4DnJEMrhmlbBuKVGEQVXRA8kSpR4GG5waNx0me
vCjMjWAwXxSwcXHEDw2yM7paDc7VgGBGQG3VgQq+4J6+QC9Bm/W7rNqmxUpUAEa1
vNx/z4d0vO4mqLaOb2Wwjbz67UTo4iFafVdvzhkFyv/1XXEFdvf35oeQ/WekwoK+
NaGgRL8gtxM7969gEzNcV+LLOuZd1nqXRLGAV81aPNiD9/2khsC6Igk5A5yS47Yc
Fhf2F/DcW3ZcQFm0/1G07PQt9pmoumJw5J0ZzcwZGv+RwwTF+mFAjkgJRSV9FxGg
PafF8YkBzDKInSmbet8UlUMdJ3SH6Sb9CvGfGXzkXKefmuHkyKRC6pwqFDZ6i+3u
efB2b/8UCIcTX+NMxQ/5pKjI9pZfhVwOEOjTEJguu5dAgSGO2rOWSXHERLpxCVsd
AAA3yhgGfFe6eL6vTtk1XqnxPz4zJXKW5Up/AjWQbEaWJdTJECGRjQKzGFrR6pBO
ElVkyUduUPrab+acBOWnnZGBxPgGJ7aIWoJ/X2xejkTOha4EfgR6Znb3rmF8QEAP
NGWuyiSjoYr7Lsur3ivPerazE6r7to/Ih4GiXhvoM3Zpyc7L3FiSv9S/v7p3bOkf
MceIhEyAX9pnqrW9QoRsWJBXnxUIdPwLBBY2hu3zKq3TTZzh6jLBRFbKiLGDq4fL
BO310SWVrto5CxkgOtA5l37pOQ7wD5VA3SsuG8kkXzz2fMNzccFHAUbHT1yu8wb4
vCrpFslV+EtOSAxxYut2jn6Ji4yCZ4bkvE0IvezbOzeHp0ehvi1llsILvtZFMClC
OhMznVSUuVu/mxNBQu0se/CLY7pfK2oBg8Zxn6zt7pHIVyt+VVuqDQAIgd3WYUA8
CHoXlN5hNtA1lA3MVsz2PCDOqxFaUY1zeZmcPZBF0Fu2wSVy72rhm4FLNHEFHQV2
XM8x1vXWXbt7kDf8Qols/CWttp83CDpCr3I66WmXlscWEo5+3r0n+6yrxp6dAkmQ
TLwjQBtBhDp1IgzBQQxbKGbGVCFEmYTqo1O0e0ZNvfSLpbffWw+D3dSR3moMfUkZ
GTRKhHM5ceMEMK6Fa3gm9CqLuGATddC/kzZImdd/0Y5VHwbpc5ILpqPAVstn4Lmo
zgQn/mRpdoNQfzwtX/CvR7GJU4eb9b7e3qgCAutPZUaP5M1+JVxnZEV4sApcQi5A
6A3NSMK8PqL75cmoeMs4Ls6ItvvWBVsHCI7LGsvgjur6VkHRZ0CNJXRyzIMwm3Bo
01heFfw67aOt8HT0L8fn5A3gjJPxrq9W19kj8HKfP0JkqJjrsYiLviEZEddRbAr0
nhIByFuNnh9MYxziBxTdxQvufJnz9AECXnnelXC6JkFOPnzGyeAgJHAf30nJfhle
hqCv9pYMHPDH+TOdcBcpUGq+zanCGPZ2jvMBmFltH+qKyLUsd5vScVWhRudyaRue
J1hvyyzBymSuM8vOoiBBYWw+Tf+hnsmt2PqNQVOq1w0deQUdcmu7zjfnqAiM8aQB
JWaLGhe0wJnM1J7hyC334Hn2suqsk0X+1bKd+whae74sENab/SfYUO3Gfcg8/+f9
RcsOYWk5XMmkFdX5RLhJfT+5/xoXUd3WyLuoAogNykf9GkdIw1b45CZo2Vb2jtg8
82f3TuuK1c9fZLh+ZMuuwfAXmktlSulEOfvpxKLeunitGK8Q7Tx7vETukR4ejXjZ
2DRwyxBB9sf0xMM8KCNm8XL7mJtlA4Fl0nGAjowQyPkFQWFvyH4jWwURA7R2y4/l
kB4GjTz0w/oGoBDa7LzYmvgKiRMOYEpE5SjmjdFmNSv8A2T5UQVUHa4qk3sCbWXO
+qMEOspwJmBRR5uy+QHvR/WtMUQTAwk5iirie7F9ijfn+KVYSF7+h6alkIENiVxC
RIqwc7RIE8Bw2J6rmboIS+EBW4k0EQ3F8zC0BqraXxvXlcy1BEF+9cHfRBbTxwb+
DHCRJ5UUdvyiOTGxTHWmJvKkpDYppBLdplKM+q2XZcEhpsquBzIILoKgw+eH9YPu
d4PsphI0bFWKS0z6cdHAWaiUctT3GUsoL1PKFV9GhqSAn9BEtP76TgrlHcItJ21h
mfv3GbVrYc7ek41x2W+Mrw7S5HriKP9REpdYtsNjyJpjoUVaB0SHpBb0OGcYEtlG
AxNUJl9v/XBYabOfg3o226mPklRcYix+aJCkLQPquQGOvbGbJJOrmPAnwKp/0ne8
9Ow58OfkO1SzBSjLCpNv54YbKaPuSMhyJzX1toiu+DpAwrtABmTugkGH0nmv6diH
EiNvLu1KuYb3u1lQw99HMmuIc37ZnmoN8iZkXo0OZ1vO99+FQQ+e+k4xQlAC2nqx
8jzI+VqiVDSVEBFYBiJAu+gmXTbJSdo0WtqnZX45nlSp5qpJYua8uAWwHj4Ol1hL
EqKVg8ln8rUtKWI6zeuDu50YfCvOvhyLqwhjQoVlB/1HypJ+Cf++X+DOc+ZSrQTq
p6BPhmUbdMyIWIkg1HRKL9iV4WE4zPPplxUpzBNGwF5sXfjlSxenjezQeEwYQGHb
/heo3+0h2eEmsZ4XnUEuX69gMJTpL/gu3sySuXn8rmop08XVaAD34wJX4OWBn+oh
9IRdGWadLdcKcBOPGVvuv870Ecx4RkQbISubG32noh6kVRY3fUZhGH3/S0O5C6Pm
U0IhDGzVpO02yIgYwC0hOW+naD81Cy1tvELdgkqv1rumvRHD7yCT+qg2szJ4+b5x
/83CtAj9jAa4/9chVfAY6WSDF2pYym1Rw3C2GSmPo4PUk8/LNRpBDJq7hO+lddQ8
w04BH798/io007p0l5kSTSrDvdGFZTkPmEMIQv4CN1aCsCkAsXrt7vdz6I5uPxSA
criLeS418LzmWcK5Ozz1xVv8lTmDMSP0cbpDznMHQRcSkOjOsU3+k/oDnGGex7e/
zbHPO83AUp8JtJTcaCTliQxdShrVwKxdOKhFzCyvLvmHKaQWM2d9IwL09IwrqDWL
OaSO6y7FKj2T4xAs1wwZKqnZm/lGPWBkU9/kNufwtvzLkHB5E4i6YuQ1zQ6XGoKc
psRauC2Dukqb95aiAqK+STgQh4wKafZUFOGzQ/q9BTkZ1GD38MM3ZE4Mx2vNPkZJ
XD25rCdwKThPKlMwxDt/z/vr/v8WBEY8OkJo1WiOfSYTC4hQcekCJPOUkQ1vfaC2
kJvsiHoJJ2Gc+b/BJHSFrOzIHn+Ntu3vIui9f1qrJguHevefu3A1JRJbyzyOJRn9
V7myHsFFqSzYnB5++iNFeWFgEYRjam0osrFuR8gQpLuddOZZWB+KU5ZEHBJD5raZ
JD+hO9Z1Wl+aCY3OBiPXIgzAZgSQ7PkoLiCrCAhhmzJIyjcFkb+I5uqcfoTIMFqE
AOMWITXA193WtTyIOwGVvmf/nZUABToBs+csLgstwyU9I4E7Z/nMUtKLBY5KKgkl
4xO3yXrL6Fqp5kJaV9w65e7XqAurJPtmiKrVxYTOcm7u8qW/B5fURFBOno//MlbY
mB3sZ7o8FD5uUfHwGltylRMrF3rPJ81w88+cSOOSGF5USKOPT60Y47NCoastsVCG
NOFVxsJV33AZdeUIXqmDr7f9gbPnM+IKR4/HXeM8P9vOZg9mPhDDCAyoBDcUS3Py
13a8M72bYmbv+W/wJssrjz6CCEzJqes3BgmuRQNIt6YAVs9+srw8jZ7t5gOCgCwu
idz6ViLCXYPHA2XKKZW3JYZiCY5IELvx6T2LoW9C3NgEPhSGPoHjJrh7pZQ6lJ3N
Xwg01BtuQmYO6GGqgSqDKVMauyzFNXAVXj5yki3WKEJL3ZNu9bu/sfBtUxiZYPu9
WN7X3ACtLTi2g1iXV4gY9NKD3lw7iviEtRFg5AZdAHNDXGVlOzNDZafSJkMZjhrN
9qAXnJMpLlAXKfd32whBwJ9JQb95fgr082yyRifyrFDGbMWdv46oax997lVzYqUU
T3pTx7QSJtaClyI0vffFk39iKSd4ZAaFtSZZKxofTMZTkIpjmHOjVljay0LxZP3S
SN1sqVbnx6E6YkD+L08LLPgLXsgBzBqapUNwgr+FyXalEhZbtimFP2vkBakYO/8k
/jCGkxNigWaxh/o/9I2ZSN5DSrnSrM9vpFt/1+iLarjXiXLjmnxyf+wTyXohvkYr
pj9F5oy60L9EcDseqdOFHd60YxZldZXdb+SMEd5PNE28R2lD2nuPNhQOLqQ/Xi+q
bm97nKX7z1RjfvcinVHOk26cY1LPVWp7cTmMJDd5PxpPMemIB8aHl27uDKl03J1/
ewKiOXFtprzmcnBUray/LMufd+cAEwNkF88wz64a7hzrrzd6pk2nnngkN8yDTqKB
PaIAro8Fc6kQok7RiPaao5BSvKuFxB7fUUJ8toBOizlmULhIPpImSeBRfULAT7tE
W4lUSeO9oOMfcIJEVzpaLe//Nt7niHzQVdw9X1qkr9PQ1fjSG4EODIQuITjZK6jO
6J5EoBdAqoh3fACdyj8tvjscvit/FaAcK60m9PSZ3Na8Tt2ifwsy11WUfYcS6IAW
VdOyMwDmNA8kzZa2TL3ihNvVWgzoSpb2NrsMuYPOpnJl14M0yAIPgVsEEOPOYScB
LnxHGrobkqcRjmLTbfyKHddZSZcxJWHxA5QIaZnssLjBPb5ubhkSgjHvxERhgYVz
YMXZ61JoSAXwk4KrLHSFgfaJvci4og/OfWPi023fsCQm97v9giMxFlAz76bWKGmP
2y04beu+FC5p85RkVRxveCaP9M1oI6ahoATau88BRmOhE3eaAAlyiwTPXV99iXEy
6IXH0xh5a+4TxewwX/StS0FJHmw4EVl87wBwIFaLpWmy4a9uhigfWdhcqssFNTVB
7S2jTQVlnDC//4/E3IEE7gWgiEgQWKGUmARzjIHhd8DjfamxWD07tsAMThgy9NGH
0XGvOGi0gZrEd6Dfib3a45Q0jPYaxBf6APDGb92qfJZIDdThT+EJU5OIxAno9msK
sj5xx7PYDS1eD30J3QCTsYBm4AhET8d3wWY6d4GYmgIzdChHyol3Oxxf+JzhIDCm
MGf8tgcYwJvCOv+qz2y4P4qWn5zQ767FYlh9qAVBITVTP9FrDnWQd+lX7XMQjmAm
95Lo1kC2WHl79bvVePHRpDeXmX+636Ydppywzqqdv2YepCBCk5RJ9CKauXejLwT+
4loa9AG5yniWkD6wNVMKdEbsvel7cvqp2KouMOGQ9qQ1ng2ry9ycZWVlu5jhsBkt
uZ9JTEYkRZYyp00BWSUtyi5wdmujicbf2WDBdSVjGQoTsoypM4dcPb/amKHDEsgd
Jz+zI2UQY3RkFql6VPtGLZb2fLcP8a1SJf7eS0Gi6K7TUV//8sR4vIohau6PN8vp
xFWebRVkw575PvZZPcnGibENCXqQ4iZRXlWUOIRq3jz/XVPRKKH3DpM+aGkHDID3
j7G8h4RBTDb+HqecZXJANefxJYa54Zbj7Dx+7lceHt7TuvdB+ggQjqXTN3Jaqhtw
dJB56tfbCOgbX0/ObtFGKOH3wfkhbJ2CsaYgCgBd/9HcKR18kLBnf3pFPAm/SwNV
kbzbTjGllpoU0jBDAWeVdDUrLGuteT2b92RJ308fHTrtk+M5IAFnTa29KbqzGGZo
/oQQhZDB99v5niEAD2asaufq4Z869Xa6uJ+TbCU3/F8ISQBDOwsR0lagClb9XuYD
R+8iVZlXkROZTkjPIvJb89R2jIJu+tn1dwKjqln4aRfdsmeDG4crnwkB4uu2UDr5
q3w7D5eaEKQ0CUKZkiIiHFuvsPESmmHf6eWYxoIxvvEK9copfOSwigi2DVHU7ild
qHUbV6i9/wrl0GC98vSDLA6UYDqyyN4dLji6GKDXURBmS3DwHyo2p8i/rok0SRHR
p534YNmVl/RoIlGw8lRgt0TtT6WTEp7p9dix4THtotQqoCDIwZ6tYrpWLKyGjQfW
tPhZyxD7E2iTkstfvZG4dmQPBp2kpFbYQtlhaJwn8D2+kyn45q3dbmrPwLNDO9Md
qbyFUfanl4Xmh9vV++AeTXdH6WdAvnmMbrfXKurHNgRQCbT1SL/1PHfWOvB+zcLX
9/uuYfr6Y9ElRy5bmqulK6YPz39kBUdFAkMoZ4YWwv/MixAfvoyS7b6Gs3EWpTq/
E8KNeIk0twkSpGU5eh6szIHq/OX/a4BWyf8iElLC7Ff+059UL35V8zlL7eAFtK6p
jjeaD1V+A2avx9FJy5tGAKAFJaLKX1PZ+1YSi6omREuBQDEDJzjYQCkDm7o1Gcc8
plG2zkpd7KO1oaTziididyv1ZFzq2GP71OM7wyEoo0VYSPtXzOUigE73dm2hSTvq
rl2jqB0YSmFpD65m/ngG/kc4pVYpvPjHNdRRwfaD+OjMtEP/NlRHGRH2zhXlHA3k
ciC73L3S+QGl4DnZdbb38DZNqqAIrYvj7mK7zguvUTwniZM+1uCYruRm8JPJSUH9
32qCE9ZWlVM/SPuHeKMQMB2SNB4PFnha+AuPkJvUv5OUsBQJokw+wnnCLrPnK3Dn
0jlPfnWtG0r18S5J7RGRN7FPzUlLX9Z/VnW7KYhposE3F6kCEgBaGZXN5JN4eCZl
wQZv3ge1P9bD10XGEGVNtLB28H0gkOkXCxJ3YKq3pU8Gbb+6WYStSq4OAWuGT3I0
0T5ZZIrCDsorjErQnuLLOqW3vxlhV6mrGniNE4GVNdkBuxj/kfyxYAG0Vw9v+9lp
GELJ5gkclFt9eiqQ1uzECXG9cJavirwJi1CzkS+Pm/zraf1gtbGUCQ26vYWfcWwH
BL7zPtlM3WuGL+G6NhH/uDEefnvpu6RD3wTWmM/sXLuyKx6unYd7aJPA7pkGlZNq
2r9cSpBrzLsNqPhCWvmHNFREhTxRXW4nDkQzSM7tDqNrA/QEqjx4ecudhv1lxSGe
Ge3EfA0GCLLyF5tDLrg0rJMPBbnxyPzy15x/EUk+MFAGx8Iq+GnwQAIgiZ1pVMMZ
mobtEYpOK5xPNA+y3nT30z0UkD6QUB3R9Z7KmLVQ6PwGPp+TTH1xhcXIwuZM0oZo
7ZSEQPNm5i7Tdttlrf7qrQOnYAz7aOKCKbPdKQwYBxqgxJgxV9tRvNksp32hjGfw
o0LR3KQmAgpDkraVJvysCBH8NRzJldB5jT0W0WXnSiK8nYhkie+u93IvxAQGnE55
oRy0XHgzA1EsAVgtynVfZHgmrKA6xG9PyvEH1F0W8FAzWnIbKJBnLWwxsOuMoYxO
ezCPjcQnKP9qy8Gk6krs4x8H1ALq4oiTWZDf2/R7zr1F1UrV6DcDtMTdb7y3lwvm
EM0gFDXXZqb0BPgBg6i3OeeIt0axJlxfLLXOeA7oVDiZbjKyjzCUxLpvmyOry6Db
WMRod24m4U4j4zu+xgBun1OJqkHcs7lHVHOoiXEBRQobx7AOK7pStrTmrIpCnjWO
r2nMauURMLyH36i4E+eyZtTwwXlOBHiIcn1gXNbJk+xB15LggvOF2GMwN8MWxjy8
4Oy0HepB0OfYd+94ufLIfWymkfPM38biO1RhXm/LR/GjaGD/8NnFH52qzTviZMKD
bkeCO2We07vhu/sIjPNjSIBOi8ADm8pp2eFlzJzB/cUfls7k08t0VuXgwwBW7r6L
jwR3gFOUQAJgpYet1J+5buZkv5w59EKgydxWyOn1WdLq0TWQhemO5q7rmojHLz32
xenRqP1m9Qz4GXyZvUbIbHfvysqoRBolL5olI2/XbFTgGVWL4hLa0Bt2Xql6nvh2
kyM9H1fmiXWOMqWBD/z25m5Fo7B2dnHFecYvzBnY6kM+POfl1dPIxKycHpsnbWCT
Afezpxuk+iQz8iDdEGAFolQq80AJe67tEv4mtdCkCSuA/IWoldUkRivOFMbJzirx
euTHnt5Ag1eMdQEBPXEJcrde0p38zI5RW1XvwZz18Sp+M1GJuGS+zP22GiLb0FRW
BaubNds8EBJtyXuaLrPgiYy8w4NpgRyf3Bsq6PIo84OLRJZtWw0mmeAA8cjzXT/+
cnU2x8Hoi2rzuLJ0IadXSBPB3K5AHn14M2yJ9/8UPxKaoiV1V4mptINjBmMfFei9
+fYfHLLyRjtSng0HMwJNTpVtlAAo+rSVugnWndeoE5PCLiiRpowLdj+YYoIKqMMM
/eLL8C8X37oXti6E7gPBoo3bTAICv34CQ8fLTUTVGNWdMakz+C+unhS+x0mQAA1c
uz0ui2OKWlbi1ZF3FAqhpMS2mu4g5NWGj0Hf9pKIP7n14m1XsNWVOp5FtmdXPTjL
B5+c3/qqdU+BZm6rh4cSKySgnFqq+pej/spO+PQR/1sBJ9LwPuYwcUuHt0G1RSvE
eBuhQRyxNC6UrZSBjsw0/zPYcEfxFzr0UMv5aCy8CkiJPLtaJayITWVbLpELCx+4
0nEq87LWJLiNZe3FGHpQ/tGz39fhv3rTpW+kHt5whOo7votD5pWPZc5goq6IHepK
eukXJUrZhl4WwAJ3njVHxOUcrUjtb2M8KPc75o2REUxBS7KYTqXAnJWGfyrBRZ3G
lJ+15p+xyWUGm3fF6FGaEJbcCJVPvJQ5f2KQEwn1ZO4wHh4VYHZiEZmYkvoWpQ4j
`protect END_PROTECTED
