`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYHo3e8zW+uVXdrVqXAS442++oxcRgrUWP22Tlnb5Nvgg/2ZkHGA2eUtFgi2TNFe
mkUdoP8IYtOvCbZHSNsyzS2MUjKvezYOSSdxtcuKkYhxYAE4s/TW5T6c6+aqJ1aZ
J503C8D5mttfvar72IVwcEql7xphpA9REbVHnAxbAZeBigbAEbDD7LOLg71U35IP
O5pXwQY++0nfDaYBBtCVdAzzyPxThV+sdWdf0hL/V0cT69D9BROD5WWjpAqLR4n4
HwdkH9izgmBq3+aQD2CbmoU5/kaJvZCpqp3DkcD1WImB9Z9Q7E8YQwYevkdMvYhk
Wu60/5cmEeZAY37WnU/vJtaZeeogO87es2S1nvuU3OLkPAZctWlRluQUl7epYuQx
hEWJEH+1ti8ZLSTZ91ecQLzt29f9HjOgZ/Y441aN6rIp8svGyOv9q9/T74LymrxE
jUEGtaiUvQY0wcAa+CfM+fTpBCTblXcpUIY1gcDhc83+zn/D3dP0i4lctacyMP+I
OMhqdSu+UqCKoljk25zA7/4yx9c0FHHDuaA8O+gBJetubCcyO3/e0k6Ce7BAEq5M
ygmKSrpr/d9ngTf6F3B5hCnlpniued4T8bHhBoUDy5A1yBdz00OesS2Pb+R0cKKh
ruuR1xIx9h4ouXYaqDQ++N385FpsutNGh6ERe8QX8HSVqsuuAMua299KCHEWI1NJ
HNqJkVjKcFIl+z6Ca2WB48e3ukZp8cTkRwzqd3cNspKD48vcydZI01m+b5goffty
QfdQQdIn7eX9sGGLvKJ7hPjSjL1n4Zfxo6QHHqdHUlf+aNIeXVWsA4I+kPfZUrcL
FVcYbsTrdJScOqbJIuTRvw==
`protect END_PROTECTED
