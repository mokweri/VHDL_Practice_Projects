`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GTnqccxeed4E66+G1wr6EvVq34LHRSa+Q72M/KVblJovQNjkdfKwIAeWjmB3Hh0G
z9PJsFRtMdkwhtQI5Q3mon2zyCv3V88S2ksiIgOjoKyPwbK98U19qBvVSBTJvVio
0JrxM6cWmq0WJAPAtSCnt9TD9VxeT7M1Iy/HKGXfhV8VeqqT0JJRE6riRBeZaOt/
7iG1g6we0upZi2jh/Fz0Rrgq83xxdviHd2rRJCXps+bDUFYgQjK8gEaxqz8R2Fse
sY4yW1QUHOK0jnksch0NkJX0q8fHYpnFIhWr2jYj6cLUGZ2XXbQCRhKIZByi9jPx
LsbFZlRmczhCg/032/f0j9c8FO/uuQY7UU5guwdz4F+xqn6XnvRGAB/ukMctcT9f
Akp79Ji0WIBmrgrT6VRqgW2lNMn7myIDqsAQB0Qnj4q1ETFtXJYTn7DALpWd0dXS
RyZrXfmmrraPmMgI5IjI6fUUqA0ntC3UL6nkC9Q1uLR6jXW+3ZeDbP3eyoUwW66N
/U9tVIog3f5TXnT8YQAhf21Qt9KvbZfc79plkx0EUwugejiYBI1+NOZzHE7YXKqR
lPtUDck6kLTdKGJ1dySbdrd/LXYTe0hDb52rdPIflzOLZFX6M2vp+IxrZLIrOBs1
R0C62fuxusErTbMu/IGD3RQMCNY/B/P90guxnSu8ONmyeHc2iEEUv0d6RLzbBHpp
WFTtPpkP18v1UA1RVsSNrf4TcuGwTvU/+sdKIEMGq1AtAKfJ4JOgrJ84S2qpGR+a
izOX22J4CJlRKY0YWogknxtNAY+1zMXzhH63iQ2mePzzKz0g+Iist9ST3B0RMsYb
xEE24klKJZRGMqhSo9uEHB/o0JcD9X5Zmoop6u2pgLMgc4qk/oa0HP7mkheY3Pos
9ros3qLlfjl7QAz9LVXtkVq8OPqZTSbJWgdDFFbPzIsUH9+zLH9nWAzFSP9OD87s
alMKuDuFVry9ADZgCYsY7zPfV/RelF0RM90cbgEzBGgBFar2zqk9FQ8GVcZCC5tW
BjFhrV44RcFf6ja/VM3D0dpinuCGm1uT8vMunFDpaVAnVQZ52xyVxEfiwxyc09Pi
wj/eXdvrrHjlHyHLRB8yYbo/FiPhNI0WLVXgbebcVnOj2pnAMf2aTWIgDpbMOfSP
l1q0+YkjKzZQqMGJ03Rzc/zVG/XtqXQGVuHBh4Jv9mYXML6Hi2z6x6tUOAh8S5rd
ItEANg01hffirznq5pl++tU/Jx+mZmmSTBslAtmCi30Z8kZReBG+WfoYoDeMEsMs
1Vni9krNIAZHqqZbBWfwEYgOXIT2yCA2Odkz/RdJHTbG3eYHY93rsTKO8GJ0iS0s
hJw+hEp/ebl0dpeFdS8jM6hz7j2gC8M/qfeVusKP1cgBCCJ1yYBs2d9mR/iBA91U
S6hRSGl0A4UGM5GnYBayofo+X4UseP0dCbff6LBTcOmmD4hhdgenTMd2hZB/Fp/M
gz8bA6xmqT2bOz1Umu9MYuwCdhH8cd2LeJraKwVzXwQpdArPMrpvtv8mAoj3mJ/1
`protect END_PROTECTED
