`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLXkPkK+ORie8404/TtNMZqu7f9xOntz9u4ffIdZmL24nFzkdzoiF5OqbQPzS2Kd
lpTGnSjp5Zt2dn8+BZPrYXR0ynyAGNoPBoEeFm8fBYYsx98ckBtrpj7u69rXtOIK
rHm0upmmrDRXRHU51ZW5fxRiy41WgiJ8kYTqjw39wcIqDHrB4l8KxDm7Io5AJfW+
bAOQefELvx3CO64db6oaJ7hsxRqAPYn7oPC6DWHeXC+GNAO0dEkxCuwOtos8aZcU
6tH5k1InghscsMcXMVo9uYx7WZjzgSK4k3/hhI7Oo8MoU5VvBKTSShDuCyu3eeZU
9qvfmbV7xCiXP+sD9XMIPBRwyL7RkO/OP1auCjktcI5r2TDM98bXVkjKGRlbJYgt
+4mmh4OsWvT/2SXPC4pQ8sZVFWOX4gBHmDf1GpjwGiQgTdmuN2zPOy4fHUDa5rrN
cUdrYOalLgBv9fmsSoYulncgE22EpOsHRhVivRIgyJkQ1ci78isUaN6J9uETpY1E
9dxPvu8VjmKATlqXnn1kKeKvzKUW5Pu2iAGmU1PhJ1yTgycTNA5kvO5N2izPox2k
+bEbnUU8Ys/NQlxhziS2oYGRWCi6WH4D6keLEtCsi0DDYhuEPoJuk7mrcpbRNMfg
wCODAP/DUEFWjVkAS3fkuAYa1CdcteS3LVdWNEakLbtM5UCtoTqLfRhOlYnhvqKU
FGx+NOKUvY1GBqw7DELHqoxo6Vf/ZC2VKtLSGxPrmI180RNdMJfb2QVbqSOZ/uFo
64ur43UrViLUHhMk1H1TXqV30E7tWuUcFVlemJXob2loBz6aDD5v8mFPk0sBvy8r
OShqXrVXFcTgfjYk+gPYcISD3Ua727nckQYNb0t1srfQjSleun7G0eTmDsbiWAL7
OVY7lQT4CiCNxecq8mPe+MCs3WHoVwxb/W2X3sfMQRdayQfy5rLscGdEAligtC0J
E0q8g0H8KLI4GeRoDMiI3+paYfSGkMmOIXHJq0lPB8ujffOzME/OtaSjEzEJiGlD
fWEWIlJUoCsFZMYWN6eU41ir3zz/+xKDo6TTM4RVulfH/NrZpzemmxh4yTK7b5w6
SRXjoTRK7jM+WL7+GTw5/K4/ybWxffrdPvM7F4H75iNl/RYFI4HtN7S2GO079My0
9L8KFRsWXXkIO7pgLahGhfHRTa3HT/j7lDBBHkCSenpFxbraDzB9r0S3lx2ohyvS
0b6I0EUWh9SnDy3JQCbarqkiiEdrahRCDSZnIHcPbTonjxVp0WSDbOLuxNUZDNwV
83HAUdIuol9zOarwTaZwupy6Z7l4nAc+i9CAGxxnDxUUMvOGY8u6oYhCYRdYiUDu
6KwH7voGDLZVNTyjrfI+Qk6SOBPA5obMXL7psl94odHdMDvF/RfoluVzfVtLHy6P
b1aaKpn+LQnqNt2dRN6AYKeUhZw4M7R073jVkCxSS3USG5G21FcOpyFjkiNAr1lb
vh+qLoezPE+ll5vBtbmTh6cJc8eicVwC1XtDZHAN06AccnCpiTMFvnM4q/rx2R/c
JVMHZ8Pk0wnZT7SxEJI+utJQ9pn8XvDtUeGDgq3y+BjWpFO1bYRvm0mvtWHsE+2g
w7OYnuILb6IUmheEtYjoSPFuZAF3cmR6agYBA3EUtJmugWTxumG8839+dmfwFuCT
E7GQGtO18SnA2jY1vlN2e3rV3hHqPNJBC265nd1AokPriyQ5uZ0zNzDH1D/Xgj7e
80IQafsQW9IQoHdnXsIP55wQwRu4RpVFyrTx6zRZQ5FjPojQrzPndWg2QIG4ERCd
2PUXXTnLPoMG+M1339bDDLipBLaS9IxD3GI3ecv/G0J7dTkoc0kpvjDZndCwn8MJ
93ynKYsvTrQ9n+8UKwVQDCVqKSZN+T8rfxQrSu4kLnrfYrWhQgQU/y1exE30MCib
x7x6AcdLdqUewmlni+dVFw6O0lKYvBR8DxWDaiYoGsSjSdzvDpcCS1XY8vdAtwN1
xu9BVZMcjHZ+i4q9xLU2vh52/kYjUZElCalNMNvPPc+eIbUeucQ8CIHkWDT/FhPr
Qyi8mVdSpN43KW/wpFeo7ZVwEQykLeZ7s6nbZbudeixer7X1wKObXw1yf7VGvOW9
vHRBj+mWUzLZSTaOzZtTSOQ8HXrhbPn4YuFPNoQDcpDdXZPw5w2e1EpZpS4r2PY+
1PyomBDk4d2mB8w+fTnOj59wssyOqfepV1bbO1pmhvWHKA2fa9kmPamON9bYWZMm
kZhrBkFdzBmoQgWbIsS28Mn9vBmgc8rqCXdg+4OKxUML/RjY+Xdi/DuaZNZfn+uV
g4nqiObZNEjFSPYFknjAbZuoM3INvCEzOG2AfNh7xvg0Gz+N5cNfvHqa1NrJ9opb
aTdPdyW2H+E+xT6JylJ9OEWiBrKPok7uowLExuRV7BhmZ900iRnJES+S/gLhow2s
rhMUQvFM1CJB+jCD7yYW/hV+uGQQw+BIv426REQ4R68FT6dwJGlOv9Sl/4Z5saab
T5tTwfhRefbdrA0JbrJYgkbA6T6UcwLDBTElv6WIhvOs9m4QD1ejb8Hme4pEWr17
SD2ebkfBsKf4M33Ohx+XH2VEhUFj8VV6FMitJ0/Hv6Xx37KzhLMM1qepc/Efewpx
Ih4FhwLygh/xXz0tdx9gWrdfuacPugTL97OIqXr8G1m2eXj5FfpdasbOMbQKZyS4
oXqwMG/42HTdWJHPZ/OxngfUXdT6r/rTISgYEa07v0XombiV8Hv9uZjSc/pkGy3w
KMkUndjFMUvHN9Y01Cza9WfWrQdfOdbn/dNzErK07O4BkbBwyfm3yOEwLJY9qK6E
atVwzxT8Xv3I38lb3UQnbzu7zKtzbVujZWz3w5xWpQigP7kNUUsjWyE4M+dLKcxU
I2I9cNTQZvDVGVB7vvW6YV439CgK9gkyDtI2f1ATeDJ1taTOGQZAN4VEoc9QWFxx
z77b13NMEnj0pA4fHmOzIhIpkHdW2EP7RwHjE3IVWKPKunRzmg4LLTxsVAHmkk7b
CIXsI9rgCoP0YHq7otigoYf92Sy/LyTJuyya+ZLQ7/QOqpXbAejINE+vODp0jdu6
BC9HrEl27NOm+9UIbiE6QDGxHL7SoMev8faE8YFdZ+4CUj0kbKU6DIz5GpYKAYIl
cl7Hw5dogWMvO3NIT3g16VN67kDC4atyU9JjcFBgBk6wMHMd1BZkPLZ6BTt4EZlK
OPuq/g3RGbjiVqqEv5OfBiWSXT89Ahq9A92N4xpbW8XF98pySCv0HOEDqIV6xD1h
E1R1qCsWv4dafa/67R77uDKqYlGLyf2JVtAaP0pt2u+5RYoy+ViyVFIrpwcOkNsR
CaIXv0hOuQzEbQZzwF0RXQCVbDHCVAzTZtOBJSS7FKCFPHTYt/vJAolbZPssWm//
MkgdKVNm09xrm+R3VG5eNxkCySEGKpRWOO/LPhLJydMbTMMADkffddbWqfPW/1s6
Zi6t6vtaoxvn7Ht739nG474OxpMiBTyuFXymFXqXgjPnwGI3pC7Dt4beft4egImm
E0C7IL4nrc0X2AhZdmz2W+FDmb+v/vCvgpq9stb0eWgtQczaB5ll2HtkUC5sTgqu
i0GLSV1uKSnbZKNUYl8oa0cTcBxeapTuMqOUtJpV0ieucjTa/qXGAZDfkAtbVcqo
ctWbU/5ghdE5/jiICtcA9nil/B8J81xlMM1zF3lzRNMBIr4Ldh+iZzHPN1R8TNaS
yYe2vXW9OCXhQ33dQtyecNYirXiGQ4f+YCAgHruhVScz4JXvBKDO9jOEIELRP46z
wH00IFJpbfWUmu8WIlISOD90TrCyYDqfM1EPfRdvWdA3DpjqJUkvMIwHsQpn82lf
wPW04j7/GOdAcTc7qB6452XhRH3Oz2AHzEjoJ8GfWoJtfPZiV3lDBzI/MAxpFoKX
dwKCfynUf8MvbPxKjyfF99ncPq+SufgmSDRJgaVrEiD5rJ/kUtrJc5PIzoIKJkm5
4RPJbWPL60NvWOGq26t8+m8rSlllh0Zhh/4eKbIdw90Gr01nz2CTh5PRzOV2CuPl
j/thCwrTBRXY4YJVc1eBupOyWHRHVyXgFs+Vi37jz0HLLnOFGPuZZTdTPnf/6f8w
3FdNiCjWEOsvfcDEiXIdK8QVquVfmfEKD5dw89urYmZOXeGmBc6czLMTpk8OPE/c
Vd71wwVCd81iIX3/Tx3rvHIhUqr7Jy26lBnmm2GM/vsE5CTQugMBshbLb/HDx8Fh
+gOo8NbE2+BS3jInXTC2qOn7JlLQd2k/U+7YD4U31H1V9s5jCi47g2WThjB+DwWv
GhZaI/EXdCYE9hFHnCmEe6q6LwTeilMcW9bXkVWKZCCxD7wZ5SfdknYvw+BBbTfP
cMjEBDVtIzyLrtObROkDeeql+a1EnE/oQjWLIbntdo3YJ5Ik4CSfTPZcaFXhcgUZ
IAikQdjwTTfn1uKjbX0ylc3TsOHb8vB5/zVbihuWj286Zt6PTeg3r88nz2BrUoxh
vOtYlEUMw/RmMvs/OPEl22bw0zHzfHPwXvSkkgBWdOGaikiB76jhCxYUwxul0tno
chZYsxYSoe+7+s80ZR5ookC1bn/JaII93qRPdBlt1phAIIvWHN6TeVYkYn3tinW0
`protect END_PROTECTED
