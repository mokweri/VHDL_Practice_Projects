`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMzUrGUyqWJBTQc90I4IF2sqH5Xo9iRX2Q2idiyBQ1pb9WXWc1UrEfGCRCmSPMUL
DUH43C7mZ5v2LNLNyVSj6dES3I8zx9H7oGTnaWoAbx1C7J9sW/Mvr2T97bA+RoLm
8f0/9uSmkViEXHrA4yJMMj9OXm+0HsgndkVFlZx9baKOhqRgwhnVgh5BIpAUnMrq
eziaXibvsJsLNy1GtzUcaU1q84hc0Whi7ZoSCF8fYD8KvQmaVv2gZVxM99alqnLj
2cfqxmiFIsYOjG1fEYEBrOXqf7nNJUqfKOsHjTqRpdg64lq6xHLqVcWDrjMV2F+2
lTz7c0kaTlZSrWmSRn+E68lzaS2ispWOxXcH5V8ZkGTnq29iEPsSXLOMuOV019Zu
XMC2MgPdj2nNfy6JkZFKj57NWDdTf1tMlWk9J+FTpoz5WlHP/IBYaBGxz6Bw2q13
SuOyzQnqqhKROpWT7F84RfUpPsMT+Q0/EE0jOjTaOdg=
`protect END_PROTECTED
