`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E2ZUsiDjIDjAdHPtK2jVPa21C9IGRUSZf6qU4sRbxKDuzx6/kHQ3diy4Y4Wp7Y6W
fI54o3/ps61MBIOfVKbWmNFPbMhn+w3P6BqoVZnShXZ535DF7cjfEGksotkL+7is
K/0nEpBt8VvGel9weaVzAEIqWAtX76be2L6ngqqlyL9lJlbBT9AiWXZ99C2NJ+I7
7bSECBi/VYvf3igwqgn7j+pyxlTznPmkdq91pLJljP1B8FbxBMy92Rduv2cNYv6q
HiERC9ca8y+1z+wPs7zMBRZg81h/N/T+3t2LRD3BewImyPqPKUDDGvO/2s/VNIAE
od2a/7iPVmwh5s/yDwYaOtHgO3sDtPl+NUJtUTzM/zCa3i0BzuB74stjMZF833YU
cENnzyw+XDY+8XQ40GT03L0EXJJTCnYJpuOwg+SVuBwlhwLWgL7EHKu64nwbZ58f
GNJHzC92qL4+8oPy3mOZu5v3WH/Zt5OQCUDP6uDLUCnPUkQAwzq8ZeyPtdUlIaBn
j2WbHCEt7Y+tPAmxmryQL628M0tFyBfRycKsfrXL0njoNJ9187Y6G9gplK2YwLW7
VAupQ7DaibUbVcdCy/2V4h38bNXNVpBjlBj1jMw9XJL5w5v+Ojns8tTEH4cQ4cPs
zCVK4pTwdlVj1yhAIqMUj4XLoNhvRItkDRsbQQjqo/+k3OWaO8FnACBU0uoqhcB8
0u05IGQxwCtZKq7wpnJSEDxBZO8XXzM7b0oGhNubbvyAPfj/41V2lnGvwHjblw5d
0sl35yuRuxH+IFRRqSU7ghEV93EmY7l48rzLr2hlrnhTkkhiqivhSxD5Crc6lrLA
qaY4tU06BVMTU1fyWS3mGLXp8aPTB/x7vmaVtbO/E2HwUpuFKS9fWY655y5JbK3t
pBVc2lnXPcIAC+mKh9kWYNZejT1iYKda1hYynZry3Ot1MbzuZtFugNPI7xntl0uX
zb2w41hYecneEm4Bd+n2qobtGOyAI9PNX6D34Nii04410iC+IJJQE8DS+jMZD2NL
qEPPmLVAXCcjCH21RlgoISRrkbU3tvIinZ285eOE7J2nI1Tp5DsjzCAxIHQtLRrf
XPcLGxSTySSxsTcY2J9VllIZyTizUSg4EoWKJv0IxvdjjGrruP13w/l9AIcPg2A7
hzpsuIpVWEo1okEMb/34Pey01JmQRIO5Ri4eRK3SMrAKrTL72p2LZCdkrMYuCfa8
JVMK0EyjF5H7mPwVegNbJjkSMk3iUQTw48Na1AGcoHwdMBAFlVpTlLGGMcvXINBT
B4Ut/E4lfr3VDUtZc0t91V+xL7A/Akegpo9hjOyBq+gg5FVNaGzYOYRH2urYYx9j
JK1oNrAscuhS36JkMS5Jwg/4ZyCMc5fYSAXJWRIUVNgPkT2LvXDZwtTyIYlXE2/m
PoRwxpXzw97qd/cxpI3WIRQMuhyTJgmpKDhR2ut+z2rWt1YK+M9u+AXgLHVprNyB
CMCmNCfoAQv3jnH6yvYD2pI//TQgv9md1CqOh8foRszS/6FXofIwqNlH4rrG1DKf
p+SUQ2JyQEWRTSeMrb+8sBiDmh/mFxtDD51b/9EKI0C6AgTn8dmEpDc0uQgIZlme
e6YGMhzADOXMB5IrFYFIzru5p8ljCb4JV233Yo+5AHvzUch3KnYmDIc2TJ4FmuiF
8k+OYq2ZCYld8j8D0ZLZvmHO0AtmmcNaGniHTSlvMdixunlI5AGSyGFfEN4y/Sr6
XkMpenkXSe4raKQ+ktqQVk8iLN34vo4MINhBk6SNpEIHo5B8G6muGpU3iCHepEGs
mikrpYmLvaNQ5HRyVKPNiDqQeaqighERFhacumgTJ4PlrI3EaAsTOE+Sj7FMVpeN
aNcd99GvG2OY/WP8bNKTvg==
`protect END_PROTECTED
