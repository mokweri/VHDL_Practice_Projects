`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NuUBSgETIPSPMuJKt9ypJ6ybS/zLY2pATVKUowowMfZApewLcvcI4SY5Mbz/EX4
LYYTSSu/nPslE5ufBIfjTnFX3CBLmdCfg9u97uDcyQ9L9vAmjwmwUnDN+5Gbo8JA
PFcgMykLIFOVAUsz3m4+IwZRbxzmeU6Qebiyt2vFm8CAetGWcHKaORM3eNzmXhir
YqEVjhhVBe8fRezN5F4L2fW3NCwOWyUGC0DO4nLVff/raYlKGTVQH6W63BgFJzxu
do8/dmkZMsseBEPYy+7KtgT/QdHkEozJmMcZqJfefVBflFvHAqTdAbVcDzudgChi
ZQ4WX21XI0daJ/5OcHGuDR489qcHVXjh3Z8QNJ1y8Gdl1C3r7wWJwRHClWDrP3n9
9IuDzlwGt2EggGA6c54Ei4oD9zA0m7aUMpnT270QKB37xLtI28Rm1NNQPKkdTx0e
9KeRgRT6IHIHYNeUq4S7CfN7FpaecdPamVOfaT1OX9KUraN5OsjLAFSCslPjYNG8
S+84GwXRHNFc19bWk4fZ+Te7VYlms3sV2BmZmNE1Swp14j20XH1UmmIEhQls4woQ
CONbgUu8YWzzBlqY7wKuh0bbAHXXtOb4066d5A+DHpNdj3atIX5fj3xK01633yjK
6Iq+eVRhbZkSlKVhqTVSS/6m9y8DGpczWI4/KN/oi017mzMIHJyp+OdLzkBNWxX3
G72KRI22FZrwYEE0bC6+YyHFRIujXlxPhPPGCrHStwS/uFFyoUJg8Q7f1rPUhLw/
EE3X1Dxk+2eLxq76x2JmOQj1OEdDM3a74EgCyTxEl72posAVwQEI65Spe8dBHNkc
+Japwa/Qh++6/eBWcFQmCBRVbb27n36kemYBSv4k1viwNnRX8JHuFzG/B/OFcnnG
9b3EhZg8kmemhCfHqdXdIxRkCWyjuMZaQySd2BDrsWtHkGhGhhcAexsITiu6IK20
J2YMWI33y9YODiy7Sh+OlxdF0tF6Y8SmQUXlqw7i0CGJDP94koWDpd4G6lyGmR+Q
ZARIC6m06/dnJ9NKv/D2oP7HWXWIIY0gEo0NbSYgjKyEEDzN7yJV/nIenkXudAeK
wQh4JPsnUWOzyCD8TXJ3XgF88TeKtOcDkoqiX3HrXkCrAT304vJ+zi024+gvw0qR
11kSWPJXAhRcQXKMF4Y1V6XQE0dbGf7NHQpqWdfbHVni81my614jK7tEBVf8uZXt
NGSwgDorLBPyNwaI0EzZitS1/R8yU3WEDLYwkkaXJqAS8VU+dv27MNsog9Lf50SD
/AVNydQFJ321PkSvUdSNGL4kf5OG21KuYSA4tXX0fvSma/FLUL3jupVkf+h8lvBu
UIM9Syqb76VRKquN0MnvRcJ5qwfMshr2dlKoCWLz1lmKdFdl7f159wSFujUedWFW
cS2pB7Ls8mPPiP5AzoCsvh9aeqV3Gf9hEvci8EpMppnew2vRrXBLw7H9bO95uH8o
8P/XIRdDHJh2DVCwjjEtEUBaaWWP8Doz9Z9j0fVCJ8PvdBf+TxPGiZUMlgbRU1C7
rNi6r8mJ1pcpgtloM1nkj8ZL+0TjDo7qqAyCg79Dhs+2Cr19Ay3LCIpxvBZ6vqfX
PTkKiKeEbP4+sQntvSa/1UOUnH8Wcc9hVvXuKLgXlFSTwKdNeiz69dkgBFE66Heo
ZyeZVWMCSw21KtHcVyo0lgnukFSHUfitZmf2fTCuCQniz2xTedi90y/brlQC/xwr
VQj68/A2ke7mAum39VheWnz5yS7K2itZPHeOO+0r69tlJj+OQ+dcVYPlBfZraAkW
mjlGjpPumKQMoO0O+el2njmBcNElpXS3Egu7vkyn1zZNYp6YrYPlmi23rSYnZ2w7
U6DXQUHyCY5elwIy0oKcFohDvWvF0fXL7L/Bh8aNc921AepceamKIVPrlcikaCI4
GWFEArcngY7mIIPhwJR7Hv0ZhQgpb+SImUTl0eTzCgE=
`protect END_PROTECTED
