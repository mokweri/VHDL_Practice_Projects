`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ5oH/sJwqIs8BEE+9iyG22hXwHqrcPAztC/53bdV47O8bfBsoI6X9U74BxoG7+d
qJSkeYOPPnHixAKf+wdJbxIMgHUi/iV0Lpx6BHbFwVhalj64rGJ/UZ5vH8UVb53U
Jc/w3P6KCql7eluAop1xameMusL62F5tzZbY8HecCrahU6am6OR77A/qvWa6hpII
OJbcumGxubmpEpQ3OyN1J0QJh/i/2bmEOwKgk9UsTYf1Jdyf0OJRPk+Cs/8RCQR6
4II+PduTJO1iOdyVUGUCjAh96uJmo5oruBbnFI/rQ2J5TpGumhq2dPkJoV4QO8e6
pO3rM9+iaDSQYgc0j4rY7bxIh5yd3IkUKoNOBmr6wLHy9bB+Fjz90q1yhJKog7Q4
WNDf676w4YdeMQqAXS04xJJgewbRQRxm/WdxWYFAKce3HhCnAINiSCPyrw9WjfXv
YYi1uSyf6nYtmX+5YV3dTuS7zowXqLwCCTPqeXED8EjSJTnVT49HiykISNsX8beH
rDy4fgendM+TUxJXTKKoIiHZiInR0UdOXo4BmNH6kcyTwCAhjlWndYQo8ckhmtbk
XKhZQ3OskgMrczP2NpLuT740uP4wws2/q3AxUa1hSBWtmjrvuEYmYQ721dLLjdNL
y7Dmr/wkudue4TOjOBv4ruOPsO5S/sNqK0umf5wTZIL9ZyL4N1g7atPkPlI1x8lM
ZD6vR6z5wnInT5Vhl+2Qhebm8LQSzMVOSXrPU8buOG+W7Z7S1r15hM7RsmlORCiF
ZFlU1L3nzbwtE6CNVGV7n1lTtapju1bvmuMF52kxXYUbE1z6f3AKkBi+KLk1n7p5
OEvhEnKoF83pd94N1DG5hl/QCfzPBvvDD6ee1AFv4s6d8encCJyM0qmt1X7V3NOA
E+uicY5tc2Mbb5igupm4to7oTwj40YvXa/DWOF9sgGQpZzv1UJm1nFCSiyWaj2IJ
DSHMvAJLCxb88LjB0RKQaMyZtyrxU2Rv524JdctSyA7Hz6GL7n1w63Gkn9GFXRNG
FuTou4C624Ji/8HvTygmrIhyIjkyxUYtk5QCzKRNjdpdipD7xlZ2TFnYn5Ea5z+e
YaIhf26FPSEn/PSx5+9VMvxFodB3EeDol3yT5zX86TvKAv9GSTztvAvwgicQELwl
jSJZ4EQWIiSqP81dEiHYzQjJGADVKg19Pe4cHL3aKv+XxthTyVx25J69hk0PPka6
`protect END_PROTECTED
