`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
swHsnaI922/VrROFzxFB/sPYmN3CynUPJenPGwQb7MDFjNS9jlq5xhuDOyKJ4mQn
TG9AcSOFOx8/NPZ9up2lTc+47rn2wEnjYGRjB+m/xKyAnzzmh8G5Vgy3hqOe8eTe
4gAHkCmj5SuXPU5lKox7I1tQtVsQROoPgMElBYtjT7DVGXcxIw0O0iyF1JbwEpUt
h2BBKj2AV5J85dy28HXOU9F0+2EPaAGMobO7NhSVIP8Q/lmB1BnWerz8pbbzAKiq
JdZ3v0KhzdpNSPfVdrqCGyUhDZTkGlAtovTCu7JpY4QqY75323ls3ptSqpgLCW/n
S/x5jB93hRgz+V3hbQOyG6xzu8xVglVsW3D2FbfhyXtJS+/NPi5iVAPXbIv0Hp8k
gC6TihJ8q+i8OS2GJPOB0JJjTayro+3gMejHzUO1xsTYpn5GGw16LYnkY9LREgho
ezQJbi4IvGJNuweMHc2xMVnmeY0n8sQx21sY4litcq7YKj2RmJVfXjY4z/xSPYvq
D2CknWZB/P4eMakUKlbCdXWB/BSnxv24cMCiBbdbQ91ACI76vi+e8CBDnHquEp/n
MLJCAz615TjxsEyHcRYS42BUoUjUTKXGmgXp/UwOoi9pRoTt2I0Zv8vpVNqz9acw
c9FIh7UYfwpuvDghFlNR3OfKF5pa3DZODuyoamlUG19ZGymk09YdQNnUu6Ki0OXU
224JGyyhV1Mj8x5COioBWgEnvGIjXPpHxd0Zrl1194JIeQtw3wBk7ucrhRnC9Pj4
j3Ih0l0MvXtmzRiYmWzmFsnFQsHl6dRHRM+EGeTVCJiXCCvJDb5zUVSjIIDCT6oA
bNJ1FNfK9d1aulVlJgeRbi0w6YiMNMIl55DpjT42k6Ny8SqliIzCzIg+lTnX8QOM
hCTYccT/NQeDOyYu5gg/JJUVitE80m2/s0mqZX0DM1ueiRmwutjTf3yzGKjuNuN+
5al3OdyV/ewSonLQub0f31UWw9mJu9WkMVPsnCjNonTz0oVZwfsFoF1mgePaiUYx
39OSZ9Qt3qq65D+xunxcRWTh+7hRG2ruowzH16UnOWhJIKMbtzrAxVYOFM54sYk5
D45BLmholjspf7OAHImXPAL6d9DDMHcBbfOD6sQJ55ruu9oFqjTwz/uI57eoCPo8
Bn5pRt8dPoBW9BBDrdb0XQ+yDIDD6OKIHb3+Eq5jeXxt38lok0mYVczuYONpaUjE
NM4blgHi20IPdDLr5uE8jnM2j77W3BukN9GjS6tpHewGBY9FlamLBmtIHJ07a1gB
brrf5V8KIw9QCLBiYUfoWKDCSP+FyI4GEI1quZlZfTryjO/kI/3mgMfP+9iL8OzZ
O0gwpl0S2DFVzy9Ux+jIeuajk6cizO9bG8jmb020XTjkywRbPDDxxW9ppzTZEGPv
rtnWnKzCMNiHrSMknKCoYSDsV6p5gcOIpA3Kmn8tLdXVW1l6xsSqz42Fr38bjLfM
DuTUhMVderrFFfNhLf8Vadq6VfEwgkTcSqzy/C8dq12szHBUOMOH2K6r+jTwKbTb
BVp1jCPT3g602pA5htfTI3Uz/vWwomybHuGlMtyT7HehxsMnuNMT+SwVKQYZ4gSA
idtJ11J4Hb1ASqSNDJ3NpWNAUAy4bY+fjdexNH7TjwzmZPaU0QJvlgZcGbrtA+K1
q3Pmdbj84ZivG5i5g88/sGzXJSQpALV/+B0HmS9ONdVP+FFTjKARvq3Rku7cVZ1q
exqCIrlVREoL6xhXsp8ZBQa4ALV6l4G9vfGItEU3d5u38l5gxp6RhcYZDMnmHqLL
KoUTJ9B8DEQ1SXmHmeOrq/FjR5DUGNtqCwq5ADNQ8GKY33OFCsbkxyEB/KQejl6O
p/ZpVoH3crSbPZkECOHmdImM1vm8kRa3YyJ5aSEAoZe80XTrSkhAypKz9fieHRV9
gSGUN+cS0M4niSWoZMaDGZOAGyqe0Q9OwyNC+YN8vdv49sFQKgZJJ2hAcar0oE2K
EWyyJSPMXhnKlSv8GXS06lXWeWbtV8jdVwRoT2u1AKum3E/nw8uPMeFuvavJAfq2
zCcMKnzeCC3YcinGM2e+Funq1Fc2ft8Pqx2jdHWqT975PpUStTpHVuwkt7hezP+f
//6Gt9i/3ZNAI1VGPfVDi8QNceiVYwvkpm6b8ew/jrpXwqSPPvrVDYCrUB48cOio
ZHMSLOzExu2DcjozDTbNFj4Bme7U66KRQJEOQ9cBscwPGawYzRxcnrA777B+d3IH
py3Eug5wWCHgpmGndpYfITLH5EP2QDvyhQr5rCpNEpxb5V549GwQaNFO7v1Nfwnb
UuOsXQQvHbWTPIfZFAqMfX0MKAKf0rlotFQvdCFR6UR9X5DyimMa+3ZlcCPXqisF
m72tZykYwKpRgB+fvNgbIsnUer2oMdBGwE305B2YLEyYAE++OIunpiaUyTsI0byq
lqJl9ThuvN11/zB2+qmKxiDU3ecEPnj9LRbOeZq/AcfZceHCnbR5vdXKgeoHuKWS
+SqNzQQpDGMIPs7+6HSkOlKyFxEPoDVmi2P29qbs9O2gE4e/lliVJ9CIKIiAsRrj
S3y4ONke4xbG6MHRyWYbV4sgWO6w5XJf/+AR8U90eO3Wb9j05mutE/tgf5qbEmsm
zvALcZ2TTrOwjwfK+bcQ9O4tFFcgOzHouUFoGSWlqSBzdJVnHuiW/U8OmlJ0DRl5
JOk6j53UqZexek2SOtIVc8sbWmHT3qgUMtSPww5+WSbu3XXSbCGWTot1P9Y5dit9
6SeRNxKrBudCXhLX52QqZmU+4W2bMSa1sKR5mXnaYrnn5HyRPOburbykl9PLLOFR
SakqGQ2Lh/3aHnhLI45DapbQ2LqjwGkK6MHSoow8HMY4ED0VlD9PRXuO0GXfsuVU
bK2oltQKmW7BP//5gDutk5xaUWoOeQASUar/IAbvicNSusjbVop8f3i54/lW3drv
DsE0DWeEVyOFyjtWJYzAR1LNJl6LAs/Ea5ZkoO3ZgGiGDd8QoskhfIBAigKGIoWT
ZvJWsrDwKMcBqaRytXSeEQViKfUh74XwamQ7MbJPXPIXn6ODsNfszWV9ZH1ZJHps
Y7Im3Q4OFw0aR7Vkh8jvbvu3jTPqbnnylG1cTnOuHZzsC8xwk6ADT7k9+q568z2W
CkhK4HkZ+JnoiLlGQhKM2KKfLsi93d4qI7xpPrIQlRF2vlXvEyG9KDbOal7aFH/Y
trCVPTcROhyxFD6sNhZ/2ZBHa7pylHXSlUKkeV1SdiUDbPIv7gOouhe1QnMrobUE
GaFKYgkTNc5Ld6TZSN3GLwP/7UZ0Zg7zPK/ibALOfYd7h+7d2U9Kgnn9toZW8XQJ
2Rzl1H3CSAS9XFWW0XOEUMCUSM8vqEk/S9ma8V7zZZxoi0Fx0X2s5OJo84QQbYyy
aex51VBlcmgicbCh5PwHlDojhMSB/WgMul6fxn830K4rGPi038OOKL7SzRkMr0HD
tpI5gED87vmz1wZ67qHTg/X5c76W5K9iPCUqtbDVaZyfc1HvC/m8s8Kcz6+oitco
wSNRo92Kfmkzq2FIBaS0T90XnNnESjsgkq6U5nICxpeUDTha1jq2Oht5FgxSViKN
gRpw+aoG+yvI9Hn+hbQO/eM4QcK/7+vq/wrea4p77ocCKEveC+kptFIPoAWPfQSc
SzrDetgFtXKxR1EZ4MsK+qiCMiJ8URCJUp3DpkJKZJ3m1HhZodvAvP2wfgFNexbj
57LcO94BLbw1Vq9ZCvEcOrbaHCyPA0R8jyrZO5jJmEjSxVhNm3G6+tWwHrZ0Xypg
mqUnn8EbRG9h71WCn6aLmN1IQ4Wc4l2y0y/Rbb+UplEjSgz8V2zi6uKaDeI896d6
A+39fbIMylJUjlvM8N0Ajz/zV/YKeqN81TF+lGmLfxHX4vw7RcAu15YpnFrx/FKG
5Rw1XoewJVVhW4ziDAIm/q5XecMV6ShXiMxniKsBVZKZ0vsoetMCpGWMsN0xz6Km
6hwshEiWeGteJA4iq1QuS7WlaCww3c3ZxB+YcvfbJXPtwG6auxZhlpOujrrjDfIt
b+EljOVuSoD1NRhFk7fpTQ==
`protect END_PROTECTED
