`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+pJR8jkdVKttTQM7BQZQeqHkL6AEUEOpcJ4NdO0CLZji2xF1UdOnsZhr/y/+1xN
h6TMdDWoBGGQvIX8cifRSrnoAmRiYPoaHokaZL9dZlxTyyOfHa6Dqt2WwByDSDFj
X0v+s4FeGSEGeUvoAvPyMePteC03YOlhG3hAwksEBOhUaQXMZRZ7rm/vMuG2InMe
RjY3PSWYpSQ0R1+MVCcx+hoHsK0K9XVV29piPoG064Z2GcsopX00kkjrqmVIBw8h
xD7R78jtMwfjHeBePebK43J8nOE7MEUpURFdKb0W7I2orfUxC1xvGoAImi5OePJH
PhKKuZHm1dysOcWH/Rxk3/g3eB10QNSncyTBJ+9Eoq9qKngxRGNK8P0XwMvNYkSt
Ni8+g/PEIU9EF+ENP+DatalJ4XIQSNRrL9+s6t1P7b6B9QYoNC5v7Ax4CIJWuF69
Pm7t1k4/OWvMYdOpAmRzfpY6Bal/rCSbUjMv3aYlGMf1THnGerLhVbXA/0yeFTm4
uYjYqXVgm0vGa30pDDzycgtnibAJyMbGvdRR/3l3kr4VU02f6iI3g+eRzR110dEJ
gCtnGjsPcWzkHcxfC0TLnSUaPkNKMQBoad1DUy2ZItSGgYy+3MKvGF8p3d74MZBJ
DmMKBQ4xysHttWAS27WeUcfCpIEnsFcPiPeLbOw2eLFkV8PVPEmnJ+dXuCUqPeYM
NQBrBBrRn8aowwcIrtcYHdovokSEgHv/jPgVP0jeckxleH9FLZtXqb+IaZyiv4VM
WjJ+XrJWy9HQiSdApAsFarOD2yB/DkuvFbbT0CqChC7/aXVf8DtZOmjcevGqKyEy
JlTyDvYNz3vpLp7Z1sDeU+TqpaBJC5R45DmtCyLsk0MUiuM0GM2mUB7VjIjTdmkw
BFPpQ5gWaaLLdOq3yzaGilie+ipf1JiEcWLGXD/WVjeV8eWM3klMvPlEOQ/4FsRE
rG0QXUz0KYucq4UW8opsycOl6CLWsozp/ZEorqpTvqVPJpSaYB7V+IipBQYX1JiS
tspnukXzF/hYQJo51jtCgxJa14GaE4/jpXoFC25NHSX4tYif29IBwb99h7kVGOC7
j7VNfhJOnyYaFps7mSbPd/KYss060gYrQwYJr56xUsCUl7BZuGXPBO4HjuhaXNYq
YpcA+DkcdHApdD6RCN0OKSwamlWhQROh7EVrsTioW+Koy0yPjGI5YOn14+xyqJCn
R0vAqZhg/WiEknhXOXGiiaWBOtYImvfsK6X5Lwgq8FhZjL73QhdpMqiH4GAuFSfE
FhAcfYlZ8QW0Hh5YieeyGGHsTBLyBmMp0MZjJ50ygbcofrxKWO2wrxwaNz4d8nmV
3K7GOYYV0Er/q584rO96NpUg+L9/k/Ffa+pTF2nre7JMMpcM8kC0lvayGstMbsHf
6gWrdLUpGplUGf43fsTEBy9GIM1U1m5xxkssc/WVjWAc52vnA4QaNVvxnU3jDajY
kmebN+nebH/vReMXn7hl98D3kxm5oD3e1aCT4i7+u9aXZhCFXin1a+Po7DpRMrFP
gMsqg+01lFcpea3HTtBAPSs6LPUfXlu3sNNusIv7mNO/VHJgWsY0eHGedozB7iiW
YxWatgPl7vC0+nBWTnIbX7NbO6ZeFCkQyfzyXoM1grby8Qq8ERjVc93h/fnsr/WZ
/8NqmcQrvHhoZ5EuTMGrdfAcVm61LrIEFocTL53g8QL5bLNuxk9GSdBqO6RtL60u
ZkRzK5X2HSU6ifvG0RXhbPhsNYBBSHN0uHiEU8Ayt2pTKBMZh98U8EV52NiCNfac
DFNsIj64t+DI9sluipPRiMdyaJd93VZLnG3clNXBEigf8xzVyMBiB0dZOgnJ8agq
VZuF5A5tUFF0jqXBNSDb9nvOR+T7ZuWHZkrMWU4uuXt0RdPgCM1BGwHjFuiNF8gG
JSwcnn7rkH+vhSfZJ1rlLAvMMMBmB0xVGkp68uqTp+HutWLo9YPVmaaBRTxZC2S5
9cXvBUNtpXb73us54GzUcpvlWudaSpaZtCXtT+aUzKEY7paAuOSHGBkgjDc6VhC1
GpfzeLhX16mo+oBk/2tklBljmSvkXNZ3YXei15CSx0wTk0vwE+Oveu8qZi0b/Cbu
ZqGehwQyIXbDRlWfolLYjiDyZ2Ho55Kl+j/XyBjDQWn6wy/iyXDksMjBliqBPFVT
mQgvym7s1pNVGwZU7gN8If9BRGTXDHTd6c2keO/xlAXtgn32z+pOSL2Z9dRaAFFr
PR5vanXOlLOiAQTLYuT+c86TqOGiLherRaHHq91xv2wzCMAJoHXoaSEFO+IZn5Jq
IeJz6kslkLI60fVVned9HgZvj0ZTaqajOqHhKg4ZQOz+1hDhMi1XqEDARBcrbqQP
2y4WC3HupcC1xcimIBwzUMBAPuVGpOsPHT9XAky3lGv3zLdpzdXI6qMiNdO3eV+o
ppO/Ez64Wm1H6BQpyNmoBUyLmgYltQ1cjejqD5/917ZvETfF55AIdanB64wrh+Rg
mIDQw9Tb3wjVF4kwNeu8opj2NnTsUmTTJjJluWgQK0gD9PQYjfEFF0xVyM1T8F7m
NM+DXAH/Sgc5RpOqE80u0MYuGmSXI2ojbWarsK9PuucZ26N3hRvNzNEPRuKE7u/L
bcDOtpBDGNURqs595E01YNYLRLJRqdWf7ITCXSXobvQLUktJWieulSJfIP/raUqd
QgbDEJMN/udeU9C3D1sR+F67TJ0HXUUvtCSbgM1IsqeBv4lxWSmKVjIyd3kGr1PK
u3Rg3sd+lsCRxA/ADg1ONCEelW43oyW9fVPjqdgFBqNl34JL+SdkenmKDvEknJGe
RYFiwhgay0iJZ4FcTJmEspf8c3Ff5hngOGGjKtalSBUUueXynUn1BYwytRxHCJye
j13bn+Hy5FzJukckI/mHwktZpNUR+WQ1Ui68x06tGNXiZLQck9MoofSfcHgSUm2d
xzFO6VdRbefXeGM8f6JQn2UJEy3UXMtPJrFn7rtW+/FFpLJgz5yDGzl62gWFjOR3
H81PqqBhFY6uJUmhH+fH47F6F4qsHjvJXho5yS58q5ixXqQHVEk4VGLST5mNnYG5
jhqZwVNoJnY/kqQyTB8c0Pai6Trwpj40dyqTPBKj0huBD8icUy+4o0gFOH4s5oaG
ssh7rCtcLg5DfXrid/Jg5gIMyPy8zgLY0V8cQhqtm5AWSxDg1dcdyLrpAou+f5yL
eL1/pz6mCuvcorm4VORoP233Yjsw3HiE1YaeF0g5pjDYDMAMToZ+a1FM7V+Rv6xW
yE/sJxKXmDelPRYbdcFHHKS1t/wrQ07Vx57EFAS0a6oLEsY1QHa/pFmTxtgvONoG
L0YnKry2tr2dVxuKvSOSQwAorFT4Yfs4xphUkAxYI7hW7Iw52Yldff6Hu7TuqSxM
XXbTYPDZ9e7xnyLxu0Ba0n+GCJ0eJglPhhzxZ+hbws8rTZsSO26MTuq0rAp/p15F
PWrRdswr5NKpydACS2m7h0kcBBgfB469HRAA8vUSXj+jopQK4LSb+sxfcLGWiqWZ
EcaGUfOz1qCzcTKJSBpBdUpwdc2SVA6/nUdn2lsfZLlMN5nKB5sg4B09+znWQbHs
sQvUrQXGAE1erYSuZRd3Mf+cZBJU7hw9848r+Mzs88EkBM3yGFdFxPeYxii0RZJj
+pDRYK/eRkclBMPBqcc87/pCcEOQyP8y+S63UsVsI3UtJTWNNPzJoCcGH7TlFtTb
fA4wEXTu8RtApF1joRJbaGXSLpc5UeaninUgYFEZ6O6w+isq3i0/SnmK0SlI3qnk
UBSp3dSDM4eS1zHdTynZyM0qSqr1dMv+uXV5FhqKW3HCZ87dIMIvma5TvrcKz53I
kitdQEgnrwfAu807i8RAtCjMKGfTDmLZUjvnjPg3+7hey8cvqC4J/9z9ypuxXvC1
3oPCKdaNxhn5kML8faVk3wDE62dNgAkfXtBL+dcfVsntrODhUOjqMmbebVXv1rpt
T5JPx6W0KUenud+g40ku876bcJVx+omwpIOzwLtn5bc6wsx3uJxs/mCOcog55uRa
lnAovxBeO123Ed+JxLc6Lg2uZ9SaSgAmm9lIDYyy9l2BLAz9mIi9W1S3+3J415ko
SKttCkyF8KjtPKCLUoO1j69GjPsuF+4+ElEi0PEGUXHFJg4dX6sT1d8R2ng8bO4p
GGTntvUDPZJnUk4Ap61mhAFBAQRUrdjsbhTZ5DIjoWfi80dbkAq49m8M/M2MAxM4
T/R9bnthxuc52GZgLAWn58EauvSfm2eBzlXM6eiZvAwRVjxwuQ9yx8RhGDb2nNLq
f3DLf0EHieBMwk5PKJ3fYF7Nmz7OqA1K1SOvozBKL4Ucdlr0sX2iQAub12M3ZZbt
FKEWN3KD/T5zeYQEiQQOqGczH32MNtQKGPTnLTxqetgo4h8fZfqONAXB6tImw78T
vv5zfT54c3WM211CzIKaALXgZJgbJX2xsfJbPtjGEs/G39EaYQYTOGukZLlgULqP
YIohNVSZNyToK/LfS7UlUjalaqk6a7VPL0Q6xjdolGZy/6UQkqLdbIZNHQcyI6Kg
EatsBCRDfCVl3cDkVwrI3kv08UA6zT5/GJUSoKUepqooBdgXTqfa3zfuRDrMNsaY
UQDytbm7niWM/FxYVy4oJkQdtRKgseKDIBLoWnlZrSetedwp+dkrlXX2qu+kZU6E
E53yRN0HSUTabum9vC09/rK8Rk388A77cKN8iecb/Y4PC8yfmG6caheEnXwzSVr3
9rnOLVX/6/2Jxfba62Gc+EmSIuDnz2T2+mjP4DuibgLwKMgq0toVnTZQlTqbv75s
SUx4zweoMMD33KGjn/6hNuBG1IPzZqtSmVbnuaseb8wq41WaDuFmB7uIbsfiWqhQ
F+9J8+oMzP31oREfH2WLRO+JoINf1WRbJOcUsrIgowvktnjoPio8iicAnr5HjejT
0Rcq99dlnyVNRgGeB4dVpTJdYn/1jXnXX5T1U/NnTmzSzjFagl0IOLqKf/ktih4K
Bmatgeetbey//na3PNif5lyDs8lumrrpD6ln5lftiZpj2jm4Jl1v3bAPfS5rkzcU
sSeYoi8Ee82ayV9vvG3hJlhP/SvBexDV7fjpi+k2v7eh9fEWSGvDj3eGv7l+yXGK
0qEOPNwSHqLlcdSLwyMaVnf39IPrEbZZIeAtcajnrpwbwXRUPQSgaJzEo6yglv1B
VhgQZqIVjRb7YIxQt30s1ANhATVjZJkfU2u7jI7OsIoIp5GhSVLYn0Tg5aLUhdJh
odeRhxj3rBObe7hVCLw453tPizAVciYvzg8XKgqqgGpQAbI9/kke2VqhpKqO31Zv
zrydW325/A5XSosZIpH0iAZlhonOJKXKI85uORJhhlix1bE9qQQxzNMTu3DpeMbY
yRlFddOfQ8YuyKrqD09+yxGQcVOS+eGrwHJzZMwKhlNPv0awatUk5DEeOpzVYfKp
p4zOjT9OeQEkXAcVpAnDJaF0Qp+pJnUE/rl+a5xtGN2MtLF/fY8TtDbmfMhTkOXA
7g/lkUjQw5Rig+etUCtR57y214GTmfe5bVDIEup5M7MVxvaA9UNhHEVVoqVmUJy4
b0skP2lAGvG7hiQmz26HW+SspTzPehaVWcHDK07+pnR4Q1KmzERSclN8QVCx6vZO
evxkbRgP4TTzq5/thpGMiTqErSg/OEvITZCS6nXLxBKHdIWJ8JHvAW0eLzYqQpUE
Nmg3HwG7pPTq4DtnxFIwiCR/5g2i9yJRmQGFajq1x1xphWWaY/Gaq39ExTjk+2RY
AsLxNMs4uIqobgvxvreZYFCBiOvye/WeiKtV7bPHlUs9+rKPqS4IcUAj5aK2iHiW
ua5FK+VkN9XrtauqJ9wm6gwqtwUH/Z+biItPMxVvVSpO4eMz/a0UEwv2Umvd/LuE
3CTV7A0+6v9Og5pwhJbI+t8K/ZsBW3gyjQRj3JidSqWI5u15tue8s0CpmQiHqJwV
rqZZjlFt1VesD0qcqeW41I3bDXimnTYzsglsE6E6Coz2nRkP/g4q49qllkSJkuKK
NixZCqtjN6CzJPp7zSX2OPHstucKFihsdtGK2tj4f6ZpQ/sF5fDbDx0Rjz9nN4K5
n5m8O1bOVAv98b4gfCL8B2myM4JIjx+8AaU2y6Dtw88w3jOUIt3J7QIBUTFwmOg0
2QFycrvHqx9dS9V7fMJiwCYrEsFaVGctzsc5czGOdGSABRvxNQVn8xSpjoGlbwCe
oDi486fD7KCs+R3wt+lNt5SBr5rggM96ZmUrRZT5eb8vDKMJGJ0VTY0p6mgHT0TE
mxmGxy2SE1N5xoaOQ5wJksoXGs9ugsUtpmVB4lHwdXf3MoxJhFFtc+D8hbArbFw/
Ox5hs4zqCctCm53AZwNH+ZwiJC3eaeUQh62+xv8/aGR/Ttm0LB+epjviVxEscgsF
UEqp4gSfFEXa26qr5p24yUqpDGN0xw8uoceyM4t3qFFaFOteteY0iDSePgKo7bE9
5q3/nzlz2ZY/F/6AkC7DzOAKDM00r96uhTOAd44wOdUs36ucl+QTQiDCFsFTLiXP
YDBMpe7UdSUPoRIJQo6NbfHqOlnjyffzw5/nFSiDhO3sBpQQZLcvcwgvul7jdL2/
Pz3eHSp187p0qMJhK4kabWNHw1FLDvnc8s0bhG4VmBamwva/vxV768TQfxPj0PIO
qPWN/SUob+49HQahy8MPc6BW1PYDRAcgPDkN0BQ3e3AS3bA2XuY/MGX5kOZdGBQU
55Ol8y5pS/2E4dWt8B+KaKMMsW+bdT6737tG9DWsJlH+FLdxFSwMjZ8JOMuL4nNQ
RQVR/qSIaokSnUNvKiZL7n8KlWeVIHZCy+aSS9P73oQwJTsrQLjDpcc91C3Oe4ga
4R0snPfOECIVq9Q65RFACU2HYclsLnC+yuEwLvF+TtLM/mmSJun1g81aC1oDogBz
HWF5w5jd2oMXyCMTJ2mRlBh0jFSnvTKkYersaPgJCHNWO77Oc09B5YIodUpWzTu5
mg9PLr6hzeSSeflHgikOTrqTqs8iseYhyCWGAf+MqlUw1EkPePJENDeV0WW6lLf0
zyn0gsB9vgkTSBpQI5cGDQGQvEarFamZPhT7j0JSkhMKRGjKYTF36JMpmNE6m/K7
jxhTjUnX0G//PuPk2FXq2rDvOBnoFaIJc/pi6Y7Kd2LlT8ueU7AXHwIsjs8A2Qmw
JSRbDWb9EOY6cYLPLhthYuISZG9TqB/XMOhblLuvwloqk1r6v17dtf2X89Jf4U7X
I3y2tvnmNs7cPk3R7jGP/hmZt3ceH7A2G3cbnFYOKzZqlazWuHVaI5558b9XZW+k
lnSufFGF5zLCBGGC/k5+QwhoP8mMKKZwp1w/TyA3inDf8dBARr1HLjDn6mmW9Cg9
ODYI9sqPmSB4OvX7bo9BWJEgBMp0najLs0sVFSd5usofWmxdVyyKe0xQoBnysw4X
yb9ZFnnnHHPzheDhwZw7ZQRbvXO4ACzzxyMXmHOrrvdvzC94ncaC6uI7o9HKvPy0
2a6hR6GLRRXOlus6fjTooQlZOViS4fq9MyytWO0IEAryTFjTEQ1EtViILy2F6E82
OwHFxlNWpU4uCMMAsFKRigXKj/Z25fDu7/C1lJqKqGp0LG+juNuxWzQB5jHpDlGz
N2+IQQ+nEJh0eU/TaZ98s+uT7dTNN87Pm9xyBcNa7oT9Lx4wrIAtApZRiNOQtifa
mTkUJUehw8eaRf/CcjcMuSOEcouIv8dCoyVS+R1Id0YM1VtRdzIgJL+1F99O5X+G
Gi1a5cEAvuM0hfLL56ht1kr1j7y/UjD4jQUYXdbRTVJnKPTE9D4BX7x67/jNGBkB
fpexza+LyKAHegS5ioF0fdEXbiwMFBDEm6kXqQBsIgZz89BPI08XXCG4F3BV80sM
MqvNfVeunIy4E/Kts90+L2G6oWYF0fEGfZBOeJjot+s6JvrmjY+P8BhXov00/cHu
Se7ttNuhqlj1k391+2O0/N+W5DKVdtfACgADJGFaOBAVRM3XqW3aI/BQUBYH8S58
Y8M3OZMKe1HcGPbDudlgHwvUWGCnLW8LvUXVK/G1tH/45pj1bH9auuL7XC+55z8r
Fs3n1H/ilFbQF5bFs0DtmS3jZfLzdvlqjbVF8rZtqa1v82m0mXMTKJX/e7RMDd/E
gL8cMGhhcGttQjrEiThFqzmJwNS6humG0Y2nhXWrCXqSZkqf2W9yZdbbVskcxst5
XPTaIz/7tF0jSZVD+hMgkmPpBsxTNBQ8tqus1jvSuUeXS26FA0oe8ilVG/2EtR6a
xGVoN1RBNdCSN4vXQR51lPdq6FteUQOEr74bTlwFiE2tMwabF84dc4ky4fK1mg/u
cNxzpeP2mZhXGaENDIOfhZE90N3iso9ZGyY+ntw6H+2bbmxDXcphlYqi+RkeynWu
9ycEJuMBoVgnBJjiAvQYySCvYA7KFh45N8SYMPI8NB5pT++oah9m0dXtP9Ss+dYa
cj7ZSYEhZVAMJvxiuP48pOEe/n+ljGTopGRHjtRYbxO9T4+0rVZOSVCarhuzimN7
9QMjI2l9TfU71Z6ITParhwqfW7KWEP/PHrSo2PvO+z6lIa37iJGyq2esjVK8ixe4
ogfRt96smiJdf2TepLTI2i1qS/7iDaj/3T0/wMTm6y4jSD9JRTTSjvwnpa13l+Bc
7W8kzrMpoYNOJdKUoTKF+E7XH0QMpSbDghg6dht+Lihh1mvwQc1g9QBkON3Sk0mp
RYGgrBtrtSO9HJSvq1ioXCS6YUAeHUaAhpilw3Y2HjAIaVlxRJjoYCg3ZqUEgtdB
16Khb4I/FJSaIPXzOfigOZL8s4hdkURv0UQG7D8Xti3sefsh0PzvH9gjEWEMHirQ
kOXoR9POVcvN9mikg042bfSwNSum0wrBd8Syuo8iAmVtAbm+iLXytnwbibZR5olL
aNIxQgEVj0EEDIgQTmI3Kq2Gv8XEP9AiBieQ6FTQ2SnYj4oApbfKnNw/B4mlHfNh
qLBlc8avncfLRnEIZrWJD9b+ZSq5hiMLQ9d0j58a7NM7gZagBVpMYqr+hzBNFiAk
8kkqXPafbYjrimnkSbAue+AU67fZhk+zNFt0yYw30x9yZwhxtYA86GQbmlLVrASi
Gi3CjoMaCMzUmG85WQ5JjzzgL1yM4Cn2vDNq0nHn0GGnaUcuow4ka27gi+gxty2y
LzeGY1DE8Jg9Z1A6l0ofYZHFzZTcnyJjvkl2P0p38CCGKAfiOg62ZhxRqaGkN3P4
NHHBoWz6jlmeYTqvQjyQvyZOF3Oe5W1wlZrE2FTx86Tmz3iCBoJQLc52erwI30P7
p5gmKwjJXv5EZV6kBCAng4cAhEJh+F3a9hsVJ/gxAtPFz0NWVCku8Or64AvdoP6v
CT7jjMND8lDsMgPtRcq2m0y5RNKSBEiyvpjhf/euo33icE0dYVbHq6kNo7oq/Uo+
tGsel4mfU+1exBJaom1ijaV1TgWbtZsP3xvDo+nEkY8l92Sxrd+cNgvodxkLic9A
vgGXpWMBbhPc1azX7vtAI4wqVf0GD6EuTDPdYCkW3VxsxkTAhqik2Jvbzf7xrOqS
mffjCIYoPjc2gw2DlUc/rPFZ2dvWp0R6/+eYDw9H8DDDTUtfc78b1pkScpVrgPm/
4qZbwDnk1AOkaiMkHuBIN0pY6OWYj3XK4gCE6OR7dmd245XJRmCJ2st9eYZ753zi
9y4FErkN0pgdCWfdhSzukOF+fxvtRN6Iy6hXi1x0nuynQ3Cl1KkqFGS31xItilpO
qsGbxVihF8Z4pknVmQbDpZGQiZSXHidfGUtdeLIDsGC82ms6snGocYv+YeVF8K9v
tE1pXOxv6a0CcFhpLe/uBJmnPF7uObeavr7lFjwAxXgMJZsY9azYeO8f+DlxPGdI
RPTPiLV6yEOkGKGazClawcc3woGQlcY0dIiOq/XwgdhV/QZnb4YC+pgRxGyt8sjk
8DgUazRiVucyt5FlGoqcoj9aRAGaMcev3zD0tH5pPGxukv4vD6yKz2D2hfJEM9VH
Xwhs4C6+74BWh1KI83JsGZfIvGdQE8b6FFez+++AQcQoN26SYwvohilRbG2TPBrk
qe1NlARWp8MhGUpWsBypJ2EiCVmeGNiEUXTi3oWwG7d13Ab0IRzTuvu1AEDT12JR
UK1jeHoiUOKdWgL+urCSKQ8KT0Zyq2YU//BC24KYcSA9VKjxPCL63cyy3s0EB9Eq
i9pXJJAaAv49+AKYMxKHWwjGZ5kG7PheZUeWStyaB5e+ic3UpEFgSudoFg1jOeo4
uQ3AiINW2chAj3oZxslKjWvxFJ8IKh8JjPlF3YASjvwCIb1QaETokPQe8sWwJJjV
4+xWhcxM+AaVI4WS1FHwriSpt3hLa77LgaRZkqZGqwrFSN5EGhvJFcBB3wY06Aj4
xcTpoOpSByUvpdSXhQcmVVTAa2zqnwzoOIBI7XiZb6oB4fRULqYnZibx5mV26pJP
+gzjKeFE6oaxlxoHM35LmTN4cgIp82NVGvF+80fRjgGatkwlML95mbg8TYD06CVs
LFIrgLsRc8Fh36/wMdWpeMsjs/nqrbi+RDwxMUwCoUN2mUCqShRN4zbnwuJ5hRm8
SFehmIzMUBpHgGyOOT/sBAz/WFT8HRF29GCjmWKxQx087NklryLvaW7bXmZCZVD/
OoQtZvUBQ8nu7ECmd5CWttfxmLDf+BvJ8uki2/aNHycbILVbyVsq+UgDIQEzvsfK
pm4hKdnChA1pAKjfgQVRWChRjHnOuE9lOZUaBRQt8ysNCZl3KxLRuIuUPo/YYFTv
j0FC3TAB0rMg0sK2xTUgGtW1Dg+nKpaCmUhOr4a/B4GGc21Yl2Eo+9sGvgDX8gg1
IgjmZlxaXYnBZ8/0dKQJC5mAnbuHloUjsFaiqyVa9nNUhn2pfpbFZbQ4hu9+0yjM
4ZogwNp+s+mB8G6sdWewDftbDyUHp2q4z0xfYeV3j1RUTzzSqT+I5AmO87kHrtk3
KvdJmR1EfMrs400D+CN6qgpozqor0BR9IxzgN4r99W3mqsWlO1e/F5X3eRuXNzyV
4DiGiO7YZX36v9KgY+lLlGO3DBDa6IZTjNmHXbQ+hWK7VXbXnvpaBNYKInUB382I
LsJ24LjgkPb8uZrkGPOavNdkxS0I7YjEo0wXGLD33T1Ld/15umI5M7MXCiBOhi2w
j3facPtoJcvzEIZMdBS+rgq96Yo3ti3R1PSlmPuuuG8S6Y4+zqBNLS7KB8aIsBQZ
Rtw6PubMH7XpaGDG0ZR2gJnU/YTC3X1/BLQv9MhybPuMib1KwINaAey4YOBvtjHU
D1UKB0QXzbz0IZBnT3stWIxlcJI7cbkCIWXSAr0fceP4vLr3mwnZ/49axDMj9HcI
eSpdfsVTjkDlJ3B2ZrPc0YW22TR9HHETpdxfYx4tc9yZYdPjuMhy3RYBzIqvfdQd
87akDs1sNfxzPPAQ5BS3g7bZjUUuk8C0Gtn990z9SRSukkj+CaMzYXsURqKrGFiW
nBt0qgZjvz5ctbf15HCUG8lnVHLoS9ar/c84m/QUCo+iJo6aNLb4u33EG8Z5UG1K
iFSdPeQE2CNdCBwUgC8WgH1O+lbmn0ocslEerBrhkWBb0e1k8iC62/fVjCfbeOB5
/ehjIDxs+lBDINaxD/+DaWPH+4MjJ8/+4NGkTzmWTSDBbcQ0QqpTS0lnBJaLDOMe
p+txFOmu5NssJit7itfyZO1xqM7cxCI72La2YXdgeQfV900i2zPts6g5WdTYzU5W
pa8rsDxC4+k6hF/gAD2BKrzYYt+isEzI4XAhakqLRo3QnMagVuUD+T3Gni38ArAf
Rj8CPoQilA2GufUuoHjSliB0WzwlCseyvqQXnRMubdhY14qg+eVCa3vm582riCvo
r+eStZKg40l8kCZ3e26M+8loclJYWNoDsajwFk5/HTzaxkVP7X8b8QWZHIh/D2PM
DAJ9ea35FBGOpyMPdQ65r4Jl34CmeEVU1ImF0lpzCbOu++mVFAmAuKXyo6c6IDBi
EV+32i32RmD7TRUnL4u1sq0jIEFohfL08SgPv2eTlJlbUuIuHv2Qj1E3QIY4TTLy
j2Pa42vh5K6j/vBPDe6JZ+8VFait6Qy/l6dH/dkGWSt3Lg3AsVypr2sRLJAxgB/D
SZumP6ThwRREB/cA+bXNLGeR2mqhM4qjLyq+ZBAOSWhh5md+O24TkgLjlZGMLStY
CkkQxmqEkWJiCbadA+fdXgWmBetw3xz+pyT7XK/fgX0VqRWaChmJSjUMvzJRsRse
aWvpG9VMjZ3yD1Q35eRmKeMCw+enmXP57AkILVaSsnecMyg9lIHqCkCOTuR2I8YW
EJUFBz5iJ+S4dGLhil47U+Zst7WIIuxSGKg8vVFUkRqP2NXtEVraiUK4pwqV7rXZ
h8xvdkjMoOVOo0tMjA2+PH+kXFcTWTPlbZym9Yugcq1rf4MxKZIJqdtW9ZbSpwqC
iG/is5Kdy+iyIkH5f44W2/r1QzXcBscbwEVQs+zwt4CiU39EwWMW8+2MqAIIWza0
fHfFnG+loAHAStQ1B7BMCxQYjQQieeeLtM8G+0as32CXOjWt1/wKdi1IUReHlfD9
lDcjcOsjddWe3/vcU6hYI35sEsDlTTTgDey9mSoBsFq6ToiSPYd2xosTfHQySm9h
GKu4pEDP0EKABWuZ9regP+PWjHzcL4tvyYklEpHaJHX1ppIN4ju7xLknHH34k7p7
FhFmdIzmi51q/12eS4KHyb8Eq4J6LMroGocHLPw2+JL0LGAihmhQQDrXGbtv5fBK
yZirdoVEsXJfwdOR3YogsQozy4K1sZKRWg77CypbIh/1zdzyKXOGeSa8DdcKrtBu
3c6cQaa5l6yOT7gBaWlCZ2ydroh1TFhhbiYABIxJEg+V3igi6GYu6gxa7yZVdu6j
w07fhV6pp7UJmOG119p6ZampoV5ws8YAzB1VHdX+o25loVXZv/ewMMIvsemffYRx
K9ypKMbg/SWb2YJhjHrRYdUTQPDymA2SyaKTyOeeyXwftXMjG1ODT5zJz46lcnKB
bFGearcUGB+L2+pXM7jLXPBl+mgGSwIGD0hfC6vjxhECDw4rPbK7ZVpyDwYUSa4v
4qTFpCP70RfFOGywYbP7yfwsUYblCDiOufr05PPJ283O/6xogHI64U1jJPdl2cke
/+6lG0yqmwEkPVi+JExO2THuYTlQ1O5SmQvbS+xnA39eJOqeAepLHH2PWFdO0c+j
4WDzoCNyTkqC+7qjnITfxbkgnUrKIUa0COSegcO/msLBOb2vJgCuPCnYIA+TySW0
p5DG5WTKuYmTZWg1NQMI86VjqIjQDKuS6h2Ptsb7X4qqsoZBy456V9FqLbuGzQlb
eE1sFpR/5FefJTCMLOF444ziQxa3E57WdS2YM+Wen8OJtaJiXAo52PIfhKA59eOo
YqGnuMZkwOKYvlNQ3aZlGqHa9m74B1nA8iBbHhwTEdtodZ+dPZUPs4abZ6O/49Bm
P+9QquzWORYQYXkkg/Rm7f4aothvQOuhDsTBw1k0oTKcx9Zr4On7CQk+q/otz2tM
Xg+T6osKpOd0Pwy6j/k3MyCCElNxW7jwRwzdxTmr7BdknGR70i/JCr/r1k4TNtuo
St3niAghkOgJiRpi14UKSm1vKmskgMlOCJLNzTGrXhDCGFsqlte4/is5FSY2lm37
c9toQ2OFFRo+pQvXUwFuPzr4sC95HGaeu8rPZtfA8mYjoN1pSQxQfbqiaRoPoYcI
YGoLm9iL1MOhMZfc03cbdKRLm43TY85gBsNxpACH598IDEKNTgEERtCjqijAtnz0
XjqL2KvZ7lZn0wF0oYzqmDlVPBKSAPvByYtzRlBffiqWyO4qgr+yFwN5PaSSiC7a
4xxjX5zRSA2SHLX59Vwn4gDXturpAdeNED6dlfBUyZSchkjTIiTyeWmJFX7obNWd
9++RtV8dzBfKfDp6I116bNUnzr+C3LfOX7tNWz10Sg+wYV5bzKHQ6QnIKo8gJSb6
ekSvhKioaie1uQYYdgrWK8YR8vnE8xivWlvgwOnpqOjGVLeYAEka1nbniPGgQeCV
PuI2OweNk6TI0WOwODGN+450q7ecSTWxgfi5wy0vppx7bZWCqMdUwIlorrpjMpGm
t11djt8bdcntsTV8I4Ptw2K7PsOc9k5fntNQvYBvzzd4jVgvySpy3e6WCH97jZyY
MhXghDWkRQOZCD2h4jvQa4/LPjz5cAcimIF7i6JmRjkq/8pi59yM5JBDG163sHDT
C8mKelzqWavizmcYLHBwiZUPn7VOHumwgY0f+P+uKqyKA6U/7GS1Gg39dVhyxxU8
sTZKm8ABBvrBGXRRWX6oov84W7T0CxXLFloxGNzD2mmSCEB5u6m295G3Ssx5iW+t
yPZVD9uf8KCXv1vsb+V8QdnoqwpAe6Keoj7ptRhOosIlIz+DbtE+i0HOT7XFt398
RvHqOxuIl0ohqvvVGmdJRWlWwzfLijalzBuslJK7g+KqJEkm/MviF9uiQTIKIQxZ
3GFJxnrfgzUptDjssttpqCM0l+5KOijoFOG971zAEsBcamcfAHL2PwtJfvSMA8KN
NMXg1M2HPtUCfClMNXLaSFUtsYII2JXTvlKG1cO+GY1twQrMwkXanU3CUw/baKZu
sNQqi3eAp7obGIt276H86U06HrDaxUUR++eMmJPtBUnx0AetTaHIjJoPAz8F82an
BwJEpeAc3Q4h8fqcFdDPXgDHP9VV07jStF3l2eQeunNh3LgyVIl8UXTDM5MEJo9H
SM5FEzEBZ6KTK2QPOf1J7UDbn2rCptFsUgNK7O+w67AUQ2au5BYXauCyeirXS5JO
VfBlDFms13lNoRpA5bcuL3ejhsAyyC5w3DABqGQWWd5QC9lGoeBc3fLMPsx8zOO7
lFs896rCB34RtM/bi1ttH+62NChMfAa4gerBYUd1towiM3HBVVSWMaOUgLOAZGbt
EQhed4sRCG6yv92tqm+fMZBvJ8pQNHYXvT7wQ0n6obefGON+vxkBhqkVErrx6XZd
LcuaCWfl4gmY7iI/61EwCzy9Gzyc6820B4z4bt01AhOffYyUt64bJPdEw/E2aj+M
Urd87FhrG5NOtzIG31dw8eNtb5IrllkIx7GEuRwim2/sGu7p67EwDvpDviMGfDpp
yP1vKLvREfDRQYh010X181+huhXqaFeyG6KD7SwvNeCvNTDEKHZ/jqEMR1+X+lfp
/pZPtjAC5xC3ZYweUMdwdhnjm84j10aCBt/MpAXrv8LEQXerTjald7qR89qxEamO
mlzy85GYbd8C/WLwK3M8iOmrNUmq+YimLJqdkNvKcFPM8emxUXQMVIej8onGwYYk
EiMknZNyRxsHpb++EH3NXq9JWREVw2VjgvE0ChO/vdxplF/UYGT//xwZGQhnd2PF
dAOKl097qvRZ3VwPNvwhzP6ad9DeXao/xBlVA2jhEcFEURVr1p/gjtcfAbfeh98p
v2m0Jbr2c8rf9ouotJIH+BYDP4Zk+zGzQksos65JBIe5enSW+v+UTO1+RZ55ax4c
0P6Xc1rO45Gs1ha8JK5e52RV0PZDOyemjmjb+bl7C9EatKcliHdygpA0jzv9lOuB
CCWdJOv/TPpDSQxBLrR2z+ZCl6+N/TX4hr0Ep8pTwwFLn8Wm2bV5wpr342rKkiiM
4neVO0A2Ov8sJ9+qu9q3S4Hnj2wFWDNTQsHpPtQReJ5oE7u/Ptl2ACGY522UZzq4
U8BnEQYLmp9pzxU3ekHXKkCOlFwX+4XgPZY7AtNBvF1dDj80pggvMDIH7qrZWMkM
/kepOVDBcLuRtCuDK1IWgU4FQv0XqJ2DE2nJYZLQDGGWLis9i6D4q4o+3QD9iNNP
wMPzVy1fqixJ/hNVUCE/Z6klOIX0SDmsUWz1ZFj0rriE6XAw0Rm9dtTzaBJMEkAO
feDxlgcWAoBbjUTufs1TNylPeE+HXS8UGA37/rPxp+wko6loY1dxbjBVitiw1ZnP
8KL3gxhtcfK56u1jS0y+vWKY+X0ceGYLLrqY78UHAqZGI57eFoRwRHGyvEXz944p
s+YrMT+tIKCTsuLxc12cApYWqh5Eg76DNlVNaEvvw0lWJc92llD8A2CPlxgZj8i5
U7UBpOWbdl2v6lgO9w+YfdIvgI1V4mXi9YXN6JOn069VwVBsAmYadZzbHhn9cxoa
woAdr4kr5MsU97odtmKbhMHMCRD+bq15L04xR+B/MeHKZklXpJRZMwbooMa7C09x
RvxonHV3+7TVDcYPMZ0E5h2hyVHAQAd6ccQEc63b4dh5MRyuyZd4MSLgvgL+4L+N
wGDBgspr/qq1dNWrxSibTEsHFYcYPWSYx8No51Njo79WYDmPjnG/lnFc2+Vp1N3Y
Iqya5i5Fx3QUGss3UusvQvAgw/PUGVVUF3xIogEeIrof4VZFRGsSokWHD2kioT8Q
61wpbiERhl9z5CumOBolJLOkHQiGRnfTYqJUjB04Qss2r6Sxp7IpRAQSKyz43OVV
we5iN2mJX+lfBWRwBtHlABGw09wzkil4FuinpGSKICeRRTK1/vXyR0a/HqAJaJ00
d0LZLRaJ0KUUo3+CAMdQ83/zi7RdxL+Xl0XlI26sMK4WX0YqBet6ToV/VT2Q9jHn
uSL6LFxZEw8r9h/Cd4eGNua49fte9cFNaKHPYzWoi2fQZRBsdcSP12+wj7k73HfV
V0R8SItuNcsS8rjRAai4LQZ1zFlpgBNNq7MxMXyjM0K+MAgtsOlW26JkbB+ovFn/
mRyGbwY0w2Y6/UefaXNhk/QaEe0ovRToeL3GITJQCLPyoqUQk5htDAhIokdViDKA
murw3Ky0hj23Fg90Tz93f2AVtrm4y2k38XoH+GM4wI0QTh4A24UJktpdtowP4Y28
+dJfUlmT+P25Ju1Tw607gOSoO6s8GsfIPUfhOh8WEhSwO6VrTHInYYquIv6IqVK+
RCzUR4bdiJasV0dNoh+Fj8apqihMoXJuWzXdp2IIk0nNVy3+/GUYuoVTehGQwizz
PLlrKtMFST8uDzGclAuNRi4NzTvGfvITdSoFKUIvqEBMa4iiK7T5piCL75MmwYMO
qP2PR/ts3R0EPH1vonMhHSi11pa+zfWUrNmgNGlP0GG7EeMg+J+/QGn2umgWgMXm
LOnmWJNJsTJ1gX00T60kAlhKlKXRT+6PMIt32zp6hgV9Xze2jPWHFEZbJT24QDKl
ixVmSlpRi3tedeG0zckWZr6c2sFt9rfa+miwPICYLIcTmHow8IpaQtDKmx9UOL14
txaanlnkooRdbTupc4ZlbFhVHs0ljRzMIWx0Cow52Wfglb7f1uOcnVl8Wl7yr0bA
jCCmPcSO+khz6HXDMsQdqLWbU8pmBFeq8+NmkG7/akRJMhDNNVxsNqpBLxEWqaKG
nuj10fr9Lv+HAy+G4zjnj4lau41K/f6fXP3by99dZVJIl4BqgL9+ajxdvkpHa0ZM
HbnnAQ8Rdj9DowEpwrED/yuonA0lF9hQJhtaiQzDQN8Bb3wONlIyIiHwvHBZ0qEt
v1DS/p2G1JrHk9tDtcDMUxKu/CTn2jwhCYKA79DKZLyZykzHnUAFjsxXo/XY0uMO
DWZovckPoPLnFqQAcmM7CRvsUTPGpryKGpyDUtQddqWvuepivgGi1BsMEixLjR2N
NT7zCoUB2qRrv2+3idmsn5xCtcOaUFucWYcCpHNOU8ipAdwrVxNY4f199rztYJ2j
0F8IRMduLQ2CD5dxlrvYQdSqk8Exk2w0dJEfQ+9nySmUqpaa+T6Iv5f5yHSMGE1q
WZMudfBgkJJ2r0lB7z1QcJFF9Wn+4YrIVtE1gtQR5V/3LzRy1lz6x/IAv1C3UQkb
2YPB4ysYP/MILEcWyvAP9eGSOqYuEEvMfWi4m5waAHm9fayQ4Qw7LeOGoGYbGUAV
LUc91TgVCEBijpWrXgYEeU85r9izYqajF+ECTrt4F+olVvdOsKnDPoxhH7vCW4mO
kiUre+I/6MHwwBF/wtZ+yeNfn/0gjayRrpMAfEqXEad+Q0sec+eA+9FFjJ1xLa9G
h75WYL00L/8SNJJBHuxzSGeEDv0V8DwicRuYymF+IFoqSpywwJgLeGa/bwRhU0Vt
j03H+HR3F0G8lNaRa7PofNOlNXocJBIzFaGTl3uWBGzhhn+hk7/enmB1fK5wI1d6
em6aK4PY04wpGmHBW6R0WxMbapuq2SVXjn1WDcwl9AqXSfXo710LkJr6gR/Qb2cK
H+4EoktA9ItVWP0NOUiin1Eu2SvR1cV30ywwYwwYBDuVZxvV74RtDHGjE9V9rhuP
Gsrq6hLsBuKRJMx5Obupb6CzRswKT9tGUcGvqb6uaDzHnDSR3cHecVi6EvAfWXmw
ImkZH5k6PgmqMG5obhF+IBFnn5Xfy0PFLIEGMW5srWMqhHG017KPtqyMZ+D98mHU
tGkIUuTUnbCZzDqv48/YeOi2kdyXuGGLImUyheE5ajSOHIch+Zbw7lZc5J3AvFko
LZ585+BgVZl9sBlMiu/XeM1o/p56NhBxQxuoahKO3q669LnlqxCUDTji23b4tHDg
U9buxK/q09V8n120ONjq2V5P/PcPzYyDu9ZlVUxJBimSulvkQcIX97PEarJV9+Gk
jKi1zpy4iYtyRjmDEbfLEQljW7wLzlF1nQrroSZo5KBG/gFFkZh/+qzPW7kx5BDC
WpwOHinWBDAq5jX+YZjcNhy4ivSzo6eUJSsrP14OVNIk/uzmAH17kpUma7DiCJBL
88Wj9yDVGb+HYRE8krALMLLKJm7ccBimn4wCVN1Alf3K3/sTNSl3xAHyiUTL2aLV
P+nHDWHC9oN4Cmppc6rgeOTg8rlOWABMy25Ekmvobi2ztti5naUHAOu5qtvNebJP
R0EZb3dwIEhLDS4yJ/dgL7dMTrayKEJHVax5EQJqC/+/15y+D0hd8FjR9k775kNH
Fm5j4HVIFTrvxltTn4H57Msdxz4KH2trUq22VxJjMoDndCXVAoXPnBKa03e0sNjR
GUXTSBgaH+c0pGvpGLPOS6Bb1CMNmpoQhaoqhDyK7I5d5MYElP8dfRwlq4YA9E3E
W/63PbN3boEsK5kXZdSQGZRsyf0YQOSJKAwCkA1nYUBpbrfr0tNg2wiQAtIjeqhF
OnWLhID9xctMkUkQQxxdgzp1KQfMPpLOd9wVs+sySL/xhW9hsoGYCY3xip/xQ1HV
jlpQxF9MUH2qexb4wazAimbjm4GX2v61a8GP6R7eF8GchHYnZ25aNeG1swyD0mGM
NaySUnRSuETuqrReZucE0TMJguPCafr8ZIb6PIDeZhwNCadSRvj/9MOShnUYjrCv
qkW7arLfDlxGquzwvaB3Oz0GnGzlFekHkVFzdFcAIYMKr0F0R2H8pOH/dnIbqkaz
MsfJP3IOgFh+VcN8osBz7gBmD8GQ5YsVORHKYMPjddPhvrfSS8QYPB1ZiBInQW9J
dLzk/ALPIQVMBXPiaksv6nORY3o69+9juDBk2/UR31jpLaJA2e25/jPtMJOqMcNP
ovQSEv6qw7PlUx01B+vstQ69sJxgkb6d3lZ+K83MLjnEGITOMoD/L/MPYbJV028D
MxcWfjYr6CY6ntyLs1a48bxVzajbJB3YOAWf0z1tlgZhEH0vAYMdbWE+t+5ikHX1
LNaCBsZyYOH93bs+0f3Jla24r+5odC95qNMScrIGI7x08zJEVAlb1IkKLYGoLri7
Qu0ybUSB0I9AkBUw59SLztEtBHxt6B47BZMGR0yySHh+gemSF92psBvMXkF9fNM+
qIFNyQOoTmEIDT63lIYypVkg09Z3Xk1+4DBsLSrEIwwfHmJD39ptkDaPph428fnj
BzNyiyLxe2X4DPS+x5aamtKzSn5Q4Mt6KSL3Hl8yLYK6K/7BweFLpla6a/iYtfTM
to+Php18onDFGl0YX6nsn/RLZFN8cxfXRhaNos9LZ/isGK5XgVKZitBS3C7+AjfD
Devb/tWDUnFvE3Y0uKMqrEcect+lxOwHGuUNNCpQNbrd9GFat00MJwWNkorbDs/P
FyCyyPeauS0b8VVQfHx20HEKED2NZO97oaTpkEIuhgKhzz+MtsSovd0h2XJHQ7Qc
V6oZcIWVkpW78gFEGLLU6lnVKxrGPcyCaumvUieUKlX8TrhIawuMGpbtsWc3ij7m
HcHyp2NfkUAsppdBpr68iHYs//tYPUizBdmXi2OcxFrJoIzhf+gKb3IoJQ5pp4a5
iaS7dHhpVpk10fB0Au7my00b9liVsfo6FYMksgJY2CG8fg48Tao6FOdZoxCaQSEq
1OrNapza5frRr5VFGGx8RaY8eca4OhGVjx4Pz1pMX8p20STvr/cFXwxKdnerg3eE
uvAiPjgvovo1tXIodPMGzyLc7s8FWpzYnm00c5UR5zAwwZAm/7zAu0EItr/37MKT
OstVZI5/UW9LFMNmYZGK9cZLhE8YsGNvthV4OIXKVx/0Y8+xlJPQvo/mloH6xlIw
J/WTktPAKfj1WiwSGA1SwOJnH65rzWANLK3iWOcCXOgQ55gvzMRYow78JjaH3HHF
2gYv6hT6ZvVhSXjId2j9gVUzGcb8W6eQ0xdHo9YuyReb6gZS1Lp7KM7f0fBNrxpG
XFu7c8IwbREX6IbW1Z0bXFMPcak9fcdAHVm6H9r+sZgIAvx8zbYJfEZdP/p39VEw
UlMeB14xZ4X1+G8sB43h0GCdvC5cE7O6nuA31BG4IvcI9sh+FuziyX0DbPT9Nked
yvLptXt+htFniNAlhdkp4gLAYyjpG3qnQA/w1rxghe6rzaDI9+etlA038K7JVTYd
bwGsG176pS3XO+s1yxqlOmZW7ay7wlIFyfw7H8jcfHBxe14OU6UL05iczRNVcg57
W9Jfg/xJ3TSywQrACFgdoJpzEn20NiWHq28LQ/UbIktJSGIlQMwTtNjsSgiM9jrN
wYu3wUxJ9DD6nZQM0jZ2ZsHoDTYMTOY9IpjIWMHQjld1PW/v8JdZ7BPg9MhobmMu
NinxlcwXylyTeAIITgG4xOdIvnLmhJyWFh1y4J1sD/myMT2/Z1LjPfK/BNAU7g+D
Oct7nPW1csmrb87oaKTzsDyqr33gCqKWEOmhtS6Va/Y8AZsLobXzK5B4yWtEcUDk
yvsBnymCDXwrPyG5KPH9HbnF3DjJBPD1SDBvtnb6sE8WuMgEf2N9KiCT442g/Hye
K08Y8Or+aP8IZGSLSa7y/tD64GjewnfvLUlUNHMeR7Dg8vz8UUeAsNdegaTSnMg9
axYrN97+boSWej1WlU1EsQqAA9UvQJ+Wa2TFPVXOQOm0YcBX9ANbJEmT4gDm4QBM
HEntK5tBzKWpXx7E7AomC6kpqRBiS1pGWpIufbLTAd38HGhWKZYBN7yY11migIw1
JhQftwEC6xfBRUBrL3ybJr1DkP3BkMoo8bc3jPzMqf7akAt08QQQbQVrq9lkfkNc
xH6qwWT0cB34laDWeqwdserH9CUYyC1rYkT9SRNiinQ39/br281tkjCiBW8Wh6N3
NkgT7cedo7ar/3viRhfUUe4RQDExwayRcNm3niD1lWE67HlNMyFtcaNjL1NXqqQ4
kuy9oWXdWLKcrbus0Cl6TyVmLlX3c2NqyH3XRmJQwJvBo4tR6Jktguvl/wW5Z9b9
cucF0viZC2BoUf22PrGpbILedPUhGjqnh3ZprmzzrrzvjBmElnOQLuznPSESV40I
ZNsFtIdzNyLe4iCGu4cS22eTfrl+qlxwpgOorYwfxMlXULRpb3BbxUEHfpqHb7EI
fXolvg7HVUQXf9mwmSRCyt/MrIkjmfjC0al0WnW2V6tuXDD4QkufRsG9eN9xlKvO
EAxKZBKbz4rSzNrrPxPZ4CdYaZ0pGFrm2PN8mBSgqNy4iKn0XQvpx8LEj4DoEMFt
ls4QX3P2FaJ7dZtkPUoHtp0eCncBjfc4tdQCds9z5EBenQLzEvXPYIx3PFlrKHDl
zDpJOM2VgKTMlMnp1fMdCFVo+MULjcaB3JioOWAMUPpvlGJBOg2l4uJIWnCOlxab
05Ww1n+IuMkQsQPpmuWBf9MmQ5JwQ90EQDUqRNfqfSziIxW6dv3vnY6jQRzNcb5Z
AoQC0avK7gP1gf8Gr3VAuur3vjqDsxDtIAVAR7xevVj1a+WdofDAENg/g9anV6Ke
8Y9VYsOFTpvHKO6InR2W1M9AlSDL9WRbLqvG7Wz0QhHvnErchoYqEvPY5p47wo0w
Ya+xKdEH9/pLHbLbxa4dMuBRaTMmZn75WYs5lswfEFLCd1j009iJbEfvLzMzyAGo
tlTBtLy2enaBX69YjMzEXNSis79SrPtub6sM4nOMH7LJHz2rkqp+3z3Yxw/eygPM
F5pvwiVhuL92S+1ofu14y/VA7X8QBrRy59+RhMHfo4SNwQ0AzqJUwVTu8Wq8aw1d
Me2WcERuF5DxbSkD8+3pJz27E3ZdGRlbXhTL0iPpYdXSbMlFiOcWDTbw2Wbe322g
vvTWR/2hZ1vHDzTdJTUmlRnQDXFnBAbXOQFfP4vKNw6qwERuXHVtIXZR8g4hTvjd
4yGoKs1HsZcVvakviop9P9v3kYMcmXPC7c04lY1A5aoK06zGlZL21a56tcha2mgt
VFROPqno6rnTSjbNbQSHgIk4kTEmoeOahn2MSEYughC3umm5AEpfeQ2wuA+K14NU
chOqcpHGmzIkXKrWGQ7DDu+FCo6/ICbhmdpFSTNpo1O9qJci51I0EC/mBLd+ZTU8
E6f77wIAEHd9S46TNRgzJNyA2PyBkE9zQJatVvYSRD23Dv8WcnL6+0HOAj3d5zZO
S9Is6ZIKJFNYBV3p8wLaS4+AbGfrDH8DExBaSVB16QlqC/dKGdcont7LclGTfwQ3
kF8rbITwO5ShMzVKMUMRf45d+u+NsUcYBthTG2p7DY0j5/tphg/INFaKV68HpE2R
wUfdFlmJEmzhxHheWYWp9VEibN3IFQINo4QkzNu0+9ouPWpzr62avyDGPoAsncti
ACNaza6aTwSxCl6EIkR1jvIWFUWW/SpUhn1ic61549xuhtbBjl0/6ji6jF+wlC6l
4F93nbzHSFH+6FKENEXLSgyhl4bv5GCB5O4OQey1aakgDEysLnnfqPMTnOJgDwwL
D0qHz0BPiXJnpEVxmaeVodvdR+zEHIzh13qO6Fphlo3X3946d5sP3PIBhTmzxwUx
V6H7tHFusITJhD0nN7n5bWMNALPwzUPeTcIhnIdlrNT50dt3/hycGSC5ThhZDkbB
R0bEmvuoFdqmMRloFA6HXDnTR8DxSjFvvn72VTXZxosaXovl+FrloAEQkx0Jch3k
vzKcHjxXmrmkAtLeL/XvN+fPllQoErY6lNpwEyj2ue4QbCPODCqYyR0pINWfeq2U
WtuhTNvEqMZ3HuWQxwV+t4BG3uaWGTvcMd/WsU48okGeudMCsvwfAl2n9hcGADQn
AZwb0XXHKveEwLOboeMDiMHowtL4pUIJlxtLKfUpch56mbnb1EPxMaVgzf4v3Xbo
LTcaxuGgvwO6beXEsOYvRonRrQ7S386mlaqvdfX2sFde8sswinjlUdpmjYhlRV3R
gQzTYOoQbmbdEY8mHgz2G1PQE/D7hp7cic6hOBMVu8QUd5SxBv8rn84KA8Fe8MbI
ZGlMBYrGD5RyMB13OhKvYxbb3M93TNxe7eKyNq/8GKnDAhwLJbsPiRJJvGORz+u2
iR63iJE86aHIPGJWFdN4dPZeLJjqqdO/hv5MLKTAUOIgo5oTAGi5whVqt1hjyzlO
//sHisSh5VQeL10MUC8sfTf0tnhKxV5MM6pLe38F94/54Iv53Isn6VScplbRVwJ6
xCf7IyRH/x58hAWGFX8OLZInWQ/NPCWE8pr0GmJg/ubZuADIpslimDWptKYbuBKa
UK3B/wSP7QdA5SVMNxxuKdPHKEjlHK70CT8URy7s60PpxDGfiYOh1lQD/4LXlQED
6dsTrCGpmhrvjvvqhDslPg0ShujfmkgJHtVWeTAWyhk3rDywsp+uIiIYjMUOUlKe
xzx3f7wqS8m+PvoePBXfQps2OYQvfkAoQaN4juaOxJzCFN6nPWbh6NCA2IXc415L
5GbOzLhAz8HE3YqScQDHOPSLSxtxsV5ZDuOkd4qyKW1+38FDGWAazNdNGBTlJ8ld
WA/jMBqWOD61EsDaVoxTaxhXF1/FKuId6wkUloM8vz35r/+m5tOlQRT+lBLzhmNo
C4aMJAM39egk5vykMiXYpIA1fcA9CdCqmIAeqx/Uc9P2TOsWXs5ttclmEsDcLx1r
KCc/9OmnDprN7QkZ0WoVPYUT565sjuwVqtaTBzO/oDhqW41VfISbqWoEpAeQ5qlJ
KMoePNU2/GB9Sc2gpn1G0+rtvoxh8GwPokpZINgxuajaV4BNi1uUzAGzVG0QdUUI
ZreZrsW4azFxsygvt5qH+HI5GSmz8YesgNY4scg1Ge60YuCOiGWRFibZhbTn7Bkm
GfAH2Sl8AoRPV4Di2criBxVQBpdVaWrumAAjXEaK6meKjSu6C9ZoqD/39Cn6qHoK
8JPU8EF7koDqicHfuXzIuTQqDn8zsnJUa57kXJ4nvLQzFOLbPf0r8PjwXQOgJVSB
AQJOPB9jIVuFRvFfT/LQ1+PnETV1Et8kB7jtKSuQngH4BS4iBB66QyZPGqUmnLAL
fvFLa1/dafNYFyf79ErQAiICZSkZu4wnsOGKkwEj9GwoHHpmks5DY9wThH8kQ8O4
TAUczx69kalxkMdZo2wFDaOdbF5U1J219i39+QZe8qvxRmMTOPhF6CTaQvKcDBGj
QhSin+DycbZTj3A6y60zqQ5w0gSsdWgGjXXgJdzao9RoG+8ijXciRPU6iVQHkj4t
TqW9kJJnaSYF0k4HwffMd7+Ji4fojfouS21ERg6zX2+HvWXbvdEqa/kLb59ms6zN
KMUPnMznOHip5WmrcaAWcSisnuZ+w/ExH3lGeaGhn2RLK+9t2VySBLX8lZNh/gZq
7DV461v6KpqWLKBW0ZNYayKkX6ZeUj71jiUSouNKShnhebDhRPpbvy5H+iyYK2d5
MebpHWmN8rawWYyQagBX8PxE4L4EANmgrPKlf62HoaldiAwQ5ndatJgHmBRePMfn
yzwGsobWYakAX1x0+FilEtnrcTGwM4/rzQM1E3L1cAGNt0nv7HB7CKUPK02t4Ybl
p2AzASOZom+HhaOOxUjk+SkDIt9AlQg7Ovkm1WFiSCA0hZZ8WtHDw80Lf2QEcrxf
en5vm+12W9D1pvhlG0PlpEpQx5PDOQnoNJeGZXkJql75cg8lqa2fwkOP9+jSBObK
vWTWAAB09k3201NDyXwyjLbExJpbnl0ddCN9FVKCadTOE8MFgTkIrDUIBryWsHef
iEpLFbi2fa8aeE33pNWNg9SiEnxrjaOSEne15mzlHYeHeXK+w1e0yfTu8bd9epBl
V0yG37tUPjC3xo2YR/effPTm8WfmbdpCyYuIVvON3IQstCoB1GCRQsqwsHZvU0Wo
NifZ+95re7HqVXDMm6hY83seJfnmQR7UUdhuLwYS+wRuZYRDPdq+NXNbIiEp7T4b
9gGcTXERfp6+gyXmZBTL2enl90iTjTox4wpqs6Y5CcdDkSeQIiYlSXRuTauDK8tA
Y016bmKNQz53lEMcjJ15UMFwrED+NOrKPEF0vJlU73cnVsD+J4KKHplvpnaghF9U
AIDiaQwvcKPJ+t9TPXG8Oh2CfL28leNh4K7wP8g3z4cX+LVqSbQxvnQUzZSnujak
P0QmRu/0fhieRJ2D2SKSum9EYvZ51Rfc1bBmdQETvSQAb3WUC+bBSeyJEXu4X4eq
Rg/+2O50Ksx7rhF6NzyADbZSmp6VyoAf7nybLaVnpfhoBZnk3Wm9VcjfJLODMLU3
nGsncHsE4MjkNDdINdf+FnjvT4ekhFns8+XcoZjjBR89OjQPIoOYGZ0foHrulNqz
SUxyr/JVOTNivWCnD278lfdlKEnf5Qfo3dh+7e7MV4AICfYTrhoGHFbYj+XqfEUV
2BjTHCYA9btvi5HHXBGsR367IVh79qanNyA4yL5a0rlA0MtjzaUM1dBzzXoMd4r/
NQrKTVOiw9eC+mNNrxdb6OEBUAvd/fhRe1b6Onzmne8HUvfXkON8W43hfgMzbWrG
CftaNLvzd+SJo6PzfdhFQSCyrrrb7zpToZoN1rfalBfWLa+eGTqHnIV1anNED0CR
SuoLjYjcSzLs5NsMpTfCO3gCfSf0THQRE+oeYPegPvePUGImeijN0CxAOvo26eLt
Qwq71cc/UIIOHLJOjZ4m46S4Ml+FAQS/m322MgnhWay5MxHKbs+lE0uNM6SSbnaQ
h7QFd8vcpcD86Z6eCZiUDCj8V36kg1ABbqfcGJWmAdn7e62aU3uuF4T66UJSwQGP
JhVHqkd7ekEvq7jqzmIrHTM0haYf5HdvEk6m71ivNx4uSgfzmfo6bWk1V8QSk40a
Ap8Tl/S4Y8LryP7WPy0txENmB1eatF1k6V17HgC786R865dBFVHf2jVYJGjQHh+M
Dd9PFzozgmmSTInns7CMD9pAU8YR1B6ewVIt63rdfavZVKOXWiU2ACBRqZoERJ3V
6M4MsBmUk4xnQ3PFlKIzaRnUN78UBaMoWQMIwAbTfnPiKPRxTLS9UwHwj8A1/Ziu
6OG+3oLZCRYr1iTmn6QVwvVpTcanTGjmbZcyk1/8o/2vjiT62GXe6Wi2mlxgJrQ2
Y82VkgX5ylI/1dNxx24u0BIwJ92su2G1L90FjtuAQDvmKTEe2UpYnmq2gdJ5PmHg
fnRM2aiBGkFwfiCIk9t4sUkGIF/XKZxOcYQ3wzunkRcqhC/ob0on6IKHi+svXzxs
wQnCztaGhrHToIMei3Fpur8GnKO4FDZ6dk8If0IHVldONW4HSISj0crDz5tMf60X
W+5KMpL33Ejoc61Zcl0lFhYoLB2SRj1E+ApTOLRTIVJCperuSsjzdRehxhPMwF/r
BCbthVrAuZCbDftHtvFGGdoDRgtJr7pTqkMYF5dWI59EjDT1gvCO4HRExA1y70Hq
ZweIumiu7S/GxSHZYCOrQowOKn9s9Xg/1BBGhcRNrKGewqvVeo2msqKQsV4/Fc3W
OpR4WaOUbaBl0xtt++YHQXg/6qP63XIjV8CJqlxWohWaAnK13qCQTqFeVVghc2cs
5q87ysp8+Ini3jnql05Pbp3sGLRPsx2oGuk3LrdLC8vncptjJPKyhXFSBf4mdT4B
lwXcC2V3rMlAi52tNuxqKCV43mAsUe68JG7TDFs6JXjuXXww6dnaBOopEQaW6prR
CL+8ebOw2LUGBrc69NxMixbkfR3FZKQj13ShWe6tZjIei/W6OILEbVq/wSk5QJGS
aCSJ4rBiB6waGlHUTpt0ty0REfQq0a7wIP57O9k4fB47sj7EcEOZjtrJhLmpOdxK
nDQDhS/GdRCxKL64fFslTl9j5SFsgDLOvn9KDAiS0skh9mEVVGLkSFrSpTXYOD/j
emi0fivatrQguqs5yOp0bLf4Ro+CjlowojtwNZgtZ0gQG7Owl75WwV4tIYva5Bp0
1d7LYnQo4dr4Tac6jwLnGGy+H1EfOXnGdYkS+i6a0Uk2NjEYvtK5KFnd2T4a19Ch
M1spE4DET3fFaApO3TNknJQ5g+mzZUQLGN0JPBaoN3+ZU0p8HQ7JVahfOnSgtlUs
zvoF7KrgBmLjCuJR+6RrA8DjuOhQmU/qKfg1y3AJHyF+ZIz3KA5QEd2iF61szU4A
tGVUHA7GfUGgdduZ6Nv5Tpqyf35owIVxelfv3Gb5NB6meRqZl9GAuh6DbQlQM0zB
V42KmLm8bZl0yDJXYYRqSsr6Axas8cHvEFcrUVGUYc80G4DCfowAw0UTVAhesGfc
YBBiFZoBay/1R8k0crUwVS3DF3mcEmq7K8y1YRZRYtkf4Gp6m59OAnNNn6kIIpU5
OOrVx+VCXzAFacpb49XemNifiMoPGIPDOlBNoLcuPR/DCaUYjgkyOekDjoudP2Gs
nEZ/Mc4rMO/gdYx1nEJZALm+zxb8h73tZrTrIKR8VHUouGEeS3NwvbeUTppWxoeO
ecoptNOR6nbKa5M0j4dKzcd7+o9NX8oHrWIMq5o/rizPqj2o82x8nAtWaEKQHx2i
4b1w0bqUL9215DETqpfNkAEuSHNGEEopMrc2JfZhnsrCZF6MKRERcQWi+ISqOw3h
vM7j+mENid4QDqicGn6xJyu6z1Wuqrnuo6+UQlLU4mywdH0HsyTd90N26ipg9eLM
UgUZoDFfrunCs4q4fN0wjE8TKsLjTpKGfnt9miye8xoLsHs+GOz98+C4CJdbCIMK
HusEQiux5ix8D759amWvHAJOpxtQcZAsdHSOpWr1970CA2JN7FgPWsaCJy8oqS2R
86XYaOZPpMmGevS/5qR4DH8SJXtJtskYBKr2lp6bsvk0UOQLeBJgtKzDqUQcfL1h
l3UbDqP9TI834Zz/axei+QAqc+pTEQHmawPr1WuG4VRIdGbdUi0kfTyo4Ikx3buD
X8ZHSGEyCnZ1hZ9AktryQ5ljxWhlnw9+EF7GqONteNW3sPR+5JRHyX5rChJ1KuT7
wijhel3mz7KqRieD5ige4HCElFirwRgcz0nvZTa+xr9u6IX1QKCO4NPK9ifdNoJw
pmRSLLTKdGUwEHtKH7kVqySm0WUu3DeksYjYAk+Yo38r0yT01hzh/5/fHrAjO/c+
xVZPFN0rhcal//qdKlg4A2ipFMaAInMFDrFJWYrBMDaOW/vBDJUjLfVNQq/+/Bll
pa+Dd4VnCdhXJhrQv2FZnTGYdNjK+DAQJPZkUHC0FG7k39iJuiFAxe8koZWlVnYe
zu2XgInEkD70/ooQZiObewbv6+0gC8EfdtYrMf1MnhreE+S736MmknIMkGCSEdvY
5mQlSzfxjjGybXjQxFdQfKSjEEAjjEMR0EUFh8n6bTNXo+m4Bhm/YgSGH6GPR0f2
CEdUByDTXuRaLa/NrRLifvivv/pA53S1Qkfv7/kMQW1gTxHZRAsBC5d+wWt4ryR0
fjnCZftDA9UX+Wna90ffXvVWkC5Txrr4jiaX6E0YF+Nime1KOvuG+7Rt4xCS2Gpp
ToFfh/jGz3981Lw86pttddRj8BC38GVTH/Jjbc7hJBU3HNluqaKtfep/zpt3Cs4I
ZG1kpVZx6iP0sATSYMVaEQJoxn+j75Rr0GiHO9ehkPo+GRK1MtgN0/amWNmQhJQ8
D/ADqZjfxP6RNh6r7d6wzXh0PB72anF+ZYQ8fQNoZ5ODSOeIZkQdbL7vqX3jxiIp
9drsExqsVVWGpBlkyjExEX0DZ1bYcrKkt7hzJ0WyKAZ8s3X5+qgyrt+DS036q6/6
WQLfoTS8w2XBmb42b0bzlxAYULKuHeL722jday32a0pvOyIQUzB2br2OxofXW0fv
SB5DzVMZd/SMEDfPYScO8EqA335FBo6UQPIEzMKPJWr5MYDJG4KuVgNUufc/Rqa0
hxrLAEad5am2+e2l5aEcNVlSI7Y9AxD5HVdDXc2izGEWxZJ3Jw1UZI+v5HLWSX+a
Gv+oNmqm239EPx+rFQtgUWoUpfAJYoIynf2fxYdBNQLeV/dqzl3k7sBsd8DDTmgv
0T7quRmYelMbo3cLc4MV+/khSptXIXbiOQwaipyCF2demOCr1MWR114/GFlfFxjc
JlVuZf1yVju+K6su+bEHsBQYSWcdTeeMUkbpilQ34WkA/xu8vdrKx3DGD0srV4/1
MdlVBUAu9uloeRQsgdsW3i7M1FL7D0j0bd5HrijVZRXMfyiCAqIR7IG4pChSCPkF
MWLsuD/ahGuMb6G/vS3MbyYT3natm2Z8pDtMLOGhFNYNdqY7qV2U4lUJP/HfXGet
mBN1smD85m3zifFeVxQtzxW7rPz8fCyNBxdPJh+5DtNWdkrzM9c6ZCGvRcb/DxKE
cP6mye4ctWbwGEMNej9Cc9SXAq63a4fDWTAwqtmVS0yWCAqF+SAcq/QJ3iafh4IZ
2+vdPwgsvIKz4sQkmr4R/X3Rt4mRJKP7MDDb/2IOCfEHNrwEz+CgB/V5IqHVVeVp
74V+Aggu9SI4vzfo4sIQ+YPRxPPbcasZd8VfY9THPSO+MtEt/2wOFXnIPgko3jmX
LT9gIt+Zr1oX9UxID0kUUJWsHSzMo6Foe4AKcU9I+1LiZHNM+4xTpkVurxxd6hb4
eJBJIGYcevpgnIGLrw938DXGAYA/6R4hImxt77wkEd3cZez8JVztRqrJfvsLovDW
xbHNGiNSRe1ZuMM81Mpf7bgB/52/NnSQPaCuE8sYebKdUVw+DMpKtO6jQrbamYz0
L54Zo+wx5Xo8FBEJm7emLE2sWumU9yx1fLDQORv/bg6GJo1oCgQgAjF1YXk0xn3l
GjgJbkgC6L4uDRFq37d23/2YwN7Gx9icOBVb8yLyNv1NANMFRA9BVUWs0b6Tuf3q
l6s8P5DVYiBif0yncbVaM5/wPWq3LDuty4jqf//J2tAgapnY+yEJUX+S2Dbv/+oz
3jx75ytL+hMGXvuUVWBjrOjv285eDz71o/KveWAGR7aXsWWnQbCRUjUkJyECun6N
//fLOUIwhxnV7y/14nnK/FaojJv9O1GGB9WI7i1w0PX0v07Hr2Ni3YmsVAY6gOhG
m4JK4e6h4xOnr6hN4BCLddD/BgtMt9nD5R4wGs1i/txkplBye44NlQqsahCeXtn6
KbtmckM1qiFb0RnaHZ79aTob10ITh6mzU0BRlJr/8uBYkwxjIv8EqqdHi1Wn6nAL
/h4VECuTDxWrwt9JYPfaI04pdWH4DFJCNXS2uJg/FCyl15lKlIbhenPHBDkzqukk
KmwkIp41ZnCmqWWuBgrD1Asx3gSeeIVUFyhHCCr47gowHqz7C9nW9kbCY42TCqVZ
ryHpBvoCw1a/Ow90e0tBwcNo52lZo1j0wLUErBDpHMYKMRXkiOxgBHQXUaWNzSKM
qUYjKshm9srt6djxnzwlV7m5/GGgNRWffQ4cZ5IeSM1OK9jsjo319wn0Gj/MR64c
6tcaqFURilh5wwacrjcatyRfVyhrFmZnnmgDmkIqBS9DScBWOJ9k3DH4ZFQbZlZC
peufco21Ns4SEZQ036uCK6aAXbZF1wrBP7rIz9VObzrzZFsjzIJ+YPPXu94J4iFP
5nQOVdtqNfgAla0tcJEKkzN86VCBjnEHmX4itn4ZrzUmSiJ+YZ71hiO+4u4J4CIT
eQj7OumXf9WkqyjkLYOrkMZ2c3PR/cJnzgekIe/uJnGxxdakITyXah0bm98/BQEg
84WO0ttNKkpgsFxfLbo8KD4DHk4m1n6mMMQI7eLiRt5TUwXS55Ndy1rHXVS5yRum
EuXK66V+aarfg92XHpqo+RHer7itdmU4agTlscgcL8yiRhzvJCHSsU8uYmMKh0+5
jqQ5KZ/hKRtap5SRBVB8sU5fNVBimUdqEUVsvRfeNiGDc5Ze7q2MCBRM/rHxYvm8
m1pVazPiRIdb0BiQGcOe2pp2SNS56be/yLk6QFF3/dGePFmZbJhvV6QgCLvOTkUO
dJFLj2Q3/WojABiJJ9qtwr/HTAPmFXpZWBn+nGFMcpKIXWUiEH/Cc1MCzBZTsrpd
4y09g3XiP9bBW4fC8j/SbsWo1sfV3N/vWoYwIxwdY4aN2w/6jdOTxMKlsEe4zxmG
QzhK7MCKnyDHmNmPJEUOY8Ci1/hApT9/iV/dli9gVWkLnJ2Hyw/Kdxi6yqhUhYVh
nJgP9EdbDMcJlh+f0pXsFOnJKtkD7uuxFbVkFKyXpIkg7EDzgyyujolumwxyKS45
HMW0aR5YYaVlW/ZCW2ivjQ5lEt7p5NLqtXDjpkwA2HVPHE8pA9a9KZrHkaYHiOnu
+Mj/CvHV07SSAz0hxNKro2IrJ1q0QrP//H4Y818heyLnaAoITXUZq7kGuskAxKD0
8qIfCR/lXYlPj8INSB0lp7KD3lmFBycT9yeUfOWjjFewPxrcmN9aU1j90mnmWl4q
nFU2yoPUQB5vvtdViRfaB2ycBw+zzwx5TAS0JBk6/9e1xfUE4AsJRHX/OdHRV+gf
evlWSOx7rpkSvAkM2S4+cep9xpYHyJJzvlvobHKMjoj2lJVWq4kJVPoIV+n9qeC9
mBSJR0dDLd4ZIj+lhNmXpNTs0KnI5PtTdLczzhpIs8/CUUZBPKGJpzyb/0x/UH32
wEamRjpQ3G1CeeSgvWuhqp0dyejwqhrBjwpkt8IL+FSh7Lx9b6uoecs7Oh5rf02q
PZumsJYL6ScKukeWseHE2aepa0hTq47V6lNFTFCaX6EinWmOkTsQ0P5ThY1fr+Td
c81EBkckCmtYFVwplSs20vmghRtKZgwn0TiR4yjwPdIuAXZ5TKiSBjHz8bST07Fq
HkzQjkODSugdIbX7X75WSc3vHv2NWFFWKLDLS1VyCTVtongoK4L9Ta+IMfRTBTl5
x7489aEjP+48wFFyvq7t92jk9XpdxhWNBk8Ym8BB9l03/KcYJBT35jeXsMz2Xazx
o0sQmPEQJQRjxwIslEaLAqIGlVadnSD0RflH9GFiMyTIdAbjSidW/MkxqQsQHmrS
ktozbxgR6jSL3nGD7A6qP8ppbE+jqvr1kV9UApGPIgyf7Hmwu2WJ45fuhWM/GZWJ
/witKZI492FVE503IPbKmnQ8qgPSZ419IPBj2i3xun4cLntuRKGiwVu/UaSkGo5x
9ZdsG3q40tK4rKQmpK+oYQs4U6UPSDnn85PBJkEWm9MYaaWrvNjZm9WYxJIP4cg6
2V6Bq5ixJ+4bolOfkcsw6WQXpcyFQq0t5oljiS93CXFQsMjtXs5CQxQUnENZ4RRw
73H3QZxCpIyjwbzJZtOls7lpatT+HQzL/FbMWRXim9OZLLKzXKuq1JycG1TTcwFk
MhgFmicVYlRaiZRb65ST/kLj09gPj22CSeqnejceJ43LRKAow/WKIoKJSwZm6/V6
/awMd2HsRoySHyxTN+fdd8O69jGrfCflssIdAmS1UoRtG72mEbnwGiaJo93LwpyP
dY145jh2bvyld89JQy3EOVfEN2MzMwtghs8vlv2GtzzJeWBQVnwPM/rtr8NxG1J1
3PvAdFG9IDqg6mMVBBOK06TT3qxvRo0MHs7OFZTxtNFoLknceRRYqGIKbhEKvGMV
ilJVRVHuqdDIAViN7r8rZT8VVmPbIdDuYBVkcto3Sg/jHUx4jM3ZvvLgflaQhgQo
TQhRH4WgzPHwp/tyYKWYc642c2YHjqVxlzD344L3GqOSYfW+G5OGuDRUi2tbhtcm
xdaqTicSe6pTrIozv2id/0hSSYDsR+02qbTxG/s6rPXW9PZFdhBzjADtAm5YVBQO
tReSOBI5m27IcTlmXAFU5kcHWGT5vTMJ638RY4W71BP6p3kLZdohqRlmveqTx6uo
j8BAGpOvPAcA0A88wGndDS+SjuHE8FeTbQ7skezianugDii4vT9JdNVg1UE0fvwY
AYCjhBL1eQPP5fTocf/XhQHF2vQFVJ/vofsY5EM7iwlsBuv7Wz6FQKgAh8F0oRPD
h11SdQxWRqVfmehwelnN27lDRr/cqv36B/XndPBMB+39h/iCmDULWwW0LkSCSv3/
M6RgpmjMquENf1+hHIpgmwS2HOap5vu0gIhhHy2i1clGjrWPy+QWTDvpXG7X3lEE
W21uR0I2V/obB4wMqIyDwO6ld3sj4Kz0bZR5ojdotPUddiI1HGZI7VeqtN5dkZOM
yYuiWtxh+MTETyJdXuHxSlvPqXkdaV2DY/e23m7/Lza+YkT89S9TZu6F3lBVHqYo
K1Em9WFSzjEEZmiNpGXepQDuL3UB2tAALTiZ9dVEx0z9NJ5DFzJ4orioOCJx6S6r
6u74PJo2yYcvH779FFwT/2uwUKg0rY9zCYYvPlEBeH+mFrnDSWcBKr+niw4rB0E8
aEfFliZXRPj5gvW2qHmZtiTbLGedkaHe30WwV9PfYEo3lLihqUGEFiX7yKLxHMiL
+9Hx1j8qb78588ieLKVpHJyS4uc/r9PfqbwqkFATYiGlhyfz8PfcEuVaxz29eaPk
VSPDd1c6PDWXjjkDe10TQYdwGZCd1QROgP0RTYVxPWfVX/JBhjChM8cEZKIuEezW
TbwQMEtl1qbYHEOsRCJOWQZSrzdH+JrPcPaafhK3UWoZFlNFAX0f1ODi11rS1Rt1
KdNYTiie5sGoLbYwe8hQeJGqRO6XC/tQPlPInUcwkAE/Cbktrp1kT53gvFP2asib
OpDzeJ+3DMJZm8Y9pCDHlUX65rWCPj30Hk0FFkf4SqywXyBd1ehB4Czc61+nBDLZ
06ZRnrvLCirYkqDSwMiWIAN60ddxibPJ+205WCi+6mK1Q3qWtFMOUyOb7mNV+aT4
lDgLXQzYtr4AGewRs6TDGku+fliqrJibEYRH5iJIfmQSpdU6P/OkX1y9vtW/5DCR
5MzqAyPeE51mMqjAoYNRGPTOHZaeeGK2D+XhRvQjxFblKbO7EG7QIcv218vJShFW
kQD/RTA7pj++O0uTsNDlbK3awjYp8/l2O1KU+98lqXCdUtp9txjgJ76A9yzd2BJp
BSCdJdjeE63vuGbTQdG6r99buNngq+GTM7OfebZ4JilkSQBXmDpprWjKGEHrQ9d2
6AJU4vOXlqvuZiJA2w2K7ZUJP6qsmevMIONAISwV6uNclnXwrwBlJmUPGHPDDZWW
+WPbDySma6LUrdlkjt5veZUKSXSsadXJJx8uTRLc6ktpEqyk2X8PDdXmPpup6xe3
+Mf4aj0KrgygM7SZVG1DH3iPWx8ZWfOYRL5eZWbmvMSw7zNtNh4UxUXTE39ZeFRD
6xLNp9ubrNS0RHDIpaD35EOdkPSvWxChHbost4mPZ03CC6qUwCnlNB1xyUH+lpxl
ANbS5ofwEDI2eZJmrxGbVH+i6P7hu5KeKfHPVuhrg8gx9z4RlQgGhy87rtmdeLGo
R4EQVWMKmA41jKqve4wKSyKhg8scYwVmFpcY2EiiDBD5djpCj0LiHpbp7RIlQ7G8
mmXjXf8EM5Tdh7axyGTYIXB52Lngo7Ga1li0CjglrZSqnYNKFXMDssctAqhfy9gQ
EIurcMPK3qwsS6TOqyBXsS36mn2bZ4/Z2CuMpCChIw8aq94qHiZTEnQb6wb9EcHx
mBGBUOoJjNxsROAuKUB9IG+KMvdhrCfKc0ns1rdXLJZ5xWZULY1nh7fCMGwBjBB9
WVbxlC+feSzYtK9rgV9fAY6ot7TbPrRbNeKswh5/Wz67xvywJ+/yDVtdHnpmgfxT
1BQtpMD+Zw3LuNtPFT5TMbrouQLtLa88JvFmzbgTiskTJTOJsTh6VL5dqA2fsobm
/nUeJLiskmrHlzNaIgyDhAIBmazdAhwycXVGDZYIsWEKmIsGYjrytcBY8BSMJ+Pg
VG5ESBNdW2Ng4ejfRi5WT/u/DjTzCHTmDA7XmWVfyjsC2U39R+KrYDo09MY5StiS
YY9MWWhVrkhKaBBIbyQESO1gSVjgs0REYdR7JK83vP+fTYALWuEVC9aDlQaeRKdi
rrjLd6Nd9r4X3ki1kguMypJnIlliAF6NIV6NwXf4HHop4D6HaQxtWbVJWfqntDI+
02OSSsLDhh3cOyDEe2sfqn8uxKuZ+bSFxzFxE7aQx9G3/NSAl8vSREzX1wO+gPEl
fiKxLZbQ6/vCsnG/TtbGdGBY3m/PUwhCxz9U40sKZWVITUQotxVPcqVLaNIdrDR/
oTmY7ySTShemv9IKtHGxnpD+JwbDbTpQ2grjQyg5+Vp5Bk6YZaq8XD3t6QjMg5+w
pXcDVQOO0fLPY44EMsS0gbahzga6UIhTV3g1TgCodaUVJ0KmxubiJjTwwf6Psn+J
M+DdOWaim01ZO6crcqpfMGKrnatWXVdayyB2DnHmPM2wTF8NIiDiAvXPMcz7j4BO
wYxvY6F5hnpISlUe2sYqpOFB4Iy3o8VNID4jXcP+Y9YKGcoTHni7vDFFrI0TQvVG
j6NheqjpH/hYihZuXJCHM0CrfW12BbEVfDI1jaLu2SNKLx4ZdG14F2jtQBarKUO/
ueM8IPgC6bNRc1GgXhMCRsI7iQ4Cr37iFzkdtdeJszMTCzYZ0yTU/Rftz2w/ZdpH
scMjLtKDfHJKSatV/gLszhD3ixWpb1jioZuMiddqJcfd54bhJJ6TnD8tz4pvCAHU
yGS9w1PpAfAi+ip+kjjs2zsqn9N0UE6/2+frQ5/eKrgFpszkNGm3z/So0qF9IpTk
aX1KP0l3S4cS3JfT6KCrhL/+WtAU18CsTWPsi4XcQNfzG15n5SREEuE5gM/hj0t/
+VNKsaBjPgqXJymlrsprT4ABRjj6QTf6EJS2WrepCZQgLxLrz9pQGmZyEBHmNxN8
6sAUqm4H2Un1TIQkPglj0emlwXVF/S+O9GtkWJQASF3xjh2rmT61DkSmTZEmZ+3t
txTzVbS2HMFKLp+9uvySks7BKFAMzXpVUjzeFDEc0BdY2alMVw0VSZcYQ5vAR969
29aL913VCnOs6zyTc7+Nmy+eVXC24+mdby8C4Uj1ZOIFGBXafchi22JZhwVt5wZs
TMj8zXdy59u2tRlO7u3THAjBAAT/8Pt2g+wTiyRm+6Y14UmtgsIuuEEGENc+I0Zw
HEKQ7Wm3ni2AIPGIaArEeMsYRLl6cKsfeO+JXQtz6Y3hIL2FZ6/PBf7X4Ylf32vZ
U+8B+wr/ixFUeiXV2QfJKm82U75KM+LLf8WSzhtCwAcl3svrqTa+98LsQvsPxdzk
W4sE7nevyLtdb31EP6e2v/AWLRk5JGZvkdewJkpM4wKsumiJRuuSPrqpubVTeTw5
svaOz0dyap1ui1bJ2TRPzCTckvvxtI4/iChEPDC1/H9AxQv4487wlYSSjSpw6jCR
AM7sdtDwLzsDle5dxhGznAMRF2e9cXUhf7YI3aFpPYmMw8mokr+mmeN5S9rx06mJ
PSsfQ8f3kHRJX6PeRo2JK+chbo6ZZ0nJfk2CXD0ptn8Ager0x6+6I8XRv6+rgErC
7rJBLLgiS75XkEYzZRBk9Qpe3sPhrjjwWYv4SpayJOlTFv8dn2/6POSuRC/ae+2V
4LpVImHzorMmQRrDZZ9Df9ARrQdNvCaPfd2FdZyPCi/rdeNCyIEL/8RK3kIDv6Of
NxAX3dDH723+xaYVPCAROpm5FEbgrkztZWdkgs2tUr0IOWbNeo1AInZtNhzSXzFt
7kdmo+9XPj+wxyIAfzWw7d3x8selxMAeFH9WETPZUWnussTQTacVpXpmVprUHCWO
2gbfWMDy/n8sPc5YCtaoQk4lpPfaUN1Z5ApyZgdEKf32yCg2r4ILpboFPVn8I7Ut
Hh6FOhC2cpMjB1WKn+5PAniP7tOZsnmIzH65lNmBh534HvLEJsu1cWx/QI+1AE9a
soSY8YDYaqMqdd4HLNaq1IhSB27Tquvl359sTT1OGxwV8cJMkIxCCrIy3HFmxanq
pql5Q0yatkoTJ4A/0IUvVIOMIudo3b/QICFBalJTSiXI8a2ZddmLDFQ26mMxPdy/
HiatTHYvIZax7a0VqnY+3AQXd/CIQosqDOPkw3OK1g5vDlELu71EicL82B85Ylbe
m4DW0qsXpBTT6cukT+wjTQaN0ouJKFOy9QMS7WV5TFGqrvbLEdqfZ/692VEAaeR+
32oGKbDvVh3OQI0VIQoHYJ34SCNGt7gTi6Ykhi8dNHu6kpq30SUyoLyexBP4gkmd
/a4um/iYRKL8WW8welEHLnvxgyhq9ZcSaZpzEGfHHlMX0g2XnbXZuhwP9A//6Uac
X9dvBK6qHN2J4PGLLJyte/ul5Yopj2j+4pK6bJpsp+eWgFGQfoDLt5peNdZrVRG+
0jT6DHKzQqhMJja7Hn4GpIIVdKoIX70QGVeq6kq3ObUTRNAXqzTSYc8Z80xA3jeh
uw2SMC/iBbscbAtkk96sxE+KcEjzGrVDJn5DB+MVR1stUqyDvlXe50R39tW2BjJq
p6sFGcAOTozwqNHxx5YoYSj8S7/yJtL5ON24rU4K9ZnPbI38LtcQsPl4Pzjuvkny
I72LafDYAcH3ZvtmxW4n+K1KjlyVHWmSiW8IN+OUz3OemmMM7YqmdbbwrWKeUb8y
Iqiv2UtvwLowZLWdr0quqJXpo5c3Gv5yKy48a9Vd7JsHDo7VMSxcyJ4wD2Idyizt
AdHsk5XqtBbMSv5P979lEm8F6ShkPf0m1rfPgCh9oSo6eufzj/HMEMhl79j7ywqU
hrrgh31TkNabamFdf9ojlQkJWpNaVkxoWLRC/jlWQU++1hKlDMzl05x/iaBNbWho
f8XPIrI2z+9Ne9iXlng7RW+beE+l4ZxMjDc5gtY+ed6Gny5j3i8G7tI6tDGLe2LV
lIUdU2uF4ARrU33zGjDWcKpJYp4NHLsRrxiQkiGgkDsIUAmMwZJ+nVUITTed5wlo
YtBIzGpFHplQfjaWRrieHkhsUPU27i8ZHhDOaTCrxTXxR8pnmxBz4/JtDZ84EF93
19HXRXB8YmePSyfT9w/PtyfzcpnymT45nMWw3O7qD3tnPZIJbRMKz/pVBVUtj3ny
6TxK3R58w+PLdQaFHrje01pbsgL4Jl7sadegTXkPPT1gql80eBjGmSuH/lyPdyv6
e4bnyuQ6qmtckLn0qQZPBTSt2F4TybMTKMmUmYayZQXBUKolwBlvDg0UXwbCTnvc
Ati/3nDT/2g9+UCHzT0kKZX4TNnlxVfYtyIrQbA/PYb8akLlXlFbi3RgdjrFKmDy
iXVRnhYPVdyR6uMBBxSRE+Jr3uquHKIoWSzdr0CBaJBNkNB4msq4/7WOjJ/PNhah
HzfwDMSlnsOQfaUOCpq4QkMe1+wzVh8m/6AMV9tdnVhuu+sNTxmx1OplfoDWovrz
+XvOM+a5L46XhTKjI6aE8wesX/RBesdW18W4hzeUMpx7jF9HnE9/wZLeX/ZiST5d
qxYCjZKU5a0aIYAbLYn4iW7qtDewxQ18C6g0FLimWUSKgQtxQvcepnHLLgXv+Bor
MHZBOTb5r2x4HhpFGo6FF8mCdsjZD/TyG+oNMa9XOCbpBDF3DXK9tPIavwDgalLU
CvQHrXCmRr4i6UVxzgoWuNCVojcc2oC/Ch3FpVDYt18Uw2oNCPRJRO3FWX0q1xid
etff6K08UGxuzLTrIJdcVJmWQi8lbmzBBwK6t58CMAggJ96HnbRFXOWpo1fQqDth
7us2outmXZmdOVfOQt1zUsCzchtcb8Z4BYS0SLcAaYn+lbrpS2gldF0pH+ylQrXE
KA2dQEzAOkZXgYTq11l0NkIVpWPjblcJx6vKN6ta4G358A7t6XLFOaWdZZpWCkHn
nYj+ZFsP0QSKT0nN4AHSCtkWXxW09K0KQrRZMqiu7olbgpVSQUoxamoZC5Rn4n70
z+laexvk67NNMmsomrFIKf/8jqvm51KBXWN3+8/eRj5KsIGbcyqaBXE65GZHRpED
Qi3f5e3vVr8jI6dvK41aKZ8rPI5ln963dp1pa4THKNlPB0ythbnB4nVerDzKhR9e
zHgZdd3RQb+anpyGEQUFOvi35l2PlJJ96XXlJz/fwBsAdnHlP6lJZwaNOAtj8N2k
yoCnWfwNpoWTBGl8KK6p/5tBTJJMtHrmi+ZTQ6v9gnwKCnD2z2m7fzvxcQcZJOyO
NStjBbGalopYF2Kpv39hbZQ4vFdLA+AjA35geXx91I6ODIq6eZlEfeUdBN8o+Lcu
W1EFnSOupf3vHqd5f9GvuBiZC3nkOxl0v0QeiMVKL40Eh8JHMWGJsY/+UgTns8gI
ijJmrBGmTY+31Khq3MU84TQ7bfI7A6bAiSdl70VnPLn4TIRFRPmoIMOsPZB7KWpp
1h8aOSsRaERHYvPrqyS3UyQnTuZzbkJ1cd1qjGrzzx94Td9SI1Iin1cvkmrmPfOf
fn/dcuLrwHi9/imbcm4sa+JLX5r6MkmBUMSgFuvxAo1wTtYV2Cmdj41/i/u5X9Op
ElTaDLc6ADIIlctq1sp7U38Hb2iC5PcH8EJOCN58+OiQozsa3UtKbiI5hHQGCLwx
+mAaLx9JRhzsQrwR3wcOMgoal2Hc/lPM4hD84pBJlfrMIQBU+yBqtI2JkG7dHfdJ
mQptZVWkmTwFD/iYLTFHr9w5o9b8Q3OLzGwBO3pNeUHywvPAvdcjFM7ruC4a05I0
HeeDfJH5H3HD2Y4c0qKBA1tWyrbA5aIBZ5DcJoNGu8sCFpxFzo48VnWBaJjtvQ9Z
JoFb4d4oLY+tZCS/dEVGKrVfsQbCaGTXzpBVKQXPhwQYjqshWvefG+YtLpnqp0CK
8F/BAz+WwF79WQpCdmRuILBFmV2bZZhW6pZP0r6+rXdARPQcRY8nJooa31A2bsYv
OePVt5t6VOUSzr5HJq7CR874jaGgSjtovsrdCoPrc0ndlkuRflKMGtNIyRFSO9/N
aAHglhKt03PzcdFgKcMsIjcZd75YHa5cc153ja+agI8VOpp3ct4/M2ax+adi2EzU
BZb5rjBy5MLqOH0RedsduSZBeLt7O6RUXqPXfjqH/7edUmSdTlZew9zLVJEwwqKf
6P6lZFZ3O0tnAgHdH87BodxiquALNKdnxIn21EHpIAWtmVlwsJ9myBUGVuzmqtap
2NJjrBhB/nUBoQ+XJtBvq7p8De1vmU6xRkvC5VghGuf4VwHVwbkMez67tBQfA3WY
OdpCqkfanDTLI/TJcQcn5gq/Fa51Hmjz9TZiwHzDgzBd0QLyDC2+9O6I+hSSKYmC
8kp7yhgGs3nkPEYVAr76esoHpApKe9Bq+rH68d5/ek5mRhH41YyvvojA74ZoJf2h
WNQ0Gam5CHYBbPOHS9O3IUX3wSAcTduxTGccoie1QRGxS7B4nuXYSUlCHpr27iup
Fs3rD5aOGTTo9rQ7MDTzp3n5ai+Tx230CO/G8SHW4zUxr7MgBIk6b2dl18iGVCgC
xFKoe+ZPcEDpPFweBMtgewjaXTCQbLJ3I+3bE+Ez5eE6ClZAm1K0FJl8t9GpDwdV
aqw8wZy2sxioKoBHSLoJR17wNAZVM7HNE+VFTWqljQzAAh9EuXJMno8/c7Qqv2LZ
X3OLUHDyvLO6UeAfZMkPlKh95bahyE7pXU0C1bFP4bMdtRZf/9LWlDZwNhYXzh8g
AnXmVG39cevXQVK1nnNcY4HofmHxG0gcrPwOCXx9Fg8IDvTXxa6uY3lo7Y4dUbdO
BhV38T3c8hYIeIc05/MTHpzPYe/pCVOKj4aJwANWv9lpirlSG8FOjxWXiWT6Mrhf
2FH98spqjQPsPEFZtx1qAXbZvatMga88l9AWfzr1/BFpHPnWSsPPh3oKziJ7nSLf
wcoBghHjlMRl9++Kg+6oJmQ3LQfriNV4eXZFX6DwMHLHvxYQFagFjEEL4BwpXWx2
nRLZLKPXqxVoca8XBnulHmn1vM/ZOtHBjeXpUEBr9f8q6wrMZXxMn8N9V8nM/aEY
4lyiByVRbI3Aa37tVgKxR0qBjs3Ivtc6YOpEpe2kSWsS9knizYwlbwYUKm9xLBSR
8RHCdb5wDUO9yhwKkkHo7FF+WACH9+qzfrf8vLW7I+/VDXBJPycWJYnhAGYDEjjC
o1xBumuoWemZkkzlrIXOqElIl2tBpOLNieCxA+hNlPZ1eMh89/ex3SJSnNcdh0Vs
eHZ6xQrYSG6riJJr2efdbaKx8k16YUlCJIsIpaBlgtgx1IwqJUXIxQO9if1jfATW
M4pEQ0GaHbmT1qChqQhqrDiLG66hZvPdUm6EqBzlHHbF9DIn7BHEkDKSSGrE6iXD
+WbRZ1flCVq2/TKt7CZ2paUjA7v98ZN5ojdDJD4YVDHWyY1T7A6LqcCMHKQp8QwU
zGiKhX+TtorXatXSPgREarPwD17WqON7oV8K3w7b9RSeUbp3paf3YtjkYzKHdhEd
/PO6ocUrGzM375FACAtWCvT1QNp01RD7cXm5jC1pvZN9g+BZDP4sBeOJMsN+Opml
u/VFASyTh/8Isp495VjfCmbKHCogEJxohdP2RvpDEuANPoGi1zhS7ddBh4hrjhhz
Uz1lCjgk1C/wdttrVPbzBJisPxuPSRM2sLZFjWGwpfl0xnttO4wh/lLoNPy1riuM
Hnp6XyBzIa8G+HaaWB10XfXutahhmilBCUKD7pfGIY16BIN/rtiSijNAlL37DPK0
WI0gozgtDkaufQkbq+4kOz2bgLYzqEKuQtdaVMdsHaZKDukPq7NslNQQFDQEsc4A
Z9ocglYchP6sRUMSeU/gC3u9QtqALmqd4XftKvNwT3xff0qFXX6W0F2tzbj5JVoy
3f1Ul+dCIMQXxW5OCYU74sN39Ew9P66N6KAFAoEjyVH+arSSf80RzfxZzBrfgyND
h/rz++tG7EAWAXaOuzozNtT8dWOUe5iHArYN4LDnPUCjCMZGQy9uqlvG6F0HTWCR
OhRSHvR99ocLoSLAjQPUNC8vJ+nc0pBlJEYWlLUUAqx8xr1GwZZ8UBiBqoeiG41h
rWo9Pts5jY/e/tYv8Pqdsbxxj5uorgt7zrFxUvo9OQLOakU8vJzdtUTzV0I/SR7S
GU0sHgUr91lv1lgKHNSz+jDKmQx7voXi2o2g/O/f3FtUTWXilBEbD4qSqSHwLE3B
jn+ZyBAnaLWI4xZiRrZjIGY8nSaYARvd1kFiUpI8l1fQ0aosbZjee2iiJyhTKnY6
XGtCq8v56TYRQYUUh+RBVW//F8BrYRiS8fV1iEEvRBPNLc6lG8/irOvltbiIU/T0
UYwcQXvEl3aY2BUugNEtLcCTXEruw8JX5Qgqb82Qzv0MjFlvEf2vdzSjR8+gylRO
QD8wYt61aKUKS7i5DNUuMAGDXk15yAzuiAxXUmYrWqVhILvxnDfHwA+7YHy7SJqF
qwnxRHlphxqPCrYrid7forUZDsA877DymJaMJSwA9VGNTgbOOIgyv818PbUKh8kS
y8x2pNH+NYXp2kHwydU53WKQMMf3813gdTDkRZoucOevidnudxvhMdTK3tAdDaxU
950sIB17THLAiuT9vDnZDs8oXJ25ME+WiwoYTt7BSQNCr9Xam5u//37UY0drn2L4
/DPSv4FK0TT1zwbOV6AhSBHskLrtJ+EI8uJD7M5pFTWWUw7KY8WfONIWXjqzmmQH
dRqM+qOJHvqnQYt3finLhlAXKv3v1iNR/6e6KEZbEiGFnxlJQjub8o0yKpI7o4Tu
/pl6b9cfx7mznhTScOMeGqQeyzDsj10FuZeICM9d2mt6i2FAdGFe84Wt420sZLVp
CPevhte+QJ5OXyBwRQUbMqaJklp19Pxhgnkh87dqF9/4fa+fqS5JnBhfH5NScDa4
QU4CK5gozIBzXeTA8haJ0XjZfFZ7xa21U6CaHAziflhJsinXvDoGouHohYZyg1cw
mCz6rOtABXwVIzHgvo6fIXvMsIa13Is+PpzjqMdxs2CzX4kRR+LlBKk5Ouk9rNY6
QA0H43hI0TzccJGuf/I9hRagzoET2FSrRbfKsrDHfpWVbgIlItDoTcFoLjGC2eQi
j3eLGg6A1Wmi7CSfbc0GeftiOkuChIyoZIpWA7NUQul7svW8fT06r+NEaLCNFKzR
iEY5xuNwiS2Alwd2pXds1tHIx2EjNUckcp8Sq8pFXWn5uyqTvQ+aLwPO15tYdC7y
JWO/m8R1vqUx8J9e0YXupCQg9xIoK30OWSwbzX2oSkGyIB4jaZ/B5Nye9PMcOtu8
JVZ8J0KE0YnQb7Y38KAuRZqHYHDRbDYofD5BdpQjR4AovYhmyuuvRGp056g6IoxP
8QNxyh1TWrS2KZBkE6477tdCK4HDUSYbiCi8v8Q8xrYDP4OwNWfeeO1jPE4zEQm5
29b+/4L1QvFqqeEx7kFN7L/KcX0mrRiuNlptb3Z4+IwSUs4NPlXKgk6nUWPdkCku
JXpgXgRNmz91rigkBraXLusqdNQFLE0jlb1HOQRjCz81wZuoOXdemRqhHWyEOJhv
AlF9hMYguC+YCBve4cMRODa+nSe1RRrsrcLrlZ47uo0K3RleLdNMFxT6ppjANXaD
UzoqOo5qyc6nDsketV4pABMrY7YbP+V8+rjaO7xyS0NWUwVwrT+r+a5vT57ZBG1+
UG/8sIB8IlaQnQkm/ywpq5e9MyPDBayqEY2u9zV0U0qylk30sXHCvwsR1M9LDV3R
v/Iz5TeXtpnNOrZ/uFiCMQzPrG2HEXuw1sRawFXERuDouJgaqGvV+moaa6DfGPEp
JJD47ShRsd2GkTih4Svfgv7eOPXHoD/3VLGi746+GoM+UglQxEQ1cOmQTW4N8oN5
wIa1OMadl82DnwjpQmXlxqFo5uiPG9TtqnvR6dyaBr2vXYfLweG5r+IobE/LffsF
4MK++GBHzCa9hPYCPx9Vqg==
`protect END_PROTECTED
