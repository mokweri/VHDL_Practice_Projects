`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HES6XWcJ06xPgRDaJ6l5GdNy+iUt7a/k8CY33/XOdTGWHRowHRsZGkoRsGhPqBaJ
Nagc67ie6DOPofWC89we2bJ59/b+saStu0vcDHW3e26ORmz12UHKe+iBbBPfn/oH
kmBg3HRj3XlutglQUoDnjl0GVduzYw8ayVgDfF8oYEt8PZKdtRHbIq3urSAevwmI
dtPcH9cP3vqIVMA4BGG7Dthq/QTj8ED31rWHktvJ0KupJSzIj8wOCtEAw0oLtz4x
x4dEnq/IkpPKHT7aQqs2x5jAxh9Rf55BAtnZYX4SigmPXNkpqXd5FkVn54Cj2aYS
w7Go4lo1p5zlnO9peiWBVEgS8X9hnIsFOuhps8EcdrUu80z+56suns/58QQzlBDB
RjpIhKRiGvpdhLqg80JbN/DvTUoJXTTTEQEHQ/nrR8Prz6i2kqbYWmF0Oygrs0TG
3Anf3664aj4Z0bYy6Rb15y4V1XHBuRM6xvT2G340KgA18lIsbnYkkDNUnPSdfvSB
Bx6bJ+3nvao7g/VoxKR4J4FG9Ea677h1/M5ouoFJpsxFQQxKzseIXqcgUIPSp8/l
qsybSJZ5akE8DO9H3av+eeEMLm/HOXF2PQ3KPcfYedRjZflsUaUtQp2KyBlQCie1
2WCxR5/q5u7+7UK7WBDEv0e/ahekU8Hsx95m3o1ZQjZhEdGSsAbNIpfC+/P9G938
xb4v1cQwDQP2sYCZ8ODbpwqBIq285mLIX2BHzLZDscH1bo5z3NMpPg2lOSRSaHJX
NBJBO3QsmR0afAxR9SiN7kOEGagVV1W8Zk5Vjzupox1JE1E/j0OMekepi6iGvc3f
ZrQBofS7+4SnujubrKyR/imSm+EYNO2yC0pa4ADAlZyyL+j9S7vgz/4H51PepGuB
LIWP7ycA1W3czwthHgTcvdy31wSh1N3/b61ztsXpNG+19kgSx2MFHqLOh5UlOBNN
X+zpnb3Ikv9FOIF7ARUASyHwlvGDv6FAwn1d0xtTRGqKSF5gtFUid9SZ+aJkG+ai
2WIlg1b3hJ7z83/oMsY9+jvRWRw4WfBwuD2xPgLnbAN/nnV9Zq7YKaHp05I0nuaO
Q1cPtU2M4qKZMwTfcZVwTRP6NyK67LdV/S/J8h/W2BdjpFHzu2cBJjqrKKhDFO0H
lSgktcvGVVlbopVJwuveMCqNxcYG5PQgzlWGXeGMQC7P+AyglVrA4oQASMlohus/
3AhfF4+27Lkz9NAcw8LmH29tV52CItVqr8U2Ejj1d4/4ou1s98YVuEFi5bz3pHic
XncRh9HyO/arW3dIRkxB++RQCmn1AHdXrVeStS4IWiTPQORrpFUqXnZOGM9Ryn3Q
BW9dxgsvdXaCUbhKdPNwnpCK6AwWOQ9v96RSBY26Iq4f/pjj7Oxv8uqeBuHWFhys
+JGJvX7AAtwecwxe1Fc0fhW5RSMOIFHGZtrPiOlXFB1jYHNq7oNwmVCJ9A/+Ojdr
1KIG5b7ppUK4UKtCULuoJhRBJbDz+4F5kO62Cs11kc0DVlofA68Dzgx6ZexuIvjQ
8TY3HwM3OCEU6dOcPJognvGRPqBxdkhVj8cnN+J3O4OOmZvte4xi/th+LT/beFKK
jK4uW3/tLeZss5hPUQfKK03T1fsFcJQn3kUN3CyzBUfDoASQcp6UzaWmPra+9wxs
7TfkXdCiKP1x/tYnNk6haeGUuS9fYMcJOOFP9Zvi11F92hzx7Ed9y/qyJKRCTRyN
r/WXDt2k2u08wWx+jIAZD7yFRNamj6mKsInpDxOF1qF4uOGbv9+jn6qgrpqgPSo7
dV+SrDZCx04C5BxixR+3ogldUQoS7emWsWiqmk8sADq4YC+DiPoaUKvuUf7tiVvC
8H0FPfxdfjHa/neUoILLwztXZB6dDFXH7mn+T4YP8Uoy2iCfIZMQYle/WXnZk/Cg
oaBOu4ggydIMOTwESDtFjT06TpuRN0mPxPvVIAJLwTehFVQVe8iIrCaUjru45oPL
vvlxmyenPw5IU8zGoDi+3mSL0rNeMvBBWnrqZ+Vn+ooun6qfGpq8/5HKZ/JrJohp
+XoD/wzqqoRe1K43oudtYKSfk3zy4Tl01x6bdvulsIQnKUnD+oZTFNOzoW1zyvi6
AGdf276DwgjVrnIG7o72NPoWcEy/rFXiny6U+J+JJclvmrf+RiidhmSTAIYQdxlR
0B/IsZgbXU/5oucPa29F1mpS2EZyllAQb2E5GCMeqFx0cJd4YMxO87+QocsZVY4i
yFvOfrOlhwe5ovBagpP3+ukN5CC9+0ekfHe4sE2H0SMxXjM6k/uUGzdWf8GU7FOD
9vTDvIbDQzimmty7vQyvfmYOBdHt5lvVpWdQDTj8+rP4gIW0QsvQddR8kvFYS42v
pkrnnVOPp4ktE7RWW2R/JMQyHb7xblkitzui+Y5r08t0cwHpwkKqLi6gccDELfEu
SW5Inz3uwSpY3yd++iZP44ceSuWMLYPvrW1W/TNXF2uea01pZVbkfjcCSJO3Y7tt
ULylM4NbXgerG+zvqzWSsr146R8R+kMqQuTFV4GtDxvxCbiPUCl67XUiVaAtm3C9
XoWPYUhOAdERqTHgMyf8DyZxG45IFli/xt5rKs8zokOPvAxJz+YWdb5YR8V39iMU
gs3yQJSUdjyu7qWVFWUTkK5v3Y0IfcH9Q88tsDVnw8Jy4rOQPche744cb+k6g2d5
Ph75qXyw9/WQAI7jRTS4nqfCna/hg5Hf1QrPWcaAiLKtwKbq6UXx0kw3AV1fNl6R
K28b14CLe1EzHz4o2URfpvxMOsYkcPuR6WsO8Ghpa/JIIFtTaHPehrhDbJTtpxcF
0aTQQ2BILJQD3sY4FAWKUzUJLxeftHm0CWf3fDWLhcPMsmW/Y2061EvDxteiedJS
JpDTLwIFbz6GS6VE3JjfRBy0n4kHXACqpbeiqGLadcFg7ygkJKvZtFIRyYEFRCaD
AOsiX+or0hzxXN4CNY5JDxk/+6YEdiv/qLHewGxAle+R6zu2rJ/NK+vh2zy6fdWU
tFAL2Xun+OZwlxAn0hTk0DPX4vzvO/fRvPdTDUfeEaBnOU6kIQyM253JE583h1JF
QgN9O8RGtSIWrMUxsYl9tCyvHeILfcLbq9tkE6Y/MSLJwigbBCGaUiEZV5TGNwql
k3goFosmeUAJuuUK/My6f8MvId4LfbGI5WAXLO9SB+am/Bp+m0g7jDN0+iUwXTqY
154zLCqvfISABoFIK/1IoBA0w46YMs9JeQIrtoj16+qvuzVcUzLTKjfvES64bsdQ
EzqjT/UQoasthzUAn8fpSDNnPFhrzpws4rKlK/6tbFAWrMEXdGYhOL7eOhQHE1NC
ScjemVtEFdEX9bVhNGQNCHDa7bWiinCctmAyyoOc2BM/UDP9lB2gBhdY3DtQowwv
j/CV0RNRur++2Wg6gmmgM6hb25GPUU9KUSGsNlw3M5IaZOJBki+vIRXhWZXWNdj4
UbpyrjDDkUyAnlw6fmxzS4prlKptnfDtpN5uo1oCoiRmawxK3VYwIiwt7Y+YCEpR
eDGfMRfpq6X1J6kQUBuaZxDsUT/M9dnlRtJU2lBZpHZxuLbKCgSXER3ufUW42MEf
9lNe384WyNHUzqniLjxwcK9fkyCpq94E5UIVGL4YRSgdCHl8+HwVa0EE84QQ1X7y
fQg79lpUpl77Q9fq2Bm3il59gZY2pHn9L2P6oSgY4OEQmBC5qPvW5kewMhWdioy1
H3VSCnuI6kpP5pQFWZES1v8kimIPewAhWho5XOetYaMnk62CmH+3aWkfGhK4jF/X
BDFMPzAxRhuz4aD3bW8b4L+JZtcf1RHcN0zfzr4ZWVZkMGUvqJzd8NPnjQ9dzOC6
n3CZAjSw4Flv9t/tKv3R41YoU74VQeHQ34jF2kDb5LcjITFt5wA6mXOWT5jiam7L
1paVRDDkKpwc0QrLc7kHr22C3s44t9kym8S1TFTvbnGYhbp10pXrJmNK6EQ49ZvC
To2iMirMIfkdGcVi5ej1b1VkhOyVYupf3ir5H11wxx17LGeg9pP674q1UBatjC8y
trLPnbegnWMQ6GaPTx81BQOIoAhXSLLUCCyBweJjpOMLF0E46NGH63PJxC5DG8P6
MZ95qkp5RWX6Wp/CDEUcKECxnnOhVgZGl2ecIc3AZc4a2lX98psDWfZJ3tBWsHiN
t9SHLTMjTfa0UWfPV5FY5DulkaFP574/gwoBF/ZhM0QmuWljxxYj/G+UbgoGw+UG
gvSU6nhfZYLcI4G7+KjCBeohyLbQOgWuqDA4Yrh3syUAdcCfAtcy2/A1waEzAYZ4
DvgDKxTgbBpQFChjI3KbrpRi5x58+q3+/M/wNLO5CBC+F3+mi7HC38ZJ/ayv91ht
WQTA6fr6eNR2P9lRTe/Qt/iuy3QzXmIJk8JpkV3XoOVTbh0U9MAPUZk25AL5aLKY
oSlTptOkNuOMSlUq3ydF6s42JjgqMAIB0JEo0FtzjU0od4Hxn8C5biFRVjSzqPrL
JNf0DqcrvEzoIefaoArAABRohEwsOseZ0qhVoLh8xjtFVmuTSOtLbElRQehBkEQf
ZDRolELL5yigTlrbFUVC2gPTdZbFd19e+/dJZ26gWFj8gAxMoYqCudRYL0BmN9Gx
7RdiXHssa2zhvuFwFTxBGEGxuDTDLBQI0pICKdUjG4ZbTApeUwC6xPDm4W78s3YH
+H4Pz01MYto9i63JNpXZziXqcvNfVts4bWYP5LcbOHd/+WO9x/axHstGv7n2z68w
l1lprbsTcYfzKKZvBoLDDRjfUECqUAhbvbt6ev2/HZnQTkB7iubJpDD1prv731WU
2rIEqBEUuLGoLb+6PoA0gMyC4gMfEyU2pr+1aTxldsdpIqSO3RWmWxAfLH0hGkdo
OJo3A2NLHz1wLVhu7LQ7alCqPbMtS/fOhKaoRCEEosOfvu5Nq0dn7GEoJPOHIm5n
gztklqTSfds2T5xeCUBlL5U3WwAkPWgU51sKkOrD7vZH1QSKsCTl0hNS7mdPhuZP
SFturhn+x/IAKlgtQ4eRuO0W7I5a2aLOpRg46deGeWVKJewq1zjnYnplCfv5kqKZ
rIzs9TwUZ9oME4PAe9GK+mBXRc6+K5Sk1m1YdJB0W0bMxq5Mg2ftI+unqWBKtMZx
hiak+BGj+wRmQhijvXHK9ooWyZzULf6k1VDcKdLqqOR9YkuhaljQvGNH5QvTxJHo
2B2kwZmd7/qLe3XqdBTqIY3PoD+kGlU8ldSuCEb+0h+8vdJSusfzDGg3tNnUyjco
EJnTTwUaYpK95YI4bvOOYmmMXmFkmiVCJpSi3tZ0/VDzE6RSryIi4wy7ySe2FPkK
VP4rFUlvUujLr/CT0O+Hu4jAPLhVUHH+9LUCUYPw+XEAfGXIHy8uBXyk7DJtEwaL
eClEY3sB/RxO3+G6gVj8P8LWjCJoTRx3MAA+tHwRPGd5BjxUHjfLd9qwkvB/ccTA
CtFE5fo4IfUOFuTPEEJMOfjEN1UzvMnN3UsUgq9yrQeR7ViU0Ygi/oXGjzPm9V+Q
d1R0oFb2liZ5E5WqaU9bZ6/G4hTKgaXHd9dXtJu4VDVCAlp2oY7hD+W8vL48XaeY
j/LpNa2l/VP5ad4bHjA1rytnQiG8asBVuropNB37x5A2qdq9gAxwzzSeNFPRjjYy
mD4ZnTptJKPjjo1QNSgEeHrOcm2NmNgY13DaVEUjBAOWK/ZZOBsJlWniYjpqbesY
h3aj8t/Krhaho5Ww90P521jUqzdTOxCM0rMTPLt7GHiRWSitBB60eNL5KjjERHGw
V4NiM7006sf+mJ7Bbopq3NbM6tjSWP81AyuAe4/vOGCZTpqxpPBLygUezL9z6YJ+
p2+ApQB2gh0HgduAKZ8sMPGpmNffDxpu7QkC9k3WOj2K2JKmzyzmV1rKcq0yeYYI
KipRspPeDfP9iS7o7KvXyO4LxrHsklGq/q8/lQiNEwIZC0IKduh/GC9j9EZK31vJ
ceBscIchwiK0g9QD8dey32R2g5MKZoK79f6mIMLoMfxbOjtOWisNWnKeMdQ4H3Bw
dTef4Cv3Lta5slM96pSPqbC3qcg3aKyjGOYOqU+dsPq13dIXNo2uziZcwvbwy1z7
cHy+daH9NjfV/1tRZZcGnYMkaVzTVBPAs9kG2Qg5u1GSfRbYHQZhAOBk2VSa90a6
9QsEmn/Ft0qu3b0+hPaRH1n4Zdrnx6TdoH91SqVqnfqKfkGoUfjsv9Bn2fQtFXMP
fphYkYXC025wAPJIQkl87yOhvWP/oNANR4dJvZCUx6wGk+ooWIsNQ2HgqAgEQ4QS
LXYlpPtFRqqZt4+uilwcowRhSZeQ0PPVM+zxqHb7mP1ae6MlSxZnis57ZDhzddix
edBwJzARf+bJ4YqXDcC1sZ4YdhaOGBAwoLbAD4YlmmwhU2cSZeZ/y+NiVW26C5wb
/n5B+9WOmmK0ZboK+oNuyy2tlpafJT1wWIajd+G5zi1iRep97e2sP/p52ZVtugaA
NI4LcG0ILqAnz2o+bN87g4Vs2OJ3TBMgGFnwrF4ehAP2KWYvWoEdz0pC+RYbJhIU
ijQQlBF2bk82J9UC4/lozB+oCrNbMbX8VM/J19N93FBuDLxWS1Gq+ywzSiJkSSj2
T6eeGESeBVNDmiD7EhGklrGkQGXOD1ZvAy2883PfLFdV6JQeCOcqCfQiy0eQpVnz
Fw2L8ZDkEmsIozzXQ9PaPUaKFHFaz7X6+RheOcLT5GWfaTcTCHecMIU2Gtef1vTZ
tvrQ3cXqv8qnYgHEksDKz9h4tosnNBg6FpsoiQhRHvnRQNMuKlyYu5Z1xyFx0acr
22X/lGvq3V8GSzMyRTJfjGMPZOXXyeqD8sn9gMNBbXji3CzHun/z7tlYFHs95Wxe
RPzKYN2GsL+hdS5NK3E+Tdfn+B+jYrMeNlNTl5YUigcTgKpMsLMXz0EqRMSJbU2b
jU2Eq2EvtR8Yw0zd5gOvcA9mfbnOAXQBdZnnabSPktzFcqlb1eQuDtxHpK/zrtYs
`protect END_PROTECTED
