`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AmmJWuQknWat2CQOfIMp413J5NxFczp1SHrCvx8N3apoz12/SUXAMzaj4vvLLAXb
MU8fCS+pKX4dPz8NZ8ZcUigwpOa38VirfEqM34owssgv7F9THKsvMUgEpjSzbYZ8
qijxmCeRVzsYUX5hw+J96r2d7R/lRy3TV71rnbnS4Tj/lVBr1I7RirbPyMfdUilC
SX5tSx7E2oFCSa0sCCjf4diKSYQBG9ppWG2EwqTHRsXJtrKwFH446q3Q4mtSHdaf
5SHI/BM/b4wyiQUXPSfnbTVReDyRtHYYhCNEufLG26d1IlS4Yblg5VwV/PFuRYx+
tXQM2HqXT+MHIoflGXncGauRF92WzW/Qbt8IJpiNVVceE4VilASXAzxEOV+5TnQ0
I4c2Uo3QHnFTq6urwOSCrA3mGMaMq6ezIJgO47iaaFuE2CAdmMMwTwxVL9r+c/TA
O/dNxAYnM56Cm+2nKhL9zlhXi+9u+/Lvk3vQXh/csH+4CkPrBRQRIS7DFHXfGaIU
6q8thd7mbYT3UJLxRWRpJBE2YQ/uJgg68pVUyM8zZUNI1gZtjqFNw1oV0LoVeVg2
44WZGP5TofaQ8Zi2hOBXdslF2zoEWeUgPMpcN8LERzGNeBzVkFkUj7eiT3m+j4XU
YW7Ul4B2vRtGqzR4GJkXqc3p9pY1gPlzSqtJb8qkXX0=
`protect END_PROTECTED
