`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cHYzpXA8SuITgTilzVhOV84MfGX44h012LYZEI3nrZnxrHuDW6/yHFFEKsx11lxP
6afHaol00G3zzcpoAGJYgq4VGjvw+Q6b/r2wkRBGekustPMHBcrTDeX1ijMx03lr
rVGh02JSfuHBVAMCX7VxPJcItZJ/RpaT3/nTKrRAZOuiToArdgSyN+Xm9PmzS/72
PQu/VnS5cgWokAZhOm3u2REfTXGJBHzyNBaXoXsJ0gTh9/VSeV5qC7RpylsKCyWo
ovT0pOszL/T9W0bPB4ezVbZoZDikK95Qcp8GxYTqaMdMnP0pUGnPcdahGvZOAJ7T
snI0MtAJQdIVQoor1NPeZyrMozrz3aacWaTrVUn86cEvtdUyBhjj19xxkPvnW1NW
7Wri+cuZpM6k04eZoEphEzqHxx0vtUnIzLd80onv1LtkfNkhE64LCTVJYOwu9qJ/
98FUWvLm5TEa5HZj7XPEKxXn4ZBYBLoVJqSHy/7DiAJj8zgQ0r6/cdcaqmfYRQBR
xS4zYAWNb3BsJlW783O4Q0RAgr53uecE91Dn0Hz6qiO2Mye4+iks+v3UIH2IMaC4
ep7gH0ow93n/WryPX16xPmXVjIO9kGNBOlnCc350h/GEEE++7YGqKBXc1c2VCNIm
AAJzpOxVNJ2/8Tw7Kq8CdxgP12yoFMc+Vy+/W12yX4oG17mpmiUJSR4DEZrwTA9+
pY4ZYK4L0iLWq/ooB9Rb43LRhv+5G5lvlDwsnSj9hRuoPkwm9rhoMPGHcaMXc9vY
72/peQ/QxE/DiQHf3aFI2Ljg9j6bmDy4g56WOn8tD7aTzobRgbzbzbGbqjDkbBs7
gMGOjwNTjFnM6hHgJhn121qrkHHKoDy5Oaq0HDjFhNsHcPGD/5NrmZjX9f2ZUskp
Ljd0t+k5xpBMlFcjGsGPBVC6DeTPMgNxPZvuizlZd7ThOL3BNI1GkmjSIONNVklT
VIkfMZYaiZD/7msooh9VKhUYr5hpl8PrwGjDBa2MgYNjOUrvCj17L9OXVYi8yXjm
AoaQdJFSXAr4kzs8UmFZR8sqKd8MIxc3mnwz8he+EW4zQdHUBH+zI5fU18MoSnFM
rzTyOYWWxllMgyo9PGwDPaJec+t4yKPC98jPpYj6A2NH+lQvbUCpifUcSYBePjka
+LGHSiTWZ7iJGDFt7JgUJYYluh13PX7084irGOpEvPE4F15Uupgt9pcYJhcZyEKy
6Ukadpq56tEwyEN+WbI3qA==
`protect END_PROTECTED
