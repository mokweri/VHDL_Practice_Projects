`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vf8DTQGmzn97AfWJGjJCt7g1T5uFlZg0yS1YHEpyEef6A0Es2SVj1aw1kycD9/7
iD5djyuk3NmZ1DwmoUyGQxJGdqoex5aQven4R2+ILxMsU1u+cOmEmWnSwh2PCK3Y
l17iKnQbbe8iHBB14nMNf7osY4M0a7Iav+/7VJMYUSrzyC33fUF7wzri9ZSmBR07
l1rrh8mJglu55jcmJBFFGK3lS2AyazROf6xb98zVZRISMytws9K1Du0Ylb1sYnzx
DVFHkDiDiFZ5/6J5H2a5h50xlLrGrcChE6BEk0u7/Zv5xvtw8Gdw7mvRXCzHJLYf
CRfdXp3NUD/amF8HIhyazex+4YFpU2yzRgH0PdW2KfnuEh3QOIWFJDwOI3TbxQHt
fCg6SzWu4hTypIljjF5O+LTjGnQ1Tlq8PILlUWITeoj7CJ0QNAY/nj6ldt24Nb92
EEBnlJvqRFjKFejApZ8zqNhchTLEpYDfrTd4MLnAgZV3MFyM2+cxdod86/kA+MKf
mwBKt/STjSgVtXBnRK+iGywxEgWhMy6kFuuzn17wTcQI5/eJaTMD1nk0o571V9h0
EYm52Qj5d4aPWaU7+F6Mh9bNsOgQZMoPgelarkZ3BJxjUWyHb/gvdR8ke0OwdZe6
1C3s/Mf2K2q240WwubpvvQ2YMJwuzF6PlUZq38MS1gHUDDxntWeyXg/s2SMKSVdG
UApotE4bQz1wTqVFcyjjq1vbsZsOOP55ly+A1pHUBgJweBPVhV5JYuhfmW01bcmH
uh+ChTVVRfWyn+c4N8RQnM5fHI6NXGiyuLdvL8ABZbFz94uRGGSKNqP0fIDW1pQf
NGsvpL/8zK0fspG3nVV8tDn5ZFMrXbsfrI0fAVnyBVuTML8ejwhupRei4PasY4gk
d5w3BJrHRp9TFrB/dPGmyuFbeyolZJX5ByogIwMWgcaB8REZ7VufLZ9dLjYn0oGN
zkTU4rlesGYZPYz21QXlq+AMzxwQ7uy3kTwOtvEXUC1Z/aVN3r+5E+mqylZaAIwn
jSEfzyC9FpF27nyp1vqEOiUoiSvpZMsRiwawpCdKy0A0wSpRUnhJ9XO0h5AQlHJF
xOq1Wy6abVsHuUm3VquHRjbkUi5DiJzfq9MdQ52qYgFflbMGYT5oY00KlAvdHvuG
75hL59tGw0QyPZAiDFLRiuzEgTjbwhFXEhbYZmsMAy2XhsbZUpkMC2cwHGp79Pfq
6lWB3N1/yXgnPlbNftX2Mcb+06/L5Q8kG3j0PvbtN6P/fN4xidBCngxlkLIgnVs2
wZv5II9H0yW+txvZh2od11w4GEgeMw+fIn2X2uFfdfkZr6SUkhchS59U6nvzr8NN
Qvq916jdZaG06RJRFy63ONhpDjsqGy2UFBCGO+2E8EWhw2t0UJnAgQFzY2VRJ6BM
KBeWmxoUmIvUfACX9LpSxRBWnrnsKhrs8LRWTjQd1p/10k5wcTrvtRO/X8kMz3Pi
xSzpBMaxBDXw+ctXA2pS/wBViMddsHdckjxzSkWkPvZbJbPoIQTA1nDjmkls4bEP
hbyRiVXaWm/UVqsADzcszZ8XOMPE/hlcwtyt17JHAdyINvgJstflo1iT3ypBCq5C
ARlH86j/nXekwZ1BMN6SPFJcYEEO/cNTEMLyA02w3iERqdb85DYRkumSPioxvgjX
oWRE7jMogIYtrxs5e4up95V16njGsCZb9Y4ZaW0Q+AqM8l8Kbg/h8N6tSoMAEvHZ
aTh9zzW7udwveQFQWbmSYhGvlQ7TSnyshXvGftSepfRZrQOWQNoplLFRgWRC/NIQ
AUNVqKNVGgM/a26MGZOSmNW1HyLgnYJdPzZPUtOnnhiCLeJJHzasK1hBjCx6PeQo
sPneJGETPOpY+2bO+6gE4otTyuj/NFXmbTIPn65J5tcD6CUwQL2PRim6wPQpPT/V
tYxC1NBsI7zGRmVO7ysC4n+47j5EA3fqVplBG25gvUPQ9szMichummNi4BqRmiOy
ycJuEMZ+hZTzpxqX1pK4MTgDoy37MweYdyfwoQEQZmaBnjtUJI/dR38lwX3rno5Z
wYMKoWa/yYj2FIqs/0RL6HyHfLCfWtV6MUiOrDlz7QQof3B6QVJ8UVTjoqfVd4zA
xvmXuRqMHB+VrtVTM7GOx7g0AJlY/pLNNk0FvnM6ntwR5jVpZax7k/f3MUtWT9OQ
5q5aATQxV9e5kx2UbGPRVU54O5yQ66vPmDQucth8vbGLyrIPhZ3daLslboFoiPyH
VfeuzV/SY/liIuIiYoHb2mG05ieVbPWlFmFSwQwwt8QSrUwDalyyPvyDEL8SrhO0
yyhWCMVlKux44ls/59gtLoK+hyJxk1ZXUGcbsT3ZzYqPi3cvgiSfrxEg+8rbsmeB
kAI1qaBdM8NxIxaL+8jTFTg8Stce1MgiYqSpYvyOADGAW67dqkgchwUVEhCJcZ6J
gx/KMaX6lxGxOck5Lw7P734Q4dWnjnVHPB2/EHCUc0w6ozo0/F6PR/AfksmJQHnQ
zGDQFuxM0xPF9uZ16v5snnGuNpIVg7/+BWL1Dzy8u3Qg8kR2KFRYaIbi8XNihI1b
ZTZuDSvnfGlPI11H9EWVyYlGyfh2WsQw2Bs5nB02dSBwcyNQMIyIEkERLIA0KI88
1SVr4/S7LJ8hVTkLkphb6uicrr4Zo7PrQHCbR+kWrQIWFRLPUIJ0Nsc9Ke5TboOF
H7VPUq0x3qfL37OBRD9/j3U7+IqKZv8muWk3sU5vIjUqneD24nfJKDYg3qSvlBG3
o9daF4gzFtg1wr7RQ1u/Xl+pE2RYJIz0ICOoQla5o9AHKQk07S8EwXgnxdbsRMKO
RsCGeMdmetbkVsn57nxnkS7B5tebllq+eRJWFln5W4cTxllspuZJGKDZxCkQKW86
+acmzhcvr2jXEmUOMdkfDnTI+/dsQuExyY2vPJN2UZM7wq2WPOq1O7Y//LPARZGI
9z2rOOOg7UhUY7U3iSYRQ3H7kMYT4Eoj/6mGH39orwchDfFe0FEk6J3+9yFQgykn
r7vi7HY6gWhlp2MqqGcy7WVz0dHkplfi/vklX2S8ws9yfTAxbki3eWOk44ArNlP5
wYbtzMH5+YJKUP9gjoZIEWgDeoBtBTQhXtl0veoxnBHCu9aVIHG43dy0K8aou+eg
DB6pW2Jzl3hTcFknqHAp+dqItYBaw0+GFDdGhQ5eiWczuoWA3k8ra7bATPZtI9TY
VIR7edgBzk6a8816eMJASKNIKu10XgvWZk7ze262p9KJqrTBw6JLic8CHh6sn4HQ
FrKEnwbYyTddDJ48f26qvDiLhpioAEKeql2eZLkp+7tVZV/Y+DfkRPUyuAPqomlu
xO7BCYaglgyXzUUWlAicYGnUa7q7m48ZjmSkBgZAgu+8m/bKumQQYqe/PIBGgDB5
9JF+OOb44XkUJa9eXx1RfE00l+mB1CMzGBkAhurOqN7hHC6H3QjB9QQYRtQg1RBt
Gr2Nvfm92jhp7BX3cV3Hd19OCysp76RPfdm9fToRPzPMHY7a6nfInWNbiVUo0i1L
aZ/EWU2h91nchFE1LJaw4LfjFFtpEz9Od7DjZgDbv3+MkBMXi25IKmuxRFvxhsT4
1drUazsultbBPV2dxv5wAG9eS+XmgioiO+Q+DkUQMWg54ug7XiYQGCCNzbIoTQAj
2VEdlXRRfXhbZcQ/NkbZyaCP6JELbnsyKiSUT/I2LvMwd3NZPXX7mLFmmDt932yO
ekkjoX/80LO2jg28zzA2Kdqp1F/XBT61nL3AVn2yyUI7oaJBFrzHXTpC97frxc14
/73BKRgbiaSiVtwuUjFNDkZy3ylEndx6SvlOpiEsiImUUOQFEdlMLoDNNflVZoX6
LSRujfVlgkGhC0dKJhYqtFpXRg/NuHe25c58jeO9kFieaC0g8zxy9Y1WTOJ4g7C5
z6vkTn7l+KYpnvQGRVT4f31KocIPTeVZeXVAB+7EdnNoHVzm/Q9U1ctXZZYlp0Vs
x/Ch1puzqu/HNopWKvPpIWnBS7E4UlqgBI1oHdQNMtMlqKsWuxC3q9rU7mKn2zw6
b43XCpEGIIxCi8n7a8DUtDTck+E0E9jrEjK3GEzf7zHz4GTkL1MCrVhzqyi97+Dm
ejC6bg2bH+2M6aNLNYGPPlisA+etx/z/Yte6+PXObiJWYbyQbl96d5hGKHs6fDPp
l+uy+pPuBg+t6oMk+rKJiFZWGqokUWNO/HActWsBsq8VQk5gFrSp872KhSdmnizN
QogpwcAwIvPTNMS67Rc6vTJH6HHLuWM3GQME6UJfy+AMYgm49Qgj7wV9pP5uPt9V
f7d5xnxvKi9i0an7XxXJvev2TKmcidhOwpZl/Jpskwlts1iyEhAsh/qNAQPikY4j
vREX2RPsIqUrRruHeWJDvHT6YgSOdTul5uNAmVzTINQwUWHmhK3S3+EJol8jr7eq
6yvoJ/MqysM1MzQDhnd4jQ9SWJyhJvdFcKBZXy4rA7JXQ1ZhYCEla1z4DZP5qS02
us6W3TIuDgpPi2hFuefh+Y4M/jgP9mewKP+7q7mnskxjqcsGRe2g7llM+DY0TWSX
qG0YgyqxlsY1AM+qroVt38ifQUxiF6Z3kvpVtxFeS2RVr2FqNcbZh616ph3guAcl
/oPx/z1xZx0G/LXjpi2+XA4WFeEZFURmnb6SA/wfOsLVMCgG5zorNTdKhW8/DehK
F65tW5xsZXfF/q4GyPDSrJaG5KVnjQqFG7zJY1EVdXVyp49VKZHDG1qHH5UX6fHg
othPGnoReVSR1rvLXNMuLGGdLAsOVaLrr2KTsjpgrn2mv6mB+DWwL9YseyG4MR+R
vdwAOTyV+eMBhHZBj1gl48c2gipl7wUyLpSTpoHvaXbRf2Sr9Nw9jhntAY5kmOd8
vB5149u8+XpGIdQUXCoN+N9cV6Ynp2V5Qk1aSBJ9xqb/W4a+dC8tB3+NANVZjLb7
1n1mkYuINUZHFBmeAg2ewCbwENRMr7nUcaJB4Z6CQ8sbC0MjU6XXaTaD7lbtx4ED
fY3M8t61kTHmnmeDzsLNtqb3cNQ7HTxUGJ9Rin11/n+pBRVQpLcw3HD8eALGjxkE
OfPO5iL+O0JvGWzK6EAGuQ4WDzdYydomNGAQVhsImIFrrp3CiJ9O4UlbI9r1mhhc
CjrL5jDwzO8p3MH59ZCgCyHCZHZdPdaJMnkK8VyVzGJJtiophbI2FLqh29xlNKON
HhquQeZgAI+HvWtvVF6UsHzl7kL2Oy1YFoE0vMlMo/ImJHIwLGifBzRVB4oaMeGZ
zB5KJW+Q64oF04APkBU38I1up0zRnXENQwdvVoNDMci95hpqxDmmbel1yP8HEfsC
ysGVD7xXdFPFLQY8pDeJ29GLfEpJO1fvJAZmzPhGfdMv+MYBK+UdvwINVhwrXI6g
39EnFxyxMzjWoNimqhb5hs/phso4Z0yITcnXd/9HvDNF0Qq8VBDq6JsrVoWuYUY7
CuJTDj+lEHv9R/XhLeEysR39QuwvD/FAPaa44n3Q94mgnrUaOgFVeWL2l9JXyjlZ
C8r/QlDXPqDHcLzvM7snscer+o+fFZWGiaaviXPuGQr9GF40WcnggSCfTZ2FFDoA
BYXufJmBhXgvdBxPxyyyXZjkZypCmG+HI8DxUgRWoEcBbnU2DxQGIKXuIEEeR08J
xGKAqIZIRccCE6PI1QRGbE1WOnvZxVYe9OT0J554XggL2blGLdjfSuMZx/0FF/oa
D1UmUWgG9V5oWWUl9szfRORk8+SoqvAF6CUxgW1FrJ99Di1T+YCsmZ/fvddEU2Ah
oWuLNcgvyQKurcByl5SylrNFpd0as537P3xwY/Sv9QlIbZxiw8pJRERc8dv8pl6x
iQvFb0wRCvK0OSSYGDqOfkA/FJnE4W1dfxqJei7b/zaPMo6LhrCnwN5/iftMQ9ob
0kmr10zJinbISZXb3mBGIIxTO3swT8tmNXZDDZZshrvVnCEvanp/aIQmsewoHPcZ
n6nZq2GvXCcPtDm1MfXNdjzcjEnY/Q6Ik/GX7ziNvPXy5PsoAId5Xv9gnlxPmDFQ
W/mS+9x75kmBU6H5pmpe6PvctEzsy++Y68s1ljr38ishA8p6BGwjdqEVqx1UXj/6
IdGUfpRX5s+8lMeIZu2A+2QZ8SEtFvECX3pQFrjXl74Xxe2C6EQVR2ErrR73mixA
P6KbC5FRl/JNvxzs9Fr0uBk5K8hRHuMKgHZ998ravjFUWod5ACsIeBt63y00AD9w
48kgOf0VzC7Os+CS4EY7cP1r5m51c7Aer4oAgwrawhLtyyEZKCPEPzj3Nu2dJkEY
K7MrbOLm6a3a9c32u8Vd2P26tP1QgcyVxHJuiBJtz80IEuuFQbyTu79ZEdnOZEx8
yplLHtdkOKqp8+5kMwYnRYL56XqXcf2MB7sFcrQo64CbvCdPRMtW0x/Veq/NU30L
82qz8vDrvQrqpbYM1Ve/rFZ2tZm5ko2kQz9+dJEk7Ktj9O/vQDubQX+/ZSIwl1mS
6VSR6HIwllTm0ECel6tl4xIinOLOZkSa50wtGoMFtNJgO8udruUwAHNa1VlAdVZ6
CJZtV7JxnrcIX8TIY3DRPoJlWBk8YMNkzeHuoNm5GANVB4vGsCGmX47D0bjl7OXl
YBUKIytu124A/U2hnJRQRRc3+GstQeJn3JI6LHmEnGyrD2EVZNKlMyrZ0vha5VZ/
f6RtySOpZEqAr9bn9P1CPLzw3kCmgJjUzPO1dFf10Gr82y+s1fNg3vrewr+HEoTh
THB/O3VPD6nPxxmykeOltHOf717SjJJi2J5hMruYQH0M7qaHsfJBl2U7SeehpO9j
qLgbQCzHwZbHRWHIHaj4k73PkGqOnfSpp8lDhdhvneEk4P6j59uYNxU1W+i75Mc6
v3cWaTeT84v7brSxDX2Yfqj1PcmvnvVEjn3G76nsSafVkYw8VT1egzNFL0q9+GMp
lr/8uPRWPVIRozcF0u54EO90T6q2tjsvXBXjfIA5xjd9+hnrV+UKeIOgGQco4PGF
bldXVNIRf4Rak8EeBH1j/lHDGn2knzk4JAJWQQZFcQhuFkmQcyaXISTKP6SRcx+O
xiWQvsuXSmdy4fRpMaX+L5XkBNP4b3iVl3PtQSGgA0QAD47T+c6gdYEvI+jujEAv
+IjpLVPHIq7Wv6fabTc69awb4h31BTJH+XxXcU/8sW/xBNGXUkw29+WxG5yRDZAE
4nNM4PgK5uERE/GN4b+FVAw25FG9qKjl9InfFCEJNA2JPgjK1bdRBW3zogiChLpx
NDFof/gg5Jc0P6GpwzbqzMiwqk9zLPZ0SfgMho9XICuxUR/3SNShwsPfk+XwPkfM
DavQnkzprHVrQZehPNVn1AZ46E3luJiV81WAvCfQD78xcZHZ/ZhYZ2kNzHPR0gtQ
lO+mgvHl1wRCBPMEGC6yfXWeeEY8RjltG3uIGgk+0Bl8UOrb9X9+8JtMRVUGhksD
t6MsLfD2ubvuXHot2U67HPaNndYv2hMWL0rgr9GX06g1CE2QnIu5Rd44vtFIRpwo
L7Le/fyLM+vZXzLL5nQtpwKj5/qbjtu+PBA5Y5JHDY/voEF6JwJExOT03eU8ZLJ6
AQRn1prOdWA7D5lE0LPkUusKjqiDrC9GUH/pyk99gN72IHiIQe7e+6w1NfD8PS3q
rCQU18DPvwKMSYV64i1JQ+blWr0MF3WAjxOnuyKeoZozOG1sI7nQq22/HHrD0FOd
JwXnuUkc3cJzgBDiSsUqTVkMxbJqQH6kJqkAx6s/q6Vd7kp/KLca2issSqESjW16
z70Ax5KVJ8kLeCX/M7/KhIIq4vwQprzXHZB/Tr7rFmnJYQDpslUdBC5v8+Jxs7jG
0YzPk5zjIu20owDfTXcRzYiUV5zhj0XYqzS5OpL6u/O8Gi5+fC9uYDtNNfSZM4sE
LQPipw6KLPA69ELHCCEC3amJ0n2OXQ03ohOuk+2zjltSPuSNpPuPbY8QgeXuw6ji
zJH7ff6gc3tulztlkRg7TJlEEK0BicZdMDOFgVnTKu5hS9TR81qMQXgpvZWEDQ0J
vIVuS6OhSlvRrKowqw/xtY8hmHKGz0mAPaOqwWs7RVntCnnVoVMQfSHN98sRub2y
BGUFeftIbLWsuYI5NrzmfkXfP8rFuBt7QzpcblhErWWD1I+EL4/K+DxtKYf1qpGN
5hyu4Vo+vP85u+9nDcIim0vrkXLBz7afPCTB6c2SnUE29xUNAr3mqAwdo0dPg7Bs
Gqtflb3Zgc0P0qd0t/u74SP8d6a5mjBkVV8BXGqGf84xuxwzFi8GGUGBYD++DUyI
bP/9h69mcd67/1jBpDyzm5ZNI/WAlEXyjq4PlHkrBj+KVxwUHJjZXFLdZrvSEyqD
zSF4dPLEowQBs982W2f8qSrMvTbd/eFadgUz+08WbxgLUL97G+i3RRe05AXaaOKC
H0mJtensEMFgf3WI1wvLIVvEUHaFVGNhqjXxoDc1QVx72NQ1R84il+BCMWywpysL
iWGP7D87kRPhcBsnDnw/mOFW9bjhACm4tbjscxb2X0AFSodSwEnzVecujmv//44k
9Dm0uMfce9c3lJVfsxXHhfRCE2OjT8u3syIVd2VHHt+NYmOO6sy5Y7q3/OxFeFql
bU3ybn4RPeWlcqEaUcH84PAtqxTpOXMqr1jxFxx01wUQpIEQWJ+fiKO+5GEA6bc5
Rh4eFUKeiQtJVlQEzLkt4e/1FW4rROtOJ/iRhxpmfMR/BsTVXhHjtA/YC9sSjEo2
h5aMmxPsb2Tgn2+lnBQTVPGZMWW2Mv+5D+7FLB+hNetoyhEnikvjUZtCsrUXR7jD
ceAL+xB2Zbrd+McAci/HYoviA+FikpMgLvKFdvt0dnvWEMF9i2NTU1XwBTwcYlmn
L61xYl/w6zlRmSwGMfiXTTnVFQuOf3gkAKIdu8N+xRHWoqBj3VCPhoB3kKsFLkQK
Bas5t1b3Nr4m3ihp02UtxKAEQ6R0DsqHZ1bkjsfJoFRRF2Mq0shbR23v6nbyiSEe
7eiqfng1GqNEP3XtOP4IAmPUhf1Jo/1aViqkag8ASWP/Wn4vIy2c20ogOApQ+r3u
oHKgzhER4Ur89hgk7JbSpwP8yVftKUbLg69wVnSyEY7Rk5GTT5YPzUKnqUvC2LOh
bL5mD7o0QmQfQsO7seyQ+T/PGU++W9rdBNUHgtberb2Ojf/LiUfTlJG8+3H/MFN+
MTb7g5knQGo1S9U1gAI/k1MfUZaXpmU2VjJyMo00GOnUFtAC6WFSveGkA/C9feyA
6Kvxz0nLOZYJHw8DG6jFeqOsHQjDzkN0W1mOnBh6xKwtCyfyiO2pIDz0LuPck3u2
nCpur4nuIMXHEvmL8kzd9TxSLPsel+UgM+LiX19eJ6smsXd4G0TJypi1UoiW6f7z
Il9vtuTXIav4oWDoqdiBMnBQyF5nUpIeUS9/h5TRSSKLO55QERX+I28Me/o2S0rp
XdshrVYU57f4M+jcnxubbQ6GWETlUZmT11m1uVQxzjIbpTTW3Coy/wqGgbJP+3nv
itYStl1ook99oZMovfKqrAsEZpKFEhoSFzxHOR4k2cGJNowJGfLUlVmbKcrvWm6z
vp5T+iu1f13K9xAvR1weABl67uiLVgqKLRiGNNzc0vbU6Nrz8kg2bn04ygT1fGcJ
ZGtuE4OEvxHPEZ6oc8/v7AyTYhcLS/Doz153yyt7WXVPaXuurZH4mKRT+oCtk8pO
x6oFwTce1iPzi2odXgRSJ6nQmxIfiKcXW+rnjL2Pah4NFghbHXHHl5gFRagW2Mnl
F49m41hJDdEIRLWOOmIJR6MCL7POVunV4bqP0/fdd+IDLz+uqfana2sc7C6LGeBs
33UytNqPZrDA34aV35dsagINm0NWnaeLgxFZYNrYjsvg3Zv9mHcR7QPiwsnVLxQU
b38CwgdeIfaLDezKwBir9Rs97w1icjODYM7rHFxWkaW6HbF92G5NIMV0QegzK09R
SugMaMLFlarMTx6j6na1zmiyKBRXEtkAP2zCUWYBEqdqVr7NqIVoAXqXSntihtEq
ayPVPJkyKpfMTpJqDwYkgecKNEnq6btPylDx2NxGcDMdwljtshvhECeGa7p73Y2p
lQazTj/wEofTg8l5ee93yMPIWSIhRaTtoJbIgh9CCqPZuk3g+R0pwM5l5gVcAeFT
FMNPFLcda7VAJgTOks26g4CcUs4o0xfNx/NqN4yjU8mJ7oyXCGXhgUH2+WSUIQi4
cISi5QiKsoDuJxg9xHPa0eKG9z82/3Yp3T2BcQrT1UNxmWeS7NY+Aa1FBcvKKeCF
1dYLSJH1SiHH8ZtKexd4M9/WS9/wcGJp+akvS6en1yGk+0EMV3Mvt6stJvMzNCIG
Hu6ERHoLjDW3MJa0rJEuqpaZihUMw4T6Ur/is3JxCffmaVaih8aRoWPK/ci4Pyx0
qzk0ZWsn3JFUoj0hfph6y0hQfA/f7LJhh6Z0FKJ12VHWcCk6JKWTcRUy94oItkWe
kdj4YoOj/iWwlrw4ZqpX0GTs2pickm9k4Kr3oW0uuO/8SNfB2YwiSke/iVBUJ/0X
6y1YquVJxm2ipsjVYigvoSt/1DVThi1smmbVswaM2bF+GJyqAF+mOA75VcyeSpEI
dEhgMxuGQvMK42kkBUzc6vp1B9vXZ9+Yi/rHcDYoGae+tSW1SC9SLcd3fMdiEZwM
PEHru44LKn0XeNyqp1RTbFYf1qK3jlhPxUCy+AsIBTg/MY8iUfG08K7UzgzJ1V9W
21eFasKgoLbtGeOUXyJZYvmspXolUIC3VGObOxiMhyevNhQ0UJ1YBlFH68h/b90I
MMyUQK/D2Zb7/np3r/MMFgvDvnxX9ikBBrh7KDYRLRWEZYOxQ7feXbT/namTFYsW
LDRc9d+TqHXdSTNFPhifuHWauTHD/FtxtrKvkl5z3eKdItbJPFfAXImEQawt3n2D
3/V2NGXv/2kV0MqLu0YbMFSc+TzQAV0ah4YduYFb63R1iPW5BWHA2wlbwdgENjw9
xwpMF0wfT761NKzYvcE40M1x7xVdfNBGQNIoUJh2098E4JuUxc+0wJEF0Oa98/40
io9Fyg75ksSLxtufse9abCQxfEC257ZLW6Zqoc3AGKEVXcaUARTjies1iFVbe4AI
R4rp3LhoUQxpYaX3JR0TV/LnJ/9QwLvCp4FrP3aopXqF/0y8l0PlPAr9i2IRo9XH
d1+jh8dHHW/ne+HtP8Xl6tL90DWoE+eAezq6r1a+UF4Tq9974vUpVVLJndJ25DRU
HBwRPA9jMeHEJhA9eBePEZNy96+wXdJRJVGUeHSP+uLjqHEEgBKiLrvxxNW3qRWB
NmU/AtMANWI5jCBDkHNVS4aAnnujyORWzJJDL9qgiUteV4f2OitX1j3hoSDZXTzt
QvWMMSpQxuji0wRiug2smXMxgpG7fEBY11N0r9obSYCoCLdu2PnNjV8fxXyq/t65
hw9JPAO4hkrO3MDPfcibYs+JbpqIAZd4BRmb9ebeA9bg3VQxL2Wvtcl/4hfOsPRN
I5/6QkaVl53xHt9iQzzMy5lPwae5vnS2z3lBrCbUSdbVMkDyHJbIU46v69QhuC/V
EXjoDRidqfN579Zr0dGXgnxOwag6R2I40YYfrX2Wfc4nAjB1j6kvsWGErU7hFgF5
6qZHhbHd1Zf1DPKvq5/1n0QpVwvJTHtcEhhrEOuUderladMhxdu232N58lku7KUW
x8S4mByGshcgN+Vx9JgX6beF7xjJFlP6JtGZB5XNBZ09wBqxcivY1cvln8HbJ5Ey
yQTvVvJyxW/J5NlpuCsIl9XpNFwacR492ibh9IjrxQpq0ckVya0KTq7+c3KA+PTx
i0CVCHZE3TafraRevrLeaMbh/5rbvM62kMjGj/zmJuSzvBQjUM/7HJOt2UKEARgb
XqxWGP6J/qF6xmGy+SMJG5LhoOZaNd85mTVKx6A4bRDr5nAjHoYwYM9BRgpVET+j
qhtv6WJR4GhZJzWyihAr8yFrcxFhdjl2f1bJ5Z0AoBDP2s4lD73ISUNeAgW+xVfh
G+GKSUdx9ebSyaiRVAgOjx9kJWkyMcnMqyjVrBlvWGyUH0V/Ryro3H9UVa13enMy
2DaKzYpX4Blt53lkdAzzW7Jyxi65bXI1IN9DSWsv7CVSJctAHSl2JUH6fJ6dUhz7
MMHG2Uf+lNP6IQMMLkyKqJrOfpaD3GEm1maMvELbP6rqtTMaqw0iBFUNtTgpBp6k
IfDls/DRWkkn1H8LzZ1PEPpm539BzN0KbEoIdDCNBVSIoaS037duWvIbM1tWSXJe
uevEDADc+NbqGse1o96rydr0UuGzBcJT9RWQ/fIexVwPlt1/ja14nzflMriYI7tI
3920JebcEb+5Q9vzIGLg8s+1AAewHbnymUvikuWbq34/x+dDUgS/29k1cTkuUDh+
uQ+nTEO2W4x0Rob6SC3SX39UHCPfL9f6nU3i8Xu4pncBDrJ0SzI9P/UkVuOab8LM
XWYaG27LVFScdwpG6LLqBXqEqCu35BdhxWGabbnhRAvLDQ1LrJ+jIoCcj7nVkRKp
jV5lEpjWcE/KKRXn0chx9+le20cHmryL08BjmZCKQxqrN4ccJxjKMNQDTfc73at1
Xjhp5sr0SBPg49mi9JuJgRwgJzO91RIY84kgUx+elIIBaGFcjceITRkEypsHmxcg
FJLm5hpcBtAH8F6G7FA85tkwYa/2nF2e9AN74RTABrOobIODG7oqHcrGPYe/tdXv
zDNAcQ5MvZ37WwY4Fufp3jWP3xkgJ+mZ+seE27HD6Ur6TG56fJDgXKUPAjd0bWFY
Z1rH3Cx/jf1MOVZqH6yQJ4qg6ZgCtkFWPU7Cji8HWnVXEyEW2jCqtJlITSEMfvQM
Ucqbl0q/nZ8u6k5zu7B9VhHoAbuGfKOz6fYRT2O9X+Yvfo94hgW5NpPvsFK7GlXf
Tdpo/inND4ruWKabab5rTdkvoQXsoiHnOMZVdmkWDkykaLZFTlMnAXwNV709bH9B
OuPtpXxOwmRwYdo4VV668bYmJRnGcT9OWE+H1HtbFdrTBt3Lx5SMaDdb2ljna0IK
/p8EHghHWa/MD7u5NloFVdzgnLnnHEDuIF9D3dNkBvqP9N1JZ6d2LUIwv2DHd4I0
C7ywhHGsx2B5MRv3qU0fcU2xPuB+9Yrm6qTE/z7xApJPOF/Mqo7pqtgKqC00pxnL
Z8eY4VlVBSFeNnxwZnCNrBxeJc5y0rQVKM2rc0clXbniAS8nlg3ZsPUWDn+UCgA4
2ppxexEqU7vg4TyDq0GYdAQLerP2D2piW/I118dC2O3thF67DtxM97Vk3fthkQDf
WRtgDKtv/y5nGojOSiHxa5LkPu/FP0CNMgGCCda5CjpnLJGWDgD7Us8YK46H17IM
fMk/b12QlFaQv9BYjLKHz3Y3scDKFs3MvsFM6bU/LyL8vcZYFH/5jpnu810OM8NX
D1ZVn5Dr/g0szfDjLfD6lHA8q62KTy8/79rRzRwPV9yq/hFMgPin7KtRMGa5Z4ul
V2SMXppQgubw6879TyKblBR0/LIyqmil4E+scU+TUDdSTpLzGiEmTaumthYyyZ/c
6kYn/lyyklAbdjnBt7EzwpqdJ/9ylsdRXEsJvtUN+LdzL4Vphse7RKGB/1aVr0m2
IPa0Wdk7P9xY85l4xLENaRE52QEizAFz62GzkUzCIfWpHnitmGlfv45Ep505x1xC
uhXJk1EJ0CctpIztcpg6aiw1XvoyWWAU9p71jUbeFbj/LF+JVVenMqIiCjzoGbiN
lMkMhPtU6izG2bdtgIRkxuE60XtUuV3Hrrwq4fSK7LEGX7HkUakkG1AgTNvBsa6/
ffhQjn0UzZwhOTLQqQV1Hx65KmG9MJzl9xhirQKOmR23JbHm46+N6IQ+Fim5aQaJ
A6DyWw7moaH5YDbQJvLjsH1NdPUFkspV59hwIKgdF5KZdkp3jMgcOUOpITJXUdYB
/Akpu1F5cE5IA5H4ODLKfM11S4LQIcQLO4+05F16DoU0naC86kqYYuDHRKSD8LA6
WmHdOnkc+aVyAb6cJynfbocamGuiPflLtomisJIMkTQp/UrdUq2PgJ0uu7n6eI5h
HVUhJiHXYGuTMGOdeOEt6aAss3j8o9KT9djM/ZwG4nDGplVxMMO8C8H8BBMYg7Gv
tVVsSjZR+GmKG88xF5NPX45puOru14p5126p8vSmdYP48WEDXBQL6uk794v1OlBU
QDRtL9G4g6Kj6FGt33iFI1E3RGPDGKkchVuyXi5GH1ILBkD6sSWEPpGFjcWSZprD
w2zlBSPLgNt65yNuP+GVUAIHIQ+2lRDFHno/iBpkiBnLwuAw8mwnWSU1mYvY9mIh
OQupXFdDEYpV69FL6X8Da4Uz2um9AffnpfhqKcPZzH0t0fknzVhEnds807LkD0S3
62DHZ3cl5ePM7wpH82Kvi7hFzxe2cS7xHR17wc0/aBEKxJg0Yl6PzfE8oD65gFg5
DF6D5EUpfo7Of98wUmztFFZ3uSVuAcGupU68VQVqx4hvhEw2ldFTb4q0ebxXmWlL
oQFd+FtPk8hHZSSj+m9sDSlCqjiEOI0FNwlcrGySMtlcUzfq06vFJe0PW24PGlcf
JUvBrg3wxhbKzTpePhOvMp7cSe0yRG2gB4gEqVvd4CCpYS6t4c9Rv/qPCQB8vgYE
oaaQzpx0Ppx+lkgKdCW7ZOBCHy33osz2Vm59durDRqcDMEqq0XSIH+zVxfxYkJwj
hSNeOvij2SuMchFyirMoyx1E3B6NpXQiTMkox+S6wxGu1m/5JcqhGjZaST0J/d4Q
iNJ88OefubNmMCmMQksH/Pu/yqXaunBA2v540xlez7X9Kiqh46o333C3MluCgkTb
8uljJxcrk/35rs8Z2IjtGKWW9N7S87Pp7210OI+Novild2yaZRTZQQr2j3SgHecO
wjrQaHPIpns6a1n0Kd5ZxwIs+l2NqnZkWTEtGtqEF11lexFG5uOgU2/XpHOdb9P0
6rvfLtwXvMQ98f7BNh7j5dTEEdEKg1Vdu+LulmLnRyTELVpUD1DkFcqeqLoyAXnR
vrqbP3MC8x4Bki1ac/OGw/p5rXKgWvwNSMCptu6NG7dqk3L3RzCeL69uZrNLJMIl
ZTKMiVAYdCvN7HkgKoYqe9y7MVdEAHWZKBIrDVZeYhCf3IH12Ahe/0ROZbHRgo3l
7kIWntpikXNU6vqTt9BRBQsuqEgsU8e8d4ydHGLdHelKOeRmtKm/CL0vkIXmi1+Q
G5fOGr21oh2OPxIIqKo68hZvQC7MXhCpxM7ucgIWfV9ETpEvkOD+x+LQ27Wk/9SJ
f/qTEgAyQ/ZYaT2DnukkSfAgofGKFbxxK9f2Ncq8ISu4MVDTFxUJX1nrAoxNAymY
VmkFRLcDMipPYoN4ar/1odNYGCom5ZZI0RQYSkguvtgA1w7V4VQvaloK6Kn/pv5x
lx66lsS4uqCosGvjfpn8UgUmHd3dRG7KXHHct+Y5EjTluwz7ysr3RFhrSwMNpEaM
B5gk2EyaZRZhtuXXHrKRsgUmNfjFXe0m1BIrT9UaX7YF4s4RGeVj2gtfyzagx7cZ
TVY7MP60eGjAjdeufQcVokL3HiGWQwddQ6fNaz/ddfzzSicFt4e7MZT1rrCNPu+l
rou3LC9eDbFqE87TnHDddYx5rVscXkVzYE60oCxZvqhT0CGV8cvyjZFAcrnT260U
KZHE4AKzWSfotUNXKnHU9/xYmaokHk1M8/Q09+D4pahszJj4cNW0wWyub2YIKcNg
N31812BNIRSjOkxWjSxsbrgOjhkz56zUWNucfdWFegfDzQ4/Bcn5SubyYt9Clej4
bGM0yTE3A491O8YniLUVCnPweFiN7clby7e+dqRaFNc902fa2rF1ykVtLKNDzx+N
74tN3XXT45TKqYgPJRcVDJd+ZA3irRt3XwpOaO8ZZ88ZggL2OL4puFpjWop55hOF
HqEOuG7NNf59HCf8UNhzydXXLP79u89YUHCWmEqzTnC5SKswecVKx4PfjjJpuk0L
XpwQQIZ0ZTfbVcSdzU8SJiyBBY1vrtcImMa0Jf1EuJgdK8ljrOaVi0PPquosMRQu
R9OKDYuZA4RO5+t3KFu5ulYLt1vYRw2MaHst6j7xOMdbQ9FofwudA90V0pgAuXAy
VYSovA6xHZWz+BsJmH88lMDDXEKtNtsyRhGk5btCvKp+RqtFlJNyEB7ZVqjOvBmN
jUCmSQ7gAIHyMI4o4wUslwCdfJHSQ+PgkaXV7Y9GAyM5RcBFIvXs+5CzOazXHzeg
Qu4Edue4uwR9vsa61eiT1gnmGgenA9hhIpp9cqfmQG0ZIQzIYOKlm9fa/aUP1AUv
R+D55BeU2nh+dl27WBcTe7ai3oOQltQpTcfMMqo/GKPdnLVY8HamwsD5CkffR+8d
6QReNjCw6uQByMcugE2OFfQGLtHeO/stG/8UE02h9pOaymNTvncNa6+S4ZnnaTES
nwyzhQNHsy85YnJ+0TuMaTDQ+ZZPPbDz+5XDoeOyjQx7fWg7mNXKHuKmAnkfF+KN
suxV6YzNZo6F5RDrb6I5S+Nbp2fafTSvyX1q6W9g2beRsLU80QFXUaVfGywkhWvr
/jQmdV44MdDomTYEE7Xx9N9R1NMVYpaO07SlZOpxikLuXX+DPoomMwKaU7ymMR/E
QfWzlo312emYu1p3VcxQTj/haQuT0U/kGlrOlvUwHcyZMuDBOraAUdg3uLC2yqpE
A9sfi1Ew4vjRyHZZDXHQp/9F9Y4c+qj2+9LKid7An/PyBOq3UuNz2vNAQrjeXbDl
PYceHGllLBg5ZrOWHEWudIIvu7gq4/Bi6JQ7Y0RykKpZcvuej4r67gmRNURF/GJp
p4RSoPaF/jaE/RaWdd5vl5ZlvCJhjM6E1uwicgs7he7IiZC4r985Qu0uVfR52Nnt
wwam7FEDwIIRMduYGsVotIWWpMjarc4c72yIwqGr43CURTKFDIyL2nvBeZwgseoB
mzsjQlMIewFste87WHflD3xtPXR+pRDnPE75GR45xZ0LMrjWqGdokAdhM8qA9Gw9
0lwWbRg1cjlySyyQy9DaXzxOTYYsfehWx3FTO7/7tIi27r7UHAgUKs9dMP+9cDv5
0D3M6gSVQtNR116vmqgSqLIitdQf5wR3kiJ0FkAU6VTfKbAquAci6xqFf/yWCY/3
fBVioWUh3k+yOZPXBM8lKvcLWZb5HxefPlVrAwflTPMBNIlwQhRkg94jTIEloWff
xnChdnTUItQVXQj9Z3OPri+Z1YNWUvt0kVq0cI5SrKYdOmjZwzgE/Q4PKBQFNgJV
Yz+O+O8cs266WvsjSvBn//D9jTNLPsWifPoJ6S7nGKtmro8pRziD937Glp39BU6P
JJ+UR4Gfu0WARxgtlyZfeIW4YC/hzVqrPUM5kmsFvqtbd52ZGrC4QVv0emk6igAt
Nwdj8TPSOUVk/GArAt3rk4nmYf+YK9sfowCp4TPOYvQbJocCEzADbv+Dgctdo1Du
gFwMwcTb/8oB0x5ZOYSjfBcybrjsWMlfsgHxp1f69fmkVfqD30j35DTjEGE0X4yx
VotUlJS4JkVex3QrOv9+q8w49a/CRPG2qX1Wk3PkIpFTPsTNNvwo48su8RKhUwh7
zssNLAueK8FZCd1wrEtu3Y7dMxr8hy32VSdEEwbcaAii+pWzn3MMRF8bEM6S+Msk
/ZICyQ/Jhj7V+Lorh3WrPgl8VOrxZLwHRANTOGSq7NRop14sdoWFYTFWyPTyOsON
vIqzl1fKC6e1POYzQhrb9RSfuKXz6uqcLbjBy6JMv1F43fq86bfrfTQZVFw6LAGc
NoIU8GrBacPiefuCLDIUBOorZJqCWEAf7Jdu9KpfIQuXy/+5Y2fY5Lae/gBx6CPy
4jGgCo+6MtrhxlPDMDdpsYOggCPu1hUiOm3POI3SKJtVSGPq6gLfcBUya1zq03+s
ER93vHkUKWHwd449fut30BAWwckc5n0WG1r2A8HFaeawu++2wdhgYfySYsY2zcvu
wVWT3Hm3TSgmQlxoveiV5GiAq+flnRB1bSR2HzyLR8/YwiI87QWkZHLfhiur3QNq
y/z71NkEbqWNA3j/0wIWOP462nJ/qv3uAXTm8MN77rMHSi+8ts9k5IXSJcWvdBWr
a1JJrsPRVxJCDRcCc803V9l+8yXF9nh9orf+EpF93M3RDeIAgdSEIGgFa5LvZd69
E4r9kC/oNVajJ8HqknKj4xB5zIkB4JIv2MCJiuyQF3A7K3bAa8SkApkUXZOYxePK
Ri9sF66kV2xdp9Pj7tLTsrguvOvhw6j6LDaZvf+a7ks4qOMD+PinKa9ouYFJO1hw
MSJ3GI9RRcahNUCzxA8XdbbDyeX2rTBP5NF7ER7kMdLCZM+nPyOyZfR1xFGdy3qS
ZrNvXJh+phZ3K6beAjMsEeA0zuo/Qzhvn1UP/cbN5BXjgDyEIYTUD4qQqYFHCok9
ks+ti8/9AU3NEQQHckUn1H4o1plyx3/FYO/B1pcAaRUnsv9XRZnUOT7Zr6NpTKmC
1lZttwHiUbyW5iiJfyCWDYdFX685V95Ax3FTp6yBDcLtty9x45Sp1M2WuA3eSMHd
A9yI1kT+rR+LYvhbtgDSQNTp8Ry8JuC4v9ao/4XIHQn+v+xHr+W2k2RMaqtTnCUl
F+YtiLa0xmQ2p/JVeoCRYVpTTiZsNFfJzL0EAjA7LMWbzNe7LjNpAH67DyelUlLC
fwIobyiEGFS4Ak6xl1RdOskVuRcafog8gPdnu//t0NwmKGEfszzgKf+orGP5DNAn
FuUTHyi3Rc+aD+NzvDBsjzhXc88PSWlwLowNdPy9rKo1fNIl2LRpq5eXV7e1o4au
0PBktok6+/pUbp7vEtrYJq7Nx7nOrOov+o0QNHjEigqZANpo3HjNxKbWdLc3gEUZ
VCuv+uHDPUQwACSXSjnNpSCC3qaNEaTPWMLzGpDwRKFPRu1FROHCus/x2/yhDhg8
+fuvXLeYccqaLWIBbCVoXChM1VhkqrU3nmUBPmfFWtV/D89KI3iNASfyeCSsyhT0
zZBPEmz+fmThL6KWHk/wOgEPaThxz9w5xQOr6ioxYmpxJoeY9MC7kdytN/ZJDKJl
RJzwwTsuAunaAmBO8PKJ1PQGylnCAfOJKzDeNyI4POAtxZ4B954DGuWFIod2c5+s
RsjKo6Yan6COmf8RhoViN6S7DVkjvXzS0EMCBem8Ych1nFz8cbVkQPL4vu9/VX4s
jRQfsJSwOcNGqeeQEvssJ59g6+WNmOvAMd7b/UKR9YcXU+SnJwM5GTJo6tTHtUUs
LiPM7yKBVW6CtQCWorJS2IOuXP6rkz6Q6WQsWzw6usT5MOk8UuvDfu5DKmAfbPSt
PjYq4bIb5In/hcOCQcDFWTM0SylhDsWvip5vBC2AhKR4zmGObwmS1kSmYY+QRaz0
U3uGn0t/+0LjMQ/q0BI6lBEaR2ZQdG5xraEFxP7zxz3vcEFkuI4Ozv3S1StZjLHC
AeE/XDmc2YvQPpho1UsAm53Wee0CjLSHUuPXwcovNpmXMwG92O/1vdtfQq7nFmyy
KRJqhZnHw6snnQZPI/HQqOnWZGt8Evh8WJR1WfteH/R+Lrr7f8ZNcMWelLi1hZn2
VxW1dbzgwFuRdJFJbSf2ip/AWQe03s1jU4eyp4xq2gqN1WNPU67Oxq8XJntPcaXe
j1nsewuhg7uEORWR+hm43msvU/PKq1uEdy8TcJMAffEVyRZ8t860zBeK68Il7J/C
xjJ4pAaCgm2+A89sEqsVpMFVuu/QwTnmK4kNT9anvryQ/YtTBOnGGM2R0akchtOX
sguJINIjz3RbMVfUVqu+0zD+ctlzVcp1FdAViR3K6U3Fylk/+svrpW83VhELe2qy
EGX84+Ex7vcMltbDzEhbE/0cVYVcJPwapCS9J0PFH8ioxHQdQTZChJaFYUgUpzj0
NR22r43csWRq2LosDP3YHcQS11JjLDoQ5wi+BnO75SMCldPNUHsLWAGukAl/9iwG
T71BCGYZ6uDLuDO5XZtXrXHBoVoajEgtjt3k1k6btTeqrhqXpbkspvvdakHrpyuS
kvgvzIcPuVsgNnN+ZdKNmWthOmufOiwKJfxKMoDbT7mYg5yqFthI2bWojkNO2Q++
AQHbg+JI1Ili4DHeHaU59A9HdZc8XbR0+FsRaPBcK/oQytXVUt+1jR8cgOdmoBjJ
ltXVUaCAQYjAs6u8ie1IoNtrNgnpL+jCkmJcYAfCsJiG2iLpCcXHh1b3bVSX1vKa
0Urm1bEwdJyVziThn+lsJdvBLRu8nsJT/KZVEO64/t7+8sOPIrHUSAlXye7JTw1B
Xli6KWzWsje9I8bBPj/i+reVCnJ/saUlCPvICoHNZOoUItWmfIVZ90UQZQRWjyVw
mvF2gUIKZs4wgDgXooB4tZ2h99VsSSiWx/gJpCjLbhtEbtpxFov61+ihiyaVsQao
mAJb7J5CTxfVPZZFmIrEry5JvHANxFmwEJ4IzYlwRuIiCFe6rtLq2GmEU441nfHW
FxwftYpjS05sVRg15lScfP2odaXCY7KfJ3eaRgrPBdqN0X3QXk1ehdwHtYUVL+ci
eJHlt9vEGDcPUHBdWbYE09NgFtccYfwjkmlSmKyGeb1eAaC1bVAirhIXLasI5E4n
rR1X7mQdhJYmDQM97x81Vb9up8KdpVLsSLVg20xgDx72R0haptK+DuKQ5yEZSH1P
VQeAS/zQI6HhwHOnNXWI3CvmjfHdt1au4CP0PhL5lxj6z3ZS3QABGZsze/Ovv2fc
IRcwW7DmFHFeQs+U3XcJpeiGohNxgnjbbxMxp4OuS9OsvM52fJU0BsYwxjpD9++b
SVt2pkaUQ8cinhwqhYDipNg6/Pr0PIzLb23lgxlQ/gIzsjErtmWRkIciO3E/RjK/
0CseUyIADJykarLjlsJUUwBxBqwdgyChFilIddUwmcgqD0ukvRNaJOrO5lgC+cjn
T2UpeLBLFMvYKmyuehf8WUG27OtlmzIDyZ56rb2ozJJwwJEJkMm3MBmRX2gBnsfT
LV5fwVO4Jrq6wOr6UDwXBw/EvrbJXnKyh0PCp+MhntjnzbICGE5MakTkjd6lgicL
B8Lp1rYM1WvpAkblemgSx/IsBoHQVUK9TCiw9XjT0CT3EWsZ8V02BtJo3rhE6v0n
DLQjsxZpi45THxk5H35qo5Kb/YbWnVX2vcwHR451HVNDXh95T9bhe7Zf2gkL9ZFT
s8baQKRTkKFQnF1j4T+3d4WmUtegUJWBOr/BEI2c7CP4JU9CGOsiZ/8rtvjm4bD1
tWXTgb+qD8SLLf057FKWmwuxu2HycjUar8gsKN7l5h5q3hNMYDBNnHbyCncKcZF4
2ASSIeRcX6lRJJoImSW8GOPBSy47tW8ruOuQTur5ok1OOp5kg9IXf/sSN8oPYzze
Amo/P3E9sl2lWmc7tDYR5XeQB2KQsfpDreT0WMA798CDd5NVR3KmNafkg+UAISEY
yMuPgX2q1xO68EINNlPfYeVbAo9/8SwALpEMK3xfF+iEbVsHHV4op2hETig2khg8
VNMYSw4OQhCkQmfqJzhhDuE2jRr3l9eckeeSFBKmhNdf4ZFN1osXhFp4If3f7HWX
04JN2r+oazBBC7hnB0CNrTMTkDnVHk4otQI9gYYemR4NrZROqeko/AfvPrFHE2j/
B/k44IcLbz5Zoyv1Ig/iKu/hZBPoXdffzIjDOwoJVWvKj+8xgBaZrighJYm4Ukr/
mcKmBry1S+U6q7t+F+/vCGaSUoW28ixhlXI/U31rfhUEAx6+ultk+QOp4r1WmpwK
4+/wNN36lrN+NjtZPh+Z5u64blZRdUMjhi4m8Hxcn0ct9UXoZcKX3mbGgnyDDKfc
yce4K1vrK1AYDoxRU5UHKDxbM+tqUVD5vT8uxe6Lz/Kbj/7o+EeIh4iR9q7iw8sg
uJFJVzjDiPxUOpbc4Pmu54vkmkJ0FpEONdNmiPTfByoJ9h1s7frWlPLttzhLCIVQ
xigT+Qux1sLdQ/Ycn/1lfeY48UoNSK2dnEGEwxss0mmaV5WAwLeUAJIYgPPr+7QU
lU9ZJA8iR6wNo6izutPEvI9/Ff4iQRAhbJUkTg7NFgTXC+Ghf4DxeSZD+SSB7FqV
mlWk0sCXhvOuCOiDQrC4/MOh9GzQE113P8W78lyqNF1/ifZ6tlMCMaU/8kJyej+U
FDBJYKIGcHRB5JO5IKCrCfiDo4NBVy8c63dmWepz7sjeFuiSyi5RQwqlAxnF2sAW
tHtmiKECVC2bAkpqL6PE9ON/B2CqLm69waFuu8+C87ojehVrkOwEEDt3AFSoVmlS
YmoGc3jykNI2+6lmMrngEuv4B+ehI7B457J311kK7hwTiMj9l4NVbtxRlYH936at
3dBmDvaIO0uNUcXX6xXsLfxavwljq7gBQ8q2rLPDvKw+Z7I5gh4sJRDHVPW7ZWH6
YdJaOZbMuwZPuNz3f4DnsdvllWCEdoWfO2eRUmHskw+niVw1CBUnVsiKCDbv/aVF
Nqlg1tXjz76mZ4rWcEpQqKVeI8SP6KK9mLl8cUkhss2ZVisOuEYaVmrqf8FS/NLq
KtY5CMsMQqNCrbeg1SY7QKYLlzFcohZSgWZSbsYToHZ4LHb3XW3b4eqeM4CMf4DJ
d4p/jk0ARNPUCh0RtHrwZk+1Kjhreb9/RhBqujFfySCX0r2XOcRv3d343GLZOWM7
DU7LFSMtXFKfhDpDFAIaDDyhNFnZbxnU+9n0ypD8XZJQm1XRD2I0yN+s9YYs3EU8
d+vs/dKaOvztOf9qiMjAXyFUxYH9wFz5UliH/JoTCbSqq+KVfLjSnR89zBQ2vgud
WJP5rjB6IP3nzItDrDeCLn9LTqT5b2nnSS5EvdFpi0etjRgq542fo2SJ0EANtoKP
lhokyG3I4+1NhUAVp2NT471VuDieDvmL3MEcJxxoNXTAVvqgYlFlGsu18a1OYB9X
4hTwtUyxbeM1FkgB1dPgTGhhYMkbtalCD0YKEcwMbOmsBNlnYC704QFJmY7uz2Gj
i1+Crkh8AjEi3ZXMxUPuzG0TU4gqXT6YC8dgKV1zwttgL7sf6jNg1HkxZSbDMeDM
bySgp9lK86s0cI0rDHWJX8SphS8oyY9ZeIZS5D9C9vVLDaEOFo9Blgmz6Mk8epfk
y220ghpAFmVe33jR6BmSYZlWM+XuRWfg1XbdjZzR2VQFOypZYwSv1kw6Xbqn4fn8
Tiokizm1Oyf/p+T1qJBArSrohEODNMwaGhB/90/dKI2P0vGsMv2cVYtq2/cU/H79
PS+5Yd9QpSGgKxtaZ2HMrBER+sSCYYrlGktnAAkZS9WLSGIXNaJkO4SeIhh2sOrG
jprb/Mll5aU3mXR9arhkBQmIALTKOcs64I8GYp+zKb54oXK12E127LcfOmSN7BUV
Xm9938ZbKtbAOkzegj+k9Cjm9HcbPYEPwbcPz1LjECjI8WQFYSAqZEj+hVTqk2kp
CBFoC7TET6mhhHGpMgekDRl7Y3EFMJQRtMm3QO56T4ciue356eGrvKRN90hbK81F
GoVqCMxygT6ael2hnr13uCmje+dgJhBonlA8hrBpt9woAK8HJkrtGijI7M658zm/
Kegia0NAcccWKxR7FjISgkwcKIRx/JZyPHAYl2aeAGJxiviNqrM7dSYfOFmurBlr
tUmYtQJGDncYVgBXq4f0p0Df9sUgiBVkpITcrVBtlIvYTtf8NeJF1dN/V1dqMRKL
BCYeCOIZHeDgnmlFxWuY27dVG3D+3Mh4D54l77V5Xd+bgmAMeuMYqGSOdTUf10lQ
5tniP81Nz0a4jgmKblhzN6eTR/yJWk2qpv8kcpJ5OhOaC6xmy8xG60oCCph1jilW
eNE3kOp3nwHIrOgVarwKRweu4ObTKMhcTsi1nVuwLin6yUzN0CZfXuvnZSC/KeLV
3uNUCYOk15mn8wxd89/maxSIML+HEN1ZXBBgStPSjxfSR+vyU0kWUMnUCpqwRbw3
yOGdOq6nSLT0ZRXTv33w1fWnZu1ZFTAvnkKyBx/C6/FEnBu7iErkAQCgGIUddJLj
QfLb1DuXhUhzLURuO+0Tu6A0mjudCL4/TJXNl4HO2c1lhDqpvksaU4FCNc1Rtco/
DfNyPZjvxO7V4JlFLlDuKRiF5+DxkViQMREvaDW8C659mTPtNCgQhvQGOG8gqQT/
lLaJErc9ujEgyEq+U+abjrwMmNnj8xj0PaoOvtIL/sj+eGd8xuB/j8V6L4HkXjXM
lBcT+UssayWuI7QiNWWzHYY6M2hQRYnCNiRCz2UBepAHcSJeVmVZUykS2WKeqemQ
6ILcWeMFc5nxehGdPqh1yM8ZbWo15WcIyyp4NIvfh8Li6I3tHoVsiSn0iiF8naLq
esOeymo4eyUxoXPKaQF19/6EoagnIQHG6DEyCYvO19fNEWSojXj5CEhwoLqN1r+2
MdJ4b6dimfUd87jZUDWyJZAtR/h8tKZ5J/PXFaftK3oOmR3Db72pS3MmyHuTnre+
UxlZgRCgulH3PfQP+vNfOvgF04soXDHzGa3ldFHH/BTFSYXnCnte+BmyHhGdox07
q96kkrfpEsJA7OMHKCPZ3Ui7qZFmUUxnWVaCO+5KDXwFAemPoy7g8aeMQAfowyq/
kOJ8RImm8/RhW7uvzOE9MQWgAxx6esfEAn51OHXJhjKFb2aCFpZVfdOACXjXKaIp
Fa7TxCJXHtq90TCs5RKUjWGpNdlARu+DErXIR9syondzl4ULUR7Biy+CM1oHrvxc
JV0dw60Mkzzm5UHdWDERrHUONddDBdP5oo8KPenvOA9YHqv/SB0/6y8yivQSQQY2
d6v95MpOEIwiXpPKoMx7XYdVZBw0bEVOosW/k8HRAWRDXE0ByZa181q9VzykZ1Ih
3Bqq7/G9Yxaidw97b2QZN3AkMUsuEuIidAmMJORGZbiMeSlV+S/yXzTBbfVibfPU
a6WrSDCWIG8bEqQEgm3Up4mQ648HdojqcS2EY5L7ls7sq8gNqyq04Lyn1a2FOFmS
iM3RrcILdBKuCgiAqYqyk44GiGLvcY8R1HXVei3beiWZTf99mULX69SYOeoFgS8X
+RbZt0EFZRn88HmuNFYpBlA1SfGxX9R2SNqcYZveDYjSfQ+uYV66mWPv9Bc7OYBs
zWhM7oGnsMtkJwvYHSFbrue9Dxr7+JY/zPeshTIseLsXRv+NqTkxtMU3+3hJrzTX
przfxu9ad+GGJ1b6G6d0ozgF3s39p43dyCJfs5rI0jk0w8yO+wBsucZtHjmX7uNK
KRG1GSoM8AFPnNQZgrvY8BCQWxtc8q/wO2KJhlwS+m5U220k744HZmXLbMkjN4y7
a82u63kreymA6Zep3t72kwx1LhdQcHXx45KNOOef8u+9AoyMYwwJvmgOsEHCmdO6
UiZv15s2QJbdCFeBvTVPm2BfOU2twJg1+lHbeeyYQoUPrihjvkvXP3yIvFWkCRhK
ONLWDN+BV06ffwHdV4g9vLCyKUdjvEz9mCjnZUZ69m1AgSuqGsP6GHhiT0K3Wyyc
1rnWwhY15uotECj+NwGlqRd5Bbmdl6/wDpcBnfubMZQ3sW/gamPNNJXLlFgjsDbr
axNBAXs3/3BmPvaKNZwnmneMW7vzLaKz4bphOTL6ncFmzgppR9IUcZb9MbcjzTeq
MV3anvLO/JSFKyviswLHb8NR50hrrutC6aBu9LK93oEYYe/sP2gDCBa7s/pUUZ3k
2eYJ1VMyVpEHNjgRsgAudxGgwfXq+aCpdpHDbPXpfcclpiFSBd55jIgPa691FGl+
rfsGh4rtXAS/8feUOQE0mG04ImGl/j0riDXrrnHT8/i8fsY74TbiV4u5sFHERFSB
xn8VVkl4EKiwLqu2+rrubsUxpm3OSGRYQrYU1fwYcME6t3VE5VGYsfZ0t/brfetn
Et7nGyRoBVcC8hi6Msp0sM6AGfaXOjO+pljHEwCNs7wuivMqOKdv5xUods11rWlB
cw6CYe/Ui2uyClxPujE8JYNYdoLNYQnc62Q/rF132p+N2r07gmIx0bRM8o0ai81e
oR39TjbsLWs04jlA2x2J3dbHgON2CZPAGhYl/wN9BCOZaHNW9iUp0YxkYgEWaRBd
+NyiuIKAILY4Wa6amVLR/DzCvGVksKer0SLZN2/wfxRHdlHJFe3hdJG0GgUIsS0J
J6tOruZtNYhY342GS6ajDduM0BY2zx6+W44dAw/cna10Rv96YjIX84vKmBKJzGS1
bB98iyh0e0+DA7RcCS+X88WYrOHSqivEPQhsT9Kzgx38U5z+bj87Q5rjqa8CuEfF
PRl8cI5Vs557XBmC7Q7I5h8zIB/c2T0/AggHFedoq40U+LuWmOokPwpROTGBERIM
7pGyxjxeSXrh8y3IFendpsOzB34SAve0+LfFbvcLUSpHxNP9tEFcSzc3qXxkC2Fl
lxTTAUTXGLJFHzJM7JEjM3a8pEcuhw4hSFkzjs47EePknGfanlM3Bsk1WGtOwLqZ
zq98v6PynjKGFmlCKI5u2VCxljUbX/AQbM7yRRIie5qzcRTXnMOztaSEkVE3VzSI
00+nOAqaGcW9XBJ1Guh1tkqEoG63xc+iRU52JVBIz5X5uNh2kx8Y6eo8PjS2QSv+
0J3VG2pYsrChtBdVdCbdWwxn6E/6Yru0bM2BTNK6SYr+BGT7uq2e1S8oNv3OCE/c
4GJeiM8x7/4dX0ggbD4h2MFDaTJCvHLpVMa0TtTIxkeIn/hsW0NyTvhbAtwVdIAm
JCngAF55wBe6IF8tQtPhjq5okmbz80e8qQbNGWWnOpQyvL378KTajYhTSWHg7zRT
wbLXdvk/CHtLpx0wqhRFlV4tgQyy/Y9zacKXc+njWQVFr2o1X4CXYS4HQZ/UqhLY
4VzTpRcLGPfBTerLz6QEvzO5ReHl2XB6xfPh3QeO+I/eg0IXboed67YJvnaJ5UO6
8biNgHKJVKMA6GC2zjtCuLKl7jU6UMV2fsBKamooTF1aHS1sGPt02mxAK9SONkPP
IBKC6AjzY8e4XQ9RLifysMBBqUbnoEXr0to1Gjbqi/J7302xckCLnOx6AoD4GHTn
XLP3xa5EuJWAnl6IMb914NTwpiL4LelWLTsFgMA+LPIt+MhJIt4DrDZ4tNm4xxA3
NvzFVTxT+jSZaeDY4UWdi1HuIVlSqqmvl3ccmi1rjlxAuxQafYr5adlQ21X7xvf1
NDALahzRj7ZKYrl5p/l1iHmpQWPl5RoEwkMsWxyiu5VCkNW5LGCzpIP57WUcRV71
GOBVILOFegY4eLzZXu3Goh0mjfcGLUMKu8Tr540k/wAmxGcTBgvjlGtyKVdvQAFB
NU88Llx7iOOlh2bfkKenTGBxr06XA5MeGLMhSzmG321xeRSdKoz40WH61GaeITN/
ZgaexhVCEKwuxKqQk7SUj4x/5AxpYFAqwpoje6U16e8OfMxFoOyNU6nsTMVcCfPd
mZCPpYUBl4lPoMEc3qaTAzW/l8BcZ88GoAyr4wWZN1N6BbjgIWWoym2MvRvi9ccp
2LyTQFCNBsVWuIEF7cF5YXIINtoinMPEZ8fgKTZtFCIpQYJpwJSAdXrj7xtw/cav
oxq2YnLem2ZtyayndC08Zs2mBCCzIErJQ8i6tq5FMAcFDAmoB5y8JRKOqa3wVxfq
hc3e4Mi8NJdUjQKw2iU8+WNZHZtkfTlanwUGdTFi2alTWXjvSITHtmKOXS2FjjVT
mCh7x6WqEinYQORNsNfM5DLtQaL3QBiZtsMZcLzAzDNs69SuHv7OeJ77+hYfR7R2
UALKLT7HTlNOYJLzfNo0u3uGEQ0wiS+419AA4Wq73UFjLQygajyDpFYEtS/+ZGn6
qBpPFa+Ao7Vnsx+v0vdFUmUYUIGgSLNpdKtA44DBols7CahZ/uB9l8nvvg27+6Jg
HRfa+uz9rFQw23NSz/JEHyJ60fCBxDL3Zx5k/bGcOLGGN+pFunOjznlZiD1ZD5w9
SYnOPF2NY6x0i32t+slnZCiRjoMKxjUwHlftYbC38G1Ybrr67enPQ32M8D5Oc6++
WNoDIxGXnCemexVNh1VSwjk3sEXiVhDigEURXt5S6mMORrIJlg/NHHxP+B3LH1Uw
hqVO/H6Lj2QlC/Nin3k6hw1WoUQbmqb5PQpgV90toJz2NwcpADWY01DfaJJntw+1
dEYvRdIcmmOR72ug6ImuNOQqZiBAbHBIDdr1M1bkm5xWd6gyFJ4nPIVkHOtbKrbH
Zs0P8WObfvGfsBByxp7kqiYRVUT6D6+RBIt8E0Y7R1OmI66+WhPM/gSeOBm69b7e
OvMoOBRIa8Lj6oQtZ8nUqstVnI1IaqvyDqoAfVzMUmPYoff3QrXWdfH6ZbVjOqTZ
xJfL5hLbSvCgxJOgm1uyMSePmf5f87Hcidzg/doWXne0DK/dADSfWnLOHyIfwxR3
bKVQ86CPKdXQ/Gm5U7AeHIbLhS8eCspxYboy0aRJPCnlpWpoV699mhekoL+yACZ9
zExo/rdk4dDME1aTFxxfFYLKULtXKlGlqztrENfKE16nKwIYbMTKZrUAo/blrrcq
QknBEl4ymw3UXuXvq5P5HrAiR+BhgAmJmYp7vVMdKueBobfWSXDSg1+u1cQl1jMZ
qFM/WCnclSYTW0eXduOEjD3GVAESn0qWuwsUD9e/dPzbdtUp5cptH4ImJwUfFe6W
1GTkMZXLznLjb9C8ZHAqcJ5qk3kpqtHn+wNEPAK8IjMiGa6mnZEU8bxcSsPxhPfN
IEfesI8X6zEWYwSDEAgHPOqPCzkw3NZUg05mO5wfjRflwx/t6m0UciFG+yF3c/Kg
OXiYbt0KoiBERT8ACW7x39Pn2QaIClg1gwVYzjKBE72evj0BBqxeS+z9Aw3CMDNf
M2ABGLPauHJ2KXJEdviVBWLwUiBl3LNyDgN6wva+kb9OPd4RcX+a5cCOP/Mgt6B5
194OnMfTid8/on8/l7OkEdj4mgjVj4ryeVx+ge1JywGN9JGqdzlhFu5MugBGYDyx
wiFOizp7EaCwMh733/KY1z6qTe9yVr7YOkGjkFkHi7naciu0PK/pueCKIZ6yKprc
83Lni2sc17gJy2eJLh8EUkYgER1ePYL2S7QQxGRyrCfx9SZhjPWqrgSPc/+IOJ3x
72bPfK9x8v5zdNYAyyZLI0UihraI8ZyC5v0kh2p7xufNcsaG1qt84uA9Dr+3sRH9
qDRkIVHE49fXetbYMYDfsY3/zk41J77PpgxYU1gJngeZlQGeKk3UPJbu2PgK8Od3
FxRX1iN6Z4eozSa4s2ERc2eKLx6JCZhadWSwASKnNpaktv6bmxUE5w8sHFMxxM0o
d6w9mCLI8V3CAq7M+2eIE+Gigdh1AWnvryHyepL6ayv0V0jtO8jSlSkqsZkIwB/+
wupQC7BBzGnFu1JKWkXt2kkm4MpaUDqmhzYZNd428M0z0KgM/oGeckwU2LnbmD75
fhfchsXMq+6p3DIH6QG+ukYq6LjGvcnzyMzByj81/araoXgKHCAL5KO83DbQuNGO
ViF8NrCfE39IEEFrNaNuEHSq4p+KkW+rT2Z/0dvHk8k/HWWoBxWQgsOaX82Y62pe
wW5aLYpA+cpBE3wsMmG7I33c7l49t0mNUE3nMXf0i9X8DJZgN241ru7Y8icB67fJ
6XlF6sVBJVKZIB8K/tLs8soK//LKvzlqNwZlULXNGTDGuKko/xw2PrW5r4YrFN6h
36L4F8zfZOCccgzVRfJi5GN4t96GQu2lvT17c1oBBL2ZsKKw3IwscCgcPGDgDekO
uTQ/Hv39doZhwofoBZtb/6XODJX0XcSsbFz/Kpi8Joza7PaU+2vtmHJc7ETn4ImP
rWEcd6x1zA4rG9bhQIH9aUNpE7mu71dFmNh596er6jtrJRnr5cRzPa7bUex75yvS
8oLqdaYwGrmfHgAg2iB9gnTCr2RMfKMZAxR20MX+O/rSEu+nP1P3wzjLhV3SVUHM
F1e2WLiwLxKlTyyfsg4Xahcuo9iCZRkECVi6n7wvSyh6ApZOxL8B8MpuXA1NHgfU
Ii1A+F3Y+SVX6B62MuH9lq5IjK0vv5qPrBdCSg04g5mDMEgVLVJ1eqysmH3uOXQo
roFfVtWRdlun5v3ku/PLiPhlqSI11E4umD+T9NAjbLUlW98ckiIpuPS7kRnxYeND
VoHrF72Za17wLddgUdEHoj+84WHvitf4D1C2SMMCbmMSHuQw97CEG4pRmPPRcpXK
+XBK4p1LMwU21a8PL6u8YzyVCHwXptOFelt7ohgn0X73QxDm52Fcf5YURpMLZ5Kf
Qa9cjCxbNSJPCVEHfSz8Inq0GC08ODD7EbI7f2oRTWQBWrqvlxi6kqxQM841DWlL
aPhawOYBm9QvaPYqYkOWn51pHu3qOqiJmuj9L6VWPgozGWwV4fR0J5xr2QFMpmnM
C894loM7wYJh9cB14SGpWaT2S39qW1lNrSFsdMxeGSOkQHIwf1Er/cF78MlAnMz/
2jmQQPqG+lwIlGKTNJYZIgOuF41iboTMO6GlXw4TLuJ7thRGHbCfCaTWwg3TJ/iH
c/+p717ip7JZkWS7brSqPGHvvC9wK3nCV+IGAGOZsdkawuCDImf/lsZMQm94BhHW
xiAaAF3bmVq/wAbActRDrPv/jBXo2UaKBBaB+UacfkZQt9osQvbR893YXML47zhA
Kx5lUR59NEMoylvW5/fUdrA/MfHXD5acBlWnOTB0JThgWved+BM/kKonLG5KSpef
RA+IlzDLKCNqeckvQ0En7FKQVy65sdn5eUNAYJhvcJVxw1MFStEnHJiY6k2qzaKM
1CRVuAwNI79xi6MHlGTqYEihby5yIND7o1ORUEiyvZXkHjNNAi1U9TG7IK85ys7x
ZoBErJmBxYH4+CYbdGlKQxnvxOTrfOF5qB7WolTgsqlZTu4GyE3vaCMjKtDEdGIf
3b8n2UtJvd4OqeqWuex2ange7y7zZgwmPqBZ4Na4AC+qIxW4RGsK93I3tFJ0yx/O
uMlewvcCm0Y1fdTmFnvvpTlsVW3nlztuW2dwFIg/xkvA0yQKzhHuxJWDHXJmfHYw
wa03zmRVXQcVsgm4DhIukEYvONlbto9Cg0vx7QxcfkBKDi/sg+Bh9HSLULpV2Tuf
jFVfMjEa+KtyfvOOh852CiCk6knDNkpov8thzWzDs7U5pP9iBNyNAcp1+rDtqzfY
pgX2IZXJnuuDkSPbhRxnQg92ty+05ny1PvTYxsx0/0r0i9zXbPP7zeVnBE/sw6tQ
Z+KCrGX9iSr6xu7c1mbAExOmrM9aQ1oU7rSfkoBUOLJuOVWwBTkXV2u2STcJdU19
bbG4BPtFVgJJEhRAY2mWCKahdbCNhESVG6zyxXD8WTYbMa7zrQROiEQikumdSAIO
ZyUXL3JLro6pjx7beBArd3Ym9prKDirT0m6d3+OX2aIA7WtBcM0qBDka4DuzfG69
RSVei59JguA0FsVfF+iA3wjDfoFW2Qz020T3vaaxqySme2YgaH/scoEAir7yUyuU
KmoFP7KNm0+Ne546uwvfobnyfobNFITT4/9tRJLhipRSeFW0TvKJQUcnZ5PU8q2F
wcEWQT3FgoFI+34jdR0ODremIXj3N6eXyrumKeHxHAyFiASqmmPrBq/QU3wQoDYx
wIA0dQrwmuWHfs2wwrCp9nN5VE5W1f3ApedrWhvk6V+hk39DhTixGjxnLUjGDiBT
k6KaTfW5SstfLVw8Y3GY8fgxFBhMK6xmyU7c8MaXiPNoMU/5OnZz3eiXI+VYlv6g
v+yu9+4TxzhAnbsDDplbj9FhEuishizijaKKQDlnCeXoqAvCQiFArSlk9Go6eRjq
DMxocxitN9pmtzyQnrNAQ8qKA6DV7NnSLwbMsffeaKn4G6LQJttuR9i1yPQ8haeu
6IPMO+TtOWcQxBcJmGCL0L29doEDolfTzczLBolS+ClwnjaiSuLfE9PNQmgucNUP
tuNq11VVgygOPlZUrYaK+/mMpCrhr5oAoeGMZ7yGMXWWgxs0sX6pqc3YODNQGL9P
12SvVOn7qCG/wcjxcY9qExb6nTBV7kiksegNlHAlNM7Y98C07+5W//7C4vKJHCJr
PKlrsBgGohVFTb8W/O7sLR591zgIFL31ctXk3VgE7a1r2taok9loZaG8PEAmoXyP
Mm8+FsLe7ygjlOqns/V9LInLpY2ZdO/t3/gSDuJ6gEBrOWn5J/uhTX2r9WqwOiAj
0YoTCJKurGOMPXLULmL0cOzzZJiomS1hJ4Pv661GdnjgXP3+EMGVnVf17kcWC/fK
fMn/GlM7IEmwjOJBygrQS2gpnWCJzoQvmYNdXZiCsR5z/4OcIEvf+uv//NMHkLLF
launAGUwXSFjk5Rzgz1RrBk7Wi2c1vUAzmHznkD0oFhFMcdjBGxjEg+WIKakupi5
GFrrvBKGVs5tlKXc6T+67Z1F6fYYGh1A38gu+37pnEUpSVchMj1xSAwliRoVPgKo
ck1SlKq6/J5mtRYMTM4pB94LRqkjnP2pDJAxWCep6bi2tKiWMaZh8rvzMprJyOqa
AC1Glb6hX9XzHU5Sg7eeAtcGKr0e5iRj7R6x6yknvrDIcS/YFpQ5yGzS31e2Unep
v7YKGs8d/GjZCbY7UyMPo9bHMZQh8Lnl1w8MipGCpwcahdtNH/XVm4Mi4RrtMZ59
3OKVI8IqBCq2AdVMcw+hkhy0te8iDTbDel/d1h5x8+vRYW23xboPejBASzufQVR+
eXytblP02VjKjIYu+2zNbUc9tRpeDxMTynV3VmjqhdvPvWqIay9uW9irM2R1UwOj
77VjwyRxrAUIob/8tQuv5MObOreTuZQiiBPSJCLy9a/RVVW/O6nBqV7tRL8GBxtC
wl0sFQBw8/78FD9FxxrqwdAeY+WIxOAOVhyIvCf+KZi9k5PSkajyLqU4Y8FRfDEf
xiweBqpVkQ6R36a/ng5WzAdx4ehiOR+3azwwTB7n97S0u3n5R84ttrcpJ21g9Tpp
ZaTchUomXGO+7Pw+iZmt5nuC0q9MBf49Wg2Mw7qAQqGd5DsA8ldyUvC2tmUAGAuR
OdPej50l0LeWIui+Vun5llYjHOsLeF3SoNllxCAmU50hZ6btW8+qph2L92U6wlxi
AR9EKcjXsfHda3pBFLHbWgzRmIz1dRFqWWyKaPeeR1KF8ghICgG8iXbRlsZayabh
xEhKNWWmk0EkJH3l3aGZuXvJZ/ROZ9FZJkwVeMdQ4Yth8DcsvFU9Gh1Kj6LQ0uhF
z2qkGzbZlgkwsIWZy4z29E66EGf234vUBjiAwOglg25ksah2pMeKrXSoLGTLXady
40WokrddvUGN/XgklwPtkB/u8UdmHO0aDvUg4yHNACc5Vn98bWFw29r/XyFVQ0DL
ZPauRjKSLZ9xahqSGwtZYSu1FByRTj1tdWiOh8Wv5SJXCB6b8XJg2JVcSgvCFoI0
6688aDZXaI6UyGxrJOK7ikiFXsFF3FBFhdh/4Tx9MHJfMdSm6X6QWSX52b0HyPYY
He8sxCDFCLjYEoAkSskL7E38TcXffivef87K1scQI7rWkyMCIXUGUx0ZZtp9S/9l
jIuVgjXzWjjBm8P46pPeQ2zbtdRFG70RKcti7TAQwLHJfyVGmOgM5gjwWybl18a3
sLIZCzk9EQc7m/DJiUWtENzY4rjHP9yq2JQabzNdInvV8Z1+sxezNrIRfOlETqMX
lbvKK/djeVOOuY4YLGnaMIMUKtoetywxHAZw8D0wWErC87NOc+qOJDXcEwQnLnOR
jwX36k9ST1ei9CtVdLv/6LDsn61qZNKhkYRgea0j6Et2NKj/jseqISGg/ZiwzVCb
D3hylOJSAQxNB4FP6uuWizln/9kVA3JDO5R261Ww2tA9IJ1hxVt3wlI9VLRuP2rd
kvayFQSs3qQzNHNC8U3R0mWzvLNaKUqRryhRbjyThJJHc1Nu4E9omqBlLTZEgL1M
Uj8+Kfly7gLFTY9C9/byMLxc9yoqWBbuUfnYfZKzeeR33YRWu8ttf7DzLxhOit3I
FX65Zqez52V5w6RduauGlYgvvoK6jdztW+Qq2iWDnuQipEJT3nYaLWpQwkw7AF0Q
ywJUWSZ8No06D2Li7LI/P1fNmc8qPIFoAEYLCxMfRP6I6mmB/YV3/zruU3hbXUGg
ZesUvRFLkoM0niAObY37ihbEgkvFPzwN1eVN5bV/j3BHyvAZTyuV8Z/npuuKksyk
9BFdDGWxYKW/2jWMfPs+epIp5e9g77WJ1UcQZItoW9fGyBhT6ZUdB1y6+y/jlFLH
L/VkApcgZJzcyO0ISx6WjbTM8kRdmBLXazbTd/G4CPPydyUY1WDUmo0u4KP37x6E
6ohpEEzH3uwmd/TX3iflwkGDs30C5VSt0hBfcxvLMvD1MDLYueRhFtoYXZ7sCzHR
aqjolGyBTshf0r+/UNaPeFjeft2EVIQ3HxQH3TYs7pPTi0D688PY+6WQDOgC837R
AzsRaGzt0wXarZysKAdPYxXIwIMwJCo88rk/hEXny4691HSyUeUy7HmeHKvhvtNh
RYiltQmWsX1qYs6aCWIQAP3axWHU9XToRFJUZB7ffQGpGhb6UAuVHlyN4vhriBVO
UpYghy+JafsTtwtSs9OUJx72JWJoLH+sYoQJUxPVdweXqxsGGBj0YKOGb+v1dv4G
Z3AlWwSOB3fTI7Qkty2PtEC7fzBsvYN88xLEANqmJxyOaq2rg7e6Y/HxJDz8VYcu
8Xgl6E0zvF+H3m86b4xyg1lmAG6ZM8FPbCk+G4AXOvtqr3UbK3EIPR9hymIgxS8W
Vl6OS3+BVNEWRuO6fyOeGCil+HKQovLWoUjwPD29/iF/SIk8WEI4RokFCGXqilsX
WXJwyzXIXLJ/0GHqnRqMBYEw75p9HHF0ozBSh3DQBSfOj0twlETTLVUfen3NROYc
N3qe8k6a+Tpgq6WknnO/jg3inMgGEtdQlmWfJBQKKapwPuD0qsijiRCjXR5whOe+
3cvn4XPDihY8APxP9ig6jB6bztHCXIJyH4vlTqosK2BervgMk+FzWh+Pd0GBn3il
UqVV53ImRYrDT/IRE/+AfFFNoezxwfIPdKrEY1xcjD+uf/AR6S2z0XDb8Ua/p5UC
99hA+UvGmISOADmi7uQTWKM6zlX5I5C6YvcQLLAu26nYUlwLu4+B8112M9+skabf
66MDcIXvf43vrkWGHm1yFOb6J0IoIKejJarWzojNRKhvmV1ohSIa9ocdtaF/XQhg
GGqYUdk3PeyyaKtb5BNmlueIT9T7aa/Pdg14304UKoOAi7Ib4X3nOWQWSquJJV9X
tY/tl3MlSzUt++nVOs65jKmm42Xfg6PGPEjcEVNiOPoDrvnbGNL60+5qs1/A3Jbv
7a2lpgMQ0UJSYWMVt4LbjTn40Pqy/O/F8A5KV4oJ+5H2E4+ocnnSpiZuuunnBI8h
XDw1egUUATO02YW7uYlcq0HzueYHVCk0cCtxynE+tj4iheAVZdVExcyNDHPdHqAK
WvXCaEyyy5n4swYoivGqL6qxV1A2D9+z7e1AburXFyw9O+w5hkz8SPfkTb/CQ0YI
MWDml4kyLcRfxmdljrkvPLRXj9QAErcGluMWEGlwhxvSqjELa//qQWezSbrmG9FM
kb6bTm9Z23DGsQHbqUuI5PME8pQtIRQpZdRUGpRGcl6uGJa35LyKBKj6qQo1uyDd
YbABvp9Kat5acZp3GGnuuIStjFqEbDuehwQwc8PlhUG1wV5CLhnDMAWanfcFrqBb
08Qd9dcCGItho2UI7jhq5BK3Ans4CerKZ0QinMDMz7a8Hey0MFrj6Pjmd97ZzbAq
3Xk/fhd3ac29rME8Fe5gesFl/XcU/YGiumS4dftlMxWtKIshUmvKOqYy70cQMORn
57MUKtB1Y6OzZsinI/X1WUvohSTjAiJOuy21QZsuStNb84w/79DlyuFco4yZtr4K
QeVHItZCKmCt31R2BDipaEnibzmZH70pMBlm35aMCog9jIRndkLE/nCmM9/Tw6nz
vbO0kU7b5+eKLrmMUPSDnbH8mg7tzrSfByLzTDLNKYd3gMnQhZv7+C7Uqbs32Akb
14aKNmkp42BUxLF8x/YjDKxqYQy3UJ0zNAHugICDIBytzYO5VEPJYEwQZ8Jte9TC
Wok8pAncYiJsk59mGA8xvsvWAS+hivFJYN3N7GFFXuM5JAiH8ireCsboXcWwAxG4
6l4CF1Z6/i7PUwj7nPwkVkipObBDPf2wsQBbIn2zm1yPfdf5K+oAM5BeR4FoJJPS
lqUe542wC3ZgCk4aPpW3qUzI5pWQZ+7fT1zyWBsNBLsIVascjUkVCY5Fd//1TXNE
FUhCxUvuIsJC89MxVWjeF16VAhV3J6Eown9c++ruWp68Jv+RPdrhKO3WNFVQ45KD
u53YpAMAjBcVgLStEQtP/CJNYKGnSLd2QWKuH3uTSQZnthAYJ3EiZlq8Wx+tsGNO
qU+ax5ie+e0frsCRQS2OhIBB7FzUE0fz4vIVtZs8IKOW1MAZcaLeVu+5XoywbDqx
Gp+tQ49J41XPEpcYI3Yzqz02Z+egVGdUJizEJ0KC3YxXM2flmoPf/du7QGG11fiZ
LgVtin8KEYF5fGUW4WngTFaLgmV9U+kguI7eUpWZ0QByAfmwtUs9M+HJiVuaM/Tv
12AoLzSjumSCJV76UF7Vfm1aoUIZTgQw5emmOqWSbHEHC3nYs3ZPHrKAsnkmj++D
jqnnUCeZ7mh+fojlrm4MAKr6g0DRglUbxCYtXD8pN9+WCagML0FlwjXGB05c4w6s
Q86ECdhIQ9Ke8GSrJYM+mtd/65nOImoARn6q8rzKm6BprV1YH1jaA5t5UtU+Jyzw
d/9praeOiLsw2GiI8iH1xRRmybQF8/8WGvLtJvRsZW7XXAh9tT/qMVOdEVckX5VU
Lbi5IZfXDiEupJ5puofaMDu0SWsQ0ZruwQXpp8tcQv+6HwKBEr30sAgoIfeaHxkO
CPi7HMtJkoYdqNY1tXhshEVwe12whVV/p3JtP8MWrraLxwHdwQdlKMMnUpxMhWi2
WBi4w377+qhcFzXCopOzFHpRNas+K+PGwCfrrQKj0lGjToWNlXjy47bOx8qwhzG/
He2dmnVrF/mvmdQaCLdezwvA0QDbfw8Gx39gLp44cGg7k/R1Svq8w5auMN2HcKac
YMmLnzp5CZ6bgfRJqnL82/Nmr6S76TncuFFzU8wZGNx6OdQwnoCxCYeeZNOoq2Pr
u7wRNXl3nPJNDQH2CphTY2Y1OptOozB64Yfgs89QbOeNg7zwjLMAwz7JpywHtbSA
D2drVPoJFd6WM7+egMKx1kMN0PRYEKA7SUMb4Qx7DTyzPhzugE8m+bBveKhGEBQA
fFcRkHRZhyUGovmbjzJE2KBHJGaJRcmZf6/wMW4+tQf4T/iBvmZYbmfQYyZ2hX9W
yKLA8CCJDi9Pc4DhhvsEYJWEKoLGuc1EtbfaiwpIdO8yt4NwYun8rXhkQdQRWT0K
fhv2kQDEZ691SQrF39GPZ9ynGqCpMGxoLe1SnLbFgft/kc1HL0t7NtS1BZ496unT
Gs7KHC5oUrlcibiYDrpaYRyiio0Auxg5XlUy3M+0eHhocf/VOPq/3xCnpFdvk6JS
8KZ0klxz2G910CkhuUpebXUYGa6QPxL7Rkq0pdIb1bb6/iz4Qq8aHw3jMYTmG7Xe
tdWVB4hEuysxwHU/cf1DVWlesdq9OAMRSiyoTRfUEVxreD2B0fVYXTAhi1bxZBme
JIyU9QYj8oI25l681sH/wVXsZ0rloXQXDCUJyvlfSSkOzt85jOZQFF4ZGeHo7pvl
DpAEJuNbQ3zC9AmashWpazb5sa+rsAfYFj4j3BOJr7h4DYBzGaU/flaJpZJU474n
nflBLL062OwpmrXHYGTRB9rLG6/5NOCe9086YRNGBZThDeCC2j3jcek4ddsXGlmb
Gz2GnZO29mdXWD+4xHBIxReka+VYImEmvFlosMAECrmnUhdkyTcIC43z/Wv0Twyb
skmZy8m6zVailj9GgsUnBhvSBmD7mH1DWbrBmpB4C5gsyfC1UTwnMY6dfuY68yYi
F1497kY2X22SlyP5kSoRvxMaKv28RXk1px0Wbjd+BKqisecnucAi6bTi2OklkXWn
JbkK2AAq6DtLde7sTivaDzN+E5EuqpZiwhUqgEs3RtPfGMyYV10qbtU1odXMa5Hw
EZpbgsRKfD8TaUk6rqQwSvt9X2j5kHtS4kRs/Qk+Ci57g8hwYitGoYg/GLWoIg6V
8PMWFgMx+b28sMP1pcYeupZZ7A9gKC+uI2BiI0aq0XgF7wOHUJdEYVbb3FdkZ6b0
c/DbqK1AkyTz2o8sVB/cytZG/NsWa1UsTgH6ez+5Eyf8+GHAgaR4z+o2nqBnoAwS
fgun9EScC48ohgpV68m0gRiIT7735RTNYXnsH2SetclL4FKtfIGJVsZ/kp9g96s4
WrHiH2/012Lym5qXa5FkyeCjaDOCOzJdp6D16i14n1i31xM9fShCHQrtK0BO14l4
A0RiF0kywe0J1Zke8Wz5rsvjZQT3H8A75Fpww/ljuiVi65jbnXTT6QvaPR15Z8gu
GVtfRhWrj2/gQIlwxx94997YvseP2RBX7hlokRNKi3N4J/YoBw8qJoPeVJmJ8HA8
cTuaNzw4TJ2244CFdwF9Qm5/RbCudiup1BVY80rKhUB5Y+KdwlDwI5z0ZIW5PseN
u/B93iUu58WQkpGf/p1+F1uHv5lxK4F1jbGWoEeIe14lse/XJMEhy+/B6GADz42Y
mAvROnHZyZhPCR4prDIftBmptylWSVvcQb3xe+0tFgRgDSMhlFAfv5e/WcPH+z3o
TxwAHdg3DkvFdSTHmxUBdMgZi9f8a4Oaigsxm5L0HloUJ7pNIhNirwaPu8CXEmNp
RZuI7+rDbYqTzKqOccojM33dsfL/FvXIxZrzfjc0shZLW45sQJSFYz1GSCBHBddS
r17wDx6aVDWNkd2MhzFUGOq9tg/OcsndLS2/wkgc/IkuoDKbiBqlt2lUd/Tp3dlp
Z/tL4QwmpUDHCDBzx8lzBkcYwlPgKVertPTsl1iib7REiKn9FCDzTVwmMW4eDrtj
+xfZ1egl0uWnqfnxpof5lzqZNHOGebfUQ14QtJynRfPl8P0G3APVMBtwLnJ1DQ8n
SvFwai5nfo01YTQRF7HK0KtiUZYFSbCCO3u4UQM1oWWsqSKoBAI9qCUTXighVahk
6ZM0w6iZ4XEueYN+a2LzcOBXHiUKIzACYaZDkX6JbW2glLZKNXbN3cWZJAP7TabM
CbcsNgp0Q26YXBnWnKyFNKhutG1dx8djva1kfkneGHkld6zesqxfeLUk2a+RRPNG
ZSCavRYAsK7aEzW4HTaUjP5UZqL6RlNOkd7FZX/lpdCeglSjctXY/YlIs66wTkZi
/wEp4xk5gpkZ0KFGmWQ3SO2UHXHKaMRhz7e2TBZKwYnenXrq6xY9zI6q1fMscPcK
4TcN9aVhcW5KBWgFc8LwmNq2vAHqlxKDNIt4O1PhaYt3yb2Vdsya5pJNmQ8rfKFr
CU6v63YMvywabxxo9GQM6XjX1jLqo6qFW0kkHy9C5TOgSRHAxKJCdfVU5ILNTIyg
ju10g4bT0TS7xk/0isBusxsSR+RHQiAjk14DM25YH8Nf+34Tt1ti1y6EgV/FAJTw
`protect END_PROTECTED
