`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOB9bTk+NWx3RStXwcywIie1+Bz+HL1jFPE+lmolgxHT9QIkiAMkeEnpUok3mUwp
SBUKC0nYqSiB2j84YlbtmG3SBaPJVOrYVqip18hcGFprzWKhgFO+x+LA8JlZbBWZ
yicN9BxLN138OY8F3CqWS1nJLRnIwFErOsJGVr2OV6AMyq/tqRtpA0R3cP2C8iNK
rQ2KxRnbm7z90gh1hXNNK2LJTHoadlIKRcNohFeLS77BUbOhROoF4o+Di00lIa78
/StxtAZKZSveyCgT6AOfvI+6KxeC8VLui6BZrCwnG+POI4WlytdwVTGOQY8Qecwb
wPwYzaeV65B/dmHBZGRtIcn0LkabF1voaIydchnUGDg1UGvpI8RaeF+4927ApHu/
1cAROxHyr1tKwQnecfG2of83ITEjQ4jes1FJkZaaS6Ehgdhvwe7b4Il1oj1Co6nX
BWs0YH+mzVTzkskgXxhOAO5LjXkO9o58gjFxkEWW4voDdSqYszPbVOrE8xutSfWp
chV3KdSizwNEE+u8C/R1PY3gw4uUoJG6IHiPVXrb5ZjZLwWac68bgBMVsDAYZzSg
ukM7czEDEZHwBbktFBSe9WUM99Km+iVydF5GMePL0RB/R4Y77uLWle8nM6Auphiz
UntjXKptec61HAOhrHCGh8IGKYvW98ojlVSUDK0KEJ+GzZMJVqEJssJc70N6AqBY
9+UDFfXgM7FV2NWol6RVqTturqmxYNY9T5ijUfXwLA8QDuP3FVas0+QI92vJjBoQ
7s0ossRMumkIBsnHhBxw5pQmiYXRzKwn+9niO2e94j0oMsLQBeOFKIDuErIzypFN
BWEGGc2k3fqX7b/i2R+NuzALoXOgz/VmXDHXT2GYZWIWWjZa5G6cw20M05yAzO9e
dKy19boiqFZ9utllfIuiAvT4Pvm3MSiVGuQGiOqr+nHg6VB/tazY7xQo8P9KxEUv
Ya3/rs0RnK5QWZXyVn3ffXk5p5MoihTohjI+lqspWgrP0kXYAKTmM0yqDsE94qN3
zQpMavWdvgYnOTfaWr+ZPmpFlxaIrKL57MaUD2QpKShwKnOd79OezmDWhad/GwiO
s/Rk/MaSW5v1+ssZRL4NHkf8c3jI6JT1HqmvcvsZfYwco92iySpsf8ai/4npc0Qd
0SGpb7Z4hwBqC4lwbBq5vTJRxVV+6thgD9cuYwVcd1jl4CiyO+YXJXngpam9MT8k
3WcTKOJODN/jehyVtOzQnHNc1HxVzDQXfDO2VZAAujYYLmo6/Wu7DT0Yf4X4EH24
8L2nSyg0uiLbkTIlbClKKpibr7VmBKX0hIbgAsSJP+gFmrLINKdDv7bZhl7WY7Ux
wZBF55Y4A4jYxYOQGcKRSvx71X/kM+zENY9SH061IETP3bvyIzhoqfWHWY5VnvoM
Ku+ys0hqrDmi0Bv0Ne8MU0EXXPuaQiLZWB/p2HcGBqtPN2GyOZ8xb2OXUJSpCAxx
lV0iujstkYgXmwo1MjjOhO8Bx5jUnM/2n5j2aOcaoIU=
`protect END_PROTECTED
