`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kHX2hO6jnykPl+3yvc9kW0X5yj3pfo9WH840Tm26jpC4v85Dvk3tTkl+GWWzGtXy
ZgXCPloLSe2fDsR9pPtjP0BxZw4/RwFlNYsZyE3j/dca7wIuxCu843zc/zaf9kc7
baKvASkwTtCpfQYvmFTbc9ZmB0TOBfgWgQ/68UDlnDPVLBI5RzbeFTPLPbgW9NQR
K6bbT/qdRAiARW9hdpDeNPJApgeoIMu3AvR6VPl5MC0DGpfF72KRi7gS4gMstI8m
Mm+Jz3gJX/qeAnIsazmtLauPEynKjkOM+MGvTS51DRttRyqfE1h9y4D3+fqCPzwl
USFJEKqtv49H78kruA/5IV0MshxcU659qO8f8+gXPaphkIMndruSiJ6t/IAqRPN2
NhfIfVsckWvMFrmL5CbO2KgvzXdHjNjMNiZwTXqH7Aw5MhAXH5ZKlMQ9fdYqmst7
ruGhOr4S0sisnFSq5frd8hGADRptBGXxOFSTxr+5mamRqupJshdJhPez/72ex3HC
eM2CO0XZMlRkE6w5UxSk/cGwfmLZRDVfvHGLpDyQzmy3WSYb+lsmLYZuTIojM9eP
VmFn7n+7eleLhrGfhG5lk+CJB18PzaIzPK6SMIKqXhUsMaikwBmK/bY8hUZyh/8p
N9+5UE9vCMxq+e84Cy3deTQ2SW2XJmTdlVNZuqeiu4/6Tja03KijwwWWTHZaLxov
OnWb+wJeWXDqbWXrwnqASBiPQSEH3ySpW6RyOrtoNmaHf/Rq0h9oDPaLReVeC+8L
6UywntnEpL4LmerGOSokW3lbKkOMJgxhg/R4jY9uttCL0YrFESmJJJvSWUpw3JKk
d1gACGTCtqAC1fPdg/epzRsIjOFfjux5ErpSDwqcaeVhdybdg0iukcIZVWStsa0n
ESsAguWBbts2+vSbTxW3bO36KU9k2Rp81Z7iqQARx+QIe/0I3Asj//YjKU0EJNoH
FIm/VPg87pHhcjA+X18zaNHCnf6aT45ntM1mNWAnYz4eBon/JItTVF8JVTEmsfjH
csTbaBFgpeQy645RB6vl8M8I/IcjnE+n8TahVNmQoQ0g5oR4vvnFjKBOaOk1JGG2
a1CXNdFwZHFRfji6Hucx4C2EQrjvlZfQ2vMa4ei6EWzhfK7svmdCHBYYA7ckk5Np
roZjoSNLLyOfJ2aZizvnMAXSbtFSwN+ZzH7kvgwoU8/DFfJKhR33h9T56vAU8QfC
WoZTzXInsteTtbP+aoF1zxZ4TnLMMmUzoDTnKwE0zua9SveobLFFyyPMKoZop2a2
gP/KG7J+6OahWZMS+PLq+UsXI3yxkSz+YttsrleZV5A/yn2x2jGyHzqLaF4Lm2do
NyixXOfXM0n1Dyn0Vxf+jLPZ39oT9zm6FmL6VddhCk4evfKe7Rf+7tB/Nyn7nPFL
/wlPKa8S2o+gAbpLSZBY6TSE58F++4jeWOFHvjCEaSNLU6mEp13IiCDptXiaqqOx
aqIG9KY2L1X99CJ13MkMRw==
`protect END_PROTECTED
