`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
df8ZDMR0cpRTlGrG4XVqi2Wwoci6jlU99ydVD75DRsKtKQSyDxT7DhIflZL9Gr+N
qGlEKHjjVhXLpyWNqBtkaegUVzCJMvnOuDqFRwsQ0BWYgbAWEJ9RqVWGuljTBBeH
f8socnPIOVVceqHumQL8Roh9E4beI6t/SfkXSAfeQbEbU7yZ0LinWPCWiaqx7Yth
H4csxqUtqnQKhULcGf7YanrHL1tDYgcgPCZpyFLnlEhCt3APdQCqVJ89F1tarKK7
72EA6OlchEf/FM9CXG9rFyHk+VtD2Ifp+DG8AnXtqJ43zhEMLDvleUjoEggcgjd2
PF97Ltpwu6QCLtufN8rxmulkZ1quABApabhusaPrUS5XKjHjiMnQImEVk14NvQE6
wD2XFzbYHRwaPemhmaoh/fyBIfqg/86RrhtbZ6hJq8tDxE1zNek9dhwub/8QNezD
oB0aVF3g1s7EohVavBxom3sNDf7B5XgQhMO+37ejit0=
`protect END_PROTECTED
