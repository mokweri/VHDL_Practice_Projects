`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vV4xG9qagco4M/efJTuO8pEvcyS9tjeKbboLhllQaCC/O4dKK69jMnLqexaKYrk7
+9JfG4aWKNCLwBExRJ0yzH5QAO63dHckgw96QnZSwlmkYnb+hk1Gysc+qF3YU6ma
fEthaE0OjZWzOcUNrQhWkpAHNvtMkpFu1PD0TMXyjy6UnSFBy4t+FnBQNyeFE388
LE0IYY+IUXBk+2kXMoVZSQrI6p9oN2FjQBOag093wk2zBjksqL1pSGPO76j/AVZ9
ixYu62R1TEi0RJQGWeS45vP9nW4A5q2bfMjTOcFw4uUW9lxl6z11/JfTUxk1L2Oj
Lr/DFydcLJpTlaF8ef0rQ2wZE7Foj3/+jAp1LjVNH4IT1AUmcvh2juNvD/I7k4wX
NABkackQfAJraPWEXag7bDz7rKeSWd/ItT6ICtrsx7IdCB5qywKC3Urqo+YRV2mO
YETJlEj8U+csed8PHVtaeMcwVE6OTfusdqeeB7FFR9N5p3oRBFcjOO4snJT+V9FS
mhZmZz0MOpH0M4Cpv7VMGVJvoiJBZLLw+znnGhmMO7T456g/uEI6Xf2aGaWEo0u0
MFI7svCos3yHl/eW5X5iOjcX9hYflpDKBsmTsIxw+k+zttTMwns9MHbmcyAZD2ec
hrz8iOV0pr4FJpABvPgAKRaLydlB1E1wAkDmkwcHy4TW31CRVfIQ8dsbUDKxhVKG
ZWB3Xtzs4+yjWNkSMYS4jzC6fFbRJOaUKtkcE+f4rDml8aWfdsV8R5rRpwVeGS5W
BMQvtZuzlNUKbXH2XD8rwX7nHpzQlIzSuYWR2i/BnOuqt58mcgj+d4s5GriHZRo4
DJPzsS4lvvmvvgkCWBY40BfNaKwLXlvh+tyD2mcVNWnXyP247XnbwDUzpUKr8vzY
1BiaHsWiZYVodf2AncO9DsictF0irGUGa+aMjZ1HlmiwIJ/gYbXpXmVT3kelZy+n
BBMXwRCdgPI9XW5LcDgwptJnBSnoLHQkjNbHJd8G10hqTtN+aNoCgPbzi4kU4sNE
MGCveMJZGC5f3BGoXSgB5LLwEQQf231pv4LOuTnN6eMwF5TKiZkyRf9lc+G0oUNI
j4aTQhG2WW00k3apK5apv4dIerzaKKodsr8zkIfVXL3lHe58SFgzQQv4ijhTf03L
FSBsgqkD9jyq+2zeG2dST/N0CJkvL/91Wzfvbqsj+RQTV1E0pFxZQT2tysrk+8O+
momMxcngmJuxxvEEGZAc6lP3sXzmnOFpN+jj0HK7HIIX0jbOqQi1c7dsrWaATDZM
g3wPwAyHvP/Y0DxB9wFZmrU0HsioDkU8YPbfOReCPrOb+Z+k0vOTcLiALUvETQ8F
GOcPPJVVHRpULBM6kWTxlE8Hu7k5KUmabrl4q+THFAkN+/ceF+6aUpw2AIMmlMOA
tbASS1GFL9x4TtqsXnZQ4QwfS1lEZ4ptNAbc/rfLC8+1f4880WtllV1Y3C/PafoA
9nltYCr2T4O0Qw00h48YE+DL2rsRlQ6jUSI5XK3t9NB2BEQvZxXxNNDkxQGa/jif
57UfzXs0Us5W4S/ue9wkRx3Q+qLfjvi3OlTIeluWFVd9yqH2JCCBbkzWDroNMjdv
lgsOln+K5QYrPchIbSzaTm6GoBuItpWZwoDjuTzJid+FlY/2IrL8jA0sWPyId95y
0h8o2S6roL4KRcmaHYoimFA1JrPjNZjaqkqbpo7cwxTcnup88sobVED4mtz3hnZF
`protect END_PROTECTED
