`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gwReZGiWMGsFeHSyaIGJ+4zgvrxaXDASjFsiPToZTaKFFEyrcKwtr/VBoNiSRd8I
2DNAx4uPIx7cvi96RC6k3VhULDzHcb8G38W5GcdAKByxKQkbGZtNEBAgSyYZz4kM
VCZMR6eHPngMRtEQf2t3fdYcymcSoPlr48i01pZ5qOKffZidZXAa/8XLme8SnGER
TLg9ASZ4RfXD2bqkaqWeDN5RqNgt9or77INcHaduub2oRg6JhwFNKmnaBNBgJL7J
jSU8vNHO7b3by2Yd+2mx7XGBlSM+n85KprK4NBui/uuGiTuG+JOQOFNqywkhTmxr
38QIp+O0lPMq1yqinXhcxhGxxkWDF4CsfhreUVuYKSwZ5pXWxmhrFit2xL/EepDk
fUXHOgshf8hu714XlakeA5Bagvdvzckh3dMXxtaA4xlrse592HSVcywLwM434kJm
zQ186hxJR4sN1WasrtWNvc4lJKDohrA64HWpTPypoO6kCpqBpWDOVj9hWk7DWvr2
4kTPxLOSlIjmaAxyqSb8KLtFo1c7TPEiEvNzKYRxnmS8vQNj5fO8eMNOMSE+H20S
dwEcnmBX0vO34u9OHb4vUg2OTBQc4Sz/ofYE+wsMmFJsJhxBJezAHqJ21R9CS72I
9ufYCQBqSrwUFKDakwOfcE+17ntkbouiyvw5msxPWuYHT+w83LE52/0UXZTgskMh
N4ryxpt8EBHnjsuatJ0BQUDusWHkN0nqTvnHHycxE3PpJGw/eFvjXiAEk6D7ohiU
tT/hz5qI91mZFlSxGy/TEVpTwMkXHfkvPLXf3Shbw3+b1ZAthhwrffW+4zDc9NYd
rO0h9r7D5CIwFjeKzqO56aVPfpZUBfYVDfpa5W6a3vv1L9H5ziMbSl/3NI+URWqC
ZCaJxJYtJhegs+TLKfCDMfeg4W3bEQlZYTM6JBbwsGZ1up4KZBHjevm2FUBUnnbu
9nwrRPWXz5GqDNZ+jkfYLVoXYS7u7fjXeP7LBhSRO5klvfHLnJgI28iH2iUMLmh7
u6qVCTNHmk72K9mqkZyvuOj0lAfasnwb/eGuoRxe1w3vz4HkCe+H1uFumMCX0On6
DSSH8CzZ1PFgRYCkonMuqegZwMfSa66XnW8SuMLF1UZTbKwWnDIZrPluoExWFGZW
UE10EZVLy8/EWpj08PVX3YbCpalTvggn1kpSiKbnIuNoEkR3wWYysXWwTUO60Eq3
AZL+C4cY4gGy1e60pOAeAeTKiU8SlFcQCWgiPw3S/jQi0Oo+9Gh5oLarFs1uN6Up
gILII/DGbtiBqIaN67lj0gchvNbsjW8mco/GkdpMqsC/XIRtXu5ls+YxjtbaR7GV
tCiNmLi/bgQYwtmxGtMWKyikp3qyDCnt4Caxs9pCdau3NjDdWkb3PNOGtXJebly1
/lSRVrMD6WnMN4IZqAOZ51npUuHNytdpG7gajG2ttKX0jLfChM/FFViARo1o/eD9
7zpFWP096bOOsJmnxufAZ/a/LlEijk6feukOJlpw2eq0mDHgUmBewk8CiaxUgc7z
ftYMRo6DfUSX6JOqPLQA3SXQyTt10KrF5GBcjdFTnYhNtbWJfUUSIXP7oKndGwMI
XrP7/X6aOAEOtvIJPeXu1tn1Vj+b3Xkq1fmPDpyOOzAIRY6GtTk/DS24arlQ1QWi
/fpcQrWrNS/7DW41xitDQIMsBFztEwieAXzgcN3zgVKaqyn4Npm/zqAT5575CqbR
h/O5+DEHyp04oRxQyoi/Cm4NBAByCVi0zzjAnTCPe+SMJvwWNHsDYy1RPV93DH+b
VbytS/g4IqMk7ILtCOsLsVDo3533MNr06LUufnwHKz+YnKkdmXCArIKnX5a1xvnD
tIjidXRg0RKMlUWmixyOgt1/B2DoR5zUkJOJDAMAJGv6RlDcx+xOtW286t+WQQKO
LO6Hj2szTa0CmggB9ziIrRp91BBI2juNo7CQ+vJzvWISWAF2mx5dnORg5BHn7gcu
biUVRAFT71nwrArmF6B567X21hjUUxAgKV4AUKaZpcmUP8oxtPpb5WhHp5lXtQ57
83cgSluI7MSIsmn+cLUnqErtkumWJxpgb9p2HyGBSCc/KHJEVaFQULOfvQkdAP7b
fhSwgw8UsWrb/Jd8+orI6Mxkj3MWvzP+jMUBDf0HzdrpjU0MG/HnlPRdItAEYXYq
burt/t7kGzmKF5tMj/Jev4D7kZcEuo8VN5kfPhNpLZ42/92deURKY0S0B4FRtGY2
2w0DrIjRojqqw+udJf3yjBFqlbm8+bvBeCNtjBwPBgBj2LJA9f54ltfRq1knoFSB
mp3erBN4y4EITnzNTtthwC+A3Y4GbWS7JyUBht9SXidJvYA8j5Fsc1YtPoTVsuMv
8g7ay0/uXMDYwQriL4INmHUtG9LOQONFFWNqf1HiPnbkd/sernAi89WN+5ejUTrc
iAT9IDfB+lP5bQw2ptBh7qXOgWJK0POqGx3rAFjW4OMzR0HPvkV9KkhJaZiI4A3e
braCGveZxykhTkYB7qFNjYq67YnEnNI2eVpXEadyJULzKikULnagSC9Y2yiEj+NQ
0+b10xWr709O6OweO1p1PchITvu5zsiLRzeFIj9/+eJ3wrOiOduGDsz5jc7Lx2rM
QmHsMFJ2SuFq16Oin2ikYWUnXUjyDFucoPhxTuzuxS+Gjh1yQNmDDaKpJQYvuRkw
mjqQEU27EpQ2Qv02QAEQPusuvQNNie5VhNSXWFz4EQSCRYHMRRNhMYKXYyxziyEO
6bD04z7FU+B5y76HEwqmspeqJllC8qDxnn/994aEdMEqXjNFQQSQG3dmHxLXSvRe
O91K+Urj6b/0UOV4MqhP76gUar29Mn64IEdWyA2k6NbN7dMkkmUZC8xlpdxQ/UYj
Ka4rV5McdIKpUgTD/W0noVDjNgdLfHJMc5SkiCFuQjjps8Rz3BGauAyoyikjcdRl
YLxIHAYwclVv+2nFlLzWntANFJ3OJYIqKII3bQkCGHr+wEWWRxDZas2nwKWfnjiq
vNIU0bGO53nzl0L1/7sGH6/oisu3wva7VnwSq73hhfsp1HCJoXC3Psfhwhiuhr5I
YpX3+YjusowLNJKUITqJDnatkLmJoj5/fQXJlXMTExwfUgCbuaDrbU67+cSaWzDo
LHiVGiDz60O2pbj6D5n8RYkg78r0BIMCRyk3zqijupvtEYnoO3YSUHgtTIGao4y4
P+WBvJTYvmTkCmDMfj6fTqPO8cjEloBz33tn25iJTNaMWasAFEphXmcJH49EC4LX
2TJwTUbaTFmu4/xAZhOKtpuJR/uCMA0RCO31XowoON7z7y/DwlvWUqnCIrl9s/Fy
MkOcn2HsOI+dwmcBFK02Qgu0nd4MMAQnFj6onXadLpI4UVI1S/ntZobJlR+gI/yO
ksyQfEuDwzBKbdDCj0lqssUfxm5dN9zxMuTQqVYhL+X2wQFRPrLv8Paxaaq0GQML
eOFd81JbnXR6WpVE07JZU00HUYLn+0br0i4DtedrXR5tUqBCm3URWBgWybf0KmqF
x9P/C+UUfK9zOHW69ILQdJD6CUoNjH49cpvWdtEz41+szO6jp1HAwMCkw897KUzK
auGI+/1kCGaTy89lE2HKH3z8NoJJo9m6La2YDOvui3Rvf2WQEpQgayL3kTlaJ1Qz
i8UYSNClWNrbEaij/W/JEnhrGH776CbSo8kc7zF+BIZT32lvIk8i0g5bJxfC+ml5
nPUcT29N57yECIQmDkzD51lrX55EotlJqdt4hJ5HetMLSQlThPY/w9n7wrim//pv
R+w/zoGm/r/2KMJFZpFiQosmsgNU+8AKDrgURz8dzHLguw6b3rodTUE27x2QMWul
qrwKj6ISQnAUIGfEri+WwR+XbdtcABp5w492MWUlZg3hJMyekatQeGDY4maausS2
aHFO2VDweS1e0VMx2vq7XM2Sz6NTwAvB83hSJ9n3h0IDCiN4RLmAyDSRGgJ4CLJG
sinJf2qA3qQS5kn6fJNpeVLQS94LRmv7OpWS8aWnUk60LdwGuZ+wH/OJjSBAFsgs
wb8sYTSJojvufOszg9ugKa37x6RQJm7TDKOwI/VkfEU256nMvEVMcI1oTeW8w07d
EheKuvmxuzybjx5o2WDKOyX1+Ps7HCGVEV98zjv3mxgh1E/QpcYYGvZualOf/9mS
h42799ZkMwtbufOYf+pIyGrZIqAqgZuUtT99ArulwwiJePDzdmKly0nNB1aeHTqN
AfZfSVtOsM98TZMjMhv/nYlBu0BraP4FnHvdihrHYflo5eTTJONxql0K7Ew/ipXM
CM1piv41ExcneSBlt+P/SXA8CrAzQg3mYTTIvmd1Sv1rAiwu7Fr+dpzQpehqW3QF
hE8wAQRiQVPuEdr9JxaR9XTq+tKKF0zJ5p5ffH1X/kIEYkIsDv1B6puTYIfpsddm
sUYzJp9rNkzg1NIO8AykLsf6G9NdoC9dtaXn5I2cExJdhb22Lg4EhD8Bjo+BNwyH
dUnZS8tw95Beghn8pFT0KG1fU8eOzNOoGDp2v7udAXJEt6LbzvgbHffjA3RgBWrk
76Qk3jEKYOYIDCgXtVLSB+5vWKel2jXwCw8A3W3F41V48obrcmwDxBkgIZMJmogt
AMeS3faAMVS8tduM/B7UoYAgS5if4J/jGXPGoDy+DXPXj7bbL83+0+xsbZ3Mcc0A
IsvfbvYXux70ByoZZKZS0yhr4ZEKv6S5DUVlAoSBv5P1ibdHAA4Ri04YnEzDkkbc
hyvqcnObAFwvRYkTUAGLEPIDhgZzRsbOagmvJKIsuyWmFgp+ezhHnTNKCzM71Bu0
vcx2+xfAz6Hw0wXCF6xbcqDCHVjaEbvUIBVXx/V+7lcKzDW7Ac/608Fg18M0RVO7
zcbaNXa4OKbDb775Xj/CbYu5nvV/l848d/wDVmuhOGAbbS5p1clnSLGs+OD+dpFM
JQREjBZcGuKwqNaorsusHlAlh1c++cZrJmwev6IZLUhuSCVOp6H9IdagYJLaWlc5
m8KnMkXJ41VvoTbr+wb/2v7y5h1YeiGtXIadgcoipJKFBHMUk/7SdVB5cxqnS4dw
l9JqfGzSFIbqCcWO3kAqhpTE8nHmytkczX+1sKfykCDZ6Yb+mStU+T8h8OmIqbjx
ViLR6f1QH2sybI+gCCwcnx7ZwNNefDTRuPpPXkJFlCZ5M8Z+p/fAyDe3iX3dFHfz
5H+l/+T1pbB+FsUFxSuW/8uxOxNBevBQ7dgV0F3l4BA0Teh2caSXLC6SHV1Wl4MY
pdKsQtb6ES3SbmKB+74IPgcUVvCKi068hY/7aE80+fRVlMFxU3lPUmORo79fAqId
gHDnFd0pQe2FJHikq4euTbNqruGTPAQDZ3cUAq0qqZzCyUft80cRVsCZ/cOiGU37
yBGwfM/xles26BTf/8GEU1ftmtIJKeoFJjz57+D+v2wAYbnAGi4DaRX2mGeUcFm+
3CTWhFN5oc36v8nQVrMFZ4LcWyTJ3vQ//mSfG4Btf4kHhARHABFMahmsOz/DviDX
A+q8b1aMQsNuwra0fJrtH7lMoPPvCxEZOhhppfacn5l2yCiQsvmCCYnkOURPGGX3
iLJec5qQe/ZXp8jDVrJWMfCy6lyLrg7l676hFfkw5F4X1vhv1iwUwhSuChF19eWI
4L/HDDAX0ii/TnwlXubLcTFoI25LZMnRreqZBm7Sqfj3zD0umbVWXwYxpCfX1xnp
YPd1T/w8YEk8AmKS30+1c1FQawgdngRuOhYjlwpIIDs/5/Kdp+bCykCp43WK7X8Q
4INlBNJUvORs8uwTaCkwQcxUm/3sK+nMTl+PmfgkpuY8cK0vjvrfarudnax1TTqM
PZurMFqUus0igOgvv2D/Btc+E6obWjO0oBUz3fveLg449+w3ku8YQkfP0GtK4CBr
IAgBC7LelkBBXS5IbOYDFfbDfsDUO9bW7/RW0GgMeT+Ehh6eXoVEKknTz3/ou8fA
skmwa5y8Lx34I4YwB5D5N+Ta/lf2kE+Ta3oBkhKtlO07vVAmEUl0T6qepubpQqdC
Ng2k+gAOZm3ulF5IepFwbQF87Y69NJDlPOuylJhFwJXleg76Indln5P5GlPryEqI
ReGa2DC94MqLl4dYbZxlE4BYJWMO0yyGa8+tQ++D+EI6FqQ/q+0l3AhP6Githr6y
nZjZf1ltXwhb/zDnpc8G1Kq+0+qwjXrZoeesUy0NFk+VE05rO/iR47cu0MkFWLC5
YclWevFDg68cX/ZGtHppOizWMRfIgPKabozo0SJRZ+3iXCO47XoHIyvHqZLxlrmN
ywAciPfjE1JbQIACZTcpEBwOXO8YQyzBb4/2BdgrLo5qZj/JBP9luh1lj3f8yXbe
evtevg+DaIhM1EH1mqZ+t63ioDsVt1pCXsi3lfjPSRtek7x/gwHHD91oCDV8/tbX
tQmbt8HeCtD9ZN/dx/Xx6WwgaaQVTTHgJ9Bvitv7Hk6yvfgr5YTBtw8zi+li2SQ8
TgdpwSnAhNRWDaZpMzmej6TDkX3+rnUnPC55Xl5ktlOup5BBi0EBd4Hj4gHE5tfj
5QwVO16pRVWVfK8uepz0mK/gH/huTP5aRpXmbwVvG/KefdQJystn1BwC5TDgpDVx
HV1M9/t/Yaol9NvsVPEG5CDh73p0/YUvJa9hYeRshEuvdaVJipd8brk9MvpONFs4
65K06qB1SfrsqG9l1xiQX7uqg7yGHmM37vqvSecpFvMakH40Mv99feMaUkLvu56t
qJaSrXX4SZkyqqoDLiSeccJ4vfmP/0zQp8F5E4NG/KunTMi9H+A3i2YhcLDiAqOz
elP8TSKnz+q563mCpS/3dN2FNKo9ceHxTrdR3eDiZxxaIwQQT7rLm+G8k5giH+0O
ii4Fs3zWoUWe/ZmoNW8EiKfjrGr2ahgqrbg5c0jniwyZSXx5uC3Gu2E+/LNwJPxt
UV0aZbQxfxOve6g5jbw9DKZtJQpEqc6LqASLFPLK7qftn85IuygOReR5UfDouwfD
pbp2esTAR8hCYKOEnb+vKLq80cbOccRfkOcWZ3Ir89Ub8yK9coxbCAggyefANFXs
Oup33XTBY9Ot/j8MAV+aXqeflLSNeNAEVXT1XTPbcrkgUIhffS1BuO4pA3XFHvGL
hgGVG6TYc9DK3xBxXa1dJ8F2QEa9mjYxwZ4F0/8caAGMprsi8fP+9fGBBuCpc4zL
ECQVVskQ5hdR0UES0vx1NMBBGZhYMP+YNZSz5chdfNyvTXch10xCbPtemv29hF3H
Bd5PpHjGPi3LzTHE9eF9nDZ5Ib8/CAJ/xp0EVa9veP91v9os2A3xcoJBhuRdnMdt
zH5zcWoJDzLu6xLiDRJ8TTZIyccabGu70hkyUMSmZ0nzwC7SEyherqVd4oSKSUY/
+eqazWf+Sgi6rQ2DpSUkQ5UShunGmicdWrgfUPpRKhKf8mvNhtPErmbtfGTwBNXO
XMrcRUZgjrcT7fGNsCAQPcZbvRAS4cgPlMMZ+7m8+SdUn+tKsKMd/+pFXrDLXq8o
cMxzbenDw/AB6NIMzfsJ143N1fF792Dl46YTIE4wNXf7jUCdgfmjCb+3dTukd/Ei
XL+gMvU5Hku1HvsbSusNsOJt7epbYbHsddIdGk0UX0Bmt4ZhZsnnve9cbC7ReOnR
Ocqrc0nVLn893cvNLhA96wSMjKBlZEWcH0QbAV3OEF0AHfikn8pUxRZ8KrxMwib+
UU71+4tEydmIhrP3J4AumlgKY0Tu9iqvYL+VHoRIzYlMK/DFj+M3JNxGkw5udt9h
LTmtJer25s/Q1lph8XWVAvXF7L5PQto5DdS/uzGrK7Hmwf37QJr4WvijipAX8IFw
tLZd1e/zVyR6B9lwgQ5BOkoSSUEAtp7YLnCxR/bTo30smogq1wnakeB7iI2he8TS
MDlNc/YDZv9pvXRFF/IsH1p+1yGRT+k+i13uEEhYdhM45gU5JBIiAhw7JM4gR/iv
bDGG+yCOHk1S6vfLgUKljPVGdhUDFWjJOeAS9TPq4FqlB6v4uVnKoFJHLaxjj88O
vsp+4NFhXy5kmW19eaZcBEt9GOzRnADiHIyofvxrjqZFKV18Q9MPbj7dXtDZSeSR
mXk2OP2D5foKm+UgHoZ5EUu0nUpJf5ooJS5+ubQLs5SVZJVnIjjIaGkmdhnPgsqL
1K3riw7vyevUKzmCrq4qRdcUpAyVncfW5bPMK4usgUnG1+ULFYpxfmBf4NaU5opN
Zj9b0dT5oBvYU9k8Reo4ehL7COpgcYNJFux53nVC8m3MfNIzsW8E1T3FSVNlLz6E
4hlPs/0qsdsjsS9ExKmrep5+2y5oUBbdZ4AdtyI0vfPNYVxbhpW6ZLnxZpX5Z2x1
yykQ5765ecEJJ07bVo98Yj8ke7rQVJQvOwfcxlswXdjrNoAFAXL9n0wW3UsC7RoF
cJkXMT6wVKDKeSZRIJOTsrCiqxMlaMUPzEF6WK3xlwSephY6+YLAIFiRUKg5wnE9
JirUANuOKNXd0aQ/wLL4Jzep5ducwd9Vq9JJjWW6LOlxB1IMhm6MGLqlb66gpVTc
C0Uqr4tD9Zj2jxq+pR1QeMePvjImbOa+mZ/jFAxtRmuSXNKMXWqSdGdmwIWDUrN+
q+yWm0lKqXjOm9td6G25HORB6IE3ilHtAjnqLGJdkqX8H65l8fNFnRXesTSbb0Ey
uUYf+ffwDJksBicg5IIBBAy8Tx/m48AYF+xbLKXStTK6NytyC8Bb8w0oQZYh86dg
0KQBvxXdtzZ/RFgOev77L8lzKi2qdgWFjzZuenNQL6icbtRiOm/+pqK02t10QztD
pOMn8smjxhYZCrKRlwtma02fxf6XsFpEItjrhxEVxuWJ+opPCYifSzpJG5EAs5DY
TaP3i4tVpj6Mwue2Xlhz2F0Z/eTnv4RBjqk32D1Ze+7krJzX79wAopu/Z/QHJkmR
8AmmSAtJLshAQl8B5lMpYsDom2C9FYbDMO9YgVE3k9S9lXUuv38njkvd//8gA8WV
gaYm6mb/eP0t0nmx4oqlDseJno5SZgehHMRi26nZtJHpaTCAzodYJ4NqIDOv69nN
f3x9IgtpQLwgHUmz12GxC/C07kmL6npsnMSP2RYm3NCdtjp8dZuIWmQKiHaib0BL
3mAWCbn6o3s/dnBT0jDOA7aEQe2tVKqfpM/3dAB9XkgvXkWTZLLoIjQ3LQsq7wls
rdQdrfbEDuz2tAxUnil4dbP37Wx1y+2/SkZz1p9jcg9SKKjFBMQKC53a50ko96lJ
wLzfe4QaUcoKVsaxfWkxPuXc4xlEOrUcTu0jv+MqvXI/myyXAgbJ16m69ZLppqLD
1RJX/Xx5Hf0+D52GHanELRfyi7waF/Ymj4HDimWUXRjtbHn6Dum5y5p8S6EhjSri
N+1GIEs2i5A12h4p+d3nuX7JOHSdSHP+FtFK3S9ltX0iS9UMzc3ci1TheeRYQi2L
a+ySxEX0IiOQF5RY30CBbGMtjDh8ReIRzU4NEBzb+j7Sjss/v+9nIv1810B4B3hb
9vpIBLrBLeNgCbeUrTNn5P4s3tSfT7CggIR+R8Dwb2BWeRIyOoeVmgw5YBTksPOa
qCxzjS8UY9DVn+mSOP+RAszPMM0ULb8BpAh7P0v/s6xhcxZONnk+w2UoOK5io+OW
Pchhdkjuc+phssDbuDxkiFozQ8L9aDfB9GQsJIX3jXcgcXcG+nqUmOfk8jCFzJXL
l1RqYJu5+m78ZTPcPUU3Owx1TL3eSrio1rCAGGuPlvgLwMxd9tfe47rBsXNTj7hw
206oT6AvmslLKH+Tu/rQONsA/64Er1SG3f1nAPa4ThsT/pzA5FXAM5C+o75wrfl3
Oo26PFBkjDEaBXQ000DOzfH3LpyCVc2S/BtVSYOaxPUOC3o7MSBKtnmUBr9BnbQ4
aZiZzpZUlAd0iijeB98B6ztgnfJ/AS5ZBR6uu8x69npNMluqUtC9nGGpkQScPlqf
k19wbvGxmGVFOoBw1lr3cjb+rbKk5jOsa02bkUWHMMY6Ek8Ic29kRmyK7S8AH8Gl
Sr4c11f0JjOb79qlFAnR9/8QyFZrATTG4iUA9kVlep5CNYCW3tSrXb0bgBfHO+V3
wT8kSHoYa2iyxE8Bs5WQdyjl4Pubn8FYLmOgMOm2n7zbVNmFSannc62eSpZyVNBK
yL7aPLOhH7vWsC/Uqwtx0YHj3tp6VMwYOtOV4QELLjFTT6lNNI+kUqyGrdSSO6ft
uRQ6UUYahqDLVqazyQwwcUY6/Cz9Os3+jZ3NMx4ilL1SAtC/6XYB5y7GZmfMvOo7
wRrcn1CVE2hZbv2WbOQVsRX4RXZx++TwS350x1c4y4SuJb2DHVukNLM44rXjgrBw
LlzXoPWmYXmuXxAcv5HOi+pDY9hrO8eheL4Np0zeXA3zUB0RmgYjBJisccJYImDf
F+rC2ymJ1Ug6avalARb5YAbSSO6d3/UOT5SZV/2FRvCOQach3uEIMWlSUVCCiT1H
U+oeHAEbpEX6jusl9bvdIA0XPzSDTHZ+oNXMw2lpljNCy9l8qYs1WgsAlcHXBgyX
ZxQl4W9rVjiKWizIuCOAHwDwUc4s2qJpYIP0iZb3gIa0xudDwlc4AcxwbCcPr7wp
KwVZbStpH9aQhiFDB5GPtMAizaZYVTRKY9SUWjM/yuVqtQR+YC/slPoTDit0kfia
06ZeY+4GJIVJFAOwIr1udDzdAAYFVKAYd2GrvYm9zaYPdi5tJq0yGM2ojthNYPu2
EIlVA6SSc7ZndVWyUTIq1g9GeIsEbK4Sqg0P38tjZ98i/ITW/3HIuKqoR+x1GxuB
ymqGSehXJfNwjI9MPeBhdqTgiLpHw1mOtUcMiR8cPFfdItwiSvLwfQmHAz6QItvT
hVm2yfINieoU5uo4yr03tB1YPuR1jSYOasB7yvGclNNQJV5vEwtRY6uifXCTU7YI
XS+qTtWrtHsfIQba/Ed9Tvf8VYYbRnZ8weiMSv5BZE1jtFQW7c3X09QR1Z9dZ9O+
B80oDGptZNxm0ne52q53zKCamGrAH5Y7y8A9h6v+8w8rahpuAr+08j4Y5qwyTHqR
CourJ/sF3NhhePF2eR8AgsmFwsQi2cLOVuOXM1yeRCzgywv3ZJQS/GGF2xGoGPWB
sNq67Vs+OqRdnPxnmn5sGPo494FyQLIQKWzpjAnjo2YppAHl+Ca2VIC/bc1pn0Iu
8lpqssuP428aiNd2FW+ZZ+/e+53WcF9eTak3LmkfxxIngxrNGdFmfv8+ezDApQWP
7QZUtspzNNfsX9YitOg9qBUlehOdyH1SEIVEfZbkFomKBmptrSepqye9T+xp1U4o
3DetTMD7f6JhZw8VDxW7ggpLbmy/qKjIvB4BoNpySBkpueOYNfH8n4PiqwgHr0xI
trErl0jYJo5jzvM5a7B83YjtUNTNXeR+5AeacBTUDNUBuDsLCPEvuVyGOiRRoRDy
khqh7oDrrACLMgcYg8WvC6RcRLj5sQKZGBMUw38NwqmILC68Rckl1nW18iyN9qPB
cyNn+d6zL5wha+wFBvhcFxiuKVFL3wMWYQthBf6HqBFCx653GYQx3cYRCa3isi3X
ppz/wpzDoM6fr8qkA4v3+jyNMgAL4lCP980FP22d+jOrSFUAeiIsmqO56IJ3A4HX
pDJAV9wUUDc1WF+SG5QnaL9oIjZHfQcoEi3bZS0eDGufGDz7zHrigSV0GMzGH6cH
21OVck6kiP9wEwC9D4oY9S2Y/YSKfr0nP7nOyAiTXPd7Yxx02ZdoC3HHSF9mVdGO
J9SF5XN3qccrtHbTNT83zRMfGotFXLhTnPaWnWBOnlgj+ozoIdjjthcnbKzy7aJJ
2RGFZB46E30M5Mu/qCAQFloZZl/XooY9VjX3xLBELnnXHaNGC5zl9jgYKsLZRykI
KlOQCZh4OLi4wklNO3znujiNLkZTI4ZigAIrQVNPGAlSSJi4d0FgrRmGoeap02AK
1YVNSQB6onJ8VS19Hr+Vs9NCzmDMlMQitUe2jzGnsNiC6tR1IvsesRHRuAtKieRd
z5VH61ir4dB3sDfYzA67/0o7tHNUIb3Er/zilLHJVlWXC15zx8w9CpRrwdwV3S6B
V013MbdhzWtp8DwbLrGCaSwwykMc6z7VlLacda8bx2gIs84JfKlivQV8yq1OMe09
IJV4tUUohiVig9fgjHGyzP6BxWOD9XtaOi4RT7FupiPKsuGrTrPWzXYA1fgdsqjN
k28zVKJZh1G4BiaY9bK7U2+Bi26alGSAsQqYUNUgsYZIN8F5uuBYzobUKATtKbe7
0Yhrnq5wMXfV4A+C+9zDKtwTF7f4RW2l5d0GqvH5mOzEp/HJAvebX7vRooS0HCW0
M3miVMnWU4QmKfQQiM9DTDHyZsn1/XkdxYsrV7RsMugQdW+ElwDTKNUR8YfCtGbR
HX4JiBuo+bYqi9RTHBoGg2pbNm2mPwdwmOfMzTRZhwoyzAFOcC2QY+zx3ogawcTm
Vu77pzVV1wCtr0xqkD8DbuRrRJ+ckMTyjeBwGRXVMpZe1FQRVoTojU+0+7/q8EOH
9XSD1xk9riR2Zyc4M1gmxTstWQBfvb2s1eFmnP6A/5EmT/TC7hAF6go7oR8HcvB5
OTjJ94puG89UgPzAtVCxTK7U14oiNZrIiae7iT+0WMxRiP3M49I9tNJUzVrTvQsj
A+wAZGrBpGlBBcQVjxsJz16/yyIopQz8SC8pzOtgr8cETPt3BkQ4uIdmeMMcQYJZ
DtEYGZwHxw0KvkugliaWnQ==
`protect END_PROTECTED
