`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukoD7Npv4MbJ6ugzP9WnygHQ0VxT0kBnSG/P/4OjAdwVWpxLeLyMKDerbp7aFosy
eOW23kjYrNHmAQ6nqxsjluYdHgW+OijkUC3KeUfqxAJwnQCqesYEjR89u0+zNvB4
St1NgXDZupmbwiXYVW4zM7eC3qJJd3lEpmUoigsiT3JtxfdP2bpOy4z0to+x2n3d
xU+Zc7Bu8hY4qEazKnImgvsKO8FgsAHbG9Dsn9iUiGWjcs9VYe+UD3zIAc1/RsYT
nYtfMOlRY5D0e1IUMX+mkWM1DBMykPIMHaa4FknzUrTX3L91LYUGXk24p4xJ9MOy
Qwdg7j0skhTqWdrAeeV48STfWgvbUWV9XEnN54V2fnHlcGdnrI9ai3TFtWwU4DyW
HGpH52uQEAtPKbuGUug75SdCmqqq9Wuex2AlQ2vXmX2pa4YGSxG9XWww6nLspuhn
E0tYyITra1tqkYqv2mgqQhSuTGJ/vuMqTY4BRgPz4ck2rHDn2uVnIfi2YcOsRVFe
z0bmJjqS2MhrUjm3vw7Fx+FwK7jBA1wkdF9RLdJbr/SIixVMA+gDFZnXF92/ex7Y
HcPb7duBXPVEzqvOWTqLmgvoffYRpZWyZBEDflJlMd1ISVtA7sdNDpcJxreQt823
MfAOeANY8qv7bxuu1UTcM7NMN9x3J9iqFI5J/Zj+SSZYtULhXQkjwyaq7Op0YxLy
QCywRsAuS0vn5uclbfZvDEg0T1QjKvmV7LXBubAp3uDbs4crChnuR+gy7xCtR05M
jL/rB7HSeWdIBnPvemur6P+liZYdePJtw88NKnMhinOtwNJ0bDF8HN78llnzZCPs
kLKlBRQzNmfZCo3TO3NXt1aZAhJMnkjYKusOqEMNkPYYlCqZGOsAoRCJK+mj/wWF
QxUwAmVv7wOe9Ifc8M7Z5QjOlmFhwhS0rWlGTLeWCLguiJjUkd9UVgO57i4t7lDl
S8YcYHhsH7xwHmbkWiYCe8moilbZurpSoPUAjyIaMpNMdSAqU8/+Ms8IOm7B668T
2uXXPbiVL5YsWhlQPDgEQ6wkZnQbg2wbGvoWuHRt/n3VVP1jRfXn4V1g3nPP/X7K
hpZoGU3q19GhXcMA0GtTAkxP+SpQZIk0eNFXKi5k20SYq4VItWR0DlMfQPYcylFi
+HZcrdCqk553z4xHyMQwY4q4mmn8EDH6i61m/43WEuUgSpT8NsSYzbT/u7CK3n0l
MaooIHqYz5+u6sQ6lesD28y4r2AEUwM27XBL/81xNfMQ+yMj3YtlQAHHB1MhJM5n
CIjGO6vVN4RoBRHz7xRb8kAlLvoqR3tjJaCKNGDjBWUkGOJnXtB8OnDklV+rInto
lm4sg7h8VptZjAVCUbp7SJldrRvXWXengHHyL50nAMQX9pePPBu/sSuWf7yaj9iR
Kz6uAJO5wI/IhhKi1kHDlNSqXmutZRc5z1w8pGyV9l2QuBDMZLuLf3uTUeIPTZH5
d0Fcumrg0YmIWxAJTauk02aOXRrSyTd9nwZKidve/52Hs+5gfOU73FlZQphyYXwJ
fZM9KQaK08HXBua9kwsU0auL4jrXgFXKyvRrf2pI4FisFYqv0r4DpBhCUTWkO14x
IAFgXVK8MvrIxJ0O/Hnf/EOOEV9rM5p4QX14ZaQAvR+kBFqqi9RTdnF6MDqs8c20
OLD6un//PxOEGh7LOt8qPA==
`protect END_PROTECTED
