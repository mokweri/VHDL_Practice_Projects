`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FXdj7DMcuHj1/GC5tVHAFgEM0kk+1YlSD72aVYj//0NVxQAJS0zBE9j3ObLbqbkw
gN5oVIL7BuGVPzQMSExFT1UflmaEMoQDl9DPwuWi8cElnHiWaoLrEAt/hK31f/ek
5rlY0WmTzyf5pvIX61L1v2hrYaxoP29aeEGYInvFngXTcZFs9qzjlTn5+XeUXzhz
9/c256r7dKS0bYoTn98qJqG2JbURH5rQiJx/8RHF2n8YUB8GIDwHIW5Pkq/E5uwN
qfrdAFIGdecMhPISDl56EhAo8d6cf8ccVZByAo8xdcBFK2JS1vjIGl9+JICFq4yg
XbHGzIcL+3T2wFU8Q7TvfdRX33e1I+i8gHnB5MRGT4bE1m9polwDu3Qwb7d7ZdJW
1H8PQtEqyN90BHyeCouH9kHG/Sl794oi0OBj8HAnMng2Gx7G++NnOZfU6g2Tdd4q
e7bMwXItK1/fXMqawyu1m+8J+SGeaOC97Z6Qzp36oev6ZrDktjmuqdkEDDTy7uwc
jV2gtNAU3uHHlbE2Mde7E+5AMbkMCzHGVvxFGyGyNsKPhlfkfFAMKc4OApkoEigI
WpUlfLyBTpdtTtDJ0F/4kNmadwpT1LAE7v5c44C8c0dWjsyMR4i4GzOyX7QmZZXp
qF2bjl/Z+0CnSdeZx7h2I+lFh5zMxZ9MVrMCAAs+FMDKQFZOgNahsbzornxkb/Uy
5WdEEKBr/xw3MU5oWxT+CP+fe3N3E85trvb4lBBgkKlJFR04fA874ayRzL7Ai+3G
Cpb6tHURBB6izvTCJYPBMhMWiEFS4zFNtrUiztm5drx8yB/UwoxrmYxuTURkImrL
ImFnYrGGW9JXu0UNc+LTWtdMY25hgzWDkq6FreGjriSnySQOigfWclm9Ju9wYKnC
Dl1G5LBDHcEwk13Zqct+4FI24WpYtO3V0mtGl0B4UVGeNor6S2mZtG9ixK8aYzst
z5SyJnW1ito8B0qUeoqfc7TjMUVIz2Vsg2WjC7nCZcKBtKQ32C1x165q76LZ4Al7
71MZvhk3Zxp14JvPEs7aIsa54S95j39o+yylgI/s91n9zSgTdpKGQi8C9L3ntRD5
o7XncEw+H0sY+CojDKaCx9BJZl7FAKzso0wq1sIJ3+k=
`protect END_PROTECTED
