`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+reuIyDUC5LdniMpCAhV5yBYj9YbDADKF66u17Wwxs/3vPlha+2ZpqluGuMFot52
2E3PrPIm+QoJVio1SGxduvBu4SGxD2V6SAggS4nkLMlqJv1F8RV4rRjnzimyt90h
vxIjU7pbM7gHzet4kfkLCZZTSAnrJnigCjaPFClQfFX4bkGoM7sZ/4TGo9UnuFfK
9aIfCJT+98CSEXuA2hx6AcOER0yiRZtrM0rDfjNJr5TGzVPYzmL+mA8CuuTMCdzC
7rys1GgbbCnBgbXwGt6If9wgF+54kqGocd7/QWm0uB6iRUpSuT/bqrk+3+ktZPuI
WWUQp68zLvA/18gKypCK0xdayX6ckWRIZYFbGcUc4MQCO2GWbRKLqheqIhbVhrBm
3dAyzr2i0i3GraJCye8Q7m7427I8HnQSun6I3Bv1fJ66vXiLykjZnGqZfAS/Vlg/
oLGImK0ZIPSxiMYLtCaVmdNeTX/ijP4hrbyP2g72rliZ+JiiUp83AjEedJoAin7/
ElBEatC3zDeS+FpeR46XothBduUHKMZkl9yh9jIU5+38GEQwuHAaoG+KjePvoMw1
dP2EFQm3qQEXS6b6wmZNKe+JfC3TZnX1+90pRlT64RQUtwcDEIyvUmvcxDkmFDWR
k9zx2o+msP4WyusiTocTBESBqy3dblNh5Y9LRDOqvHGy7Tn62w2Cj7s40/ORt+E4
eejVrnZHK8yDe5mQESd9p5FuTCrIGY1rHl5QmFgQJ3VPBQJEt6cLeWw8scvmYZn2
3H18gt7eL7SbDVCZNR4ZLvg8I3gSUpV7/+tLDbyZdEfchOyDW1k7D2bvKMxQ439j
1ce6PE8ng/bPZcr00pM76Y87PJyPk32H3Dvm+97lfIZQsyzG6zEaVVCfhxOeunTF
`protect END_PROTECTED
