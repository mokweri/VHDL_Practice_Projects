`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mp+9aJRJ5hlx2Obl4ujd1rbWc3+c71bjpGtOOnESPP95tAerbn7Lse/SKXlZmBua
a4eX2YfDFKqM2XGdcDYUogv4GbsKTPmv1ieOL6QFuhP6gbslQ+4f4lV7AFkyzLcT
eGHOLrAT+4PGWPCR79dA1WmFoIAI2RcYPeaXrW1wymjB+7pBnNQXvl4vSwlt82TQ
HhwcuxQTiFKycyYfcQogfx75kM5lyIYmf8stdJohijgzP20PwBO7GrWulTTp7ddD
Dw9o7vkvoX1VEJgz4K9hU23dE/iYy2DypiRpVIaR4NxOJaJExgkk4SXRhILcoTFX
hVpyUOhbSwPk8PnBHwU9hNy9ibnwDmzo006oRItlsqu+oEM3fWAr1igN1efeK/8P
FX5UyiriM2EYbjk+8Wfr02qq/D6TFOAnpnohqshHl5YJ2FnDxJEeJqThKb2TuRXn
ixEL/YqVOtp8cKfyGBwtS/6jcQmSEAKmGg1aSLSnex0ll/+DYdmLkRq6d4lTulFo
SLJ3li0TKb0VooVeDLP/vxZ/4cjDAHaI0s1DlqVsXAA=
`protect END_PROTECTED
