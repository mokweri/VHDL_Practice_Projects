`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GTbRtl3lvuByx1HXfhbjct1ywHC8WjKgmRqZi2s0d3DBEJ1pvXo5xT32qQTtyxv
8NrHVMXnZMuWFlrezufjRGApL6GeED4Mg7Qn5XQsyC9lTbtQAMVEdBFHbnM4kjVc
Lhrb5y4nP+rayHrsh5CRvYIYh3gBsbvL3xCADVpgQ64ejH7tjxZj9+iwmqtbmpmW
SaJpU04dH8CkgIm56XxgioN1YeB6g8LQUQi7V/VwhvZS+FKTXyy7zKAFYkjiBvHN
t6ab6By3rS7Uxe/C8fTCQOyFZhW4PkIDT2EsfPkTBpVTt7TdOzQcIkHq80qvt/5J
cN4A0AOnPJkuOLiHY3SO/zjmB3ljPN6l66kXwcSm4t4KZ5X/B07XwK/35fRt8Cvk
TD4EI4NZ6C4hmxZn7+v8XbkjVuE8lT3TIK3imBaHzmhe5nYH+GcHEMd8088VCkkm
HmqI8ku6waFaPKKTYApwJDB4J6rK3yB1hfkNLkBVIxYbiXZO0QvC2NrgiQZhNBop
1mInyDFfBhHQvlCF2/UaIRmvao7S5boZyjEahrU4zlCubv3URPE/kcrclvq0VbAa
iRfZcz92+ghM7h4ib689h9o5hA/6CcHL722B/x6cOeOL22o1HNVkqva6afJYNo7F
pirAYfYc05xuXwbxFcwNF/uyhS5+673MFcRKhIJtYZfBMA8XDBvEdzbLxKYHAkf8
D+DClmYI8XMNrNEFjgCoKBol8qVrEryha0G5WCpmrWyWOf1T3d64O2tQosVf0NfH
Zp+DB9+0w7MEENhpq/a9aR3orYYXrcYyfAw3jmlyhsAGVor+tZW4PcWQIB3nZXp6
esNMR3xcs2U87ndeIN5T4vPLJvdAfLORF+TjUa+SRY1/Lc4GVWbgOsjMUuZ5V2dA
CmbDXWqJf4gwq4sCJ+xRqoFqnO4lm3UVknj9X5zrsthuoXN35+eSjUGGwpBY2QYb
n3cHc0p51ORSYKf23TO82Onl0BMXTUz0wnWIPcwDlpZdaOugcHh/Ciz8PvEyW9KO
2P1YXRKPSUeTyyyYSCQsaaQp3MWcDi8H/sGMtDY/Ml/vCHMgrkGSUiHwwGMzFxqL
1eeLWA4rye1s8Qy6IyLxmGoci9U1eCX4NvTsIr4v8pTdJn7c1hIfeJhj3hflyOfC
GBXq550HNWyvR7Yzouo4Rpi5I2i6CYUKMzEYvbIrqhR7hA4vn9YHkk3WNYvZkKze
q12jAVksfzNDdZUwG1yJmNGfPguwQa7suTrhaLiYqrvNj4Wv0pSPiVtdoosKvpwm
6kW/Nfzjvh+pAH5hukxdoloR3iIirjsQZ3rrKOfjoA1NnZ9HwUIuTLmw3RrM44Dj
w5nVr0KQJbjqB3LoMXZw8upaN0tDJqzV8F8bincyRlASHQ2cTeoxqyQGkOJDxhcj
4iqQ8trPtvG+qune6kiYzAn5NW4IZKgyHCS1+46fIRtQswzMk8UERUOLV/EAeY3k
EiTELhZyG/Kb+tknD1DEDSa+OTg5g3acGinl9a2qt63BOUIh70WApmLHrUMYxYCq
ZCWatv6UUgogr9kSU78NFWUiOx5hzEzYrRIei9Sm59iD37I+4eaADideUpfo47bD
unl7TpxKel67g/leleT8QiUE47IzCdA5NuOxhoTRt+Nc8DUbXwkRi2kP7ZmjaWpV
tXgKH7FCFyYbmDJmfjxnJ+o+Fi+vy2e9h2ianS9dYG7z6uiGcvVgaYhGvfHbBuUg
iYxaJsq/5EdvZts+1NeGzzyZt7D/em1LffoE7fCp2OOiinoNrJ32zOryky7CcPdW
15dADkEDApm4yFMko67tTeXpVh8KdDLs+PtU7r2MfS/AULQR40nJl0rbsqQdpz0A
ztgbKT0v5sZkH1hxuHAGZwsQvkDkRVcB27KLdQwuWDW9OwSvMLzcsn3mQuKSGWrv
NN8SCuBtfPNU7uNCJy9X17gw/w8tbrf+gnjxSSQSwCzEzkiu5AdlrQHvCB2AWsO2
IbIjPOt9aKaFRyZauUO+qmCnLE8jl5QJRyAPRd59BeARC0jTn7ziRnr+60iWXlue
1Dt9gmAo0eAtUJt7G7oM3jz3EvX+9NshErTV9BjKRsatdVKLIMKvHzDzGLDOnbTg
vb2NBa2KLqZbWKEj50GcgCH7RHun/GHn4cpBVlMsp8+LX+a1x5CPifIMsc1Qx/e6
lX0gizUHuZceGtU39eBOci0S6oS7dDxLT6HmlKxrwmJG+8Aq4whQ8FGimLqQ96Vb
jNfvVjTSnpD8gJL1Sq/sVfC0/8Cl6vA0Os9dGB2oqXep8nTjoIBiGSiWxuDwK0lz
Fwn2Fgb6Y4XgZhrs2BMsYVbguf4XhuTigb030GFlif+uwwuFZEDj7xnHOpP5zkdf
Mzdo4RDyGFtrNC2vwcCGrk/O7auStAGk9y1ueSFXREuoTR+L0vkhjaW0fKc8J+Xv
6NL4cIFy1FJx6mYOdXIUd7AjxXIlqEEK0AkObklYBHYQy3+so18dYHk+yMQR33rL
FgiVEb/A9HXuD5JxBvDXJe7gV/qyBVMZhHgJmJeko+ece146NgtbQpUw24tJ8fCe
gtCogz57vMKwa/EhobcV6kUxVhVU1tyZuW72klrdlv+WR72npjjhStz3wqemEn1i
q3iqg9lomINBOeMHQvaP/0V4vETW9jw5i1/P1Ry9m5YrE42ccXR5/9clD12QVo81
setdfoVgeF53MH9g484Xnk72tdl1kA/bhASPPNP2GUvirlNEbE0WOHiEcFcIg830
cgqI8WGWqykS5SJ4CrMuQtdti2L23Xfh/3FbRdLw8c+nmejuxP0MaHIxpp5D0pvg
QAhAv3ag09i4KX6iHim8D2PlE4in9NNA1JxRNKSiMO+2fgaR7iaYCyPqP5qvgAQo
ahFyR1R0PMqAwAcwb0rP97s3KYgLY3/6CzmnU2G5F+tBlIxsJiYnAKNFbAYJ+tYI
MwydfTVXaWUjYe6rqePKSbF+sCWIbRe1afC5sys5c7CSkRLMtv7qnm+q5JZLCZm4
Ha3GbkMkahqIxemoxCyvFkSfGsvNKE0FK9fD0jg8DKtzC+QUXp7sk0h8EbFOx+FI
Zz03GBhMTuOs1OPn8OmUKMDYUAIEw2s+Tt+rcQcIa1HITuyVYWXl6vlzi/AlwNhL
a0sKcQSauZ/b3IeHPS8j6/vXXiMgzs3A73jP+QyPqWnDcdpmLdSqDR+IFN+wQtm2
m5wlGEKN1oNNmBLFuVgAMEKlSMoYbDYVIi6ky/S4/LnyhRLYMO82FWXGu265kUDX
Gsjvm+8tbZzW91wJzMj7gYB37+PUl/ouceEo7EbektEbkDvOyWkMOao7kbzg+m+e
4hthm5dWviSZ67KSOGwQCK1a+7NaFDjF646sTE0rrBt9A+YQBszuI6op6zKevtu9
KLCeNRLsNUBrPPDOFSNyTp0C7dF/+rBybRhlznGX+39rXKrtrbVh7m8wCLpO4ri5
j3D8N18+OSAtFDFK+dWazg==
`protect END_PROTECTED
