`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LHgsfESpLrQ32UquwphxSg+GdYQ9+cFM96mMFm4TnjSpkow0rPVKNM1QxaK0SEiX
fkonYfojyPTeyJMnjMgvMxuDBxizbYo1j58S9un2tTYMubOVfz/Fch/IUMZcadXk
wFc+1pZQaMaUEkA4IyUy3gZFkM1AivJbgeps4t/L6Z5FvN79wEueCuZcELczGRuM
T2O5GE4aGF8uz+n+EnBfz+l9aMaq5XU1T1LGr2oAFJtu6PwZUiVIpz0v4NQS/HSx
wAp+QrmDf913I6FPjbHW5SdqrBO++hwKvNhvFUHSrULsBvtbL/p8OZFrvKeMbnnP
dGfKycrFYxIJoLG8TBoosKNMwetm9LKv34LRZ7i8SrihkOWNct79aebkSo2PylIB
DL2gwuw8U9VSIrLwCiRdIiWs3YNoon/C9rbILdV558TrLpLVCe96PVah28M7Xscu
VJRm/zVNxlB5KNdHJdkcVUDh8FIjXeW+5XSSfT2LZ6HqgSlNuQNvxRyNWvGdFppv
8aqJhPWfA4mCnLFVeZHmh/TbrwpuKacERnLU22mDjlGJmeNOJYQS+T/5lFcdNBiA
2D2Nf3y3cl0ZRP+j5XKmlBrcAixBbhZKmgCbnv7IkI/8piXH7KaYJqDTIxoxBp84
GTcAag6C4V70pTsOpMWNeH/7ubmCoqUtBB0JS4tgVzPHNbjJ+MCzD2HRDVabRky2
J/20AstJ157ZiHhUs/CYSl87n6rrRshSV5hhuXECULb/y6Xyjm2uWFZJOkxLy52C
clypCEPRl4bA7t2yTH61LyWTk6oHR5aGRXPmfUK+14y2A+RBePJBJq560rbpPQKo
fvwStqE34ENXriqOHkII2N+yNagT/HvAQsJGIuUv4XEdK0tJaVCEYyi09B8ZTdv9
zsvPjnusSALgr4IWPF3Tmaqc22seN9TUPs6rlRJ+Wfvq/mnkJvAU8fdUe8xEoPRa
`protect END_PROTECTED
