`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cw2wJ8BqRlWmZ6R3+kph5BCJk5YFRyIXzyOZv/TKGZSCrnjuRKVN91TNpmXSAGCT
Gf13DPL/Aofc0BHvexPfB5U2XsOrcegUK4WFrYeTQ3AymS9MKo/MHIXFo0O7i8aN
qGY8CiFOvi9KC7dLXRmXsxhGDzJw7Z3ldb9PE9C23+Z1IiPUZw36F/ycC6Gfjao0
MEmHD6r6HHkAfdalCuwHjPuYTns972mp4U7q6LAl+FOeT7m2GV1f2YDTqcLHwVuu
1QCMoa1j/HsQX0Qmo1gdFR5mDB1XvC8Kj177R3Tc915VopC676FLJOF5ei8U6hk3
1O5VxK5LigF5a8610ZBH5eDs08yeFwYka8VJbpEAHYmgfc6UwcVk/oqmnzMvVmvp
WzDHVdOoGdy10856IyWwwyW4b0rRf7JNHe/q2bJ/mblwUbcGnS4MgbwV9pWvxfyp
pt4LcE5AvJoUH3I9kYrEt9HmTbtKK/Sh3R1ccummogZQFYBxfILYwZfVydyXoxpg
VbRujcGurcnq17kc6BKE9HRkav6Js59hfGvDnS+8W/iCHtGNKRf+1r8SKFHrGVQZ
wjD9Q5LHceIqQH8/oKe0EsB+kXI7mEVE1G21x/Iho9RmvOODcaJYKpqeQh6ReIeU
r7VsI2D0YqRi6pL6i84cYOpKgLDqqG6czD0Ab+sRwHWTbKCKknHUTn8HIiPLHn69
dMMDZU3fVar7ark1OVz1kdASrjQgVBj3LcE5wRF8G6q6sxF2EnzTqbbmuBIC0+FQ
BCb0eVxXqCwp1Y//aw6vg3r087QIh+LeepDgXKlVHJy+k2hS7bFFpPKEQPgqC5sQ
liFsGO9FH6u2d7uZQfa4UB7S35hQjwPwrvozI/s7v9dzfF7dbf2UT8C27cvaTgky
u7u7GT4/X+UMQhteW+J1f5cu5CZ9DOlu4lYW3xGwEfdTHd904ZhuNZjSyS0cmafv
im8QrG5iUfOiijxQJ5PXyr7y2HgK7XXnsvVGL/gAJ5koWCZldM1cLxBGNGVjmvQQ
1k0lq0oH0fojTgYqtQbK9p7/a54AW6XgMmY/kT4fH0BKxVv26ZSdyo52pYokzq64
k/B8rMRt+XPOK/mh0dFVFOjvCeYhBoOOAYyagOGcFTXHVskEBmzjzlIE3k+2ndtd
ImpFw/AhcMTOP43Z8zddlvClpepZREatFSIexoGIpCKNtwwF2oexNT7Gcoea9FUZ
YIPTbWXyF8gfNBRkfzUC+1D/tZCqcnZ/zOGqkk5uCaxMylWg6ld1qoua65xz87w9
9fAHbTmvRdX4bQ6k1jN9CrO2cPdT8DugJ7t8ERBtrCXj5twoAzgQGNjhOr5wyeZR
Fz59tFWlXi5ySO7Avlm2vcUUBTsjJVaVjRMd7DVT41HyPdNLEPWHDMeT6n8heC91
4OiAjxNXXcOCPfeh/WVAVrQ9g6rNWHxN/HuShYxnpdJPNmNhgmmAhvVWc68Ln82+
B0CN8rj7ZXiOQ0PlcTHBBMKmEaQXyfx9GCRU3DiB7xY/63zvO8zEchl+G5X1UX1r
F6FA7VyOq2Mn2vCiRsHOqWrecKqreplHNVbpIOivXlFXjvm3XgbrkxZNOXGwxeG6
b8B75cUyNTVwLtjT5Yo5ooeBNKa6aKr0oqeQdrV9midRErIu2IUZ1pNNXD9SLJTT
OGdOchN5ujm66SfI1/aZ+rrzUUAy2N7QUelQMzTuyI6imzkg1cESloOAEXBin8ga
elh4OZxEGSOvywLqUhrMaHZv0+/XXCmyP3VOInZN0Hkqn5bxjGzm5tmDo74kQgHJ
pg0jLyHzrfy8+SRVN88LDYvu7vBHX12poI3j8Smic9/Tyj7ZX0F3oCSzy9cJT252
/IJuIFgLPU/toLaAskLsweB7Vcn9+cVPyO++1SPdT8eqKdTHGdgJACRMhSEcX5fK
lIIvC+MJKRfQ/1/iOlPXW/jvvl7ZBIdoJdpdORiIEzZpdJ0ri0WJeT4kMLh55rba
Iu5YYsT3dQKF5Tnk7K5Zf/7TF62ulu7qhfU6LujWVICCWNBMUUC5+k13ZEgzIc3N
gDKlUOIWEHk4SYjgg4uEvNCxV6kHxTAeprFXALnkrYf479BnJC01bLJDq9r4Q1O6
MGxXyhQB8E291lWe6JpsZYgfKqv2orTwPVd5oiJKAUXegIqDXRpo9cp1+x0UkYv3
WOdSGg8Jj0YQNt04pVKVXk4sKFCjNMJQVGIzhIrkuWf0Ubzp2suQ7G5XDkarhUXS
i+0io+2SiZXGK8w07NFmlO0BZPmzIIr8OOETd4Ah7ij2qGiOMpEWxWZskEWR4MWC
F3eTykpbOI+ftLHhsqt8zyB+bQzK1G0tlq931cyb4qdGhZJjnort7xO/n6ByThuo
cWv7ay7MpKm/4LxN5c22WhEflx5wMhrfXoGa1DvHNXSfZnV9b9GSV8otxDebYI79
7tPg2UN3MnOWPyQUpU4W/ElZgR1yQBrseVXvHhzBDz1KXbBKF5DWgFdVroqBgi0O
z9w266iSLbbN1wuigHI5KFvu4fSW40c9hYuYDra4SjFf7DXC9Fx+A9IECkbeIpRP
pMAr29+ppKSLCUyFL2thPw0fDVQXmEKsvHrjvFW9KzBvmBshFkSCb/MNlnzk4Odg
KTF3TvuztwVZpey7K4CTu/FMXu/wYeDoLDnY4S63De48UVtkoXw22TaWr5JptIPF
L9tqo1c3g+wDOuFQBxvfJt8FwLlx25n1Mfcor1+9O0FiqrCG1Yysk40nPZf3ASoc
Q7IWjxin8jvisZ+uFSG54RGhEJTrzuwk77s5kK2DaeLBs6+WV93/I9IHKr5lWSlm
fMWinQlsmJzBdr1N/AbhSpY7qMVQnv2AWlF5mMLHJU5R3Gb2VgLE2iJx2WUhStdw
bnWrnQ0P3cR9cnlqpcCY9qNPKZ/Sy4wb4w++DT9bmq5PkoE/AW2Kq0UPwpn9hb+d
LrERIbo4MiV9jkZmYasuVWn3TKuzLxVLYV4KN+6+KUW/xAuXnv03GFkBp9EMldLc
52i46iz/t/SNByg/98IgvXMsTUVGzTewbdFJwMnft20h2tdS/mGDKbK/ya+29vSA
zqqyA7EWgZXvUvIZWUKwpNfhuwEh4TrtZuHxXQin5lFa7mwWGlQ3S2xxAmrYjbGI
edRN1PDS2YKfe+d1Iyc8N+4wv7IzEgkGAbUvB5xx0QWJae1lHsl/H8w2KmDV1f/k
HoaoUJN8GhXFxPNF5P2ds/JXTp0ZkXk9uUKIgSipBD4QlwFbfdRmre5tyx2NMpo9
mKq1Qe7enHQceXRU1XqH/fqlgSyXH8ZJQ2usQ72u3uMX6FbkFcRv+ke6kmoVlhAR
8wtPwZP3JJupK6nV5/cXgW5YBnwNDpaNdM6IcZPNZu4qZSxttBmDtvWh9z1BoLUg
t7dtZ68WYm5aoFjNAGV8K/WnwKjEDePAhpVSfkEThrYjMxk5ESJKbkAFWNlIcbnR
DhLF8CIq75Sb18kFJsWwivqDLlsRpYhJdZU9OjWUsPDx6VYqacCR4SPJzQtfcV2H
JhYidSl+LH6JOWm7hcil41U4Hsb4O0bEu7amUwlD2aJWGUKbyX1zVhTC2YY0mi3j
hLSQV+sWNdB3VPehm7EofD4Cgga3Wx62ZP3kNJwvk+Ts8nvCCM9IMfIOTVr456PV
E1EHLYXatYEgzsWKRfqPnUF0iRg80XpUVIK+G3niZIZDRUG/ylFx6yz7B9arR1Ih
C+A88KKKRuosxaIXY5AWeRHNoYHUgXUW/eTrBjZEuSZlzQihLW2lmNXANL5LkZVp
cirak6akVmS9ifoE9f9dsJCPSXraRSmlv85JOVFs+1zx/EjkOa2tm8AG/XGxZOPn
GIOcZcya5pi9n1yQW9dV2X5KxIgjoL4grAewOMN27rGcvvC9AOtb5CPoomINH3KP
HgQfLOuJvw0z5g5u0UlFBxafdFYjmld1QZelOSYx7oZZUUX25XjchVaO95rC6jdv
6NTjQl/JRIcUGY5aZJCerl9DG11KOSjEH1WgI2f2gChQsQuBo/g57CioQlCGnjVx
f/hmv3vgjG3PBB0NnvlXm6tA6QLxMyZf6eNiirv+N7j8efNzmnFWiZhTKEu6+yYt
Jv4WyS/KhHMaru7Hs6LhTD9HWaiAAz7Jkqh0VsBaWAUDgplxHu7yj72PLxoUNL8d
pO9Y4oRMX7IXIW4EYNsui716XXCiFdkG5OD4HFS1GiD818jjGRh2o9Dgs7TA3B6E
FRB/kLDRuyRbFQjtiv0OB+HHRhBTB7FlJD0/bUPlrYnNcGCP+1OSFHgnu/4O3uCJ
5hjY0AyfoucDLxEdhVU86nKEptS1VtiGwCuyb+lMt40mocqHVkR8D+6IVD08OHWv
82HC72e//q12ZwSO13cFEn5TlVr/BcVQv3y3ESEqE/ylre+IuzYY41u73RRLXLsB
1zqua6uAXwjyLVVLuPS2evljBfiWBERLCcNFnjd12QPJTvOeRlaPgcppaBhRxcFP
Ac3228SkRt0wJ1gjocWNl5olNgXJiVb/ynMwxYD3DB3WmB+KvLfLlFKn8fTZ9vr1
cTDWODRsmEYizkz0QKAu+7Si9UGNdoJv5G/MNBCEgfyRYjt9k9Ypjycd9RJe1khv
SZSsFR/pb6njK4RRAAx6KvLKH40X78jmrwds1l2GEv6y2rMWP5RuNo8C2i9v5Kik
NnqN49587NzOfp4m2VBJsfLKU4lGXWB06XMSVey3W5bQ0D7topX1lFtwNqFQbQQq
gA8IFExO0xPmS1U+peuiJh21PAxSei/3oy9Hy9VrsbeuHuwT/uRh5socCZvehnfD
KOwUm4u+vPzEDfdxgl0jqIZCXf9vWHGmVXrX5duMlOCrcyFI/0tdWYthQxq/2B5K
Gs8t2PXVnAxiBl8leeStXv+ZzXPd1PHLqL/KADPSoPVuSqwS3WdqIQgFT4M1E+LY
teLV7mLX+BTT2PQLxXsVdhuSlDJYMxD3iTAD9xjVCBb6BRLRot2aQTjewgqFkQAj
bwIOMiVK986pzvenUQ32e7DKdBqwO++H8Fyk7CeJ0QgDWmHfNq6On4FVzVg0sAxp
l3jCi0UxCAITPoQjtiSkFEX7ecHgJIrudu4Jdi893eeuyeu15bzrDwL/QVb9gYfd
OOVtiGzKUKdmMxxIglHc6o/gel6LW0TJwuN77NvKvnHkYkr8kkXMUqlduyvzzzhD
/fT1dzvsT+AeuZAiKkZuHcL239zZRpo8zSGTUbelieGhE6511jhohTxlfyhgmFun
flLO59/fJtwA02qlMjCL/UuLkBcl82xHJj4Qj0kNhBz+NfSY2Z00QflNjViK3/fy
NWPmiBzOQ4bGmCCw/noRo4dchGdOOx9EdSOaLu3PbGsQDxTKfZbZrTpHJsOHI0EL
gIjECxDae6Jys8B/LGlu9OG/xhqzQpjinOqz8fTCqYWCoKtzjscw68EISDG59qkQ
DVH7I6YkgfwvrQmxpf8jbmxlJV/PTRCn9oQCHR4DHsf12y/yi6jt/OIPPmItFMU2
twndhKaSE5JExzGRVyIQqtAhODPQ65JcCG0gxslLSgHePCihAB1EnNFU8nkuq5/8
oVK3Zn335kZfiGBJpg+FxggQICo8bg5lN+/XV/JuKw4dMpxLIy/TXawMUEFvm843
OR050BXTFiV5GjrlvoDACGil7k9aMsoqyFV8vChiyLWSnQHfMX/Msn3qOlAJnpLG
HFG6g+jq/83NkoW6LlxH5TvJksPjdQaw9zd+zGGHjAXmYCfSih5LFakmuQjtNEam
PMFPBe0trRZ80XW9TUNFhyEp4dcneJp0HjIKSplEWkaGeD6Ue9cbxw82VoBqpiRv
O3uMTkb3a6kjbE0em3ZMQumVp2Bw1XpqguF4rNooDjKWcyJRHdtHqOiUSd9NQT65
0b222fU/AEvbUZ12S3w9//krJzM7B5qQPBE1XQUC0j/pwPp8paC98XSrcsM6+jzh
3XCymQvDIVG90TV3BaZXqG05CXRdZ9J1l5ZZlQY6A6NnH3VzoE1I6cCbS1Kzx2J8
RluTePWyJTIvFZs2VUYPeNa4Uu6P1pTiJXt/JrXEQrh5H7JdUJH9xMwLqdRU3faC
KEuTTp86Q9HcWl+cXpaZHMTESVi1N6dPyhQ+VCQWGAQTsEPXGdiXOAUSuerMxuqd
DIdgM+A05DuyISCybUllZ0bkNRgQngUc0fIKyx88LJMxmDLwbIOUtPL0McqLW3lj
C8pHSG21sLtgA0Xq/RLLQh1MRaOIK+wylQR9NO6IjoAi0vFjhp29BuheEfm4koLO
tUlhz9tYX9/IeXojZSclEx9uT7Sn17TNIL+8ER/K6ZFLT4sIeoBQFiIxj2WnSBRU
/9m1+wJJNpquc3WlEXxynjMaSIYaVMieWGjl6RferHrzhMKylQwHmWNxqbFSJVLB
3ME8/kjI5yQzkaB7oIV2wC58ApmL5dc14L93ikAKqS8V5m5XmvYx4NTmbIb/hsYz
lgPX7LRFvB5t0zh3Ip2TG3tr1rgCuJ3LWZbD09WoiIRIEu8Jdu69lCxfFAqCGfdc
NOxnqhKemepqobdjm7pi1Y0e8j+1rqCE46ivBTqfeB53ctDvBs1HKq/NbxcGQPGo
53ev5lYqCVrmXCX/AHRDJwFYXognEa9B8wev+HwU0rkHLpyJ57rg5gho5PU9aArL
s70EWpSMNRTsvzxC5m9p+st6G44NwBsxE0JPT2NOXw55d0D6ayGIo9ZVEc3DX8pp
ae6RbFnYr81Xm06hzd3slJC3YL9lpKRBmhdzhXC0yZelkMu1lXkYe4Wif3Uv+4Mk
QFiid/OcI6TR/M5ZEBbqyxlU6aVsqg6Gzr5xoZF4b3knImZHuEUQ0IznH2bmsu/w
sHBCZGb/U/WNwKxsG5G7m4whE1YYvpgHRNj7S5f6I/lkxuPDpCluXS5dAZZt+3/9
nx31SKV3l3KfP5tm0Ywl94MIMxX//HTIScV5Myu7HwjDkzXm4Pc1rK+XaCwZq9Hf
`protect END_PROTECTED
