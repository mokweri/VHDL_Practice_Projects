`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ffz9D5wCq6g5+h5t7z1dfCJEN0klcqa42mExT6fjpd73jVJ+472x2HEuhUxY0BRF
tvQzfthbU7ixXAIY2xlQzakhuHk0+ZujCd6c0zqNlENxE2h90uI07BXUhy8sxDkH
dvrR6cPrqOt0TRrAJTlN4kelbnqenKCNj1psRMMbDUq7r3T/eNNK+V+pl8XmM8Wj
54DCjGvK2ESAG0a99WrJe3rogTnC7wRvEeEhJcSXGD6h5H4IbRrrw1wy1bBGMmEw
e04sC++lH5sMcK5OArvVRVTcoVAFfm8KNgCLJke2TlOmbw/kvNhVl+JaYaRXTeHp
VkmJAQJvuxp/WrU/b5/W2sRPObd3/mYnSMHO8U6/vS8PY+5rN7uSW/zplhK8Sc3a
48PHDRtfdfDF166vJVtNpsyvZugjI5NcTAEpFs2ff7DBtrizNeIuZptGgiq298zl
4I6xrtK2hk5K/1P83yUrrre2RuLjeN1WDsAIveHDYqEQP6hINxzW+trjzrwU6bno
zZDnVLzocrKhGrTHr+gXhxft7p3yPhJFRC/CwgExi6+O3iEYH7WVYEY07Llobrm2
uqm3SVr22u5LlN+R3IdBbScmg7yceD+k+wsYu6f0okAbNpM8IgzNeOSM0CBMSnvI
c8nPavzDjIQycLp3kHV0XVo0tjy5jlu9fWISq5UisNcVne0Iyf3xPq4CoauWc9cj
5oXQQyDIDA6vtCUDYHHPrVve2A5MMry4ywwdhZHMsR4wx4ihzShOr3NOy8BC229V
bw/k3bY59FUBf1RzM7aJVwVVHYCS6zFN14CMzA5NZZ1X1TxhfjiSxSnujHVbpimw
Kf+WMI0tQ6RrydDDvAy6RwrLEhhiW0yzACx+QWxwQd4G8fuSmTkxzMKd/2wSb1al
1omzeca72lHpl0PgyB9oiPFexO8WxisiZoiNJ/Ak4OzA+8vtwFpspRUbp4/WY04p
4Y1UhEmtWbzpmpI8xJLmW8N9iJFQqIm7059yMp0JtnAHFqy8qusvHWLb28YfUx/n
Ar+DkW94HPmzfBHFkdmE0jgG3by6BZBDq0uHd/AbA7hfoQmkUvgFnxS2WII+0ycp
EZu7FBybJxgKQ48YOTjhmxQWdCz00vl+aa8lGJT+6LzygK4wafVt85vZd4EX83vJ
zRgejgvr8IEUuvdzBMxokbuHF5LZRaglW8YmOj6VzuzVW+pQewSNLBiUbMPpohxf
iVWZYLN5TwKpR+8tD0hXrLyRPLeKsnNx59L10A4nfBZJivUXwNnU0r9RLH3l2iNW
iDE/sZG7r29Zti3PHcAkypNwDQqMa3Zw/CRD3X15IORXtyNqKYqvFzhBnH4YI9R+
h/STnp0awi8ATSpbaePoZ3M13KPpAkQEd+Fix6xWN5BTgzEpUcEt7CNfL+2EZAoc
I5uC+7L1ovc+Phn4l2v5kefK3S8F3f+YvT+qT9Kx9wUdvWd4Cu1mEWwRxKRDjzCb
ZoREICb/SEFD2cAoikeKUCAjPYsQafbSfFnYh4gvcQPpYRCiKTrBAhhR6tFYy6YZ
g3oCXkcC2qgbv6N7iS6yI2f+QCAyNZDvnbR4ytVqUlowsR2r0YJBSY49N1/Lipv1
HdGgL2b5Ka3dvcrwcQCdd4qxyaTNbK1PDoGS5JuGn91jC3VIbX//O0n+PpK6S/fU
/pbA/gdLOcQQQ9271IoaHMYrfTvBmcapNDcsSjZJCxtqCYtNohW6n0eaQT9ETLEu
U3S7mv/Qv/owN3mr7zpy+hm7+S9O7VnuxkjHdStlJAbG+iNBMzchH424ITqXmbJ9
7uH1pWwpzPw4iQfFl4OPMx6lx2X33jhTWtOJM1bDPtMOZBNzn2roc6Kjm1FqCTva
9L7PAi5Cz/xuHfR7UqamJPQgko1FNBDd0aNrfyCmVikptE1qAh5ykEpqOEvqK4TF
X7+fS1U/uc9rcGv1iXhh/zHKbMilk7H3gHU+6KhSj0+FA/z8iKY2soJcCTP2V6Bp
1+RfwCOudz5jLV59/JsQwNKa3a8COQNR7go6ipve8NHHYnenb1SgPY2XWjpPkfcp
QpQ53S0Xui8dT2UGEO6LQNcmWreqniQWs2fgHq1iQONzr2bB+vxC94r/J6B5YAFy
G3XtjNKXPYYCL92dmGo906hfPI2OFcXqQ8ynq36U/8qPH0Jb3Fssxg2yaiVMQM6P
ZRXK1e4cka3Mha6bM8DKjjdV5pmc9ud6gEi4mHOwQaOMNa4bqgrfjoKoGDl/rwT6
y+7wSGRJvbe1u10Ot8uj9AEBpo4MG5t79SsltZDubBDyZGsylJu1L2sGIEuG833o
Z4XB1PfcUNZJqriKCLMeeM3Wrr/TtO4TM/tJybiGPp4E8FNQjZED2MS8f7wg2TbG
xz1Ca9IHR5G2Ewj3rwNaePj4jonmzi7rvwiYgGjC/9XVzTvD45kvchWFIdMRIdkt
`protect END_PROTECTED
