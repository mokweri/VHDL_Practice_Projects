`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RP1ketkw+QMwPpLcP2XDxIosg7ljK7o8J7qP/3bi6MBuqwLcsfgLSjsj5FKaeIvZ
r1425gQb9c2qtIDzktVwwEjbMvIvDn9XHHTSAkZtOslPq7sR8+4tJMzzF3XPpNz4
UIm9fqV+iLNVE+oxVgifTYecbcw8+UKdwyJPuhi+ppyXJ0xNfQ6vET+d8O42CB+C
5mFqTHXkmb/kVav5IPXXoJWE1cfZCLbXsK+jtJwGl8iLNupCxrzPHy8aQCPJNoSk
jqru8NMipXDGgEwNTsN363TSXxEokBoeUnlIb7bXU3CD1+rRxJPvhsePcMr8XxlX
ZBqBWfsNSVBhV71sLLibXpcmepGzKknLeXJKDvammr8zCep7K/q98zLIuOZPzj4u
BmUkDzu/IbvgyaGF7nhAyYKjnJe1Ol0TVQcEZ4tekIHZMOCEw2ytPq/B9qZ40TFg
W23KbfEpxJ6u5fBkMZLhoDiKEdBp+FTwiVb9tr1wvSyT7x43oQ7iRE+2wISJgIPb
suYkPo58bpzQqQlKayqSsqgaL+jxb4+w7H/siQTEK6VRRi4U448m97Go1l2R9b1t
4OI9HuG06Wci2LWfgIdToeu3HSKxSNyB+aEeTTCG0wsq9VdGh0H+QTU2rBpaIYL9
8IDzM1hv6hCvuHK22sfjAGOS3DB5RcX46rpifr9HmKy7E+btfe9Bxq1ooGWXFgLk
L9cYNg+/RaI0UCCrhrhEjDVF1yQBwptT7RFGpFKZCMPeoVzv6nY3B9jaOPHGfOL6
Vebxz8Kc95WVluUYtz6tf6UDkdpkrw7uh4P2gTq/1doUMEihGYYlD0k5DJKGsQfy
zmC3nYI4IwWaKeG1/3ebQ21OM/t53kWbVn5JbLP/glq+sCuLuDzJ1bVhquI8IiSc
KDeD70GnFHBv88xY+5Xmu/nnT5hlNIKWsMZ6Ai2eKRtfiG0OkU4PqGvwoKzLve8b
eVZGONydz6QKxJ+no3dk2vS1/T7HHkXMh64nxd6ZDqrcpRD5G5lCSEbk0A8VADnU
DMnr/YKY4aG9CGU5G6dQbjWuMzdGPzd+S4+Zn26LrzuilULBWuLW0LQTQbnIwYV3
/809Kcc8n4iRENxLDMwHoECDE4wPvjqiSazauMauKzT2TGGTChF1t9Ozsa9EiR79
8xPygixwAsyap0MvbyaKrtt0ZZiwzVxokOhCpenDiJSgtgEWFie6wbT17AnyUHjr
k1gbZc1rZWOLzajXEnRZ3oLZfPqsKwd24FkjxumPtDU=
`protect END_PROTECTED
