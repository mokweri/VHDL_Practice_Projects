`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hvIl3DAw52I7k0Zklg9WtJaUUmJ1dyrAVFms9RovH2OTGITPdGefSKNu11CPL6Sb
CcNVjVyTbiGMrUqU+wAYaJwQmvb8qkHvQ2hhmzZbtE5mzRDV2Rog7Uy3Z/XO/UJ7
EySMT8G5i47PcQVSxDX6UrH7gxwnbNrr/c02XXArPg6WEORu6yOwvMVy4Xdq41p7
pdpuXGBDP6CrMJMzPNbTLvCxS7O6VVZE5kDoXwGMgNTIr/BJ1LREK5iCMqwOnAue
al8aHloS5nBNO7cLPxpyVVBKBiuUJOSgBvvyNuJZCNg+jfTzXMwF11VT6b6gq4uq
X9ucPsTe3nsLxUU6BbcZ3HxDhoVH5moPnnNHWB2WvowBxaHEG3wuhvE34YIa7aPJ
krp7QlBMb7TY9Jenvkcj5KNTeqWpCytu9JGMl0XFNE8iGZVwiC/O6ENSlUsP+fCc
wmokIXKMBCZVwTotQAa82V6xGGV/hWy/3bK/vwMRNL1sFP3HGj3d+DSvhr3O7DGy
BLc0LABF63tvNrEBUo8OHUHtrbcpyDbkMS2hb/wCFWusJR5hUK2RGpOA/tbMqk8H
ch1zBGUOgyd7SILrgiqvTPdbEeoMzcbM4H3NwDevMVcT7CEwa8FYp7RaiMOXKsWn
2meBQUHuqKYJuwwzPlDzi1PTO/8OkEpss3mENtRWasNaQtTHt3AkzoszyEtPfkJu
O5OHJtNMJJicVSdt+Qxe16XRSdvEBmG5uydmEmfIllbIEIkYuYxA/OV0uQk4U4wR
uPEYUjcwR2nK8ZrdYNPc5BwocQZXdJ8+x+Yp5MgLWCj5JJR9CKtx93fH49JV4j2b
S+9hEVTuEAlu+unDx3bfYsrF10wfbPO9OAnz/zBRV3zMCcYW1z90OyMP8VPmghLd
JP/VvWDIy5eoC7eHthHZKh32EGhPUCy6L1+vnMEtaoSjThZCae4ZnwctkFyB+9MA
kHkSbwrqzjWSf2BJCt+q1Z1ytM8K3TIuF0s2r2fY/6C3h351PXrz/xldplstabDt
0OfagH7pO4wE1XD8rOE1zyRzw/VSDlcJUVpi9KLpH973QYrhKBdO2BoKsDfBM6bn
bOQwGDlmOe+PlnoirgWRKSKzoUFG4sxfdSEZgHX9M1KQkyMxm5b3Xlq9IXfVz3Qy
usAYN4Ziyl5vzxP3vLc6xdCXyLw0zBAlrCmVSZRQ0nUD/FSo65dNN3i57gHumByO
pCnzUfuIyCgq7UFMxiHN78DnN3MvDlevhYAXnPFjJaGMm8qbiEJFp/HDNERJ2cL8
Ea15isLQ4w69+oBzI2CrkjIOQqWPB/jc7KJz077tyXOwSasSlgvkekzx2s8as2ic
0zXZP98CRiPYS549BLFm4mnvwZ0z0Y99TVzDhskyzLcgjFLatRJkqUV66gtIbjFW
+H88gQZ705kwVkQfyUC5cXa0dErzNEn1uv21EbSV74N+QY03vB/NAkei7j89wUFj
6ccAqiNEVWaBv9zXTmS656G01ac1uxbdwN+k7qY8XZe6cVwCecyQSYVxfR6rf9qU
NvRizI731BPc/wOuhJYQutDKcE5pKoums7RN0TXluss2TIBNPbS8uJ53IdyiB6W+
P5CenrmFzEl/Yfok/v2k90O27bhupoyticYI8Br4dKZbvE1J/QWEy9HN+057Cihr
VZaiGWsuUBqV87Go02efAc25+o0rNDdNEkXSEGDhVyFIqmkUfylil+diqZfT5fTF
WjkuKx8Qv9i5WTjORG/K+hE6giFE7wCu5TsAYMIyfn0vHp5T3xfgpWNnbUtFqyoi
eEnvHwizNxECQhaaRC/OgxgnJJ1Ar121DVa8Q5JV07Mfu8eQ1jy+a3AwW2S/+QTH
tbKrMASrQREbZMR1pXS+cPKQrKVya/740v8M2HCIz7ebNTbxbV79CT8qw7whWqQ6
3RxzLQsDq5hOHr0O5rl+QxXxnklsD40/WZ89veR8YS8SRj9blRak33sjaDEAUaVU
QWGZAUBPrCEl/Ajq4zdYDgFFRIj8UerQ69hm8/02yELaMIczqPJLv0O4ENxPdnQs
2oXa21KYDPBQ9ntgRITJ4d3B2p8MEz7+wt9b1/JT1bwJT+KQsDMVKgxcQdmsOSPE
1tf8LgAcZO/gkN5PvZrQHIyUi8CoeczPQD+iN5ZgsvnhxRXryywnMSzkyqESDmsU
PDDuYDNpEVbPRwaNqQD2V10M6N59eQteQaIJtBk26CpVOTQ0DbSZWaIZpcsCyOlY
tqJ6ZONkZtQ7ka9EgXictRIVBb/aaltI9An9I33R6nAE5dkWSIyDmMzgWbgIaU1l
usYoz1o7BiESeaWuUYQ/pHKXpKUaKkgZzC/IUgzHH+YgVMCvd31NUDlHsMsTbAAx
+IZ/sFY0ciskJ8LUEO153JA02XILNG7WTJ79gx3vW+FCvYjoJhRO+QKfeqHd+NjB
F5qNZ9lD/v6RICIv4fBx1Pu6z03lO34P1tnoddSUjD9Lev4ZewxwwOKOpEBGkyRV
ReKTPzshHTmzYgUTB/pq5ln4rijqJmnr4+jm3/9EuxnK4wHdQv0MEbguYZcUZKzA
utHT6iI3INHriYYNvdPgBA==
`protect END_PROTECTED
