`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5qwjmqCjHM81M65ntNiUwT75AKuu5Hh7Qqzqs5uNF1P86ETDqF4rc8vppcrbfa3
iblx+LfgLtwsdJC4GuOlOp6P4zm98uEkXZEu9corab952ysgKDkzlAT1HTpEia8V
VJgoY+YRLUdvN+8dxuG+fhZzsFu81y4X2w5jY6JD6RoFAmf8ICGW1r4lhGFac1eB
RNZ1LwxYl94Vtb2h5FPH7YkxISzsce8TS7UFfJyZdKZp0iofSUzEfIb6SXF8h27V
83Iv8TsGn+feRII/F9N0Hik8kmZLVbvLssmhkgywtpLoBXIZGTxAXfEP+eyFzorr
8CaDvTqMSgyWyZuJfL+QHDsWagKCO3M944/FgebALeSDBWADtaYmZ5W3jM++qpQy
Var4zdq6pR0Y/emMfla5s5TYmcWKjEN/O4uc6sGLV1sYcbNwXEQJ8jxuhYtbUbAZ
Vyip/q209JbMs4uRTnWXPWOUUhqOyM7cXvEty+C2yLFR2fe2zmRvoeINBEEIbJIy
bq+JTwgHB5ENOCB/P1fK9B1+APCb2Po6Cp7WNXUeo4ydmPrWTyr0yPfHyYh5nFGc
iYASiqE2yto9yjqqzeFaA80yxoJpfDIuAyNQ8GqUI62dfT1So9iLGmJnS6F/iRra
FUIbyHayAzKnBWBsBnnRWC0J/Mb65YYxhwPMLOihTZD2k53RJ7KdVVzhsz2H8UXj
kLOD5c2iUI9Qk4BtskplI0khJth2uZ1VMtyYBnHPY/JEItEqFR9Gdo0t6oprBIhI
u3OvzQmiFPb3/pE46OgCXJcv4VkyrewfZRSnTkd++i0MlYKA/slCEW/WxpEixJ1L
mVOphmF4yBEXwn2sZynLjppZbJ97HX7qb+wreahXraNcguoxy/3/SW8/euIuGkH7
8gWlXPEekNqN+7d8bKfskDP/rETJXiaqfHWvebokKxn58rhrtoByLzcn1R7E8uv/
n1egke9tmjjZ5YIpz7If8d1DpfKGobfIpib0p+UMlGoguFXAddjZFLBEShC6Y3IW
RY840q/LCpQbVmk7gaTW2g2gFpukCoY+VDoC2KE1m4OJOgmsb+9QCfO3RuwbQzOV
7C+qYtF+eJXzuS+uOXQfRDoHdahN8qTJ7D5s/LzTGWi8qYx8LKXr21VitnVKZCNt
tQtQKcx52RRC16+xomiGR/iC5zZSAnRMOL67hmkRtfMhqBukxw0r8jlhm6IXz6Z0
cP8lypbRHX/wlOFCQI3zjSEwYR5KFpN8HemcbK5mVIapgEGx0ApWjk7Xd9dxAe5M
aozPjA6tyklaV9qcEEkTgLCaxUqfUPXGnMbAkUVGXWCjuaaUEYEKxizzoBCYKpGO
AZsHMiVnDJwZtI0AvDTszQEF4yN8wO1275yaozq8+w8kaLcgkIZcl/ehFizYpAHu
yyhLqkSwG5b6nQEZU2h2e0WEiCquwLzJHDdX4a7vFzee6xkolOxWHSpcw8vG9msd
0lpe0hMGGgGQf+9AsVejyWBrwFJZOlzXZWLMfdPS3M/KvoOMjXf2Lsx118FTVdqx
iNFcniMou37rB3Y0D0GI3vw1UYdmYYSHr7lGLwKlNUQgYQd9UMDqXw5vW6vwLQ/2
FQlCE/d82/EGFmFKlAkHQaYy3ly/UvXqvSqZI/g1+r5Cbp0E6W8jBFWsiZE8eijy
Cfa5OZsdGYRAtJSxZoDI3mIamgouQVIMY/A4/u9IZlbPOPf3yKV1ChNSIcLMhTPa
EmnRXycIn7HYOmGpHV5i4Newpcb0k6XZOa5b8XlSw8zMNN21teWZmVXIBrEBFILE
OBVGX+qwRniAYd1Shr5st5diCQpGPamAkUXBx99AcmPmk58WcHH0N1yOGgf62GkI
RlMYi0uaBros1MfGE/34mObhz/XJ3BGrLJNALuVoVbXPQHtxpz3ZThXRWdaRQ6lw
WqIplMUgL4kuit5hEKZmvhOJHBgwLuLfEsQh3lpQAlc5aYbrYfIoTG9i+qbVAaWN
YfkYL276ep37vMu+0tqaK48i8DZJK0d+UP6AcQ8QMBwmbw4mwBUoNqVXntK3mGpv
2hx9A5KPx/llSS71aQ2Ke+nSGwKquhHHj7P4iYtQTiQpfPEWbFYkpb+22GOVPwOs
zniTAQIj5BSTcgFbPJSSOgcXjJ50gvRbB8BxJ9/CdAjWg5J9GtI4zVEj3hni98Tu
0X7BFKvc77q9DYiHlCO1FWovgpwrK/7blIxCvcNTDFDceey6+AUyai3pvIJJ9WCl
xSJ4GpUEjOqVwvJudSkV7/d+ksyBKHmPpO+Dj0XlhlOpTNQE4HND1yFyZV4oaMIp
VhFLCPjlSRPV4G5f4XM1uu02g1YIK+BJIBt2Mg8EYn4im28dlW71Lvzdh8iRSZct
zB7EGITMbRAeBknxZxFlPkrIvQDf1gKqitXyEHaql178wwhUEbnsHZVZGgO7aOsc
ubLh/gDqFEeHnVs7HgVNniyRiAvxzTl7XbCUFN7xrm7b+POFSSXVlcOqDHuoK22r
Ug0/y7nV4AJ/RI1yk6vqTuYIgW9L+VHhuK5SUVqIBrW5vQaMAkC6Y7jqKPr+MeRx
TiRTKtpO/I4vRloE08sfsUMn1QWbxbCgkfWB3Ad9HcffHCw3oScjk4CtDMf4e8JR
gIl91jqzoh5NdKbYnCXJsBJgqmmIBpXplTcVQ815nh2pn42nddCFfh8H0/3GewbL
q4PYOKIu/OrcJn+X0UZfrssDGx4LdNPmUSCvlAKAscCobK8GPASRF1smjBrsd2eP
NpTyv1K33Tc7Jalek7TmtKZPZiFR3Sdic2XLVpiUVpjjq3IejpONiepxwB7Hi6SW
7tddzc/EAaLbVJ45hRXa/Mr16g9IgE7vzRBFcx0/jzsksH2H0IjJUAQEm85IgY6f
RAtzhDVIjA2GiT0qaB3rfMjbWGRGf4afoS+/uullkuRnisfUFLxO85s9Okkrev1t
LRACMwBAy0k7b3FNUDARequNBWonDWQcCg3CDrUXjT9jmyyLBU9uNnzL5GMLFo53
UlN4dNTTsSezhtTqfh5mg7IiA5QGf/lk/lZbCIcuHXVgloriZfx/tTe8t+r2UHA+
M4SCNN2rQLSjeYK5d9ioaQjzuiTIjfiz+OsrDKAOmp72UFuXsot0TDqRckDTmxuI
YXDEtgi0Nou9MbHoTIRn3SqdnM1CGap585++j0BvPHiYtvZY6HL/smhiLMOFlCIB
xK0cC3TDXyB2vCIt9+tAfNSztMPpSQAAvO6s8nZ41OypM5A0ZrBe/X9uosZ3y0IE
1QpWqUfZyohsAcP3HNR88ygVa8pvmDfDw6yFApgokmyun+WHqMyLA/qHbrIZCzQo
LhvkiNp2eCPt8bD6ROthvQv8fZnYIdwpUWIpyWjLmI65O9mxLzj2NNHrcZFvtf0y
f386K6il64RZsRyyE5L04MelQ3ORsoDDJe1VG/g2IfdHlEpPf8P8Zyw9xWstPfec
Ld8qk8s9e3y4PmcTBwg+0lmkn1RKU4hNV7QCu4vKeO6OkF5+frmVW06IGl3Umi/l
`protect END_PROTECTED
