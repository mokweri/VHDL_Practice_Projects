`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CREA8R/vk7vTqV7CB/TvYatVaNAOtxOrB1Um94YS6HgIdooMWLbcbN+bKa0VGDzh
NPRFrB3Z9Yk06Z+o4tSUsa30NipOGCmHWZo7uCJA5f18qs1b5jVEByLkErEay1de
CtE3ICQrEmhGI6ctd2LBPo4up/0N5b0pRhKwIcr8CX5onvnJzYkYGdprPZh3PFhn
bdEVCR60mI/otoQHIgf/Z0Mrz+0F5SCA6tClOcmTElgKGezBAN9OLhjBKoq/yhnl
FuhMoKQdeMMmYIvx0VmakYzW7g0zk3PzEIVXKj+3EsJ4BBL6+BhZhHhEjxSsGzId
QoaF7IgAOS5xG5Qy9hbVGTVpV551DnVOvLFmVlX4rPuLgOJlScihFSod7TL6o7lm
ys/lTGB4Vw30d3VydEEcQa5a96+6f0RK+wTraMhDidWLXJ6lOCUiFhlXlgwEPDKQ
MjGbW9vV3l5ZWZUWu0H9bbLm3s+BVrOo2hszTcmGEtA0uuzUoeVOYth3pkAyWFX3
5KKTc7ZXv25gruARCN98vCu8hG+bsjcjwA25B1beNz0aNDsS1ew06YBgNjKDNcj8
yee/DWX6eD8htNRqFM8+Xg/P/JHnij64dQFcO4RdFDbtlO+win5fYOmMqTq+f7Mm
/nR83ogLpxc0PCpUewXqFrcB5jwaX+sON9gGurEbPMSpYfwe3M9MXiFpmueRXOEc
nGzsXk6tIJhybRkos+2ftabA/qnqwgRTYpxRWjIdY40W9rFQFheDXKra+im7iuk/
5drTPW/oPDRHu2/Q9UFEIg==
`protect END_PROTECTED
