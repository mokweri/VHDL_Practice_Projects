`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0Y11I3TVHTEO7NiC0GIhLWpmi5ZIUjMyxaJUiRdNo2lGmrLVBAOg7F5wrQ8am2R
fV1FqAvmSPB97QDA79uYoEGMQc+lyD5HG3gHRiqe4blXbzz9iK2cbA6q8qlZOmnE
wXVRB4SIuaDjnIVG4uGs7mk9DBO4r7ZS902f3Nrs2RibLk8kcaD/769IXg+Kyltd
JMI42aJdux4gKdnyQHNe/OmTDo6z5DfHQZ65aO5e29FIypaiN1yXuWPPxwuOjYgq
NqTD6xrZl1bTkSkcOlPOe2XAdwZPGKLTW7vq/wN5FLSwgmePoAlPeWPuvOWVPbyE
ob/QoOjBYQIZ4DxbEnyGwmQ+xdYmTApci1SR66xgNneDrUjxybIo6Jy9gvIHis0j
N5tBDQBc8sYRIpctJg32ARPqfClXyq6XkicodXBf6x8uFyJ1co9y7X/CwCkozHDj
2wf+RCRLHkHGiXnmuAGG+DPr9ptNVlIkV24xeJoEpu1V03qbvLR5KTmwSXMZcU1g
4U8g4rzIFQ3BA4T295lhgtox9/9DmqQwVzuKoeNysCVCHsBXSy5+BHhUo4wkgYCN
t8N1kSNZ+MEWkxwfnBhjUJtacRIyqc26pfTV+Hh4FMXFQ1wVw4c2vzxn2G67W6tr
cof+wB0hZJIjLEnM34p1w/FnPXbc1ZqbcUwAHJyrJAmDwnmfRday4I2cUCQlBUwq
ScWfmQG52KXTi8rleGmtPmeDqDvi8V4eargElYC4Jia9sOaEqTCFaN5bK1zvHbta
vvUBu+GKuB83+OWCoBW40GZi9D9oELvlSA5+SGp2tFM1oqJooOqAq2fWlblE85gz
u7wCpGne0yoAhXZf0+SbYmETageSp5iBREUDk5XvK5l6Be7M73nQ6Jt/d0gLzrVO
/4Z76/vnOoiW9ihqqvTWClkigraYHK/iq4NjRub/sCSKNP+ZCX7NVJKS68+2JL2B
QN3t11MVUm3T/nJpDVAYPujFeE3kNGp2tdDrQjgC21KTR6PWcyJiSV6QFpi7EXfQ
piQ3Rm2pOzoPTNAPUWnZOSm0bMrExeKBWVL0EdRhmI86DbpMTmQlTDbNwhwnGPd0
iZCsDRJoZJKGkHJJ5a9TNpEsyArBd9CdaOTopY2SfvHKigUDE+2n61IDgG/mG2qg
2i50P4k7jqfokp5lMTtLqha2dZpySV8n9veAuwNvQpOftLha1apAxRf1S3qxmsXA
XWsNzG1NlWfGMDJJCIsmjZD7u7IwubgnhgSa5JBxgovDD1trR4ErvE5bqFEmLduT
UJeLjZtc82gkF/TyV+FljEO/tHLkqW+05F4k+qJlhz2iappbLhsWr/ZWaOgUR7bh
YjiY07kcOas0Q9kxV1WoPY6NN1Xb8PZsMl77Sob/SBdsvpl+/yDeiuTjyDmGpKb2
utMJ4txiVE7Li09WBwQiSXCjk9h2d9EhlJGwOouRn3g9Yt0RLWHak7z6sQNejq3M
7UQKljPA90h0tkuLEeiF361IprRsm9pU307PWJfrkETgVFcBBfL09K10BsmrywGz
mLa4HtFHEkEuNthIQWiHSasuSd4Zmazz/fdI++FtcPPIkCUmZuV9Ur0yXmMXXAUj
JFMsZ3jB9+BnJbZxxy8K/1460WZyFqTL7HiMXdNjFErqKec8kMJyxKpBMrqzeD0h
fAo/Lf6GSWojwitR0H+dBTx8P2ujQxHqiOjPAhGjDSNd/CYeskM/eGlcZlQClcph
FxLNW5+1TmkW/ATwPXE14+/LRHTuShVg8p45HP+S+4Ytt03GXb+/tSRxDFdGYwth
I1VJiznSxM4rEnnvsX8h/n5iSKimsQmZC7HPRezHRYw7FDjQ3rhkD5ZCvdmrE7ZM
pscC/ivmpQfA91aE1YsMfCOg68gy+dtroh9cp6AeBbubpOyWlg0ouGm2YxtX9SdQ
80iEmcznraN9bsCj/ZFhjmho+YKPwH88iSkA08zjSrGVxzZc6RROIFvlJKqnwbaz
MF3aISlQIx7zIxbYYKESQt1DTCed6YB27Iij3iSjZZ/tvtKmcDvd8nX7NONGm9/H
Q8hbXovm4tjGdLMPvWVi3MzxTNO8EUFTkTg0X8N/Fn6DXVnsB/pBRYDsbbTIqzsu
ztSyBK00V8+FaaRWxI9cVXSW/4XUvoEygfbZs/PBryDV4HDh1nu3Vf+Nj18RnpS1
N5sO8dINjznBTg0XdhL0r221aQq5ZyyDFWrtTwra9oSGoR636VLyrxr/8AJV2hpp
dak7nISLjVMmxwS/NQAtUVAj465L/qqyqjEqK2xPVxYd7Ka8qprcAord5NXOisvA
8jMbhSCwaKqYub7sLjP+ylJrkv4UieJyevXH7YRHLiiLodzbBd1lCRKJpC3T+NWA
ZhN7akZPtn6pS4pLmlIJ8DDCm5yPAH924QgXbYSRx6LCt8RokGg+7WCpAu15KwcK
+ablrMh+QhwvoPjEFUW+r9YsWGg75qAZdTg+IDNB+fASAk5syPfrF5ArgarazGS3
XtJwbcUeOvApYvCFR7xTK3ITW+pdI4ZpeB5kRt2Fj5KLrHJZJC1ZRIC1ZGjpSYSm
AKN5cekjAJCHUrCDKl8TzqeJr4ZQAuypj2KbuArGhIEmcRnwc0rAuZKFFUGhgyvs
PSp4DtPxJgf2VvhkmJikkZStEtDB44TI27g71ArNEJRnYT+0qURXVc/cJXgwnb6A
w+UBQinx4WnJFgICN6hGL2aUpzV7fFludYkDtyR/5uFtuDhqW4f0J7KrPFKIDF+R
u83MHxTNfJW6gne6MT6VIqZegEctOhqe44vKFBZyMyzb0AnzcGJIP1xfOK1eLGpe
zwXv8ZWxY95rwxCIVG/hwtTsjSRrm6rxPph7fP+NWwvaWDKftQ0NAbmX6oZB1nxW
y/QeyzcWPUOGOWwmdtSdlg+AdH6WFOFG0JfmZzAUSu+NgQnB16AzvuSVY5wUYq8Q
KpK/w4r9zTqy4LU/jz1dKijJtpia3dMi8b8r1/OBwfsu0Cc51YkgGpUhsZ3G0aS0
Mw4AqrVy2Hcti32G3PfsBATG9G/w8YZJeSyE2m+dFfsPzYTcRYEe9YkT3YyhsnlP
KBszSFc5qOqTuNq6R7/3qcrB3Q9mT58qg8YUdBwScJlWY2OPHGS58FB0CjsRvJoR
nI+u4PfJlu5wSSK3ViSqxYCAgSXaa7iZP9f/lvJoAsF5fVhI+Hf4WxKDfRUaBuCm
SmgS+blOewz7G8WttAKJ06f6QBVb8kzS5hAiIUxS0Gs2BAa7SpEa9ErpHCwEIMFb
egyzkzrC5plCgcGKZEto6yvgLkBwtAk74PnXT4u6xBrhpf3RNZQz/7IXU7MSIJ2B
ylVkJIGGzseyg5buYrdZc8zJLGJz5zv2epal/ZO1sAHSDBm/zJ4HsabF6RGV1VVR
tF8IQlHkICVXWs7cp9x9KdqtYeEZlMTQhBuhuNQt2Tps/0JH2/le4bImfiOD+LvL
Vh1SQdtwLxWA8K29+lDOHxKHcbpKHuRI2xK9EF+3V4apvvZ8nqm5hHWejNfkWShq
0gQCMaZ2iGx0DNBMza1UjVr+EGgKyoD1BRtVRSye7ma7/8RQBwduY78PWOj268Xk
1XJcLv652MFEgFvWHUEuwoHMshyZLSjbwpbP5wibjqv84sjZWeyIDAuesrae8ugq
YlyAdDOZ1UG6jHcJa/pn36k3S6OVGssYHq82WBY06CT6FfLJDlE81IUaYLedlzNU
lD/ZMD98K+VFhnkjWu4wA7N/hYjB23cVzHUXjzuWfk8EHW8yrJ0iC5NB71G1g5MQ
cd4A89g6zd0V001b/hQrXRKD9tMycnAGdH0tzJg8TRXefhrYEioeLRXt3XX6lfEV
xC6k+njDhaOZ7t4dU6Sswv5t0IFI1OnB/aoImLDGVWJuJhzXTz4br86Gxa9jl+o8
v3Js69uIOmthb1TP49sS4FSs2ubqLtUexhxZWntl7IXFmwxryGCi+1MeCgoBUYyx
PJVoW/SCfz62w5nAC4iCBDnXOh2taA9dNkaeDAut0wvwIhDJSooy+vqunZ0o2lzW
MgkYFBZga5gQ9aL7i/8b0ARr2wZ/0YldDopNoNsTZh1u4Dx7GNF9MD2yts9OuwIz
BTmfuuAzPR3ZOArzTlkdPSKgXAz2iVEC746pks1Ydkg6tcucOVOyjgqed7q9Wacb
br/LAGTjO4qy9OT++p0uIGOEcHN1Jj1y9Tx2x8BvzsdOj7tYlWQS4lhdfNFsCsyT
y37BJ++XViLc1ELQAk9BrLHiXc+IhFpOKUrxl1fNqYifNVnK8UQd5nJQa97xBk77
DqJHrpQXo4kIg+HM1Y4/js0pFIahlKVp/bmFpVnYW+DCrPYlcikz/9aFDAWRZMvF
mnCpfIWS04pgnU2JpEkM0bMm3xHA3G5Uh34O/WU5+zgL35ZXuMHS1mCJ/ZAFbMj7
bODSkwguqqInoSftulJdWYtnKX65s9sGNMcx/5dB2gCYbBtjo/1ZrXti9S39vkY6
muks9I7PxTV1B+GuhYHzxVWX5unAlW1wmGpUrI3MBlsVib//3S+7+dvOwfKqiP9U
VMgiSEa68CXo6GM7CPlhtgkSfLoR65ZIhDoOLjyeIATqHeoFPaU6qFh1OKT3S30E
lL6zd+tEa/9Eow9+BC41cV52B4+CxVQo8fS0dSloghb7MVgSKdTzXllwvEfH/Jvv
VrBbrgpAlJ4lgvFeG4v+egBnPdv/ICZM/vTfsqjGZFYw7QbfARnlqdLiiLnCINGZ
6HlS2xVvW2yrAtDMzXvk53XvyCMAEsPJZ5uqKmymRkw56EEj97pi57j6rO8UXdyZ
gJiZHqkXxZz7oAiETSA8ytUdQ2BpQ0GI3cyB5Xz2LhejO8QkIlE55xRDoBtUEyvg
teTutp9AOECErPVJWqL+C68Lnq1FlfpcUuwzv8xTyxWovXlqZOxeHPmdElFcs4ZO
iim8RKlpErfJctfEktkwVZNViF5BdVcwO+Z5hPtGyNLQDMhQ+CwJiCA7RpWyjzXi
cRhZq1cp5YYoD7GSGId2aswoFGf8aCHpnDeeRVOobPgEDRlS3qf225dyf01trmuN
tF9hxM5wm+MelP+B3aGdnbj1GZpNDZgnTOsQaP0Awu4UQlFpOGMSVoLMOvr9Daj6
6Zyq5nGyUYLbntL6te6yD6diJXVTYfU/N0RgTUHWwg6C3TbdcMoF5avqL+ChWZrz
Iv7rj3f3MXLFwhXvPR0RtKJ7ycvE97RThk394958DRViQTSm9AJsvckywyoDi46m
OvM9oQXef6mZ/k7YbZ3/mZy8EMmOUhFHBg33rJjvNbuu2pAH+rsNRb4ARzzKON+P
uwYUHuyn0E56NbeGgjBl3Vv9jPafj0+pAyI6FhdBiF3H66E/Umc33jUlp15saVWz
mQLgrO6ZXlxqG5vOXHb9QOqsZfKFxHX1/x/wZBTF3JyI2RQj6gkFBjt97r8QTjAa
sS6v9ibtWQz3s82QOF7m4g8TKOo5q8aQxOxdG9iJRgHHk9VIyYkX7BeoJBokzDYh
TgBZQpbEkwfvtLzgyHUQCxLp7pM8CmJKFsjwwkxe9vXQdilEcgozejrQMlmPx0FA
loZIqL/F+CY95M0q/iDWU7iFuqBVRqIrmf6YVvDu0LHWAGuRYWogEkUtOcj3LvE8
9fEmLoa5BHkfjzrilZ0Ta8SBXhiw9I1XrifYBhz0QPb+u60aR6W581SUfAiDXlPo
4TGbhNvh4P3srKRSWP5o5xiK+4PphvIVhxuWUipS4JZEecuWoqsU8K/THvsQLycl
8XlrOfUuVjXCX9EKeu8a8kwf7nxqcmshYYwV8u7L/HBRLTughvBW3I5XrEbLL+in
Z936O7om9ORB2myXtIpqnwYbgXrV57jAjk/gkpxuQHtdwe+DradXyAEs68KxQWnQ
tKJukd7QuEF0ERBQBXRoE/eOD/WswvEMaZqnJ0yl2r6qRkngSr1RSB5kVQoUbQDz
+lMfQSQqmIsvM2aSL0koN/rj7MXXj3tHgiWU7ELDsaakAH1FWHFMOe3a0nJmrIzn
7IihXbKOiVkSW1J72yOpaXgZsl0eEkAWa5wamj5Zhg5BfA7FkSGmSti+PF2IQEiy
IfMgBFTCADqL3SnwA/ZQgoCoNwGO12rHGX4/UsiZrCuMz09oQ2ZYAHe6pxkbuUDG
UqJTAJ7PapJUNmGjtYpMR07B1YSM+bo6rMQIeGl6jxKcn053ByLuHvJVrR/KZRiA
Om2huwcgd7dnvJu2y9WLUABRwxZXaTUOYRQPgTB4SPpO6Vf07/9Ec4wizGVDaHtc
ODpFmwL7SBA8HaC8XHP9O5wOx0Jv2L1CIxhJKcaKDAlYT8yXRm0zxEfDjH4ZVPEX
Pp2sM/rzq39kLkXBeUJRIyF7m1CZLyZNPd+JLzAUJXkOUZ+cjLS++WGkJ6ZwlWIO
KJYEjjfkBPAjnZPrCtrtghmNa2kogzc6xAa/0zb55ZB8iBstdunbnL2kxMOABGyu
6oT9g5FLbpzP2cv9VBKHdlk0aN+I9aJe1P0s2TojmkQ9pte5dFIwBynZTd+yUFWa
cZvKy7pgkPRid++buxy+ISEaCoqEuPtF2QJwbHe7c9Fp/Pli094zLCAH01fJI1e1
PAaPvrwtobpw1U+5NjmsT67bNREEr0VJhNGMGOkP1IDdGL9fg7WUOyo2yJsg6hjB
on8VOJSKJoKK2M6DEkbzBiHFD8E/g9nXaYrsX92pLXfskTpiyHi/UOUq3tBfpZtK
Mt5+CgfiC+FqjAlfupaDlizklgCmskTuC6wwirVJpL0NsEuKceZmHF6NugjYTY9Y
HvGOtpZQaivDM0tqWJ97S0wMsG5HE+PlPcXSi7RDmPeL5+NqROVcIMxRXKX9VIc1
kZRgkoor4fpCsPAvq1AALjx1NuL7qmX+h5PV1utMv3RG+7YpF94CRR1MCKJANuOQ
/Vqe3BuDJVpaGPiX0KaZE7vcmm4cMOAE7C7SwsGrmtWvtN6imn51df0/627aqGdd
ehU08E847OqHsHBn6HrPHG9sguoY8VohUlrkOwZ4ponk07SDy2PoAZBJL+/xu3R0
KpbbbPz9NTTM7Gxn0vuBrnBxonhiSssvhgLTwj64B3J7jAx5tTqN646rGfjn08HL
PGCdSo77gqY0Mso5zjzc9g71te/wgmmMl3sn/5lpg7bNaLTsMjZ23/4VtCjhiTAo
rsaZXTNgiZ9VhOm2G1qhBcJ+TuiYskzQ0Zdl+gYi4h5+dVPve4bg7k0jbTwccMUh
KmPT75H53ORDmDC/xZAIyzE5gXijD6QjmcfxIJG8D9XELpfAJz7N+24NfpVz2jfb
siQUOomhY37FYR0ncYuO694zHushLIIZTb5m7aotmZvrTbW/xcfHgB3EzjDEdKKG
4Di5Ca5ZvJSulgPSypLHTWCN2e6780tF+BUdermzjH1/DZmL1VC5+R6/Y4BFWaPm
/qGTNiyGSv0obAeDnDIkXDgCPhi2vliSrqwtg3AJGsBwEUNa34YkFrzW8Zc5ts+e
GlPJAM8q+kqoTpbWefHlEvjrlVde0vCNS1gcZWypHgf8szVCoc/euMF9imH0h1Sq
0Mnk40GdmJAXMMITYHITvcRDQsN5a6gBN4MxZbOyqV9k0ZpaVdEZwKU+OODI7JRR
BU+osU/Zxl/+YdfSuNNKqj+KlKFSRkWB7Ke9sVOJ9ArLekxQk03wG4HnQROYEeAR
veAOqDbbpCSTWFIzkCauSrKqyW/UZwEqYO0vf9OakN9tHu0qzx0d2Grv5PokkIT2
TOVNX+Wo6cS92ELI9Y6asiunmpr4wSX2aToefb77r5tYtkKvFLaQpIwgN65HADSW
2/WN8ekzTTXCebK+hNFF9SCHm1KiDdfb72aJApp/19W90/XYpx7kiM/c3RSf8SfY
T9tRZAUy9G9ehQkdFzgzTpr3WBOR6oYzGXhcHODM7GW5MMdWYi7/OmyOHMG9dgiw
jhOjthZZCmr8VaPyGLQyutz3xn2zM4h6ET+12QJloFIFAR+aLaO3lp4JAzNGky8L
zUKPRNHUM6wspCZeJUjXqO7ImHhqozRLwGS41nn/V7ITzB4k9NLAY7td55QXHssu
xRCtQHsKNhqG74YaTN43rll7Ahom51tr0kaMcV3/nUmQ4GmLNDsvXQoK3tLx1CYT
VevuVW2oY4UlM6LP8GsNem31do/DMP1VfpIbmZx8WE7BjsCTC3q2KQzdud4jHnWq
ZNE9WaNTZoWtl1bdax6egr1+bohE73b+7ARylcAOq+HRmauHc15zGB0Nwz2W9sSY
1F4rYPuCXOVHW8tmadUrEVIvT9fNjSp6jebtwHQ0BBO7s5xjEqNaIYfou6q5mpwQ
EJ3dJ2TGaUaPc6Ft/3SKSur9KDczVtDdjMEefmsoEwzO9fFxWxuk6v5KevD7RQTa
/oaTSWvQnHqq7n8i1AGJiDpGMirgwJMiOXi+QLIxObqEEWM5tnnRaYNLAei0uKS5
YfBLfMGuLHqFY8L0EGXPaIHCdOmjvAPpLaulLktIWCA/zSGoMfQTQYSjcdjkpIRG
qcREhgSQ8nei25nzKzEDJuw8a04wkIihFuBOBkmuDsp+MyAJPkXtJ+7AVgsH8Z3h
VT2vgmaIYLMoFh38am0cssMGdFEcBk1ExBxT9AAL9tsA5lLSTZRbzInjb13DRHVv
UoOZO2PdZjNGoDk7JtbJTO7WZHKu3gYpCubiEy904ebFPALp1YUPSEg5Yfwp3wg4
Oo4zWKzVZ2a+bQ+auYIIwu9DDx3Znk0q8Vi1nV5OlhOHgvHlzNuEJszBO+TsFTyP
bmMjGusUC3EIJ6ESwjZqoV8oUTRqisiV/VP3TFDJcg3mmFJIhsJjfyV5Vc48nMdV
9NM/PwRDvCyULLa9+Sn3FA3CSKVg3p6AGZ4dZ69s5k3s12Qj/V76N+5laXcLu4Or
fa6GGbgWmrYmIi4LZFLngfvVoW/vyioejYJeWXCK/TslAw+8gzQJUEkvux5jb/Cm
E5NKoUgQJzB870iYHX0fe8NLnpQDeZEb0AlIjGIf/Yo3o2RptGVbRdqZJdDWHSjX
3m/PTheFgTUM8nXiHu1XGylS7/OX31V0VzLCzXlPJFCKvNXkt7y+iYWV9gnDbJJQ
ZoiZayQXh+AIBp0W2JUQi0/G4GPCr+ecbMF2alKqmsmRzA+8nZNRqtjWOzfthVVE
/VoKrVcd70aEgg7ntJvnDEvrIhb9x2j2qrkHxTLFeuCNmc4GHej1GuDn9mU1lULP
LTsZ7a8/1Odba2wF6hMdBqgp1xqh8Y1bgRiQgcv9VPavCBWYHP/sKop41dYu+KTo
BAEU6VPionCnfxZbjuqTQnJdbP6eQt4L1/l8+2RNyH9H5pLlbdc8TPc/lHrW6Gs+
gwtz22U+9x0c/qB31F1dIMk2iTF4klY10rfwRjA+u96bf+WpZLddFlkoJ1ofLxN3
PkESBM805fveRRx7AUlf+YvV84r1iFRVU6nasnM7HHenggGF+P6GI8jFhznJ6hrW
vOd4w5NZzeNYqlD3NRFoWmG7iatm95bS+yw/D2EjB/CLcVkuwvDKJL8AtNIyj4Xq
ckU41HTTpgVlvjGs5LN3E5B8TOzQjELtCKlfrWhmQhrvBn7X8hLCCM/QXjj8YnlM
bIJVbrkWoLSBDJXjFoXuNIfCEBekQbBZb46sswWoVqOSZsMUdWC4YIQb9G7LeNCZ
ulLj5UNL8oYUkfwMFVXMVIroetsYouzY3imZ7NZ4/y5y1Bu1bkzwerInP5qrfTX0
SF8qu+WaQvuSM4yQbCo0DIo8OYaRgmoFezAxCTzOSHa6QMT1aLPcIrk41tazLYml
S24NlVVwAwlAP8Jh/Wtxt+DpDaGDc2yDAmdFul8Ma3iz0+t9bcVr1hlHN7KgTePD
lK1M4XsIL0PYhWskNu1++V0/aFiyt+kicDv/xkrZM5ShG9rPx4XjSMac2WoNLrPu
zxVvrty12GtIkAc1Svu0UxLj6TEkizeYDAPysEvjKFmX4xpJkykV0fZuxBRcl6Sb
8jNmsvdBDbUac6Ybc+XVxrs3DFKjBgKtELXUarlqvr8PUhfXrBT2g0LKmQ/25mak
oWVVvviXM0xbojNT5pMShjgT12QDGdYDy0OfdqS52FcJsTP10W4X3rgMVD8ddkcn
Dyvjyl6czi+TeSrhk1BRcLAaJBrp04RwznAvFdkmbD4rdVmM2IvPRBVkEa1RNApb
sUZWPxVe19YeZUZF+VQceOU7r7k3gW+8E2bzvP1x/WC28jeOJKRJr6YF+9RVgjCg
8M/WUmPNkSbi3PxbO1c9bz80SAqoKSI9ugkJ2XUYBxgZ1LG2Gs+JCVi+qBuWfB0N
U9zYEpgwdkllMdXAfezMFY3QKNmX9LszzHscLbFmCzaxFy8Ol2uud2fNZbUKd32l
uKyOU3tlOA+mTNH9+uI/7yyVTI8n6uk5v5lZGRiQZROPfFhqHTz7VGRAFqawYjRs
/xciEzsSAm7WmBnXmW6ZzxX/bGJxjjY3ISzuW2REnoWEpEFzrWJmfj3oU7heSOpG
Qj3GNomrHDEI8W65wW/oUSgP6A6Vpvh8bUk5cYL8r61EC19xTNLyvgXjLHHoTMnK
2GuIL9SX/FPPrc0gvThQqlJXe3/DJzApwUVHVqtceusBpt4ZxUkWaDReCbyVVEPN
iAm6QO/Jo2qbniXHTRaGIkFZ/AOC9geCVs4fOnMpA6dEis0L2Y4nIYdHgCO/KFPF
K0w/87BiSt5kvAIWYw37BZVR8L0aqbEFBoFWoNyEaHlxku509jixcRg+vJtYK2Ab
+Te72TakiXs7ZuRJqDL/H5aASOyJlBQJz/E5k0wae6tK14TG34XV6JX5kmvHhkwy
Yq56/IVxzXz70L/EvyiDl0i5ePY7nGtClABvm0qo8bGVHTjSDF3rhnIq2oADKk7i
p2/6UCz8dMgVxRwOEtkJ1QFe8dQp3FEJhJF2xSTxSAhmRMBNs1t8MfwhOYG1Y8bQ
eV7a4Xdq7rc4J1UhFrKDccNLQY7mIil/Cy53TfdBEk7R/XKw+wEpTXocBtPCTZJK
ad3UllTBm3XSgKiOlMQaOx93A+af5rhco+OsI+s66VgONwBLezxXuSPXCFZGQf91
7sVMNOOZGhKazQl80i68yWZ7Osx6RniO7K6ENvIm8TjrPJ+zlPknEZj99Ig1Fl/T
2MYkXHdp4NY5czSkTnje6/QljX5QcRrNU6IVK6AgWzcVqdJWlQQtlVPJtEoZ6XN5
JgDmtmq0o4xknSObtKaGOm5+/APoyoe4+1cWl59m9CZvXyk3hkvrN4Wa0OSb/nn0
mgx9aBwbZxUOEdG7/oBhPtwSfG8wVR4qbjTnDZmROx/K09BAO3/ct3Sa/6efHOQL
CjnECzkWzSE4Omevk/Nr++iy+5/jKeotRJFLOP6Ss06c/OkUstWEsC6t46WUKku2
WKme051Q9ykLOTZoerZOmtJNe8WNs74wlfmfaa/3gHUDQRPDnLXDlwYxwoSxfAYA
qKdTZ+5ULkYRJetpae0J/jzJbtPql74h3aViG5WAenLI94gMovGOadPT6liPjQXF
dn61CjWgtRes4gaX4Ju3SQLQUGh1EZfwBua7Wd3GgGopVO6Mkl92vFEnqlr8WFjv
D5bQYSe671EHgmFvSltzd2YvIr5GPJuSEprglvqsC44cyVSzFZ3N6OcH9AVPuQVW
0nxkuDU2yRd3aIGlbxPGqLgFV6I2YqLKdVT4Yosg0hxcQJhaZ90s5uMSXRnUp20c
TkwW9rObeBAhMnEElMORkJGIgBVG1GCy+NvQbwcBe3imR2gZBidGk6Er9r3vQgpw
aZ8laY2WcqhXCqwuYOopt8ZF09LClqvd6rtOY2ocXgVpr9ONHpWsgbfgiQiYLnaN
7OYw1JQaVPCo7yxIrgwqgWq0hQRFmlRC4fxc+eUktUm0Pq+KlmuEP9KkSgafq1VI
MftKHT6nL5qbVeyHjU+W1n++O+w8+XXK65WNoP4o2Sc33V3T1OroF3vYgnInLbHh
AsXESBdpYhPnSSg8l4sIeWCrqm2IYYQc9SfV7hjcq7lBYu1Bl65wzUQAdGNRD/Hv
UMWEkWrs/WSEiSta6qb7tmGFKOOrzweqVfGjjflVW7o8EbswcClDEn6WewfpEjeS
H5mShIRChJcmxOOXt5F3KyIuT7maFDic4j7tTUIjBi7Rg0fmQlgiaQurWC/MNu8p
7zidzvTEVaqWhO8S+pdszoTGT/teRUoR78BJzDyUqeGvyX7NRgxjzXFTgnzxwsb1
LzPlHhwZ36LWb4Wxtkx8SGLg+98XymUvD6QqGP6IHmbAO7l3MDGzD/aklkKraNcQ
28pg3DWX+owvF4s/dvHcaf0GRsTLuiqAjGVPjyhPK/Bcf/ABExHnPGRXmQPLMlch
fbSB69P3krPVjHiwpKYtiB6GdFdzAbhBU9VpB50/2UIG8mBv/lctWnlRNvfpruLg
/FQLKFXY+4fZAabyKzCYOx+NzyIXpBu/Xglc7w/wOsD1jiCU56YSA9jEA2MeDjOh
8O8GrbVgySlrbr+m0HGjecvSmBSrPkS/+KE4EbVkUrrTUFNmjwgJu2Rfsdw4f8cK
8Lv5WkJ8QiwOf9iK0RTr0zDcfDCh1EAaIshNBkgDIQ5K6Ii7n05v9jF56J33zb+Z
LtdryoXS2Sid3z6y+L6pfGx1QQBmQ7aJ+5AST6f1ER+eQPYFm4Bpmyi/mLWcI2kY
U3wdzg5YvV5r/Qd98FevUIND57JSMxcn9Zi541N8iZ7a1JL5hK15Yd3Is7hWWbvm
lxD7qH1NLtYEy4tWizqMoWoH27nbgXgp//ah7zz/BCSPwPJfk/031vEtDjq6Wtkd
fYl3kJ49EK3njocMAeY139vA+fmOry8ppOMycz95QJQG7+rfZ2VsOA/mJzDb1UZm
rh7/DP873E9UmenbtV3v6BnY+Cfk4D/6E9CVdaqnf0sT8oNBS3Fy0rJQb40leJCD
tHDH8E1XEDC023c2TGnui5m1NQFzkMtS4iboXt/CJ1OT4cWNBOPxSlqGMXSlhSk1
hyYEAItSy8ykor8h0ps06YEoFNWgkn4jwzKhYCX8PTz68Gn6FsBx/YUew+ivN3mw
rnwqljSZEAMDQQJdLeVeAU66DMFtemYOvAXvXWwJht8Lbbl70LIN3PP0hBE64LYm
wRPG/MaknqTAgG4YFrH7oTBfwLPVm6Igse+NFjlXXbjzFJrb7ShgX9V4PwKxcWiX
dKTkCZt0dPPQN/Kt7DEPbd3DotxNL4uU1n8df20y2LZ/8dLgZC9TDhaGWMhNBXmJ
otSPtJtkbJFJuM7xuJO4CPTwmSrLwNOJZeHCQQcLm5dKy0eAmZDzjQ/0iZfNS8uh
oY67wgzngIDXSw15k2WE9P6dC4IkZey+C5nPt78bnsiwJw8MhZ0KQlgABnr6pZmk
YLbQEKcBOw5stCb0hAjOSfqCqGGKQuuX86Dj/zElts6wDkCzctlLQg9vmsPMqsJw
v70+TJLPAWl9QVjLlfUOqKJjQsqVwExKtzfKDsP2B6GynEA5KJnVLiKosw5aUbkj
1ktknO2TecYnmxq56eL975wEDRdn4e8pRby2pzti2qTo+D9p5TO02Lpg7babzbH8
gILTvrwLTgWjbPIK5psoQXbTZBsRNvrWF5ZJIDkAytfWZjInv3r6UBI7qMSanQEF
r64YLTEjQ7JS0GxX7OBumj3x/6QifXEJwJEMISBQ2C1nCH2OWpy1UhHkOOQYtm3N
O1aQTwFoYEPxDPgPribHHC0r2kaNqNASPSwxt6KZg9+kHIX3kzE9t6cU21eNmbGR
BlO8Df3HlDIKMZ0pKDWWR9RreYUr0VYdfLg/GJwbhgGnHnqoYJVkm0jY5KPy8Ga0
M22/FK86tIBXZllrGKQSvseJLo3GIybMxa2NgkyHtMI7PJrZzQ400T8y0ctmfYAJ
P59Mquy9tkt35dK+KFnjlK1moSlr4wVfwH7LZgZeNwYejHlTfljM76JNpBkpJew7
kz/D/itC9XW3RAqDuXBMN0eE0o+Yqh+DnnHAPqe01FaZ290g4nMXxJXRhERPNJxp
S3Ir1S+0iDC5P84h7GCJiaPvfuVINqIUr+r6JrtY5zmSGZy040+AaTHyQdxCDJCN
xhuAUG2CNIVd8sXpOFXbgPTMqD7NHA6vuaAlVmd5a2yNz237gNA/9Wg9dJiN+w/8
cQ7qnkbleSzB706Rf0NZNxJfvPxLjTrn9nexL3aSVsQh130ybknjQJztZHPVI+Gb
ssMlx3cQDcnLgRl0d7i05xW7xTgWAdoHdMYP/If3dutvVX8NUjfjgvNe8Zqa2+xc
fC/WY1BjCLM+0uCObilWXll7JxCdY5BTSmOr0hVshHPzMj9clOK1kJaUzedc2gFj
BHPPe014mSDCoDqBJHSJ8V3eJwSiZD1M6IqshQ8B54xzfKvLdu/U1I8u0TLXPhxN
kgK0JI7WQF5z4cs02oogMxxB0M5ddbt9N8fuCMbOclmWDryg0AS75mU7lNizEw9j
7hw1m27evnmoFoqoRIDKyT/J8GkRGYR14JWm8G6Y7N+jYy1zG5KL+T2RLMtqP2Vp
XFyYb5bubgpcEJ9f+1u2ogE2upR3dZmrmjPNEOzmEd5sFXQEyrexHscapx9tpyM2
5Odcu0Od+lwKw/dgXoX5MG4hUOSmX9D2/G02oWJuHpf8ces6YBr4Vi+gLzW+tUEg
EKrRBa4/ZKpiNGimErPd7mgkwxwZIh+3iMrVEufvC9Scg0QIvCnRVz5XTKc+Tju2
7WzGjVcoOeelc2JiHlHY20iWMvUQwCjc0iyWPy5YhdCmR7Se4N8vfs1IvioHIrxG
7UYFbttg7G/K+JjH26vBy0eoEC+g2L471SWkyvZmlqaA1pX9IO4tebJIZQfosFr/
IfGdd4fNfs6IgVY9dyqCJZeGnNsf3YcalGi2/XKqkJZU5PiekWgFtSlIZOYF9NmU
jaXVbsRtKvoCtJYWZ+VidIwK+TsxvAjvTuzV7wSbCoD8P4FSNQcm9LJvrhHK7re3
YQQXbNcuNzz9T3nBIOWYVCglPOxetQmTTxCaVqHS8FOE/usJJTSrAs0KhWun8HB6
WWei08b1D/KPV2XXf3Rf11+0GpZSGLtLkIPt81+/vyExiIe7LLzQIWO2nZAJCchQ
Oo1JgW7vSM4A/K2mLRPx/xeJf8+xU/0GaBQM9qiZOGn1j+Q4Dl6ZboB7I4SXplSb
j8xqGGvE4qBhrbbqSUhy1j0vy2xrb8t+v4bB2r4ZKV1Hsrh5lO0wyUeeYFFp7JT7
Xzb18QTD9P0K43y/piRMBmKkzFJ9p2psL/CAhuG/1TTQfEsu6qeyn39P/AmJFFGf
Iv+/d+wohvy31CgCAXsX9FDrFPSFwQdoclQotwIP54que3lVivnvMDedMCwAQUlh
8aIkXgHSIF+cQVi8pc3zHpQs5gmyBcTu/hdxRwUcF3AmQQT7eV2pbttGBlwhuozu
9K2AA18mN71UeTsHP9m0/tl2ym3paZ4qhwqV/4HWug+pVSmNPMOK5MVYeh+5PQV3
lv6UC+bMzqNr7ogtE5JfDjqHgJi8vOwocgZZnaTP881TGmo/uK2Po/4amkVeQaO7
qxt6IGFzsoUmhpjetKhZ56EgSfHOA+ugybzazZfLPbOuJX//ftJE4GzQQiwVWZhW
YQHgw8Svm3QayZ0DbSsMiDph9o3P9NN0KLl+fPt0kjM7yAugY48YnKac2FGOvLM2
J4A057oD+hHR/rC5KK6bfwmok6W5tA1/83A6kOzezZoBNwKG6yEdiZ35RlFovpwA
f3rbRXx3CWH2MnYVGhdvHCE5Q/BshuiPgzLcPCxLG2/crdLc/deg28xqXHB7vQsf
PsBdp7bngN84W3hd3xPy5uDNE/DcQkDl6lDtvVunAjGnRUJrmtwAejG7xjKD276N
nmH2h9GPiJ5p5xIo/IAwrMrQ5USD34ErLc4Yb4szBMDjOFZ65HSXdH1/OJdkzOqy
anDWKoVku3ovOwoKnYTQSV+fronZZr+kQgJ1T8sVNVZ/hpd8tva+wMO+me8hS+lj
6qvRSQ7acEuAoXlSBiSrrpMNiPLZgMBAbNfW/+d5tSzfFLWfyb22raIImuauXEbD
Th3szLGPvAkmzni8FpTwT5PBgvF7UYktEX7J24pqp4E4zmcwGEwQNiV+YTxCZ+Kg
r5aXJsZwzkIZHBeJKs81lJTz/mYmQgqlvAM09M8ymzoGnLap71RGwjRuwHwa8d1+
kgLBDochMCO+YgTJMyihXHKT2PNxTJGvwrNiG2TlhSxtRgdp9KWMJAcNRY291mbE
kSJf0uSgb/UJ1AzCp20TGoZYXjkxNDFLHZubQ+gBpHfy0LCX2fOniJj5BoyMsapp
CwWqa6nz4nsjPadkLhdKX5QZrgn2aT1kv+6lHOsStoy6++f1uQbgCCRb6AfEvb6M
og47P7qrSnm1fomI6XGzn4polFTrUsMZ00L6+ucgigY+Q7hPtqhaJsdJYJcJ9BOf
TEV+pHZzjG6I9agnBHKv9GmjWgDNID9AY3TJjpR2QSGYdD92knp25ETw91PTsmSF
zHskL4w9SZKvMVEkqkBVN7w16JN4nWSiojsHfzxm0o1f4wDS/2T5YtQvmlq3SdqI
4ijDYmPG2rh8ZSXxd4gQWIOzo/Vv01ULrB2Ml2K6RBxThq1z/3+qZiSKty2DHdyr
akoZC08mW77q8Ncq2IZ6yhFoPr+E1UW/RjWQw8p5vUR3WBOPwI0MtfxNgHSd904V
nAXwrubklVfh/Rd8fMAQpAouGv/yLeQquEx7Xo46yzmQ4Esb8y0GV4udl9ZF2phZ
+nf5dJ0lqlVRSL6tDfXuqCfTsYwhu8fuPBht1nY/4dqVHmzffJz296RfN5KjF9Sr
VkrSRUvYSrmG9fCYWZZOka2HxHhQXdTa6udbTy8eVAjnRuEjUJwrz8Nb1tEXPjKJ
m9Gm/DaLap4gWtbni0k60HZbXlMF+4pm8mS/9EidCRROdSFH6o0iMdhidBv6L8Ie
d9mgqG5H3o0UquJAQ6zOvq8RQlLX8s0aiqjrdkPeFRxVWA4Kg1VzWdPeyTYemroG
uH3U2fQrS/iEQcQTeAjdbxOjGLYL/sPMGIWTwfsPHC26i2ch2CFU49hHij/p9H0D
Pu5oJV108efEQcXr3h5UaMecAr5a4ZcwFEg16md/P6nknsCkTskhgLgkEKGniRwh
K7NzeFMPu6KutXDYTIVt1yFofpWwv0N1rrBwoILTZ9RHfwzSDH0G6ew5FZ16PYDp
EIvWsfDTMtcsBKhMlnLMtZohvvBHVLHT4BQfGQb0wpKrgs3F2vCFg6u/v8doSnil
vgW2GA7eVRBSFqXmR6+oHrtzrkuOuoKTz6kE+jNnbRjHZ31epPQKZDXX//jhoEtz
PZIBlkkatMk6Dy91yeIL1h6W6STBzKe1A4Kxyp38Z58dq+jrKOiwfHUlATS8cjJ7
jg9tduuPHY1MXywkHc3+wY0vObyOyKVimNVtg4/XQY2svq1wXT/WljJWO4aVbZYn
ppJZ//7IegpKW0uarhkFmoqnD3YYK4mstHt+A3fwe1dhZLFYfQ5aWO9WW1wr0ZN6
yEOkPdkTaQp32cZfWEoUo0SKIhxHBrHs9n3j70YWVHjbrRjXpsMzL7Cj0JD8zndx
iNDJRdA5J8eZEpASM24gVk6UUWDppDR2d0ci3rHkmpXnJXmmTWrsCTlwKfv+D5KN
LT4ewUDKMvaBTUksOzB0RKNtP5bMI6Pee6akfWKqF1BZ6wzQUZshKkbwIM3BFKI/
SOSiD7kbvamOBfaGXciK2uHNYxmKiOxgXiSQsDsX/X02KuO2KYp9QDqrfsaKVE4R
8rPxYqm6MJb4Q3dU6EhGOE0am2LfLwqW/viR3sefsIdIZbNkksEdJKceXpG+8+L4
JllMLVd4gXU9m7nYAkvzvxEkhB/zE2I0kBTrRHmB7qQDvJ4Q+B0rJO+uvH3I6tbq
alLdqVwbb6HQgPnffRduI69LLiptMY8FOS3tW/OjjtnnZtz54oHeg0JSGTnQhWrd
iXwboPKCV6Y6nosrhrkbe7feWF+E0fNaHy8+cl3ntymTFvEc7CikvFnYWIuJ+T/X
zJHjNLDRccL021LsWMxLzfkP9KFF/mKABYbdQ0GVYRQsHgEZePcFqdjISRX3b+02
7xWYirdEQ+MvTltAm6EwemN5SH+lyblQf9M8TAcTCtMTvgpovnPNughpk9t7dS16
+nHEhZtY1RtyhenVJzUEgzE6xspe2AkuYkgr0/H6Q2hSf/4NPTS9nZQjH+Iwvxe9
hsG/pihNG4NGJMLOOLE1b/ryeY9+jYKzRD9zMt9TXY2Qu1k5LDtThYvrhq4t5TJt
A9DspWGP9UODejcA3r6cOJgEDzk4ykGgZEfUoULRUOXC1wkb8q0ccoRkPZ5JvK7k
jpYwvI6PTGzTQ2ib45J52xbUOV0dCCbA2Frtx+3fghsJ7/sOemQQzsQ6oTxVWCf3
ZJE9HmvtwdfYxYyqOyGsL6n4R1LnkiNHWXd7hBO2awRchjWfW9b82v614lXpN34A
Hzm/X/fKkZ1uK+J3ZLxtfVrnfv3Y4P4hDf243zD5ZSZT32OSEPyOpqeraivsuQK7
xldtNVt1WNqSRks2slXVWdi2/PsROR8V8CNOey48CnMKtQmFhZL6R9w/oixwYCmW
ZgjhIBpBa3T214OsnUh3DziYknaw2LijjYMDf5Y+7MNcHrLqaxGBzUMS0tg1yPfW
np5FCK0sed6fb/mL32bPeT0zB4XLCU1XOObU8G+2n6j5fcUQPLLO0kdwKsqAiC3D
FCtRLUGr2qINWl8k9J64UJxigaGJiYBXsiMIVIaF9AUUOAQdbUwqFfOoy4CY9EOd
dB98jqvYssPUoc9FcEXmvmrVlsEk4Fchke5IBJiUkkkqYx2Yb0NGXXNWkW5nv4hJ
HjGpq5X9K/A7eZMWKL5DIpB+fOLcVnSPgd/ie/C8Z92x4gruCl2P75r2sMwdxLgQ
CeYQw2AeFT3mtb4zpZtfYbDN49WbATKgf8aO2xUn8tJJgc49AoFv5haPidNpXSY7
5BmTbZHY25tL7MU5zrTC7qYOTO4kLE5NSM8ClHPGfXVelZ3jYatomhzK+a6/Mj0Z
xsz+ofzg4GzE8CGP3cC1o/4YpiMtDDm5gEOupgBhxDQMI2C+OjkBj75yMeOMivQh
+78dgvVc0crHKjc/aRhNekbweqwaZkz7RVQsQeia2pmx9UJzQaGeH7o92PrCmhSw
70D4FFJ8cm0JrXYJI8hAW66zU0o0pWrTy9ypxmmMsu9pVCUndY43uOyZHd2G77i8
MeoG/6ro5mmRshFkUcGKlGG26uFSyjZU7LsXONcmLWNNKgzouybqqITnYQg7/lq1
oSBKpWwoiWShz3bgmSMFklokd7JofGk/cbld4fhnYKj4j/mABFF6oDebqGpfTQTn
2mhTdUqkBjjDQEGWHulOgisBytWNf5OhN3FB93gt8Mm+kkEypr4YRpu1E0ifIp9v
+aKJ7bzJer3tBmFPUNSeZbBq0CJuU0iUYI8dzL0qRpCOHjTTKREiIYGGsMwucLXu
3H5Ab4pkZ5+1fMxOiT/eLdOub7D3/Rn+4VrBui8yl47tU3AGpW1XkzkYDYifcGHl
KAK0vTvWNrjxbQL7zd8zk7DZ5ebwrslXlY6VR+UpaBn1BwB7cMUK5Al68sFtchux
snmpey/7gxe27/EAZkKVz+zl82nWv+rJIrfyQuoqhqq5thy+b+wnRjx9pw0/ESzM
6A/y4ii1RK4BRAnJ3DN/zE+Lck06wSquYKNGpoqsiyklgyE5VWR8+mR4NLZvNW0p
QUrlHdiT6QOC8IE+xTjA0go7N1AQW6TpohAtIZaq52aRjAMLsNXBqWhDqNqdoTWv
WwyO4KqgMcCL5+xQ8oxukgLbehiqcG6XGDDT2Vwgmy4lBMgUlFS12kznNFbnPFOZ
x9tVkobpdR+R3xOUFqwMP3U34/sLGa5+TfTGZkR8EosmpJ57SqPWWsMHPX6a/Yd6
FjZ+yh25vMsfYMqSSCmRcOkAZECqF8ED5vr4jBdt4CH0imMeWf0uLwM4KcVdafpW
t1IjnXebgwBrKmzSd8w7YTPrPNYiCG7YwYeH0dgLViuo5H1oyAJf9+HovcSDwRw3
88OzFGNT2AH0a96gqaQVWvGRjoMgv4p/xfWKgoJllYoTwCaNIpqEocCRpKHvHnMb
RkZN8QQTYTs0ViyQzkbyEZPOixq1KVabTqxNpW3ngnQXhhnxmNHQmrNi4gDFxY80
ffuVnovoS6FPx4qEGj3IMUVOVO4WAhSHJPPq8n1WXWWoFQiX/WQkGjnsiJzYwwTD
3WCAevXdJ34fN5HU6IKWw/KOJFmRotx+mbOZe1MHNveoRL/dgfMM3gr5VQ3mkNLn
F5RMXHyVsJgo4jHxYkCWUznaSdBriWu+vWtvwr2EbjDoROcnzBCuyBv3Xoy0Nhkr
o8gIjo1ocbSQ/bK5kmfT+IG1pUTufKbTF5CRHIEpReLQTt2coh2t1DfCVi1TrOAR
j/fRarohVJuzPcG/TE9ttyHAYCJqtgBnZKbUvgVmsMPnsHCnD4XcO+/AWc0YHu5Q
nOc8mu3NAe5WCJKvLvzeLOaTTDc4iEjiczrh3JUyT65/yOni5NkFQ1IqUcpwB5sX
m5cVxCM1Mzt8ybxbRdR9QL7LAPWVnyBgbLmGsK/jDUPZx41Jah9ZOCyO6ic69/l2
jdnM910JVFSI0gJzs+sfrtWx8t/iCzxtFTrKouf5eiBiazNN4AVw2AA9XDsDiE0b
j0CBbw5zoAV9Un2Z6sR0j8WXzKhaKc9rEZ3IP1VliYyjnoWvkNPXiVg3HsdIKjZa
dso02xMJDKYIeKGj5UJZsYnK5HqGc9vjkn08PyWKiaL2maE/qiwmewITlA2D3n16
wj7/ci50zenD1tGz+eoNv4uvRQsqPT2ZXU2bvK7IhdSsCUsYir9emu6jBgb014IU
Oe1RCh2PFOWYXRxx0dWTZXIU8aFKLdf7Cm4Y+mR0eHPmdgpeMSnUonYQkVMEjHoE
6ehppS7M0YsytUBZVOtijVILFBxrgJQca3+qgs0mJ5H/3QYeCgxnP2jJcSAXLoKJ
0XcWQ8z7P/WOcswpUbPGswByCRQNlXk7s9WEErf4iCS7Tao12pSboktM5vW2S76O
Wj53NtVYFqBGLax7iHnd7N2Gx76FpG1j0bCLqZF3I/ZHktShRNT5hYHUIZCK1q9X
Gb77bmbQk858g8Xn9yBZEtwRoFJUjuDuB9p3rUvVc/V8mifkU+dStgGfHjq53k5B
YB6Z+G8EeqqcBe4ap8ngfhjLftPhfqSyErieor3RRz4=
`protect END_PROTECTED
