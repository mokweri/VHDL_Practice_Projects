`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXKollZ4y+Nkq/OlHVwWTyPwYX1Ba+FMpfFfSXsRKM7jN6rhl/nBzYL/uDRgkPda
rRh7pc/sfx0w3pnHIG+jHmfV/6XorNrIJaBT0CS9SvH4vPfLC/Ad7MgQ8hfj1xLW
JrjfmdqvA+LKWcrZS2/Tx+7UWawUe1UpiLxawsuug/iml0vmVAyz8APCyWKk9ruB
gMaKBnBAmq2BRZo86oGACSi996XmSloIorfI9FgSMkKAyxruhCG9I3yI1Dfs/A6m
up85zq7wUfHjz3a0mjsbkCYUpcWo6J7mlu4c0BOYxfOCkylmS5ERJU/Nrpruzb2L
kSJxVQfnSdEmZ/24eO1oST0BIGxGmsITRwPvTkdiSCsrKKLC9YlYekeNCc7a97Ug
A895J80SK5GS5Z0P9/5pKf5KOFrqTwAI4DoH6kCa94n55xD8A+FadI+pXkO17+Kb
8kPJM0DtahrUQTgO89yxVAL94ARtqteED7+CLUOsGBUQkPy6LtRCTlVhDQ/LAGT6
YLSmkaVykUmiIc8sasU6r/WCJlL+7od/vpUcdRtMcjO863tGSozO+X3GvGkqQYZu
8O6L0I5OWRW8Tqv7wCqC3YZonLHxulfffIsLeXMS4WmT/XrWYAeiCNorFvVlRECS
SiJM5alMqq9VXlVrrXVy5UUhfzykcPFyO668zbxQjV/uzRmzoH7Nt1OBKvyLCwC2
UouVDf9Gbzi3wffUwpXJg9qeIkG0WEzljz7uksMzhg7Rmh0uTHD33y1S1H7QGupb
zKdt8YO6DAAx5GWz2rijZeGeLNoHl5G0qm77FvYTxDgJV57n8cuU6K+qK/LF3Tsx
VYsDw40y53kz/VQ2BiJU95tYl7aIXn+uMy2cqLpZ+pMTHQ3dnELnuMA7iGyvGK5z
ur+RptagvVNweDe7Cz3drpVLzBpn5BOYqD8ArSOcXjl1dDX231Mb7br/og+go87D
+muknTbLE4YAIcoHCTR6/B6UApZDfdkl6+OaC1a2vAecvJLqJgQVAu+IzPFq8SpY
joWMnm2lBdNTUFv9t0AWAgsc5W68s0GOWdxIH4oyx+na+aHdiuIdCRY36yFGOQd7
NwlS1E+5ppW4D6kzDZcrBMk+masxCgsDpPLG9VMNam8EoVAUshUVXse5DYXUEwY7
yG+IMdXW4njklyRjmb/iLliAoI/bqCpcwZE6nwEPhop2I+aHRXyHMC4XePFUChXz
iv0QktMSBc+tJyF44Qoo8P74t754ocxsa2ks1lB2zFPQ5SjXUiq/H9LsRo7RMdlY
ljv1N3QJd0kx57RMeCcdwczJnkQBPh6PJTruVRMk0zVtjfn0eZoX4q3LumMHI0fN
n+8NV2JT1aI2QJAq+VxOMwCi6CNVU6+EuM3ObwCNBDw=
`protect END_PROTECTED
