`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlJBKb6Djqt/onb/ZQLKuY5xhVsp+pMuilLJm4xXv1fRMQOG9jRFCve319sJcKXD
VPfwPfKs5Z2pTKh3s3RbU4LCk7fHsIBWIjNQPLXDQD59higbcr2+s0xfGHuN73dP
BLcTWFlAxIFP/VLUJMawqdeVGw8PHuC2sT3Pm5AbnB0cqOwiizROovz1bjYx89im
qETZJGFl5T0J67nbVq9QCuI6REHC251ke6uAeAtlPiNUwHaQJPVr8TNKymmzKaIo
f3VF6zS28CgZblOAmlSupBDbSG8K1HMiHRXPiwNMWtVd878YR3fw1J2mUzt4aRKE
iAFrE+xBm/DuocRKWFLZpXLgs/Me7I9fGkH8kLC517hH4V/4ZmAb9DCylLnQe80s
nZUEuhxieIvwyofCDgDigsQaxC6s8q9I0Bs+pCYMWiM8ywLdZGq37X2hTKPA3Umf
tChbFGJa/Z6iaMczE6vJdqU3EYnalUh4v0KQ9O/KXAa5/JZQF+vU+a8ng58dHjLI
gmR80Eth2/UjsMSESeSStEaVsA/BlDV8MGMRXL/XZGHFx50wL+J3v3KNA7PgLXf9
3o/82UbF4OOh27cwWdco3zU/fdH+eukt5lB28ueWYeY7N9vS9m1znMt0+qyG775O
SH6YSB5LCRIhNrd7BH78ydaKn9pao4pX0SBDYE+Mko1hr50EYVg7PZ/28IPfhPwO
8+ebqH3oqVL5nfhnD82dmaGVnStcu7N/H5bUKF5bU4G8eSDj28NPBqolXjdeKkj1
gSNX/xD/QRm0M457EI4iICbYIjG20gMwj3vRe7Yg9cM0X9NIu6cCnx9fftR8/SOr
wZx5VuGC5kqiwrj3grplMjeyDdW7IBqtM/iaug6JTtzhmPSViB//uH5AfplNQvQc
TL53BFj9IswMXVlsxgg63xJ9d/GLZIuLEYtKYTjSttgr/AT7fKDo3BntVoFCjaUo
0GXGMlkw2ZCxpetDOk5hlwS5wbXYVyGBivyx/KdHu8F/Mwl7wcfriClF+eGGsFfy
T/DY0t3RjemQLU/okVVzWqUIjvK3bJLQlqs6Twn0RNQWD/TWL5vEuQi7W14d4G3O
e2hYVO9yWkyFgx5JrJNl+sWVaQblsT93bLVBmsUii8jhb9bEy/LHjSOTRRNUBn/m
oENRk/d4n9OPD8fhU53Sd4zjIQrNSL7nBsxu2DiYalzI6OY6Gc211vtoDMT+yJx3
XeinWpTlJqVTnhwrMCfR2MEeuUkIvo7I1dZiSaw3h10=
`protect END_PROTECTED
