`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjquZiNhXnGDrpd1MiLW2QjSZQda8gg9PXfqdTOIRXhP6jwaEliNaYp7+pxAZHS3
IPVpFIjhw3T0emwXHAzUb+ZfU40jXI93FXdv7m3Cbpi2zb6ba0skaBQwaFy4HAx0
n4io/UT+yYTde/Arn2XuQ7ZJwxbpf+enNj58ULT71dpyvk/1XByVCdpw9FuRN/Bi
cRa8b3GtQSsIXR4Bt9HAJQbNgrus1ECnA6rMLA/2hy2l7iehjplh3qYZJ+IllfSy
qt+Ccfu+Rep2/Pkjg0/wgh7lCQbSYnLArrQGuWFjnbtjkYxtEPKLCI8FJ9tIJ6k0
A2nXVmS0HqfRJwVfHti/U/GkQ9cpkXZBc4ZrLl3JoZ5UYkbDdyFUKha15M4qM4+c
z3v/1QsMFpBkvgJZ5tP3Eb9YgjMGjCUWcJPaiOf5y/zcwPpImwUsOuiA4yM6fmQs
DJZGAwq+/pgpz+mvDmZZOxw+eLiI8lbOjXN4+qeb0AIsAmqRilKa4OYof7bb+3FW
0GWN6y0IU4VRe3pW3ww2g7374aZyXaNVV+UXAJsumdPQybxtqgaS8gbPSdZUWdSd
lBk703uO9R3Rg5Y7OakWKByJnl6fvIZ76BcK7RK7/vbOMirejWXh3ULhMNSoJxDj
6z7rY19dFedA2D53/Fc3H++1vNYOL03h1RW1p5gsSpx/k7UcQlSW5d9DrLsgrYZk
3Tzq/LflLzmzg6gz/1QhZashU8i0etAIjIja/pwCWmbrHNvGsfbJkkSyYb73PhzW
nPAOV8wi8teETy3w7mTZBAPAJn1rwnaLqEbRLJsUe4eyXB/iwePTDQuCnRGSkELy
mLLgE3ukLsikjtsN25VfC2suOmfUuOB4q3ubWO75EhsgclLkSlvkvyhfhkD4li7I
aCUfwJ0E5p9Wi8ukWr8EqUncHsBRh5bPsa76riBqKBf7oN4RFNWla+i5BS326W3z
AAZOmhiWm6GoK5Z3BD7llplAJqXBKAR0pqITIf+3bGR2YgUjRXHIHYfggUrydhIb
ToeT1KLMN+bS88DeZ+/LWvVdCyu62019WexAm5Iuk9pShHqJZ6w9/B5U1cN8C2GW
0ApRYDu5I5jcQKNiqgjOX51SWIE+Ty8kYTY7+S56UHI+d/mVfJZ1d8HCWsyjzS7X
naYNpA02szhw5p6tYV/DP4RX5aoRRnYN+dvguPQ0SeQ4SQybiDFsuviz+5oOFrho
iLTPmWyvLOsfPNm9Ad6OMA4b+4B6DxgoaWHXUF69/1njLh2vRLLIfGewYrQ9fCl/
H6cJFtKNOqGWm2DgPMiMFDCoiPwhVn2fFwbK+3ccULVslxQeHBbMF8qC8j6dJHEp
f/82nAr7RYkFfIeQgyRfj1BPekPThuqe4HqSla5RogdvNTh5N2nCriK85EmoGM1u
EUb6lo7Dg56d/Z54mWrvdmWtssaCOd2qqIHqg5ve92px2iIJaD3gLfaaJKgdWvK0
0K8L4/g1iBBmrLXgnsFJvXxoM4zpPdeGM4K5kF7JAHMm2WOo5bx2ifXn3GgEgIQG
KlkKLkNeOGD6r73xkb/VBZRb4rSItBLEYZaJnDlynt9c+BOwtM3S0dikzsuZbg4R
273v+fdQE/L0veY/bM50zcsCEW4ebMyvjgHazVLlOo2hC/z6+NKPQXAN2Wf5Q6sO
DevLymi74TCZXG5hx7aKyMA7cQdOoZ1L0QeNucJOLw3F9np4yBuonoB9hSZP6KHg
MkEyfW2LppYAooogf/4kf7lCCYM+l2IJFX7VQnSv2AI=
`protect END_PROTECTED
