`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fk7vt5DXWdRAPMnaWY7VKBkvGl+6+NwAXcXdyecEjhTG7/5nrmlLm/sxhfZFjIzV
evOY3rrFW8bTseYIqj/GmKQ+rFGv/QXrj5TBg25VgAnEd8e8jd/fPV3SEOr9aWcd
rMwjEX3oLun249fbJs0IcGV4nZhpvQwbfCe5vHxn75BKuPC1pxQBKI/fwqs5mcQD
eq2l0oGyLLQE+g5coK4AxDqeN/PXdmaHLBbEAtsMV5wnGaz+Vc+/Gre5Tcn35Dqh
knHA5PPSu8jZjIQX9G7mOJGzf91JekHUpt3f4CPqMCt8iAEGs47PaXtpO4YW0V4t
1d24TR6va0lgQ/U+GHK8g10l7R1ri5u2kfHDTkH/fdACFp3DJqjSHPUJ6UdXMjbj
WR1/P6GDBtIkOOqZUjb26bmRQi7bMc4f7pg9nYNcSUmFw/HTboQLn2P8gg1Ut0+k
NVbecc/1XvuFWgZFGmLtoQCfv9nT0WbFdFA5AZltgM/Wva26wwomW5hDhdtYx+x4
ufNurS1J9aUxXq4mMZ2rI8yxvheUFk2hmPPIBXsJE0iC5i4/Oq8fSWTp1pTkG3ce
gF2jpcesGUBOUgMvLWWlgIW2u652nUzK9vKkW9f/dd61Jnl/nLxHWV2pEJzeyJFV
lWTLhcW9FEO5pIJVVcoJIq+IUFIozaVQ/ZJALgNpylFb7Vg1HVTJ6pCMuKiIyrZx
fNB8S1VHOwCrymGlHaKt4ow7sJeGu5q/qIphIcysa9hnixLRUS2Hd4lgRkyCYOac
6Z0mBiLwhdjC4j/iUIpPJqbH5DWm82Lut3VAjpAeumOA7CSEYP3QLzcbhbggpydn
IDDIVyEEwPTLw9E4twLFKhIZnEyjipVQKXulqPp6WXvcw/+9+icnjCHpw9pZZkMU
w4O2cvi0uw12ssl7t1ZaZ2Un6hd+eL6Df7F6T3k6RZ9eG1rsffJqOt9tmrZLNa+I
4ebVQD4SQe4hjLVHZzkUf9geu3GxyhXVKRxoFrYewVQZ35OjNgjx/7dYKibFj+6a
ilkqgtmvzPOBaXL82MIDYmRX8/aexiOQVVcz4ZVDteeRYGiHZm8Ja/+oPGdY3iwt
qOF84NHQ4XbuzCyl+6BEKPELCckvOpJGcL6/33Z8syV0YxvjfVFo0Oc7I4bI3MfK
QXkAqBidKdLOVHRMA7AFZETL/i1Vf1v1yVj4RhTgI35M04SkSERqXm+uUCT7slFL
YVVvH/HRP8Je1/QDuGaAfti/GbkV0qflUkqgNZa2zg7Wwjx5TN7o3bD+9rvuo2d2
vFHRbIqHqDFLtSYjA/QmWpTqeBnIX34xyZdOLwm5fSqwp/AAGW8WseOAFnQmM81y
JduxF1Dj0gsOPt1Tb4EiKtasn4c0RWj/QYZvjr33pXWz98F0NvfLKAnIwL/tzd/G
zJ9a+kgrDy1Fdlm7+lJ/0BVkZH8A78CXoN3htQrK7K7dCesyE2tRh8gT1WbKtTjr
e8b6CjBcUXm1K2vLnvcrlgivOP+ZVDFqS47CarEe6Vw=
`protect END_PROTECTED
