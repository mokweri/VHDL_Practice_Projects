`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhej83UQtTdglgUPmuIFxbdTu1wIU7MQc879Do6fzjMPkycttLhgHGHyNWKmgvY9
Lc05tjHFK7btT6dEtApTIFRT254LgXX5G8p8x2L5sIzY8m5woeQRKczYcX21LQ6A
Ab2hqE0lDAws+BW27rIvvU+SDh4Dxslfdm5PA0mnlthuSnIRrMHhh27+3DhE/Kzw
UXWo81QeUry6iooVWNFUXQt3LCeKoMiR988BKcanlIq3m+bTWm0RQ2AWvt73Ayhg
VURC3FJXEQkq+AN+ot7slnIIBlPzqBxDltyEOlRpO84sA03tVB4cZkJJxznkr/BW
2Ia/UZa8lbEFrvxG6ZBL4wxzSAc9jk1EMEunfSPKNZFbA7zvKWFvegr7nSo05rxd
HLKj4SHi6xspApRqU2WgGR7Vq1x6xklOQtIGCUnzRXKtK8RhXunIuZOkrc4eTd0t
0cMV100/qZBTTnbuOqkvc4pK9URXnSkShrrl2VVfrkQcZ5sU3EMjkp/qD+1XoREt
J3x88A7WEbwpmRjE7LmZTbTpJiu99It+EXKks2NW2+JqndRU0CoeLfaYh5AgnTAB
QLmJZCmSgeKG08xasaPrgjLqV6jesJCvn2qSNbh4zYogO355S2j1nDli1h/gyebt
LJnR+EecJM/7dvdAx7COgcSmMs0w7H1haHdGLvVEr1ckVrTDMc38Z64M1aA0ylUv
eI42StOgNxVipKRBAL1OW3G1ySjG4cXsadU0pRoH/F9QFiv/0nNnCuZ0/LIMMUps
YyeFYtayPzxiMgq4cKK+CQ0aXXccFOWxGsZHn+8jRAniRDPegCYJcQrrK3ZI23qP
0u55VQ5FxCOOOHsAJZlTG+O0jx6JytCjygon5ZXk5zxsMALrIGOc9BegRo/j9Kd8
Fom39J/YkdmEKyjfGx4ahSt4ltR/PLjKtUjOTojtvZXj/2CnprMU4+hn3V8lRL2w
k4ylymwMFncj0thgMEIiYKgJ0GLf3XgI9jmzlnZb/qdHPYGUfoT3ZrJH9nbMCPgN
YX5O7jKQrxxwpWVa0WaCOpDEMCvBYp2HNGWNCdOblYXz2e9OwP4dpXPEmfW7Lu38
YiE9h2btrREJxAAvmXGfjUumpfzjt+RFPHl76RdxLgnAQrS36eDrKjbvPRk2rKSG
y01qRqaORbeET5fLBdvu2SFDX4fP37K30IzFsmy81gAEGd7lWOOV3MjnfherAwAq
FcVY25wALEDQMyeIsnBRjwTQTS+7QY+dL2vZISG1p+18ABf7/JXkHZWGf5OAubp2
U4y7fBCEhx3VIUeFXcqPN0XK10dpawZPRoigvnOpjv4zRVSjcfYphfeJpu9CvAnD
Tjfb+w/+liOEE6V0qN9lXBuQWM4ocfmfFPSbrNZtEGdixFKUim5pH1cAP7ycFTAa
OMRBB7HTP14QAXgvRFxHuz3Kf/6RgULdbwl2Xw7NOCZM8IArvYGz64ZAdSzDpTIE
sRbRNFnHeLh7Cui7dehZ780PhnBllGa9jjBsaQ8pjSAcG6Qx0i++dLTeFLm94yPH
ZT8LW8ORrm0Qspkf8SH8yX+LCOkC53jFI0fWhZHEFt+gfHqoUv+aT0MMJByubFGW
yYmGhFjlkwnsNFCO3VBRcKtTbkkAAnvqRzURJP6GrTFFDkIfRe7z1Ve2+S7S/2UB
06bMD56GMy4PcKGwsskPvfEXWJpqMcrGDiYmoZMN64wmoqn17EyGVAOT7ITbSBBv
nTua0fSe76T8ZRD9vIjfbqVXZ9vLDHC2MpFseg21tg+3JhheS0bL0zeqKFnod9nL
Bj0qIfDyGFMCwaNZZoNY5MgtmxWP9Zt+VLrS/kEW5BMg/zb1CBHbbimY2Y1UpmD+
1hfVh5Ce1t0ZDnDXCX6abOhCeCjKEjFBYqVB40C2z27HuT/tdOr6WnXD3jrJk9pt
Vo3saDLPwaV0g7JA4sFiohT5kZuCjZYSC0DETlTpF+Ub1szeA/yWhbFaE5iMLnNS
Mf91IR0zkHUzCvihw+WqMKcX1ZoZEo803q26zXa6tRSPu9AM7SZTJ++86BJsUMK8
vCS65uK7u0ObMvNS7RhFB8dsV4fNfuBMULBGQiBqwEJ7SkWoNYYzcQMj3/4y3Mb8
eCaG5G0LT0tHFZWRMFy4jeh3G0xjpfE3ri6dPJVIjCe4iEImgEGnpYz31KObZ5fe
hNzcGAZYAB4SR7h/VVcK9NjXVr1xfBaIEyZbgkL7T6tf0vR69vxkWODDsdFUldaw
BFBT3A20q/AyVgE8RbNiyJnGSZojau5u/kCxMAEHwg9rNkV2Fzxyzfwmtt473t9f
92PGxV1INxIOxnK/wc9og+cm/33kp93fQ23cWuPba/odNZLlXfiJ6B467qqWNVSg
FoFZaSPYIh6BohCGrge8ICE/A05uJ597mu/ANngEOYPf62f7JuRKWP1I9kltgGK+
dEdnpy9IDx8uf/n7gpIcVwBDD93h8p6jPYDarcfg0Z7A2fgeIADhQuanZEE/xSx5
7Pn+mT6ebmiMemRXyylOyPlyjeOG8vGuHMeVjwEdefHrYcsTaop6Mcy7bWwpxtXr
z/GGJhiNSE8UudHoFmatlb/X18zFvHXoZ/d6Nl+J4wbUCK2KdPmimrbgcFNEQ/cW
OGwUWjBa8P9vYDSpTMlLoFT+g3zuVTZw3kJR7AVuawB1ApcuSSUgJ19yuu9UmH8g
0q0MSTtobf8FulS5IRPe9Of6nU5Njava/BYy0Xg7BHF876/kZV47pc8zax+WnU1w
fLhl4Va4NuQP1mIjHgHbg47SCQ92VUKVhPCsnyCcP2QTawkuI4X/m40r7ueEdh9w
JoQm0PiY6N9KRBevHVqOIjyLTuolPDS1SHllPODOo4Mphn8yvhgBRL6CPAAOASD5
PAlGexTCeWBO2YLIie5FsiyAa6l5AjtpV7KalgEME3Jyr3FA2qLjZXJCZ8/qJ+Ba
9SPl/NDm16ier2DFaLApzgZj3YmOdGRxbTyXCW40UduzhDW5FE9+PGCqLnM6kmlB
lWjq7of9ByDjiamL1hdsMfUwtJUJtC9FWNaLKToroAZCZPA+8uTDP6+if3isPyZh
BiGl3PjzDC4IRF/9KFcECS2Kg7rHSmdg97ytSx3z0U1pRJ/xLG2jMrs3yNdWlJVr
wfIBAtHhqNykvwVh931KoDOoxFzIMXMvNlEsC4UTMmU5xSGvErs0TJ66yN+cAuNL
sU50eaEU/qBLMGST1JH1Jo+ZmaPN3pU8+w3Afm/2I8P1R0qwB6hawcBuAzCojaNW
DpKNlJTxjpfwkVlhScM+SzQFt1lY9uap/G/+bReQwZai6wQrwZ8qI0DX07BGqqgs
nMe1LKiqPx3vmg7o1hxop//n//vyZFhfcOj7AaYwBbu4oZjJjkafx3wC7gB/1vCb
bZJYWGaD6AWApHtS+HfAVSNg9r4jvp5J91JfJMHXUAS20lLYUMOVxS9hO34XPCgX
KLZER+JDAvRKPYAVvx78ScYb+KdvuvA2KAM9I0cmFBSRHaTtdD8g0Bs1WmO61nqm
wRevrNBq77UjTuBnRGdMkUhABeKQnW+Hpqf5W0ZMBOFw+esHoUfFO5Nbs3TdzQh0
UHwkEXqiOrRgD+byOts1piRooPCbW4/ZJlEWzbPHkHRd1xWCs5ndNu9s5q0ejobM
fAhsHDUbJwcJoGM967a7hXepT/gBM1q6D+Ud6e6xAbfUQ+ZnrL8ptlhft1zU7enl
qpNQ3LSaLjG09NLMAkAQMLkl9zphceHEl8c97XIUT0uP8X9pa08IFVqEdgWvjHwA
dxzRHa8zHEd84pYOyCKvGVnlAWBlw1+2TEAM3uQPOULmOV3fI/ICjFxllIkTgSCo
o/AuDdapp3EKop+YqXxmJfM57J32JDmPvW+lq1yMBxyjKujibovHU4C2/upFJVtU
ZVW1aXG7eYI2o++7KfqbymrZDVIYw5MfE7oXQzEXgfCWIS0r2ddyb8awIQsQJlQB
hoSkd3zZBedO/+iYlIs3AF4r6quHJI8nGboV6UUKjBzjLLSVb4V+z8cU9FabwZDR
RBUcshl4ijiPTNhAqxueeChfZ9Jb58Pvm3+EUEFFcTLBBW1SrMawMia3EtpC9I3B
0arvVBJsojVXOpAMHwVn7BzlnPB6xRl/M+iwGY/7bjXgAFyJR1zegVZx23zIIQlG
DIxklxt6N8BtVjYG89pLoUpXYqEEohldSDr03xSCHCh8wX7X1CL6mMnMkwF2cvKM
JNXkqFjId242RryuY5zCdv7YhssYAgPAuc+hSSVRplO8H9W/YtjpNKWMgSoaKFo3
54bPXb4jl9V43QEpsbkP/jAkakaLpOfmVaHmSVOxA5YRP4BPv53L0thackQO0yQ6
dXemq/7Jh3stjn5j7UA6nctcWnIKIJExsmAlXjJ0zsuOqZNTLgtImh7wa6lbqkE7
zvb1DaSukb0tTbyKkku51c12+VRblN3R/3i0fmjUOhvDX6bf7bbY1LTx5mBomzlY
IkC8YktXTOlAkAt3CDBvFeb4yW3M94ho/TuvpUktkgjFpMwOflTveKrDm20tij5U
rug0I17yLd9gZufDCT8CDqyw7gIAWJOA+qENc9VhgJzJpvN7QaNkZS6e4eKUzfHl
wfso5sMAn52/Oy5wn5PxW6zhILJhJrLRLz3GymyEgN9xD/4y2ip+pZxt2d9egsWu
kVI2mJt8/9blONclIeXtJIhavlbsd9eH2ZP6c687hTZLnt9CG5v2NTzeYcAkvzSW
XG4WyyjYjiC93uTPZ8YzzGO6raRJwFGumFc3KCZg19Qlavs017yP/0gTFdwZoOgv
t1eXF0Mz9duT5EAnao+Tx+UjhJ9YygwJfBZMNi20Bpnpp6aUflp1FbyDouijTj6U
VtzOD49zcEvJRoHFDRZEZOG0Z9Xykh30GFhmGreZrXAaAokHWee9As3pNkOEgP+n
rPdc9GkXxNXRXOK5xtha24Qz73hxFdk6z6JbJg+AQ3xTwF77MYNXcnZXhLzaBQsJ
LajK01m3hdoQuKtKJ/xfk2wb9VJmivhkp27PLENxSXEGgRqM02HyHrGNRCVVQJXE
MwUQi0OEoq7HNGzpy+aNSKiWpsPoIbHRIM0yUpJWNSOlVwiwSxz+Q5TsOHzedMm7
LEWkCQ05mNuqRiKlXE45OIQYNZUeRlAxmGdwmMt1mdF4K6hC0DTfrDuJ0gtkrlZq
BZyff1zdKcKXXf1uze7ERnEXrw/rWO7XGvIBSaGZJ9+0xNF14mB0816fIZM0bV7E
WUxzUBBAeK2/BXtNO/3PWfUAa/L0vpyjJZe7N07HPqDx3k76qrOrO1rWNRnzzmM0
rTuGpWICBiFJmnBKCcpHfAd4Ardb+3DkkFv7LY53NlEdVbhCbBzvZn4902lAiVkU
q7s82evJ1pjUB1jEAHLrsWssadReDxtkuwIiN80wSClGZ1QSp3N9nNeYDr4esK96
0RnW5Q1BJYEn0vqqOb2UETUpxxA7zH/kTtooD2nS57yW7SAAfFIXk5mYA4yDU5kr
to7rVj6t0XuINT18a9GimBo2NtvvGFmNr9AUC8zBHd+E0jNeCH2/dlxKk2IoP3Rv
9AgrmiXQOPh8cE/vq2SVunRcZKb9u1dHNWEo3YuCL35Ug8o2cKnNtpQhP2t49PG+
JKALo8aYEkdxvxMD0cjqxAkyZubcEnJ/uvCP6e93jQVpJAxWt9CYgeKnIIUf0SVg
9gWIWm/WuPaZsCbZwEvf3X9UISmge7vVYwj8Dpq1KgtqYHLPH9vUDXawa9hIQjML
mBRMGqwZYyiPWdyUPSKmJRlnB9LAXrCcYRsa5XOrphiF7cTwQ5WwLGOfXyJEdhMF
79lOMQQbcNgmKB0Bdz4fHQp6hEFeTIp6pr+XaTc8cTbXCPN7H6DjCouX8N4gycrf
pfKoBkPgOkgh8myj59+VosSqpRmHmO2RZH6Z1ZA0UcrfwDjhi5IpYW6wJbFPdrkD
InZdKy5OIZWnIEXe8EGQzhMad3pYTzQ/4FJ6bFckEz15uJljUn0NUqgVvq0F4v2t
um5W279O63SKfBEHOLFLecLkEemK/HvrEtPZD+XeJnwwSAe86ZUpHxrVy8BZ8Snf
lmOPGzLTVytWsBiFWlyWUeSRDTcxI/t6VvJduxGP4UivE0OY7JnzaPhl2SA/O475
jtxA4GzVGPWRrRxBRSZ1tZsnsdgVhG4XoJhY17W29QpHlRqnI6opaK4vykpYZtnR
4uN8GWG4ukufwhNeRX57wN/nNousb47ydYOPz3b0MeqV2fhAGyKDP1cOjAPUsNgJ
+G7s92uZaHGb0kB3ivv3tCXoCR7OVOCXZRMAQUgsH4UqbzTKaeEK1WzBCXDxvxHx
YBdUyjN+99DA4MVWFFaeTq8tRI2fW+tEiW4itNUNI1KEDL2aBmWwb+8iTPKjMG8Q
eVZVnr3YtmjBO8v5huBA188riNLrSxxlkIKz9urJY/Uezp7RA2WgLAV3xxnjroUo
E392dlPlomkM4lmpDE1K7xDA3z9swjAilMu6XWZZSmDxBEjJ/xOUUSOnU2DWb3BY
Bz28rqA54xrw53K1H9NlFpayLj2bJ8JDfqjrrA8z/+Glo9VFwbgKaoNdlNbnrTPw
hnCeljz29wOsKlH+CuOEhIU4NLMnTJn3dajLw/6YmexYaTUThxaMouXcGBuBwMBr
u/M5Rfvgzl/8IuYwiacTXC7C0mtLczTyl75jkF9UG0gRfgddPLDbiC+Hd/bIRVSP
xUW4WN/CJUSsY4ExFQacwW8MdLJ/BcXFzFlymUPhWQSWQ+WPZcbS+Y7BjCY+gbnK
HyEPU8CGejfn8Xdjq3/CY1dxAiFvPjNn2IoDLYgnZLjKD5W6TKvwk6PRND+/KdRL
Ilqn1NVh5GekUliGOLAF9ItiLzldanukY+62UJ/gerKVxEmlGQ1z9vNaJ99k30Et
cBG3nUrCmUOv8mMaxyZt+/7/s61yTlFrh0Q4couZV/8KRaBwp5moBxfKBDEhYeEA
a4dOdpDRFcbddCsUiOj62jIydlhornb+68AcDgZ8Zlq5dkvmJqgh0QjBCAi4yt4p
ChyhSBjI3YZyB3e/VsQG6EtXQiJmyZ8wVCJT9p0NtcmD1ae+//hSJZNaDFQbrjKl
dYvv+gTEZ5xEjxZ6slCl/Xw19D0fRJRRaZzGZs2PelDkjWShZwTfOXowK9uxDWTt
zTXUBWypgn2JNSSBsxXcpvDzcLSeOKESXznxZek7+nJgZ9lmg2oKRTR2+s4lBsU5
sTD/WKnO+C7v1y0X5BAoJn1An+OgGvqmETumUDy7a8wgpA8jJgjDwXsyr+CI9vnU
PcZ/yw5EIT6qKKxFXy7sViwxEJizIxl+zLHCF2ovvUAtuwsrS/V6cWBUBlGjDTnd
TO/RzrwO61Jgop0ngIIC9nJSWOiG/lukOW4uhYxiVQ5ZsdIEe+JEH3FohfW/aHC0
UNzjCH/aHvH0nMpwvNmPF/98H5bpKZE4wChy4OKxXYTtTF+Xmjn1g/uxUlHaNMMB
OyP306hLO+ZZUVrUfYw2S+wHCm0bTuaAterXrtY7WzWPhW6OjpWNypInd6tYWx5s
qyUjgOK5c4z8zWxmkKlTATNq5n3bfn7UPTZrwHOJqI4I7UgWGccEH7v51pyn+0cx
8V3gQ5+42SF0y1Loy7XyICDlJgxO4yruHXzhHhu1ofQfaHS09HiRfbEFpbMcsgY8
WRP7h5dNJ1qFzA6uUhKRABHsMp5i731UUvCZt0BuETJqT/AwAZS0Nwte4ZyP00gN
UNC1V4WpvarQI5VeT3aPG2remzQHywTeYF+p9B2aKwlU+DEnbN8XP6Tz7uBJNw1M
WfszW6r5VuEg4TzEBDWnjv6Xr+Qn969AckEdeecRFmu8ENFzF7RXu9YtVRrwEVzT
/AGwtr1wTEzxNFNzkz94cOHqaPZ7Y0pdDP9uDpbQLluD4El39Hk72R8OJL3TbTL2
jU/WJlo/B4qsreLMkkRmI13U/2AnOHS1FSJEdwQ/SzTaI41/XiN/dV3+YKC02MYl
+4N8xrBfAR2NUO2unmG0lXUiP9ilpDTkg1r22zzPkgNhKv5ty5bPiKK7IoT/bULr
ePwGrMaOdR/O2Ou3mTMVfz4btwkMMKm1V5tkXJCIIeOV70b58zUe6bx1tr7fp21u
2XXeAw4M9EJBSrkyoRe8jZT+xW6mcpd875paSwECnFAZeZNZ+rEK5Y1uhZMO4RvS
ywQm9ZCzbuwh2x/pb3Fz3t9amzUjqNR002W+vmndsMm0zanmk27++FyZF90bY85M
qWoynwcLZMWoy8uomh5X10mpCvSi8NspRwoQJxSQRHTF6Az5wvGhkDpJ0ppokn/a
d9yi0kyCGeucITJMyryRkfeD6xzeIzBGhZCy0LlX6/KePhGB5HBFOttbDyHnQDwF
RAsnG8oBz6vw1m/dZbi2hYvpkDjFQ1szYHOm5GrKqFcva1n9YF48g2gai8Ea6NP+
6rwbe2cK9oUXE6yKL1v4sJ7pCzP9666R+D6Y/haivkJ++A/I7z2KuulIfLyEAbW2
uNsSVKUCooj87vgSp2CYVk+dAG69lfW+tItoSB11G5YBQAogvi7qxK5DPzBoZ+N8
hmqBePNTGWJjHvTD5l9w6L9DboegroOCzxmqWuM42U2f2ymlegIMxsd7OP894A/6
MZ5lidWvnMuBcFb43lRoHwZAU0zMxeRFtFPX/OKHGbYZKYGanNejD0NQ3f4konxc
yB2eSPOWWE5Fro5fjr1A71kULH7DXbTSTgejfPBlX9Le5Gd3n4Mir0kBOQrLH5q7
iTrKWaUJhhlN2rdshDxeNG0QkQ0DZLwcL+F2Om2J1fPyqFBkxk0k2p2U6OE3SiWv
FYImTfiFuji3thwK3bLvcfTQuRr3cgmBxzTaVDkg2PRGHIUNwA3ixFGh9AD86Ybe
0yCNqcyzZC/qanM/ReBfG9D6m19N+O0SHRmQyrKpUvlt+vo+QgLCXLPa/Cpbx5ZC
+0TwnZlbMQA/s0kZgipgAJPbZRSmT17WG/5b0nrCQbqmaCFn/h/M1WHXlx74HAYO
Y16pvCmEJGiWha5kA7el5tjziMnRJVTxjh7N42udGtDAiX6AyCnSy1mepX98qTco
1Qf/o31/jDhVpYPQTN8YySpkSqfpD9qGLFBE1fmQdkzq4SWLMwTKGropyKox/tiY
3ho2Ls/edKCFqqu7rX4NdI5jUJHWn1CTY2BbRaD10VihA09N5++ru9KmQnjAC7XZ
Y5ULi2xSzQQUTW37AZAUWZSDlLAp0sCCyquOtglSOrHYSP6SyGyGzpIreAYrNKzn
DFJpFPPueJsII8yhVv0hFHELqqQzLbGUqm43/9nEteI7dpMgetCOiWeVNnLv411I
WfgCvl3UPiU+XTaEw8iGRkQ1Gt2nfUJnG+GDMScKielVhzJQlSx9KiLkolZP76VB
q1EvuNl+jAXiqs7yR1eOnHO+3W2C816XepVIcfiEId9KtLfA1+SdLQS1T3zWADeq
3MVhmPpHx7kbeV5VaJi9l71lOWHLOEVo9THDhh+1a2Ui6rDcjPMM10T8uB5pelKk
WUFZl59KZPNHkCzrHAtbhmgZUd+yyx3v5fK/7AvErP1hEm9zVTyi1eCTC/RtQJ3L
IrFj0OrVKSU1GkpzCPVEPt6wFTG8L3GL1Qcdm/568Q2oyCXGlEn2LpsXvEIgDL55
TVENvNehcL4kUO6PD/qCYmAZKskbmxbqVtAFKDHX2/3XEu1flYjoOhauskDhFAlP
OTEEEtG1L+mMjQw16tGnyHnmS51Q/cbLcX9Bxjk+0lBg6czqzPTgZpQ62GafpuhC
5D5d3FsVmciW7V2HfVqoKeQG+LP1wgTMRVgY/0YHB75nCcrbO1EWibZbxbep8fwb
QUTeH/fjxL1ZrcgoCgeDJuciD+88t5Ix7xYlKjmkNRFw3trJQyf1TH1zd5plV6Yq
WPrwyOKrM8jStieNQOYlRjt1fSGSDgdgxl9KwzokFKkA9pvPjL/+h53SxvxYno+m
uue7Z5AV14zIsVSQU/V6P7uKXmnOeoiP39lBhWjESvjJcORfxh77fnhGTXiPLgYR
2dYyCFLTKD+kax7nCaehzMeHQdn3MgAIXcsoy7OiBeUZCoB/BWieqbssbOK8oMhq
5VFc72UEqyAueN6AKv5SZTJWXa6TsQ7LO0W/5G3mKY+lJ/xgNf/JeeZTtzrwTAOQ
bc56UPZChhGB+hpMr6kmHpek1grOLiaQo94s+8mqfFSoYdTADQTKZn7iUgmib//h
ic2LocOueXvG7TxoC87JKniAv2MRc5UXlYlEJmr1/YeSI33MAq/yv6VdIKVv79EV
mhtyM19H2Hb73Cny+8n++mUTcMdbHjy6vDnn3kj/mxUP8bAv8oUsmyNflITD/kCJ
R+wA6MgYgHj7gRKZNYuktcEoSsGAq87gZKEFDmq8BypyrWFBJ/8/FROMxpOaBUBR
5tVpcMoY2QDLUi7O6JIqFxBo4waqwc8wFxesYHocvueIF25nu9OK4Bi2Fgzo+xrd
0xFvUKK216uRug4o7cBA9YdBGUoI77fnMJkaSViF6hUPdPlq0uxgK2JLPrwi2YgW
om5mIFZq2GhXzjCMU/DGsX1l7Sh1PirmHedUlnJRJ0R2jKhTb2LgMymoEnNdvdvW
hFTe8yp8LpHCAU+pfsdDWjLhEcoCnQzDh7gpN/nmrVBJUySIRjXvrirCJ5XHo754
YhBsOG6Lmh49/Fdjc4U1B7+9NjTUNcygtkFRfHQq52IxIh+JRgXXdBfTAH9PlYrS
YvTzkJTWC554/eDLGE0z2HHHQvZEXHVj4cwWnzXaHSAaed2+3EsRSQ2yJZWVb1w9
gybAcgpi6cfweMT01YUlyQ09V5JqNiJ8RRBARz8yKSY00psbFwkB4yvQZhXDvscm
3UYSNtQo7LVgwT2FgqoP2c32tgDi+df/BG19VNve9xB1KU/qmb7eyrLfPXdsAaIP
2KTzJ7n4an0guIVx1APVvMWLBh+RCcNQcjYnOjqVMzl7Bx6puX1U83JzLNnYgczq
HITZ3I6JrAeTaxQ1ac/9g5ztWgRUpuYYFIvTZr9kceLBFbxr6+khOie07YSm/VhT
O2MiXphHdY4q2bEyWfUH9PV200h81FyUX+LMxN4pzeWTmMll9rDG4ZrYlqp7FdGt
rpN+5q8IjClu53v5oQwdV/oLuYQzLMAX9XsLAsopCpXn8F4zv6OJPV9XJgqw3u2c
Jf7Uufl6Yz9pcdXJsUQAOlvi2KFrI6/vePWZYdHVp7YiN9pPxTLiCa5LRNVHiawb
myQROe2jRQwHZ8dzg25ECCstbX4qysTki2ZeciR+dK1GI9ojNyGjqdICZ0yl48ut
TBp+N9rr1zROyFwM9G2U242fjqyVgzjoIcV/+BKLhyvT0XBbECP+W/CQ9VArnYPU
kVlkdAZRCYWYROM1MOJeOIFIm9DQxxpt9cswoIYO3MAtMderpAiPB0amrdtSH/gp
QcTuCmMOTSGD2PuI3iqZlZSa28JJdTvJvMv/ZQIEE8ioPaV/Sl7sQWyvLWM7ioFh
URD85nGGq+sgU1EOcdBkI/4vlo0E2noQpJmqH9tTRU0VdjTn42LKLN/tPwtat6rU
FC2DCL+rtdVEfcMCIZ/G+WNKWCfRnkHWKRf47K+ru+TKofopUPROWYfeN1E7A9Cv
nsr9+ANZ4rDT5HAIxNt/jlZLzOozt/E4uoDn29P0KdcJXFe46JonrC++abAwtT4b
nA6K/Dia4H2XegqYIkOX/npF8m451hh9lARBA5zwBWTF4Vs//X0IY27eoEEGfuUY
VJqk3mjfHdPc2jwNttTDlBsimGiOa+fRIIjV/J6Pklm0l1OkV7NlL08hgq9w5sS+
kcSmSGBQNRk4xU//2IaaEJk3fz3m52kyJRzzBtkUYCWr5oryVMDcOdaph2RyPJvx
ywlfycPs+ifa0BEQUbZ/AlsaZ8BpBY9R4gsrurSOkO0810pGa1lZvHupDrviOnwr
vUOzwNMRuIP2xQJAr7S83eRdiUAGM0tViqeKP9bovI8nVC4zLN/ooXSh50yx2K0A
t4boXWva8+BSunu/W0zMioEKwEncUsdupXQcoB27Si77qPV160sjq4/Lc/4LTrUl
NXPaggdKgoJNoF6qBNze8coVb9P7DDyNqyVuBczG7E7oob0NCF5I1lLspTRY8onS
WUKpQvf1caNzQs6YLeZloHYt3VQGAlnPG6+hZ2hGGulyFl/UZn6sbsmSVp3VW0r1
UqXzncyKBJfRY+eIE/gFY254iCci9ym/5M6eCWuMbE/5J1IrzO31xdwV5MzNRmvP
YMwA0pcopYQS18DTBgtjO3BhC6DQ4EhSOSm5KsDNkw5lcEmqRZhYWprRvAY3ajzv
dvjiLCVz3xFsBZ0plakL7UUThFSiOcex4XD8yEpUevaguDHypwm/JyrJVRzGtkx4
3W0P6YlJGVR57CCzwML8M1NcJIkUgqqFNT8XEonA7MXH2vvjSfh9Lb0tdW3/XDYt
sDnc4Kk668FaSfYMcQHrlmzJrrSbvYhcByr0udEXyIevZGXH9c5KaU1PpNclYo2M
Acq8VsEQmlp5KMG5+b3yWsEzPYReZoriqZvLcJZs3ZLXcMibU72BO83zKDJYraF0
uxG8U8AKvn/12C66bcRhh8PcrPRQDuuNOZ7ENO7j1WkYub57NRkC5XcnNIXPpF5L
9PxRgrIn3BsyOyIWrHfQmaRJXvgFJXM0RwPhWdh/URSqX7PxM6OJDIvkOUeoxUlZ
E5jdVeO4IUWvSmXIjPGLbFwexXp+VXc6raxxYTurUfLsrz3Ejbk7uncb4rfaV+tj
xaNWEivS+4T2UgBlkefI1+ZzYQzviHIFafuFRryXj/37f7lCaeCRsCmdDNbxaKtx
uKQEgruMSSlr6yo+sodr/dxvCi/LCwE6GcWBJA3bfBdD6GEQXfEnWafs/itbRRUF
WaiY9pSuRlZ/3Ochy1T3bfhusUsL+fYdcFQS4cbx6KqoY530QzNUVThL/Xyroslm
RRU9058nPHmGGiPXZML3g2cWSQETF+zMRZ5Fy9wa31mQEblix4XQTQh9QViwewKY
YbyLarHtid5YfCRhNw+D5h/Ov84bc7Vuzx0ac9XzkriD9lLZF53sbwVoYJOzD0CD
GtB5ewj3h0fl0mjI4A+fYgEKKYEV3QvNj0uE+UPCi5T8X9mNq4pXO5rF79RSg4WQ
5N7E2ylEPzgW7qNugqpyw2EXSErrUT9GfW1E3KiiMN7RmtM3IbQyZg5EpKyYDQVc
VAzIAZWAI6jtdz3KpG5aVjbdVLZ55M/9Ga1Rlc6zpZYEq8E4mD33rt79AnAYLzb9
QgzwBy89HIbHw3GguHyVhBNXJotxREJ5O7FWq9bf1cPsChCfW/kpW10C5SdwJz3N
d32g/QST7RehDFPnwgvECFTmTfyGE7XS9UQiha088+hGolCX43m6GEEy+DlmF3LX
Q9bvlddJHLLniVitSiLxJC9jscVKkBOcD1AuyNU7Y3IY5KnHht5ifFXFq/LeH2Qs
sni+AdHhC8hTVHXAJWVSi6V4d2jpYuOdHF/p5IP39FsaYeD5mQysv+7Tgg3kdC68
SgP8JKMx62Ct0ZE1H4Ptu0Xkvp7f1j7qsGc+7awi9PkZi6R9ynu86MlVeKwdp4UX
1lE1okYuqu5rhd8LXfszMsr2ue1ir23sKy/s8EBN0q7rwHXtliahxUz9fKcBguMb
wdBNk3S1/xslMSARlIl1ghdMo6CPKxfD2XTARo98FzaUdARA8SmvIUwxdaTavjFP
VHTO4BfeCMxnffPcJGyOgYsJuWOu5QqSTAtKobLwWZSbb/LjUv/xOAn1afxWu3Dg
XGi4CEuCieKKEwVNwXXrqKGOamHoJET9GYmEven+EJ/rCFW1lKuYt0vk5AW09R26
KHNlxFOkQ95mQc+ArlLJz29jtq/3KH+oS+YYxoU8xPaiHx+BmWwRKMerjU2DxnrO
crDYRjNhXI7QooYdRVBNM4yKcqKG7Aq7m8TNmLT6CoOrmo3qvtC/Bi1jkj79yw+E
z/yxJcXJ2lHq/GcaNkpIRNiUyLKy6f/XihnFaM1VuVq3kNVT83U7vD2+ZzapM34l
RzRw5VClaCpbQE3TLwvpJ0w5Ogk4dUnE15/4gZjCuC+BKGQvEC03VtyTk+P76ir7
s5EDshMTt/z2jZZP1nHTFgon2TGnEN4RRDwy7NqQfGKmwULZb2bHBCLWV+5ybow/
fIQkR+OBBCryxwYXsRBX4OUARgjFO/LgT4P3RcoHJnIrlB8jJAwch+5LU/NpjklX
mgCKRNQQywjcazOGABgilKxLwKc2T2bVGGEv5afem+NPvu5ed/aF6DXtiNyLaqrb
NIcypiSzZymDYw0qs4Wd+l1tG3sKVOFCJzIjXecr0rI+GSa9i+wUWpcdSQzLliKi
Zn76vg5JaSquc0atlD8V6W8bcvs8KwtW9x/gu2Hm1rrio63pKkmrp38NBPAy4Y0Y
ucYWI7VUoTdN7huc/9lUo8hFOO25sMVFH7vqohyfkHu3xLv3hMFDRy1Wu0CUm7ar
g7SKhU21GgimC3hOfR1pt0/qJoz9A/mffYfRPScRgEaV4VBHDEL0Fqa2uGqXvzZF
Yi1iOE7ULjVg9109EnOxUIb1sP4Ws8Ohjcrph0FG4W2mhKoWLIbGZOs00hKIuWe4
Cse11vtQQ+YCY+VEYrE68aixLaWDPWNx+UKWM4apbk87QZ2uXOXmG3q2XQpqpeKv
iLlzOaKPgu/Zckrxrr0V0o25Xm3H1A/nODyHGgcaRckrBJgAyVoSUMdjB9ozZDL7
kslg4qMzs38C5e8fiVHAtTiMg7hw8bN7TLjIr7ZLvq6sOISUpT9QY37J0Kbqfdc3
b7iFh6xTsYLNMaWBnC5fJubmeHE40hnkPXUC1XqZqIHbeXzvgaaz43c2B2kcGBuM
IfE2R32iP/KG7IJxY/EgClR+55Kt5NzerzJ6vyu7gsea1io0C2hWIG0ywY2Y8KLj
`protect END_PROTECTED
