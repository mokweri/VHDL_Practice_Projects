`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LlVQvFl+MmfO++b1VR9SAuIRUqKwXQyhN2ZDsJkplzvxXptDZ42TgzD2rZlymJ0H
5cA4tLmc0w0qyBKiTAOvMnoK6Qabrb97aQ7TYStVuS/8L2Bfy3rT5f1e8pmeFhgO
46KLJD5z/V2UxnyNGMb+Ep9HlHPaDmWtR7foHys+cwkOnVZgSn2oYqzgqPsgzLLf
13J9mWSLfTxVzEPu7U9HhYGLSqQBMSgUvAFSxs7yEmV/KTFemq3+VRFwzVkUeXQm
I477WKSgePYNoyzTP/UL+ljHbiQ6jLZ2yYN1+v2HsUYexkmn0hXSk8D7yO6rYZKP
EBZQtADZ/9wDtFf/HAa+7+cIymHdAw5WjKo6pHgjE/7v4IYPIlbjto91rseYVYJi
O4F5/EH93OH/I3dnqiCtrHYwKyq2spqel8/503mDy15yQl/EPcfsePAl/HyOGE3d
uhJmvtyoNhqPfhsXO4a65uRuPCxX2qgOgkTBs1p61XlIhojo5emSLOaM4MtdxC4y
RFfC9fDn9pqeiKGVEZOM0fAZxJ4OXppVLCr/D1TErTdL3cupdvD9R00Ym/lh93TD
2i1dR1l7VIsC0/WlPNA+Jxj2GM94Y1927pvPGNjJsivd44Flkn5Z7ljpbsO2Fh42
ACJx3mfsHBUf2uRWs9o+tyIrhCXZDK+692AS91r6IF+ulw9tSXNblWMDyqqjOokY
RJa90MZoYfp/vpTHzlThXLTpYK/RRwUHTUhFxNXZdjb4lTZn0bnfVp27Pwihwz09
96R9zZJaurna6IiDk9+zAGtLVuy78FUjyT8j3m0TDyz3TahRRqUiqvaI2LDnurvw
0PpFrhPk4TlaK3arL66O+QTN52w4++X6OixMabnvAagHAMD39Hce+oP8O/qyB1Mx
c4k+fFstuj4nLAhedioVD3SBmZu6YRSwR2mH/WVK0nwr/ylaCeXT1V60VGo/8ScX
SRcZm8DH1pfvclCllJnxy0TWv8m/QDhCgZxp2zenx9oJ0kHO4Jbt+kxrGotBv99i
r1c3D5M/MRimuxVqeGjSZ3SoD2DL47SqhAYJldf9789APwyeZJwqnu6U404v+OoJ
Etsg76qag56cQePqw5h8gYngEjZotOVccWnI9HdUcGm3CjMM+pldVaS6O1WiJY1c
1on9+PX9dPx9qV2D4unwavLnrJFcYLfaUOhj7q6Am+EQA3pDnGIraROn2ENP48Mr
AYeO0MmOzVI4MRH4ojxInxRovrpJSmzFUHkp/CvIeCRdyjNmsACKayojRl9qLFWd
WiLW8WykVALtB+c9zzbhSFhffPNJP5jrL5HNfduLYrTYvuaxgADfvsP9d6YQV3AH
sqeBCANH/wCwYbwCinzIrXkVIVEFQsyELRL/dL7BVhV58a5lY6FuuIxMpNWaxjZw
EpiYa41uT6EwCyuv4MAkpKYbUY4zj9MgtJkExvMawJPO0LpngKI7UmbAiVjCzDVR
CgbLrGBTRhXpHfU6onkdiqANbUjFlcG9TISwvbC4X2A00+bEH2njjSW0uRZfCqOQ
QixYeuzD2ydVuEyAH2KnwubMq1OTqKfPbZNqhM7QxVKAbOc8VKJqwMEbe+STwF2b
XuFY3Im9IIpEd7grlBINFhWu9WcNglJV9L7XyaRo+LaZSM4EUqYEq49y0sumQ70D
yLkg6uB71XXX/pla4RAF6wZ/SjmherjyRRDAFlTJ+fyL9kw1KA3y1lTyX0lUlVuM
AofpkLJHZZpunjq06fO1EDN4+IaLwehbsErMMIzhf2kk7dqUx3Qj3UEAUa7/24tA
McThBjugL5u4CnDlIhVc47Aocu8F1xyTrUSRVp0lJ7r28lAmbOqpWJAhL8gXKPMW
dz1Ut6ZJJEM8hw/Mp5NiwyHxpwqp3NmmVmRHCrHRCa+hgm7httCezNfWIwH16nc5
L+SoLTknWGkLjwUlQd9ZtY4xXMTQrYo+273yTplBuIvxUTP7aam1j4lKl6RuBJRc
eYz/P1S4puW6upTtACgrQQ2h6eFV5Ywwn44boVMUcP1vCUwpnSVlyF7AWAkxHM+w
eRrWtPQQjnhgkS+CH+DQol4ht4LnjOBiBFPd/fHq7y4E+irRnvjR0FMWeuvQUkAF
q8mPa8xOINyA2sGiBkPkO62qWJgcZDZ6Vb+AJlPlb+bgttgmTX3Q0TPOmv8+dNc+
jecsi9VwGZlBTq+r+vTCqOYZbrXLaQE/gTXp0f4bSDt67cvc8pDJimVfkJBetbdH
ar1JGuk9rzkCW3V6PGyzctwVattE0aWqoo7b3yvG6QFsSzzKkWiov9ANbN0Peqrd
wjUOFuFY/4sYRprsps+8XTii717WYx+hhjZqmYseF91wQiQVl0KMoT8pit9FZ1OG
fdwppzoZWyzMnr6qOxXfICe9o2mM0rw4uFAZkLc3XUbKPoepZGOMHDQ7VP42rDOO
APoHyPZIn4G4VomdhfZqx7Gh5WAJLuZ2NkwWZCtGpNYDCHsQZ0UesOiluqS4hXh1
onHfy0Poz1RxLgBa8Dn72hj0Y5BwCT5yti3arncxKCUOvHaE4GCmspdi4wbVCwON
L22vQiwBQ58xtIrRmO087WpzFGYWqLoPRcLl2+aO4MinPAxKbgOAqodFBsHzp8zz
jf7mbv+fhgfl7wxLz9XzHHpQpgkFr5F5PbHs//dRJ7SVUu+fxR6WfBUnwZnlEVhs
TYFpL20g71rezfRs/KyJ+qze12Pj7MaS8uOd74DXUQaBKCcuwSqLnCxkpvTB/wns
EFGSDrRYrWjQd6cs/mdQIr7tJAM35NgstsE9rXi49Dee8/+zlXNv1+qMRKu0yl6s
pLwMpgRF1vcKbblrmikS+PP1wJS3sMpP3wEoZiPItwI=
`protect END_PROTECTED
