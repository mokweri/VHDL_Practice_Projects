`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmT5CS69wkmhuT0Swl3AVfRqHNwibO284B5Hi4uhMIhDvUQjYtaesAK3IukdDsbf
KJj+gNHiD9XwMrrJf9c2VFMzM/65QcMQlltlhpdEeJvpfYkebYAaxk9WFYuD6Fj2
GA+Hfqfn7fE46r5PNADmT3+kkHNKJaUipoqax5gUyiw/cYaGJ4qmmnT/w7zGF8rx
LkSk4nUWXzd+pDvAwqIMHpobvoVvALV9eYHEWZ2sMTjyh96F41/qWZqXMtG+qCKW
O4zC0naryWQdqIriIhgcYJ54rOGY3KyYOwcSE+ZF+Gvh0T+i0p+aRj8xMt5gaqAh
HsjzcfqdY+rQa913HJDvWsu6DzhHr7q3Upa5F3nYLaigvmZ9w0VxlN3mi1GanQqM
vnUDXnx3fpz/QTv1hChF4rh5hrYV//2UUvUNZt0aMOJdkBHTANpp8OKPr8N37wyh
hVE6DoM+vHpwvLHb5JAIN6O2eWNnXU/Nt5zoBwixir8=
`protect END_PROTECTED
