`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OV/TjV6aDNTuaQ+TmXxqPyKXqZQIiE3nERiWZDpxJXj/T+w9+YIQVV1FkpoL1ogQ
4CrxJ+VK/0eAk2mikADyJGOj5VGakIgzlEdBje2Lyf/l7UUJkRB/zCNkLS5wzybu
JjpPefzgc/uLgJ/HpwDuxo9igWfzWzcyvvpOD5REBELfqPWNCajb1PBRHT/Vk63I
OXoiMeK9EbTtuf6rWvKN3tRjPdPvElEZ/6G9PHQYb+hcjhcNkpoez/P3HldAgBh5
ZBqcM5DKg1L2myMq+WRAw9FiHN48B2O73Hb0LEYMlLhHPYBWdtfG1RuuHxDiSFWi
bxiod/u1HkgP/ZCP8YqXs1My5XKt/1Py8Fotxax5les/B6L6NKKH8cPHqh/6vrNh
A8Z/pVb1aEGErkAGR66XoRVDuXTo4y1kqC6l7tklMP5ZEnxaqpZ0wMcqrSlo5LgE
fCZGXEQ3Isfw+Aek4SbGI9uvhv5si+QCFF3PCZ3tngbubCX7LQQc567Bu6XAG2J0
V+2nhnRE4OoQEHmJdLjAjzIgygReX/4Xizplx5vY3DUyNbewbCmufVKXiEZwtFvK
KZ6usJXbSovVdDuqrgwIhTPuMXshDpU4VL+0c8zFzKBWj5JYeLCIxATeHxJ8NOHf
kUoDR/8yhnxm3k/cNc6IlUV0VT3x/nDlHeuojOrT58Wnsb1WnPsRVMt4icd0NCkz
FcA6NPHcNycCCK2Ra6Z59k4ZSdX6QO+3vKVnQ/yI0YvEUOJWdlKjCrSBZGLEYisX
TeJrpJGdvzkpSnt4NCIXRx1lZgwb4YpFwUUnLsAKhq3g4AH/lCnjNX9hsZkBEnNk
vkuWD7lW6DFfPfP9kR70uTb8Kd2nd74H5GuHUjYU7nypmsQnnMHt4hoy1CgbG3TR
cjDOdMEfyI/n+OQ2N8CiqKJ7Oa4NzW83XvDEwCcUcpC+wcUSYZQVbbb787wbZQE/
Dp8JjmFtcNOxkSDJpIziyhsqKJCXeyM5bzzHMFmQxVHDNNKBtt7gQGbsZozV6GFu
qVis9NMquhDtVbJ1PYD5neRGy1oZbxsQehVu6UiLmysENq+xkJXexQPCiSKSVTGj
xce2DvrGzuzV4eQzRmHXrvc74Pwj7lCffOCbUzARnjGK6k8nY3sEyXeeG3YmkGpn
gH9PAHhoGDQ6itmQHCEkC6wtmXoHEzkWfWPgnlmV/z7UAwtgdJXHfZM0C7FlJko6
u8BwcxIiRQZEMRul9NDtHxNfM0nislRsDdgGjVhQeROuIkaixoMpY2n6kSQ3UJcb
/nYdTA1/hCUqMoJPTmxgQVB1XJ1jughZdmDZL8S2Zn8czvPn4NXlqiWhyJjFWtzp
odSEttUiQOzMnhNWTto77T4lzVD+h7E5vvDVdF0I1ghwkMURH9I7gpczR7dM8RcF
Ivr5W5A2+OIA1Ar08jWE1hWvaXYR9WA+WYhh/lk3i7OiMfBEdAQftuGC/JHoa0EZ
Fat98/vb8Fc+0+JeD2HlFw==
`protect END_PROTECTED
