`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQvnNZ0oUW4MD9Jt/YlbH0QqG0VGToQQ8AprOtsLdyZU/kfEC5PnR4D0RbNuU3VJ
pxSsHHVZsEMM4I7gTM2UULFue7CgIpNmvMyGvJ50C757Ru7CTkwlECnOJw92gHmG
LwjvxF3DL/MPOFpGalC+2w9RsY5lk4ZJT+v2zyF4JAPaDWWNf3EzCeArb6i3hkmC
nFPW8jeuQVmBACPsXA24J2dx8nPQ2FT+eWMzrl6XZMWT8QF8VdOjgAjpW8bWJuYI
6abxY96OEDstZ7U4OQnP2qqRscvMaumLZ4RYQOVj3h1c67XMLGqoEt30AwZEtMd7
vrh0qjjfORpp80JplNyvYR96KfxTsRIXFk8KFCBEEVD6os7eux0BPqNgvgFU8ay1
Qj0F/aaQ+ASV3lH3ezTVj3cscHPnRfsmshCZ1idnm5PloxTibtA4E0sk+Pj1O4fV
RRhNnvosfDMQuD3UdHSLE/ybl9b+gd8vvs9R4BpwM/o=
`protect END_PROTECTED
