`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
edHop/3TayMmgnFeLjZYivAkxpJ/KeaWdRpK9pt42IcQ59SOljaBQ2MrrNPuFNjY
qK/Oi9nFHLWX6bgDnWYdl7Ahe5lzjp7VsuZNoRmjTxKPXXQtdjAndfRPcPxhA3Uq
0XtKBWGqhx5C9o21LSKp2mshCGyRoDHGyRzNLVp8xzZ4g2mXvSrIffeYiohB5Njj
ZCYoSbysB9Wj7VHDhCKL9r/TcI/o8vTiSprA34BjsdJ8n+KAWkZp3LBk8DUQJ7Th
P4D9K/lsAss5RMJtujIVX+Lc16q6BPFNagOE0/2//jVuPGmxESa3ESdJLFHi3yKx
VJJBi7lOd+ZNP7JddRYvOSI8Ve8QQlQoT7jbSms20ene0NjNjkohuibMEc9qL2LF
`protect END_PROTECTED
