`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
olB/FPwKm/XFI7kmTrjiMATZrDnBpcRZ97TugXqjL9x8CVpT/5PI4EWalxQ/1TVK
X3l4AGtv96GyCF1nAtIlJfZsv53gaVm8VdB5VUHHyuoHtLdvMznz1+Ygh9lmN+qm
0G8b8XLYArHyQlXnlRIoNoPyXuQ8yJNRnscXhhY5ZlhJibYEIhieqscSXzhbGwrh
TZOYisuqfLJYjY3R2Rd0FTkiM1SdLvDANfwHSMeCx52Nu2QnyUoHs10mL5kViesk
gnqyCEVThZRKFSGNWjwBP5fo7pijj4omLDeKhhfeMehMWjfF9UYiprIVoFAvCmxD
QJtFjw3hmJ7TVrfn27IxPreqFfjuzivFXG8Dmh9D4U6hclTAJYOIDcNy4eUyiJPj
e72uHc0jspBMLsStAPOGphg87WfGYeveWKJjDhIuFJlfaxp9KPkc2IUHU5ATe6Sq
aQJp4WG0mRhrPUJj8y/oPK4+V8qIu0UIrDfdMGraCoTs+f70jL0ZGCfuKWrrDhyy
vUaoWTjVfWInvOkqLFfjuXBUA2DldMicUvn2hChjm+0DDpNDy+mz6ZGz2edD7D3j
LN5jNX1dTkCMRjXkClhjf1otGFnrrGsMnZppAN9ON7Hhfvu4m0+lGlP4fJHSE+Lj
BGQLNkifyJVbqZBUS8xDJb9B4/1eCnFKgWEFG0BXFPEXesMCaG8zW2NXZw6n/Od1
8FFwhyTKsfmH1zBbrg4Mk+D/qYiiL93DmhL2U6ywi686nKWnxU8yJlqIPu+f1Smj
26OIxW1jPE+YE/hCYRK4FHR26uDz3NaIHnGzul1wGZkbK2kE7euN/Z5t96CMBLHk
JyygQkccPkqrvKSf7jW3sjoROhIa48v+kYmieg6ICCeBVZT89DkF4Nv8O7Pbg0Q6
3M5+iijTKNAuA6gyUPAhtkAC6aQBN11zAtffEU5pI6MXfhDnXjZg5/DhH+0v6jnd
BQSGOYg7Vrsp+xO/hRqCBKysTwaIBgl+zdR5ZUnHfhM6HYjBXk9mObaN6/3SsUH9
Sfcsp5Vh4zELnGcpEOAEjqjozfeMqWDCY30Bxd/wPMqp1+VOrjjMjXAPUPM7Jk2h
FvLrKOO0/1DkaTPKJ/FdBvGBacJKJpKMKzqAWZMk9MtYbgashglHP93PCZwHZkSc
KGl+iXDRMhQJ5ZOudJM85J+j7fxrFo/sHljp9vq3AFDDUKFc3iztEqC/duT5XgWV
HTHYgXtG4/OvVS+Rg2tCLhSIiNvoPvtyvBd/PkUYoPpWhkE8UKOF6ftjXbBo7suT
6hHCgRDBYuM/CpJH+6fLhjSjKQdHVKbsOQKjVnDYPNNBkmSbbW3Osv30lHNzioaR
8jzpNsHPLU6SL+qp8zCNKuVq1Y14JHCPF0B7WY+bXqPV3JzRt14XzALBU+Q+5af6
Gs4buSzid14yoaStSQeFpLxyvZO8GIMJ/PwWUtsADgxsFYSspkcoto31RYW0z2CA
TbMsCEzHY7P/kNaQ2kC5/eTaUeEOBhIe8j9aVx+TYbYldMnVnpNphjGqQ9Qh/jYp
KrUUWUFWAtRD7RGFfI8y7eQMikrBrrPLHYjVC9jCw6mMFWu0Nu8PLkFdoBoPSq7/
VzBi4Jzg1L0MNk9Od6E1F1WOdLKbfmKgdRg4ivaTUNXA3QmCFHArsyTFF2e03Gkd
Zkx0Dc7e7hoLS5152/1YHlwHnc540lhmuZlgnRxq5LPOaYNEVPNrNd3ERo7G6U44
P0MlMsGeipRo6RLKflb6kA7+BFgUYfZRYyMw5VPn4a+izuhIVvNztuGoaCpzNExI
ju44ZL2vsVHC6rIu4pu3vu12UCxBT6UYt+b91FO6/YuWapZ0wdA0uwbwcsthaexu
jCwS/z+SJyLBXPwHz8xd6mf+Fu3EYlLRZn+92NScI2iIMA7XLfXeT5ZRCSC2P2So
X9J+Cuhucc3YucJYXgrtg+FKTBGNwIQUEhfvQ09/ogMWfucCz+M2FWl4eBVNY0K6
8sAvcj0GUrFA2JWvgySjlmdG0lhayXarpINEYoUeccBTMpC++Jwt2n4R0iLKID0I
MPLlnrm365W+LEPEVY4YFkMcJQPsag1+pbbnZyp1mS4vyvRRVZXX0xpLNTLcUowA
PapXfGzIDlvG/h8FHYDCM8wvY6g/QkfXCF5JFlonj9S0U2+D3ML3zWa+2/pmAAiS
8xNdDI6yjgJFb495FQMkDGf9lJimeiBmZKpGYYylhHshsX7R9dn99xmTI0mkXDHE
fUijCwJRuJO3IL6wFf6QfliUJ+sU6P/LhQKGsSAQIUVkrtAu//kzgP1pSbfzcjrp
7VjnVGA/6ksFJu8wH1p9nC41vVxVI009K4oMKUMpGSq7wj88prlJ3di+wDfLsXQQ
B8DX9sttN2p98zD0UuSNpQ==
`protect END_PROTECTED
