`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wI5sT4ia241uocwmhun4PRpH/VskUjRRqVJcl3X65B0TDPA/XbVXGQP9leX0ZW4b
joYio2hX+eWK3mCwc3srKcslqF20RXZvDcOEyYqEPojQ72mJluCkUKD/qlkqgzCx
bxVavdOMwMcXEvdnmcNiFpdb/DIGjUNMuKvm+GNDjjOpC5ni2iGdSHaVElJmWGrl
ekk4XzB3GXMXD6rff3PJmynD76i2pgf/VLQva6cw/ozK5/Dc50GdRAMHWUT1wFyJ
1tinb4bgAdUg1Op619rd0gtvQ2yOgoXKZoQsdDw9WQZqj9HlqbBjZqLubw8Tc522
Q42OAvQW7rAp/0PK/e3HjMvCafBVklu3srglbXrTzCXKNaDz9YRpY0es6MjUAawB
yTVYd47TH/SvJk9agBnpoxeJaIohYCQ6jLUxJXi3uMVzXAVYxYLnpHHr2UthcIzd
WWE5zIq0A5MIYxlFujVu7lX8MZQgSPXrrebztgyjpwnN3EW8+qXARdyzOUoUXLFG
vhurSRQ5gokw6TDzD0Zn73MCPvC9uJ5R4Au7VaMtrXADTf4hoXEsB/zMi0Knas9Y
FtRrcTbaWygX61xoxnvuq5zc9magc2BLq2OCBtgipAwWWa3Btvz5JoZasHwT13Ei
KL+RmxMxlTyoBYDZ5oRs2EQuJM4UCXPOHCxhGSPP8H3+Kci9wBGyx+mgKhmTVyVP
/B4afy+O0GvlsojHZByI5tKnMkhjjztKIumrfRLc9ptiEvpmiHZy7PjS3Vja4h5K
iD3AuA4QU7ryYIih4aAAToWG4OqVCdPaStVPOfcPNYhzLYVCuwPQ7ApsJyxYR6nl
pZQnD+ygEQGzc1vSNyPFR9b42aASHSlnUyJ8f/35cgJ+w7v6D7fIO5DSBGNEjK5t
k7a15vMde8h19q7ZAVf6aOO42OQNUgQtGBCiNfHPzEe6jPI+VylAPr2Yps4fwkFC
34f1JyFivFmExPE+/5KM5xDGUCWt1Etzxv+Nc58h/R0q5WYwFcsbRHRv9gJM/bFy
WYwVIoBGTK7AbUSOoQD6EhsQLYpOASFv4pUgMPE5lIAAkK2H4/FZJbsafq6G4wzl
hQa+DrwikCM7jW01QPOhPPzfCWbR5VUbv+RLAA1Ous7yE7Aq3S7qzpfUj9kFtr0j
nyDdJbWq2H0DHmN9hfQkyVACZPeabF/yZho1cJ8tOOwCacrR9zaJAQs8v7cl9DX8
FDLVkurYRjCadamJIybBl0F6RtXcestUp4wmUmPzExvh7rOTImhgFm5+VcJa8Htd
oNdoGN0OYsShh6NpY5yYGOkjURSUYUGpUnfLgmP+ZWFffyc6Qfd4UJM3YpxqBRRG
PDCBMfLXx0TsfYHFzAUfk068giv8BLY+MPQOp8ruQQNJBEDWfle1jmlXxZ9a5GsA
RQZcThbZCTkLGJ9otYHov2sMVtI8pCBCC7BK7zRVjtKWitV+WsvIq+NpQdRtuUI9
YnR+Te+H8Dnf2bxEob1rrc5YJ/QRVx7p1XYuc5a+DXvyO5ciJpER8OB/bJpW8NlH
NYOieCYiWb9JiOdlnfhQ7BVhgntDX5XX0QIxghvjqZQy0l5umx1tO+lIIRLrHuR1
/AweGAmow9yKK1d85PBOgTBXfpEXDvC6qm5bjdjpG0M0KLAmRUCQ89UHv4OKwcN7
wC9km4DXFDOooH7Nkd7p3h1w3hNwr/IMDXoZigNpPw2WT7N1y/4xy/u2k5/C4QKZ
Oo3X/55DSScSWK6NAbPYRJwhXAiFto56kDYg2CvwKDsHpW3wsd4J0T7gZ28+A0Pm
33mUVA+v0cnrDmpCaTMv8YiKgDHzESuxgPfLOVjt2rzE3kUiSOI3Eo/ZiMQuYvTo
SrB2VmsGkfyWfXj6DgNzMSSzgfhBMMPezZYTfE7XLHUTmw99lhCDKB/6sFQUw0WM
JB/SHw6Tg9MOrg8Q0gew+3vafsr1e92xTvA9fm/amEuCCUy7FUQcoFfalj0FxFZZ
0LaEEjDOx+AfvciH/u+gCwMR/aqAQ9gkOpSbmD/qwiAGtZ+H8ZdVKx6pmv9X+YQ2
2VXaBZMjZMvZor9k5WqjBU6NII6Q+9X39W1ciOOgStSF1pgMDUBmfXgYLicHWo/V
mMC9m3K9eUuhxv2kQSxjiLMXUjMgwtr5GBHCaFPT0fMgBLFMA60SzzU6DUMK5FBW
4ufPiFTr3Ma1L8g6Q5f1ttla1dSGfMoLCeZ26Ce1m5p8DQgpX+07Bao0VQU+vj5Q
NuxkUkxYwTfAPkI19KjeBlqztEsN79gmbjZP1KhDvjmOJyH0d6JTmWLoGjy0YY4j
7gKp5epZ0ejcg9LIWX5wEnZyPnXc3lb2Iq552eEdhAtuci39BRBvjqS+FxGu7zaL
C/7VVSO4hyJVDPDYNv0D97DIPR9gMX5Pn3Y66te4lV0eF3YkecD7zMny1ZoRN4Gf
CYmIIEseB0IHYidxTnjEFT8DJL75bf4qzZmwvjqim4CKah3t8U0239uT4dmi1TIY
5wlnFIRHZwNKDc2IkosNfGvv2DJ+NfXH65lbiCRq+t4FBYF1v1M7tZAI09E7v+k+
dHdInMcpnS7fXdRLwVnN3l7CGi7uBOkI4L6r+dhbulQUJE/iQHUCfACIjk3wcSEB
M8EOA9bFYvWmff0jdrLFe78cVJJCwEO95HdAlmcFDFk=
`protect END_PROTECTED
