`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMKJmbPGaE9MipoklvusDcu1batWNGplvB8/p8zIoM5vw46IMC54+nVAjBfcJaK2
z0wa9kgJU78padJLwC8DkLDcjFGHcZaqdOZlVxf7o16qnjSRBIu5lWZCIAzc/RuO
wqHScuoECgwDV2Z08hIlWYB9MhSO+M+OfHbzvHWAh/QVnpjymCWHsjgBBDrtbY9p
IBYA0sW18OeZfxsWZoEBNFxmDIUE8QQ4EBefN9AGfXQXVAWMYCzJKT0GAc+pTyZj
hrylMx0pWYYZcosLdwSOMo0xmmvzYrflOGZmj4qLdBTJ6dpo/MoBH1E40ybey5PH
VE8v3PFLdq9DkR/wBrfi/9BnXohzVb7RnuOL6F8vLGhVV6I5hmcPGuVLZ7d/IMIN
/S+kHxzdGtSS/srwrzeGbtsdDMWniFEZ+wFehLXVTgsbWmXZFq8I7dJAFJbvisyy
9GD0drCKhuvAn4RelMW1fH+gVSo2GimuzbY92qpIFWlzSVi5KVS04uNBoGJmHJNx
QCbnzONaA0HxsZb74bKxrsW55DrPTuIWDpVsfUu5qjkesNNSAEGzNsxjpQpdYSnp
BNJzrqPUqsvby5MxS0iwAuprh2txhOOs+aUKEQ3CKdZ6D7H91wvuh6LfmOFC3i09
bKtD7+kIReGbyfWnCxPl4CY6RYa8cFaYL81zt/DMSPbYcU6MT/mJlh+BqB5hVRgQ
`protect END_PROTECTED
