`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwNdZ1Qy+oKsKUshPCxU6k/26N4Sh71AC/qvmDVo6sEU0YoGjdDaoWKgEBipwbCm
pQAykK2AOnntjnm3IU97nviSqz0OD/nkq3qIlNSrayn4UIbdPS0os9EhdjmT87ND
blSWca0qHOMsV+Ko307hunUC9xmAlpimL4KLRdZ56HlSEw7Oe57HSbbYqY6eWeyu
H6kKDvN6urWNSHSBH+kk7hc6/SMpk43PEjmb9b36NhFmLPl85vCi6Z8FI0Bm0wUG
21al+FJt3fAPDPsUpRqTJKlnJGB0gr4+f/ACuM4LNp1M3iVsu9JbTR2OqrFvuxSq
fgqf/ltEzV4dyhu2CJ5zIvoN6NZ30He0N1UJYjhweYhHAYqaEaRsMv0P5/R++nqK
TYCPdELN8WMwtwv6TjBOlT3VGC81+ytfmCs0XtOMgR1x72d3d1WPd4GIkj18Nw0V
Nd8kXEhbmpRHq19CXIreZnTMeSaQ7p1Dr02bZo4gaLQ4fWOa6pbfSK9inX6/xJOE
b5X3Wk3XAtM8L1Le6zVH/ovDqIBqxIZfgE0Zbs1nTxSVdX0wVR4WxNG2EYMrPMvC
D3YeYsnFowBqw/ZgghaZNXvTwCVO868EU/+KqQmmWZJcgC7I1hpnunWCBHirOo6i
Zog0XuiAIHvZGIZ6uAbxAPt5cQiFzijM44OxGx5WbNrEVkdiYkG4e7EQN0n8b9Is
PoRl/i13aeYGk3uT0pa/wQeUHnz8iHntiluaMtKyeG1DQFmYekqbcAoJPMzvCeeW
sLn5noTCeeXaJi3uO/pXED9lo377ozY3yuQFpseWNWrmlhxYQSpHe8PdTXAIs1nf
nhfwo6uQgBR+oJ0u2TBhnjwk6Tqkn6l5wAZD+4HKEvyzGUI6/T6baaq/PjTWggdH
qOO9+mV7A0u1ShmR/B62u4JQTUIKXiQ7B02Ai0IViHFvA8Xc3v0H0Esk+vd5Bbiu
MKdk9QRVgIMoDro2HnihIyJhXdyrVYxDCWXaKoYCOgJIwOrCysp9iGMXQiVIPBzB
1tdiTECPx6afvV2ks9kRQOTKH1O3Qd1dUgztbmaB8vabzGGRtFUjRR6IV8Rjs16M
`protect END_PROTECTED
