`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFqNmSZ9/Tnn3JokypepIVTjtEDqQSgy+NY0ldW7bgK19GA+gJqbMXKz/nUX99+n
elNOJW+OvC6qeeNPc+zcFgKuBGuBlqpsYy69ZFfdsJkjJoNur0zZ5/oqdA6BUan2
b2vXYd9YLCqBW/274fTtr3hLDphePC8JIP6CnM0bEIfNxCtTUWFDmjqYD92Tfy+z
bSHAaeOq2A+OB+ed1FpPh3rwIl0Y9dS1yAWcJOKkO1H96q5mHFBjzBfTdw0iw17u
gIf7naAdBb0vbEN20POMGVnqdIfuHQ7yUOOc5iTuBMHvgScUMhi+eZfgHlfkO9kT
D43m0ffTLKXt7vTLWxKtGwwNiq5QPQP3Pp891d7m3SmQvifY+f3+SFyFXzK7/ZUK
VrrhyO/4xCrMVxMCnweaemc47IT4KwmueSA4JGfGbFjE31RSFgaXEs0hV+CAXAuh
JjwVSw7FMJjVtf0/cd5hvoG8kPAdBtiTthrDo9c7IP4M/tyKKAB87qemLlH9Ln+h
bqbqgHZ2NauWjU4JABcmvF6j1LCKFX3A7QhB0kBVHK5ppiNFnHm0T924p7NmIVuq
DluDV08ykpR4pjJ+L6Z8gZfrX42Gj9Ibnp8nIzDYCJjuvd55LK0sA5pUVGYbOvg0
TlLRqObHxJ5Ac5Gp1D7t0gfru56TLd90ZNmCSOxsWv8C4uWSPw2F0lT9EGRe8nxo
jxc2LskFSj/vxWTa9YhwsqnxEShMBG8ahnSOXXlXOwHHvKrRud5dQBuymQRWuKj4
An8b2zEm9cLEpszjsAgJjLhl1t7MWwhfcZp6piU9POVdHq1kQofuut9Var24B7dY
U4KJn0swIqyFN+1ORs8L0oRh7UYSOSt/WFheRVntS5BbcGaFM3HzJIdapTfICqlM
8LT1NqgnzzriRQf7DCv8w7+jMbivGGbwp8jZNMOf26c1spEooFqmZ74Y8P7P/hvF
Q3Hvlm3oFcSODyKNb2S4Q9BHJfCmRiICOytiRPvfPqzmQxdsM7fx6v95LGb5XSir
EUMjJ035dVuGvwjs+SoEkMVDEaBToYKA2+1+WaF78H6XHVMGflqKUgQzueMQ6ZqU
72FGYMZh/E/PJURmhqxhsg==
`protect END_PROTECTED
