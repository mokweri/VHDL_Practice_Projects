`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETbpntVxVygGXclQAwr0kZ7IWtHLYqqIBqu1wguaB8A8UMP+2nFvtARxX9wCd2Sl
RTIwZraNnP4MW5vMK0H+yvN5xwidUb8kxgkmsIqYDGXLZe0IkChllIazA9Rx8E1Q
0S1TJhPELN5hO9PrIYWsTo9OF7S4QWfV5SnoXJTCao2aQbaHLiQo7h0VerbVigee
LYZK507GYYJ3I7KqFlCcDcUbGxSQwGKK9GG81FBX327H0Mw+5514D91LmRbExP/N
MOqCvsFkM5fYIKwG94iJlKjq48z08IazCM/s/u51pll0wVQivs8z9kqYdJskFiYO
egjneB4FdtBAqWHvdy8XVSMxON5f/BM++Z4pflpevtnb9T89widEd7isuXSYz1HW
mg4VwnD272kaCnQhPE211L/vygUH+nTwe5RkgPsT7Y3lcjo6obx2+BRcWxjxOFRk
to4G34sszChaPl+eDLUFFXPQSPfleQ6924vuu7i6prqCh9PwJp9mHmbJDiZwacWe
vahHgGjVtQ40lZlGRfXlKOFUZUnxoNO9yVrIJOO0Cu/mCXUIB2FPQAtSQYd/0+qU
DLRqa9Ywo2ixkv40jwGTqknUttjKuUB3y9zOxijSn5FrkFwZI/bl7tbNz3ln9BTa
2USdTUuXt+1Kh9efXjFKgcEwgKDTXNoQg37VXZFEZYrOqSvKASfQwtFJMpHb/AzX
vtVi+SK2quo5wt2etuPUUYpLohl5EXGyD5IoaaB/JxACL+wkoiP7W4fAVvP29zqx
83K7EwDWrN1JehKRZY5k7CQGdez/w1My8q3gRVLv4ORhoT/VlV8iN+NuEWMPMwea
0rffXn6C+KXe1XwKzPRRxr+QynaCNf1e/mYsj0YAkCO9DwjqXMTd2hEEyfSaNDQ+
JaGrMLP8oPnZN+3Ll2ADRX07GYxbbuAeSTYHRKROvmiQ+rwJgcxzmbSete4ciYgF
Y2L52pK8nA6yCe1wenoPZS2P/GVeaYQq0ZHSfBGK2PXirmAH04KfAVmmn6Cxj6dm
1c4OXaxXBTEXbPufAZdii69hZkQsIllt/OYsmZhktgOa+PliPycbv5eB7T1ujrF1
TU2Ed1/e+6CEg4V/atHS9kaGThQ5bmjBS06tUL/s+cK4Mxst2Q4heLsBBahlZpQX
S07UuM9JOg7Jwuh8qIEUb/Aah8IiZfWP7NS42xIHJWFevpiZbw1eOJUwLZ9EhH2C
ZBDYC6zMn4mJG7yJw8nuOqXTXAGSChLMkkIL3u7rrK0cfPnwydSDi1668lGYV/Uk
H65pqUV0VWq5wHAqTajNWI/NRXJ70jHprbXVZrR4744gGdUUmxXlZfQz9LWGuCrb
WlMZMqbYROplikUNYM6EMTQ79iH7docPRbporRA0r/BRia+UHE9yMvXwinLMI4UI
hcEasBMyG7VoioA3MQvbK2pteZZFphPStPw7xO5QkNtktC3EhqWNwqXWERW6Nrxd
1pWdA/r3c/iBX59s6eNtBHrdWGn3h5xagPWFJq/oZH+xmg5MCDRLgUlEkWiE9ZZS
X9/ZevjAAfOsvTH9mJ6eY48pQhQ2BD9s+bylppDtm1pTEKkfSSuofE6bSb9aQl/d
vjsSSMJl1orfo3FCZ693FxuxN/7uriR3YYEPfN3+xwUDyxzf35Z+nFsJmvjawSCW
oQSAbyJBORPXxiP7nx8TdkDeBbxDiGV6jybDDo7kqXlNm0NlZEX6mAsGxb5cmBWq
tt7nxfLD7OA1hCCtzRG/4D+DtrjeC+pKWmf2XF1CIUcX91f7fRB+CF8tNxVPPrkv
gANFTy1FButMvPwQlXUla7vniyxmDgXb5Bd2IwuPFOLAoruJwZlokY8FS9f3stv2
JbwmCxUTHu4xRvOHvEvXcGURX4Z6ePov1LPYERtikbs00FUWfzX0sZ39TW7wCtaU
27UB+AeEZm+BGkdVmWB0rLZpjBwB0bEKgjfoq5bN78deUcbhk2d/NAU/Y/+oD7iK
ZEoJNaJXQLR7pwFy/xlXrDNZauNeRw3XLPUNFh6mdiWdw+1sd8nuVUo4i3mqTzUB
d20LDmEDZNEJEWry9MsnZw/3lqaruKlh0lO7boKEwE2wwpzsla/A5a/hUIGJmKnl
ue3UD5j0FfKblICX/cC3YomaIyeifAlZltiPlmKgCtug8dpl52yhATj27oZUDC33
wsjvfeT7Cp3Rfyq0JbJp/RXG34bt4SX3Rht10kTHALQ=
`protect END_PROTECTED
