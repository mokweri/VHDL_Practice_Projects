`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gO1Qshu6aBS3HCW/Lgpjjjrf+Z2Mjebntm01QaVHHj0anSntHRH1LAcBqmIG1j4A
z7C7wOS00FPNQycrzE9mRqSfYk/H/qdopnYiEMGfRp3zq3Y/wsygmsy1UhzL2hu1
eG9fj8P02LOKzdBO0RzbglgqTXK/cqYHD6dyN7ILGzx/3iHTA8rOnOWHB5LJehx7
OWsTKWCaZmhXDcl/nySxNKflAcGfsijOt5cFSTdWM/Edna7w3cw0UZCSNr9APjhx
4OcN1oGD3QQFfPxnAbum5qsmniwevXsfxAk1Man1X8ZwyNM5qUHJEP//Vq+JcQ6W
yxTcnUTYkE+5qSM3ooHUW6nw24jyM3yZfXStEjEaIujfZ61Q7Ucy0BdOASLCqFDF
qfCzaX0GYdbYh+XejPvuhb9CyaaqTSykBzzUpLhlnD814POYWdFLBkNVdHf2ZgvV
rrE8AieHd4Gg74tuq2B4aCYVhutfxf5gx5q6VyOd/DJUrGDzvdg6JuhSAjTNB2ue
f2s5rLfk2iW76D6Ger6ANirTQSTaOlYQDSSLF4+z8E0+cwnicX9qucR2XMhcsLMB
yQ4nOBSrsrJyAdO7ExrGzaEX5NmKmee2cmGfpk//fqwplKCJCLC0NvF6w83Arc4q
ZeoKKtcm5dvlK8dX0kmRdBMuI1yP2ojgZpiQPsm+X5fHzoJ4Nm73jXPq71Og6xGu
F4ttc57uj4TYwont9LY93q2XJV6PoxPcBzPscezY08cmVOf69DAyhs26nJTC9yqG
4iR1jpRplotyD0ia6q5+0Q==
`protect END_PROTECTED
