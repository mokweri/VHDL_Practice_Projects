`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xa5sfZBJCQR6ZrkOsDrSeVZXEssKrk5cE7JS/64lUTiO8RgbxigRtHOstVNq4Dwr
9WFmjrlvIHlMoOcdW0emBbZ8cmd31gM4DriaKhhPw7jtPec0MjoX6wZ3CTu/O2Ni
y2s0xl1JPcCNhu2mOg+WaucsCZIwFJmjo+h0OIj/XDq2FlY10hFY7r8F6bweb8w2
M+22g17wTOZg3QofWFj17TWqqs2eLr/E9Hk7OLtm6u6ntzXXcXtUymwnirJFZlZH
uDxsDE4MmNGzga3lmY7lwNlwxeG1YN71PZKW4vIP/erIpGlIpMM9Bs0exa1Og+SL
EWt4wjht49do5UVueFrAG+ga6vlR2+cG9YvtksfQBqO49uhKaz+q1SQGP9leRBt3
njxHazuHi8D+NR8D6PpGw40udWBKqDh5wNuYUdOngRveL8zPFHmz5NyTCFW4iMiL
QZTELEpDp8fa8LLyeiFkyCuMoJATYQUZ2G2A7ndJghhJjD7g8fVHpj2W9Ij64ZMe
aFNTbcOmLTPNMpg5UNUihxKmpsYqCvTK/WLbxL4FKF7+zXOn4hiws7bmvTEy2CI9
J67yVerXtkMWAZjdVnZpiS+ueCgUoURKny3hNI0K9rblNcox6Bs+YQEBgluxOEes
RTDctpDIL+x54QvFrC01rRvg5AKSa2diZXDrgkJcGp0kb4EzqNbjK+vmERz3bjwo
qAz45aYNMVlYugRRZme3Ol5xSGk9i13gB2aIR/ft1U8=
`protect END_PROTECTED
