`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRvWNPi/1/XC2Gjq37E99ZbP0dohcANSLdchYSrU4b1pYQBCxWBH/2GZ9TL6GGcr
hkfANnLUBhsE+a7iLwulzoS/2SZjpnEwrvAEsVD25vzIXnHIquqbiRv97wbL4Qms
iftymw7RL2SNjRR/iL75d+hR8Lx6J9PQ8y598Pie5mDD5xk/cIPpYC6WX/YH0EZd
X3HerJbDYsjmFvXhvKLI915kfa2HHAWmYZ91J16cPSf0tV7FHNDE5z/NuNgLwaA0
TkadwQAGslULvfB6MlcX9DqrXLnkg59MSc9kOroj0hXxDIhWTFqQSB5yppcrXDtd
mQxL4UHyklIQFKn2dVn4vUrXLq0WXdWQZmLnERz3VhWx/pxbqai6RJ3fqFoQETUL
ZMXJEFraHwPPP7gy/PEIeevzUgXMqg5Ry0OK1HKCyMaLw+VKRYmwEuwByuP9ptxO
8v4nMXXIyswwn1HAa+1YwsWltP0oHV5utEg0bbxOIuqJnKGnTFOIhYViXZIuQLNM
MA68asLDeu1pHDSuj5DGn3ILTUid7JF1twXlHKP2AFUEYI5IR/0WB2xxCJgAz+AD
NXDF46fRU+t17KwC4K242q8OyOrcO060K0s6TbIeM2d3APzgtqadIbQqZQ5pfkwt
aETgWLaXQHUlDmT/Pn6io+M0PPuhHMIJ6SQYdXnRp0J4fJGkxFGX3sWHEQvHOdRZ
/l9WDJ7VyLnVnSFh3YO+/CwO1V0njsPIZCz6pXUHTePImMK2CcWeCgnjbum+PItp
5nr2VmheYV8/2yzui1vjKQks0g4ChhcEjX8glaZyEv6X3/BR/FL2+eqFEpbhxKQl
LyziN2hUcMKUk5z5uZTsSi4G4CIrfRjoAtv1pj76lL8=
`protect END_PROTECTED
