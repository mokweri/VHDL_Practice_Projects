`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2GG8y4ZU7Jec4ERy/b0I5yVI17w4el9AhJHKre0KtqaDxxqPT7PxS5rtSAJfmDx
wTvmU7bi9FEuFQgw/6bR7wasMbHhbwlSz9eVxtqIJkeYem/z2tGNiPjuFPd+n2Ha
Jo6VKD7BEkbvzJKP+HXyShuQuZuKNoD2DU5/3Iy9SVI+fI2u2mgid6B45R4Rkhfw
hT2YN/mbTkghuyXdCfzFSs6WzxuJ7bPWygvamP8Nm2Foalb/JEFV/CygOzZJ2eDd
+QhLCLLubDh3eCjhCLGTP7S2+/IBM9Ov84AGBD+lp1o/tDwnDbZzR5xewJdfJxXT
cJro+U4cB3Ny55prESGuA8ouauhk3oVjzqwmNGiJzNna9voZAUzknWqwxWM8WDFD
paP91r8PHWIL3ZJAPfsfAMtgytQFWCWuZyD9Pi10xIS4gRzcwaawJF62PsdWNK+A
Ups7pKqmsL2ZOa0mr6u2rbSqi7zyEhSgXpz5SAzll9L6g0aeKxNvOhZ5ZVtos7f8
dRbsFDH0XM5t3DYeVHw/5k0l++/AkZ5bgNJ+OuN75Jd0CvyNFe+8PzfvfANwuRot
AJBYzpDcQ87CV9ytN7Xqoi0WzK1NqmuiaJ6gOQawhly6BIYr2wfIWSYTKBFpRaAM
fsRVKyQCWz0SKjsM/RT6Xe601Pw1DQGLTv0vxlQxYNk/AnPjy0aXRyHSR6guusiJ
qjlo0bYqfxluyWX29ZUN97mxvB0hQmkKVcXxHanpGP2KmlASRWIdErStbVUxtsTl
x8DH3CigxARnDozWHYluVblTkvrHBhDAdTKyimQ/Ej9VUwwZ6FZ29C7RejLdqlXK
NxyE9D65DvcEn5yj0ktbHCWhthAGw/RjudQKihUirqBIrAXht2bMayqBjgnIIDdZ
ZIurlevMeq2+64Ep29m/I0EARlZGjCa9F/qx90L6GfjRywVu3hP7SPrQOSDDAD0R
4zuwfZOI7IdTYRXXKnyTKzrPh1ZJ5Jat8meLyv6KXaM3juTe8YjxEE11/4M4qWF8
sY9JN/y9SqYMBO9I+xIB8EzlrRDJF4F/SHuw0nyNIzt/BIDcfNblrIypgXhh8sbo
37NUfUPq3Q7cZvC59aeZFAX9hWMzVTofozHYmp9h2E2HD1SY6u+gxoM3g7QUm5Lh
gxxD4koXy0dWJnaYLB8LWGGEaJWPi4rAe2vMEFtK1ZmKn0UZqt0PlMB2CHtqcuDx
yHKcp735B24qFR2KPcZucDEREKrOn5d/vY3zQOqyTzRqE73iWbYR8eWkVbJfn4Th
bsCwKNBUuFnPPgt60txbjO3dhdlv7I+HI+AOeePTzcyziUYwjgrVKWZSdg3iBfv5
LAKQyCUhVXFHyMsmY5ceKxtXGORsh+VVf/W4VOcAv9wXhq7AOfngKio/oIoDLed2
BFOL223xo7Kn+zi93K50/b26S8eUYNfNS1WtVwhHBWrP77t2Xe1CVSapyvew0mGl
MRmMA+wkTRu9CbIrVl7H2PAmjVFzcYpxZ/0pxr+Q2NK5Gbwxc+MNYabQuE5FMy/H
MQCD8Tn7X3iix7rO5Jdz+lKsRagn/n7Cm5tK7Bys1b6MmQPMNCqPAwvVK6VXc8z3
63mfWlgSQi2Fo9FcohHQwGYtxbjS5TCgMP3RPtCe72PGU9o7tuMOm5b8EeswSRYk
NwUqnwrtLFoktazZhOwfH+NrvwUmYqoZDHqXdjYBhUkHxkuIFuJdOz0nAW7Zx3bC
K2kB7tKfyqRufznYov+ETuC8ZS+/iDi6z7oxJWDc/1xoaSd1f4UBo+b+jdUcdN88
wXszkCkl8gPNU+PO8YL/tPz+eeKVa7yKlGFIjDInIbHZJXtHMMnZOrwsURf2PTQ1
WN7hTXnoZH9Bpj7j1CfMJhO6hPe0jnS9pHZktpx4C1GIu93iI0jHMXYKwyAU80HA
PVWhFXul/mTatifSH27MGb5Wadqw2SlAygjHpd99bDpq+VPNE8CA2bWx7WV2nv08
gEFeDei+Z4pq1zgIQwgJv98eXUXmB3wWhFULa6dnhTUdOXpSJ8QjVtc54W/rWSgo
R0T9Rgb7FbSIiQjjlSEkGTcnHYOcBxVRFYTFawVrJMNE4SnYO+M26Ri54UqAJOIo
EbNbT2FkvvFgxJtiwR46wNtxbJ9SdOaGFm1MewX0/pQthJ6tOCUyGCYF+UAiUeI0
3bC8k0u8xbTOBwdgXDYSBQE/YhAexW3Qm79Pb6C5x/ew9Weko+vmv7GQymdBd11m
dmM3il4yKHZL//qEFvXuYMOJDLwsqBgLHKBu+11pDwMjW/nIn93TudAOk102BAWy
zed0iz1A8plP9JVV0B5vBpjRciajrlQB1BdXo1K473IDUwFpTWAmBPc0ZTTQuz9j
J9MYGBdyVaJLntUozeGNEOPr/ZenNx0BXZVIe/UbM9GuUNd1Nd7knv+b3Mtg+Nnx
mhAKt2tCHeZz0AFsv3UrwAqs/mUCfN3KD0Wf4vkwCOZx2t0Ao7KU0/rkCqrX21D8
bQuZ2iA/KQSwlQP0b0FR5ZPNGrLXQtM5TtzAyzNbtRugwYhSf+O7IOtOoqzg/Smj
qia65p3ctiKDGyXOHRhOG7qHDoGz/2ab02aiks7YajclhIrhihpQTXDlHN41QTHz
zlhgoH2yzZuCWgSKOocfCLyEWOlyX6WkW+Bdvxvj7hUitmNc2mPmrDY+jTzGFi8N
X+AT+UIZwslZkFbPvy8+7V4IE9rKPWBX+Iq7R2aPr/+smVtGL4gluE2GJSi1tQvp
sSdyPOtHAI0AZT8uclG+URBhf3l/AIF7OYHHmcW4b8yQTC59oy1n768A8lje4NUi
Eut+uHCtx8T1DPgjluSQOD43nhy7rJgPg3ZDXyVFeqGbgUeyEUluHmgZpd1Tfkwi
4DBkY7NaY1xrXvs8lIWkpCrUOxVBVpJx8FXfMx3DZqikKWAbPGiK8Dih5R91AZRz
y4KhHbng/i31tzWr8CqVMwQk3j5xxCGOU/bFSK07czTZz7aK5vU8CYISwKSvyLKE
ER9T9MuqeYVsDvRUAfO/LL4/UitcYgt2ejCxH3tuW2oqQ/UczQfgqDAsZk3dU0Ge
4AkVKe14GQcf//04D5Azmn5WOiz840E07KfacnNmbClWs4BX33Q4LPiN/EvLRqSm
AMbCrMOXCUfuEeT7EowL5F7SwWCIjTBMxjPBHxccMxd9XLK8vswhN2fOoxorqgYn
3oGgVu9dzLc0V9dJ/dDHMXjzb86/IU7L/sd7BX4wqGviq5XkKTBPA8GW1qDG/HVQ
GfpFuHnSWSHCTM5UVBB+9GBxrzuGT9+LqA7P4mojlysN1F9CZvVTpnbvbECy/xCV
uTwFpml9d/Faa92DOJk1h1K4K+avsGVpxfWVeV2RzpLk1gHIeeyLNkIOBhme5+Xp
aD/fJfG3KXQjG5jp5hEpFVLC74LF6frvOft85Z2Nszmo0ds/EphKRTcMq2koXXR4
ItA7d5bRVD6tMmzL3/MXvwXT6yf9clQGx1XN8Xq4yR0d7jpJI1j8c6qTUAUll/wG
3+KmU5IknFltqNNDXgck5Vm/zY8thL0O8VRSp20gWIpkTAoc0nFOvisJ4+gQbfUU
MmTV+EQF4rzxJ9oaFIA4UON30HVdIdBsnlYJNq51DDR2PJvMRZHWn2QyjooYtzwN
ytQaddeZ+iJsgf8IUaiTbYQNc3e1KTIr1uoWIfwaN40AevFlPHx28GrRfGj1SbZY
VRIJBGRjGxCfqPoowmL5Vuy9hAeznxqGZDgUUuqkuqHbPBfOP4RkWNOooCwvVKiU
RdITCg6e01+xaHmkXJnwjEcSN0BQ+0HoPt3jcTTs+iMx0n5REL+LgHNMHePxlkWw
oEpLobTSUhWuSOW/a1x96COYpkdtOfx8IYmBWP/V/i6Je82Tp4kPplAJE7fJd36k
DqFj0tSn+9MfGNJXqbSv1XRrzZ00sghQsfbMa8lvSH1yMorDwmIBuw3uq++Z3w3D
uzuAxffurINY3xiqtXz6zO6/8Q6PmEn5JyNhjQgKYPtVbcYFB296Q2gk7C3cEqr+
kE4VEnjvHBseyJ0EVfhBZjDoupAv+AuipsXFGlsiP1w15CBZhdQ1ahnBkcYVIq3V
r79SomrRd4HATCGvhuW326mV//XOe/PRhsR3gjoQcea23o/IxEsRbqHimfLsmq2z
gdwOrdeGdZcO0SBOAD5BmgENzYa/g2lDtL6vF4Fg0Z/jROqk1b9hXi8dqYb7iwab
bfkBuVyLYUbxUlwsmf+wHuWA8d4caJm1qoF90IAmVUpX5uwQco6PGUf6UtUldpXN
RSv8dSw42IXB0a0eZHhxQfP4ysZhGqWVjYFprdgIq3No3Mj+UrII9vTAF0sl43Gi
dUgKPmzDHV2fW9XbBfKK6Sm3ytPNHKLujzZ3/gHXaFgl/GmiJ0RRjDsxQMKGq589
02NEJb2O5/zCovrZ8hfPYGC2owB8OK3DsHGfdTRXppo=
`protect END_PROTECTED
