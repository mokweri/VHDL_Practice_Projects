`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H7M92pHwnBXo7FcyKvAts90/s/V6ygEZIDgPV1nsvJ+tvmme57wnn14+ldoFBGil
YSN6WVDZCgijn6zIKw1pmGdXF7KMMySOQEOERFk8Dr11ucZQUFyc7vAwqGHVFaM+
NYpRP7Q3xi7p+0o+bUxuMEjHrTQCxBSlry3P/TxjAq1yFk7LPMfB8Z4QydiAYbv7
gpa0ZW7sQOKfTMJg/V7RrES9v2trJNi34i+28gfwP3LhHRl8TG05Bkcce59kEbtf
7+RWT0N+7dvcnuUggDCQmWgUjZ85UMScA4SVD2OVIAQdWtRE8TQOo358uHS+od/a
0n+mH9w0xV4tzc/Nob/eAjMdR1/2enELxFcWBCLWWTkKantzPCSlqnbUJZnMsaQ/
Za4MP+bKzwvIgY2tVQD91j9grz8bayUTwFJXdhisVWLrFAd6sUplnw9LrfTf4NtN
C9sI6d99gwUtEA5TUolbyrItmLHY6KgcFytfnNvZoct/g7OM1I0O5JbeDo55siWn
ASTIicj2iNDZC948vU+dDnV7xQ0w+rt76RRl8fIxsmxpZFBzKEIm1sYzeF2gTG7l
BU3DZKVgyWl9UPJPtdly1IqAOOg8pmBS+lGXE3Opm9EDebPxrze3ZAR2zNoxElCL
N67CT8QkKi1iJW4Q0/OmLSCtfNd8WOMEAn6PdleVj4iZOTot8CPZjc6hzCVrtV7g
YXihtR2SK0eZBjdpCRlpGey+3qBpeXCrWy605aXq+4Mjo0jBakDBgpF7iWYWGT/4
QT4R0IV2Z4wvkoy5HtIVz/J152csAImCdptPsDNnR70wDjmQwZd+6yj2WB7cpj7r
VBArPVC/cNvDHqBJYkvswCqHr32gTRm9zVQMUHQCYVDtoFu9DgN2VsTawI1pi90n
EItY0uLA+zGYPs+vymkftmi00I4mr+ND7jSfb9gi4Jp6CSv+KB1fkY9OnRLa9Ea4
QlQ7Wo1hhWYab450dxocYvPi7Rg5/5ZXvS/9Y7QqWosu9643tVF/uqm1FPAEsQuT
1srB8ZldtVTo2isI5GbMsbrH0BVlnKuSuyT6nbp15ALJr2CyrwswJLLzoXcFmX+4
2RXCd72nMt3jFwFdODp3zFu7ce6gzxv6heX9NphVjNSQctmTg2dQRxO3bE8vwWW0
dLvU7EJx5xnF5g7yITW6eTc9CsJ5ZaH+TJz22NVIwiw2Zt+lOusfK10sXC0lQZUI
Z8ExYMwTrkU5okNZQkRhJ13pkorhH2jOXinQYTvOhY1D/DHDxafRv1HlX5JwMH4f
nnY/nHgr2weEKhSogSz+Fq/5ZfAd6ieaPafQUH07EkORNZbdz+u7eQRZTH97G7tA
EnEbydDMaUOrVGkvzeL4ctSneA+9CzQksZDyO7SdwMWLMKE7thKxug0uiY8byR1Q
jAKUmv7aCgmWwNwPmRtbL8WCuPWv+LSavIDg93mJcJK9UH6qVsMqipDsoC28vTu8
R1hoLfDNaxkHwgm6fs8X1GUVtrkJMY0lgiAWBE+ft8UNMcRlm1MZAWYQb2TtDg7n
Rm3RBFt7Pv4wOoG7rnkjGcqmiaRuEM6PV7eyhEGLqguDm9ZAe730GZdyhus9/Sz7
z/x4IOGE1O0lijzXwSJpSId8IVRSASjyp0ZSBYpWOVaac2DmBOub8B6QyvHyshfs
FxsNCh0UIys2gOq03ku4sVmtuXv7tFMUyLECg8idBBENz/oM6gZ0RVpCzdrAmOW5
FZ8JCYXFYIZZGiZ9chi4RlBznjlgLj0xJayKtp1a3PULmeVbY5i6gzX8uABkgAbK
Ud7bTyvyWFD4bYoKdouXNxNCiK+/X/Xn/sKLqZOcdNuAbSr+ky7ukchdWEs4K4wr
JuRvl7jDu/Dq9FjVPIC5tJESx0g9tH/bwQxg9R36PNwT0GG9APleKIb7lF8uLvWl
4qUshi4TIiWJ3t3S6GwCsQucmkbXapocPFzJDrqdOnkvuHC5X4YRgkFwcID5T8k2
vGutlHtayeVQsdeN4SM80AG/Lfmm3veb4fZg6ewog8n5rTBHT7L680drQ8plWZh6
KPYYD/lt21qnoTtBwABCd3eXO6lzDfmhhd62ib6Ijw0S7/LTZsiOf9vIgfVGRf1z
XyFEInivL7eh9lPhiVZpTdrVDw7uVDKPHqmi9h1OSf/Kwl8F+yVYcH2GQiE6EA/H
mrNBQD+iCzwSv7cQaxJYd44CTmXkgSBxvgZSOLGJasZWAVFKGFKBtmRgoOU/U/l/
CKzoCYGvONMMU+C197zzQazRQO5fE64pPxaP5Cy+r91NYEmyov20ZXlzNWyY4SUs
pJ91wxk4uPtluNCUgaCVHTOrLGYRZtLmjQcQQlsuL9Eg7PiqGefM+iDVNj98Q5S9
n4L1Cmqyo8hKmPGNOpwsVbPlHA36ZS2EttWtbSQIj2yysv79JY/9euJnWdtFT1CL
RFc/+fUR5SPQffljDaklUAjPOonEJjs9j/u8D/FkY3LNuGECelkR1sPMpI9Rb8C2
vdZ7AIph4pPS3TzLcgvM+XRVFUQ+I0n9oxHfQrOKMQV9VXKl+JgR4KVTTlaSW7lt
T6V9e5IIByTsiWF5lpMVZ0VVdnOdVYUvU4sP3u8Hd7mWMRxg5PiOnHNcmnw7vVYY
5usC2712xwMHb2nbMOP2BrSWdxgHX8NF3VhvAeugg+mOhra871IROkl7ubBb4Eoo
J4d2nhVnEBKIT8z0R7cguAERzfPQwhrvDgvtlsKyhLjiGSeODRs6Imucnt8a+HkR
/R5xPPSN7CxoC2oTwmof6O11wtX3s7chVepPaSoSt8l166g3MwMAWnOu41G/sjdr
rMlpU9/cC+qgLkGXHkxMmsZl3B3zOh+kzCyUMrIPngNc2dTIlwMyPx7Y1+qPFNTJ
iesq1dReY75mewj35pP2wAMcD6SA26J32w8dZ2KgepxMd56XC6FLGs1VttsAg5zF
IAIte4SKmyZpiXkAQ/el5xA3sBCgqb+SzskZRCRuzh70MRB5YZY3ToGuvCqCuO5r
l2qKStmljRVgwLQoNPhJha3u6ZWXYSBZUXpD0000etcjji2hndz308V7SI6DjEph
yiNaxqKbMruD8QeRVu25nfIxcESIS72un2Wh0d7IiqtNLBrFtUUJ7W2fWY9bnU4X
h2oQSaj85aHM3FfpkiaPGl68iY1m5agr+7p+53THKvMYY4fNRSexGKAZa5yC+olp
fpb/TFGDsQ2RLSsWqgZxt8ysvuAbSwVrfBoW/MfWRjQXeXfWZiHsOAud8ZQVZrDt
69rFZmku7QC/HMn3T5SDEbFdK4r3iPH2U6v0yfH7MVz8v/bSazFm5AIJpsYkhRm0
tXpUOSaWQekiztROj/ttfaqMS7acUUxez3d4AxZDwNFR/bXN46q2jyY2fZyEi2/P
hDoLoG0ei8aLrMyaH0IHhO3jKIjZuPcUDsCtMxxl6O/fJAqFC5PB6L/VNsU0WWQX
ukj1jROEsAd+UpJQnCIyb3bRX1oUkWYRnc4xkRUAZyw8fHCN7ksXnLMFmk1sbP2q
qwVJcysKz7JTjmSxtuCNSkXsUtNZO/8K8GunKZ0iVfdPXYjZp82YMvkv/nQC/9SY
ma35knHU/Z+FsAX+Vzwu893jEXz2s6FsxJtToMWzWSAMMp6K40AR/Q3pR5ZjJwtt
yIpsc3dCHzmwMZ2OYVrLA9U0NPOR+ANE9TQ96oiKemo9kYA56zf0KIOw0m6GEY8U
6XOL8gZ07wf6MNf1ZZSvsbZk0BgVPotAk8kIlFNoSieniYJHDkXGRSzhXYyLT+d1
J6tKVruV74Tu215y9uk5y91K9OO/UCNc/47cBvSnRKmENPKSlm1tHIFDueAvtiT+
IDj5ck28Goa1RoqsE4VTAFJb/IdBw8RJh9fbf82J+0zajDjd51IgIVT2clR15eUT
h7x25Ruchv0t3LHLCBXzqFyW/qlHUKcDgkuwJXaAGgi9gh2Y2nE3jPwGio2TIFIQ
GTtcClZKhba4O8HgUS20cd/r+1kwfP/HyQljRaOCfXi+xJ7/i8wrODBB3Z88cxJO
tQ/muNX+U8EnMnF70XIVJYgYnpUq6U8pfI0UYdtAE+aj4P1uc/6GS6/tlWC6yzxv
hA7w+s0MJhxDAQBDVILWrfyRY5Eqm/vVI0/JXP7obzud4kR9E3IB6yG4re4I/8x4
SjsUGMtE+BdC9M8h2j1ahA9+l5n4fnRxLaIbelamLo5Il6CDvy+PuZ+h8Whl0a6S
JPGBQ8xwOjyApbGx7tWBGI3c/XENAaNauZtVIkuagJceIlTSNKglqcQ35R+soCG/
TQUXf1H+3UuF6uuiyhn7V10hspfbYJg6ayFDHt2cPTeM9T77i+dXRZuN4Tik370q
1/4oQFgzxWwFSXxLnNLsLIrVxB5eyol5HM72KxKnT7PWyd6+POra2I8jmhNdj/Rl
gPcxaCQViHhdAqgpkWi+9dLRVIoII7VbxEMfMsKsL2Gbz8FJA/cfaRmLLdNc1/Pr
GsSn6pdac+wIDHia4a9ZsATiZ7pwgBKlGp8x/GjeAi3auTH8h19QRR8GO4BBOa2F
xT0RDVRp4H9s7B9pKAG3wgyOgiIhym1cbmdwWI0oMa1xfZD9w8kYWqkJvvnT6TaP
e+XepzWSuJV3cZBRf937hW7Fpx21so8fM+ZtkBm2XJpkdqyhdFqTx46g0+b9yPTb
RxEw4geecmoEymGWUK4ZmMBUmXxDbAbU6I7J6NWso9gxwm4avjRsyjsIGj8V2en0
wHGEgJ9D5ttHGAfAbMeMqn7OHWHNtuNz4afCBR6qrTvxl5bjrkIPGl/Z3ARgamSc
MZxVo4GBVrKzfc4cdQwdxmkHWXaThohPNUPqHh5mDMU8SwOBm6P7eAG4nt022Wdl
px55tMBuFQK5JqajxHtyzzNAwiLglQZdOcAxeNYnia2vzRWOmme18SM9n2OZWJMn
X3KiJVkQC5P8Z4EJWAo5GIA+kzk1qLLVUZHgX2kOFCAHsNpYyFA7z1/1HRntKgy1
XyshRBFOyl6dCAPw33O0CLRY6RprDfnOn/f6ptZ0zDD6NK5RjAESH4JXO7IP1Afx
Z35OuYABbS4gEknF41UcyRTpkQQg0WYKoJxHpiS0chkyfAigPTTYMIJ63zLd8e5I
WoeNu075JC45U2z6/om+UBHCuTURV5dtOilTqALsKtlfI8atz/I3p9AJMC/HEVrQ
N5DlwyL+tlgow0bRKM0oMSr1XG0FKTZ2zFPtreJ9IEL6Hk8QNZqWf3+5UNJT9P9d
cY5r12GF66Jad6xOMoFKbpUKeR919v60cfzsecX/4VDAngImHmTHvhVZkUZgR803
ovoYjfbHWRUE+W3hy2eawTshCIoJ4bOKQuEkmQmeGWs9A2ZDA2LLusGW4XhFBYqP
c34K4oUDQuaMvnzp9WswEPTJ6pguxqnMTjZHRPAZkibJMzecE7Aree03UslR7bY5
VX5D/r8HQc3K4BBJFvaHHGzrQxhI7vwk2tdULCkccENkCkfX3bafwGSRpqPi2T03
I/7lFr5gK94Y3jDc3Yj7E7T1Ctt/je9ZFOTLxLe34J0aPD0JaedEpcublyW8seqv
HUtqGbV+Oy6Herupi7JldAYxUBDkmH6HjIXukLwfqCb35p4nFJniVUZXKVeCXPEf
Y/ybO6KCCVp6jr6eI228RFz+qzfGrqy70IPj9Ryb2IvFYxEf94d8mxKCFN8DotT+
43kFFbRnCjBwbQ1GZmrYAG0An4+q1Mt0pZaMLICutv+froqA4MTS+zy1XgcrIyTl
qJr8oDg2pYq0fjSayE2MjK+pmhRX8iYnTpinVcpc1n6vhURPXHL+QIFnJrsoeOA7
R97oT2YCUgylK0ijuADgbDBMf4Xg1+trOkOTItGgkat+H9ODpMApgPbuMVLSbMtu
0BNzK4eCVgZWzQ3gwppZnRagqMP+H7dGdZgMnJi9HoGfAPgSN/WLugtaD2HJ9OJu
y/PpJUZjev1Ink4qc1TOAGTgkFC9Uyr7T3E54BfJMaI9mbs9f6Twp10shleuFfBp
cOzLQVsoMGibk6kXyFTVHqczbPjlhXkv5qdF3QokkpKMtOaSokU1Tpc3gR7fnm9d
`protect END_PROTECTED
