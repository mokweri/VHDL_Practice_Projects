`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AVgF/fN/99TaNjJxwPBNML1/dcnCSAD32oq7ZbtM2UjACwyhUY7r/zNTYZmy77Nd
DdALfzjv7PhaJAe3FDuzCXHzzH5CJvQVbOaZRlNxAmIuJCyNKXGqIHsYqoGCPW60
73Mf+gT8Oy2y2DmP3Z9SsgAj8wacGSOWUdIm8lWfijsQeVWJr2hrGSabDahv9ioN
y6tDDrF23kVW6J3kedQdFUej4OWvFHpeFFsJFHvhIJGOJD4qIJ5BxKlnnYGbboSX
Fa+uGKJEnIr2fTOW7rFNRQPvPGjEEgJGWpgOlXpq+Of6d5ms9kexPqkGMDEbarV0
W8THCbjFKajkRoxkybrkHnHjYR99jXikWt3qg60zuGjrLlhxtW3xN7ULQZS3P9dF
XFjKQgoLLkBbEj4yv4fcE3ZmRMDwsvURyb6YA4ERuh6PxplZ74Y++9eShQprKJPv
OuZFRBp1hrcUIsLMYp6PCr6JC4L5HJ18if0cTHaUCXMjKbeyzkAnGakhBzJ/kYzB
HSxQVegRT0VBOOuWAxO+hrjaui6REmkl9zKDVpPIxSSl1I0Nw6Rp3LOy0XLYADbL
IEW6hWxnTlFNUn2c6obLbaj/GofYtiBHwqdCdPl1Pi/XX6sDyK3Cw2WB8FKPtiyN
9kQjiAWqvKNOxFC0GNBFT6HCYx4n9JQ6gyHTa9ktZFOPdIMjooDYkanHfa7OFKxM
36rNPnWjU7OSYlJtEf/0IUOLsCVveUo8yomz+yX8SRxO1Gm4WUrtAutNwQQgmzPX
pBF3fYXoR9VvG1CFx4CNE36oiy5rwawc+qDyq/I8aEi5bL+CwgVhICEQGWGv7wJp
v+PNLqzoJmQbOjiihWviDu5hCYbEARbohsboqZj1yeTwOHOFKy7PvXYFIC1ubZGJ
v38JBrmOyuTuldpljoCeoGSgyhvGmmExqxS7B/cGibL06aRpxX9GLJ+zx9OPegnM
3NnqZUpa0VjM8dufbiTFM4tUA5TE1JULDmoG28rkbJPaWhkj+5BEYDC1g98qGNEe
vpYtmax3kOxMMx5ehrUF4HxY5tod1FPm5nD4LrC2EbOI7b5P2A8SRZk5uWN3lF6Y
jrgFH6xZOLiVj/M+2pilR7cVgDcai30Gyh4EUupukJ0+r8MeKoNgyHmfvm9m3NhJ
LK76Bdu6xkI8dVaM+sFiKG3HbVNFYsASBGWnmhqAZmjMFA60fyuWlbc5ua+AiuVI
2UGGlzHuX087KOVr0NoVSF3ovoz77X80s6cm2Bo86ZF7JzlaLrp9FfmV0dMi2SuJ
TlvCGpF/HgVjiqL/MufC2PWBf48k9ykp+U2dHRSxayn2jEsHKCmfvSVDgXtsVJaI
pBdTrGt3Jp8he//jM1mrxgsUPfL5PftbBeRoVFh1bt9sQtbbaaU+19oIol4vadmr
+j1VHEdFEov3EvoO8nm0nOEmZmx0b1/tlA1azrTjt6tv0vBa9Ft4i1yTzX+qdkm/
`protect END_PROTECTED
