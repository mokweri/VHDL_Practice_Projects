`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFWK2gc7AXzwTtjrcK+J+vfCTYVWljQDZQEujSm6xeTR3wu8rCEpoc2wOCkhRg2F
FD0EtORK54VryL9wAhu7ajry2CEU6YST0W1JcHfIVp2o43EkeJkxgZ+AcA8Ojzj5
7fLoCyuQC3Q7X/DkYcgMBveolYvlVQOfEwKbzpd8saNBBjASsEloLS7quCfWPFPd
obxFfJw8BwmPrQkT8EH8gkVW8qvVQ4jMxcwphYwI5GUAKOvADNTD9MiMll4lvurN
l1JVgF9g00sYl0DISTjNAr0hijvG+zk72RdevnW5J9mLt/rb8PQ022XaO7lU1VGL
9go1t6kusTFhRKHNvpbU2pBzORLe8YnrXwj6It+R37diSwQ7DR5RwJS4UItiRSOz
9OFw8EAgwHHk4gdp8jEd/rsJhRl4aTYS9C6msLoA9vLJsVwJ+vdHrInbDBaGGA8k
k5rhrRoU4A+Fkuz4ESgh8ShtIQOE+AZ7xxOpyY8nbz2F+aKpCW5hDWpxlRAPXSxC
yJCrFc3440koRIo/xHrXImbhH5GqvLzCP+Q72tGUD2rJfJfVl56FWoh7lftg8InJ
eZkaqcrTyjA/UPBwFHPE+/pkbnTTBkT4/u2OvSyYomlFsHjN+2QCnsqiexEEa5O7
pivCFPRFJwc2SlmSqS9hD5QAW3k2UOtXSKc3c0ZxLSexZc58IMn1wQKdIjjnGhRx
n/HhIRDsu1wDoOKZuq2SgK558S9D5nTwYAvr7XVwGcqzdYGUn7+6AJQA0uRr+mpr
SDTtbUpOUluABmN7smUXTXhsAqwck9AtaoRzR/t1S2bQQrLvtmcuPKDQQ9XA7Va9
cxvJI82WXtInFE9zOc1pFP2iyo/UmyZrKhLp/gk287wAdcmpVIzgnaznUybPlxXY
XtWMgAHMb5wU6XhfktiDeGJPS/WKTUIgxTXgb1mPvrjREOSQnpfWlhRbrCJOUwXI
63lsDpV0m0LqOzn5oXQk+Nw7cF8TB5WJLVcyYuO5mqgltKtlqI3ht11rlVy5mnIS
LOOSL9AHON0zjWVe3EwVG1+yOn2BpAov+7xXg/RfTQBD0UdHZNAyfIUIYYG3mPJX
afIitNKi9E+OCJgczjRjUM/q63khdfD8kTYKNqsyyjPcRcPa6zmaaZVNpFAMkbBH
Qt3E07fhfhyE30Tjr4+5DPolu4FQOrNyynjtPPPT/7Mk9Vidxdk3XcFc5oXHVBP+
birwg2NFsn/jf41EmMFv5gTpLIqbTO+marMmASLkrvw8yXQiI3YQdR8oPS3rNGe+
Uppq2gF0aG3dxlQVAP3P7i93m0dZOgTU5ij0Nh4H6tEr2u6aKtvWCtquRgIbGHhw
LMk+ZbfxEvMFEM0CG4NN/PMFUwLUHm1PQNOgN2lgc4eCSjSJO7aStcBW4xm7zagj
UIlLYutJVi+oM+05KeklzCLLQ7defGjfz2ZYhZNnnqBKzGufpMWMIJEcMXYV1kFB
`protect END_PROTECTED
