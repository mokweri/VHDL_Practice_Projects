`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2tRSHABNkun4Xn+utNDB93TUpoHE/xN1zwQD6ZoBbsBXoq14n2X1d5O8wKiMzE1
1Fm/xJooLjgvzxED+MESWrLFjWRKtr5qUOqzg4W/Mg/L/e9UdcUNulPBi3BCQB7d
zpycrL7PqeXh+PVrl9gZ81leQWyi4Ejvao7NyBV0uBTk3mHX0O45kkjEucRFSK8q
/MOd73K2zrzgeO6i8yWHPVQ2C+E6wUixzjQ+zFVJn52nTaaH4eKAZBUJrbsFovFB
OOau9AM6JMCJvcRH1616MjpAB3sLN1rTB60ScnD7x1hlDlnenLIk7motuRSlvLDP
MwC2gusW+lpvbIGr7rW4CcaEbty3HxaoTuhOTs14FGlJopnby2LAnG3NIOoHQ/Sw
2zvyDqvjIrDkFYWscaFZVHLgGcqBZ5F3jCoH/0EYMu9mqpmTDxl/TbFyLt/0BVog
oTyH8GIaS1m1LUu36VSi5YjTS/IM1kZzYJajt6GEsyrOr02XC0OFapl2mhCRXP7h
lMDXDNN7ICbXgnoi87LRtd6iIzuuP/xxj9Ad00vpvUPqTtNMYVenIfMfwDd3Hf44
fcjtuJQiY6k4S4sWVm+5uBjLEPvLtqaRYIClg7W+qV9lrHoAXPo3uycWaNATzQqe
HEi9Q5yu4EcxfV6522henyCa/7QwwNhRch7RXHJaX6BAsN/5cd4zC8EKyVIKfP5y
Q1aQKd7FVMiQ92Z1lS/0JUIw8X47l/7JSQPI42+eRrJxodQo7NmOCJb3IIY/qDic
F8ajudTMCJQ64qlmWFVLtjCb2l+/A/C09Jz7bP2eXyM+nWtmyOK6CWBqBj6F8AYn
fWPBqKzV2HS4RmES0CQk0uuo/zY7aNlXZ9YZw2dvhzdPrFEAa7Ft7zJRHyCrcwWG
rtEFcWgEeRDGm417Jgy+nA==
`protect END_PROTECTED
