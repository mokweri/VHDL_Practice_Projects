`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIL2AhdWpYFyZapm5fOJxe8euSwbJI4isPEsC5yrWrfImdfS6687LoEcYnZtLiFc
O30PVuqaq/VhNLofjbaZXUWjDTJMZR/qQh7511sZg/hwdpasaw4tVmDGYHNmxgYm
4PNMP3Hxg+PvywyBMMBUEWfOdm9MZ987D9jje2ASK9OnfsQosnvhJNSi9lp7weWe
WTk5KfE40XxJEzbI01BUs0Z12WC6gFHnZ2+48N0WMfUVYt9G+fnEIQ39gdYExTHn
mJnzGwyF56yz3m1VeM7xkrD9on7MrqfiTxpBqmF7SL4ZO6g+4TDcX0NxzL2CYqa4
HeMn5xO8et2nxhr2yJNMqHd2jld6C3hK3s1cy5tFFzoCS8k4CEc2GD6R1SIk+eJ5
zz7T67cHioK6W7X/VvjxXiryb3kLhYuCwYuNBMKgs/aDyPtOHW9chTeWy11f2ByW
jMLRYsz6PFYuiCdo8DI5jW2NCwZ3ptnBh77l4ixTu9jcHPcxLvuYX5y921vzQstL
tuST4T0SBwWmv7FltcRhWdTGqzxCMLOqus3jZAFlJDY4vvI+bPo1SetwY5Bmr4Pb
AwLS8CjUCHpghM9L8cJ7lQxg9Tr/ueUDN24cObpodCYYEC+3xTDRLoK/rW6FcrYd
h/lBbM9EMeqmcq8lGw/L7W2hHKnDBozh6yVeRIDk+GRY8nDJQfphdPKXwyDddq8f
h2ExqM4srtsfGv5OnVhec0XjQVPnqvKvmTvAuoXMmvEmRRzoG4K66KA0AT7FqsRY
lnmjJsx6u/RjJiSwYAHftdmgMxMnccI5+opA1vlMf/OqcEeQgsSSnDTA0yFC4aWE
NA2VJDhOqiUScJiLZtPWqD2oDbfW9TGHPVfeqALRcz4hDmmPwCVjUtyruZTk8jYM
wSemDVJMgekkXSpDliB4NsABEsOwr+xogndDxrTKsnGSHAfW7mH4mDKgbwCKqV+p
FUZRWBbkEARPr9qHYrpuvX6Dwd0lBcF5NE5w07yOTAF1kq9TXwHQYQBwpORW4l1e
25RHI7UWI91nGKtO28ctVt7XX456r0avNKtGA16amJkl0v7pWnYxoZErgp/XUbR4
5+4x0PonsqWEB177/RlNECKa5LlghJRxQzq0bOYg0G8x385W7GaOIRCE9vn0zU6o
NBeeHg9+z66KPqhosUvOj1BOEndh+LjKRTuJJe06lER0FKWd+3o8H13t7K6LJvaw
71KUzWguLcfzfON9GZ3XRXsr84NyKVDCDEeAuGzJg99De7UI1UrMH4vghuga10V6
ue6t+OCeEEM2TuVxJOFIyLjIGlIsEnHW98w2K94Xzl90TGppR1Go26hH6kvW+fxQ
9HenpUYj2PDKRKC9v3cO99/1ycTGUx98d6xTA2tccqKzyXlyCkOFHcx6pBePvG/b
yTo4LyJOvZCPByWDQfSBL+/UajtHFw5BxNdXOJFEo6L0NiH+/0I/YpWZUG+qpPuS
pmVv+6y9QoCFH3mgcTJ4GofKVm1DWxEM3by4JoXOOk0=
`protect END_PROTECTED
