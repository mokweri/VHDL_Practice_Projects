`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aySzNLYWOtkDi+nCbbkrJ9G6fCZHMEemx5TgpkItqxhUEsWIIj8grbhuNhYzCC7z
eu7IV5D1/akDS5CKOdNOECd2pf5HoaBBMB1hpLw9tv3ff+3PfmOp1R3RLvpyFtlj
4kyLjO+gDleocAHKT2zQtEqyvr7FlJ/2wLU8lv8gwZpkaQbMb8zhYopcxUHitgMt
8ZC9AlAgfMbeQ0KeZqpmNct+Xh+8GQoBEs61rj3erECg8ns0txBEvWd+1P6WGIV7
+XL+WQLOfJZq+yatBlxZu3VDHmQ29PKCEJ+3uua8l0MTDD6GPVdNha6tK5SlwNWM
NX8dRGKSUEDpuefo5JPYqz9GxyAVs5Y3pkXm0DGIuI420fru+UyyoFgUT2pERwJP
oNg2LFgLZ+OYa/5rhVwITP259yxjaenEHDzeHeFrq2OEtxRfLpw7bmJpEH5IEKxu
Sgk3k+Y0t2mjGF9aXFr+fBp73VtFyHB/SV1SyM1wi01w5C2gwLNswOpdCGV6IO43
owSWIrSLMO/3x46BcgqkPxDxJRo2hKiVWkRY7f+tJ0SbpFkh85vClAXO0gLlSF8S
SD1MUHPtB+A/getYhBuIEYusPA7ykHXmw62liYa/k0OGqLSUELiqf2HDAtA1g80i
F1fVRDDeu7f1sKAzhdxA6KsR3uvg2MdlC0pyffhKSElczw2ARiVnhJ+8HXuzUm4n
Wt7idCrcvkF58LluhMHl3U2qbL0FNE+z+BOHFhv3o/IpeJjyi49IDbTkDo5zq9DY
nHtyDo5M5n1K5A+/bTL6EAjbRpP5OuuBRTmdHwZ4yzcqA+H4I+DdkKorMPXVracz
eTSD13EpAscN9VwHC05VclJkee4/wtC/h01lGR9QtZWpjM7iLRdJfKChyl7KWak6
XNo0CR6vlahT4H11vDBo/mJTHYH7b2gitjqWlaTHzzXaUP0wG+bDPkwy32MqikaG
7XKysxDXZPjQR1hhua7LC1IDOTliPNeIxH3172fCSbCdj4a9bpPIz7usclxNqYVC
gZojD1O5FpqX29HWVtddSHNAWtDQ+bvY+9KVUVCUR9ugsu7SunMAqkTPEqKGOqT/
l2qAg6B0JJqPq44pdgUwB7uG9KN8DzJf7nOtCeWauJMyD4GVMrlQ2JO4/sGoR9hn
XfcROMEyWk049jDTDzquh14wHC/Xov+QI87Dw7JgiyNJKOnNmRoUL8kjCJpZil/w
rpSp3w5gPtBVefFVORWVeL8I8+UXfJEi8X85UXmeYJI/6q9yyteX0ImTkQyqa+Hl
qzqWUw7ue6Sf5CG9DLKIqGmg0sSG2shwmOYTK48KpzmO8yW9RWfNCNb6o0x3l0pY
Zl3pxQ9K6UZA53psDX267KUlj9ocaN4fOclZPbrymFA6EjGfFL8gv8dB2Te2eOXb
3SfsHobYOPAtts1TQJGaQVD+KLQPUjI55Ea+EezsS6sfKjKZHUJGeYG8+fvnsmyC
SNfrfS1t2PTEqnBJJ+yNw06lWffzRThNX4Ugz4texd6642zDpyng59/SmpGQrkDC
HeDzacNAu/39AsgWDzt141Tli1tDF3icL7ExoGMpSRA/AaV6lShe0KMUeArbWzbE
bm8HKssancJUJ4/Md/ewTZFog+Xga2uNmtPGzomLmvuQN4Xah2kaNJvgWGKS3oH4
AgMPhsjnMARXNtAgUKb/vOZuVRTHR8G16SLMr/lo8nO0iBr2ukFg/OqhyPQUrzL4
DAzfWvG/ub8jPXccdaqZIkE0XBsrcYnqY4VPIsSzOgqbbWe59zEKbDn04bX4oa8N
T6NG78pvxByLWcAffZ1AZCIXO6uxmMqJbpv5dxEoLGZjK4/miTPXq/IrKzXtnWlJ
kCvIC4cZWoKTZg0Y7ukDtCp5mjfi8f/8yuKpg3A0aG8LQCmwpHt1Lh/MSN560Sgu
ugymtllM1Si4reswvto90vDe8vE6zTufi4KWB3kAj2Cfcd+IYgf7VhpXy6y/Kf4s
DEmhMZC+0UI1E5j+1UyZcqb2DvBPKI9KnSNie5/qFTUzfBXCUvNDw9R0qQnCIVW7
n3BU0xOq5QxvDD/m95wYnzXjYZEA6u8K8YPbRKen4JY8ceGVX4lZ1O/Os7/3JvuR
DMf0ddJXqMNP99XuK7ELix1/4XTU3zOkWv6KJbaWz0Bi4njkNm4IQi7qwj5pbfwy
GzUwf0CIHdItPlf4vRZbUZ+fQpxV2eJ/oCEs5D8gs3orfgMzpR5FxuPVO7S7WdLc
ysHRsSkk0HxCCzyVJnL42RgDte2c1w6F6XT5yT4bqmRBntHBWk2gfPzjubVrx3sm
4YTSCgpPcEkwFVEIQ0IKfVGvSiENt68RLxQreqbX3moQ2toVltCFu4SGd7iqSwQ1
6mYO5xsJUc0lQsIIdJxQbLuZrl3e2FgwhtgcrjEztVX0BvuGXO1TMZ+FbmNWwIBc
wljIl4k6TPcStqhHBA3mxF0K/0UuDfPXJ8W/PpPTny9j4RM8ZrJJBk07Oykt1jT3
38BLaOCPwXlx8vi2wzjfiVTHclhk5vEEV/cbyF93kBakdQ0Q0+KuzRARZexrD9Qd
Je+/wJSYxB2e+CQMiF1Af9deu+Pk6jgbS347eMg5DBk8ytBF0pvIT2PQa7AuqTKy
ngT5NE45RycH8djoVn5Blykb4wuaAatXkxWCt0aU/FIiXjRq00tuC977k5AV5NWB
PDIbDBxDGY80ZXzaNptFQaj6ayS6tK5PI76P0RYBhp5udx2mI3F8W61b5Dqs8YpX
aGodzg3oCNBwWFr8AVWwvp2agHMG9lAi2NkbociUA/owVfMNstxYsvW1mCd8QsFL
uXGiNapsEWdrPU/E3z4/ip0kpT+Tc+ORsgwc6ROuNj+YBHpB064i/RK7gV7i/O53
emYsMT7iquv/YaYogF32S4iFlHM/uDXwGqRX6PD4PCfsTIc4hLKCFK3AT/w/jW7q
im3LyedfzfH7ic2X8E6lYK2DpcD5k/kNtj+/tjOs2TiuHb5v5VJSWucMrlizcPXb
IEk+m+2S5pyVJKrFfb6PYwmV9uv98NQ2tl07H84qQtC6bLdsmfdlYjMinj4y2KU8
g7fTPOQDpsFZ7p37okoMPkktk3/Sd8KphxJISY50JSYVfl2wNdNXYkxOiveNb277
/CuxGjaya8EUHrxRQBFlcTSXv6OJuRK3rfMe8Ed4gltUQF+MXK4KWLCWrYrYLc6h
FrT6F45u+40BC/E6ZmPKpH/2AUcSl8Gdcfzwryb/sPWbUtA6Jev9nT/hbK5xcYA2
EHnABKYVx6XCvbUvhb+BjqWZLpE2KDnAFzGcUrMIGjWc1jIKF5BpBqru1qFH69wW
8+IvRa5kJ+R4O8q+jJ2WYtyGJmUpUngG0T+r+IeLH4ojHCnLK9SvDLuYXysO3uv5
4/XoDwe/iKCHMY8Byz0shHvgdwkpIr/Oc9nSKvEGej2Bqx2VXycH+7f6+mzaAd3g
E9taU4N6Bu42MaRvyJcc7x5Q3QaWjDVZx+18eBGb/LbWjITeuyZDtTgltkhQ8snz
sKQSpJQsx4QgsLJamUI3epgMmubs6HqL77NaLSMUrV0ZJ/pqXm0e+nA1ktGqraiV
ZlxsQ6ZdE54gDtWTjJGMeLzLMkW10PWM5k4+LU680AfNdZp/ilvJwhfZldqnPDWH
vQh19Xv8l+q0NoZ09Wdaa6NqPyXeVRK7eq9IAy5q21jIauFo+7eRlLTxe4Ucf4On
58C/sjMhB/1NG9nifs4lQN24JKFUY03R9P0YKDseNwm1PY7jLbZezRLX/6lO7yyL
J1AlE1R9sPhDVFfmot755g3JrjNN6E/DKLv2PEjrQobk0XanxsY7Zmswik1kXBDz
VkLsI1HIMGkTDM17Dlobupw58FQPPTAsHRBS1FL4eM0tqDNqmyixM8ph2I9106D2
Qnas0hvFobBclKSCg3m+X3GTRrOzPqPH3mfVlCtfNTB/SgeM6WrRvD98LICj+N8r
u0QiqpsVvqqH4pfvGMdptqGtjF+XLjR9WOF6n7/JpT6KSPEn3NUUJ6+oItQZnxQN
WIGrUr/wXRvip7HIiuL923Y35+u+DZvMnl6kS4gXL0wt/Xlzr/k3aROw9U8s64FF
/1goVw7ueQ+jnR0I7IQnFStue/E0GKmLuioNwrwdoRMDhmivgR7PZ+wLamRccIhI
2HO42AahZDtuuByIqucLYE0ueg/wiCj/doAq0xUk4B3WAVoBbyGRc77vMNFGWKeX
RxuInvjnSetKAxn2em4dmNsWk2UBn9of9bHCnU4wXlWUyqLxsUxKjZbB9qWRL80P
JS//qf193ZNbmJ9sxM1uxBLOVZXKEhJ4TuRk0nX7HKhZo/a4t0ifqY4JWn/NcWPa
89xJZnRj0hpfY4VtNX7esTxSREe9nAHY4RdOumI6WCYhnO/cMi3XMOH7E/H8ORmJ
UKLg2eVBTDbWitcKqdeRVhd3BRO4ObgGTytVKoy8mrT5JOtz7ayDnH6ljV6uT4qY
vQjE2jPtbXFtrLKPIFA+H64wfv7kK+UW27Ven8SThomuS8R4Ozpfms7gHjQdf3Ky
tlPHsdnC1+c4b3IAzBonYI1QZ168rWy+Yr/nZGwRADhkeX4OCGlfxp5fUd8DNZMD
01K//MZkTbfPFn1xgHpqtkjlRecqZlH9ecCATOw9askKYR6YmDpQMi3vDuyL4AAs
dHqUWRsr29EARAAb07PvQcpacylJFmQB+V+VEKDHB+EgNXJOXWkdsd6YklwWmD5a
fMUyxZWdUOGNEgqBY6gqYN4ubMZukjEwrwttW4Ip7IGGhzK6UvF8B1mFJ4aF3P0i
uEIPDRJZE31TzZxP+RDjalQfzPaigG78h+Iu4mNb5lzjnrQPTW2v0hLYGaeOqPZE
FWvSKPnsquvNisVaaZqu0KWt/ilvOaT58SoYq5N6yp7Qkp+rgGEBFZBpiCzKcPq9
mYF16Iri8mon/am9HrouLSpQvLKANZDXSOR+xk3T+69bLSe9pNICVLUSbymzm4v3
RPUgZ0OgWz21hct9B0XXCQQqw9JyQISI3txaUVslxvIMYvKvNYsp3kfwLuyFBbtI
WU5kHQJ2FJCB/0WMVW7sduidrM4+EIOb+7MKmMancExyJumymmd228//hrk+CQ0G
WUlxmtSrsw2WBZg6her53wswkTlvNnazQL/4ZL5ycDAOpPWd1sDas3q8mcVsDD26
6Epf1JsqIzvjZ//dY9uYVe2NYK+ymep9aoyE/7TDX2HTdpt8vrYF4xmAKkSRVEao
2KN8093Tlyt/wUJs4pZL9minGxcqmLJXXElOEWOQwnr4Bvy69RqRHIeFo9hqtqZB
6i25Kj/9vy7nRt6+dvoWjbS4jOoT6ulviW+MVdSm32d1/ga+qCuSnbrhsgiAg5sV
QsZ4NM+/vmXvI2Q2Vj7cZZ9Hq0gPslM8Sz/9XGApVaeXj+ChqVjC+Y9ywWlgDR5x
3HtvFajG5DimcSxMWd839ZUORCo2+6PJER8rr7kvzbucw6zcmPmfBDDSP7B8QKvU
ow8aPOG9h/vzCTNg31AN+moA0GmcrE465sd4PBr7naNYnAkeUbHzRXwSGFDgMUpg
BUT8bHlwimhWk5/SJZqr3MDcNH7FaVuDcHXJ15DG88u/y9Dh44FcaZ0K82ACAjQH
2pAqy+rhM2lY+n17UsDu2YX/MMFMxLEpop678hCipUo9F+MxSpfDLJcdukapxTB2
N4g1Yji6NyqNPUqSRuCCwHazdV/9d3zivkRcqCwwV2uEFJMSmSm6CjSH+A4vMQqW
EfYQTpkHuoLv3W95ImCFJ/Lz/1ng36GY0oIsqx0RWCnjCncJEE7OYRekhhQQqphX
e9U1iVtdTYasUAzzlpIcDbNP3vlF5/eUsGFSe61MVUFELnToPHdaWtWOZzaD1gwl
WliyYfTHu9sRcQdWT/TotC9A4AMbpN2MTLSNqE5dlHKa8YTWsXLe2YyBreg8awXO
0kzJ/Hl2jc+nK/WqqrdMV0I+80SIGc0/95clp+5gZhlahTBvir8hT2DEASvz59DF
rb8FfBrtVKDCSj6kIEH/58D0W66BLJOIc2xE66OAGE/ofi6lRouyXJ5lVbBiv8NL
NbFxOPgk+dxlLur7imy9EhfuR5rxcD6RDCgefZYe5HW4prfnkqflsr4TWXVJ5nMX
DDZRmSMlF0oQV8vne3VSOxJUJZ3cDdc7XbMy1tqY1W+DZ6OeacegNdSy28KqlnmP
0Ssbjv32JXusZ8i0+i4KCvxvNjg4aRVxEyp7BN45l2Z3W/XT15NRUtp/eIsX/sU5
ypIhZBZ8ROwCpdnGKvmi9/2MrpZibkMkn4gmol8vM+cNzrr4aN1MDonyZfRFNnf9
aexm9e4nSYgYKoMfoPYpoDOK3tPWJVyaNpCB50uI2ViJLV67jnpseMBp0T/Iszhf
ZHqRLqQloDkYm0rrgeHNfu8FgJBP5N8SmmKdO9r8dUFWunFb9Agim6mmHXESaolw
q6zlhLhVuOm5qmcH7Ki5EoUSI0TP37pY5U2fcadLCzERqGOOVMPBLuXHsmVAGwVG
UGGjlKTsqFTi1rly//qHK1DXvaqAE96dAxyIfA5TLpdGIC/jahtWHjKIahj7dOET
xF9j2LyUAp/Nxp9/m5WfnzCBCSuw2hoLDsuUGi+sK/1VpM+Q3jwNzqUekjWbGuNI
5376wBh3IX0m+uZLO+66OarTIC0+COQ4V19gcEJRb/7FSyYWNJKUG7O1YJWYYSsR
bhp3YEn8Q3DWd+qbYZ88Yce9jPXTdR0FFEC+/04UXi0YDdQLCA0rRoxWe3c8QYgd
GUrDxYetb2urGukeOxOk7hY2BDnlSguy7GhyvhHYNLRYDIsNB7c4HixgzCV5LH3C
YqkwpHvmB/j962OV2NyeKu2SwWU+Yh6+12fhqeGUwujMiSeFoagU2qZk4ptNU4sT
SNkGcb7X1ycCmSAy8LwveD9acgMMC3KizxbriUsT3G/yLFfQt7R+W/5fVGeML5XL
adcQWwbG0b6Lr64WatMHgY8jYvqCrhFw09r+I5E2etttBeM5Y1FE7+fCM+e7nPYT
ROZGUmoMdOioBOfqmUrN6Bw7r+wMCRgkFoBmLfRtCRHUQM1faQDu05BgQkbDiG15
r8JY5sHLGJMcDG3m3D05KILKHvzcnkzPUDJE1E6pkwdsL1ENo5HJLiNdc3Om8pPb
oH3pihDKDqN57ntPTJ0Iq53YbHJCMqtkH2lWh07V3I5pQk1IPelSqqM1QHyLFnsV
MRL/zJKfpeYa4g9OEF9yXqDBj+HZcfbGASqwUocay1aElJtZ5mMPTad7QWkxhk9G
PKIL7wrSwXEMXphQfLQ/ZPteEIUL9ruvmiIkZ26k4WvKZKgcPZla8OLk1SFr7VoS
KjJGk9cnJ7eP2STiEWR/jVr7LkKniOPHPnl1+pMBQCABPON5ZbCcLMCV/YifWwZk
A5ABecduCzANetHUxGyoGsc4CG8kvCaqAmCHpNrFqwXSSEqReOzVM2yUVtRWCH3m
KHbOODiV5e6UDxSYigYSPDifvkKS2tSQR2PYfuKQLNne3bJklhShVCkSL56QpjPy
mTdwae80nxldXtoOaxCKEwlfAQrKLbEi9f+P9GDxXQ7u/LSvhs7KknKyOq5WRcJx
NGEPM1pVwit+MM9kJqUl08NZ0Y2xdPiLHFxdicQPEdCI/eZ+chmzXbErw60avJuS
9+XiWbdsVCU1uT75OmDQP6Yq0gQwb5hw0vfARXjHEpMblgDFGirtjniMfrjS1R2r
DfhOpby3T45XjuQuYTPArlDryI+4BeEhx577TvGWIw1d8e0ufxKD+eVqmFCyAIqg
hhHdfOGcT74YL2jO3S+YzFb7HVsu9xN+TvPCmf8t9dUWxAqjdIgoWBxX986HvYyD
dJv7N2Sy8ukbRwlzlzE5aaweg5MUPjTSRLyKrpHbZGdiBgAlK4zdnkYbvJTB8Xwj
8qT754C77mTLRzMyEzTIC+s19b9qfjiuTWPMCTD0ygxwrHs4XdQDfgEuDuJ/exdT
pfmCW8fMSkrVw9wUtPXBWevUbgprLFtxDWxXt/B0PJ8Nix8P0L7f39uHze7xIS6o
a0B6UhR9W2smpdSG1IFFIZrZ+Vuh6+Kb2CrCkMv2/nFmP7Wy+lRaFUIt9nH8gzI/
+Zr5sU4pI5SnwTADwxA0aISTKHFh7O3sPxTuiarEPfqvWWYAHBE91cw/Ps8EIDAB
3Ak3bTbU+z12Z5hdjvTry6MewyEJhaSAf2NFaB0waa31QoSLc+zJ77xEQgXrzA+2
mttA3Ky0ksle7au+2HmELlNJOQjqwHKb3NQ0GwMlqCMgWLjctg+/3/vNKNQenC4x
o6YpFyR5V7QgHz23O+R9SZTypVcPkU+OiIr7KiRYjn8wTs2JWxJOG1NyNE/tX3bD
4Uamahhg2CgsJdUoXlciD664gN3HeE0MungEko3dXEI3iTjroz4OCtH+dn/YdP50
Grqk5dIYSOMbQmVmatdvtXmmQPub4SKr231DIKq70baWy4mwysbAazgjkij9c5XQ
D75i5YfZv2d+vF8WKkLRIdAU/wNolf1idXA+kG8Qx8hw7CdNM5Pfklpv/Kqx4tng
lUWi2a7JztE29D5TFuiNP/m4w1xz6vUIL3LjZoh+injPBVL7ZbwhzbeZpXvOrU/R
P8DNjT3M79kV9J+ktxFEc8NOWCZGaZPUV7JrUH464AH2IcrDKIsMGbfhT4fQwZp1
i8SVkVqYt8RDFlHYuid3XTquE3g5YyTvHOAXtekc9tNYx+bBogkgP5TaXXVlD13L
BzqHouleDhNQ3MIn5RlzVsFIWx2jyuOM9DDqGqWrbPSaBxsNLdEIHQ5xZj8aTY32
2jtqFnvFxZchCfwkBlIU+Wrjeofbxm4CRou6XRUE1AqqAL7oFaDSiz0sQLqAeih8
q5Py7q0R+fK/mXjXO5TnoQmvYIG2yGCVT39B2By1YMTEZHPCT53myE+miF/AdwjV
sFsVkn9gf2bAPEuD4+/G11einh8/ewLFKohe20lLv8Bmk6rHxudI4ej82DvtDOhp
DN4t3yctwdPMeQR8POWGNYAI68BE5ywmSFWMr5hG5YmgwO8a3l2UXJ8PJHVGCJml
Tb9gtDw43zbeH/o/3mtbpFM0V5K082PKs+h1eI2riVvJSFiVHpZApHyE0vnHV+wg
gQvFfDyGtwZ+MCPYMWLKQEeXDf4NlYZUKn4q9rogxsOdtgutwnBDtYqb2qgS2p1w
5pFb4zv4Y3wqzvEsYVMj3Jez88jOLN2XSM2JVD4K1VgwoWCjxNRJaedVg8jaFOTZ
zfszSrEXbuN4XXNWmphNZQSmvEgrU6jtkJQLpYAHy+QJYZludemBhXs9KzoyQmkK
+lvcisz0fWYhhhL31zopwZ5m7uG+qHB1iqXUSv0+x1n04Lx51gIxYUY3P0dhayZi
29TqHPtgGegSFefYjdaSE0D3FXAgPDMu1FbqrcFQ7saa+5XwTGsQOssv4uHA0YYK
nAaycp1bHYsHxHttA/JELvMYObXDOq2g3I283lr/GPLE1gf9hWQ8iaPJ2T+NQMdO
/5uCf47k1hjo4LjjcBEB3YLKwofQjFeMcftidUhiQx+AYp6AroHEs5tqUnC7YzOt
kIbZ6CVwXnqE70zksrKBnV5qyPgt90LFnSPLcrCgqWHZYAOblj7aXJPVw0l0p6Ae
E3KCgljnJjLf/nKxUxv+cT/oZWvkVVSSbdpqIfhgcj0v2215q3Lkc9aypcd+vX38
JE+Jfpr6uhrmNUialwKXy0MyBNzfBE7dUhCdf27iGK5XIJKRVfrnHIW75u8XQP10
CeGCZZW7S++qgiFKc7QKRo62q1TWfqieEhARSctMWf2i3KtcvOPx1kxhRcvu+CN7
E2oFNXdIroEtceFdYdCt8KU49x3gBAXxvp2BSpfHMXYzwYzWYfmyON72w6qQC7qx
6PSiq1TcDnzjGbwr8LU4xTgfVszeFWsWrqV3kxvS1ZuAS9gAlHrXuZwVnx4/oI41
MmuJVQbh0pipiwllfl4fYsQb0WyEZi/0qvDr/8RouwJm8hkIZ6EngAZ9w31uvapb
NK12m8rCQYIi+6ZWYeJjNPnrBAnaBBaT2RDDLkQxzXmos1IHRRv9ZEV44k+zMGxX
kjT/nFtrmpXLkwyVRCc3Nd87jxtNQol8roYqOdpntJ8ZFi+q7AjeM84OzvRZsgY/
+/PCT/97A6g5PEr+P2GcnocwM+ttiqKclqB8h7OSpCY03NpiCeHg0Dl9KJT8ITpn
pbdCsR6v0WVPxudQFfEnTRlVlhOCFfqv9pPkzcqLyYPEUDQsJrzc96bJxE+voQca
BBBaDPGrWJHEd13iFRpoTs4OvmUWQ38utl0b8c5Cl7JGUDKAL65FY64+g9ZAUSfC
l0bqVUZIIcMgCEvZK9SeIkA5dU4jCVk0hK3f5gJdT+UL6ftjcrhguCOWSFPP4QO3
M+BxsrG26sNQOb5kzGOvmgOR20ynK0Eq30r8cwkRKE0/1drs3ADqM9YCdmP7DAiW
XdsYLWTjSe+b5rSb/c1sIXaKQD+iYBa5+p4XUMusRu3gcIM8Ht1J2ndg03eIoYVX
UVYCn5iMlfzFrTdvTe6Ao+JVA5gGWFbgd7XhAivRoyXsAWd+x9tsyFnJYsbi1rvG
cBD4mUGCrlbOfkQmRgCyg1rgyt7MHQZX2nf+Q83vG1CxdC7kwmdNnxJ2FicJcEic
iAL6TbxlpYWXaiymt9p92RahstZ4IYQLMsCOqA0h0ItMlyYK8LKLUiO36M5KR3s6
PkkndVBAg+DWSH8WWcKn2UrC8LDZNsm4Df+Z0jSyjwUVSxzrJtxRy0sjJ+aSfAMb
jDyNqMoaiAj3KZtH52jjFYslg2R3vuPKKqvuuUr+PYdCgJh0YkT6lgBuybkA9VkH
/F3VHP28um5gdca+FUJ1D4p7UWlG3Dhp4UW2/DL0IZbBKSFQ1yJ73Sb8Uv4rhTy4
7WJFgmKdLleM6Q72VnIbZl7FnAD8OE4wgwyiipl1iiK4hLp9/QlxZhV0j/Wx0qbj
guFytbbvNxvwB22VlKVBl/E260j9Fj4N2rJYUPw34sBXO8OJDdt4JyRw2ODGDj9R
+w+lVuu8D9frQbuUukk79PzJHcmoUXmNPyNGTNd7UnCwdvwpR1zTmxHVNPXtez5I
XuylpMY0L5JjSW3KdjnwLjspZCj+8218OvrmCerfuBtAhv/1eBNNk9OTGoTu1R2x
ymR8uXY92njUYN9cdSX33trvOxWo7e2tf2IIsNnp0jSNJ4+H5b0s7KbAoZ8Tq67/
ZIhF3N3ndcvbYX+Ju0jrNxJwva3ZHiiMDr7Mba5Q/tQR6A5fnqL2wDtOLvVJDvW+
7HzCvP9VtzMIXUVMabLiDw9rcWOWLxR52lt/R2ofGOJSUu/dvPv0Nh3F2eEcP131
RnBnovc5zEB/+6earFYoDI6wW7A+j1EmD4Bpm6Nua1qvtKorrabhgX1fZuGqNU1q
aXw1Tm8yAyolDo3myHktjutTPeW0kWPujN2tUUaiwgpf2J14h7XSAUIBCDSse+7r
VqdKecjAt5BtdmhR5wXDr3IFlxs3Rc70idtk0vqPdmy+0R0wuFutXAsnciM69rIM
YaPIqY6bdabl7xuOshXD68q4q2F+Yj+lSaLA9dphgfkljVAABP7nZBkjR+GvasdE
vWN11VzfGWpaMtqgGv/BZlSODVm/S3JADfU91LbOah6Vu1XX7xZvPnoYGVt3ivhZ
9sDGpJ4Y9GVrOg5TfpY4p2525mxsVjHQyO7GdQqnh8UWYtybQ2LRgN9wl4tjOKqj
9snOaN7rAIJDfpMKUejMoxTCfg+gcrFlurzYXzpWtUB+xf781LCKM1oFHoXHYLZL
i1vMLE5Ku51U35+mKhC094rA4OTsba+fsc2JyWYc4Ht8MM8151ROJXZxdV4hBwT+
7OnNiZDeaX8r1rOj0dowgezfmAJbVJYUTFhBFI/EwZaSeBg1PTUZiYXHfwP9Kaof
vcpF5ZbljRLHBygkqVNNnHC5kJv62d4Q99mBxzUetHGcfG7H6M6IBwJDEDAD01Gq
hPztiMiLHbSLBr3ZJ7DzrQhFXOI61s2pWyux7am+f7T0sHxb5ln+TZ4sKnZr31BK
xbTXkusCq/kZuo9kU+lMtH6UYhp9miKp3C17ejSCc97oauXr+k1VrV0iys38/nbP
nfBEO0NaAWGoUKGsyRB1lU8RmL4PR4560L02iVu1/sC2+icJtF2bpam+tnvV5Ht8
OClhlCmBbl+3AWAykk+mV2xFAa+dMgXj1VY0WpW7e+NfJ3OT+yn/GQCWu9L8ZyAU
zERzvr1vGf98bEdcMrPIBgG6uS2LQr+FtiFlC0jQmHH7Z5+nL4vTrRYFApXBduof
GXhtaQC/Ydezl4tvl8XETL1tUxendCYQQD20/h+GHlJYQ/+rX70mf0a1vLNIkFTS
5CCyv4mYiG6stiUVvybNxtwsY3gh9VofXolUoRgedBTVDrycRUCI+/Lju28YzCUh
4ORJSCLwRNLOewPmxB8KassupdO6kQDBTUYAD/zpcP6HufWw76aTBCdq53flPUjz
/1ZzLhxbRKo5jiOzzRg5LLr3UUiMPm0ct7F4FM1TIFKVXsAw+VRDYRco1PRggGKI
UKW3YU45aCA2HH0ws6hKx+CKeFrcn0qROExOMi1dFaI2kVeQsnZ+n6Jyu+lAnOTB
rTvCANNWi3+HmF7yE74/+yKPxRO+a2SZLlgY78EoZGbTryciWb4u39S0iy1HKmL6
p1OwzloskEaoCYg22G/xKD0Z0yL4xzZYkAq3T/RNLXZwkA/V5BwiW8nPJTEy5iqp
ba7GJPxC8kXKsO916jM03O9O4pqv/xpARJ+H5ayCQeoZPcY+E5o4laAiPuB5T0mk
su5ZCfknR9uSCYmKQf+KSQJ6v5hxKSalBrCHLNNuFbu8uMkD3OpTSeoJ1o1CeKb+
M0g3jJoGI8Yb9NUY8zE8BSKaRmTcDrU+vwDaMQH/OtZVx+IcQqbgz/FA+HlyIfMg
NwL7LNmcni4PqLHPypddUkXhZ4TaPYLzxp4YwurhsHmM6dtAwSGQd8InoLw9cAtv
KSxkh1loD3+dc4+r7yOkhKR770B8ZXs0hqb7UDE+S1+yFtSIwGic1IurtXcakFNc
0XQZMsMSN/eslNodNor6KI6h2JgAAjPr3JBpFVBbCrBg8k7nJPrFD+vj7DwadDu2
EtiR1xqp3oeiuqRL6UnNh4dLt6Anv0dtwYhL7ZCVar+8X8Nw1evEU3aAu4beuePD
e1tDQwYx969TbGDn3EZmLs+KmVf3RWAVOb6zXBwHxPSh4zgjjqj/5ovOt0ltJTHM
iy6JG2bzAbpujvrffhv34W/6T6MkBW6nOsjGdBCcl8N3/aXCvSrM9nbsnGuSGi+k
5WeCH+fSZlCg3cxDCbGd7dgrNWkrKE278fYh/MsIVZ/b9n3p5GoTuyx3ldZQdcZL
sqjFcomx38gDCt708I+dYsDbJmt6jM6JsqyFEs+4E4Po71U0Xdqy1nJRlEP0KoE4
wNQsoRgt58otC+I8mEaBUQvP/9XA+FUbxti3CCrxI//MLMoeY+Ujd/i1ulNnkM7y
qzyYk9aMhO7/zoeNGAPZiwBnkcU1II2izPWCgn3Ch5/KkRrfLNNMh7mQckXJeDQm
ptA/L8kYfyCRCep3QEcCv9X8Y7k6Cv0qtlKaeZnGLNPXue+Rv6ITFR2GSpfnqXxq
zfq2Y4KBPCDbbVYZMTAPuQaOEhZZtv942KrvXIGIppot5IwZngiQ578JszWAt/wV
oK1vs38fAIAjerkboHYX3fJEvHqcfn07psJ5idxXcm+GMfieiZbOnoPKTjH6EsIq
OgofPrpDxDML2OIsKtvuQA4HTUUumWRbP+r6RZGO3Lix/1zxbLJfZXJt7BFK0pci
UZOl0PVRa0aROHcj04zW3XFTSqRoHC/4PdYJjMXJVvTcmz2kiP4PLLUVQcFPojIC
c8y2KQqxHwFID+PMFKa1slWvH19SdJtkuIy4uT4Rqd0T3KcMmJXaRDIcndwhVksI
8Y3M+beEOxR2Z2GqTl9eHgQg/w5RMbGp7mbe/EsIKvIsM/fKwn770cekKl/I9HEH
eAyvab980IiCncuN7s3A0exspM3or8FeSeQDC1uxrKU3vFwiYak3pd19kKtVt1Cq
wEqWTYkJJ4vXS7gUenPt+UaBtDa/0qzNubBoK6TZkEEpaxs+hSN7vse1RbTNVvxh
ANn4nhsVfq121mqWilLvgdebMSszMM2lY27RhG7j0l1CGq31PJ0/gA61m42c7xex
N5tDi0EKcY2U8tdKfGtarmSBz+GpoHC8lVosnvLlVErz7xJWP4r+pVZ2nBreYmP4
giDl6xunzHOH8YguoK/MjrFrIbtc/+4yTNHWSssyWdObd+OlEvn78h6rvJJO3IPy
b5CRHXqQ18yqPAH6IqRAev2s13qHY3cIcOz9E7aehQBCthWhw5/sro0jDG04xiRd
igW+sdWFlMv8NgNh80Pq0QJQMIvma38BJfnPb+5xRfA9J+0O6cGu6BN8WOe63w7+
ijrK6JixS4u5qi4H4Kl1SMkxk7ytLTEN9EPLgqtxBedx1Qn1Bn9mNxO7GoyMCRDs
PjsNXJqXxKzjKxPXoUrwifP/AV7w8zQk9Fvtut6/w41DuJRtXp1iuhHcwpjgx+tO
6hynApTDhsUcKEE1jLBkuXRNy1H5CpxUkFrX5UOlyicp7zKDzTm6tmzBRwhcbmGp
9Hg9VbYNy65NPvitbKZ8XmxZeawMXDPVUPHyEGDpL/LhAL+BorYJhGjukPX5IBEK
q6NydBNvO+p2V5w4od2SYDmTcz7tQEvniv3ssOZBATjtsLhQjtDj5ObcNXuoXbup
8DeAhBMq59VM+wjRHUVgXecHzpNnYM/R9Vo7TxgijOvMjKPLyr5HvYI8LEMylD97
FIYu9r10Dg9+PDpm0Glo0Hog0aWgYuK163sz8YTGLe6oh7EwbC/Ph1QGS5Lp1U64
uuxP9+3W7VlwzhDf6UGNbQIeHbIqCeMecTCETckILdx/6E6eRJzMsCFkvzn7xSuy
cJkfmabmL+cLoLH/stxMU6pdcyj4w58Jn0EO1SPRuDdiuVILyiTbP8jdBUsNX1sh
ZApkqvck47hrnXRKv+5U+d0EzzZqcyuZ8DUAHLzPW9JriCWL9U+fE5+A4FfnkVsJ
o3s32K780X60W7lZ2S+9PYd1yMhT0Pg+trYJ+mnSvOhJbiy9BolqJnhcvBwWtnYV
IjyqwgONmpns6Av7Oc/4vVKH4xSA88yOjQpjT4BbpDiDgf51M2SBq36QQsCPc4BA
rGcC/HMFDzv38Omvis4QhVuvA0xH+jzDQdreOGiYMzGOIHz1fdB0YvLZQEaLOJ4e
TSjQy8IMqIeVoavbM+dgWy8aHDCmXTYacXoNoQL6x7xmK7+xG9PRjn7Od4Ua7tBn
qOnUYIEvePK/xXsag2H4botIODssYuRadGmMiev757fbwZbATYw5f/aXYR86KHM4
JoQNoS401kr4bQmj13qe6SCkGlbeQsiH4v4ztlGhyaKF0jsRr+BqQkBGA/im9px8
p5BetwontZZFOOLM0q6KzkTApVt5U6po9HPwiaJ0OlO8D1OcVbOW9hVLHeOZ52GQ
6WZyHOmF8FfEeNIGEuj1V2Mj8IScpmjtgxzz1Hp+HGsvjtZnHpRp9+LaxuZUDYfE
gMmqSxoWn3jeY9WXfLyiWcHsQVajVWBdgWnLfssJ9y/5GfK6VoKhEqG2aPGQUevc
r3W5K6LzpHNnazxmGLnt30RD9vuMTtZpLVR19OzrPxIrtK1GPdn+owy8+HBvfhKM
AJnf6BBgIQF8G6QYXCa5xEyetmy+UDTOFWDQMQzjVNikOsiZcm40kjcTe+HcaR1E
+C5+WlanthHHSyu56XuBc/I2cyhNrFaSWarOC+9fpjZnz19rruQi0mK865gDJav/
Kw3h73H+nrpJr9R7AgdC0oHnhOCV9ZYVVyVlTy1rIzVWFPUO9KyX78sGTEQJqc7L
585YJQ2GPHp6FbYB5pmTLrCZxHO1Hw6srMYr5uCaTOmTjKirsJ/VoyPAAkHsPJ+I
pYd0dFWjdDim3aIvd1J41wsM1KqppaDGp4JcKWoj3G3wfdm1gY+IJBWQGGqwCOaj
+fWuGAzBv6OcgIfF3IK7m945mlCy/IaQq2TQrw4ryUOJPAYSz7It+YMDbCD+xxbz
RB84uWipm33ZECXcMwu6SDy3YGVSN0g/RT5WIC2UCHe2gl+NoVwKOLZdNtSe0rq+
Q2djcAQlWAupfKauQ3yiMrrtgfiVqAFQv5Am8jQVqOzEHmN8FRqoD8l8iAEsA3NL
8rfGynu9964btTRJMyxPoDeECoydyqjpkMNUr7ezs5TiWyQShXGcjP9GYDVUSUmr
tfFg5dhROq97zi0Abclj/vWS/UDh/46I5Htexy+6/0cto8rT6zeH+nzkGhobXg5S
2vuP9XjdfREFbJiaGAeQJBg0ReSefX2z5foC5+QXY5mMqtEl/H0TRgnVUsLgMbGk
VcqKHHl76zQMaIRp9gjaGsbR/RUyiPIRm7/py6NHQSiakPF1shP2r4OyXZ1Hn1mj
yPN7chsqX3puM6K5k41nwP2pcG0I161NKJ29Pwy1jWGO0xbe6fjOtH0KBfE480gY
clsPFw1C7k+kWq5lyAW2VwlRDClCW/SqkQXU+/twxoyNl9OAJtuVWEj6eXrx+OO2
GFgfsjOPO35RRpG8mujIr3avvY3SX4G8rs/stE0rydRuXaWjc8HBK6/fXkzCC+3i
pOwJwNw/0ortbzExb4l0KpyGM5oWRnk2FC6JhI1UoGZzIJfTr5Hhg7qq2bsIsR7T
jOYcovP1xFCaETBniDssk3sQUtRO3FgA2V7O3MSOyesgymyMnLRfau9Mbuon+rPp
kqFwJ9FkU/yysRi2jbSFgxhWgnCRR3pf/wppoPsgqNjXMhECTV8mSMwhVEtXuR+6
HAu73SlcqRY1bZrO6gPQLe6rwofvVlgNTstSeQJvZ2GXTOzdXUgnjNvITEx8KNfO
7yUI3NDtbbHaL/3nrMjjCSZDaZOtPTJPHTpMps5+CRXZyD/fezwdDOkKpDVRREZq
IvDJko9fTJpTt+v8ZVB5bBods3psmy2A04QF6kTrb6L2eOQaIlSxhYBqseW9IBhn
oYrLP1fB8aaEjWwdNt/OTIYkDfKi9ejFLLKiGvZ7Bf9/cJVTKGtMDRcBmumX2yV/
A1pQG4wzD8mLZrKuCn1Scr26bWmemXUz1/8SLmbltAfna3jLUfrGSdXHRszgyvFF
giBd6T1Cyv5JWv0ih0i8lr0OpKtfSXNSSInrwG2BYVlCRSG3UZKrWCVor/AVqdwZ
ZZfRNLdbtZLPfd7VfldgIjE2BVhYuUx/+JDv8qMVvJSjQuKQkZg8AHjoztrkViys
O4RRwt5z/Xox4deEqGZtXJsp2+Dso0Re0zZpa4IqsO15dTYB3vlTGHaIHbE8XToQ
dRLvZF433X/lw1OK88HTyabLG6/Xd+RpBzjn6Sd5sOLTrXg+DKrBh+22cVRQCAkj
eIjTKFnFT2kdcHdGa0zIaDurnCn40MUkT2sAMu2dsLfTgXobGEne74zryiFT7/kt
m2BLpyXEQthpfXLRqUcRj5ib8onhsQl54lh6cIFKGGtZ/1KsqlERIKQKWmc/ijVg
UtMYHFhNHIgADZ92gRlbIV026++zTHukR9/ifABj6dtm0zHlAx3LRpjSa70SVK6v
VgtD1XBNHLI6P9a0/ph2iQ120ZphesBKGya14vxlAWHu0oumN+PHFTNkUUEfxlM1
KgODpkRY9K9n/Hz4c1inN0E0Vq6oa5hITOeUYwyPcvoNBc+Hw6r28NJSO85quCt+
/iP0e4vgw/Q9EJKpQ7yr4N9OdA4TTwoox97E5qg5K8SrkdprfZl6kC97X/kiWisf
cY9dQ5v1hbPWyuwm6I5ZSEk8ar+ZA9pFurQQJI3GcBgjZBlmfTc7oqE5KbddaZ0p
J5a7ZvB7b0AAKuhOmTKsmPRqtVOh1Vr3RyNwLlOvQCyunJebjFdUVWKaT8Dli7r5
WS8Wga9NJck2gCvXL8o7BcEqIy5pe0RHljvQ/RPxYUYTJlQvHhNJT4SITFpStCv7
7NTFnQncryOueiSHJWNizzQwEJCMaQZM2MHTmMvIEd9LxhH27Z3Gw1YAb5pP7vbS
P0MKCtm5cOAmERGQYycw2bOiuYMDLiiMnkVez2NxLRGPgDeuhprhLBd+jkMPH9av
2PxKBRSWVB36WZHVheXekUjRfB+qoyTu9q6GDbEZtR/lx4KaSak/rhbtDwjtVcMn
j8ErpI+Ey/IcSt9kxMqgcUQOoyUETl5qLy+ZpqtOC6Pd1P5FuRG46SFGHc8N8RUo
h3FHrbg8I3MEtU2ggzDLeBlbkBYpJYFOPuSZs3HEGZ2UeXWKWc5exY79HVwd6vtv
+jBUBo4Y9XqOooeTFLaih7kQnutFgsR+mYgfv35buP7Uaws5NBqzwWJqCecdLrRt
rujeRH4qesfTrMNELOzz2Q8f+jbFhnT9zD3r2jfWQdI3RHcD/NL4DO7fRuj5rjAA
66CEhYEKO16tm8QWdPUabiWNJYQTkBnZUAnekdjQh+n6ISCpue2mesa4XBVEh6DC
Hn1gWloBAYhVz47zB9hDXx0HXSAPZDLSNMdI8T/cepw0EhdErn3NGa6VF1gZHPwL
aB3lhBTMzTWKwwrHX77dn+w9rJZODWboNQkXWdMzYzJ+NGHCMDzQ+Oz2kxPGoWjA
KpiCAemZvUux6OcS0+urK/4ihcSbrk4wEaR3J1I0kBKmzMMI8cStKKyChnZORNhB
3SFYnYPuDH7a7dFr20jjbXk0hW9A3cWwLKqQS7uqFHFwiBpFpBevh7QQP4rH13+R
wnjyHjUjpk+6JfMvbL068F3i76OwRhnNFg9wNQjgITIB4ttRAwwIPACwRfc4fMmG
Z0E3PVtZFV46D8R0/SiZoOFWEX4PYvN0qAO1lgVECKSO4tRkW4ANJ12+jbTAFeKD
OZBBWZq7nvZsDBxVa8C5NNRZUaBJ1Fe2CuGyjRIgzHRyxfrOKJH0PNDogSZLDf9j
geMfRra4t0NFRowmlaehz0SVzFbjdSgFwTMQP9ErGosD1kxApEIovwWwy5cmWuVL
zyiPGHty/KPBqqXkBHThGSgc83EZoyhj+K3/j9nEftcLOcBB7Y7Q1LRW3iQ8wpQ1
ChzgU0dHot9KdH24QKu2RKhdXQh9W6jsjD7mbDpskTug/zme+8jSGYwWNcvpizLn
hTl/sq+0RpG664svXOCdFvfxKzqee1eIDwVW65e6vhZ5f/hg6g/bTLc3rdbTiylv
zgX+dZJrUSXB3lNfQpARqfwd89b42KWQPCKsFYgTmwtQKl+obbYrD+aKZnnQ3lq/
zGNmeyCdpDf2HXJFTCVlGaX22Scf7FSb0wvEmliPybQmULCIA974KrH8jYOurXp9
nQ1XEtroky8vNB1+Ri5FkJ8ABxd0Q38dNIztYmWgiT3DWHsdfGMU3e3oxxy88FT0
A7AaxNdKTsU/RJaHL4Dlts7eochC/xq5esUIyAyCQFHyniQTZyOEGcAdVhiyKMNG
CKnPZwSvjIjtaqJLIS8FtCWeJkp2M4eXxmmhuUGRExL7Ws/nIYli5dQ3PS69ENEa
petO9qgnPiL10s3BgrtK/uzAgU050Z1ijnISalqxFyt7FLp+I+hHGtTqj8MKJPGp
zQXE1DW8i/qUkc5eQv+RLCnABidKp+1fQDXwXTGcU4hv7rvBqDJs98VV8UT8fQmx
TKF6AIeNJDcljuBiXlaj1QIUCxchDC2y+IUaa2Rf2PyVs1IB+oZdpekqNX0IMNef
jLMsZCusAN82D+nZ0E/S2Wn/C5uj3uxxTE6t+8s9BnApBfMsVZ2waq/FH7fgxgKn
SKCZ0tXY4mekQID0hO4j1nv3qdfI1yBC6Ln0CBjJYSGH7h3Fu7XF98rp+b0n4Q1R
GKpLHnh1XRlFDhzotGQ3ccQLKKdGlLMDL+BYL9mdrdukrT7NXwS4PqWp+6qvMEgz
+TOIOqe+Mm/bU3EMMF9CQvhaBLCf2gMHFrq0nquPC43AAVh4SeGeKlj7fQ6t/cb+
ecoQCTvK7SxoMpz9oTWyx6TAe+yuxDhuVg8Q8+NHOH8R4T5nARRtzJYe1nRKignB
oQleIQ9RxUgElcJaat/u+ikZXS/u+zMQczzmwQmxNhra4rqq56GXIoxfrHOJ7Iub
e/nzzuBap2zgw/8yL4jGHMVRSybLHztn7UVOfoLyl7QGAn42FXlnmlr5nISYwItT
lVHFEKVYRrS+2UyCiBMJJuBpRgiX0COHTopFRzwDHQZ3vnmwFWBsJ1t74+egshRN
cDb0jl7Qm0+7acFVQITUaKNWJ9HwDWgUcqN8BH3+SYY7U0yFFwkuLPcpKUw+IF7Z
5q23EZuUH/mxqlAwsO7aZFTc7HtMngjJGv2cLRlDNFRK2w1iRS15i4KvXi9rOAsg
dq6Mx2LfKIpIY4BrXMIhBkw+QFfwKVNnMktnJS/IX/50a/sfEVVuZh8BozAcQ1me
/1HRhdGJns+q7P8SpAE9z8TJ4goepTZuwEmXYwQ7VueQ2BFuduL/++y/kVk/efVH
FrrbyCdFrTaeirykq8joOfY8Ore8+BwMk2lRYsBLa65ce33t5ZZGlR08nlEE00jd
CcZjI3+vtCSZM9xgwUv/f4UsndWEep0ghusfrQJ6DiW1K08fL6QoZtUw7A9pT1Od
ExtECpFphN7D1KbytVXUmVo4lUu2LCumoTHc8GEZWYt0nVYwo3ea1aD6qoyjDyi/
s/MdQlGrZLmFV0yL8RJtUATBHCLLQnx8IUhD8OfGD/18TBt2N3Cgi40Yc1sSzMot
UjkaklEdqRVotYFo59ZBJY6ay7a3tRzyE09HniECQnNy7ybbw10bX7fuIBtCjJsd
juPSlpLTlAJ5nbwBr7nOTVYhhrweLH0R0KKdWA7pi+d2gsSDuqrP+65vzModCUlT
kwrcPsyiWNMmK7wG1ZvS1m7Y40HL7L7lMPU5cByF5DPqyT4UtFs18f9o4yjLReIY
7/vAb17KAGyCCseNYBhRGbDxI1i/cf2Qd5OTKANQXXH1zE2YDkgZj94g46yCHbQb
eCxjZbgDCTtioJTrjfG9rNaQpxCm4Ku0ws17t1IK7KlS5zw1s7C8pjSfZXWIa1of
VGHHmrf6INRM3mMMJORWZO6O4xMfVPTqGFPKBKQC9GdQD5Lctw/CIQUp6vHvLxtR
EgYXi0tP73+D1uTIJ8GozGl1uueOOEQ11ibBkiTBcDNZNG7NFzDPL/dHO8e3Zqyo
3N/Tejv2PhMzcxKYM+6rZ+AvR7FTnO27wLpm7LSsPrFavsehnt8AuDnpIWAp0DUi
xCoOpcOozEuRYhsVydUrLIKjKdBRXSENCt3N17ejBr7PeazE5JeVmdgVTTL0O3LV
ukdDnsvlQIzo1tiEeetdpJJ1WlabXs3McPOmDwrO13d69WADROYnjP3x04oAha3g
xeXJ24S4mBAeNiBaQlvulboKN36C6BV/I9jWXBlQmVmbyK15YJ7upEo1lFnA/tHw
HVp15SARPC8KaYOYBmuKYQa4NY5nv+l2rHVHBfbdEFtwYKw6NYF9L+B1c6Xz3aHQ
b+VWlFRccGj0nsv1zLi9BWyNJ2srNB21JziUEiuIuB/88wKi8ybqp6yLTxR9sw6h
QPct8mA2bNczAg8j+02oDqNUuyViBLOB+nxJgYikR7rQmFP+s1vWknr2zoinwnRm
ZmgTi3pe2IUzWFCeemeLZ/mmthsMs9hb1k1VUVUNCwNegv81JUBzKkgjqUpbycTG
CN6y3vbvGZIzyYUh02BcmZJr4fBI7pxek2jgH9t0sVLWNBeuDVvlgtlpUXb8DICs
d0Sa+oNMVeXif+18ZkcP/eoRb4akfFI0UPkbZ84oJUMKWIMnhwMIaGCEIaf3CJgj
jmwPor9jnK3OCR1C9WNsWdJ7wHyIadLFekl0Vmusv7Di25HIGppwNxOGQU7OuRFb
J53TNjDe/VVM1PjjQE6d4f+KYmJCaLkkhINPyE2LFps14d04qvuKy5Td29ytQFCx
UpmrvWC4zOq84bdBN/eY3acO1IyHGh8rwlX0rEXzCD3hTgS6IbExKP25GP6BKB4G
2por/HbbURBocNkgD+QRyyOvwqwJkIfYVqcc+cjpLnUPwzhrl9uX8PJB898Iiy8h
9xPeZo4TJC0jKceO9FSINumSJ5G+KDnNKof2Q/Z+M0UibA5ZeReJxylyNJcNh4vp
zfDHfZTm3Z2VMIYDlad1UN2IHftLLz7/lSzYIx8Wc8y/OySS4AXP9WvhEk6OartB
nC88jERDnxOjXH/1wouTSDvqY10X7sTOZBetY25HADCcXIhcuSk27RGt987jasT1
zm1FGVS5QApZfB/FPzYE1b5MWNDCf+pW6ox0eItVL/QIuBkMJk7ZCLvPnU4zPoq9
Vi/OPiZR0aYDVpEe7tDyMdGbovcg8oJrTXNq4aBDO/hhTN98s90F6QHmptQQJKBj
QPJVnWc/fs4GeSsF3WGLSCdiuymmhduAsUMZun73dpUlwVLGV3yL0RTlAhDdKhTr
+XnXeCmDhf82eya2eZ1Cl1eTeK7Uvi8goyqav2/mcAQtfC7qe/TqtRdjLmjcJGp4
HZ+MqbpVPoVSBNZ58aQBq72Qg+3uc86VXqA90etQ7CiOTSx5S3jLTwH7HtRiQHrd
JvCLr9FmCTWJyqFjBugtReKg7H3gLhcO3Z3/2v3vn0QY4JIR9hSd0LQrrHi6SHDk
HFdYOVEgh2KNE0ZzmYGjCE8cSNCcgTfDy3LyZfir0z0cUSQIye6veh1eg0dH4O15
37VDxab3075js+fOZiKjmObwQRgWq5EquH2eEnecSgAdmVoxee9KuX3cO2ATmLOY
HSe8mr3AzF4SKQ4dVdoax9+RrB+PS5g6n0X8KllCPX0dKmBRZrdmGFXRGQ62ddgM
WJgwiXf/NDnA+XpTVh7RDF2YFjVQ5/aTiEJOV9l7xsvoIv+bLrJcVhHROizmp50l
AEMM8dz/elP6dMLahVrdz62Qha5z/p8qAiIi/YRkBIjTQbz7X1v9tHx7WLyD9USq
LM7ZVEdIDXigWpF3KJ5VHlakV1XeVwaRE2FIZ+RmXjBaoHyhbxDIkciIyDe0o9Yd
g9bw+GU43DMOMaMsDIOAMCZyqfTbewdwuIjsrCSWxQEQQC/OlPBkwzuHdf+7eC/6
PWYBWwHC4bPzKnBAQrtp4VkGPJ6r3NUtvv7aUMNmFb72Cgn0fv2H+h011242ZGKu
kVNsFmyls8vV3O9OwMNAVkl5WWCSLaR+RcU/97JS/c+JRuvi1U71BKpQtowPG21z
fbaLLW9gy1gwOBTf0R+hO219BwKS3U7QrNPFH452uIKQ9SaLPFXg+Y+k8or73OlN
KZy8bVI0DnT91R2PSMWQjdzLJtwybq/auhPNhtgDEgWVTzEDDVL3jTuEo4VDx5TG
LX04cFzAPYY1/2dsBoE/8WK153pmAXQy1XNiXjfGdeYgyraFhtiDdy8GAsZTTsCZ
StGk9on14vnrYQZYH+q3JNDStwYWQSzaPXQ5JChh40Qk0eLW/veOVKoCUftwu27O
+xq2p7eHm1hqIUyXSMAyadtY6HIHfXRUhDPc86N2pVB5dfBBYHd846003+Wah9Qv
gADmTy3qDsdfigZqIbnzcMsFpCJfNbjhCqZdjlhU67QsoZUq2kltPeyJ3x7c76lI
rvqbLIqwy15PQ3BEbvspQP3dqfdafwnjEe6O/J0zvbO4DT5WG2S/W+jAq3UJM7KW
17Qq3sGQEOV9vfKMUxLmC5hK/52WVkm+eZ3ua8SS5XwnegflF7myA4uux5yC87se
6kp7FGFytsSLWcCOL+chD0QlM/T0gt2Vrmy75LA/imZL7RcIaXz/rF7dQdVsyjtG
pYNrS5KUDdTamfUKjbkNDmf3f9VkkBaoiw7jJmxJR6FomK9xYQ8X1jeJgRCcEhFi
Vi18n32sNHj9iWsS2LoKbZlgFrRAPDkoZAiWMrNxRmzeSUzdsNxzymfHggFwIszo
HzZoQRir1Q4VqGSCg+Qd26c8+ljOY2V3DCg2js8tYDRWVwKNBayTgI6qHPK1SqM4
XNBNfGzkoGQCUemvel+lzK/UP8orD4OrJjbNAEZj4vTAJOulxyiblfC4KRVjlEmT
t1yh3wxW5OdDdM3XOdHY+eWCDtA1ypgY7/EA6N6ye1FJDvXeinJ1r64l9SRB0mQ7
9L7Z94kW/fI2rzAK073JG0ABv5UXp2lvH3aFL/JbRYRl9BlunItCaTYRUsR5RHXp
GbEOf3NvvY8k7wiyzE3EtIAECRpr8mUJtSUoJvPo6Nqs/3XdM1kSHfxxtIZs0k3n
RnBmst2reYK3m3I3fK9TtmL1TAKMuF58jP7igROTB0/Oiw3QYYLe66wX5ulLhOR9
t4KK+R0xVa9cddg99wJfZIfv5j8B4KLx8dv2LTxvNIuMiTmLRIP5yGlJmofTc/I/
x8uLX8bwf1x0qpULAbGQajYjlQGC6EcwhBb7qsz6QYE0m81U9YjcOZVW381+MSds
l03/rYdudFWCUpbX/Du7IKp2Q/Cxd5ki4/XwQb3usgiHDeE8e1uiP/S5b7rRdxxg
niFEh9VmOyHZj2ifQpqv7ZFFmEbobCecP7YLQ5muvYOyGYBv1uu29KiDF2XbIJyT
U3ezkowZYf9L3fMFLpJ2VxFW2EHXjaJInZsVPC4qNahodrtxKU9VHC34BLNwg3xB
AJHiDgUgLzDsiEPWYvEtKYrYYJNueFBoOwDfqITZlYthDmHoDzGKJ3qYnqA4wwM/
UUcua1spl0wsgytixWnZYmluXQR1nIysFq2G/oe4fb5ZqHpu3yRF72WuElzzqNkU
ofXW7BW90jJajUfOCkswCTh8nudGr0adCObZll+a1blFe9w0jPNgk9zZiraOL/N4
8tl6njmSeuc7V+K5a5qXKMgkdQCf4lWxE0BslXMtTa64f/UFjYR2/NR90rTs9b10
SzKJT7PUb4WQTetCJmxc3X1aPfYN2dyG0NdA8SMnsY7Khav6PT5uqjDLdU/mLjlS
tYCLEjCEoKkZVOGhKdjT+A2DPHTgMgnhMWXVv/3xsSsNFyT4xXiU6FOJsU2uHxmC
d4613PAOhAyRKiOfoL7hQN4bbm7ALSFNeoGdsJpe5NdZPdmLyDU46IlM5GpuyT4G
KDl/TLRF0TQUm1SVKZUCs5N2q5s9UtLm/JhOQHb16ZqEzAtRaCpNzpVmLg0dMcD/
Olf1jOuq3p2zFEW/N2hqLa5sSbnAA5xSFHf6nkJ8qGIkgPAOz29JELi8sGjWvtxo
OJSfwGPemJlhZq3HbuSwoDjUeV4sSdNAfypt/u35ildzHYAcEN4armWhpmvGyVVN
YdHlJjkL4rM7HEhyJjuEz9E3v5cVrVGy8m87oXEbWH623cNMtOnsEeeaEnwBT/pB
WZjhFX7SenxlpIVWhemsbhDAqouMrQqk6hJx7trG0nBWalKXSoXcPe7sR5L5DF/t
P+LqE+YPc4a1ecxsrXd0F4NQrPSGxrB4cm60ywHm37MrBAVwMAaZp5NNbijpAzcY
quFefUbE00ltGyui4tuAe02dAuj46/TdW43EsGLpbQPSOSus5I98mNRZ8zAKp70R
JoCFc5PeZ4sIUF8OoYt7RYiZG58qRjeCFAyPPyw5mMJvR4Ma8LH8sEInwqhUkqo1
Nsn1KbAUFU0N0aei8l7MXjpX+7H1JBd4gIs4HcQb1/0QEakCvOmgpd/y+DyjAUJB
l8WtvpKWzDI2U8xzPwFvxIU3gN/8m+6ir5g/UddzBFEshREtgfnKcAovtUf8UMk+
W4Qhah0U9T08MFKeq25N04rkHgMaQ/jkEksxmjN7+XzYydBqP2ubfnfIJitSavYv
yFhL4F6uyxu7JG3UMU/4cQBOAWwXoDwyQ+SOeed6zysLQo1g2suER2tOIsXgChR2
IjXUbjcWR3eQFGbwmuyE5vVYHcKwpf1QiooRxi7vI7aF9dVhiPMx7H0D152t8L8l
B+zGA1BIODPIPEddQcWaoni7TDx+H+1bV1FaXQ5b5pN5SR0nYHp0vpAOZVXhvg8P
3Fy/HmgQBtTUCxhHgBCUIm4zO1LIvczsorGOm4QOZBgNt1Nf0EZnRhqfzDXFS5fn
beJihG2hUXkj4Uh+gxIHMm703JGc/lIVtEEkBs8t1Kx1jekd6xkLLhiX9K4q+jfP
qYHrL4P3hOZJaC7Pj9WfKenL8Q9KMB/KnpdZvHvf4/O+tGqBvuiQGNDjK25ubSez
cmVawZnHARNiK6RqpbQcV2FU4ryp44ms4CZSigg9kXpqoj1kphSm58vT9kKRjXtu
/oCq7uqG+rVHrAyKC4zCZFC2SbsZwRzNHJLDqu77pHPX2CdX8IaQy9Lu0h80EUVS
yie/5eio3rCqIB414JmiBwN0mr1YNM+B8GXtl5DIGty1uVVwcFuY/LwPWDz/h8S1
Km8iLZYEI8wxqHevJ4VbYMOy+Cz0ryR2MbHvWQ3aaOLfzXMdzt/TzCLMRCoOBlCD
wsyaU6kACGTnMO9W4QI6PAJPNxCVQ0Q+VvaBil2ixdH5EWYQdsogEYDeJraReeOO
MmUbK9Pd5j7X7FIxdr/fZ0hAS5J/xRtRsKBJAbbGQ/SiO8z9hQe2CsOJhvuXhEUY
oC9OCe1BBOZ4BpV4wjBug4B92EzYwVNQxegvhQVevjz4cnsXWO3EzWWj21m6SIcY
0NeFKxxYB4+BUHNuyDAdXV2AgOrvZcyH2/4/Z8tSOSg2M3YO+1aD5kPffI1VTfW0
MX0V44Dtw/VjmHeXL4LG1JuUGs+OIYmI/ru1442mA0ur+5RIBU2XeMRHawgS5kOu
HHjJ+dZaWUMA6kZoPswz01FnMj4Vz9Yx1UaGTVfvvk2hFukzSqX+onbngaObno+5
+zXwBCPgLBCMo7MIf4qGHBIYwiuxlQ5tf/oKFXIZ4IcEX2xJvCVzfvO0AfWEndRv
Er3zgnhtnX+HKNjJ++uY24pdUSBzyC4NlfZr4DQYlCsTfutOlD1kPmfXdgyuQ5Hp
QaqjmJGxibfrg221ItE/ZW5HgKwhYpD5VqAe9PaPGSEtsygJPo5dNw+vzppljcy6
GLMZJzOZBLdlxAI0qBU0dJ1tFrARZDLC6ZxPlh6aoj6butTXa9LmMW1h35+1pPM+
52T5ve0I5vyTgbcwMrqitKnwIGtnYkCxdrliPjG4Oe5NpOKgQS4w0zSKUBdVXslB
5EOEO42AZqTGSrEVmcawlXDFI1O2VHdtoAcyjt8aW//cuCu1UKIJ86Sq+B8d9app
TMUl8wSNBZn27DmyOOWGaBpffGwGfQy3vXv47gps55lXVtiw5+QqKNLGrECLX68S
fEH1Q/h50MHHl42OjIEbIqmGNJXCbNfWLP1sXUyhKQGq/wE5fplq/fmYdZQsG7Nh
P5oNuSm+MZi0X7+mq3jHsxbQlK7yY3qnTRw5S2m3nSHXRmV/xGcnEv+CQcJKR9LV
kj8WhJGrn++3Pjc08/rNiZcM5w6CoxQEPalDwKV5jLj8GvksNCKpwpXEhITsQAtB
qxChr3JYva0443p8VafRbwhys71GaioLqgv/Uq8W6Pm+GzUzXUte+5+cJNhY6FvB
GitmBcuQ5EWMiUVVkmGmD/dk4Rrqsviy2wUo3nPdrM1m3wX4vclC/iFKmB3/575w
2TQMH7yYloXnACKUWIJu8xGfNtPbLfjYCAJRE94eC4LYJ5+LA4qSrciRaB+cX6jt
RhxpkoUFZAh8zh/91VXCJh1c7Z2laLihNMdD3Ag5RG3g0GCfrN9vNVf5hzfMFsU+
9OEagLcvGW7Y/nFijwBYv6pqTi07rXjm4QOGxrIdBPRQuFXgA/14tTUv4Zk/z6So
5bD6qp94ev95muX03meXc85bvMaNRJSdtur7duMi2uMX7X1IgjHgJ+u6DAqCkaFu
C0KYFzMth7upTlfZsjV69VWOrpqIEt72GMVYJjHmovV/mTImXgtWh7aJ2bxyOyog
NxFMwgUdlRwLgWO3igXcdc3rCizjMsPEq65uuaFczlAn95PdJWWGT7m7a5RAy9MI
Go5WnjOMV5q+7k8lsbAWGmVMJZEdIZOkgIqlK0u4PqIMSR/OMwXQIJ+YebQVNN60
ayeXE7pJTMfUGyC392ZJ008Ue/XKP/SMkyR6k+u3XYQt+szc3EYFqmZDHXoBtSyA
4aJBbTpE5FqV9h8j4yiypSwvctf+76a7JNl/rBp4S8hQY2tuOpNg6Ywz1YFdhwXU
wRm5huPBgV05qs5FMB84eMId/4HyLN3YtX9aXpv3EZzVeMoCwr01HDRMH4y8XeN5
TARrwFsVV5xN4HroNprb8KjWcWGfGcpaPItjTMnVGKHNOSKmJIorsbrcfabE9ppw
ZNbm3jg1d1An7ZmFMy78w5vrjVXulANAPXqosRM4qpOfdAbL/fZV98CmKQwK1WRC
2RP/Dlos+I2Vw4pECghCLUQrrqnxYi88aeHTT01kDDuPRVed6E5moSPb3TEt2h/q
+JnLYGSs6fjV4GRoa/s+Cnldrr5FJuWZQBUrNmCTWred4X8R9D/b8RzwsUI0D/eb
wc/beowWf2YQuQMnW7MBHqFYaYuCOa14P4NhmfTSW33+8jtZHYn0zjgINxnJ6xRh
LNbtbM+uupfrLcPjQeWqZzjL4/Ga4izAvb/R+YPzQ4b1fh7401IkI2hmkSXXw0zf
c4VO14ThTDA0B0I8LNSMS+BkVfA57o2KYRWt+GA8g0niIcMBFpPUFa2A+Vx4GvUZ
FxC7tCrNnMcqY4r23OKNJ5MQK7dtVNlOWGJDkXhEuIQ5jcq6Z9aAAARqR/qA13W2
mM8PhmtWr4sLP9SGP6kA6si8pPMjlyurxypu4zuCxRIjbIOW021XPxX35XAKP8nm
2L10+zS+EdyBG2FX4QkdXkkaLNbNBaNO01KiU4EKu3jsrzFO1eLZ6U9azAgZA++P
AAOMMXNdae+S+Uia2XNexuwl7yrczxy08z81nmmQlDmZjjww/scHCiAMUVloTtjW
eVybRpi7/8LgvCsSpJqGtFWCxAGwXsoNGxCRQH8MitvmDkYu/CBUl1kCrrjE6oFi
L7J3ieCYVVTMcprxm3OfM0+bX7M5zjn0mkDePM+qvuBdJlol7a81+cfXYAib1LQy
SMMu/FSxUzywv06N5nL/Fdble0L3wz5+jMgtoH9cLGUMO7NEde/h8Xfn4ZZYBIUt
Zoc9lei/I3bd/7ZlTJU8EqZlw6P50tIlqlK3lbbgObFvCcNMAFHFv6vT6ZBInFWu
oboHyzXPv3T1d07t8kdPHRb2e7hBLOc9gCbat0wodBjgufJG77l7WegrLgxkWCE6
DdjdGZU6LQ1XIOIfnatAkfFovonRiSpQRpXLoyES1aaiwwCzduTP/EavoYqMXkRv
MFQMNmdZMwuA9l9KnPz2MCCwB6E2lvuzHw5n7d0OcBhBhhijrsKgU7+Y0bh47RbW
EiT26r+O2Irykr0nftbVW9UOybLi0CMceGkWFWSPkn8qtAJQ1QhLON1MiQetC859
/vvD70X5E3mrVY/ijhjYvxiWqlhLJgKnY6EXQPLtMzy6yVM8WKSxZd5GAkzdlVKz
oVMOukZbHdiLUWGrcBO10DGIJ6PQXwcaCbWGVoRBSP8DaU4t7gjIudofTKi3S4wa
bDDhPh1eHVqrQTLRPLOboL9djy6a3J8HuVy7XhfPbLwWkvxkCioLjudIrm7lQQxO
Q9w+7pYVQc7LAaHLfK+9jkto5BEUIVNWm8M+KwzUA9A2+LEXNiQgWCjG02fbSBBo
mL2NnHMZlic+t1LnEpng7lIr0sDgMR7nU6XQJNsVqhTzhxA8uU5wtNmuc96LtDAK
5yGI+BjU2JVWwDlKUbd+y1dRTOtzynEuMjUaiUjNs6k6cG+mZdG/FGd7Ieu2c1Id
E/teAlML5GTcMiUUez5ABNVCGCpFjSK5kvmxvhqad9nLsomlN2RLRxZRsmYGuCaJ
o+P5KRe3URYfn42Qf+s7CmpuFgLwP0+U+U7XwzguowtO7DQFWS2jDC/W4YFlxqrr
35oD/6rT4kSa7jAllL284Z7dTPijMql8ZINpJBBqusXT0Mx5R0Z5ECAff6SHteFs
4S51zgKb69/wIg1T+Wjh+8eGf3yjvNFaPi8RPBBn83D24sTFaqcbBaBy7YvwTL5Y
6q52KiWW21kdUrKKNSd6hV54rNjotzc8kjRaYCH6hn13MTxiq3FzG0gUWA593UXc
kwyg3bdJCXMkcNbZE+Xcy55WE5bAXSETMxRUZLbA1ByD5N7U5gp0Q6qRq0ktBVHu
ozwwJzfLAM0xMKjEiPZ5gZtZjZd3U+Q4SOTwLUTVbwXCv9sUSahAG60aKoVLyMpT
ee1l8j/L/X+v16f++izJE6gDxLefEEDiBYoZftwVSVXjP8hhCgDCpgETJJD6zTPQ
n4Diw/ZG0ST81+3ABxqk/EiqDolvWUldNa82m6EC5nnC9JspHrnN7d+xS6z7WPD3
I8DeLPxDE+U5tSc2FTx7xyXxVDnXKfln7HopAJbDnF1Azw5d8Jdau1vEo/E2hwaW
4r2bfS5mFw1ts3DXn5SVi7Z4ldNUxWebLEWC3k77VW7onm+u92VMAFXrStGnLsXa
5/urJ10NGdTC5TZ0dsLgY9ABdBZqiZdrtktqMm43xvySQt62M5hrw+Mj70yHrQEW
bKe6/Dd7IItYJpX0LkpXOwaGYERYw3vNXaG+FM+UbXpGhwDZoOVUTswRqWYONBd3
xVdq9ypOynmGgxT5gl840Jnh9bHNCqxA6bstKpH62/pfXASncHsC0o12xjWuCq0c
LTRZS5vMnBurLx8EENZ51SDjGbK+cUavU6xz6jsqch2IhzhK8kaxg5KU9P2rdCPQ
ClGg9MP8ibR/LtYae9A6D8wIivYv8EZ70n5c9ZMbNmKYvTYYwVGG1seCqrrqJbwS
L2DaVy98LhcuuGscMsI2TKjWBRbGM9IvaOQR1qNYy7CxiAOFhlscOHEW1w7BRXoi
LmNUwZc6jgBwEQCcHHu5D5xSjJTC/6neX1MQf8x2g9eQvNAiSNy+p2zLuO9QNFAo
ZNAaCCXpkZnQJnd6w5sQzONFCceWyNNJJpIiP+4ddwdzIwkTZUTZt5AOhNzR/lM6
xoPiKmFHJmMFlhsPQF0q+GJ9NoqirYlBIPeapfPYOV2G4hlacKeHpG/IcCvXNRB3
csxRGqnUfA8J7g2sLUzb8HCsw0qUDgvTHtLgHBG3yK0IlF+YSpr+KTYYS+x94WoL
1xpBEclV+QEV3NsXKTllWr40psgkcj3pLVDKLlRoZmdsc06iRpZMIV6hP8lF0BTu
OIujCvu53eg9BiqqT9Rt39NOQ7sleJKJGglyNWQ4fBQDnMQioirPKxlngpEvoVXF
3XVbaJpAYQAMmDTqLsxyzIOYJwQOC/rbqhttGozFlvvBjbmCiZlY5G4xcK1Wut0X
HXn4R0rMDIguFyGKJIFduTYLBDSvM6EakbnlHfLG3hQ126grqZixY/pFBiHUUORC
HPIKSGRQqWauMUR+VMZ8yuCW3iBrPG7QQOPVOq6QoMI8INEZ+kau81ZKP11wC9bM
KZJ73jCs+2ozSor8TFk1qyH9djy4jzCQ2POE3/FstQl7XyZij/ytH3U2wq8Ra3eo
S6c/52B2BYyeDAsTdhuTDqSMMx2witRjvoo6U1L+T7Zy0ev5uFRJMTD4DcyuoSkp
mkUog9pBePUkmS4AoFSUY1Pi+V+/dFWqCsFqQakh7aLY+dLWwSbhuTMzkqlq8ZKw
Oqp1qmdMHaAMgNFXgX7QQJFJspUAUxUHnlwgC60zTfkBi7dfV9bB6zL8xhM0Qk16
LOfqgF3yilqbxrA9Ntq7ZMUA/nyz/9EuZzQ6Pety9jLSHFj2bECJfiOGxZOpdu9I
w8jRm/D0nvi5mJDuI5fqof9PaMVWSTEp27bYpAnHm7BlwtigUKJCE8WRxtiBQd21
R9XqABRjLw23DeZFVO8m6QfkpvgwtDAJPv2p1+6XRHII6dvJ+ItjuSRXeay8Xv/3
VTqI4RmZwEEtD06RssJioGlHJaZHJ2SzwcLnK0oYDxzlTZAyLswLIvSENXohtTYg
cm1ChiLayGz4lTqpW78v1YY/fCDmph0Hwdw6MEry98MsvrsYLTlFZTJKq16bDO6K
7J84fFAHaruMfwMa+C9ExPxQVlUq4UaQ+u9Nqq3im0NE8gvl87SAweL6n8KhvH6w
N3B6pbkYWJL5+I6P9QxMSM/JVxnVMNfcABBEPzLzfrfSWffrBqJb56PaPnmxwnsQ
azCEB9J55dFyJc50o8zuzJQz7kX6H33eqY7pNWrg5vYiMwinjqAe0vGC/uJEpHs3
OzkvCBMFG3hdd6LVEJeE5CjWAJv8+cFX5verzJRIz3Zzzt7VqBUv8WakjtFHs/OF
L0+i1LhN6u9MijwkJXWGgdwVKB5HL7lzNLHlbNp5IL29/VQl1qz+V2L/k3dvgoNG
F19+4CLVSTKj0KxUdPIpQuLrT2lwRYBOsnf8pXRQ4ATN/onaNk0Of5i8dnLByzNz
pAB/H9b52vOJ6cOtMFe3U3vkrVKwZlaaTGFliHAOlrLINOWUT85s731m7s9y39Px
hOb9ED2A+rAuPMlEFjDcwVoKE0xmeJnEiYDb36JWG9+z2M7cVMC27QnpMfqtgYaH
7OAQFTIT8DptoOWHlAtShegDsDJC2jf8pj3r/rGsZoSeywcuyW4oIajTzfum3AqG
1uihrzkfLYxIofSHLGR1DmEYsw2zIDN1XHISukM23zl9B3jaeAyhDAnO5oQ8Fb0A
mTemTdl9DttwcsdCLMS2bIV0usSiDur+4ljG6Yqk0dGJJl455LiaZs3VP4dF3T3m
SLVt3T51txnPmzvOGzLw+wnqPFnp5DulAiUZQIAE8HivcNyQmJJaEohlBxLj1Ivr
kJT5iKsdUHRpKlGG102bHNBFpB7yKwJcK7ZoRLj59kfzgFaVQMdx9jcg1sUcjLTI
oiIIp9Ijpng9yxXDFSeMeJRQHxe6g/QKVkY7NCe1Djfmb19aKczWymfUDYrWLmHa
puK+BE2YRxF4DYV+z4pkp57Q7Dn7YKX3AXzzYKs5w/fb7m7IMyoduPENBcEwPL5i
gh4pVRtPFR605RknWyoVqJWXQXHU9zysBGjTUPBEVTiu/pWkOR1g03q7LOYVaMSM
jg/RSYXGVanBDLCtdkKp/kuHLOW9nGYu/UmvgLrI2vV2Hj6hRJIzNurpijSu5eDu
WJah2xXKELBj59lnsSLaDVqucwc0NgmAMHBObHo8qYHSC079M4zmV4YfXsPoc/MC
T4zz7aiL0LECT+/5dT0MGK2JmYGebrut7GLHnBBjZDA1AgUJ6+cJr6kRDV/Y0ZHY
Xko+fogAJPUfdMpCr44SHrZ+NVr+aB4hWAAxBwscrUhe23/ot4UA8P3d7kFA3SJS
10IaGD0SOu6qh3hC2RCpNmK85HpD1MUrcnjKRUC0vikm8gNoCkHFSZyoz4AyYtGq
vcXhCipqrouLTYDVQ2v5Ir/pqy3NJwGycN/3fzUoNEt3fnh/W4UnlEDUPwmVQDkk
26id1po+jXlyzJupcUveCjlluocMppCHN1fokj/df5sKX492TsiNH3NOcLe5d6Bo
zAg0oW3VzP58TqCTcTnhi/AsjpCR4ZQ7pvNFvtUMq47/7mLNoXt8B3TlfMUFwCWi
L3FE77wg9ZmlgCq4EYi9UbGIA0N5OFIYq3sIqt8usPLvSMMm00GEVS0Inr+nNh94
zc+SXoiy0xcwe+kBROhPswW9060Nwic4YZGXXIoPOQ7CfOs5PWjo0z7IPweywCH3
yGQEyeQ87KtGR/D+qAFnbPQuU3OQQDOQ8wOvVtLAL9PkBPrxzA5k3gFbk1TsIfoq
uQbqcaYKV7DUPfXHtWYvUSqZgdtHmHFvmxR1Dg8B3brSGYHSbygbShokqj3Vl9nd
4Tv6vLn8yG8D6GswkFvxdOpxo4xikj6NNI93tnE4XghapGZjqbCuaoLWWXkHLj4n
ddb94sa393sQjcJqgjwbfUFTgxMDcd6Iih+n0rZwNkqcO5hrogCCcesVtPJvO7nX
/KXYJLC/o4iluhngODknzTfedjDCCAIEM9o9om8NED5PEkrrl9dlsLqv1qA2x1YX
RD9V/sn/Nodz/o8I6yoXRnJR/qd71yFau+/MubdC03KR5Gdz6s3+zda5l52acf/j
pejoQRucGY5NqSRqFH8KQSTqUa/5/UzHawWkipeL6O+5lvNmyb1oOyfpdGNx0UUK
DzasHTyCfkOYEY/D0kf0LdmCvygKYM+RaBT1XCXBm6xmV+eu6WbTwsDOEvOwL2Pz
NrdzCfc2Ct881Wy8M0m9zoVnUw1xYSjOkM4DdXcJVIhVDRxDd8J/nScnlVc55u04
4+6PDALOpkFCrE+4aRUr5ic/P7U+oLUHvuma3WC4Zz1B6oz6dYMmyoSN9/EBEm/S
r7ylGxNtIcSkNEoSA2TTvHIR8FFlJDH+Z0HXoy5r1TJ+NKIFpdUsq/qVGw5Xv3xX
IHp9Sdw2WLQsGdaSAB/ujJu/8Xq093t8N0ZeV7bx76jbyUXK7Z0JRDQ5jjuqXKVN
PNPyagODs1JASG7M1aZD0RB16rMu1f1a6tbl+5uQOd4+ep4T41te8X75rdKxw1bO
afsms3HJaMs7KlJNTcT8Bpz1FI+W2KA7Bij4fhm7SHm0vjqNh6uV3Re1qlDDXzbT
Sk1F+wNutPqP5Du44/7g2qh+Y5wSy+mVczWHhHlbxirXQ/qQLrOehKO1XOmWZ9xk
BonSX1VxcJ6eaQC0UyEhDvOY1QYuny6mK0dGxRN3Q4mu9U7o6CV/VpzlXh4Hv9/0
7rZ/M8/xK/1tCmXnI+9NlC1snKXhUARhYq1R4jmAagPxTEavh6NoTiIlYdlgZKuw
CMA95I9eVxnbT08GKFZZjLDZHDIjuRNIMtG0gtz+pLeHCtKEdh0xYEb3AWwhwD7d
kOh6VDRPYFwa4XVksxC7yhxznexsarzeNMLE32Ps+siF7aeaX3nTlt4CZvFoForN
3fxxN7MG0zipJ0EKegqdi4mO1FYX1YsZgmWuOtOffVD2Ow89c7fnfXbZ0U14l5Va
LcaoBuypqohOFgAAtfKW5E6s0zInD9DNykfV/FpoybPtaMWLwLqDH/E5pQuvbR33
6SQ3Eoj/If45vkVfUKkh35XA1LpTtgMRLM4sBhKtS4zn3mm/AQ5Yxux/M+vu5L+i
+akFaF0drHMkQYO8PLv7nXvp437fRTTPAkOjMo/qgZ9xvaQZzsgL1UQwk1AgIwcq
6CUDNBWzn1K1RlQK1mMR3Fs0wE70OQAI7oEK/58SwMSekQajNKkFFVr632+3iu33
QW/1mG36Hf+4MVmG4c1/ZhafoYsn+YzLi9szOk+Y/v8ZBm0fbGIYX+HNxr7k/UPF
EZ/JjbsyljmUNzjW72cH5fjuFk+lY+V3ce9eq+/LdJEIRTrBt2sFBIR4ckV2Ezy3
Q40xH7oUKWd0T2Ho87J6ac1+ZUF3UQBXa13yt8rsjzwHAgw93NQX5+PXZX5T/YtY
fg97+T8Q8n+qvDVUCcj/YvaGxZGkUdqPxv67C5v1b473CvWRPIBRSVQjl2hcj1Kv
DElC4+qnQANMkda++6TmN3JAe7QGpaqKQgWkj4bnUKdwsngOEkYo7iIhCa9x08uj
rYbs59658Y8bpTX+58zHwpfsrhE3U0acQXDFeMaeXObwzXyToHCZc9JYmRKYgFpX
pGAhMbczqxmqonXss7uD3vBgGbYXlR/tb1jMUi5IlWYqjdsYUvTduwHIs62BGXLc
UQ4yVaQgK15cAtww8Lj7CBDH6gjtIapOCYO35PeU+SVQydtPsVVGPKq7hAaQU33I
5KWRaMb328axOE0B6wdRyIJTPj0R+26KND3G0sZgDZWEQevi+1buzV7R2ajWdhFP
s+Bb8DNaulbXN1Go/+dJ3bTroM8KWMLLjLDyRwcvOZYEH0fDX9myW/FEoG715GDv
nhObJvG4Pvw0AZ0Ow24DX275gghajGBbNEkLzNl+n3iGGmsE3Hs9wLD9YMOt0JeC
RS2M3ff8iCKNTvxq6q/QB4j0HjmAXVS9//UXewDu10TM6IXFwg7JEokX2Ok4Kego
6wHFQ0uwLGdTNfhLnJRu7y3jGKXHrsc+VLNIDblgAsFTZcdkE/R7dY/uWsh51VWo
tXULNDqJac1VWRiSKYetx4lw3EOs67qqmR/OrK94MLJhP8t0Ue9l4H0lR8hKEuc0
+0mWXZVN5aLznqADdVZYih8owmElG8GH9qku1iz7eWrEhyOYVNW5Kw0icGz1JIdM
X2oCBB1nXn7anncgYUm4aRbNJja+qIE7/JX0Jidz3INrea8PZdb6GsRHyCknRQYn
ISwwOk30lQkAEcNW6aA0UTe9i4tUfBiQJCXA/H2Ce+rXmep+hrlnv/whnilkInmy
bDAdrZhevgtmW/6ipaiu1Rdq3s/63Casz+19AcgJYcZRkzwLppKdc47FVyX4+uYb
PA7fs99fXvRwu3uqvbF3N4gQXUHdlBNI4Jd/J1o0ceHOi7lotCzHnjSWEP8khQ6O
UzTMCXT2/Q+7uhP/xswuUI5teVEoTyr3wb54MR11aojiKD4xXd5N1wz3DQI8ntyU
/HmwmDtuWS0UYXHodg391QmGONPGA8ibqoWpl+YWFLqUhzhq+3ds2bPx/XOclrhH
cJJll0QUiyP6xs+Rbo4UGjLpkW8tBY87QYfNeRBl4KzziplDuQjeLxZiig0VgGsN
HpgdbpdEKs+fex90A8ljjvw43u5xFIUrCbg/IPqhbyqI0qMc2qJ77+Dl3p5hyK/K
gTDfZ3kiygq4Gc/aCm7K9LE4aI21iwN1KGAK0o+/RbOX3pn/EEwjWuQ/7MNO2YMP
piVEzGnfCpNsLjspMfSMtPadX82q0D0YZzUquTWYq8j3if0nHnmbsXKLXmemD6lg
YLugPJE7RIa50gPgmfgXTfrebp82BKZdDvN7aJ2nCxNyIQQwPJ3yfe9TyvbQK/Xz
XiSpORBN+6eWaKhD6c1oX0JJIhXjfCd8za2BG7yGDq/2IzrKjmqbPFSsmDfJbhnk
G71AUQxBwsGFradtQ7+ySyKQV2ddGZ4D4T6cmj8Emt9FVRWG/wvUqGH0QrrNotzX
5jg2RC31+fD8TkLVdXnO5dJnow3e+1Y8OBZN0wOxS5RcgzHnfLprE7vTZthlM+EM
behfHSDgM3XCvibmvYDW3sX1+FYuPBOKgim2UN+PqhaYtaE3k5ziHRZDYqQ2nm/G
tUJbd20kl3i1wCNMwndHHzlMUzEpZTeM1QnNVxkWm3wQU1BQMu8EuCNun6VXU2g7
UDNq/wMIpqO77tFnq+GY/uoXoypEGHE2rVVhzkLoSilhZiyt7Rs6AMJ3t3rQYp8t
BRyZi7ufInSUxaRtjGP6LDk7OpYOVWY1hJCZnN4ZjLWUTFORzFroeq+ftIYgcFjN
ogyUsg0M3Wylydo+lQNDDcXf1W4fMBFdz6q+SXF7M6YHrtpfb183uNv1kODnLqP6
Awsj3hK9QnRZPSkc8uODPoKYehKYh7bbZqxqSgLuF+EXsDOznrd2nO+vWZAWdLmc
+EE/8Bpbrc2R8itM8apqEGOwCfjl/AWLWqs5+ybmA0Vydm7TxfJfc7GHPZAG8/LZ
GsTCpx8mmCOMsg3FKZ3zJ7eHpJnlGPogF+/SK07IpoaMaBvAyM1c6EagKhJwYfYb
JHiIM6H4kiW93GTHZ7diB6BO7L6yJ6Aujt9eEwFaRm9Hgd6eWaZxSUw6EqXfpfm7
8VmU3PYnbEJIlQ24Fy1W91xsg2RFCy18+4Utca0plrQFtJcRKYDGNivaqqhD9tad
D25NNPu7Dix7990hmP1wQ0BcrvOBFKR1EPNH0oECMvD6d5C3uDeCY7rVKPj00xbi
2Ljx3ouIiaG+CXEz7lbXMp/6NpdKb3GY/vYMMvI/YtkqxbKVCAtvA38PoIeTrwDX
jOSs9HOTiw+q9f0dvL/pa0x1Tz0jivGHP8VJwroME+hzjSpPmUWcvP1J6EwX2Adw
fldfzBkHr0Zq1M/2u+1/wMCJUrS7vDdmREs2SWmcDhH/0/loEIudGOpyzEDHBbbH
A27TkDPk7xmmXVPyqHfoT2KRysVcKMBcOJU3O1GOIdXXEN5+pNaEri8vfFWc1WfU
46h68SpNdNv9YgAgf0k6D7XpoajANULb7eHBP/KDTCyWykHxSVzM8DHPlfIinbFw
wXMY1sFAV0owHbY7ewNaWFUP4fKeYMlex9RLxVcqntXBfyhp+BFZmKeNG8AwN5Ff
L5IlvmvE/ixl8lYmjXw4QnzkFwTCI2kigjf4fj9vj9W0gr4tZOz42aylB80l5gEi
xLa27EUe7yVkZOolA9VTHHimYNjjceISOo84dI3xIeli/2otPVU8HlHA9MTh74f/
m9ZFERCNt4NTBrjxqJaP1gqRU/UBQTVuf+ll+sy9zKDa5ZgsRSKbCrHYhpU3GyvC
d3xgGvf4D5M0CAhiNeOLmVvwGJaY3GkrYhAXLdQgAHOlBYN/ZssCLmFY8IT6wzmJ
oFtFQeWaFl0qBy34HicXUDP5HNZ7AweiSY10CLEKTQWY1Rvzm/z6WrX+uEwl8pqb
a6d40qM+shrr2IhR0fIwaH/IGFVqRh5b6VqZ5tCKHgHwfuvVQehYQCm6IpJMFbnK
F/cysPdphk+lloOECCUd9o9R4v7xmhI4YecHXI/L+HkbKN4GPwMTNel3lgCzap2Z
4siZzXG68EbEm1m00LmY3Lr2HOdQvNfN1zaweCxtymarAWCGVKodgeiOPo/GQ71d
09Aeb6MUe7ztV9EIbZUybZl6TA2Ly7XY4DGYjjwuWXvNxBVcTAPLnuTmovOyaFbf
/OJo97WQs+kaRSBZ/o6v7YBwpLya1wLhYSN6leAnmNSrIN2UbHUqwAbanrordYPn
m2udJVOWls0dZpfXeUM2eEFLJh9b0F/E1svp0eTbs5/jmXNUHGhLCbPb66R6CUzO
qSOSqmK5dY6sstgZ1M1+rDPbA/YgR0IwY54bYQMejJwLa82eg0bhVoCKv6C9RWD/
32gulburRy2TCqMppzdHbIERFlRDaPLVvfgv2EWQqjXqATzOq2jxde2A8FDkLui5
RQU0wuFIjJceOaXN3fynVt+F9YwYfM4XYC7Q2hLOuReRbv3uJR5CFjyWOj0Fa9SU
D8pvsEmlyYe8A1cN9j5qKinyP382oAoNJCVSFim2A8TKllRGC+zvirKo3I91wS0y
230DZhAB12nZV8WbOh0/DI+gWv4vrgoRhBBKjp2rPNrUz16CVNDQxggXoiJFvPXd
uFHKIgf0oLsQ/3+HA5u46I57kRtnX6REOFUKQnyGDn638uawCAVTncb21kqnThpj
0Dp2uke/5YIm8g8rX2nAZgoSgNi0V8kD3j9c8OdLREMphskR9fWhYP61IJ7sZvOP
msIA+wur0tkSQ1yR6qknchunNCbWzbU/99O8T2Kp4BzdRCdpvT+AZXTZHl6FqaU3
fdneNp8LcnTZ0tjHSG4Dso9nFthGeUxOig7WZscOh7EPUo9YxSHa8EyDk0F0ln4/
u/8xlmhHlm+8hMDdqNHJRoD6CQfLi0qDcFwFdcSHXJo4FukYscRZjAGLLwohHDn+
tD4TKQVSm4Q14ONCAgFPlsYt/TzEokbYp2AZmS+vXvwC0bQV7LWdNne6DS2F3JXF
t/Sy8Qk7Vicv/OtTDkR1B2v9KAN7iP1IBXdALd5mpfBp+b9G5AZbw1xu8GijEgKY
ie5dFO5Tqax1re3CNLjzkSRirIndF1aJ27po+wPV9Qq1BmzXb43uLICbf2Avs9QB
jtunbCCfxkWpHLljMWeZrt0iHtHClnX6+k2oNSQ0jTEoRgYPER+yCMuXD5VfTAMp
tyAX2846OCU+2jm3RoVHpnnLJL7BXkvFdcL4F0osIqCjwg9Y+Lthu9T1AZiK3C7w
7rw1z0xC71Dr5PwCojblxaemiVSyS5cZsjQbz+M6hD74eP5KpbWMAIwOFfzn9mx4
ooz4H06VUy9Yszpm/KVn7gbVCU3frNFp2N3/JF9Sq6sNiPmw2EA9NGuiqpllefqL
y1Vf1Hignr47klG4MnRN2uXmAmveyvG6/D2p59HsjkDZb5fLLXyjK9iIHwbrgVk/
vSqymiYf5J2MMicclW2tBlpzDBzRqCVZIOmwvHqiK7t37lNpDy9ZlG8GfOa4sfmi
cQ3DeMQFCkqLj1gfsk0ancSlAfqwyCzUMppQUyZXZuqS553Y4BdKmntuXtFjcvcS
1k455RW9MWw1cQcurH0p65pYmE7pLSpQx+nT9Hyq2YUnEPBPHgsLIZItsrQDnMfW
8xJzx8Njg6A1tOM8dx20I2GBuicaYC4msM1glnK0mZidDxaN9cbEgOBZgpBioVDD
7ysWDjAl2/zgaQJJve57fGap7ixK+u2w2/7sGSu1rpq0psYQTIT+02ILS1HzNB2H
6Bf/RxfHGO0FqAAMGjOs0BaC8BZm065jrqQUkxRc6VMkRFjE6PJngXuX13SIkf37
h213nxFa89Mv5lg5n5rZAZ04V7S7WjusgDfK+VBbydwMv7AzvFIeOayIz7KMVg2K
mPYQK74kcKnkoBHoB/ZDQmQshxUf+t/s8ydYXJ8KdcvJGFklQnsojkf8KJpxSjp9
E7+Igr5rX98PnguYT87NlPKDHh2Rp+UQUt9k49CME9pHlYLT4eaP9AVXRnty8f55
Am+2RcPBSsolQD6ff5bvKIK8I/cmx87fTHgtBnI4sCAIga3+md/iITQItCVgh4W8
42gtwfdbFBnqjiOT/kz06zi2N8kuMHnDUWDAvznGnuBFABUIDwF7g3c4C7RkO8IB
WJQ8w9Pk8yjGnecEQ/wsVFH/oM2eIsVkNYSfgP9mevTz1WKcYxmtOOgwVtUpsefi
rqiU9dzpH+nSHbgmOr3bMqJyzl6R7+UxByQ2g48eOdC+9T4uaW/xaeNb0WTiRK3S
SSqROgMWzI9Sge8w9vkQPYnblIGtqZt88gW15KVgfYlBinNV31i98wNS1NUg5Sjf
yE/LEDmLxBLPvXaxlL7ByyOV0Zs7DMoi2T2M5GsOjhSc2Ts47h0UKIOzvTXua9Ok
YUUm5lu4AxHB+MJ8hFFRvVjKANEVnSRQJSu1pEDqDhekVNqRY7URskltQUzTrMH0
xfti3agQP7isfjDlAzQzZ19vKRT++EwUlmf6vi5+86Bbv9wU6r7mB7hvAZruWzGW
ererLUynxdH1EJN7DlnHj6ejPzfdWf7EWCGfV1PxOd1id/pDzzyLy3S9sWf2iZi2
qVLwoy/dz7oKexKMEVO+b/SqoC1uVNeE+K/r0oTunl+WtM1dIDOCBNXHiILd6mde
vIeq/yGcHrCllMKQB18WSnUL10OpyExJwJBjBQFIctGqwB+0AW8XojuYdyO9KkxQ
bMBVEZfMJzqEOkdoSAzKyNezU1+3x7ut5DMVkOyXwmMDTs+ZJELWmOwW3GiXFvVn
U+FdIA+WeDQtjSxf9MKqXiFmpGW8S0riCFKyOb4EzoS0eqULl4Bnm+DMDzhOivlX
nNBneDf+abt9l1mpnsAy/JkVLN0sv2bH3385qxIPLy1DdFcfhm97k40YbtEAAuwU
FcecCcoTikGPpmfQip/ivsoRD7A7yz4ZtUsF9y/2SVOItq4hoI/SdVXzeoUNbiQe
DuDJ5p3hm0gkJtWTqfza5PP6uNFRnQVu0PW7EgwT11/QESVW2m1Cw7YzhvvqozA2
Jh3ZMwpRfqMZGgT17eOBgSIc71Ryl5WtHi+yOoRmgZPbys+Q9MlDC/2D/riX6lMA
Qt4sGDRVqNYOpir7WBXoRhzp4iF21vzjhFNKD2ln+zx8Yu3Ro2XHSK/Ri9roC/qE
TFeYOQC62rqpfSMV4xEddVbKiKBGPy92gzD9gBSTKXwV1/LMPrGoTFBGmsDeDphS
l0WjA3KJLkAzK9C4BoEHp4cyvXVUJW/pzoadBKCw3Y8tB0RK4SSF6ldDvl+9mnm6
kdiW3L8tNpH0g4Dbt+acd+/6Ky2dXrjl2F/XEG9ovlv3046wxfc7KKg3GOUCi85H
03kFfAqjgh1xw0/JxZcl0dpbbKT1Ox1vCq+H14IwQdPKZ0v9YO+lwElVZnqPB5sM
aJBv+XtuO7YAF8r4ouKux+krWbg8/gT352iGzgvpQW6dDual/OtlFyeAdLblQ0mj
gAv/DoEMkUUigB+TlyRSyqFee3qRp5wRHfvLLiBE68hqXFym5hX2kP2tUzY0F5n+
Pktj6az8P0Op5AlFbXeONA428wKhXkSooa2pwoWXGzhnhCXkTKGUbRVayJ3dHEYk
W1YeThDckpapw5w+eFQ5r7VwsO4izeB7sAbwM2wLBxLlcgrqPVxSCmSEsMcBmGl1
LQmip2z2pcZIUAruPdxMvKLOWqn6fZ7hzrqPkbrkyo0d6Lw9dlq/szICSk1axN/0
VpD9gZoUhBtAtMjVcFH1CxRw7gWZQTMIopWtCmgouHRfAXy3BgYPBNwobG1G/wkC
psSeNC47GOBl13KQh5E6vjFfdFbEZ5acmAsu0Mp54wFcpZgwnWfMpSzD9gH4AtyW
VeILdDFjFCvwQfKBggcctWMt/ocQd6sY5+EePqQ70SmyWtNSwebV7+7qsPXON5GI
xkVfOsS9Rl3kgsrX9ma4GtMgnSt85bO9hT3TGlTI/NjTvsplVX10wCmldh1t2CuJ
hGnZKkOStSOmS7OQzlWAlSH55HmF5YIwAtFiTcpi88x1nch1pYTI59+DgWIyAsCE
y/vC8eVIqEELVWBhMxgHfgjsSm2VfSw6aXkEE8d/DkMzJBdvg6Y+8TZadfck2EnJ
XfwCJNseG7Me7zRVv6cE4kpRaWi11KrZOxsN7o3gB36Dgba7oKLavs4qVOgkywpK
f/+ThdKVL5OzAy5sMZ78U0DNgg9oZLe3awdcR/kosWqNQYBwDAry4I5GsvZ2Rfcr
NRXaSn11DgBpDz0yyPGScPD1n0A8O2h2AlklDgAV0dQ3PiocMNajv2ZCNfPDPeUw
dAI1a6Yl4kXjZKoJAKLgTc+ahsMeiD+Vrno2kSvu+UjueshRdtHrTawn6Iff6pIY
lIJINwA9kMKomaL3CwgJ6ZOXPHN+3HiWAsJ7MKzixqMfwpZQFldbMEMwZi6Dy1TX
2QM7bMqZbGcDtUb/3LIw310010cAFy6QKBPuqdaeBqee+3cH18NMcX6drpKxwyZk
s/taJyBGsqZrFXfFvaUTHWc7SPkv4dekr8Sr8aEBMK8dhPL3KccD9uDzVBFh0jPs
COwrANDMfXghtRZHnY/ueFSpchK30zxqdv9g4fsrCHjrXk/Odi+D1ibRWN4CRv3x
5ro8bCaC/bpyB3KBBvl898Bkgix8b5gAMMsZwqUpOxGKO7uUxT0wS0P3QdbCFvl0
gAs0nudvuWav796vfkND+PKhDrTxT4M+YdbB+dQocoyRa2wOs4Dn2DM2Qg6Qjjyu
YltdcFgrvTUXtzn2CWGvSJ6crAzyUT6nrS23s0Gf0zRQerWFYLVppTh5PEGPL9lR
TIT60qb/6LirryWq3lCFxgOCG5n3yLkdmYITb5FCCLU+SW4v+S0UDz4XFwzLjkrO
BZ+Mu9XmERoZG3IArBwumjBpSp/Na0kxioYisVzqUAKFtdKXzz6lQHVwhWvxeUXc
Tuf2nca7Qhp3SpQD7nVAUsEkM0ZMcBNMvnY60KBwHz8bW9lUuB4iWyeB+u1EEMRC
3u90fGqozff8HK7/rCs72Ad2++homH4h5V/zCWOJjPaErDkqNySryBX2T8DZUTXW
BlbgeJb+zY09DaWZdHF9Gx5O98Cl81sKO9uXLgbL2ALNUvJh19AgyJXHu+V0T5AI
91T1vkPdtb6w6cV/UPzUvL/dlE8sHRHhYYXxcgc284SlzzTHKy+q6Dgle80KWaAh
fE4t5acycGq5etTyZ6xFStpE2zPQ8WOA6Zsu+J8Ea7go91OcOm31+9/mXp5W7BPr
IRmZ6dn2LU7FF4U9HSitwNa/Qa6C5xHyVlklH/tpNSPgXfMbcZR+0b6Z6jMTqpdw
gSVV/4Y3AOGKgjxyOuhbf+75oqFaYVpnUAMRiesj0ZYB4tX8RO/d1sugj97WwuR5
YHAeI9ntFmIXCOLXLzgrjSLyB9OVIDh0SfK+UZU+llbFmvDC8Z7O6cjoKXs7pKwp
GRWK2yc68HZ6hC1PUpnHfg+az4FhhNil7vgTypnz2ddxovXi6yX/npsw5WW69Mtv
pAzQ4Rcn5abQatslQrK8I+2bZmUXEs+YoFzt0l0ZHPZOlJEH93U+5dUAu69nDEHo
y5aLj6hUl84eSQGG3bcqv6EX9rL+WoKTjhqh5xJ65H0UpOb0IL0LTSuMHUFcIFyY
KFrTxNopGlz1KHtjJFpkVzCAy3t1TslHyWur8/OUHftzcLj+cPbyBNof+W6SXaRk
TlnELa7DjyoAjDBxXqKTKwsx35ZdM/dWDW3+XP78Kwsno/a3MU1Gysqi9/EpMdbF
q8HypwTkSm6e8VZ1XDXxjFNv56QPwIvSzZWazO3mNrd4q8NZ4QWXK6rUONqAwW9b
SZqiQrEaxJTQ76w7Oq3nY9PhrYQzH6jRCtI/Z4TOtGMthmhUr5+K/ok+CLazobCi
g4VI602jrpjSc3i+wjApNqTtrv52UGdtHIGn8+AooyBVNCjhg7zYaSMZGVTVhkux
tn9mlXegg3D7wM3un0B5jhaY99VF0OWoeHsHLJOlr+55ounMVZPWcOD0iCWqNkKi
F1AlebkkzFUPARkHJdz7vJ+R3zioym/4Ll5G/jU4reZ5piTSnMrUdOE5RK/djwTm
2/je6CCmiqsvNAZ0LQh/UvO26+luES10pHMMxBi5R9XasLsUPli/nhqo/Ya8AjwZ
CQaVD1oNJZ4kLJj7sQhFfaIeZExMJIlEsH5Isf/Iqo/N8vAQUN0G4zuLBn2JLLSG
ASXRa4i0SxEhGKIuCvj+DWuOdMJ5oclQUWkq3T3M7qn1lZZkteNYnUmwvcyjzC6Y
+FvVXvz1HDdIiASwFhMY9okYUNW4C9x5Mn/XJ7pB7TI79xiI/NYkneTTpRzyzhyK
20Jc9G9T/UBJrpS7VgvCr2KzwMWb1KkxsQYbT4aw1IfQsYbZufN4kbEC6t24iNj/
duNhkptZm8iQsqH2XX0nmJJA5H4CRj24TS8vjITJxEm7N+OKUJtVuVY01n8eha3V
Cei2WxlHpTtAguO4Vxdf2hQVcXdEnEl06nywOSfKnt8Ivwj87BYxZ9BFNFj1iIqh
cNshbPE53Wo9TRCPnfaXclVbOy3kRN1nUaDb/+7RUHIrPpJB4DQcoXjbgaxnqAl1
s8bKaROo6AAVzbjc3C9LtepBjjBM3ziII4soFHAGSSaU2l5SSZv0xKNETRv7vYM4
8XD0a02VZglCCcyxgTxUqcWwpS1/U2BxYqeimcQCdPXDX2eny3gSlWkCdDk2hy/t
UXgvLh7Ta4sR9r95Fj/SsZ7aMZhnWKSBuYgmBM+HWP9Ovh0gdiPcXJqoy9ufJp53
HOZEbyZj1jpXl4Umn/YrQjy2y8EIE1o68bADNQiek2MiTOTcpdOKnZc/5uVIJOQL
O+CxoWOjzcpo5F3G5bNLMzR/6/+6e2rn4t8iYIVIywKhf+tm1dSrDd0KwQNKIIXp
7tExanPra8tTMhbTdOdU8JLQdfdubGoVF0oLOi0Ie8t6BBJafetpLDKv1tRRsVRv
A77JnFausQaAvoyZ6XVHWRAkiVc7PmEIzrc47RkSsTiIqycy2x69l/wi9K5x6ZTv
j5OSeEC1KJRjC9UrnQ8U1VDpeog31IG4bi7GQc5sGFqOIgCNzhAhmLiaUhRNgXk0
+d4PLHH8gB2Kpq20MDYp1lO6lLvfSGjVPqfFHz7TOMb6TYJDUeH3WWcZ4mGoxvgy
Xw/A3yRY3CEnxxsekLIpOCNh6aq39yEEm99P9n/jBvF7XSOJP9oERd/symw9aEkU
ICJuMT2uRsqPbt84IWcRqsxzlVtZ0LNakLO++4GeN6IZGWu4SmpqeSVeNhZX8E1A
1W5H+F03ruQ2ql5Va3RTaENPBIFrGuhxqrNx3SfLcYAnn2+//EjgzcnW21UqF5s+
YO2CxAtWLee0xryiIR4HJmDrD7stup1l3pyFNuAGMxKGZhi9NTHqDeIASq5EXouT
IKDQneXqADqAv1eQtUTeZos3lJPEk6OfDQ27suvLH9qNhPWgpiSkG98Qe54IXds9
bS9L+udozMHM4+fiCqxty8JbzeNVQmztVE7yKwv7lN1AqCGihzi+X4LfVCBBh9s7
z1+7z+0Hg6kBu5v4Jpce9u8fgB7dnQNv/hb0ng06+oJLkjQl4FBdbmKEfmBPuo3W
AYn6wDsveSvdJ0jB+elfA+gTrLS2EfwwgvCOQBX2D6gmDsGkfgyz6iVSJC3nWHlS
7485MEafRrEK/KG6H/J95bfMyJms2pIBNCmp9vr/VEgcFoEUjH5l8XRSDzDDGv3t
CsO7hFEt85kUhekjITIc5xSGZPxw0B/jCy0XXuYiWIZP460ieiG3VL7bGB2wSLJ2
ZWtDBQ3fDBDQ0FrKe4fQ1LobcGAtKkhXmSfL5E36KBx7k8hy+BRQo6n5QS0W3tZc
EGhUK2mj9eckigkxE1HG5GhzcSc0twv0V1+EzvtturQjkK3doQfhHbdiGJrHhLCX
3DcJYq2KtMvQISIAoLhwt2SEf9XNn3ynJeEbdIgtqU+pELzvutf/6xaoH18WB+/J
f/c1GUqQZW4+2ZXjovpiiOxEvx1eHoYADB8k+DX8NISgehcDjiF+YbqGifunb+iK
fvquF7aUKbe8dpWcrFnBmoswm9ZAG8zCx4JeiTJ2jtUgJIQrJjNXQJClRn4S54/s
MezqzF8t/O4q0EMtCq1em11YgjBStcRjSITAIjoqYK9N1hdoYSwY1TkNzPvBg98B
QfSrpAkSMJazcxgH8N/I426T0CjgaLdZSP1/wRMfz295ZpIc9MbS4z8Ljc7TsXvY
f+T+YfG8Q0aRZgF6Mz5WsD7vGYuFI26X3V8J93Hg4/pc03VuRC/LLycn6uc6VjOU
SGoVz4VZ1CIW14KWignaB6/95uurUybeUtKYSCeFX56/NLCwGH7A8N9Mtea7wOh3
l+EHMQdOCipDHNG0hN7BYYmo7gICE/lQIEGD8NA5n/Do7fQ0+aArIFffpLuAxVBP
9kbeI06a8kqixLkLyMiyr8ij9p/OH/+CIrNqYtSew6xUMxk7snzc0df3rdHAVUqp
Z0qYm/6bvCrRYYodrS0s8IoKr8mYCRZpAmkIB6TTKG+p9OyUA6dMSYVn649AwE8a
Ikd7zn7VJxTVhubEsx+YoyQ/rVUZYOWQdQp2hxyvsOMPV5B6q0ZnumeUCbu62d5u
JE8c9M/NpAq+L5sgANBXgJAfuaOaCqqslanyL9NUlLGzEeci8jVxutFvdk7gIIFK
Wn3X52qZhhIVgzpaBDSCW04kfjTSyOSVXxSrAYurzjm8KvqHkgEBsf0RbB1HZ0JY
EqRseihhbgeL1Jz23vc7tTe47dfG7ZwcQ6NdQQVUoAX27/oE0H7WmDKyF31q8v84
x35Jj3fHZEJ0PoWiLFcU0n55lemABOWEN+Qebmx9xNcCLTeCM+ytxHYsJlW4jSTv
n2UulrPWIi5SYp8puQ7L5ynbGNIGxfnEKb3LpuQK0NrozMqGV98tGF8e83BpVGir
T4e5aUUyKaxnlIH7dkVzgDx5T+z+oXtcieN/Oho5RK0gCtjc4WFUnhzJBtu+PiQe
CGLkR/hJLqfeHwC+bcMbtNi9W3Bxi/jXb4oVo+5963JeRbSNG8ZsCSLG1dLanndd
4im2FRkpD/aqITOguWMZUA0xkUDvn1FSIU3lXXKcTVNKudCsu9sKb/vAiyPXKqrJ
R1Cfs4b69YZdCxJb/uwwtX+E80Ot1s6p59WNQf8iGfPMQYyd/KgRr0bW8UUSfAws
az8p39m94YXpRoO4g0lJ7YvlYHLI1iSxdQTHlm2LeFxQvt76C+zT92r1UkKUgFYJ
fHcqJ/uYntO314amJMeThLykq3BJ+nzV6LqEBnoetAj4K+8bcxzEUjr/DjED0B1q
VcXuQR4KsKp2OcToIzIskDsI6oHJdRq4Hs+EmX3UIWOSWvTVcs15lO26gEoacRmQ
ROFpMoB8Tv93qCExfviVnn7tVhIKuu337qQQ29ua7pwHZSG9mLPaB7IaEPxHs8dG
JN3Ge7QAB//A+emSvkx72PHFyHzwm8rp8k03u74sIs5qnjAkIJzI2IkIQcp6fnr0
4qEdNJdpHpPPaghJG+WTozawetAjGSYI9QOPaZ7DKAhby4HcBI1BOmyGcQZzFCps
8QhGkwTrE29RZNP2RoevO7pqKEjeOlTq3M4lw3g3eoySk6vRboAk8ClB5d7x1Hew
mK1BaIqxJ+eoDnLmqBV1N/re3QzaVszK6b7jMGic+r+2TxV50Qvk5nkg+Pfi4PRz
Q1dRPtTn0a8bTPx9xvxpDO/RCTQTAgMqfc01B4iocPrraetiCgnXSWT55371Ue5u
9Dw8ObR8RjUJktVM8geb3i+Q/ghxo6eP9J5/WZXKkA1r/naOY2+VS3sC0ixnFGzm
NorC0hWcsUTFLMZ9ZVdw6KR0+VmzywyfU6WnHW0/tqrl4xoCtcQmLLU5MGhEhu9f
rsv7NPAKzhL3BAd64FO3UAHWP97CBoTMBIrjlEtKqqfyCvtfRUWNxzop/KooDQCc
aQneldtOiGUlbMd+g5pPeqQpMqjpVhjdw6Go+hEk2MMY047H9IP5uOZRGizKThwz
MprRb4BtsDLNhDYneGP5zPav9Qs8RoKEjehZPIENZnrrNfJJKYJjEgUGkRZeWdXm
azs5O1MmicctWTQnBC+/jC3zgx8AVS7ot2Yhd08vo1yE0hryOhGMTxCfvNZ5hYMK
0dWihZ+xLvmpe8HUxhqcSOG+NKfHvr1G1iY8fR0Bh1h+Ysh+6jTIrokT0q10D4i0
XjHgtn2kiRnnxEVA6mtbnz1OL97uvCoDvyeeI+uL7DTFSVoXhspfc26QT+JRF9pI
8NQ3xvnP8cZPEiD+pKTmul2t41xUlnq1VLHtRs0k3Ga+w146ZGA8tHLpIHrA2sKm
0ydITFtMI8dXu51jxe2m2MKeRM1CXF2NAX0G3/rBr4Bc1pdt7XmnCjV9kb3eZ7NL
mqNAtvTVuYYA2Asgmak3+Fib+R2TxnSmQLYvd379ZMHPxA8dfST62xNKr3eovVH0
YUgoEjzA1geApbI+gqiZmHvmmd1ISAMFXU5Sj/lAbBFiXCWkq+gjcikp3VWEHmxw
VR6N5pVT7UOvgQD/l0ilE0+VdTLTCCpvPVrKG7LuZm031K7H9jM6AzEHpYyhUjss
IipKQeTyHsc3AZCPwkSF6ynNSuZ8LKCOBfAAiFIdzT5k201u+R+Ax3ILkSLiU17P
QXdGDpevqf2gEW1J2oHMT+lgy/xmZcm0uqBONXAHfXtC6YOH/Jy4b5RpNgm/Pg41
tcwbp5f9XJ6fLdf9+ztcvdP0XgnBiYkLttUu7qJcB7YhNVxwVbxUqxClg5fg+l79
V24MFiCurmzbqOjkYIk2z4b0T5X0xsdpIC4X59V9G6f/8hCMRQ89yCgSfj7yiakm
gz9X1d7aWiubbk0m1g2AsYJF5fVdheJv/HYVkXC0SEYJ9i4WPAS3Lei/AqsYleAn
aAcf4qqx0+NiiHSiv2OQUgtNucbrCsEM/MzYwFDBmEYcpL6je39xmFfpjRYxyb53
Oc6+WKFi5NabuTHl26IpEAtOZWyH/oKZy0AIIdxSEZSvSrUw4/pSHHu5SjUZq5al
HhYKs5T4hSkjdTkrFuxyhbyjO0MyiiNHuTFb44wQ/qhFcq1zjp0hRpEDH3KDxt2Z
jZfjRGViMZd/TNNijXL9vajaYyVD8bVahVvwal15VOcwFic6m4XQdndQ6KE15+9q
iwJEaR7RYUb2zJGpOuFGEVsjYLAuxHJYRXvIUtySfyuywbhCE0exOUBmRMeifVh3
0LrHcgPEXwcv0Z/hrfZDt1MAmmfAY5JAfUmGVnRP1e2cu83EeiR0gm6Ad79AmDaS
hP7w5RbDMlNBXDVVD31lEgRr4YFPJONgxaL3UReOJjwPO9XBmlE0zMDenYOdpJjM
2wmgMbBD49XuT9BdWj79u3M8hXIRJxtbo9D4LQayZPuZnHU8KJ5IqY506UyBFdiD
bPra507jG72LsUif5z8I2+QGQZ/x0K9I0lCjFIRnruSLuUCszd7vdjbJacqLdHWw
9Qm6eIBESwTZZqvwrxTDn64J+hFFKo+zZBkuJGv/RjChp6n6/T67oqZSP/35HfMl
0VgFe7DKZAupJL+pphfaqW8ia3AGIvCyoOJ9XdMIT4LQnyMb8AmXJSmKmKUiiBmg
SxAWT1nMsMPaofXNlS/wPqEz1n73lgvYOT3AHSjuX9i0auZd6XXaLnC8xs9ijaPH
2ksu5LBqWKHQn7oCKRxSD+dzg2D2R8wCiierUzntPerRFmGN01E/cEnyrqawdCx+
4wTjyjqZjOt68smDJvYKchpht23jI07pe3ozTeuulc9yQCFR4f06Z7V+xqRFVrSP
ZGId6Eu8TPFMHhk5HoJQHlk0T8yhYVtlIidAVjKdyaL4EiRW5AazaYUBKqYZDa+2
PrIoVBS5VM2dv5ZeBAtw2yZosWxfxFkW5c8HxARDtlej8kuqDmClGof00OntDaFj
bsTQAREFi3FO3jdASBzmVfTKGX8C7BtBlj9fbB0Mw2u/G20gWLYx4u9YSzLAUTxj
/ragvQ+dT+r4mCcH7MzlMPX8QCwtWmWJlqEsyvGXwmSOmRMnVURbbIdNbUC0eWhu
6S6LUNGNW920/iaoyjVnPnTNzlWSbe8bZJZ4yDTsD1pML0G2qBOvhq4uFtUPp/hG
aq4oLutu038gvYuWLd03ttiVvbzOhgzCgEjjYkYOo5zcBJRHYRZM8p6RlhI4UYSS
by1u5VWOs1LahsxQ7VQAkO5/L4cJzDKkejT4ApK5V1OCFMAVRSVEJgR3M0i1vd5B
Rplh+BbfR61bu9Vwb9VKBEV978kDQ1LloEZzPp1j3Sj+DC8hG3IMIkCHnebfRE90
Iytii+gFl1Cs4Xd0ijO1gk6Ioivh6ctgBibasbOah9ncOG9unOY6LSwfemFwy9no
nrLnzQCFgF4nGciY9ANbntF7Nj5R8n9ABKga9SjD+tC5xrgvcB5qF3vza5byxPIc
sDKWETocGYmrXkEhN1GWJwNz7sxR821JKQvlxTVaySbH8TYdkoS4djerlofmI4Zc
tAEkh24ZdPX/QOjusYFFJsDjU7nsH5KMx7x6hoN0nwwaEwylZfkOeHQUsTOtETFq
ABJJb8IghNduU5Ea00Nz7vbDB4vOWMWPQoT3VyFI83TYXjjfAx66yUrli2WUcq3K
ibfYVDGZwjYhA1pUff4o+23fTA141O7fkE3NqzDXFpXPEyPfIHqnVdOUqBr0KyfU
rh72sQORvxym0i+TLyp0O7usOz3bEhp6hRB+cZ9lj4vyFuS36gQvIlkN0OcjgQ3V
INyCysaK1xd6Z8OS1GOfJ1yqss/ZMHePRlcXvWhXkmpFI69jxEOfqTQX+1rL7j1B
p2LWR/QUZcE8oi4UUON09t6F1PdGk+vF8T2Av7RKPNIT2uCj3V/ES4zC70SV3xrK
G9nKa2WUq1WnAphYB9TaaONu4yt8tnbo1r/NDpc8LMHxB7efk8r0VNsfBcku5THL
02TrK56NasNgKOYlt8GBy6PFuDkowwK7122ybPiqpF74lEFLTwxiE9h4tbDZKCsR
rkW1cxVK5bEKx8ghegaaTyvA0xRrjoxxWdJt42gSwYCZme7ZieKiQr4FJ4LKB/yR
NMAaryG8P7N7PP5QFbtXrh563fFBBmS79kF/F263UZUhSxTVoRAzjNBL2iHJzC28
Db2M/EBsvttbPzH39ga8lHY0k9ISsQXHkQjmc6o0uC4kEHN1ePGY3r7lk6dCsesD
rlMndMOPBdidbApGyMyUjfPCEzJWOiwSgmrgDeOkgbSpoRVjpTqBkNC7bPXxbWn/
ecLGhBBcnO2LO+eITvWfP+FrevadAwhwNuaCswir4dNBHrAD+Ab3uXvcWsfn5wtb
q6OBRIcdf/EusvzYTLnxHqAeXqOz+Rz4qxoklgXvl/fzM/mrKTD5YRo7VWZxE4Eq
q8jnRkBJ7RjjcX8i00mcTlTn47uOTHKq3rddqMe/9+dPBnSzoYuU/alQ3T6iwp5f
1590HtSCPscxDSlCWn5VmRgYFisNlh0d6Hkejr1E0wYhLmi1aX5NNNajKikdwUSP
tsKUuj6QXkaL7DLHPnKvJHww6+ymUfz8/eyzlTkpuzvOu/AMcsCiK2lqd6W2EgI+
Gws4KEqP8yyf+vW24S/ytRkbY5CzJpuwHVb9lGNJiLNIqpruSaDW44VyxtcrAoSc
cRg2igEFYp1Eo2kpghKm6OhXRmbo0qL+b4RPOE/8zvxBg/xHasPpzPtANX0n57CA
mAFJkCbOJQ5TsZMNr3BbyT9XSl0jwqKG5S+BXeO0Ioea0Tw+AiDchm9f5TDsy13t
LO8xebYoJGMYVqBbmlH0sUPuhYFBVS3PH3i8lTTb2I4SRiiHuD89tTst1zY+7QbW
mg2b/5pHmMSNev/ZW9/Se+fpWayYgEfORLf77Q6qcXnYdlNd9V9IFLopz4jDhw7m
i0+juKb9Oq5dfBoZHGq4LzUYk1c39K3RCqZfWStQjPBjnqqCJtLVyy43vDLaQxSC
DsERyGGClPN/z4FN1BeuGGBv3B7ao7ALScEhrUFCrzlHPZVHxXpnOy5fO8i/jufi
iupJ1uDbNsmZg1WVMCWjT2Z3lS9cpmfwJwHT2uGBrScktr6+2+pnF6wXh+peAa99
wTj2eDbMKfyj4BImGxthnvv8hL1fhh2ADTInML8Mw8Nawabx9N5dhjnlH6SuOmkZ
luXS5Zb9a6g5re99kCdDMIXlw+1uQsgGH1GRYcuZTCHzmzjLPuSBiLltIaZxts2k
buUDnnUB5Se5v+t162czB0wY9OFf0VGy9YdefQk42dEOpRlyqp30v5btCmA7Ns4N
1FpPIdGSjPo1hR3bzAd7S3QfItDPb5DrcNriiH5uH4PSKhvH/PvJuH8h6ypPg2NR
HSWXcA4H4tNgPJXy0zYrP9prfjekHmxrUT+LmTVe+CyBs6+HblVSpt9IRf8wImAm
PKoMuBSCDC/ZlXq9PUCSZL/169O0S+M0dTT1csFyyznNAeksCpK5sPC5NMMpp/yp
ibfJh8EEjuqimesiNh/p0dSM+kzG9+2vVLe/UJyosvQCYNjG9i2TdNRQjno1LegP
70j7eqRdOdhBwYcS5eF3MpJNmTppoyjMcZSF2F6UNoOgTCUQy5Ov+ZgI1CXTqonS
ndXENOcDB5aFSOqyxgrmAQ0W4HtvpTrj4J3p2PKxIQCoANfs2bJXDwEXNEWjtgg7
r/8woFbZCMswuEfaTZiISX/QtLSppeX8pjL+d270PY0A+LXZgpdQJm9PCwQBB0gZ
CcCW64gPAX6RWdud4ehOp66jPGCP4EFawBe0T9mffQjpqlJBaJ2N+Sr+7rQbxIm7
TzlVOe11XEHjVhJQr2a0KsFR2X78eFRr8lRLNaax0vS3YKEEcMp6JS6nGjVk+ZYw
fum9D0mtWWuyhidy8z6jeiZ3f18upR852m3YrNm4VGA1GKUwnbOZ6RpewK3GdrUV
HBsijoOBL7I3yyy3yoi6dS5Gf9hLQciL3gtV4AEEV9h6rfH1HvWfycSUnkuIQqrU
Tkogrro3aNRz6qTA2vrk9JIWBDUdDOC1mkXoLCQzW3L6gqsmQ8HhIbk2gge2cZJu
19diju6jhYHGabKpC+LCZvqrQsdyAY5OynrVpJFaLHfgIVn1b+OnOHA441+8WnHB
wkvAXRdE5hnqTeLOhMOUCPXws8N82BPjuSKbsjdZz0QGO+KD8h0InYTUcazzGYY+
GPCod9MXxPRXEX28QpgRwwYpxxWc2HclmjPHM/A7v3LLjDjAkwT4FbSUUO2zpDHg
k9kWOrv6s9dEKpDzilvkcMlIJJ6MGghJnDI7NlEQGLC568ZqqtCaPn7NZJtnNMYG
xoP3e8D4tPDN5opWHSHAodq6mIxMl2zK4zBEyvlrJ4IK0TrATMIZ3mbN+xPhTGA2
AM+Tj10PU50Dx1akclHHCRb/AvGYZHZXbblN8xP1BEFobUk12Sd4nSCIO58HAXuG
k6spLEftRhovBK5bpB/MXb9Jeng3g/QclGmCi4R+71lCcL9B5T7deRy/NNZhgv5v
+if40nbjc5vXdEBEtBLi2Cpc2oKQKq+7KVwlGQzwWHwwlkT+/uETqRudvK7HZWKq
VZaEyRwocdPo5H9/D0g3Hva2V2tm5OuQiTQ7STrqcFqGEeaFLGal7jyKhJG1zIpq
VSRlLQAM55hhT473wltk6QmNzCMf6equucMjCuMjbbWjDdauPE0WnjjbOGlMauPG
gvZZ3up2aw2yoqAtgO0rYcQ7hNDn4gqxK1G2EGVcCB+jpw4giEZUOevhU19kiwVj
xQptgrwSRcwS/4Dwm1N5a2hmDkGxB24Mt851zAKIoF2R+R6ZrkxokAmywC8Ry5FU
SN0iGIEhTXGgspEpGPpyYm7OhgGstybsN0uYHNnMeKWzFmSVYf37ltS7hF22d5K+
2M9qnI1fsRz+nqtNEOThdQlZSB6IdK612Q8mQb+jMaqcbNiys7bu5+m4qjIpcB5W
9qgWTRFfCFMiCjoakDwMKyTOSWJ4KGs9Rgk4kTNMyytrlaPCR6MQCc58+Z3dxi0G
V/Z6tameIVIVP3+3jbi9SFT8TIJ110ue84lxlwZlaeBbjwpb2s0i5Nvy8ALUoDMg
MJAlMrfuYaXs7iPRJTqw/nZePhMGKvkvlCPFr0aV9cdfPoKhn/mVuInCLEr4eyWF
8tCk2DWXYtxG0oLXmLOh2Ye1PzaFDc4OxMwa74X39CcSbprvGOJIrczFg9ddujjq
bBQ6PQ1e2eOFSg2ZOjipGvC8BJpS4vhJgxY9Kxu4N1RAr+BMKU1bas2VP3mMViYt
AJDQGldO871GzD3PRvkTnLYx3A8pUpoNgg11I4tJuBBjvSt1B1j+koWTjaNQ4M9r
GpD7LubdCBIyP7c6FH3NvxUCzkRwoVuT80VmErBucGyOpfOlaSSloShl8kXrZsN0
bWsfb2srFr5Tq05d/zpUPuCMCS4ViFgjBvRS3foG/4GX8hJI5kv2RSGQ2hADWhi5
2j325DDxH6paFNt2w4q0sCrde9B+qalLO310/p1zWx/x4Mighh0H1oue4jR4BLxO
q7PFoZgoEVWHPDKCZXdtFBIDV3jccfJxmucI6TOv6s72SkMD6ib5GQG/Gf/go/tG
AqSSBx/4rVMWFxScnTwF7pz9+zso5VNWvOoxLNf5eZTJs3lflcHFnniX8YtugDf+
kF8Ao3xjPWXum7N/RcvjIF5CJtYS4cWm50hILsN7T2scMlNd1mZ+DK7/ZcqMdWy3
h9JpMfkpXQ6f+ZGr5xq19ippGqK629oK5nJo1T3M6yroVXg8qaFtKWv9f8AOUDNt
o8upsU3Q60fI2jSAr/6mjP8zHY5CDaQFPO6GlqP1Y74pUO9rdmIBfbZmeYvQb8T1
VardW8icdjydSrnIItudFZEUlFZYuCzqrFs2Z9N58Dbmld5PdxzP0gjc/UtokUwo
SO/hGsqo/v5sLytLEl7cg87v+Fws3BjtcxOy4AVjWgJp8LPlG+8aTLSGcPmixCyM
yMXS70S0unACnIOlqHyT1DVk1JanCGfsdvFj/Fm+vKReK8xEAUY7mY58MHjdQuVO
9GuxJ6a8QmE40uCeGDm2tai+PvZ2km3Q/JNrc7cUlRidBJAjw24JAh2i0qwEscTv
155xbgdJeU0SUET+XAKJSyEglBj6HR/utWoUASWcDWRGYa14i/0JNOiG8WsOpZTW
Yx8FMaZIGkvQlybbBkTbMOMckySMnJxRzS5WykLUEyWi6mWoK3iTlyMcbv98pnPF
HgIRh3xLj+TP7Np+2qdRXEE9sj9/Mi0QTfHmQ0IUKbxAApxZw7Z7cu5sjO0liDYM
PK5zdCenC98lie4zk9P4YKUQuAFy36zOco50U3tOAQ1o7SmTH49yL3zlVVMbzw0p
/56WCi+GTnAJgl9JoA79GacHAahsM7Qmb14hdLgL0H0Igv9NcvR/IZ65yADtqDOg
Mu1768FlJfnNfUSwidM/sfFpABIRNQh3dACnxty+pxJHPV4NKtI44ITZpzgQYvEx
QUzpI8PkXoBaRbRnjf6xSDp8GVKva/wy+1W9fWFgnzCi7N076E2LVMALceArfouB
VQl2pswIQN+cXAp2YCq3GMiIyTaiBIheBFGQDV0D5VBhxWQ4+Xj86z++/Qf4zM4h
FO1N3OYN+03xjehksH/fzzdxCJc+FIviQU//BOkhVdKg8rRmr045RMW5L/Y3alZ3
S/uLPogZXh+WSoCsdWNeIbN5k6er0zfrRCJvoqTkTdw6k8KAiDfDUDwI9H9gcPgq
bFVNsxKX++ka+21kemmwQ0QpID3UgXE+ILnfCFVAM7QUx+jSXxcFfCN64gQtgcCd
1MjsaiSgl6WRAMt7zFb8v3ooQEFKGy/hmzGDa5KEQycFGAzsmWODAY0/J+qIKJVf
GaepHQPVQtro5pxOzUDRTXPNlDpaI+AbUKTcwf0dt5EW4tyK0PF3LwXHEHDe+Euz
kWw/DmcMWm6CaODNORHrbn2khHowkvReLrUAhsIcmrC1RqzXCV66e2jTuQssvue8
yvbFqnpFmbdkOMN7kn60YESeoWNPwQAW/1QtJhSwQb65EK0EESPqbG2AMqsH9ng1
nUNyIuhRmTI/xus0uCaR7jxCKVSjosrtkBCbqMwWm66OuUrmtDFMQYRInbvZkJZh
vl95n3pd8kPQhEx9fO77iwQnf8jcUPqYMI3m4lQ6qlSrJ7ksjJ/R3WkAIKtt0wj0
YDusI2maeico7sfEMPUlKNbNbNMCDk+S7rH+4An5Jb6PCFH0Ey8Sk2PoNtW2hys1
zomoFWTQHgYY2vhCOfp/F+i0aX2PyGSzlZSl3TqoCWspbgLMYHaTSfXYqtUqrQ/2
Qakvs3z9+0nHZAnRu0ZEpeJoDmQZsRMdtwwk20bY802vqDhbw/+bBMkyZ49mX8+6
Q9vzNQBKYfog0Q6eWBgl13xA+7Q7THMmTE3cKjEHQSTdm/7so3rOCf8I+bfRaasm
tL1livEgD1hX5BM5YzpisIFor3Alh19n/FDYWaC4i8yS4HOYFbl7G2b1rRsvQnmL
9k04uekgs1rrvNcvnnHIok45rdwsj4uJNspP9qOE/XeLOtJIaX6zS3U94OAyGWq7
IDwTMyNKc7wIPzXW7NG1RwPshL2vWiT/tYTWvy662ufADp/qeIZKVnOqWq3dZntU
y6bRFGPVqJ3djCXONv8wZHhRtoUCYgryTW38GIt1bpUrqKf+BD6XQdV/xEqIA1b/
frvRmmxL98Mu04wjOx0I4arLrUJdzkJZIgIFlePQWpSVC6BEmsxn1OvtZ/iQ2UIg
gkJGBn8S7jgU6YWoMqMacURfjPwv0+KVc9GT00AMnz+/k+XS8feXYcmNg1HTKKL5
EMINGatv1ZpwoGnXIruYxtXzWtoFfS3PmcJ8wZNQBM9TfiFHe9YlnHcLAz96vGZl
fO/tqJpZ3qYp81+e6aTGzUaaHLBZ2I8w8qJCIFesecEmr7yjp6yltzRYvFdiYoI3
Ha+SsgDmaCeknFkpKYY0siX/7+8H6+wqTaqGd6W9prB/wo2rozyD8oStJgaO8GVk
MNqvzqRdxNhtSLV71bIAnBVIxOk0scd8mAaByci5guzw+fehvD3b1ItfKwrRMXTi
o6jIIpcUWi7vG1Myio+VkSrkrV4a/YHwruE1IvoxjSFhtVKQpE6DoPJLHeLdiQiG
kd8YaW7HbZokxYWaNiI//dL50WRoMAw5Yj+/FK/Y6OcOhyrVaC97XprEcxlLwUDs
OrFeKOoeFBpAgPuIHhaeIYOqXV53RZUwSvMIWYkQZfob8MBy0XRdhjMFDumCa7+M
6tWmhPWro0eN3JIg6kDH2uwN/M10SbQA7nIGYc6jKjN9+hhLMNvmYuLrW+noWgX2
ZOsRpGyzQfWXafQ3vDfPEM/dhw2mgS+cGnGeDI1Dg1T4+pcOsi8Uhj7iGY8gCx7M
GgKuZsUVYseaIGVAmDPs5ZfE5pKZ2ulrb+zCDEWxlWUuy2lEJaNrzEb+gC0k1TDk
2439AuT3yo6WI/L8fKxtypFKNqejciBTuI6C6Cm+JlfSiUUUsAEq0IvSinXnPHVZ
4e3SpqhQiQaCmZoySdoUXdtnX3WMCSF+oj1M2vOXvtUIBA1jZ4GSbLKqf7SQ37rT
4gA9qu25TVwCULWJirCfeWq4I6owuzKNQLAN/DlktyHIUzZBdEpOnAf1g5lSZClg
UBFxTJcI9Jk+D3azbDDXg5fE2WORP+NlvXRkEXAydg/Dnz0uyR3TGCjqDQ8FyrLT
GJtq+xS8Ug8M4A6yjBRC7tZzhlxwdH9rWQylno2NFOANklzMNefN/bA+Y34tgOwq
vgfFYiLMcJCKIZccHTRDnXZSArYgoEzdj1sEqnEykNXRrYCYojoHyg2SGfOhzEkh
IRZ76Rx41Tnp/FcROm2dFH0KYOAE2Rltzx033Hv4TkVnGumFuIxXrKQY8MHROMYu
wMgq8SYEN/8NcvNoP2G2K/1Y4wuFafowwvLi2w4lZiijNsYmdFBYtgBLV9/GI8DK
wj2gUMjvDa5t/fvJHGjP8fUO3Hj9SiJIbq70F/+yj9gDySAzypAX9z/tWrUFe2FY
aJuLdQxIryaM8/EEJUOlcgeALTo/PnyyqoBFT5BWrqgC4hE5SeK3P/6jjPzWvIbp
EtBt+AOYfcX7meM1G3c/rjy1U3k0GM1nKybL71gIpzOJ8G3EzXqQq5zMF+/2L9of
eGABl7f+o00mCeCMdShzcOSvvVJfPIFOVM5t8hKLCw45+Ftp2vocKG9Z7vpYeGKl
3CGLwxrUQF5hYcPfWM1KGmrOhEju+rcbMlL9zD+RoShnJ+bj+DTUE2F5yss17deK
zC4AwBg2UsUfPfNxXsBzh3iTsITnzMix9e5Xel1vbbwoEIncUkNsPEFssEfCgJ0l
8buazuv5Ke+9eKq9nY3gXnnOvjxCr0eJDQTaQSQ6ESpbKYbX2a4t/FhUTwBGYxSs
uANm6R9zYacxBa/Ew/L1oxy06xZ9WstuPc/JLJKl3lsShy+wJj9k7GE1IoFS4OUz
IO/FDxBTjnEKAmESuoyRtnNqKYHMUL18Nm7Hmz2z6qb4pAbhvPUFAXo0GHWC+OjZ
jKjVACQrWZG7/LYxAoR/9QRrvxuomB9EeNteECRDUgP9Dg9XbgW20gKPw0tz/KIl
0WmxGdJN16RlY+BJ/NhfZ4V1yQyYz7ty1qSBxdjspLYanRDc71rh4dY2Z4YMXNXZ
qrmSZ9+1gkPvd8zJ/pauP+260OVPP3s3p/EjGkjsgcyBrAZ4apfYHDupkWCwzdJo
B1gMabcoZv5XR3b17ehDx29Bkh2oFgL//uibidXgFQQmONHyfR7abdbbHtdBlkoX
B5+thah091rAqyaZWUodcUaQn/jRfjwJd+hrZuPTo4dYMGxSkvxXb0qcxtw4m3tr
awWFwDWnOdVsu4DBgWQljHf8H9OXoVmN5LWMuB7CtfUmx5F7PzaBJYwvi21XnTMD
KKUV3JZComY8ITM9WRaIvo23pgRCv8zcIR7EwdlUTohCF3tqVH0HvKoBSQ/bHvFD
wwMIS4UZIIjnkwYMK/iZyJ8IX31U6wzjE2iB36qIOaVq2ja+R+awvTmF9t2eJqtD
+0v8BKZV6vSgP+Ltk6VBkqyqiB6MvcM9m1y/FeNz4+sb9WZpXgHn8KALE6iJsixr
nY8IDYEjsyxUDnH5lyfPGvVRBU++EF4Nm9lxYA4mJ9poU/9by5hrm0qW9pdRyIQf
RaolUhpoIP2M0H6XaMw95zN6MCVhnn0KPMKwVjNcBLxGarSCFcyW3y9fFDtZotQf
nqDnnfk0O4VtjDeKgygnraNYn04uaGjpTJyTT4AGWi+6mA2yCjUeoS9tBTG8pIUe
u8UEqoB0DS43G/3sl0JC9xdRYS3wMD87dt8QxaX+YHE+SkrRf4yCWRfOCQbL6wKI
eJK58wMYd3wPtueaHn9KtcRWH8XaTwNuAbNIYryMqOkK9Q1D35NGPeWByZawSpVe
EmofDOWLDdS5GjQ35iWL069nkaQpGXbAnHuGv+nUPTttd5kpfuDWYVVFqE0fCXqU
Qzd3ywDj8RQNAQbmRMwCPNBZ2YeZkxLJzRwsgF1RMsfxra5pEoJahTuhXzLx+Pc6
iWj+CW/iyDhBTUXOxASnZTaIACAfP5ffStxis5I4KKrpTpGNUJpnUh8haWhXH7a8
oDKEhVxhyv15AymPHPt4bI+Yvez1DXNkJKaCpartkubmLENp+1sVzkAeTItUPzqy
pGB+mhVHhFK54Vwp0RHxSFjWyaJIwZSzxCK9aUf2eBnfIdYmmh7MSmPez4+J/2X1
+hSqo3twnO5dtGUm2F40lBOsCUZllW8cgSfXcFxiT0uTn41l2Ih3WAcLpf2YJhPw
nSdiJlPsLj7SDkVqsSAYov9y4Ed6r4vbk6plJYCWI/qIq6Y3lY5Rg+eqOljhXPiX
nHR11ptU0iC49rf9WGfB6w4l/PsFpIyZk/l736sBPTwaAOyrpNosZ+3s1k6Gvzvr
gJUe2DxPPzFmluSVvI2yzSNh+nVB8bVPGnuHoMLQ1iqHhmbmObU6Xy/u9S1nI//L
q8kyK1FsLsG3npFAuX6eOvpReVuK9WZ7gwKXjhn/jM5Lpn+C4IRVLkD1dNowYQAG
KZJ8pZSPtG7rEX4ggndDGocNGcIh++Mlf9JOTk3LpRre0SSkBYKIpWdlsiI2WoJr
WJyKF5K0Y/aYFic8aPkvkCJZZ91RpH0IRySVlkQwZ2afykNXmtWBIj5sUjXAB4G+
zEg0O/vo3F0SMSEIaf+oZziuMosqE//utSKEyVVfKaUMWxdAWB0s3heJHwcqdsFx
5w5LYPIT4H+N9d5w77R+qeaXzL/mTw6a9XCZe1TZ+opQde7LVkS+dJOv576e0Kek
EUg20MLaosDJq/ZIdVH+M/R40KZal/6L8uxDfQgrFL1eIYLRnmjc5hehkS+Rs2Ef
md6Bqaq3PBDyIekue7D3O7M0HLmJ0krdUBB2fkiWkcckD+kIZDt/jHLf3KL9m7nR
ARqdNWkHgqPD1lIK7/jDBuoSdtX2/rm5C24MxmalOBbJHSSn8qlmnH8ea8RZH6vw
I254+M8UJLbHwd6cJAmX86fS0soR/VXgbo8g8yR3uLgDFd75bKV81o0hof2jdWJy
F22x7z/QfhIsrAUZDKiHQqpJrtnh8xSqzs393ydVVGfFAa57g7qs0uxxkNc7ozby
5Cqm7zcrWIUJk8l9S8NSyUrFyLxWr6ck1muqsPOS/qYtIeboG1/UFMHi6FwX9Mjl
fyKdrkM5uMKD7nLpgf3nU263gsxO540J8AIhuXkpJcfYhUUKZe7nq924yUfQFcjM
92IVYhH+FpTHcw0Heg+cunPX6SHzlg5QQWOGxVIDnHA80gIK8JGhqp3DSBbXp9+W
cP1he+1rWBfHAnTl6rBgLGLnc/M+v7ze4NFWiy7+FBLuiPS0vqfJTXaybeBzpyjH
Si5J/nEk7+Tb52lUSqax+Jzkdnsy6a4cyGc63y+kyMhgcBJrsIct+5yNKQnbPYda
V2PVBSDceq2hgSfcbN5mufvdCggFKq4Q4EiTCBOYmyHwcFEnG5uPBboTVMw+0qM4
UyIStVUU3fn52+dmiuqNkUbEE9SHECVuJFpaKxqbFkiRemqgCSqVaw9ZBjUqir5p
wau415uz/8VQMKok834nmTY79uZPwD/nkBDWlQrYMmJYaI153nYMyu4nEXn8s16h
89zHYuM5Qi4O7qfRdzI6Xh7Xp203VOmLOvNXAesTUotDmJzqNcb5n2b03XNHHn10
ELDBdl2a7dxm24Rr8qYzljoH13voNp4cH0i1/Q82Pi+1dGK6shvgK5sd9VGaxITo
4/KzuINj1SykXf5DJ2VFjcvi41ZMAz8hrsKzS/aUH9REMgsbokUgnruFEdEg3Hz2
/3KVedqSZ4TkPItsvCiNjXhgWJIPFRT7NrRQZtW1SeZHtb1XM8O2ncedqiSHJZtZ
RK1xQfRQqIIyhQSZyaTvMQGJ15B7FspCQsN+0JjN3d9QF6wQXkSIpveAWC2r4p9c
2NmcREIzQwLK65qYm6q1vngTikz5QHCmDp3hX8AAGAyzZzNFfG6AwC7AblDByNjm
YHXHV6ZBiJVCtPVeNTufQnZY6N1p1+zgUidnN4SMOr8STm79Kgl+4tZPFniuOxnM
NDykkt0ny9r7SOM/lfsYRUlBVz7yLSmDT4jN0TmpI8pOCXEWgPny94iqXmkXsm0Q
mU89OnfUGsfhaJ8k+YnUrrlSJSUTgZjgpdk8dFor3CsiwPCMUXqsFrrQUuH7lBEF
51pnwQOPJ0p47vOn3gVFUUb5VfZwwoRM1z+IpikbpN6GWD+AVjUjPghRB1zVyKZK
E9vv4k+YfMX+r7SjqcesBQAu2WmHR1rZWVL2eAfS0An56y7A0eL4zd2WVtZxb+DX
ppgVKYK8b0Zsc3wey8IS5zRAmF5ub0TJgl+hxdovCdZiYvzvHIiZgRQaHpqqWoVd
N9lZ+PXxTqvH94v2pdm8mdkmCNFuFzWu8OhoMMFqhZawR9i/PEKVAximwuuSZ2BO
qR0Mf7lMx1XT4vsMOF7VQzAT5+l7YnSKipp8GGWUebaZWOovLNeuyPQh9+/+1Z8v
BqxA0SECJTvPtVx3NPrnkU+PV6NaXqtoHpHbbcJn7G7S/0muYX9f/Ld7VDoELyBI
VgbQcxqCgzHvOi0oYDLBna9UU8MHO53cQ6P319bxioIfkm6WQpN6jbBwpHjDrNbb
jQcrfAYBcsWb+N/HRD+3II/sVpj+CnpuSb0QrWDNfsaIhJALpOUrbe64WoaIagco
vmfOmdw8jGIldUvcGnH8MfdZAEc3TeUKT/w/IPRU/Gg+tL3KXooQgYI20vSwIQ4e
dXh4sXm+CZJ625YJgsZ+A0cbh+kB4y8fjLqbmHlyDBWT7R7Pc3PVhO86pr6T7QfN
AEokPG35dMSj/UNedVXr882TUeUJXk0F9Rqu22VgBmm87j8D8oPqT2csiMAwsatP
rzbaSx9FKU3JukuD0LkRoAIoSdKK+jCGYcJ7lcEDWb7TaBMb9ReNXOs5KlYRsAc1
xxTQz7RLpR2C/C3w0Wpgk35/gEdQZ2r+UWcuInmKFoDnFUwMeYOPFrEYEZZOJyZg
PipBBwXZHRmsJHv8CKDVvC39Va9lEvpB6OqjO4CNet2oDQMpq5+ONdKGaIW+Xvse
8rmbvVPx45LNAXs9x8mFWEDbcGtRuGTXPVDWtdFACQWmS4IBXLjq+4a61Y+mUOMO
UcjGcpjVdVesYI5wJYWuDkvdTfbRpNxKXK2mLVgkoQMLfnsh0Ey7BKBnri348FHk
Nr7pH7gsExPhQi4H/9cHN0DVsu2Uh2k11ZMzxXClP69A+0/pa3ZiK8s9ivJqoo8t
gKZcsYwjVaKcGhiWWFSJUwNmxAAB0omhxD5dnuSsesmpcz2+ugf3h+QrkrfoOO55
2+ZCWP4+hV+b1x/PK7EWKGIgWlToAQ03fXAU0/7Lo5JUgPXFMqUaBjG25/l1QULR
seZPZDFq4GEJggX1LaJijQPqBs3Nb63DNIwSMSGLkL0z3jAao49x0fH+d/Sgbdzf
DTQd+OJgdY1ss+PtmcZ/RpDPdKQRMKkQWmUJAjNVfO2M44qwik3ZxmLXEfINEIfr
SYAcC7leRK8LF/z/Wlk85CBw9R1A1v74H6rlZpmtsWgm9x7vmuLckr1B3ticijbo
Tk04ScK2a/h2Pshc+V7OcXKd+L6NygFgU+bkSJcjZsB4qG/sODSVhDn/ytpJFoMP
zIBZ7UFCEBAS4AwWbDE9qmFlTExYieMsquL3vmLU+NYvRspfa6D9D2328yU3aKhi
NemhR6n76FdyBzbPaL+V5Cb9N+bq8S8yXkpkfBqzN2k+yjYAkf4qC913Op3NljrI
/u69t3EXmBtz7fe4RAJz72xEPBMM1/1CXJVvGbYrn3yhcH3pno8T0QWievWrH87v
wznGbFyHrBtLl47ovDxBbjgzaRJaOhztYQA12bO/S8n+TbQUOw87O72erlT+rKHU
j5pKj9Hxg6lbA2n41pHydPeG/0GL4yofWfle2xLFjtf+J4FRpYBDwoblzW8pLhiP
BE2lVanF2p3B87/P5IrMdZLsBhwfXUc+Qi1ytL9/5mkCVotOWWdqng3G4tmo7/eJ
Z66eoefkKql/JZCjKudJ4jlnzFQDt7tRNgdOqfhIXfKE5cFpTE//aYaNvrqA5crr
9fWy06YjpZMteTTSeVsbgGUequSqZ1NMHcVNGHBVGJ4te+z53a7AluxJZxfZsN1R
JqXfgU24pB31Pv5cH5trLkLvjMH+wsmgMFkzvn8gPsaYj/IChEvAmD1KXz323k5s
iRaqSZac+5igAfBkObFxw574nJVjZsMxlEa5a7gD5zBt/+1bTS05H457a30JpckW
18dvyVi/CC9lDZ1N2zVP3jQPQReTGZlgizqE3A/jKiP8dAX/GT8seRONw/9vWXGy
XkJIjbWERAu+AKXU9vbOAg6ufh2C2tULG4MeyUOcwdhkJU3sO6k+BNA8z8PI9bZY
zWSiT113vf8TpZAOXgnplGtPxUVOp+od5NEdk6spke6+z6AZ4YCxDOW+B9vhXVme
nT7CPzkYCsWz1lbkH7P3ZF09/Q6k8A+Cl5z+0R8P7XIYbcqGNmlu8Be/CdpiOukk
J1zy/E9Fb+a5LIT31cyN01LtTPHSRp87h9XbvTrclkxCLMXNk6Bi8NiNZvKH5znl
dkOAYFxBOhWgaCNqyHmEl8V8gUQa1Y9ANbn123Gg5gGTB6C0JkcBH6AKOHoctPV/
Ot6P44YVYx54zn7tnynwD0DHWMB30uvtVrc0pjzb/ICVRjpfdJlLgb9WOURuIuNV
o9z4HyDecpgTGROKe4dxdO05vKA68HW+yL56BUI8wsvl6fbTZclnNtTLPGRtjlBI
n1KT99VLKvcg0/XCBZwtODjDhfxgURO4GV5WjzAogcRkRvjBIM47kF7jqBkcOECx
yresO0rVdaekSEGB8FwY8wEz1AUTHZKV05Z8NIh5w6vXy5NA6draR+6v8dhTizCC
/tlCB4FXD2Io3jhMv+dY0zoPKrMqXDVcKFe+jiU79BoUpP1xfgrzd1ZHylqpXz4j
2EVLHqbr+zf9itYsHGZVw3B7US18qUl+Xg9vIoJe0yTInk5rRHTQBmUdX+eihB8r
N5Okgh439KMNQbSqpVKrfBFxeO/MxeMdJgI3OsswhZYIrTIxMco2i/roygQtTJY8
ZvG3uZ0bW98mO8fMuihyofoDzeloHZX8Xld1ZS0oFJx0BbSc7FQkgOdejXAY6THd
lvGJLWlWbhrKEiS5feetakudiXUTk7sy87IM3zXZ5GxxEwKmIgzjgZQ2lslxoQp5
LoPSVyDAmlLQ2QQDRkoOVotraXBwQ+achvRAP7nknjmlR+jPOek1W6ulGiP8ottK
W26Yvj8b4rAu6iLpmvTFcrfdS3drIcvBqkAkPw8vfqdVbAoTNmazGBw6L8xiAek0
ME0WUuZNJGxDEqvn/wjW5+BHeTQGOHtUPJ6JoE5GhId86EkAjr3aA5C3zGHRGRoh
kqKTYKZJpZFDvx2Z5pMF8H2lYwh2oNY82VD2Gr1StrKL17k50BACuwK8swpCWYrA
m2q7UhJGaJOUcvjP67K0C93UMMdZeMc6N5UcFUznUGKu+OQeUBbA8xHAdevOQKkk
cxQ2LRBNhD27H36u1WH8AfcMJp67FOjPpiDSDE2f0vqwCcz6mnes7Nya4aukNzng
Wu98UfhhLDlt3vq2NK3KNzZQ+APUo31UAYwCJldCNDeC8i7Pt2UN/MEsCAdHqozW
VaFB0Vl0DQVMnKJDgvv1kFzMTXuOzffzGq/QNfhMHrT5+JW9XGOL9Ux9ehk3knGu
bInR3bWK0PyR2BhBeVJRdjoF900eOt9VhNZcIFduBaNnGiG1Sd+sn5sTlflMQjej
EySImXVo/Y1cT65L/yqjHFlL53z7VvS6vf6zcDbNADJUS7sjPDnXVgNCtyoAaDfX
y7pZe9O8bYMCI3ArPRAPwZoDiigBPa6Dl2FWJPQDruhkPavkN1/veddJvk14PJUc
ef6LGS9FzTFRaCUJDOnX86EcIGDL9qsKbOZGNcOaXEtgxle0C4bGKSS/HQW6baRL
W4Xhs1/KTRByuykJ40aQYzOdOytCDSQAXeEmwBiVL09XSdLBwB1v9QMe8Cdh7m9d
1j8lYvgkwxRonASyPWYqPzdK2A/DOgLD6vhQOY3XzD/cl6Z7v+AM/GRAkeOlyp05
zSH4ulDGrPkvd3IRtaTb9hDt+Wq/W9LrwZKKwysqCseuZ/nW03My5nuaCTRoDLrb
pW9r2fDie54A5wHMVNE2D+6M8SufuE45k1DGPwSwCZLj73ZebMR9R9yXjGm5DsKV
/TTEiOGZ5vHD8IPeg1UGiWca/LAjL3lSOwklA/Qpfc3mLtxPDUhCvZEZIIPJ1gV3
Tce0FP5J7+YQq3asPU6y2v4cLMLfYL413yAi1rViLv8ETBlhdp3Cev/CU1Mees1L
eElqniXwCLYvQmn/YrcS69NCpiuMvqgiU/c00+T2MtVpnL7LMB7qIyt3F6Gpfi/K
jh3CnpfwiVQQArKPQ6CHzD+96UsudqnsfXJdEqawQa2QsIsIM2HSJcd3ggEe/YKP
krjcQpRl/Jf4QuECyYGVxB/IWE5E4U0XexAdCgcf1ReQw5ttXoL2zkptpXD2yvN0
VpW57mvPkZfVQEl8EMKUuD2TVZ8Agp4E2OUdWWLC1DUKicRfXU5wFlWrdHX6iJx6
7l2nRSdjOJHssCWYalDjLlk9MVouawYYvkRou0/HNl2ZZAUFhAm7u3yKROG5u7VG
USZDhy0/RSJwIZ+rfPSwT7Oz6zHs08hL4Aw0AnI4RYbGyhwxPzFCP6GHbhywiscb
veTsOWLbo5256FSdeuzkHSIa/x71igUL9kEC+NIlp2vgstiDUcFBM6cztDm6y9bk
b3ZVRiDpuds4iHVa/GsiItKid2LoWn7BbYdSiG1DDB/+7Hem558+nG9FE0V1edD1
+DlamSIwaNXTo20StFCMsvOhvfhlVdVEP5OTquhGBJCU88a55yIgTB7HxZCOpEQ3
L9QjbJoOMMrnWdwV2OEdlSqpOP8YD0N7d4+gaNfUiSKYtRl3VXbSc4mdHJdtuuMH
WHDIRDDss0Hc/W4x0qgL2rttXLB+O+qDJGks4zLy+JP1bIxw3ic1hPmKK3uH5edc
7l3zwhwx+Avs+9jpnLwov0ajt+YoaVk/jupU4eMI8cYROxv4zQmNdg3sJYV+b0Ax
5Or40cHlRFZdXgKvWt3M0D1njDvdlO7mAf1ANQd0CP2B5lCMcPq2GKmgHIlGuO4n
MtKsA9/9jNjdgOOR13thi1BNANy/c41zOs7Mmh9AU8wSJIfJ7go2Ti/LjroC58kf
2xMVbFKYIwM+WFk+axnpviqtkQQdEI9wj5tNmd/TlZoG3NVyAmEBQWBUVUTV4FNa
E4oxt2wFII33eRygwTK6jJRj6ElH6Yr5YdwE97iCOMCRyfvS4TRL0+nh7ZKbeR/6
v/G3ga4W4iNQj+dnj0wQYXQI00I69wq+0PpeAcb/2J68rj5noRoNuq7pPq14WLSU
BK7xpO33JoFJzlO3+0WM92+IcFkR2TsoP1a2QTC86McFsjYY+NU/WKoACdxmzUSj
K4JoqsJK+YMdiXVa10b4M0z7qexL0BEx2JX5Xs6BGpgRIiJje0Ge59sV5u62/e1s
X2q+nFjG5tYefrgaQr1P9LVdXUQsV0JhNyCa5QdU5oUOzNGmpG7hsI6ErDNoM/41
c0XMH+f3V4qQDFnKJcudAolUJbNV56oZnNY3tyqK1jf2RZEN7V79PQcTRbH2MV0f
aU0IhhCkIFvZW8H7xCcuXwz4LWR60kKBaM0iihaPesUDYW6sZZd9Qhvi1MVbozg9
JiRzGlVVKqf1pLNQobIyhFQ7Rj63XoC39K6ew3mEhH3hqmcwD+H5Cm7IKdsz1nkD
sCL4u/9jTJ90VBOiSYG7eFQFxu3CPfpztDYjiuy8sZ8SWXHlv9jm2b6+XQvPM47+
Q4LqdbC0OLuFEY/plqPb1apR7C/UoT3B1r5emXTvBXucpFMlT6a1eIBCTKdk7s82
hCFNhFwBqwH5I5xlUq56laz4WSYt6D5RqQGHnkN9QBZv2oS+hUJ3ACp5MhupSSqQ
hIwaKlGj9emf7fP0WELx3ntTKjwCxlt5ATy3/rVIx73vbP9MZcHYVXRJK1LCYAFn
GxEVQyO9VuWKPoemMxMdXVucuSZHvY/ywn2K/01xjMaevaEP/aRAoDtg77vGRc4G
ak4y1cYxVApv1VSkHANta3qGEtRLlGtAbRAg/tIH3A61wkeC+gzAhmd3kO6Ywr02
V8sNaEYe+57fWZSg2wzz85KqNrWNOOS8VX7kcxtr+5NIx8NDpO/KbcsQ3V7WlNtH
SiWQD+Ax+37h6V4sF1r51lppl8gex5quCUv4JpybgYA0UphbhnOwDLt7GsGRoUpM
2U7nv+JxcGeDpHRDz8fPToNhxa2xS1/Si1yG+y2ERcPESFr0xhzOWPUWJJdL66Kl
I2ePJydAu1khbG/TXj/4DwX3wP5qVx9Kryd4FjD34JrHB8fqCOg4XbqVRNtjnOWj
a2QfsefhDgbpebEL7BERnudqwkCfVhC0Azwp9n8KlTeM0bX42Xe0bYUKnbUNnPN2
2qypf8VU0DZV96VX36OOcLnCdEh+POQmckt81BD9zwQXBJ9GLc2WZhJcdUymVRXC
ePGEoSwjWrjHZp+6UJY7mGJlyjAZ2t170BHPUAgiR5W959J2c9K1LKtdanLWEYP9
knQH9gNo+GyjnngTeWPN1mUMti3sGC7uStSOjTomSrB2noW7/LmxEUO2IyiSaxRJ
sDVNuRLEIRbQ7hknOORKtFhbwghg1ovqu72IOQ/mjOAxAe7Bg9VKyczCytTz6uDG
diGvDp0oME7edFbeL44YfeqaV8pj/bB3hQHJH3BJhXlrweMOtZxTm8szZDnQzw2k
8Eszq48f/EeXZglYrwDly2kpTUSaKH+nhJEbTqYNVFt5D3jtmdUuNYldito9RxwK
nBfJs14QLoe//tPOz3WT/F/F7O3JCMndRzEIQwyQkxUkQltKOaR2Div9DsTUGoPt
Tz8nio+gDQAxJg0J1SHWi2Rrdvw0P3HOv+ycFtojWPZaDRmlrkIe+T8LufxMFEy+
wNL+F5oR8ejNOQe2umEH/wDcnabrVD2Zne9cf3QU0iMd0UFarrcll3U5Ql3mVJ6L
eChOaubIKTSUaXZhDGwSXW3hBNFLOaNXyI3aIpcEc2UUJE3ztbWkiMOSpDeoXVP6
XGRtDJmES8ORQmmXorFjgTXxsfUWr9nq30dLKnodHenT330OVoVxXCOo3mhrcxHJ
ba37Bx6dpMjFmo2Nb1JLAIxEdimkQ7bhkutVoEeJUmEaa1uyIWhEl1ZnDz7ntza+
leHU+Rixaypm+N/MQAt9laT3JMBC60OPZnommfO8dku8U/R3mI+ilEpZpAPtSU6m
EdcZGD/lnCmfBWdTDF4zDufOx5/wymDv0Y66oG1oS9rXE6VtgEX8rlL0dkY9tUkf
Tmq2239JpV3Fc4XpM7R3QKLpGwbHsPROOJz1XFVYOXM3A0cMxAOjk+zf5keOMFNq
GqPQljbfrZgjdMGoXpb4pMohbEi2X3qEkBQRgYbWm7iTaws1oxrrnHn9EH9Xf/jH
uYCV+nsDBRn5sPN+VAiwNEMCpLxzCpjLk5AvGuPuPEhORmbvodhmMHRJSQlzAiJr
bpwnG/SlpZmPugBl7PqBjjVRE+njOd9VRxtlX4hXAxftxEKl1NlB38QZpdTmd3hK
3zyzNy2URt7aYDSIk4ej5+vfV9JpoRrutYHxR/BlD1AL0E3Lon/6pec0y9sDo7qA
g1Fc/YtEa1f2CsJrqBgjHqtt5uLqY4+sYplth17Xm34F4cSlbMqvhACF/anXKb6O
6S14y3siyqJNHWA/H3HNkhuHlD+nQW6Te4Lno5i1vERGphsRrWVLRvN4srdN/yeQ
/Ck2+knk9sOk6Xs6mMbDCPUcpaKSzxGa7eaaoKRcgMukn2ZkkzCOYDrUzQpNrJoF
Gbi5acL2+Qk4DsY4urH4GxE28866rLPc8DK4I5NhWgcb9hOUsKArfxAC82eKXrOE
uDNUQhgtVSAXpD+KtvEAPYYD23AmgGcxxs6ZlwJ3qz590JGuS7O93rQFed2Oe7jS
GMNop2KgXsrjPhMUVAz0iwZyx9iE3t+fX++0Tt0tRGD25P7Vt1WEqs2ozxRA9m+Y
NDzioI4XNGdj1YNkBUtagCkpBVREEtCmVEL/au+0MYZnfB7zq9ZjIoKvXwtYOehS
thl7znGGE4HRjIKDduR5freinwplUJ64BqM1FMCRQ+gvPFhmV2bMtej3QaeXkEZ3
XSCEGg0ltmhV+EbGf8ICtfR8iJlDZGmAbll7b+5mYQi1F7XkmsWDf6ZvyO5/0GxK
K5YJIrLSGBit/aYe4iA1N9dKEO6Tv3HfJ+PrO2f4SxXSKTOPLBOI9rviaCmKLQw/
Cn8TuT7JXNns7/XDDddl29RN1r4f8TIHP+4lNF31hKf0/iWVthnyE/MwD/1dgLky
mBlGvfGah7OjFKbu0HZRc6RTDwJ6gPe+Nz7DZKFDoOaAa2MD+d0ANaed7I+3HdZq
sVreTXIn76mGKGb7bOW1v/fFJtTkEbG8AC1tS0WuJLIoFB7AeytIG4oNNUYJI15R
dLp+cBKfqdou5uUI02gynMZoSdybZzRsAIAkBw3QDxKgVgUVKZQ/gChVpuif1wiP
MkzPhrO2EiKOY44Z1xT0tLWQV1FMF75tGa4ktUCmi0/m6vEnaVAFITPSAiJuFkcQ
OKQTxdldZb+F4Z7hWTOTJ6olYVoZ2ZArrZS5C97R3ocD1X55XBihQKo/y2wtw3UL
C0NORI8ya2/POqby58PFfZuTKjWvwND/gKxbXdpRaV1Nsfp7fDK1A8B2whrgK/ka
k1T/4nfryYPiJ7CbIrQpN6fKX82f11+txqBoZ7PPTKsxwJrWxRLVwSi8nGWmyoot
YkWAJ26Z35cyHN015p1xfBK3VcUuORr5S5LBmzC7Ew7HTLficpadl04OE9Lo6hDU
ve4DKoccT9XJ4wlfKFMVgSRUWeup/82sAS7J746429efXac+r4IMIXW+yeJNmLSX
9bkna8NoAsrL2ZyDi3EQ76+FXFoLDmuZvF0eW27xK1ofFcbp95lb1e0NryCTgpd6
V95YBECfiWBP14rapJoC0MEhLaRw7J4iZiF5xAAOXJ4C/jYt9Y69/121PU277d7W
AcqBcG+gXyOIiFFXwOa0XiJetcS3Gt4j6LAPBpLBWmcjthtr3UHvVkuCu542KS4s
HEpmmwd+U3agG44HUcRg+3zW6e1C62NpBxMp5EapazyQTKEztmTn6t1FFl4iJbZw
XhvfQGr2d2k5mNkWRQVk6W5sSNYNvJ5xEgjrmyK8jS98qjGOuEuv1cjtWcmYGrYh
zLms5uig/fxtmP1h/2W6NwpIMi7flSk0fmvYOPTF1dPG6DcI2d9LBOQEPqmUFpMV
AMdN3QqCgE7zF+hVTs3MC2nLQYshF7ekQEXs4Cvx8La4Slcs9xYz9Ooq0m96I7iI
KWMx+ckCyurYfXyHL+YFlVpqHnd1xEwRrQjL3yQrQfsyPkKKIYGTsfqM+4aUmhfJ
/itiwiiTAJd7qCn/IKl5pZ6NWcLrAfWGO4kaaz8Rl3Oziek1NpuC470cDyg/2lW1
hirPrSguagUIJuTunuvz6t9KTkEiv1mHd1YimgPkmzbfaipT3QlZsN0iqkCCS0IM
G6O+Fmt05gS0aHUh8YrP64/giBUp4dfcEBHKqVzqA3E9Xm5tR7EaEXdqPdcYrmhU
aFD++E3DQYbj1J2Da6RWz49N9a2fftLY6u2qcs5h8ICNuUnRlZmV7LbptHqgFAAB
q6m/pmd98Xewr1wOMBaAjlmuN2dRWKJYVZjbvlDtmXy1UF49ve+7tu9de13ZX8Kw
zbziP3SUSHdV02ZXSVhpXlh2scn8I1UprxFgq0iyEiKPOC10ekCvkYqVyrfWycnS
oVsWxJXFB3eNiU0vxmaeP2TDojryt8uUkEA0ptYK/hSlswZQFiLQhtEfmm6smi3b
gCgmY2JT3wvI3+kYeD8o+4hMNWgsJy6AXk7dt64E7/RfYJN176fjy+aodEYmowIi
5bsMU2LFpoIxYDULAHS+eOf0mpbIL7RJKqvzFh7+/+9WNp0V2h9Uq89GSswQgAWm
Ha1aksU1InqxYnZjLkyKN64g8/bD99WTtBQxizimrtrxcGq4LQ7RaD+mIMXLA7nu
8XwpTrrCBC6nWk0OILWefQctHd/BS5ttR3alUP/+akJSb8KywBPbtJY9dtyowiz5
6eDaIxWb4mB5XvbiRn5+6L+dHz2RtcqKnvepsEuYvlyOVemNotOuudHkVZpmw/si
toEswaD8YM+EH0nXDh6b3X6J56fkxw8GwBJ6Wid2ZI1o+QGmm1e/8QTYNFXWKMJR
fekwPidvS8FdpQfB3uwmqzVxkedDrojOzIlvyyNdlXgyZxE20trT9lQWA3ihmwkR
yhYXoOTJoyYVEc+ago+7ttwmpdPTsIsBu2NZwi/wVEOtdt6EV23vqEbR6vfZ/tCj
eStqnCzsvr7c7OLCID7L7u7epbePqZAg9w/Bh60VHh3RhkmyEi8HzVWWqY1S3/Tl
6vvkPkgAaoqyUj9AUSGgPSYsWJV4a9AOU+rAg9IsBaAB7xZd2yJ+fMvwV8F8ClKK
/eEK/K5YZzbul151mZ6tEoGjQnb2COgLUWvx/7z2X5ZasCHbtIs3p9wQmAQ9j+DY
FfbkgmeouE9AYIDOvoSdz4yclNQ84TOTdAmV5ce/ly3Rty4AqBjOBgc0864YHI0Q
DOJ4stF9poeTOPTvCtHLiCz+iIKjj0TVptntIIeqQWDwEg1zm12+cddJmBMnyhOE
NyforZHW2sxNn19IGCeYEPhCWjqxzxPjP43Rimtj5Xn6LqY9ZUxj5OydECv65ykc
tFPBjWSQ43lThSarUBDKwOfautXyVJv7270ySh8gc0nKgd0DAx9hlMNQWQpW09DW
lMBD7sYKDv9ou+WlHq//3yaMeNhFXXW0q875vX1MvjG07asERgxSYBdwx73JO25+
G3n5t5d3O0igKbjG73ZXsw/7alPI2TzIzf7jWuAydl/T9uFQw+krwk+5CqaIuW+w
idghGrT6MaamKIBXlmJTvWG8ZkzS67KJVNXfD1A7+V9FRZBL2QlsATs7NqvK0kpJ
yhifMv2MzxTOPvBTGDCaJD7nO5XLtHLtRc1hoa76MjJ6sGLNM9D0YU3XVHY9lNa4
U4G3Y6x3NrJvOyg5QRhpLgsKAs1MkYJBmtxriypG9WBpSkx8VEt8uX3TA2U6+14C
cOCVKsPlyKN81+Tvzbfl23lKxm7KDnRyTZzqah64GJKSZIulyd3x+DBMsAHpP99c
xEj/YoFR+BdC5r4TC0BznNLyemvBSOSj7A3SyUcumqZUdKnopCO95i+Pkawe25uj
KZniGJBqFAdTOwTTZfpVGRnHCW4JQuR6sfGNLM0UenZygcHHqv13e1IUXiToycAE
LMI0EFZOInCDc+WwymH1YVMRafXjDr+YiTElqNbM96BairHIeDNHKY97v1Pm10Eq
aUWpQGjiFBgutrwJCI8cgdYA9vSrLDM4uMDDYNSkJ9l97B51G4/LmRDy8WqIl+2x
sGe7stChShSKxz0BUcMagvO2AI2uT2hkvZ8CRRJRzkeOzKw+4bWn4VJAB0pzbGqt
fXcbsV6Sk3kHBPfGbt+VXO7q95YenQlyYhyhtQQExXJErr8cSJhYNUSpNNBkNWoc
m9qcev/6JSih6o69mR/YLNaZPdtkCh0ATnbuIEWhGRdJ1LIZ3tYfTq6cgKhyXwv+
BR+yQU2CiX9FBEi0x5em3mwjN8EjTzQm0O8VlBlFerkeeApo38J3oRjT0pE0sc4N
JB7bN3Uh8hlol6VfjnHBjjhlaQIbJuZJEAME4S1o2gZakfHdYS+fLqIGYWWYOc5B
RZ70AW7StjgASNOF/GEGVOGIAXovspvIXxgBMPMzLjWnll3d4qFwd7XcQlnGKr0p
0uJH0JihKpH6IlQEpNXw9TG/FeJrKIi5So7SiXPEJiIWgNJKE/j7SDi2ZoJ0tzPf
2WRly7vJ9OuP3zHyfPg5O+0VF+LyxY/+iphHpkMiFubLfjaEveuGx1u+OyRGV/YZ
EHTmqANkzTY5b7/bNgLBIKLJhc6a4zX4V+TknuDN/Qk24i4/bScou8zDpfw7LySK
pyTzdaynPcRvgPJlVa70OCEYGfubagWzqKonan2cBxyAAipOqbAdXg7hCMtuAGFP
vAu8c3BTBl9FbpyKLapU06uqVV1qDP1F3R2KZxbzf5JPdHyaYsix/kdyuaUdI5GI
bOMg/JqP5Q72CJNQaKH+qEriNdP1HD/fkkPYjli25MUPXGp5aL8OkJ2Kfuwmd3qU
eXiy6ZRia4e4grSqeov/lTT058cEDvwA0ehGBeo5Nu7ySTZ5Pzn/YtjpCa9I/vjk
oNIJqEmp4YtlDGNQz2JakLvmi6Z3B7UkYjEsB1agaqhH6A2z2RQQaFKdJZNdxnGq
0uu6ZVG8UIH+BXprXFd1HYB2vQVevgKbwfIfI1m90oMgwfN9KP9KlUD9v4G9k6ov
qjEBFUTO7BMTesQcqoTfpyKoS/L5naWwoFRzcfHCDd+WN8WulIoQlzw5FLvyetfn
f7h7E3s5g5gAjfiA/EVWTUmwpcX9SUni2gkI/xAM45ZNTR112NkYzqfJosXmfZrz
xMnQzBSimvpNmDhwiekXDn6EdEK43jiOXZvL4I9eW/INP5EXVdQExY1mRwzm5+8f
Xs/uYvpjRMPhO07IDHpV2hOkO8AjrnMFrfvVWmthQWC9lMjGMSmjB+mvwDnu5Ll5
xDW+/JPqGSLHMFVp9Q874Kkv1hZEsn5D5tJv0aGshMqiUACiw5pLz9vNu5WUvsm9
d5vVfdhef8JXT5rjSFZwMLYJcYaA0YkeThQ5fptk+XGEtjCxYv+oC3DCM3lRs3b9
iJJMWPXBjITnUQfaJMMg2B9qQiXmpskHfWFN0UmFyC0tZoE9AqF3gF8296m7qLwP
o7gBcYxxcO9ZGke4Qrcz2fzwqJQMx0tWLtT85IR27ED8avvX5astedNRSABmxwAg
HSxESbtcbEq1bhZOwYjToddbJ84kmPTOGuHSUyQYkYKDEP/7ajle5SOieew6LjSn
ngPClLYcKklBxgjE57pHS4XqGDYK4pp68ysl9NREBEIdm7EoZ+V2pUcH80l4Telf
3cvwKPNA8Vsmxjc9RPmqcqPg+949YlgdId2PufPOC9R+e11A1sZO2U14qiMRBOzZ
vLySXb9zL+VbPQNsvumTm7s7loPx807/BiJ05HF95pa7Hxe3ceVjwRhFrq7jmJTC
7BOw0oVSrLixjUIgzG9uhiNY9erdCG7ZEUF2yQQ6+G2ggOyP1OCMFM0iOcPa4TX7
4sCz6Hzs4FS+G5x4U/EnCWpTStXVDvF/YIY1JPLAJREzOnadY99aGw6F8+5DEl11
FHvWidvuUqwEPbh4Ep0x/FpQ+u4jNLs0N90nRMvK9MzrSY8FGosu7nxTDkMyfowG
LBmOnKVks96xmmtoQmRy7rM5BvqJ2+A2hazkBwbPfyRmBvjbku2yWoSf0DlZfN4J
SQ3I15OHC+m2evlBLpnQ4x/ewliFXcY2COSZ7NLJtQ3HknFxv7Oqt3H4175KYt7S
qG6M9Gp+NIsQ0bE5FmEYkrZXdmTDbI0ojd9qjkiKcJC6ZJ+4OKyreL78sOPD4ul1
cXitJ11fsT9IeRJv25JhN5QYMgp0lnxSUPh+Y52v18YQPXyJuiyLVa4BqRqmohqr
IUTdt+9c5kLNgGNdZPkmzoZAytVhrlBnDtCDKADKFzQM5QcI3mvj4oWT7F72iNfE
H1tIx5gKl5a3xKM7QKzSDaDfwKBF74R0DJZRF1H4x3hgPRm+yn9iC7dAk3joECW4
uKNuXTMAnOPA14vg92uLFrOE6H2n+xYdgZnM6oWew4vVOiMEGNYeiU5CHzdjzjMO
ImBuLyjA4CbyWYTcl1aIBrZeGydqBYSNvJKop7omKUnf6A2Wd8DFmBS3cNqXJYNY
ceIZKgwE8Ycz+2NKAztmmNGvIpWYoJmTTWRj1mrSg+Y9pASnIpDaCZ5JTqTVvTnQ
7aFd87JN4dQu70C8j2tCJw9phGry66Fj6vv7OcK+/xdwhggs2zdMRnNTIIwZtqTo
aG0zJR1eufOm0MjbK2cd/Dbwm7+n593Lcjmq8RxVYESTZYlnX3/Mgdiz4p6uNeqC
PK/OCtnELbk++fqLAahJF7U+duQ2H5sNE/kxym2g99MctL349aH5PjrX4C+azqit
9bMjZVuFn483DKJaQ1U5Vv3vZV/f6yGq1RLuqqy3yVp2FGjVsC/EqSt5z0zLrYBy
wJs8kCi4Zscc8s7KuuMRuNx3X8V/mbRmNzM0w/UwxldhwQ8Hcmj++1/HddWYZWdj
a1PLUpW8OHlaqtb//nFe9JzpEzcFRbEaTlRvtGaf4AkEwP/m4XWKY2e5vg0XUJtt
iEyxrGKiPRlC8eJqsmwAYCHefFduCU2Y9Eqlr07pqwjKmSzJ+GaGs1/6mMsFTCpE
PYMBC/Y0Ec1DQ0eO4ZVGXiyqi0zOaMd3UpyMk4dJIwg/cyECCDpPND4tr46E/lIV
OY11CvLtjBq8wSl+OO7VuGS0OklLTXYVKLMSDbCzW+eofxvek69KktukqUbaZJyZ
WZGjSjelO/eLJvJuByYpebHHNtVkRdvj7H/hrgqxl2YGe/mVSFddKaYJegDICRlG
u11Ql1aLZVUIRl8SC9Fnb1WDjGvgSlZ8leFgI39wIwwV33Sy0PazcPTSuJmssZmd
GjSwULNfo7+I3aEcs2Yjsq+K1Esv9ilSVci82wKjwnR2lNJlvT2EeM/wD+PyKIm9
KwAqbwJ4zYy0qNWTKMCqgaOS5HFdaRWqXT/2czcvmVJezUSptks2kMP26ROQcFtk
EdgQXNhwpDGbhpbjzMUKjI8Seg9G5MRxb07Cy9OiLpO9QI+dIBwN/1xZfRX0+//I
AZEHFLUJ+TbhnVNUyTCGssBDC1NCeZOjtSGQVAWx+UU1rcEdTK8m/bOnbKV306oz
H0+BDoXxPXRIDHElogKelS/2plYIhhOy/akyOx64cRgYDpA70DSOglTeOg5C+QJ1
FoRJ53KxJO6U3+MD0GUwLTTnsnfD4S1IETcuayYtqFBto/JIiDiZEmcifNrLwxOB
gkkexwUy8j6YZvjYBPozWnWAR9V4Prz+ObGfPoOwvp8uxJ7avveexc+twldkowNn
R6H7J8zWw7Vro8qDkd8F9DlBM3JzE+N+AcuKb38jepLIW4gQRH7VKJhInLQfBjJK
s7mqc/cA/+xk+tp+zF6Wyk5Hzfc+afwAmzA1d34dYY3exkxYfkvcYksTR5MFmfOp
VkatjQoyFE4tQW0vfL1X8aaVE0joEGYEwL4SOHYfyjI74LSWWyvLefHilb0orqB4
miETXlPMWgnlZDCcqnh7oOtFucFDV0KKOhQQ4s8X9+fQE++CE3yCnnH1fKqttQlE
QPzOjlLKNzD0HqAIGi3HbU5vw2WepqVeesmYq64tczuc1dInAJXWJueimLYDea34
+AdHJHU+87hnvb4uWSOjBP/xH07IMOmNcBu2rUhSykoTl1ne56aFeawWc5CdQql5
xmbHsBUlufQHthrTvQeAK5s4KAY/Vbr7trvi7c0oRlCCFoWVfU7wqg4qgYCQHPwp
bzB75gVZL+puo/5BRY2Xz7Kj1a+YOVyZ7xTcjvrQjzYXGEzd8+3EjUWzEjOP2GFZ
kZOwc/b+hH3xBrgGNKGW0w4St3e4W/lmk9s4nMk/ZJgO+qGQvq24MxiNIwyPpNCJ
/3+6z914RaURUFz9bSeo3cekm05sUdpCpLH7XCknvZu4z9Xxe2A5hh6CBh1WYnIw
ymjg0Tki0fyRu82dM3VCD8eXHPSmAFsVquqozeXCHocidcxwCJuZnAukKRmvsM5B
n7k0tNiS68HRayk9C+YbcfeqBdLGdgusOlKKbQKf9tJOJrntEOq/dr+C27XPHTsa
15K+n5McAkZLkud8lj9x84v3/X/6j081ieAdiIjauY7de5SdvHdtIs5FYxPEn2k2
c7sm9wHXRCJ9LuGMVZEtSN/pA6x5k71hkmUghS1o5KONZp12yLJ+qL6SL90aSN7/
Tx5Ud968Fqq1rkB4OP5y/Xx8O+PNAjfY6O7f9dk84bxxMp6L8XIFPjAF4llNsz4J
eB6oeuV5xUIJhXSMGYFbFq13cPB43JhpiEj3aQGOTMiVc5eKrdF6HMbMiJbcuT5g
tuCnPVqMeBMBlv8C0F+kT4Gc3UGXOSJVeS5zWTH6rx1HLFWKecLB8Cm2vu/hjVTJ
NIgrZuRwxb6mHSd3CIHMHirSCmnpsGhCYjErDB65IwMUu3wd5nCjP+N1RZS+gpU1
CkpT4vg5EDpHT5lDQuZ/W2hkabj5LNHB4Jr7Oo3HVBRJmJDHzeC582u4odOC1AsM
HIqvG764Sq+fDzwyrheQK2kHpT+mtswTCn+Qko6alztk3LX1qYBRUtOizopup7I/
7+26eaH/GXKpy6Ws8Psa8upaVgKjP7CFw5IzL0BiT6C2dxEDUosVXkqcAdWq0APy
P87gd0d+RQHXVgEc0BcCf19DENeKNY9nfS72H5XwSeIzNgKUvtRWHeXeOpNP1iBa
R1QDzAhYw6HqfiGZBvfAiXFsgZjlYpGJ7WiOO8ZfGSj1CPg/J71VgLg7Niwizlno
mW2gd1bVymwtL51zKe/qHXTKt2dZxqwrZ1q24T6Phnq+ZZm4tUb9UI/4/yEQliz/
0vdSk5Ajaaa5yWLm5KJyQSMNB9Do3yCBg++BY7wSRfeMkiQY7stTqyLjGzSqxu7a
3pP5E0f96TpKme0ee9Vc2p3T+2/NYjQ7XIamc9p2NAKrEeoQaebSbEQpKXObECLN
VSrc1tIfnjXVKHhdNbesUxMrOC9TnpaL+puvuFo11kr9MrmfNdth+L37xE+C8/kT
DDlkZCHM3bNkoiPCJMkTqwhp4nLwZwpIapsWCTKJpItLrHKtuZPO+bCOZguVynhl
+pJ7Y2065U8V8rtGTF0874ziSsts1au0yPy7hi+2EcXktiBdHDJ/myGwDAvnlIyA
wuE39YY2scoPjxd6MhIikNIOHyG6iJSWErpcO81DIAImJ4lKVVKfT25/tmlstO+Q
KhVShE3OLYJRV9IrAg7ChiwqFkcyGstdaoNeAvecO2BbifVy48p/Cb/Zrleq5kcq
qosP/H0yCereza1VhDKDoPBha9Zk9v6e+QtDLLow3GjcIJwch+huHz2ub0fojz3H
nKpzwyAhyB9S2bBc16bmCW39wY2jBGxr690hjOHROUZF+IdEZwq0EgGfVyeNqTUo
u/V4Kf3DmFeF3AlL0OVSsHkCg6atEXevPqMATGGrZhkmiPBegqVAkE4M9VkizxFh
i5coZM53qtw6BcNMLitJZ9zHqfjVJaC98+u5/AEoeaJFdMUahuJnH8zoDhRsAFt6
N8FmfZHye/mCRyeTsWdza1QFcm8NeJxZT3ldeetMFeX7pzRqJPtEf+k5qBSzxPzu
y1yQDX0KIFIrWe9NDonNMJHIwDeO+j/XoOOzBhs9FjkC6fAJXxeb+SjQJPWjEEXS
M7tkC/YDZGE232pi5K4OZHfJHHSZQjSF2L0tvPT1mvtw/IzDpt0IOlDT3BlWy+lq
R5FuiBDmxQYB4LTXI2yTXoLkkvFcY0uAB8P9NaLIHtS4O6GY3N+AjuwhIiaFzusS
4FfhaXfSC7jA3u4quT6DULUixrnfJZY1lTJbSqScH68PLZ3I3dNAZlqXvweqGFRf
8uGskiZMaE0x2eEO13rNlo0peReqiY3IgsU1VJOR8I30+H8u6AgfmYTTDR7gihla
nF857ZKQ/bUJcCtSCWwkGIpqMhmzf1P1mzbtOso7qoZm7AJxcCJWN9owfO+o12Yq
WwAtDPSZoEggvoMONcQ1oNmGdVBmR3qolFGIvri3QAdNLYBMFVIn1Zghr/hIhd+T
yG/+Jg2rNVEQdO/s9/mLc7VXce3k6NgLNLV1uXYnmdKsrHQz/cOX4vLLIJKF0r9b
6fGgblZm419xE95Bs1JNXNHwbE4h/39UoXObKY/IGNsBzw2T8SXBwoACBT1kqJjJ
7q127AnRK9zkjFwBA32nHrt9PWMoRxiLoL4kxxHZUAROLn/t1oUFJXiilP7CvCex
fHIGVdxzyV+I1xWmvu/lNqyKVJQZrNW2GMXHZ+zT+MPE76FW4fcBz7BfWNSi4zr9
3CwjRyaRPcnhgize2rq5DSalkqqJB00I1QpPj15oERJ6YOhrlHBrObHFlAQTvJmd
/Vzr0ji2Z/6EBpLWcPOwDQrWKrYRU0BtVsjHImVYAq+QHAjJJsngn0HTHHuIENhp
AfN+rAp3BhNf8hTj5nMB15czatmhqlpM34TOLSmGDV07EgZKd1S7gq1HHTCijxrB
ShP9jqA6Hocnc29LRMNDTCPgBS02CXDCtIZ1vbnGxTWNdW2CNiC4QNFq45ytlFOf
NtlN8pPAQEbwHWawQRGk0W9N5OJK8m50SF2BB6OPARZVSt1rcqAQJYhO+LzhvkDn
VDgSfgS+Y06gYZWA8E8ymqOaZD1CDlspctAJ7hMTucexJJPFCWx0SPr/j4a9y0o4
bb91ArtN3dY7QiFvmsPnJWvXhi8POhVtDAVpy8IFI7rFCcbNCkW2LSSgl2Zd22wl
Mp0JPwS7CSbPT8nI8ljN+aPOtUVrq/ex/lLJz2asufYWStjDAn3Sgb/t680zbb36
FZ8t3TLhWgfuXghjXUDwxmoosadZZmQ+BT3pM1tr1LfS/jPp32Vy1YDo/j88KF7T
ZaTF8WkRYZhzZ1wkJVr3qUGB3BPxJ+g0xSncYmeBFoNigVe0MGrJbJQ/ne4g9GZ4
8tCxi21YBI/OnPqRG9miTkpVySiakTE4rev0xiNOPF7FO0j6v/RkUqO4tfmBu3be
X2S4jz4k73omdUWm55hjw3ulQ2NePKxAqg4HbmGzbcW+XYzmNpba3w+QS0JyX0RM
AIEvgts7qocJjC03Pjjy2WloEci2/1e+8CPeHWGzNma4+i0pdL85MslHY11oyH++
yMO6+o1mZo1y7fDOYbNlsPkbU5ojLbVRdSl9OdUiYmSo3y/UXdi4J5/jeqsc+Uh/
k7wKnb564iCugqWcOIyYz+H61S5fkVJgfkxIurdDx/+H5hH3gM4hVTZqVpBtOcrA
BrDf9pPat6F/9JvYX+gu273kr5flEWJOsIM+7fhgZroAUQoB/LpdUSTUCWhTxwgo
YxEJAwPisRk0bOnaAn/j8gkMEHFQXqvz5sFrkUNFRKDSHtNzPQ7085eGJ734lLpH
LJ9OT05dZADX4yIK8icvMGuxYc6oUoePAeC8f6nYMOt6or2/fdLTXnBaao7nkQCJ
D3Qh+c/hdKrCg0yqI/z4SaMHULCXsz6T6bYsZE44U/n2M4Bsjg6r5x9Cd08/HJ6q
Enl7N51VzlyxvBqmOfEPMVlwcR9o246UkgNtiwX2gCMUiYYyHK3SWbEHwSGyIfVx
+O43wY+HH4nXyuF4pZJecxH07hdEejblAwNsaJl2+QhLLU9RmIN4bu1P87J8A97l
ySkKfze96MC3IqXeJUMVNeC2HPzNfobaS5Rv9MGpuCpLmxSV5VaCYJmPqCI/t4Is
XptPLizpEXh/vlJq6VvlAiyY7ssGm+ivLgGz5H03kmdtC1vCx23obwjfQoQEXSWF
XUp4aWnmiw8+bqFsdICxliqANby3Q7bMSRTGza8ynyCPXh1zxzFcmRg/BSiIRXJk
xkAGnW2LdVfhIdSmii4M+6yKeqUldT4zx+0xzaagaL9Rw/lqfj+EgwRFCeFDX/GO
OEAFu75K9EAhwq85ebORo/3de0cSh+sInn2HEu71xZEhilmGgeOntU5HrM/U3zJ+
2/G00E0SDYzPMnxZRmEMkJsTsCauJW5Z3wDfn4IRn2lQ82WIk69nqMD5Bhk6B1L6
6ycJOeL+6ZV6NvVPvzVMcFa44UmhnN6yiZtq0Umug7KiuFgHmekdxG8xUPcokocr
f0+f7pIVPyfkgngCKjZtZyjy2TW6MCz0y5k7S9JPWsOX4pXJKfZnRjf/UnP0b+Gf
6SWMrYhqXKOooaG0ABjYisJOihCRHYD/+3uxMf9jDKmmKqTpM7zmbHKIe4iBFAxi
FjBUIPzXvnXIDi2vtC82rHh7tEgcP5OmpIVy6FSki94a9MISVaZ/HuFQofOzcOvN
niqrfibJmIkNNopQW3h3WswbREv5M2QPvPtWi+UTz4aLyPBFN1qBCx+gmEtCe+fj
jXBXnIGLiGvUz0hciq9y+9aWNIY3LaSS3p0XIpxnYqdqj+HQMk66g7NDnGxnL+MJ
qdic+p7tVmCFKoW6zgLP63bSmC5um8wHAdbyG0T+guPDv9N1+VXFR3RQO6GrnVuQ
zKxkDKKB8a16JapxOkE8Ca/egLZQVSQ27FUufhmAN1u1GimDOvG/D3XEIKTPO+lT
ssMwVXPO7sX2/sZit5zmYi+KClFkZkpycQOAs9wZOZfr2gUfXUCy4VT1hCcGuXCL
fCZV1iRefZC8SruFLR7i0/Qjf6+Rbi5TzZQ2j65uz9WTRk6e+LME0mZxN+33xuhP
KIt5637vOVpbA7f+P5vQZJui5Lu/D9eZ9jwoLyp+3U29QNjOri3JHawOxYYOBFaf
Y4DVM8ZaXCk+24jPlHg04+gRONVtLJWSZ+dP73avK0uHAqkZjyglXoTGSxB+4ACe
y+qXQw0ElCOogO/lnwxPrM4/II49vDDASiQvdwx8mg9bdx3Y4mvmXRExFqwmkpnc
w9oBAJeSKnu74HpOUifB3YwSAXtTqxtMwjTZr8I7T4yyl1NR4Rm/6fDFDw+O2nl0
WBNzcdzNOqDJ9k8yUG89C+N4VF19LFALQ1znqanqZkMsF/16op9Fp2Op9G8FBVoU
O4FvRL7BIW/L+He4gBo+hdazCTBNiORoLmMpiVcSe3imUkBkOMw5SO7HkcIXi4JC
APziSY6cl+jpzgppqmhcVM1JXCOln5Oqda+YqA1kKrRFsH/vEI6Np/gYReV07jIm
JPZfVpnO7TEBJOflRjhafP8yed14GKewZS67/olNWhathZtRXihLQyw0wnGci/mS
0kzOfvkJUW4bQGHthQTXnhUQ0JTLpLgicTzOoMJgGlwUgvj/2w3qzj7DsmKxmx36
LOAYa4iYtebAwzzza4dzviSX4Dh1eKQuQ43Wwdjywy4xPQ7civy4BV+MeCZNAcGV
7orHmv5CMdRLBOJuE1sFhODh9c019OKMumY0sUTNLMMywdGFYlq53fcgrbjudLqH
mgSpTH/AlPQb1r9p4diuGd9FwfkX0Q82TzShExbaRZGW0sBQwxxm+tV9fq2NMAgh
sYj3LrvqTkO9xk+BHIf6rfxm3BK8qgIC+I79txL8n2K6j35S+8e9INfp+yjwLyzF
oKSM7G8q2SRTxfKzm5lYNTU7Ny6b0DomfgiG3LogqWHreeGPpLZtunhOh1mmWtXK
LtC4kumlBWowtPiLpDzaIhCxMKLKlWuJYdwA4yTQzozkrKpDuVXEVA/Wlnzz/5Na
FQyY541teLP78dZuWeTO7hmftgGf7E3gbOPeG9ORgn2TcYTzj/A2Hz2vr7H5jYDG
xil8SZHayRNbiDcIUoob91wSE+WWi2NCuY4g1eWCCGdnBafeJX530HR3yuINzj5D
ZakdmYQrdBEA/z0TGXeBGjfD/UBhwZczkvXXKG4NUfAu/P+hZkZZ8+rxWH2D3zlQ
X3rPTgeQna0xrApHwPau7yPNtEicy+iZiwEGt31C8e8m30/HOVXjyeOpoDLCLXbR
/Y9gXN/E0YtHoLXsa0S1LCDtg/aV3D6Mn0JSLpp3MaQDm3b1jgsgNN3ilE4K3OjX
+ZH3tXiay62OxOY9OplAiVaa6C10bA8h63+LE6v6nzUTsefceQWiQGOOVZdgtoqy
6PGeUikJCWZpn7h7Yj4Z593aZXNzDGhAqVlPx09ocWgpdN21If1HzR8RhCCXQJeZ
nhSoS532jRKn3HIuy7Szal+b2nOWVh4wKf6Sz9FwWvxaoHGFJp6/IuPQlmwcbek7
jjp4hAKjiYNWEZvgfrY7Zuryza6tM0DcqBnt8J/yJLnpJkVn2hShz5yBocOF741X
Gg5Ml9Ja0mvwDtg1ZXfvT0pgEKyN+cUZWFIB4iZRJ8DdzcoTV9pfrCfAzdE3hN85
7zrsKyaw6faMRN58w/Guy+Fau0X5zVo2cSNfG0pj5m8VBwQE8w1K/hp2ETEPh/vr
O21JFbHUUS60WUyQMAP9DnybyAGxhR64Fgyvdgo2KIxYOPKXol2/oUfDF7pAUZsM
NYYivcFZgd4/TEr+CXBqav6+QYOVTyQ1KBK6ddbaEDxQUC1O049v6MDB8Y3vqQji
fVtBFP2ZOEEBr3TrsRfZ1cIRNpYe4flVubfTJdmZwFWbvfFIRWeSfU4Ai5BCqW88
hlxSP17g9Wey2bd7UEcx1XW10tkVdWQTnp3Q1j2uwWo229YOLGXmwS8a47R/v2bV
/TUGmZrhX3rreSSMHNRp8EEx2rvCZT6ob59RdjYLWfYCWY9QqmxU+S/wcbF5mFc7
rcOQl3T1nFUjIN4Mje3NzM3sB/6QtqDrmD4wPLunMNdX1aukGZlxNNaE/dJpbRLj
lr9g7D9VAAnjPOfby5Y+8a55j17eS2H2Tm7X1SRqrNax65PV/Pa7117Znp/aOjmF
9rZbdA1/270kHyeSlA9yk+A3Z9/WDx5Lqs0Q8VwY7fmdFrAIZTLKI6TgdfFuSs8j
AJpoe38/59xUC7+6davHijcmLzx/Z/c111hHe9ESRsd99lA2un2v92S3EMYYY8yL
uGqSFosk860Xaebs36Nk4rsEPEEzO4U0dcApFwgjAcHEJTmexFpCi/IETJBttWID
Kxjre/grZwaPJTrs1R/SaCli0I3ffSfiP6K86ZkentQliQRHhZCFIGHvaVy5ORRJ
8byYOt2zN90IuHibkChsnlv9ehOkbPEuTh2QJMga8rPC5ZQFYUzNCY19ORZ7idP/
Ea60yBgnHxcV1Z5ENbRFRVzl4FvisezoAItYtk7XPPrk6OZN4CS2xbNInB1o7F9U
wYMsB1NgzoZWNeaTVL0IxzBxcYtSzuu8xJXI0zwjHjyYO5EQhsqvHf7bk6vckWKR
NTIzXyfxnS6PIIviMCWdxX95gTuBKsWaIqroQFTgPV5LNmDbXUlnepsWbj91FU4A
lQth9wqWH2lJ3AaOHzc6cwzAUkV497o7D3AHX57Q8ST9Nsx7XMwc79mPGrc2sUra
8wvdvI6byrXwm07Uj8zAOl03XMgZ7UZLIvrHhTzzluk+BKlzjjZxhBUslXlXJol3
cQl00gkzHrDJIylXqvo3k7gBCytDaorl7RRV4OCXIZyXtNWbXG618FHWVWyr3GLo
INujaov6Z3Eg50W8uXydRCPyEfsYDR88sqfNlmrDa8DtNjeIRr1sgI1HpD3Ha2L1
N89UIe3aoEBIxii2Ap1eWLkPlu8YfFXL76zmT6yw9Nye431uPzTc6gAyuQBKmbBS
vFBzvWnmMp3Sh6qXwozdHHHNxpayNc9FZuvvjRJY0tAJLoqcONVrE+PXr+b2mVgB
bIIivb67BpYOa6Kq2yJnDzsxqtfkaSvRLtx+si2/iLzjyDycwCBkMbYaHxNG5mxO
F7y0NTmRlwSv/m7Seo6vB11X6EjQVDX732MC/FpzTqDV8duTVpRZsftbTNy3ginK
4Y+pNEMwQ0jlxQxQI3mr27jM9YxwEH/7OiIG93V0HpmtaJ7axkgajYDrTSmY/CjY
nIA01aspEWkegvHUpdpbQz0zMjWv17aO9q8fyfRRazrfufQCkhDZkre5Id3h03eO
HvixNv6e3n5/gBF3ugObd3aKx0vxrNLFAKweZDtu9ksKX75k6N9tkMLNPHZvMEDo
bOrKE2XCtzzAo51SVFhnr9QycKtIbC9l7goOsZKb0eKxFuMXK3krnT5d1gHDLI46
jC4zi06WsK/gMSLozlpv5kuwDYb1gHhItM6+/5mpbCdE3epmmKa45r6ImPqSzX8I
34s8Vnesp71Kmj6zhUna2NkwGEnIEYgSJ85R8bNwAeftnS/fR+zfpQSflNXB/eTb
aIgFzyJxKq0L1GZhhaLvvYtlWcprFzkgIsvXoxSXTAD5THnAgAV2ySFNXt8i/y2n
l+PUKtsTw3xZo2KC3QI8C0A6FblPY/XRL0tEXycLhUI4jmOSJWDnU00MTztMX8Gm
ZXoMCT6daEu8ZMJapEGEJqrGmcXfAJBQzwJzoInP8U5tS54RxYd5xVs7JXQv6HxH
ZPx/7Cr2xLtuetVb9x8PRns+JLSI551F++VoaG251+ATbNBsT23GwBOYuZTiV0mB
JkB9BLuEqMLju536p3/wbUUe/pvtHdThET2iBahVTwb8XzzpPBxsGfuNC7SPvj/W
m2aGxS/oFKODeI15Eondf0BozUmi3d15qVTHbCvv7qr75yCmnRmsYrRf41sK8Lyy
J5smjkrrw4HpKLIWGedmNy5bse3a+ITEE75ELSJ5J6WW6dDcqT3EOHXg0QIb66qE
1+1EM9BPDmXvEF4B/Zv6UvjX1pY6C8pbHoPmuE5YOOrCfuNgrSbTw+qVXPAcDPor
+7f3hpY7FS62B724x9NM2kdhVykwz2LV11b0jkyXweK1Z8iVi7XYoyWOzkZzEvXO
OrTGZjWrUWqh1618sJZ4oMif4+E0zdHKOQr79LN/kFYB1k9Q1gTABncA913dCyUV
QpP8VDXY17T21f1VX48nBkRklATf2F1IRKbqbusajsd5vby9RsOZuetmC54EqUWo
0J5j5wUCRpxmeZZMTDVhg9M2g75fhzu0hYv2ve4DP0GdNJpZ3c/gfx3OhTWI/D8Q
gLuGID2NgU1sSc1TJqJ6ozrEN/pqWa6NeVo0wU/sFFC5c4RdfpkitvDYZ+LMG1mZ
mPzR3q2bpwtSbChh8qeeWC8gMR4eNV9trnQ1XGSeDpMe8nc3i027hJdrv2PoiDzz
4evrgdFRKKZqJPa6UEoWtscoqLviCJrzohAq2xH2S9z7iSaNWmYE2+TCpp9Ex4Dv
EWt7MlW/vSs1o1aYCWNbrNAsCDHtuv8ifyYI84XdkRviXph5xfIO5VLWnkjXEYDm
pG/hhe0wKrpXMVip+k3BXMYeKKagZ9dGehhtVWdtXmEd2h8ASG+IlDf/Yx8okFmB
9MLE3L8LOB7T+/YuuxeNW+Aoq0r7ov3SqP20QR0ZlYeYO81CrD6GIB2fjuaX3xMq
pFBczKXGRiOnbMWGkBADcDmeJRMWVV4C/E+33+LFkt7Kpm1Bqw2Q8/lki5MU/QT/
Rm80q1LgEdg2lTGYonUX9jnR+oAvOby6zmf5fiYrvJr1auBUetMtmWq7moHOMYgi
dVDDVAzoflmX1maZ1OARIWUt5Xf5A8bTHOB9ye+SKSJpYMpavl0eFemF0i1Qx0IV
okKOmxea6OI7tCyPzREiNiTtpQr8nimSTC4uukpMnnrAmBmv1a5wqJ1DDrc37W+e
u7XExm6xuOWkPuwmRGOCr7ijsgC1yadOgxxabx3Kr4OyK5EmW5/+kRbkpSW7bJw0
1TQRwzb9rwZeIxIT8BCxqEiNLInI+ZZDGOuMGJBNXW8ZlCGhTGFf+rAPXpNjKi/q
nBe3VYgAY5W9Z/RInvyJG0KKdnaJFibrGhOjfhlmoqW/a9PBlDQYHr6ae86L4fxi
g4oZYU6YLHDJ/vsYUAAmec83io/QFq50zkctRV51L8nGkPj5cg7h61JNpKO2uj5o
g4z8/0kG4aipvcGpfMd1Evn0a5zPqZ75NIANBChPRoQp/nqEjlpuBmhf0+/H1jx9
6BrMLE0YOffByM6ewUCJfSA/uW/8WPKzn4/SnQ+j4dX7fVd+WcC5YE27j1kW7GPW
OQspeKI19R8hVTD0SelAs2PUBv6I5xqPPem/zOEUGDnwHawdR4bXHxX6wwX4IMee
7ghb/12x3GhrUBZ9v4naWZffBwJdpH6nlwkbopjSp1OU0OTlRbTFT2Tnczfmjk8v
K6zcRRrEDaiVqshJ0AwZSK38RgXapk9Emj/3TreCBMxEUmFyCMXbl6Cn7hkMSBi9
qMxSwCRI3MiprCFlYEDaWRlAq1U7ZC30HqT7eoFAkZHfxxK4GmZ6mnMu9JTly7wA
jSgVCeApmZi0J7MtxS0RWDgFuwcy/eqq8YcuvO3xOyOMW1YwJRH5o7nCikm/V2d8
dig1Dh7/n7i2a/K7FhErEQZs1FYKD9h0WDD0qwlvr+SkrngaM2czE4WxE/dTUpac
OQZ/SS2m1fctjC1NxkL913kon1vkcJEd4pTadPe+IYe1XpJDd+9n/IKz69SoDCTv
s2tc5gqKRRYBfIwRlFJ9iLF5k0DVQ9ncrTfzT7SmGATXU66Fr79UOvl4k+TCU0PE
Vkon9LrffQ0rxsuoILGY0w+Yn6IW58TZqtIeoQyFiphon27V2Q89qhepHuhwnNts
KgIgjeZkoinxeDoWlohm2uuDv5EW0ug2PRF9fMP9tyma7DNuurl6quoUSpGePD+Y
DeFTKHJ6C92zEDXSt55DAKJHTENJli6w0AuUgh59fEm926XLqDuJB49wBhk/TgYy
pbbd21vO4nEYrjhzirn0V370BDf0ubWq7XhqczJtw/twuJTSc2vQR8qZpVcGHrJG
hUzlP6gNkbzC4gZDkg6IpXtPjZn1dzqJ0ox4IKQKd3APwHWlog2l4Brd3e0e5sXS
4lf7ydrnnDW3sL2O8BN2Dqi7JU12ChKwa+t88/HQtzVTImn91rggFKIs93OVkIIb
OQ6zCjowWaXRNcNqd6u/o7aT+f3DVVXmLhvpoMwU7OE0QbFl+pe+uCnfLPRXcIVU
bszfp2p6YEdSUXV6x7OrkW63cjTwK1+62J5AinzUJHE7+SJSYc108nObFM4Xg6xs
t4ZOd2wUM+qzP/pElVwZQuAKza0ywpkviBco996+3i8GOPKH2gNSMC6zZZOs8og/
u+5Fir2lpgH8qPJUzhjPnMlc54gz7bfwHCMKW93D7EHhDu1dUDX4Z1daeMZE5qDI
tiXxG8Yp+gt4F6xo/w0CLrmoi1rSpybLBcYjj7g/8Jk0WG3bwEo3xsYO18x//+TF
vyier7ediIXvS0m7ceffJ7X+Jqc/5qYiRVBY74l5WrmrEBWImQKaWE6INJCc3td4
oz0EheCVXngygMDFbZTpBCbVS+nSMerUTGpg6NnZxuCqZ4+x4huTD5zxMSHGSG6b
3yQoxwIFErvidicGg/k49bdwChgOvQhm0kW5wzQVul+pmcmDlyR6jzEsSOIXT2bP
k8+DP8TXI9hPbv+CsaWHRMlMQtX/k6xEL22UZSsVl8V2/Kzft9+aAlTYi2Uax9zd
HuaGtrOabERXg3XoLQrlyoOzqau9OJ78s3abzzgZCwbXBsmLk+nJ6gYFGjNk2K+P
YiW4rW7UU6wXtcPZBzDWIkyVfhCpLifLkkHFcbzyOp+Z4v1jlyqQDuIC14ToqkpK
ywb9V7aJCR0F1jBcR/ptLlCAxSBXq2ZSYrVZZnZEnYb5ZbMgquJYIbAhBurhzWFH
Sm2GemUBUWxyRY3cbkMMJQWJeN6uIJDRAdBeobZe0IBgfE7xh4CLX+javvw5LzPp
HmWuIvRXjIRTEa6dGk5bFaOO34zUpbZyd691p+mPz2gEFJdit3rW0IoIxcmYFwQ8
Mdp4Oe6duR/UmHoIoqgQ0xIkJ83uISS0Fk233PvJh6EjsRili1LkCsav0iY29Wgx
7X/vIix7nj2HsLAlgfl1okWoqDqpu6Y/1Fm0UnjFnuEcFkCgMNG+znx+Omm+gCcX
S4/1yGbcFMk/70oMIBP1ybbJzULovAmYr+VPRjYirMtOnRz0muK9eGue/yIQnEhj
YNKw8gnZq7hoedV+Atldu9XxUMCh1rUMl66htXCgQdss5ozsu2+dSmaB4atxZvnQ
vfz/v3J+RP9qBjIb39g1nVgrO1yszfl/ky3+mudHlc3sO5gt28SrY9intZX2JqLr
pN1+B9Z3iubopXP6AJ28KwLMlMhvKMCoAxq0jGl2raS3guIGHno1GYkNP3ArfLkx
dTE0LFPI21V82bl5VZw2dAqgutG+bvJsXyxiir1PhOLs2Q+SuBuDk6OQKu1qFM21
B516AVnPCt8B/quHQ8Q1TzOWmUGxNkgxhmQog809LF4tFsZ2QWH/YILUPXvLoZm3
rKWb6EoNNWZ9p/8+I5FeUo1wLyl3BfxYQcbVbx9ILUOBDeoFD9K35udAcBEvi3F+
Owm11ckRa4TZfkYhqQCRVq+7LhUez0bNnva4PXwWr3ksfGdXllb7vlL8o9Rbo3Uz
Ebwm272MI3QIsCP+Arj4J6E570PrXya0vBnSj9kd6TXybLiZDpb9KYN4buotSRoa
KrNW3yhjJpuYCHUgWRbcFqLYcF3Egi3iWC9OGocQFAUmLAh1O/P9A/GOTlwIZY2E
qUeyCj/bV6aCYUP5s5cj5L6I32JwqEI8In0CHmRQDwRSj+ep7XOkhHOzw2wNLguz
F8A9Q8/IRvUuFvCfj34ctbvORV+pOeWj4v5JaqwlrvfZbCBdbVA0uVZvibsUygto
Yulp1reAm3b2/DeEcW03RfwcP27xZN1A7TrDEXgmtMjOQ3adkfMXoKV0GtEmsRH8
IJ23UeKV13d1AgosGQI5it7NtnQlk696edvKMbsWHwJT+XygsbcLgbmYTmvI/uGG
HTtGzY5AO7TG47nec+3/otcFHg0Olp8rBGVc6EKO1BFxfRUlVrQVJbHXVoAt6qz+
q+DjR8DA8HLkbvLNfeF6b/08zcckjM1dnUH7/CVjBJ1+ihkq4ZeNVKmX3a03TTJM
MujJQqHCDuPm/+HdPULhaIZQ3UaDbo+XoYwpmEgPfYtuZiSq6N7qTiq3ocYV5gTi
V2w5e+5ccTzo37bSUyQ5ebDJHLgvkIrkGKBYyyZkIwwQjzSFGLikGHrZvIc+dmEZ
H0b/4VR2y0BgjdQqkgcP23VVpc+OmE4TlK7XV/g+BwvyKEfF454s+a/4d1RkRRQo
8EPw7cjm5VBG6GqOiFBi5VsrSNZ+s40tPCCR/AVTi8GJsWEC1hF/g3h9d2G+d1vK
FeCAWVebuOgpeoQmsnJF8dheS1jga9Lo/nfgTRt8o117kB20hPI1kp5bPrhNk5Fx
73kPammzojyxNq3kzCDpz46lndOFBDIapVgI43w9y4yL6rrA0eja77U6d0uU37Nq
BBoOWq/nvS4vueq6r3BJqxsOhV/aZUnPlCy/c/7FEerqzjKM2XYMJZi8zqeJhB+J
cOo88XVr+XlwPhmckbyV/CD5YyjzVN7hkkzvhhG0fQNxSEconFhjydXK/karvxzN
B3dFFTaqG/4MFWf7Tqfrhz82R7w5sRCyy0gjyAWldkK71UitG8DhRsflZ7Ur/+pH
w3ou/5L4sd855SIH3yoVmAj9JkVkHSMLpHXfz7bfJF17dVFywkjnCe0rsxp5SN0j
VbzNAtCEa6zD6miJnFBQZQnL3YGFoCmkz1k2XBViVeiHzb5QCApA/Sh3bncUNuBV
EJd/2N2iFVzIDoT0I+LYn7RGJTagG1lTm+O0UzPCl0h4m/cejGgRwlfFgERXhbhU
2P/5Uk9D/MiqyY8i4DoP9EoZyuUBCS+J6Un8EwGL7w5S0H1lXSorr8i7WKZY0mRj
6YtSo2i7XNAcVg+M0BNjdmljPCqy4DC/O7MGFihtCv+tJThKvnOOjmooI//vD4aU
pJ44liw2l+fAZJOrltAGs4mIbDGIdIL33YACoYjlCCqCDrajTrVCXAU/ZdcudcCh
yeusEU4uOT90wqekJsrsLzWQZrADPqFye0OS5oipcNZTYCy/KTRe7NMAKKOsw5Xj
mNoMnK3IIVDACwHwyQRZ8f886UUGt6ikrNBXy494JFyzF7SO7mKnjttfUIwxaaXf
4ynsoIDCZvEW9s/IOgfIy9y+IU+LrnGYY924dQJVGttlmM3pgY2/7ql2PU7z4Hhs
yOcjGuE5Ix2HohiO2BbCf9kld0dUvn3Vd4DR9KQDg2Q/8kfs8e8+vfsTPGS0ywrD
lBcjrNIfxUEB81fj0cP03K7rjPtwVOhNqGWMAKXG2V8PgG2sjCf6Xj74M7APk8SZ
T8/I0CCNSaCjnddcxpkiyrCDpVvhoW5yFrt1QgoU4r976ZyGKFI6LPPrT0/uBqnG
Ut6djHvzL7xOfHwZFzVmfkS3sqvg0ofSh/Sdj5zaVkYNlJ1Dxs3SvKQkR3MJhEE+
ZnnFUUc19S49yeltuwZg6V7YoeJx4L63JFNWcfEC6oAMOjIJdF3+h5A2wLX1S7Ey
2iJAtYYPmzeeT7hQetmc0WbjRuRSicZbWeAGJBn83qh/p5nQTqN811DQ3N1UN13N
Dap+WnozTcaW7Srz6MCXbSele/rsobwn8fkR9M++Tml02o/I6VLHVT6XRRZno2Uj
h6XYfpTN+cOPJSkydV6UqiE3/MqbS726z0wyNj7io33TiRADpVUM8NPau6jt3YFA
9Mdiaz8eMruIpWTKface6PtEuJDeKEJ0aD3UjUrTxMObL9XBWxlX1x2yDzIhueXQ
7C+Y1OQtZ6l5meKXdiMsADLt4PHTHDmfHxibTkN0yiMQ76desjjqM3AWzFaH/CJc
yTI7EWeegg4eBf4CkK+KEWNNIczVEpsj9FAq5mG3HgiLfkLpKDfacqkci/K+BSTC
mRng0Se7jDRYlVGouHUO8kcxdJ6hKj/CQFjnzE3Pk82QM+L2FveFKbeqO4pu6cML
4lQE3lUMaKKYZ9/NxLw6NrpzpsHLqE2s4eC4iQE0rc9a3Xi6RitXz/fs6SiCLgn1
JwkPd+X5WbzapDtjgmUrXYrWIy19M8AXf/FAFalaKdSzPaubuv/1gwKfPLEn3qmG
Luer38PoITbRqyBJLwbRjMqRHZ7Z5zuIvsIVJSm1thcl4maurFqmY9jdsLfRgprX
oovIxZ7GUtMN+5hPTxi+b2f/8ceEbHgf23crNpRJraktGqxR7FNuz74hjBk64oxx
wTZyPUVFTE0rz5RYpJ4+MsfTpaFk7Sm+Bdw803zjaowIt3nJbcPmk5qJJ/EzM/0K
bm/DI5KjGndDYsiE8ZTgciNvta9d3tProWe4Z7lUqTac7mmd0lPZagA8IHbISo8j
jKjPz1i8aQU7vUENDLDno3l8ca+6T02QxUDJUMrk+C7xi2+SJlil3AHvZxqvBpnG
Z/Wwr7BVVQOtftTgN55m4u9EUMu03gJ8iXgVFaEWVKofbifkQAvbqzMjvukrF6Ma
`protect END_PROTECTED
