`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FK+pxBBzdH7DLHjOPfHaSX7ecgpybTI5L4Rd4LVhBSrkZf8JyGGUahxTeVHBW6F3
pjBmL1aLHELGwY/tNza++y1khw7k0IDgBrdhcMDNGWZrOItk+jlfuFV7HAueN+UK
0KB9xTiVH/Al6O0LqS6CJWqDxH9mhyx3Aoc5/b1GOiFq1CnQbKFRsiCctrGezmds
a4FKRmvHwy+4GQOIAVyYPP+M1csdl6gMaF4snBkC0xvqSvYoExDKyivtDnfYqnHg
NiLgeDe9P7n5FUTfxHg9VXhVL5iT5fNrU25W87QZPfdcCPxhsXNvVyZJMoq/Ytbo
xr+yK7X5xXePmI4tCKBxFloMj/0nBF3nm38LIrYIh/siwY9+8CVpFnJDEYq/iTyj
2uM0WQOASW5hK/SC7xsgYX90/tV1jmKH4/1+n3DNNHMMrRoAaVVL8Pfc4mo62ce1
mYfy06D6is/k9hPHXVo1gl6WLsWZin48qydwy+GOQhtZSJYjRwIgxZfCu0fXQPPr
7JI9YG14qpMyoVmOiQL1KjyK3ZU+8Mrqg8Rc3wesSxn292gWthvpuf6YGRRUtfpK
XOvYD9e6vGr6yGk0mRT4Otq25ZB3Y6Gn6HRPyLWUaVT8Z+Do74xjrXU60YiCNUmG
oOH6Lni/Bg9sYSM+mkfNE1ylAzBbc6lpe0AzkFDisgTssESIaX1prBbmnTPBqML9
0R45IGR99XYVJawT69enStQme3gcPZOKp27V0xNET5WJDjx8TQH8eDnm0mjxcDO4
2JwOX5liDCj8rfoYo3np0pNj2yUYze7PXfmfyRlC4h+3hC25qHCI+doVnsNZWYfU
OSg0aZd8hU+QLAG4JrJPrLHitVdL+6YyxQb4L/d3zbpX9qz83NBD8DnyNFPH0orR
mB+rKN1fpHG0XYhVnjsYCbX9uqSzcDZdNDefdJgk9C/cEIAfKtcasxboZ/l3QSOU
fjcKrhQReuWIdHKrUhVfjjqCndqgT2vXV1di8jImEVVFTyYQXt+mM/RzCYhE3LML
IF2Ke0VmmBD2ntME7Et7yoRF8aeW+lH0bndpbo5prHDrqc6iUfX2vFub30ILgbnT
4R0oaUuHr8dbIxWlBsKeJTu2a5PM9r8Dj2uQmkaHAn/lOez8+xGOn70eiM7zXeYc
XGHdYGorZwFYFcBxdY80rWyXbKuqOysiB4LetFX4g+HPtWM1xQSzhpesuy01ecaL
E2IvPY1EK3+IEcsKvobChx81Uap25NoVFxVo61pvFK8bEzTiRsYkiGNd0iYAtpZM
RgUwI6UoMMJm2R0VUxi8hrK+apwBI7B6qecn3XF5lRSS1PiGs4dfpLXyUYklpTZ9
gagyelhSYEHBXgBhuCJ0sgMsKqEOtvsEM9F6hBoxeL8NxmpH0TquMsKvrexXi/kD
OYVelmhK81JE5nNO9hh1WyRngSDfwumVRDN6Wr25hr9UK4AbJzD8b6FNFM9+d8x8
d4SC6ZL9wzuQdoELc5simCBMsOHFeFA+bq3+SXbxnVXCNRsy8TlWM5tPMgpGV48I
AJp6Ayk5gLSU2qSR0QTElmbIv+4ApxN4/+Nu2Q61jnA8AEDH3WzRoClM70Gp/yaK
iT9tHcQD/IEs7fZj9ZiH6uOhDOWttJLybZObWpw04FeKATAakf0Cov29MqhmsTcJ
PBNo5gJEnI12PNqb6piNYpO+gymdAXR9C8vLsCxxVBDl8Ci5JY4YkZzhGawxGUQ9
GNoZM2F13ctiWE8toQ+Pyrp62DnX6+Qbl8jDmj3OUAO+ya77DjG9wJxXaDaRxA9/
nqsxcjBV9zeJTFkfq23wrfqQ/Y6oLIKiEFGvfrKYFwcvm8OvWs/i0pja9LJIBFGM
Z7Xg40P1k6K9/dqNMzzFJSX2Zy0xmUd5nvlhDGhzEC/+yHTcHy4L/R2tMZF024EA
aM6UuYOG3BtNlNVNG/q2RQSzlmSVNxU2XelRGx1mUwu1A6H4FiBrr3IWmW3GAfr2
5llexxnStE6h6se21S5g5ZPIUnVQkrCqdiW/1PBnGz943m2Ycr7CRudzYSKEdlFH
GMqi19g+UOyiNGMz6mV/w6Q7nTiP4ESPp9D0unzdE+a/a8uePXfG8S7HCqb96Z3x
jYvUgdvPzdFqmnMcpChikEqGVSRED8T0KLihsEzim4C2LpOnMTaGpwxoAxVlx6ZM
2dMx5zq01I/qiHL425al7XXEgvQG0pam/M+fVAxmFNYgfqFvWVWYLwP3eIpKOAaw
TkCShuEL9J1I8DFKOYV7j+htNIyh9ydwL3OQeo9uFGfcsYXStMqn+rnb62YPYunS
TmPIFyPo7E5HzK1Z2WpQZIFiWklEIuKVOMb5ioXnUChBcJC5ybGOBomO5AMI7DwS
IjoqN9sAtbTs/Ge3wNzFM9S/xaWTiIZ2nwNZP1YnKybKsQvx4wmfvzPLqqVqEAQI
xBgZ7xU0fY+YN+/sZ+6a0jz2KpPKUZjlS5w1oMFSn3mXGlG+MsK56FtuuL1299cC
tQ57PaaW1NrGzipVeq0SGeI0fX01dQoAH9YYxVmmzz1KpA0tJp9KhjM8jABjYqXk
sYZDhvg5mtMUwLejV3iIVXIukjfCEfZi2oW5ia2r+pxYGznlK0xAibI2kcNEwk1R
ECO7wsKLD3zPQl2zcqkKFmxpA2Yc45DsAz5mFSevRlhN39M6vTQZrvViGDTFDgsk
SXdAh77wLqVSTxA6ETTfTtxcvtw+h6/LvF5tAZlduUCwGo1Q5drxDiiDl0s1L7k5
z+YiVOKCmkUWKbfJr9jB8yYK7xCGoSqs4CwmShQHfeePa/J3LBW5oCUyBJ0mvbVB
Oa8oHjHQGQcXfovykTAcET5wkYmVgBdatoJkVGQdP36Hbv/ncmf+9klZYP5M31MI
cDyb8yK+YMLl9Gy3ihFI99oojA6enl+GJaIskgukNdGgU3E2miH9iEHnMOqWuVXs
l451cArIvn6Ug0aIwFYkRvjEV2M7pI9GKFq3btPUeYN7/Ar/yDRZFy06MAE5FDdU
8lHu/gOA5st6MbZFIi2HknZZCXmaPp816BjObKps6WKQ2xcMxO4R0sPfrJ0H7EWS
CgneulsL0oS3eGrjFCKV9GOFs7xzB7l9P0o+pPHnHWZ3ddL7cI5FRZmAFfjKQjDm
I+sM83dHrPpQxDJYVMd4wK2lGJOrbBF6Y5B0da3149jqwkkDW7BubiYeQgE6PoEF
f0Ft/K3bhk/FnYOqJ25OH0NHb28bGBZRCR4axpJ0vSykwX6My/61u+iP/8tCCfG1
+L5cLMKEaj2turNq6081X6RWVYjM1LcJZ4fsnaoMwY2iqnFQLUVhQoPVkmYUhWE9
2TS/LiskXFLndABtBqbUdl+CDyeuTboSZ7e/nW7cuhRR2nxClWhZ6U7qVft0RjHY
PGU7dkmG+wTiQiMWxLGXDKLoRjXi14NdSFtDgW5lseB47gM4Ao5seLpFkY52dwZ2
80hTRg17/YX2hT8Nf0GSjNUPgazlhRLswsB/w801873IinKNfFyPz2dwHdh9sMJE
Ice6HlI+qh17wXAuohWWx2ChoeAN83ACnJ5OYcUT2+L8ehj5wDHJXPT6jmroj2Al
xmbgvl3pHvwD0lWxoNdXGEEyElJoiMwCg8CLuZyCJ1DBdA2Qn1zVkpviUuOmMAZM
5U5eUZu1NGDUQ5hAK3nXURCTjCntPq8vsrJu4ysXugiUiD8BFO4HqK4wLaJEEX15
8gRFah0yWRa6g41kR9xJPmJJb6FyAVTytei+R6j6XEW1PBqrjOecwvVHXXky49I3
/eEzF79CspBsVZrBrjSgNJBNB6y/Fxf2RTeSUkC9NKkR27kheIlYLj9zLbncRC2C
nu2Z7xTozKfYcPPCidz8MCHUZVjSmaS1VFX5WXAC97DmSY98b6E3PUixfuaiuG2t
lDUdjPDEVnwZR0joXQN40D01k0r2DEmSPL124nL4qhHKukRUU4HGNbBsHJ4XTxgp
84xfxhNmQNminFcA4WIm8bjEfiM0xikju6UemqnUIOqyOPuIOMhDd3Itj9xY1Lfv
fYx+GZ6Dp0Z2R9dWWhaU533JD+CnZye1fjhl+e9Ms62btPtK0cEtTP2BMsbf5EZO
1wv/50UCnnD/+4+ClVT8D/KXgQLWzHaT8O8+VMBgak1kZiuxs5Qd7CL/U9UENJON
YsyNffj0dBVh6efHXP808Z/qKJcxmWsgsaoL8uGy0H6xnNLA41pYbrgxPIj9uSm3
PYzracRjKAVOiCe1Ddw4/KtZEqK3AQ0+uBWj7wxXH22nVs4TKaPa7wyg4cSh2kEo
F7NGdlSSOpcNpTDwhalRGE3rwiDZJ7/0FMWqJ3MDMjS5uOFB1C5pEJ8lirqo+PUH
eNCzGo8epfMbexCa8g69KSdRjuiG7t5Yk5vTj8UrE14qN5GXU/K4rveBIildD/DK
2EhdkpWsQnutwcs8gKm2c5NwluPhOhjzh6FAKsUnma5RN5o0Fa/BgFiIS6vztj2C
XdwjfuOERrCmDjidjuN6NE8Jf7OZ7Q2V3SIjKsNqj6FZqw9Qw0eh4r/iGd5DrrAY
pv4xIIW7t6S/HkWFo641qJ8j0k4icF0qfwkymzf7n1aAR7Y/fKOTqsKjm69lRm9P
g4iT2D2N1mBRI66TCosRxJBR6ATwWs8iQ4qA8rUzyFbN6S8+8se+yjA0CziDLGGq
uqhoUNm/Q9BkB2D6ENePI2j3uj/VlKihCUKK5/fYqYwdV/eFvmrnu33SJsqVP3b+
IVt4Ay5+nB75K7uuuImrEGhZZU2eL6LcqBxMwv4Uim7zILTw4+jq1VYi3oU/uCQR
wVBkzH5cOYlRD2Md4FhZsx4fiC9QBQcpfnDV4wV2iTpjwOYbuP0bZsQzde0qCNxV
n9n3SlqAk/lBH/QOPGEaWUoWXVVf2sHbZUzDBD/GL4/i2uyjj99z/lpV/iYFttbs
1OFKYOhEuheplNkB85B/SoRcm31WjTDFQHx1VE/IMecVNK7GQwWq/nrJFukJ72z1
v1NpA4LL+HB+6qYQU/19OCYLVnfSn2Z14ZMfSPuZC7J5r8NCn2nwkiltve1/wUZH
3z6wLPkyIrktrFquZEZQ/avP6tBMw1j6FlOW8h2DixtP+KCLIA9rSBK/yRBTeaUM
tl8oAcYNeZMEdOQmCXOiygE37J25xHAzCR1dDyUKD4eJUL0J+6QT8BYyV/i0sTyV
ub668BzMlz+5ICA/dxb+19uxuOCek5yh7Kz0bqmloX093NcuqETfvGIwpoJdzQ7K
Hhu3HivqoEEv4L21cZECaOhNEK7AddBQ9JK75eVtGgHoxytTI+iV5eH1Y92GGCCX
BXZV/yTfc8AggiLEQCW2uy+71VXvUENi5xd2JD0JUubA+gNaaqN7WMSHz6M1NSri
6Qp6bk12BZDJxy/m4sw++Y5lNeM6HUe7azpGlBHoCi7wXDsAYBgFMFdUreSPLpJQ
Y3ZBPe7Ge07tCvrntF83Ea6ewrcF9ZffcAR4JsyLLmTEMjNfdkWQkmArGEUlZTp/
4rgA5rBJbCb8Z34DaG2ADu/F3W8yyt35QF8TkFb0W4u9+686f+rB2MjMFF0VtZie
8ribpS8zyQm9Ny+zeoiGmgQa3Z5FnMXEGib6KJ/FEVkgNHWFP2fIWEKOD5vRKwws
5zyw4yh3xDFMiVykOPovCYDNf+KZkehq1nune/QdIMiiBL1ILx2h/5O702IielCj
K4E1ceZmGeaiaUMrLbXdrJLanN3dvgPb2F2oZnu5PFg85Nodae4t32NPABocftwC
9n4x4Ko+BUghpjpFdq4cPPUsZVRmfk5AfZE94DkTtHbnXkdk8x4NrzEXKa8vFQ6b
0c5sPFKyAb8h7DBD1vmwaaR8+C278MWXdd8WdEQdx+Og20ob9xUrrhEMT+HXR4GX
4IhxMW99iFy/+NPkP5HvhV2m48LXucy6Xekxj6AbPFlb02KwenQ8lmxE2eCnn3yj
CtiJYw1H4B7w8rsskkzaGkxseLv2V/+a+4ZkG20JNt3+UOloQ089YGd8UH4bYZab
0fWGEkLYf+1RYP2JX0gqaLlY1yYLBg81EjzSi2fBq7I0rJZQ4m4hsWBvXWF/QeYT
BannTKvnpM8opKEMDtpwtcqe2JoTsbqMhr0m2qebp5c2M/7VNJKhOYs3SMjvdmlK
pPYftXrf1pnjp0jJJubB/83U+wROeBpUbMmfzaF2iKuEqXwMhKOzt9XXx7xz7s/A
rkqAwA3z75AYbije+UK2uT06iQJUTVHq9+jw4IS7dJWgX283Dj7UEMwBpM/UC8AB
oodr7Fg0doza2Ugz73A1f8UbqIpQheGaFd2+A1uwjuPiCN+Mfi0DDYNppSKrtZLo
kggsWdNCUbHF0IoR4+OknqWw0vDvuMgUNYx4VrHdq4sZoR2BuPlw9gZkO1nX3Ch+
K+k7Q1UMnilyEzziA5IW2XuAuUdTpkZFQCxzcZe0LDFoq7OMpUro0q45AaZeZJuN
wyD57HqE9DypexoaC+3hFK2EmBDpNmz/peqiDhAeyIIQnZHtjC413Y+SIoSlD2Br
L8qnoFXeUJzswS70R6kc46fPxI8hLY2MO/e/Lvc+NksBDOWxmM1aElAYwGbMc7NX
m8fqvzrDQVkXC9vpar5gVX8vJMf7x6rb8lpxBIZoRtcViQ3pm87tz2n3EDLS9KtB
NXXz54JZAn5EYeAZzIM/AXKY9u4a7Nw1IdoDJmlGlq/AnKgHG762ipCFKv4mmuQt
Gv4X2xiJ/dTsuJYVrNvWSjRjgcKR+aI0ZBeunVLcJ/NJn4vcInUJ9ejsWjJtwkua
rSqEOQf6qOqeD/PWgmvVQFcA+AcmNwUNhpgnz7nlTRzVUxeXIlzZAYO7X3hUGgkl
p4T+0PRJlD79Ddmynb53i9+WRKafYdTNZFhSLBK6Qm+zseT4CAvtrZA06QV867JB
8ni5n0HVPv3gbv21HdV7UxAB5TDcvnRH01NNuwl300QhKr8gwP8m1zO1WOPtVqb6
0WisyGgatOdz6o2TM9CwVMW2g2kE6YaUYr3wFgOASmgXFOzfmmJfGu5cFlhspQdU
U/bGw0IPLJJNZ0vM+vOVnPuoDlFVAXUkdyfm+DgBvvtenzZmoWe+LW29IaNA68rM
rCbmZooIt1kYW5GTmfxFXVNkR6CTXgOlhP//pgZ1efaUvJcgPEUqlGZggYepNHr4
el83FbShv98fK3gYLgmljY+tbZtxGhxNePLd03j8IQS6L+AjLY1b8tgHZejzkPTD
nHlRnD/e94Py2tnCvcQCrl6HqCYy425if1s61dkon+H5EEufvQkhe+sln/A46XOU
KVLKKlFanT0VA7q8LRflu0N0XImBzJjhjyejz4QkIyeMhgjj83wXvRQ1Jr8h5IMw
V3X/ENlptW1Zs/hoVuPxSvRFYPzent33KJWSdK0xxV2gqVI2eGnsqjlbCTUPePNN
hiRxaCeHJDxnCjq7lRP6DREcEgpJtI/7EKzy3Lfcf5PqBFPWrZHAEhuGYC6ojHeJ
X0iTebWop5TQta3l2OwsX7CO8/xir+tbQ1+T6jMR5KYkipP3kufV9RSzTBR+pT1T
2ALGMnALCReD8PmtqN0MxIUKq/70sBMKrdvCF//nQ5rdVEPYHvGoDrdj1tOiHcz6
nBTwJuZA8EE+v9r2MF9sjgOnNfVAjftWqqpv4tSyAT2JTeBqKMsqrUU7aPv/izVd
ylhf/0qGEHHh4HcEiaLJkS+EkNj5Y8Brj+PN2axhb4+bFN1gXvT2asl8VexY2qiV
QSSBBgWXlnA/MBXG32JKY09//uA1bo1XFyNMkWmQ3/pUd16m4Xfi+wwDay0Looed
S4TrZe7XYRyprly+pWGHh+78slZ0wtYwGsrPPxANgWaIbEATt6sva86x7y52RHng
SdOdNFbn39T0S+BLngK5rVqaOEZFzlDQgKtwKOaRbZ9tdOYxGRK/wJVgG/9fo6Gj
wDiI1E13//YGzmrwdnu5l7wf7+LwHkYhbfrlSx0EnWUUmJ08lz498lJz/GpImESt
XQwrIQTAe2D/BcFtSWGCRD5ohYzeLaG8AyzL5HoFd5FBjrZWBypaRr9GiDZ2+iXz
j6xIejcZ3I8ig5bpx1zBarnP3P2yDmLdDnJM/ar2vuLT4E2fzRco0G9vZNT2epWC
QPbqPuTH1zzZKC/dB/6tKvPk4nw+H7l5s45VSfdBzFeCaGqT5/52suaWPtMdnaGm
E87/2Gvo6AW3e+d7/s6Iiyz52lRygciu+wa386s6pLJu/VkpWWRffXuEtxKoYmko
W0Tb26ROu2EqE6proQO/nRb8OKsURBtOyfcFQJQS5UGwpsZeYSztcTNacwVSz+gw
w3Gynvbtfem1Aj7qrWrOVY5CseOqZfkyJvIXnktIV+v9JVNaLF/v9t5bYBkeikC0
fAxlU9zr8t6OFvCVgEs/E8J7TTv/mxaHQMWYB9BqIMDPjD74JU2u3VzM2sv+zEAV
C37zCuoUl14SvRrnihc1hv32EBR9c7vcX0z1DiX8+tGqYk/4IF3yDIftF1yqkk2R
MUxCShrydti/zdUy6q2fBSMpEbeLs2zCGWd/wYGNXE43Mz+R0h55AlwViWuJkPtM
0M5PPqTUW3rCMQ3MMEDPLPI+mspvuRbN9gU0uuoqQSs6j3zpozaDWTc4zW2654e9
lh4Ch6PkMATLLoMoWCUtKOys+k9UCqGKZXs9lbqkGGw5KxcPBHDzjYCmfLLCsJSZ
CuxNvgn7B6eRv86KK+1lxcHLjwiuHfQpwDCpmxynaZarqLso+cqMCergfcNnKP/W
/8x6BCn1+96Xi1kyNKJwb9JpKPDXTfWg8p7/z0lrX10lHsKjmbFVOP6b1PSZN1NA
fDoCiOP079qml5kHg4eOpFXFXCww5gpT3lWtA8UfHJtRGd+CPAECoOVGEzvEMhjW
SJRVSGG8Z7bi0zo7uAegv1MvmsTpBa+MVkVyauS8qDjPeXPQRYnbb4/yZ8iozA7V
tFahYwAxc4TV4+wchvKB6gixWnFtJZCq4jljAG3r5+oHVB0p8vdYWL15nFcrOv1s
v7759nqHQEiecuXbPkSKOANVji1wsp5zgYNQhymFzH5sGG7PdZq+7UM5s7ty8FRw
PUbvMctEMV5m6zOiN2Wq8rA3h+J3j4nw/dS/CV1bgBot8AH5VsoJsmd9K2fx1vi2
vo5L/a3nMw57oYuakw/YQW7LPv1aRrR9oBzqGKR8iTdJpBc56d4Ru9TEcXu7vYG3
kHCDE31M8OdCKTs0Jgmsc1p2WIukbeaySQHdhod/EfXk3kxfWQERF6tBThni8G50
Zys8zvwINJHA0UDG1J/CXOINsB5OP3UGxC6dWZ5DSBM5llv5/DWfjyZUfLtw6a4B
EZqGmQJRlHD4prKrsBtFrd8qHZgpCOnh8Ot5ld1joOqXwbo17FyOdI9eTmClXWg1
IgNTFfkQE1fzzadNqpgYARG+VY7ItwDw/qXT6ZbkMMLP2w0F6hGn6rWluZ57/qKh
bL7preEM3sHvuFXn1oFJYxx8FAQ2Rb60IU49PVsM3NDs3S+6ZxKZDJyE7ZkLDlv1
L2VFitC81nd5u+8QG/OVrTp4QS8e92vmTXbpTJ110HNWKob2t8GZJxc4vfhU9rBx
H1CyWB6Q1SqJ30rBC5a5G8JBn6634+7KPiga8a3RPE7FD12jvWdXQwfr+vorCdOJ
3SFysWzQixlAiF4F0Ur2IL55mTe/qHpbd06GcO+hszXvxDBqikjs8HChiPwmLuMj
3vI/FpCCStzGvFZmGuk9peRwgJfqeSRQ6wKieZfnSTlczObyHjdbdBwxLKbHv/Vh
H7bkkjXHKOKB0UHMiI9LLNnuYPPDwI9XtWtxL9NzJfmJq7M9BL1zjPvj7g7E8/Aq
yCqwNferpGpfcH1wPJQqjWWLtyg/rakkmQ1+rZvbGzVzfN6mnf5qndgiMABqBiCG
FwzoETBN0f1iM51WaSm2Q9eD45Ht/O1g4TAP6mo7vYm+h6MVQAwL6OBcmSEtBCdm
JJPofXofnKAWn690RW84iEou74svwlk2hUBwsGlzPD6TRWksOyz3Y+xtuzBhLfdI
midf2IJn8PhVMjQyr92LRe88AHdZkp+zvlRmqCIwEVz5OLTaSWQBpgCBUS6173/I
RVogVxrPe76w3htJEe0T1kO7hf9eA9ASP/N9WGiVlB4zhseNstl4SKi/LiWib6hr
G7TzcCo1+OUGar2vSRjEATdtxMxqtv8ibspkXCwZLomMJxRVhZ3vBIxx6ryeY/1g
8yaO3RhEJtGn3pja8FVVMhS4EABQxi5J/yW8a0ff9TbG+D9GUl/mLqz1eEU4wgKW
u+H6oGNtVFjAFJ9C4rAesQsev+GDKsDFUj0IGMUUH+znDI0ENEG+0fEtlzJMnni1
hyWtOeXXFbSNNrWGO1Ky8fB+W7DAL5IQrAsf8ruu/3PDPJCai9LjjRrdUlOxaX0/
8kCh8ZnumVWHC6xEX8E6iHt2j6ck4wNVd6XOoT2vV/mety4z4b3fsu+Id23xacoz
E8lWxGLYdB9AzFodyeUYPrnChvh3cfDCo+bL2P6YB4LELMEQTDVZjMPnnuYcsNh8
lf0rQq2Xx40yhx0Pj0i3ijTD1lezBWKUKCQmryjbyF3rjFUnZOxf8HNDS4r0XOgs
EldzWnzBhr2T+oso3bewF07mhy9Zv0DYpeJItMHWNQBlhs6R3HTfy8c0wXLRqy3Q
yC5e96J7nxZhA2P8Jx1XGULVdvWnavBWHq2dQgq3A5z53M4w2VTcXVy2aTprSW6F
kxLcqq2XwTRFB/PTFC+2Z4idQi3Tio95z6VtGJREAAUL19wsVpBrHbQLMvbcNxYH
KOslAR7g590tfE69fU0iVNC1jjiH+jIDl2VN+piPuQBmqAP337tAvuWFBmvRhsMt
debzR7C0qMElvz2YVGJLRhLMPh7ss7wwo4rKWJpZGXhtUQ6u5GjT+7mrfmEx3hi8
nJnuSWyht8OlLwPgKjsifBi77Yq2CdRqlf8j8JkfdYAEIpDjrelUn1wEVwR9SWz5
jURaOCI90JlsKGIB/T2xNoO92BFuWzg7PQeudE4fqZA6QcyjerAa55DIvNiDYVcx
54xnbQPVWTSO9qo+nxbO283wFbJOL/ovmUdZe4YvLZPqcs8naO9EsxpwBgoYV16O
vRb9e7KnUndxP+D8sc4ClSWBTWZ9D3UkiMiSfqk1/8mbeT4n/LZqhiygZwWUGsIF
8KHCYkXdg8o3NCokTViw8GbSrwxVPZaLoZGt50jI7PCbVxu8msnUszZ0Qde2Ka7r
lmuYBlXo9ULvr4xaYeMaGmLnYg1In5IULHz3+qZOFKTqvKjZGI4Wa8blLfOEy7nX
Ml0IyPsJrYPQKgfFi2PGzIrwVpbO+4Rx0UtPL5DcDCnd+UvvhYUSvZvg3arUXYOd
qaDRf1wsKwZvTqbzU6Bgr7GT6Tp4LlLlkJvOBW+my05qwN57rY5nEVmorz1ScypP
dZri2fHrd5PDLX4U4fSlAPqE9/ufRLgDWcyg9A56HsjvJU+63k4dit9RQPv6n+9K
vlafDRJ29VxjegZVVvMXCjX9jYUOZ5VNU5gomWkLhWoelIEI1Cc9/hjJUcVytQi+
F99heOGZINy5WNszrddZV6yf7jNtYVubIDSZLWdKgSZtIwX99kWeQo2+79zDPeHt
bAsUzNwzIIqqkTqKvt62RJJc2QYMBUsXcC9LT5OX6p/ArRwGiFcdoKhITPTmMZ6x
JcrH3zDNNGRaW8p67TBAeWLzik1R7HYHWkoRYLE2mA0LNjXrFj8lQevQo1Ku2yt1
smRC7+shUarfut7tOmeFWPOy3cgFbxmoshU6Z1oTfPng/RE3GoeSeSjB+shxnhqq
s6Y930GazjdhMe7ZJelhRDba2NS4got4d5s6gxgKCTKsGqmceBfxtqOd/9nOkLdI
IoBF/2+xpIQqOjTskvPwLrfYLbhzsf3um/IZNLMjP/bQK7tCsiPXJZ7MYWQSC4Hw
DLLgOsYr/RYd6IMnExLR0Je19Fs0D4gXVPXNDCItd0NOKYxUlODQysLY2HJAjBF8
OR5ESMbvO5/B7yMVf951rmDikPsBRO+ATxAXg/GOQcDFmnFCUrTR+t6R/9E1HwV0
c2kv+zYlfawYkC8azmpkOymfU5g67Rq4cIZv5G8YhbCNVRDOX59nKqifc6E7GhWA
UrcmZTeTiuI6XWbJHhtBYsjGHwvGuNYslcCUeQqzn8eWPfsMBuL8g5G31b2txjSF
/edvAyZ8JhfRlYl4ytFavn3LdWC+tXPsYjrSb6rp3lAmw1uWH1dIm9uDO5rHler/
ZzZQsRKNPCRGzrDjbroMvi5fJWeUiqqPNkXkS3UQckj5HD5b4J1PnuLzqaEcSjTd
Qre6qhL1n6PI5AikBHisUn2fiRBw4nOa/r0/jbZGQU3rsHBWb8sRN9bNNuell3RS
1MH7bGT89cmzlFK9Li/NfTtUeRmM33FfoJzmy8c+vd4YQ1mZgFlxqAoQpmZAsgPB
bmukE6DrG+NhI28v/OGvCUMuKmo9p2gDuV3uAxWquOe/zHU257dH1LSL6GDXpGLl
M25dXMTMaSG2BN3cxUT+i4RXDpaMhls5OEWHknjgXH+H+mEaWXlYNtNMfL/SKuLO
5evEtxAi+cBXpC1Otxqerlm8B8VqqHKA/UR6zNlRvx2r8I8GZijkWDH8SgxCTRlM
7DTLH0MDzoz0rLtDgSov6V9dpcykFQ7AgISAKRvG6d+YcdDFpMWjCbFF7/WoUjlq
Y85fOPTC6TIfjDPsAKmemSKQ5EeO/jYeR6dvDgHL/75kfS+P6lejA+cR5E5GPGIM
4kEKKoOOPpJ8wU7jMJz4EFVHyqhO2MEc1JWAr/Lc3QyKVHNcaFsD7b32H5lZM8gz
9MUOMCRF1cAMrTSR2jMYe7gsAn9uTA7E0g9IJCkAV46aSNgjXstt0PaxeUdyaNWv
smQXQxOQIfjnXY6b/wJfQjoqiliWqZ5dhCEEEv+kcI7/yCNXOTG+H9kJVdInD/Ry
SOActBEneR9ozqlquGFbeHKD9/yKfGZ2p/aRlDBJHNYIRzJvKKGJw+h+5SwZgpBP
siwHcWQY5Hqq8yfVYQcLrS7O50flYMFa8EXWINAt2D9Ma3r4bKTHAEqi26BGuo9H
3VAqkWyVBBu1S2HdqRfUe3vdnLgYNzOKQHA7FkanrEQMvy8pU9ej6N44ZPfXEzDd
J972uTJXQQtqfToMyDpgyFhXpWVcFUVEfkYof694GM+jqtJQKW1iAYIrB6VPXbVK
k08BkzwplSIwmyI4GEJfZIZcZ6p0sI0IK1xc4gU6VHrNxxrBULtc7YezzzqVeDOv
mShyMC8z1WtPXkP4qdP9Q+UaYKOQq75MFmgTtwwK2Ij5oIPWKgJg75VmFaqvIzP2
1hBiYmrPPHWtqGvBZ8wzC1nYcP+rsWuidSqpbB2w3XPS1X6muyEcl0Sw4/3pIJjq
r4mGW6X1PytscI/no8r5Pudmgt56fH/oNwHK0ywefxrO1OE76QKGc7Juunr/YTaG
cu29jE7vo8fR3w9rlCl5AYlqTgrnHSIlvvmM/kB61ytIXw1Bt9l0nIYGBj77KN96
k72sg5SA32AFBXf8y5hC1VMwQClDeXACUwvgfO9tEPyi0bqdlBa+iif7krEufWD/
9aZXXqlSPVKV/2IxcJ2/pvy07aUuCeKZm4mGYGeChqZru89Jfi6UhGEnrLVVeU+D
xX+Ojqk9MfgDj+wBRF34IM4CmB+8KKx7nGPolvESoncWuAOpTvkrSA9LZrgAQVzi
/sjn0PZsATojiD6mvGLSHHJ8tZoQ/sfeHzl7EnQhBh0AZ9iPHIyBCO9H8NDYzjKk
J1fwq4epf9UzIIjzmzkRAJPDf2nh2arPPu/Gl0AACJ1skdfcOlIPBS9S4aFbxsKe
bakgwE1SXPgLOpAqXB9UCqfL2iIO5evkAT6HI2JBkwhydYepE5sh8RcJK3oW86V9
ELY8770whSEUMKeqbjgLvvubm3aaqEEobHPIL9e1rcstwkdtjDoCc5VoT22IMwx3
EQuuu+zFaqxR57dNRLOVX1gVVpAQ9OS+lvytxYyTvhG02nlVCZk40taQ+zTkOSYw
I9HDwiyuTIPgQ5zNoHwikbn23xDw/+fEktkI7IRfgvVNsY8GrHHwLfs/25HPHn4L
u4JTKHK2i4VKaVO+72CAVwntxGyM2KHdOxi8bHQJHQHLmkI/JyZ1pDo+vBtAk+Cr
ERpaMbtIk+SiFvMbAU3shz/c9WX0y32sad4b3FMm0eLgmTMx26b69DRJk+nQr8Ha
E1yhW8BwpZsdeagxfMnCWvIXkISkRGwqU9qA6E6Hy05MeiqeJPdEPhlL70NlYcvx
vxK8HrgvbChbVYvF0O+SWkvAcnHFFTCoCxGyOZAOjUJLGmA1UtakkSrYWDkPv6AL
9Drs98bjW4IGtUx6Vb5sYg5JX/coxOZ6kPd3jBYeYbtIZ8NVN7fCsy2bF2KJl1kK
HMcB3MMhgDcKIkbViNQYm9iFSYRQjZQPu4s+Q+ZpMEXTQlxIg5QxGeXGUqGGVJUk
F8KFSbD4Xs4VzjzfsWxZ8mKaIqIcjscWhwLLRRKkMNaEcz9KVfK9oFaGM7M7Cm8T
XIYx1REAz57RkMBYy0DAIbZ8/BgjHFxjlWF/Q/JyhvgChsCdRnOVjgKPqDdVf770
UzV//cIyPdHPaPZcX9TU0k7QaJU1XC4/tBJ+2xpcVuEYkztQz0BAVymrid1cRqY3
G9S2rFDtH0V8VqguIFC9zvyr3RArRPXkxUHFERK4vPh9YYp0KtNnJxq0VqUPhV+W
lwGtUUvVzaMZ0/60Tth/Dfv/+3jPo0OxLm2M7Nla7uA7TWt8tMRGLGLZoVN190i3
nPh3IemdkWM0T2BsvXsDMbre5PN5sha0UZZEowYlmVv+HVqYNWyi7WmzVzKHCRvg
jngV4x0gAGXDDlPZ0Pp7TjdIYn6k1cv2djMkPv4hy/4x0nhVGRZZqc+pfxYIkxfb
VH+EXjBkwHA7jvjzqzOuawxZC2gaYraLHnswplxk9UmHInUbVLYFnAV62G3QY+RT
lovAJyn3spSrxV9pK5GflLqbtBC/QIZD3X44jdTthFFE9i7d8CGf1YxxzA4sskjq
OuInBJcYQBH3oMUMx9ChOV2NeJJstMdaU1XiLtjyhlgOHs2eEM6oKjxuQEV3ipKP
YAnWvueUOa7v7fwOAzfB4pXzMOP+bAYmOK82VP7RPPza2b2bWGixIZZQY9isdpIj
gdGG1bA8nARCSQ3T6lA2bdw8X+KESC/9SrEuyaSiflGNH47jXQnh4k4G0ofS+w54
Ae9X84te9OMyCRH+esNOIDRb+PZu+3AcS7cFI8S1g+kext5IinI6/YS+FkvMi0D8
3ww5UuPaZaMELp6A1HF/Aap7S9YO6JTzJGSI3VjkbRet6pxlcwqlRNpnjGG+V8hA
bUsW9eH9GjTRYcKL5WJYmMTkjref0vXedLSb0nQ1g5Mz8+7pNkoHNzZlcT/fnXg4
r6M9o9dZ2ydH6WbQs8LacX96YfETgSJXsOywNx5WxmGAll00EAPDTm0QTlL16P+0
8XPDLPgnWbSU58GrzaQtC/bP5M/yk1BrdZoXBMLfqaBc5/r4H3HpVYcFhFIbSMim
z/3Gif/PhxUbFjOHb6HuULGA0bjV0YNVkgoUHKVsk2JqvK/a0xGWljsc2abj8Lw2
UvNuMRWUf0rPttskfwTGK5XRdd0BMsLE2ywzpzbFE13F0ZlNfPysy6DrjC42dsNK
BoYmUdwgItmV+2KdA3mYAiFIMOiNDozBwZ1nNgmkJvrfhy4im/gkPVexPZeQSlc7
+ZPxYa5jUGiqnRVxHM+IkBjQJd/wgpqe86CF5KS/4+faoEAXCW5Ih0Qtema9o9fY
7uwy2rQcC9TGQ4kS+F9TGWkStFhUcSEJ+QnkonYJ4brv4JB5ixJ/VK+A5CCtgIqX
2Hn9RRovBBG0hZDY0ApQTi7D4Jj6JIsf8NhwlYjb234AB+/HRs3cq575ZpwaJql7
tHWasR5Uxc1V3bxPCepOsIPp8uoGQZe8N1poznuoJmkCBdLcbnxnIO0WbGJpqKo4
845WQoaTcjcGh++R1Gncsr8QnhbB4EpcDtSE/7QTuSpwqITF/1pEp+BBIrUAigKF
9f3SbjVspnnh/ptuUn3Wzufu2HN27KNJmcp0FBUM7/3stMTRKiPYBtykK7AHG8L5
OJaXZ0UneSC7T/rd9hv773WeJv+J9LdtMJKbc5wYk6B74wGX8LTYJ2+VfRs1tPWy
Jp7eKb9uAAdTHaXH5IWHkvnyxHKnA13Q6dNFMiU+87jFVPsdNJxTSaPQBM1hj8a7
MQrPsCyp0+iwsVmBgn5RKjr396/LGQ8ZYgZnZAcyr3ZwGLEflry7w4ue8byJ/hyW
q25hsqVMzuA0maICHX7C0mLHr7DBxQkLwwryThTUm9Jcf+V8bN86HV5N/MlD4goO
AX5Kl96/fbTa2dqnOjQFyzz73DqaSJmQkRgGAbEYUkce4pZU0LqYIlalwDrG06QM
mn52j4TtXoduI6S0qOZAk7DgKkGP3D97fMDqBbh+zDg50BbHT4m/C+BD59qa61iq
vVP/toULpwZWrMFTX+fug+u+Z+PKYKjowjfTuq6ZBcNfBJe4/fv9LCSGcFWQVjP0
o09Z3NBGzPNKYJPOmn5PCwCafWfid4Y5tYKf/mNfVGd/AMsRHCgXFHH/MdyM3MCp
JdQi4zgRBF0pHtVCq0YnbE2alJdG1N9yJ20X8GUaKX147QIrO7wdRMhwuZVSNvjh
s+mnzdaayjsNG7OoaZbidQYTmBeiO1Ijlrk6REv0Pf9BoaZBnhULoBqxxtX7Jqsi
VpQ/Ekba4a7etnNK0kijQF+7Ika2N5ECQOEc4XbzU8wOf+o2VJ8fquIZjuXyjl6W
YVtI6pqikYm87JhcWBcHC1Gf93WN0fzpg6HdA56DyGSgNW7zLLdwvya9hGVtYkms
XuHVlJez/mOuhWQHS0nN3AkNmSyC0XC7rvnDKhvh0XoA9qGHkEPUOuzSWuaBdjpp
Dz5dLMm7v/4p+PPMu8R23xQgWBxW8X8G9Ix65q9BIIRvrzNoH/94QYvs8HZ7fnQI
rg3UM5zaWKvj9xM8eNF4NLpNfxExN3PuhpDBpMAI3QeOzqz+bQcHAPItV5yerpkW
O2IEtABlnX9o4O1e2jTE1I8n/LOA1R7chyF4CS04M3DjlXEKk81W/7sO/BBknnO7
tTMOWwe9MCt8IH/OxnTuOgVsWmb4U7FcthE7uZEmv4ya0mIawwmrKnFARGhqsNaj
CBIHlit7J9AdrQeKwWmiSj+ae0JnzFL0XU7zVVd4a+E95rIKoqATJUJl3GMPtkvK
A3hZNsXHoEfdIJv8jUK8idAby02AwxRe87C5FJ+LGC+y7Kw//odOMgjO41F0xLtq
eGHW/HQ5YAIuonJYNWmTZpRq8fRtvtNmdXUp0jl3ExrFtLrZ6eQDyrpGT74v4Aeu
gTcWt23bhKDt3h+6rXyJXcIhZRN3qDp4mn5F5fqqtfa94NWSbCmgwfjKhs3CfmTf
V+cxNcnuHJZx5GCBn3mvD2lUZUYmKCG+iQgINDicES+KqxlZGwd3KCAljtv9owGY
VVY5/S49Dx10lNea25CdP5MF8zgC5TQnPc/8yII/EK09x4hW/19Q2kACcyf/Xuqi
rguARoep11MjAkC55T7lVUak3Qy0u3ZRcAC4P4cRD7QOVeUh+rpso0S8nJWWl0dz
SHKdgIMXaEzJBbgo3PCGO1HBaIGbtePgCW7ar/bQ7PL+CMj0dJUFo51h4RiaZzBh
pRCuS7m4SVZePoLFGOIGQz6LsM/wwZFdcN9McLZCUkn+4JVkKqsXY/BW1kzvPpyf
LSVoPmg/FNOTAaAp+giKw2hS8y/Q0vK+shnM5j9OPPUAPIZFg5RMsQ3o5Jh+PIHJ
Cg1eqNIEV5DjJXbJIhUe7cbLlY0jhCG1lWPGs4xFQvl1xaiZA1wcEtdQl+h1qoqv
XWb+BtsE55SpbBlGZ+SMGAYY4mK/fb6XJ+MgsXOOeHMPuE8d3bftALNak4CPtvXb
aotsmaFr82f6SIAU80+26Ns64EBPB+Bb07XPIJKILS8T6Pfug3G2QW69zdAyzeib
PBRYnMGJWrCD0KCQ3TpCRpYsm7sHEsFg5r4LKVq1vGm2fFLPkHQGOe5huNqQjV8s
FQe2lyYHLZDjsvkNLSgIV/HB7rMUBTbgXHqlEg1y+erV1gdmSJPaYSBGLCzIhUau
WvvivVlsizt+1oNNmGt6CzzCWkx19H11w7t/yrULaHdkkYTqY7YqPYLktcxRKQ7h
RsUL9me+aR3E02BJNfO2fPze2t1f1BDEP1IcrBX2Sf+BI9mBGtUJHDRnvY/hV3me
DGx3H6DzZQwZ5u/gXCz5RSGZgjnYOPFmEsdAjH+PYJ16XiE0pcT/2T9AnA8Wy4xg
u2MCiklIVfc7lwYMDYh2MjezHrXANE71YVBA2zu1ndl++wiPe7mNBjEm8y3BHQOL
9ER+XvE6iED5eG9gK0toX4Nn87NDnqK082HONbn1TX7+vJdLBS1G9tf+yWCTvTxp
xBI/Ys7efaY1pJpJZmk7kG1Syf/XAgpZ0Z8OAINcqX7NBtVkiLM/zqSvncbsQO+E
SgL4+TC6NQAaHLbvHp9D+xvfCMfchS9HMxI1UxJeVFnI6mM22FT7NIJcangTWXI7
UzsGJy9iCmAh1UL3FVYqSPefmd0qtH+yF/KBqFTSsn4WQLQcizBoo//xTz5xldBr
15sZYG+2JV5ON5zljEsbGqHFT3emxvL1aNcQVZU5BH5kthncSVHz0eGLnELNF7H2
JYY1t9+qZImXOZbyQCgv8q+sbTI2JKGpPFzgnRzmrDsN4hAhKpcQHDXm09Vf0aR7
nnsYhwp+Sy8RyarFxIMvB4AfFXpgSlgvF1QIBNL0PpYMThU7PLi8Cuayr9dzM/Gs
fE18fGou8RtM5cHPxGbSPu05GlVbzGZDf+Q3KDq3ECyZRwGf8C8FltqeGI4Eyzgk
w0yYB+OQNahiy26ZUrU6HVfmPBeVi7xcKXTFGewx3/oCLJ3m2sRJHVQJ+YggH8/a
1mN4m6aui+wgal9hwd3+7lwheRrjLQ9EOB4qpB5prC4cgpAJeT6q/LN6nsM8S9O2
crGvz7+/ti1BXtzrKfmKF5vPqxgVmW1aVm/7hARj+ukPCfoAJqrcwuQeqdqNZ3MW
YucbKmFWWHeaYuapu7eCbpALup0ZD418JQ2flOLlVTYNmYdhoZh97fiAK9nQ8sc2
nTRGQfGO6VDCIFNl+v5hqmKl6HupnLKsBQm1mRjnmMnas8ABpNnO0eVbcBo5yJP+
/Mlxq2tt9YGbKYDdGlXXgKTueDXq1PWqxJDB8ULiQpCCSb36oOiXvDkTv94WBYUY
yBQ7KxlV1C9dGU7hZNvl9p3L7kfT6dzHct3AURogWpAamUemHdxAz8QPS3RfJfh6
ZdYlGiYmVo8SjyZmiUYDeqR5kS4z7DZACg6CSsSwmWnAhWQcXXRzE5JUs+ZiYLtu
ms1GAiFP0QxDfXqtU61+HAyaPjdnkTsSQ10G6Prh65QKFahK5tPt0u+WOXt7XNHc
HhAt85jR0HC/eAahKGrpquvf3vIUHcGLG2gSyzJ8wH5+irDtIMktzrVIwAQp6I/T
nBhlNPGP0xAXW3a0z6170BnHo/mUci2jkmz0w9AeYm/Lbl0CDxBgRYb+dc2kLiDY
r9XuwoHManuJLfbBZLAba/d7ikqdvCMPGEZFEt2/s/+yGQKPPCpylQ3Tp4ADK9qP
fHwDs7NBtCB0dftwTlVi3ehKILqs0K5gmnlHsZIC8Y82bCNoVK04tSU/0bqu0X6E
cDH5pDXePqDEvr0eTkbDwQ==
`protect END_PROTECTED
