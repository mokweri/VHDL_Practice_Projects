`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zNHwETpxohVK5OMQsjfvEcyRXB0scwG/dVdCWyratBqjKf+FpPlLcbYpFyVpIoPP
Y6mtgDau4PaHu7d6mVln/4hDxg8cOtDB9F0gzSHGiZi3aQLztPXwn95T58GoiCsr
or2aPVn2xnu6IyLPBML8+jbsKIWZZKtBfbkqJh25zNEBuU3r/FyOAqWiYgq86hxJ
skY3LyFuqt/p1e0NE+djPkJVBsnmb7+gb9AQgYaPnAj2aabDwwkn+5zneyjsdd23
hZfvwBv5iCxT4N8I2CloMDPlQmNL4smEXmdZkL37Ba7V2gCM73o/GSMa2sliHXGD
8LUNEe6bkXxP85MOoJSE3UR06QAptSAti5O+BWyWIjGhC9cGZxQsDYNo50xPSQVZ
m1RtYzd7htyJbpO6ENNSp38NzDkUNF8vmmXqRWP4w1cgINxmL0BBK02gycWFDrwD
yFuS2cGCMa1ACzfwuX9O/xi2nmPqieI7ZwVElkoiTrQASE7AurF6uyqLlt9EF+ha
b4OCFvb0lge8dcmaXkHO4DgdIcy+14EiIrAjN7th89cGuwebGLHw53vPibcs5zp9
LvZfCKnODk9MJx+SdXGpWT/CUYyb8C97yUR5iqd9snVmBr+BFW1dBkBjOEC15UgY
7HgHDZGd6Yh3LpEqUJwFlbHKWieSrHzymlyJVOA9U0QSKx8dCjw6p7NZBfk/uABa
1KlNe/1gd7wqqvOTxf0v/IKPkKJqNjyRF188xDOpMvrmfO55FSvk2NrNYG1yF5bD
axB3fKD+sF6BbLRIOcvkbg==
`protect END_PROTECTED
