`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yFgnnu3KANM0kqhrImeW+ac/Zx7Ng3AtPJilgRkrHk/b+uL6pR8pWN2jyZduDln3
OB1BkkZ9j/cuC+5oQDmpUwYoTSDk4H7vGmGmwreNypx2IZSOEUCpfcbTtDn4VmlC
QQm7LRuzPv9c/uCq8niYqu7JtpKqszgI6ZTPJ8IgcnzUzA00J4yeDkcBpO1Ti7iV
WEXshxTMghIRcJBZMqei5llYtFnWWfHsFP28cJs5HhwRBV993RtUmR07ifVz/RgB
WA2bFBDGeguFRtszEbk8jd2it/x+PWu8T6l4kEz/wi/sgsx8+mZ28G4AKt1Kf6lU
ryZcHZ6pu1OBXGsOYIXZtKEuzHv5tY8/F5VQ6OOuJhLH2w9l/o4Eb4H10JUzBK5l
kb9SXPwSzYhp4yyLFEyev21i1i2BSMPdP7nsChKv5PNOI0kSGbTxn/ieT7o3Essd
Gv75EIlUC0Bc8xTBM56UCg5nxFRrSV51rALoEI0Ew1QQ6e0M2Gb6BCiuF/1CI9Fd
o9v3sMFPrYiOrhguauzK3k0VSIQelLTlguskSaFUzulBryTcu6WmfSKx5ie7MMnK
2SL8q3xKdBakA/SC+Ayp6Xdo3hns7naVr2Mk8ZpjGCzPxWOftdujjDoiL0O5i0Pr
k5HT3/YGC9sxCfcslFAO229CP3OfCvy1nvC2Sqb2RuCTxWK6ldFnbRtJ9+9/RffT
32LHvWjI3+UBdDePmciKPw==
`protect END_PROTECTED
