`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8j4R1KKmg8kvhyRjQct3pfy+aR97jUfuhZtZOfm/ZYr34eW5BgnXlB3Jsx/fNY7
cGBY/X2OmqPKa5UUD/X68UHbcNIjXbulQpYh73f6WgKHOjWGFYDgpo6yK7BPqQpA
myoKth1nVRIKG3SXpicbNSVlNwKi0iYvc7Xe29Fp2z3StAZHMk9lCMtmdrrphYi3
0hW0SSVqhysxo0pWDMqNrbRmU2FkTB+hUU3bh/yIqty7rSMrCY8B+BdD2wVXlPRW
V61LPESVwmIfMDhHLHs+bZW9tDS9dkoidQQHz2kHqjJPPrvSd/iXyguquXGf+I+R
/ZrCb/WvOlpoHMvR7tWQ9/IulSQsBWyOBEs7dwFwx0jSWso8+bljWEcNjNUDxFtn
MwE9PnkebDn4A12JI/v3G2oqqVLmcQgMBNHMZHV8cAwZUa6M/94a/DiYX1eaZEKH
DyjEwODVxVhwlbQ0uetjN5cibWoq7CKUVaiDVsjmMxQ2Q3ipEDxronx82sbYKtIE
6rcUZIV+IztZP9ZW7QPkfrQAhFzV5QAk6P+bD7d9YyCGpxkEVsxv9v0sHEny8Iz6
Ku3N+uCM/+Z7BJT91BMNiXa7MEeaAyzWDpsj2UAqCDg58s0IQZn/aYa7jj6qVCB/
`protect END_PROTECTED
