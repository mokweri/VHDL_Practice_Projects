`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FOEiln4iiiHvGIos/beOkwkaXVlN8Mg3riozWsyH1bjuGyJo2tIxd40pM1f1dzoE
Fg6UC8atrpuN/+Pt9R0Tw4ooFusk3QDXjiK0K4nT9ThiK7ANWI/LXtzOqETqhe/r
uJSFv1Z+UxHCdSgVlRNH9hE4nxraQ0Rvo8kMhQqZ1wt5s5OzvoNYjp9vH/EJf++4
i5WBhgH37H+hRH0QHUENs9D6UlBIes9SX/8E7EhNycJK6LKzSpDIZ9OGeyavhKLS
qmWVeedNIKLWnSA2e1S/rMcwqhbuv6QVn3naIvdAfxbpbgh6OmGaIF+RpGGiq+ED
CfS2vJR0P576dOqyXl++pmvOCNgJL0AqYgI+T0wQT8vi6EMk26LAa5pO1fkH90ui
Z6hAKN3n36MNFwVXPB8ZTIf+P1ypM5Cm/f4LNf6+iMp2xvagEAju68s6Q1tCPpFz
Of2Rg0y5YKezLRRJGRlTTnHMF4nS7o8d4Ja3cPvDlthIGWuwltqlZArx5GtHZpsY
u5hZurTnIci3K99AeB5pkoSjRXoXqqyw1K6sJ6k5CjqUkkKCL7rva4YE7yUmmjgi
hf83bmSPtIX8V0aInwWSa3blTnMOuczMyolEvEGpxX7oBwDKm62oI4YcFpy8LJ5I
t0ptZr8i16SH0JzzkefRh1G9dFESAJo9Ue2ld2xSECCxRQZutkdDS2PROaiY63aj
Su7LYbXDYda+HYalnTfx437RFEHEhD3CM6cWGgC6WYxrfcM9+X8BislU737pb7ME
VPmuaktRGpZ7rvvytZckWN2J7c+ylezUiJZZam88I3EdQRGW6UaZGvxE7XRtje5A
ZXPjsFSJrBT+rMDqoVGfTu4ujRuasiztAc0BhPO6z0PmfZCyRUWoRcHGTJZCmX+Z
13tgzoNNoDWffqyK1TZVUPy7F1M26LbTNYS/tXB8LtxxiNcDI8MvFEigm1W4S2Sv
22TaO5r3yFKoDrMt856n99Fg2rtF3jewn5zKQieBpDo/OhfhYMkAGqRj6ONWJYVr
c3Zc2tmq8tYsqYdwH+p8R/eP3xPHaGCeeQ893WaecRo4wBc68hVinBrjr250zuk0
BWsQYsbfNwV0MhAv2EcxEQftQCtCTcUq6DhwjvYX4d0Iu44IVjIbgy40ZJuuzoIa
HxLf0kyQuuoFpJZ0VvJdPM+IyPj/tAZ6+JMFSo3w1PBRbCJGAuKFGE2Y5Tc6mN/l
qXbHHw4Qf0BEaDP4piqCkQJRKldrBMa1PJoTcCgjbMbD4J2QX2syqU9HJPxseyfU
KvOX41KRxKZOY9yAZtKOqXFy+oomNmZTa/KigNm/EEALVR4qhvOSywbJvxkRInu0
m5ReCpQpPY30oBVefakQU1wUHe2gsV4f08uyb0Si6jekA22vHnlwGEgUIJN5Na97
zZSq4+K2IzCwLPrYqLG+GBIwAIi9DM72unMRT4OV4aW6MNq1SH8x16XkifOoOqkQ
IShicDiV12/J6Tjhp5B4iGMqVtCpvFtF7MIhV5dpZj1gErjOOF7uXruN5NMhreHO
9gWx6Z3FGd/1X0G7Yxl7o1zRtHWuiwAykNbgeFM5tlPkhjagrCS1DoW6tLYg/b3b
sfouhRgMmdNSGuXXQ++b0Ck2qHQwnASCyGD0tRBX3UGuT7F7ypyNgLl4maQn/t18
/O0pnUsLG3B73PaLKGvrETwfXNNd3Ay9Y51+Gx5mxu/Nkqh43XFoQauVLcQC4gr3
M76oRQBjwZGsuOTLAeknRjdBxO1R8p1+UKacktw5/jmHsXwdKEOSNmo77T+6BQDm
MLzUUlsRzuCnIAdAxZSxhTmslTiryCXVke0PUOVJKng1tZc8kI0B2DIQrVbsqtpA
cuVgNGzyYnPRCw2z4arXNVcNSbWAPFk8xdvvpeQp6J87LBDZtteg6Hvl80b8s9Ym
uJfJX+lOeHgMvL9UnA2xXuecPgqPXn1dalhjN0APF3RjDW88n1lnE5kyh0pcxXQZ
5geXGMyNwG59b6/QJ1xorZ/Y0VqkeU2Xa/sJHLFepN2V/h955u1Bvbd6mBlzqHsZ
H3x2dQw2FBeJfljXwG84lZdgxD5Ntp1fRAXjXQJVE/jZ0cN3JHQaqICL76C5GFcq
QAxcDkLeUDW2XReYeIWAf9PQv0J3NdF68RzHy7aTMjkSflA5BNreNOkhVHj12JFv
g3nDO3v8bnhFhrVV21wxT5nQRBL73juvAO70gq/fEuh56oMr39Gd7C1HcekMXovY
lWWrk5vbgd+g71+bGIbuzMl4bObeeCOcYU2ZuZ9WruGpDDE9I+xd6Y7XUhvpSKQF
xFIgOZlvY6QLhNgsGFuGcqhZ3qZuGmXS7McKO8s+p0GxeH6J2icxQH+Kc4+UGkD/
jc2AB/Cllg561ty1LTuPq1FDBRCKTBlwdkv92Gv1KwgICNwejrCcigSpSOqqo6fB
ln5eEjbX/4VyGIDrQoNgXAoSHD4j297x+p1610Cbd2wuDNapVy4C1nV0sSKdj06D
+xrmrcCxBlSdlFzBzsj9qAPTgUwdnMKXoVxfWCurPBZCQlUNSp1kWA04fxI/az/y
7bk3kd1EenNMxHNIO6Zfu9GNn3chKwoPF1oR0PbsGfreFo7NyJ6Zb4X1YI/SHhCW
00DrnRnYCdV78PpfrdTUHLmhhgxpM9DlK3WQbGVKxHWwCMYLqWG1ylbrJ+U8U0jx
cx+LkN+5txVb8qsHHZiHo5MSIT69qCilZBHI8T4C7b35ay2uPKhpDC222Lqm0bbk
0kzy1FeDMoVGhwFGAzXPClTM7BUWtrxCysluyJz5Nv/Uv1q9vs7nuGP+ODWhFm21
klCkU++DiWJgsEv9BiFmBLsuy83fn9AUQwvrSPokAfD5YRnX3WYRTS1+9RZzFhp7
W3/lP0fD2C/5OYMibb5VB8Ad7Ktc4qDlxbcG7/q/ab6+t2/CzM2dSyVZZLdEzwXh
opvXsP9Z1Cb1cw3ST7YS0C66sWT4EvqyW6y1sN7zfPpNK7SeGSG7xUdvgP8UBI25
BNNCos17GZUvPVXAVY5Jjtt8nBtXR9IWYjXfVa+gMvrDP1v6oTqsLYWmVCH65c12
CxyK1IUhXihcyN95WD9ryJ2dD89OJAl46gOtSIVBv7itJ3FEhUxh7l4pJlJqzxl/
PVwjpRQ+K0C2e+R3+lbw8jtM1dpisopSMjtjcOjQwT+tsGqdaISuQaVqNUzWOvTG
vfNUbAukHJx9SC5l0ZLTvpgxjRcMzj/+m1BlaxTl1RwdlE5yV1fW9Vc8fFWP4JWV
vRxVm9h1Rj7RQRnTGqrste2RbdU/Nr2Z4gVvVQHUoWE=
`protect END_PROTECTED
