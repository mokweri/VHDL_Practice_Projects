`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DE3bbzBrtd4ifj4WceslY2T1J/v1400uGxLWqGgKDnqW15WUhryAY0p8rQxN3lm
DDnG0aa3eJXQwYEN1QtaYPLlHw0jt/72ZjOeg+qTTVXWlV49rYiUnyY888ft8Ngv
W+Hp/rXXyUNtUryMhk9RvTVLk9pdWo1iVTFHRc+RSnVxdkdoThM80ydgi1LfszHn
vZU/h1IuQHCw4d76No+jedV2xkcBw3raAX0t6pMRGKQKtbI4dxcWsHI45trKSWvY
Sm9qtW5YALEu6HwAMGMoyrPvuGO0BVzTvVzoBKs19pGksZ7E7rCdb7cwF5UnXkv/
tItM9hM+GfHwxgWfCOFkqbdAN27d/21/daA4yLyzA3BQd+9dxdB2pXVnmlYgTAEm
vB5ySONFFvcz0xXMlt3nVLKv01ik2Gc63BU8DjEaF7QYNUU8FZYKBFhGBxjqTMGc
Y79thvXtarqmainmPPGxKqn7WMkeyuMT+/WQSKcIrllnQAFuNiPGucEZKUnBIjeT
ibpvNwqaOPigwaV39h4KltoNlBozatNCib+RXp1Lty9GXhrRE/cYRXWLFny8aY7G
CJtQG1cG174ICqfojzJLUkdkXk8DObEmBzKy90mf/SG4nYILf2o/B/IlT3ZjLq4F
FSoAWlnGNIBPzYUoLXds1S0mtvH1jdakLhmbns/s5i5TB1T1T92VOCysVPXwkgZJ
iUKdNF9a8OavHJOMRq6lViITWcrzOboLgAstKoAjLAoMlqQs60/2iQMtges/hXbK
Olip0wA+0yO6rpooYqAoo+bQE2DzdiCga28W3oOBgKQiSulg232KvjXaexh1cBOi
GeSxp7J3WA+P/5y9nHSeIt49kAjj1ueBIPaf5vFHvZNSh8NkBQrC9KrIFb+FidzH
X47Q3HTtkukv0EKtfNiuOraSE5snbu3nCEvragmNOAQK8NPQafOD63XKR12EItdL
KaxcNhDI21hY3wyCG00VyhlA4k7+a65N5tmTxTi/Od0bKolUBErJMajoOVB9u5op
G45kcMFYF0SaxR1qQ2gGJFbtFbHeBgaCiWmEPUUvM+UjSh/WSrPQZhEnQnJa7LEl
6RRdPDLZBNyYMZM/Uj9Gh8JqB3nhiut6GrpnpmNsFfuBLo3NW+ecJX7HTjkPzkU2
UvkkkQAGpl+Yopa8rJkWj9i4ze/sCHDGbMlpa0KTqUYolwF1JE+zxIzr/nyt5RJH
YoHTHEdBsx4WxVLSO3opAodj6UqiDYrLT8iSbk+jm4eQJPwmhwyxdXyc1DCUG+CE
6V6CfGlgaxbl4wTWhFI79k/z3KjU7DZBlmVNVz9iZHHJw2/2vu/Gtek5D5z3ieLS
l0i5mk4ouNS71mh6KBi7bRhIs07uVbKXv87LiuKfhtoRzLnzOo5QOPqj63N12uM0
9nzlz24EidAbk0PI02JIToIhUDnduvUUhQlIIDZ0A1a8LyJIKnghm+udv4nQmR2U
fkZSWX/d8GjvxLTNkYnkunae+2IfHvzgSmKGsCZp93KntzYgPqizhkVL6WVuJ9wn
EDhUOFLqVwr9jtU5yQYSFqbRbVp9hyM9lGY2jzz/7C9rI74XeX3aif1tYEkWasH/
Q5d4klGeen/k6OX0J8uqPHkh4k7PI/HVQiNm8bwHCcY=
`protect END_PROTECTED
