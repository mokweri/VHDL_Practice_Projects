`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z43u4k7flpQFuqqi9V2ZPZvhGVwYsiHv2pE3r7DnARF4Ly0IJ3c6SNdrBTBvtay0
QZoVAmSFGfF63FmFTbAcipK6FZxC1ytTjfC4K1LQ+9EqC0LgXazCiAXWrhKnxgag
sCIYz8PP0sUiFxkxYZcO3n+B4Cnt4si21YHMbiIkaUihZ9zh/9Cd8WE2OMlBNJ3M
iMfukuV95ceZLdPIceXD/9QqnhjzbCu2nkZb22TvZPYbOFWxsGAtA5RrF3PRr9bl
g0KL86UZkj8WA4doaJn6BrXkCrQ/Loy6AL47tn87aNu1ViD12df0kZ535E+yMSdX
71n7Eel4Ze0oMnjrOItcwGqJZUqgWnFT69pJB/3HMJaKfj5xfG80bzW4b4FjvwLe
v3XU+9kDBRYUHBG0IU0LM28I13Cmjf9QW5odszdrt4EUjSW+/HnXUZ/vS+/R+rOH
EmtsKoUfJk0dtLOfJ+bFI37UI/bycliXRtzslQ4DlvriEymmt8jmEirKVqGP/M4M
cbOL/e63NRPGfzZUuT4/uti9cgQJZZk34GJGtHYuaV3h3MQ6cmjxHNXKFP2XeOgG
u/HsraoPggFkk/9gyXwRc4tcN3tk0YK6vQ9MduOYf9PLnmOkQqJgvPIf3Me6lXFc
t7QEI1kqOYSMGBAvQ9oFreEAj2lvkszg9H9SRM1tnUFbnnMhgXtI10OqcU/CQbpU
FQgnM+SAnWpQKoMyFj76RokvnM0O3ujSWAp473NtBHvdWxzemjEJZM+4rBa/vwBc
xk9KNf2na3Cs5beKaoG2ktu9PR1D3gFfq3NjjDJdtzaxXD6o+9pLMl3r67HXUMRD
qg9ehod5InjuxyT1JtHd7SVUGr3xT+CR/GekO61Y6Wom/ncRKATXoH5LZKGadhiw
miILcHh+bZilBd2GP5VfyoAislPmE5aHiJD9wDAsI5gjTu4Em1HRLcnvar7nBDBK
0Nuq7y+4IdoZsUzd32r1KQWGzQ3Dop74XrY6mv7ScgQKmY02H2A+mHkPjNTKP7dH
PGrzhhU6NQnXapDFEmeM2au84GRDrMOO61km4cd1AkVQ+rCR67120MNy15grQE+K
t569oKWiUgxc9zis4tT/sO9RL8CZBFzjYwyBr7UwGHM1dOzDWYlGthpb/+rKSHgG
rQ+hUdRDMpuG/+7j6FAfRISUcJWM/yvV+O/W9uUaON1FO65s6v9PJ8sfAUWk8Caa
uZwx2zjUo3gg2EAIr1rINEIb3rjHVLLAuMPw9ddz80KBUztqVJ462yY1dBPYLEwE
`protect END_PROTECTED
