`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BrYuc4a5c88QfNcAluNthKacONNbVBhBDt807MRdr3Wgl/U0FEYXIwRh9AX6nPDS
4citq3iT7+HqKV3y2yO6sw35EjFwfHZ/jH/F/dx58DXRC5kV2SGFTFAj5XL6BX1e
/RLHu8RhLyffqXbrIj0Dvh/3gO68prZ0fsNlx2zyLzO/2A3e0pN9ofNEiO/odIZU
s/LwffPjnMYwuSYvEX/Qhrbx4kXf0CQLUe9zpJCfE8E7ZnaP/7jCd4sonzG95vta
b9ixkp3tKPs+SSVupRbJZcOJoEGzxiURwEPwxQ3SlERMpKAbRezX9phlVAhBeQeX
1QW2CJl5uhrmiWZa4voa1ezJqI2burypx1EUUwWNM/ceEGlwIyC+r8sHde99V9ua
lamdjwSIOyX9TXSFGCs2C8sQ386CVP0kEGWDqNkwEYFVqueMilaQnRO27F/956lD
TkFE/Hxd+WO4uPC4dsy8+AYGwUZw4HuROF6Z3JUsZKq4KAEo35lYSgQXnePS05rk
mQzPSQ7vIOvQvRIHth/slj3yUOA77poaXurs2OfPvQfqC2yJKcavzAnPp1tXlIsX
d5YlKLixSpBM+oSA0o/wRzju/5thR+oZ2s1XWhKR2oHVtWSduTQrGv4od8lh8mDT
EmV/amk06deFfSjT3KQo9NFneoTEltYB7tibrMYFz5ciyZB03DQGPpCCVGHRaQUX
dW6TMA96nIz8DVsSHYOs+yUf6yOL7dnHGoJyZCxlCXdxtIDYCpKcSqZGk5RsoYZR
40rBurSiBfqbFGTzWovtm7hDul7xPv5JVwIlZfW4xTFllchTQj4lnlsX9FYBnogn
BYAgAuqIIRo466SI5s7UvqXLzGo1liVe9uCG8Buo9XHUllECbOLPhESyaBOd/ycJ
A9ATsdx0LjueD0Q/IzSxwRJ/D2fR+elKy6NrB3cj4CsAQpvhMUMea6o0sUvpQ93+
an/uP+e5e8/3O/ar0ks0KnjYqnMuZla/eUb9B+jFsfZV7N1ibUKch8nosOuR26Mt
AI/5YcSsOMVf39ySHoF0rtA9JXoXx/HCFLFJC9rxkq7HCSwmxYlhYheGfOq4Ia+E
8BE7vvvqjemLWFCv1uZdRbIRnd9AxGdIlRslZYtJDop5NYvu5PPEGIRFVReF4OKm
ycdXhY22HYLx2CQ39awOEJRGw9f2hO9/KlNCCIDuFHIzUA3gZCOXEW76EJVVj1mv
7yDcZHpK5VGMOnAm8wUNHM8st3L3Xh12neOZR4qfmRR6Kyz64M9VZUM/2qpu2mjU
VLWxxi2n/mWdF12Nk4Gip1xutImB5TS7KTQ7XJ/G+d3qNUpcfxZX0mgNEdtDS98H
KKEIeLz1+KHYHU2vBSc4ETsaBgRlIbDxl/NvqKQHorXXBWHGoIM46PLMA0/W70V6
JfCMbHcO/c575LenmtjwQoI9wdOySP7yHywCght7XuNIeT1xlOFZdsPzUGmcmQij
te9dDM1oiJJJPf07fS9ljFBuypvMydswr1rGl/060qNWevWxoHy6fpaVVeeaGpNV
yD9ZfWPADx8/5QF8ya2CHLlkAHMJig6cm2EiCblwgdnb29vglhDOB2YyaeNnUPUj
yhLHSuMJbwd8sIyL4s/5Gvz73zn7PX54PiQn6fCePlJqumrDX12vo7ivTIjKl1i4
IyhCFuyc5Kaf0TAHAKq/D/7hCH6gnQF932CObRR2hvRu2dvImRE7ro3JikzGkqQp
BFy0hztVYPcAQ735KXfHWbGEoCWauToQ8VKj7+Yp078UkSwdui8HZlX5G8Zk6N6v
0FSx26bxFthrqnESswTILoxjWMkZ6Jmt50DpzG4JsMN7fKFR2/FhasCgZ3KMu2hw
eBPh9ICmxSYa85kCxspoKbiio0JVPZECDbKWDGxvr4a6wnCIRhkjRumCKNypP4x6
SHBniMjdyo1t5v0Z40+14qoCLjPgYnIvDvRmL2xo5ESY1w4QqiQKqgihNb9lMyJY
9B6yi8vEbSkPTLcQ9pu0ipfeKjvxP0PKUQTV41/fwK9D97IL3ICq1UYXKuCkTAV6
vdlErCSTRUvq2LofKiZxuDC5JDbMv9GKxTKhS7u9MDbZf5xM7pe9TnrwDiHo0d5/
n3HlNDq//SoEApVRmaocUZSaGKHeWbXBz4/Bfy+6YPo0WoUe9PWR7gccaqi7DyRW
ClRoo1iJ62Ee3nyN2+36ndX4MUdfO3sS8/O/bRfa4EGaXYWPoA5lfWHMod1BhpSt
R2JfI00QtiY4lYykRYyCnyDPC9OYj4u7FEGUMHn5KDNTRuIVPQ8ZLYHeOrzWBxO6
hiJrYxW02NLIjA8ItFVUsZkLTiLxtZxS5LJBdTbC/JJQ3SkoUNHHDVZlJm52oZE+
SFxnsykRLDQoeOkH85l+BG7WpSBPCpvSgcR75FONmww=
`protect END_PROTECTED
