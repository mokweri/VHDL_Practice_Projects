`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i2IbmpdosNp27Qxuy3EhurBePkDrUHSGgbbtW80L9ZmLayEZLfrY1sCQkUGa6oVX
ZCoqAbe1e9IUEBi7CXupzIpCTaF8EBBwji5YK5KWkdKQPDdjUkt531YKEbB62yBL
8gWQDhTga3zJSFJP8Qyb6Bh9sQjJL6CXVoD4sK+tY8LBX7Kj5sbSoUYvQH7CTcwP
NfbSnHU1lMQmTRqGkb/1rjzOSh+eKvhpWuM7cggqwlzlY+hcThyb3fFnvunhD4Ds
O05pBSI92lXdxCxdYkrlw4Gd1YXwS59tIqM19PZxMvXTKjozrR0pSv5g5fRa6W/L
rr/UDw8A3rrPBsVVWYdkfk83dHjlQEwaI+5iD8mJRHoxAIJ5swcdKgknnGdCrRU8
TTJcqeVVVITndo45vKFBC51hKfr1NJ6eeLj21l1ZFbkbAS7LAubeUEROeogXhoOZ
UBVxfaP3zCMx/kL9oyfXoAE23Bp3xwnPUJbshzaxFF1ET1/OhAz1Pjy3+r4xeJK2
`protect END_PROTECTED
