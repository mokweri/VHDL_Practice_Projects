`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+imA0S1ehCkZUE515MKFQP+Bqoq7q1qPCFaUyqZ5laVxpIBeozLB6OXopXe6+y2
A7PHgvChS7uyCOgNTs1ztiFa0VdxnAoKs9JrmKq6nST0idrlMIghtnFGsuCnC2Jo
kFAcV5/xhNnAOWkOXSbtwylyh9cGiiG84O2HMuj5tK07XjnapnE0LUC3bMpQeVRP
0WgTTIponsbmBjxEysG7BmDIDzHRFmDbRqCOiE2Rk+yRUBQmjNt80qHljeCX1+BG
3cgKIv7GLlWL0yuvq42x4GR723wTYULFo6w07LJa1DYbYlJgw8JGEWgykZSQ0GcH
aOhGUX3hhLziTfOjS9zBrjlQ5D0Xk9VckxvryOpIjhGbJ0qIsLme3XR+FKDgBi8z
WU7LyfqX1Yt4gjRtGcB6d4cTHxOseIidfb+9Dk90DHb2ExSie3hmerkcLJJhknZo
t33JiCf+FrsKeo9wAWm6z8nmpaRlSbqEmc5Jr+gz0+mdR4jYEyX1GExg7olXXtKH
z2w5XhDf/4dMd2e4pDqrhxxrfsJ3kNLfPky0CY8DdoB9wEP6rQKFb36HCX1XkHRm
y8pC3PBWqmkDIYbFLGtpZaebWPUh7vPfD+4SNl7/Yj4hwuVxbLjM24D42GxYDcH8
VDWFAYM6XavMMCJm2DIs98HjyEoOdE3RsqyRgNbLad6c1j2ifj5xR1MFhl0T+EdF
ydEspJLxD+puMq5XAU3jdNNSYpAf/LSehUh7LjsgOU7MsSmwYjI9W5Mi4RyoXzji
6aodfGuYeMoBUykkf9K5OBiXQsw+VYImQ2IsUWqvA0c68MSomav1C97rT3uTre2m
b6FU24s16RUvPhs63I0eM+/izDrgdKb57nzkSdbK92Fm369scvomvwjzodblZD0J
TjiQEsIlKMtVi79FDb02hx0WvBHOwVcJpL92rH0b8J3u2LIXmI/YDr+cshjq+/xi
TV2acyjKqVmShdSiCInEzzY33VQSURw0HmwQWkQxJqf7TVrXKrqh/pkY9yE5wrEB
ItiBBFFgxva6vV00v7+onw==
`protect END_PROTECTED
