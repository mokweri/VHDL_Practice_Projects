`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8QOKEbT8tWs2W/09ahbKgx8hQlLqkAZaqzpZ0oM5l2hHF4r8iszeSFntF/aNIAe
Nut0LsEbS2dAiTERt6fA1s5+JtuIzqayUTEzxcUIfkSE6AU+2VDQWWR4F4uLcI6c
I9wVoVWqlhXq9zpPOEXnuu/772k6ReH/N0czAiyBOkMZQAuMWRxqExHqOPblj+LE
dnKy1+MWVsZw0OHs+NkjQDPuDAMJfmrLPYu2H+3CBzA9izA3jm+Vo2fNvZN1AVcn
bGuN60Aqd3WfNb4I/ApbRZBzJe/4RsoGAARPaL6BPL8M35dnySBRgr8wVNgv2JI3
3aHb99kC8J4GO98cAOg57dB1C4SrQyvkX311Il8ostS26jxwVDc/UvQg24gOAWUX
JLo2zxAj4m0cwOB5+yRi5/KLevlch/hGvbBgjoAbZussIYS00t4p0BnGkbs/Kzig
73seDxUGaEEGsctkWWfkqu4OK747+JymbctGzY8xc5xZjUG0Fndoc4k6iwfdE01M
FDO+H8xZ7wn6hmIEBCdtmCknHwtAGDNb7ZCgiQ4n+jfpoB+N6vzzmUOoCldHcp8p
7S0ihcf1MBo4qyZtRVYbdqHrvQom36I8gqxrD4i18pZAzz2dsT7OUYzKmVKjBQdx
AMI5uiy4YIJW3S4yaK9uBubJ4FAbEivDZ/WESkbrAzl+cwomC9AFJExm0AG5UcwT
cA6kgXTivSURDLrUbtbWlayXhV7WXwrtYecKOUFDZYg59EOCmZkxie0iZ+3Z1a9s
0pgVg0Ce2DeYIcieQfBiLylKpGYDAWeP3EeTt6HkpkFu27UufVHL5QmM1Ul6sCOL
k4I1nXvUE9X/XpF8dqmq9sGXCYh8dBSjw9AA9twCDO/VogL+68z7wtSjVZShmclP
J8Wlgu7YUnbvZvYaG3hIS7Sxkhgf10FzbCdf3nz3LnM0GmIx17w7M0lAyndYjIHI
AS+Brtk4i/A1R/E1l0nEJBb9UftmH8QUI9bOqN9FaprKy0rNYwJlrgpHe1H1SroZ
TzNfzWw5gW/KXnT9du8OWSM4KY0w41Z1yuwTTw4HKRRkzCfST6l84MxpYVkUE+Xl
JKhh+2T3nyP2K3BwVLrLjPfVj14tk18fz6Ga+EbLT2E=
`protect END_PROTECTED
