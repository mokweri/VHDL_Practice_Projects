`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbPC1n51ZJXBAUqy+QQ+K/efShDzmVOUuLxRRBT+2ZHcyOkB/t1Q+K/aw+bVTlNW
Fwd6hMcKFHVbW4MMQZOo06obkNtuC74TT9ANJhEImmirl5elXhSxUIFxA7gOQ5xm
siZrdf/nkRhvS9spYDkzuiiFYrJrrFy1njgQNNa5idY9tT82Ni4BGLmaX97iM6dZ
S6MtF0fK+gFgadev8ST/K+y8e/IOl1617DTeC4zEVWkFrhHkJwchQVQ13Lv2Yl9v
RZPu4qWeOQQmZeTtlC1hZa3Ok1hOiefFW+mCR7zGQrMlxM/+QjgQA6zZwv8AekBj
AjdzAk25AGVlD5w8996cpjraxNu5Sww5CFxqQj2VnJdzPZukLuz+cBL7/hhO8uP8
dUp1y+zXsE+d4lH29NswkCfi3jfTnUHMt6jJz4rI+6MaolA5jkT3JEAZs5h7flvT
eLiZffoJk6GoFXKJaTcjQC6zEERpqlfUVvb4CTeFrIWyfophsFt0dO9PPjamPeNc
abBAD9D3IGqloUoMIvN66acRCswwrjQcwqatlT8QpFFjHsincU+5vHokcK2KgvCG
TX+a8HBJw3nOUfBUUshK/ij0YzCe7DfdzDbssjUhXw6CLVujq7z+fAw6+1rj9DGm
NLLgrWUsOD1b1SETt8EusAyPf+gX/GpBP4GqldpG6eKb3VCqU3HaJFiOzPPd94Am
BNsWIiwu1UU3wFx/sRVgsxHI2aMjc+dSvWbjqirpUFFiqJSjU7S7Ygqxx8AIq1PZ
ezM9TSELgfCwfYa26Ronr9dyGkAWuQedHAUk57zimnXGqrW5IqcUOqEwadGgGClU
G0DkQeT1EBVvgSi9HuaQyTMMc+Sdjz9kbYdzB4G16Y1/F/+oPy1G2Ln2q7v/nMYo
`protect END_PROTECTED
