`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1g8pb+ev124knU+ulOT5fwVGTL0EIr8W6x0Y2dxuSBcOtGwTmoJP1mvgtRjh3EQ
4gP+pK4a9cw1Usuo+v11EZ2dpSIkNalqiJAazmysTNTyNZXT/KD7vp9QK1otDAKd
HpS70igbX8mO0xUFzekG9xtrJpmG5wH4rVr9o4C3r9EFXD8gvL1d+5tojSpdfh+2
A8NvazAdebqRtiFWuH/+ePOdk7RJZX/PyFWen6RY+ajom68ufsLY8qW0Yjn/W+FR
lTokPnQoPKsGvhI3ld9ZqnmS/RMZBzwenVK0PAPPVzrbSl22H1d2ZZoJNw39Avtb
/dP8+1Ff7Afimtcm7QgT1Bk1qejaXG6rTO3i14UTQbWgsQb4vglSsPzhEX9rcHZR
xJ/oIprifnLsR3dyRTTEImJpl8KCZUFGv4PyujPihjyeJcg9UXbItKTRCIY0aLdb
OLoJ8FGhB2gmTnX7eLOz/qtymhTJbThyXIBey1Ev0N1sgru9pbmxxUhpVvgEEhxC
PAlrStVQTxv3QcDbwGq9Yn5XIfiRMxIIwBvxgQyydguRv3/zb1fks8f74HfKKCVf
`protect END_PROTECTED
