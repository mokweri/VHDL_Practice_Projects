`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+6O77L8VoPGxMHv9j1pyTjndEKAc62sX4PJtnARvo76t7Lk1+Pn7EYa91qK7z6Sj
k3nP+YmtkcFP8S6f79DBv5WFWgAt2oRItDxqzUg/ayoNar98TcmqA8tKFFwFai31
rQsQ8ikcGv7HkzH3TaH7ld/+RloD1elVO37IE8hZ5eebzNPjl5eGQxxybmBenc9O
E90Rw2JNBtN0Y20ttgpgexRkcDDlEQhPmo+mWUTR6JvQfGvsRhCYCkkZv+gOr45+
Cl7bjFebyeuen5OzZ5NN/WbVQFHDVohladmtn/G3sLceylh0jGw1vva6TMDYWZTE
KNXGrP1YviKo1jRsEjoEnsDKSLoYOycMsiJRPpVKzZVMzYW/9g1lDPJqwAQArWir
H7hkeUpVJ3kHSmb+hWej+fU6TNUZHllbfi4DPOqI1cUfVsVOFBC90MXvImyz8RQG
7EY5zcoeO9u88TLVZWexzswtmHVXBIjAJnNd6jKE2jCwe0AadCmWunFOfZ6cg1Rw
l65bBUVu7h/BUSzdymCyAfLMocf8wM/QTJI9MNyIBEh3gMnXYRocPglJMyWqTeJh
ptkbi6jZyFs4lxztzuDKJBmAQV/Jgz1eXn5PKR9vqFQzVdNqgXbSb7WdeamPEPPt
hNuYc0+g66Whpbn7EuclTAVVxvNylRcxXWrxpi7TZDph3CmFd2w32HMFWEkhPkvw
jMnmZjsune8XYAjvH7cPtCPS1U8VqrOVe/kHrmJjT2ecBz42jKB+N4mClrNxBnLK
VU9jjFR/xfRA4ZpNEua/ZquIK0tX49RsF0EqVuQYTQOqktrwjreE7j9su6xr53If
w/zkx8KHQ10nfJj41s487oGhd50iHSxjNGfOGn/OJOnhMYXQHh9E4P4t52rNgJib
/xHpCGmB8880QI01gArGWCdPYZG0swxmQYeJT9qUd1k0lldS1s7jbd8+/IjNzMfy
2fHmI1FWDlwJo6guHVQmQ+LQpRTh0eBwascrRdcFNGzsJROO7101ZiTRmMJhCyiS
mGBUuzRx7NBysOkJmVFTr+vOwmosCVal4frSda2PbT71Ob/uQXVW4use0jN6sntJ
9rK2Be4kxC2O/7fSteLL4OM2Mkv7fhXqYkPt4D6OAAsYFP5qI0uCsy0JfY90eq/c
0UGRVQ+Kzd2ITX7ddAScO3evhr/GEprzQEEJMn5Kcu4WeSpPrjwm7JCiHTBM0jOZ
41C0GCXkUjs1f0k+nurOHYEMQqQ4TJeywVYt/LRA40sOq7M+cjcyjwHH6NcNBbiF
qaYa0Syb/VyKHxbKb+yjY04aC++pwzBdxIXG6Z53/9Fqp2ACaUTdtUu0Gc6pmVxl
mI+jbW42PpJEoC+6QK8Gw0FL0jU4Dsk4CXx0oGu1X1CEifKl0cOLvEnwHONMedpB
exz1+ZZzTGacXvVFUjYEwAQyyLQ+xpR40yWd1IkfxMXy8vECBzo2dcy8qpYOlxfl
16X/41hHD4rfkMnhlmDarRaNqrEfGKloyqugusvAM2rjzUh3VDHnlcOBSFArV7YY
GdsAwAv0ddj6jzsyO44PAsNAyI3hDy5eYoXI12mEiay0YtLTJCE+vv4DBLeeYgVS
TIXsEvMB+F6f+uqHMxmESL6HY9ekEormhvJWZUF+0UWjZvXGEDfuUFrK/ziJxwP3
c1JArMJY1FaA9+7Q2avGuEv1xlZW8Mk9FmLF+WSp53DmZFBVCpnh+HjQsWD/FdM/
1EDsgV3uYWCVvNQ+zxY1zXg3ypdBEdmtjtLBxxGhwNWu8HrXMU2UNhV9BWVgPm/t
aZGzOCJGB87RBtmmbi0II9ugdF7970iwPMbkHtOXLt3/u+rlfjzj/3ZUnTyyHGSq
LtVMQ0CUFaVOGnnLH/n1ffR688+PZFyd0aP6RDVNKRoZZc8D4PsVVbv3ORbpV4O/
NAm6FnSfmEMx/xY88cJ2RlVgjpqz9+IAbjmTzWqpt9nqDZ7Tp6zIZJheTe4bkYhb
1S0yf2K6GmWCTZKkHP7Q55/JSRaykUmjhPloj7a4TBG43RhcL4foukcTPxQtmZsw
uineyAOwpFsekcKlCEfpkrdy+jwuqJ5MdQeoLZdb4aGup6z+FOtsfFFSV/WjjL3H
6FonvFfTEoBqbbVDjgcsnGla+o1Z/HgFiAZ/iRqP6pQ6e9qo4gIqfJ7oyQqL7YOM
nK+a3Cr+jZaOvv+OvCPec+BM+bA5Az34ZjrYXt5Rhc0mCC1OMh897FrSot67O7P6
5eXXP7sPsDVqngMDFUcUEHeLVKVIiWVRIdAC1CPubrco7fed1Q5/m1g8wzlWreT8
bgVWMy9cy1kioK513+VPM0KhJ9LXTAI2BDPLBa56PztJ10S4uL8hGjqH4MAnjGNr
uTZzPwRm4LRLphmIWWbV/BClxoy+K5lp8ERVT0As9Q0kLl5lhtCtoFcuRVYIh0Wm
x1oV/CSpKQFWaPXGc5oGjorVvwoBWKlKyhE2dYpJlIPfhZsYCD2bNrnaP5LzIVNZ
m5b0CSQC7nk6ryTSPdnbxm6pagL1DdQA4kjA/B/zjDlh5Ww6X+JHU/o4E6sGpeYl
cUbCLQ9nSejQA8Z5INFkj7HkFJI2fB5Ul7airkSP/wL7vsqQRVU6jj2pNIVLlJO+
5VDS5PDBx4C3+6Ky/GkilbZmVUndpGAiKsmJLWNbQyl0HwIT9p3GCOMJm05srqgT
TjNPpfMUi6rK6B/EIWWtQO6t03+10nuLXkM9eXqDuJMOQZlw4phj1A844/FW2hYh
d/975D/xAeeMPjDNT485YH9y006yxzbrmhwq9b3uooYLXrv9jXWy9DqhXYa1IXIQ
+IhUUAxN70sYtjEn6uU46wiiW5BgKlstmwobTBspGLeDOqRp6ouQ3katSXKF9BxF
aOF2Vfw/8G9xtIheM4E2kLPlM44sHflvvRWaLkcUNKKOWk90KWc++mxJrPiCklZe
/5g1TogaXpuYllIfzs0ueD790gcubvdf1Znp34Qoeiw=
`protect END_PROTECTED
