`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EMys3gbXFI8/9qIY15W1GkYxe0vjSoM654MuFV82gtTcHCitztrnSvuwFfBfQum
hvA6ST8JzYYMu6UepEoEhFj0LaJwBpJ7BRBnbHiI+nGaYtKvsX8yEO6KpgFmjsgF
rJhMZdVYcsef+YKnQEjTou4OiKLZUuCWmpFSxgSyCPRLWlPeUsQV+9Wunz5KCLF1
ykqSkSu94q0AZJSIB57kuPoq1OLTP8F8svjx28uOcTFB314ZEcaaMBXhtBdTg9Iq
DQQ9Gy34ehc7RjGMvLm6ha3WFThIRHf3ViV2E0GEOIAzX4Xk03yIzr1/CTuzlihO
YesDt77RA068KmJCjmer4AWhB5FnB1cegpMRFsnhdIcteC97rmLz2latSlLwv6Gs
wKTJsLutUv8FpZVGmhsrtdj5rw+noKWQimoWX2A33NWJqtVybFux7Ahl9uwFUAo1
pSuYoLfhm2kI62h/SK1+zaq1mYxbZPp4REdlw1f/OTXuZQ2aHY5mEsBtp5FnJpR+
P0lomusXlHlZkUVAj7USu/x2r4lvSqQwsa8a5RWFTWfGkopGaPW3kT0DVJnABiq/
gxXDoxGISJflAcn54Y8+yxYWjAHqgL56kTeVUn4d44AVGLP9ggXpSWulByEhbs/V
Doez4c9QFAXAgyksakP22u237xZY72nfjg9bjJOfL7m1sp1xVP2FSMzu5WxnFVTV
Ke+Sh0sTZYR5TDyhtrhV6TB4MWNXdf4jHmcX+1ifi35RKoo4bMrPX1o1MkafTY+Q
zNaXYCwkLWKz/Z8uI7wklJOwH6JxOxk1NNGHm77tvW5S7w3mX6YlkdMJS9DxYTLv
+qigj0XA1Dsp0aj8UnZPNqehhhbdnyTdcvZrZ+ARPhsg7wGasyJ8UY2TIP8SNXJE
UGf66XS1/9OX8JIVbr0yB64rUqYq3ll8P4m2017WSr0fBRkdkOpec3MTl8tEd0uk
`protect END_PROTECTED
