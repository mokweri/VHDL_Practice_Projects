`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WmcG0iKZ6RDsiT1sviodcfZT/8TAEdwncPiIZeIbjasTlxbu4wxA/af2lMN2c2lK
qK4jm5OkW7fDtmQ/f/emUMRDGyRATpYqHZfFWXBLpg+zu4ZlHba9lb4OtAa+GXsg
MsodS/jFdAmuthldgY4huCNd9hYLtRfGCJ0GjAqErtyUSCVgSmiVWQB2DPqktHDk
NAo5Mj3BqY6G61jzEnMfNFzppXUgCKzsilEbrcEI8Y1gdfh5L8X8NPVA9lMnJU+s
9up0pjt2psTdABJrUiJu9m0uTuXf5wA+bPSaMYLkEDoxp6gU+usKm6BipTKRFtiV
MnAazpw4SzcNzXMwfWtzpvXLrxfRp2varh9SY9ECL/7Qu8g3mRoY9nFlgghsGG1Q
69AFkxsO2u/CyMS2oTpIeXrjzxWkFL8LmFNJBNtrt+/yODOeU8oPowFxa1vQ1//U
dFCdxo79wap+EjnH89VY2+xCabsPifH2Uh0D23EkYvuts8O6Xnbxbp13S7bZw29G
VB5LXd3LwtBp+suzDOGuoe70+TzsOVBkKRTM3PRRK5Cm6KWSy1cXnJ2PHcruqXPQ
FAcurGtyJe5OyZp7GQJuWB05/7BuV3fScGnv0ZOM7Ujv3rU9RPn9TRpxnIx4xs/r
aLGfzJznS2zyNdNt9OjEogKnODUOeqpna7YCBJWJvTyG0EIipo2g0jL6hmE7Qn4W
rEZwUaVmSORNGZ9NZjZVZAIPYjYCV2/k8UnrjMP/1SXQLOTwObqSbzwxjbeSJm/q
sc0oN2f1S0OLd+ITGh3Rc4fM49J4KCUYAKFjzWRKQzbwV0l0B4PCk0HyGpBUvnLn
`protect END_PROTECTED
