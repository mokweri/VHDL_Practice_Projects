`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1rCoz5SQeGP9DK5S7aV07ZP/NgEEuFWZJ2wXqMx74ixDuqW8kG6/QvJeHcjGaIc
BmGtYoyUsdxLiBanvABimAQerD1PgJNiwNz6jyBUc/8HjY6b8r5DEdW4zcZagwEh
MucaycNRS0cZC3ijO9gfn7VRhyzVl4RwbxPTfI39KJXwZhuTl0dYxL2vuoOwaKFV
dVCNOG/ZP43CKLVQhPnmByPg6wRJpG7WCeMdU4Qb/7g5fr9EWnqGTDyOfSFh4pvo
zcegH37VCmgZ+dZDuZhevhKjLFZ+YgD1ajBPMw9KdCshH3r/vim7UfT4kBWAMwcX
84TGQgBqa/b5uZ/WIvqL8+Els67h7UEoSkzQVZ4WXxwNHmEaP8Ss4YNoG74Ybwho
p9LdKeEZEya2q5IMEldqzjrnns3MKG8brup4fMhaknpVrnlCa+5/aO7a/EikOgzU
0qbxm7UfHPBr1usxpmXgToDS75Ru/osruwoyEwSne5lFMonXTAssIf9Qw+wyj6Ua
gBxW96CE5w98cTy4VWwYiz1I1jDGatxEEynSpXWQOq/KmiXClZo9PCSqKD4ffaQO
BDD6jM5Bw/9EsXfvphUPMFSacLx9v/3g/oSED4u8uxXWgWG5qdoevRAJ8ZNTtQEs
5tfpfddKxf7wrtyw/W0vghbEvsipp/AGloFrJofIZvv/6B9IIkW+qY33Xq56UTjl
bSZsOjGMw4WVtZFD5/XwMDeubhvFYC1Q1Zmi64xpVlW5EBBQHgO4+bU3+PvwiVjN
UwXJATgEFEnO9QVDK5GgNpZV0tlUIZlTrkbsT6Z+wPLoC4Cjx7438eW9trtVVOir
DuxdTRpdtS9TZV13YxtQ3O3uwAhKeDnsLkIEBzZVW8bpFdAprzRwWhTbOSgXPv22
jLnw48XZi4EMW9CfBYkyJc7vP0R/apEkzvnSd9EPGF3IadlGzzlHBO5Cv/jK3Cey
2cGtIudKNiXGfg4DylXnnb7XVxpY6TmPmkAKKQaL1bHdYcHQydHGfomNRmqZ66yL
GZL13jMnN9XWxu7I9gD0UoAgoXipVgSzSkPmhQ/TGDXtVAKBnhnbsVPpxwdc2v/Q
iH91hTr80/9S0gJmqs0o3QdtID45p4XN+WTRHhGjYumoxMkfvYFgkQ5jhD40QmTb
3UXf5/1R0RaxTVOzqPXYCq8YM1uClV6JSUIQaq2eqb5j1DOw9ouHVVk9H1/j8lmh
`protect END_PROTECTED
