`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SDjRCy1U1cEpRt911me/780o4e89QEqqQbQoSPDXJIEHOhH+m3oCNuH7Gd9s/4q
RktcEPuHamek/pkDHmWBJdqpFVNCcImDiF3GLvBntlhfwfSlJdF88Co/IaUq3fI2
GV2ntGzIpb0+t+uhVyO4pgfiJne01RMImfZY+Jc1rvgiVrY6mnSSgl9PvWaQUM+p
pbN1rMYOhEC9DW1aezPODMU7MGqsTTOlIyTAr2WI3ScLPpQ/wcSj4NAkalLHD6AY
TIsy+8B5WbmJnpm2wXSjPz9ZrAmCRB8xUJJEVNx6MbLbOurAc/AnQKw7m+A8lwP5
GDMQq/w1IYnEs9ivA0bz8dikg6utrd3lOHXeb2QAOoHqinkxsyegAMxuTPoSNTkw
azctZVGtgyuGEmrL1jKelUra8tfTCk1GriI4Qgs4jK+pxvGRhCC0PlQEWIW76Ayr
gao7b5GQB7px+Kw06zFkF6c7JRah+hWOvbubnPiLANynqeSxYHk1G6mfbvLs3dmz
MB7u0hd4lu3gVJ3z9TtpsD4qTR465H84tmtVzRrofsiEuXqw8iPktK4i72xx5qHO
hHp/6srYtdZAX9Im3giwheLzf8gZJYY5BN5N1GjVWheUDkoXN8WTURnR8uwny5mh
QwNRLOowwbLOZRLAOLRF7eOZ2eU3Jabbxj10FmdO3XNBPG3qQAqBGJaTqrqCZk5N
BY3B6nmVqU+KYMr8MRaBCNyiVdJwsiolac4BBSgCuzEVCnAmm12nSLc1SjUWaEJN
ewUthysdaQDJO5VTVX/6+P5pd/MiptGaubrWR43phF8Xt70opcz94i9EgA4hPAnL
cyHqdNx9Npjjyp1jVUKpZtVMvec4YSg5WEb2UoFu7mrWbjU1nl6KTHWSMGKaAQn/
B0feDqLF6amxA0d5x5qrPdn1UaHp4Azt/Nub3+GTP679OeBfWeZAU5758ri9e1/2
ksu0NEX5XYfMPX4DWe2fB+Qyd4PW9I8/ZqcjvgqGYQO9bg4wobSSFDUc6BupSN2R
YF6JHBimBQeeOStmVBohwfImYXOAJhG1p2XTdmtiZW8yp4d/SKT8GfXNF28RAklc
+cHXJ6l/OYVry1S7qrhbmn5JqAyGiG9HMoFPStHzLK/eZPdCZHqsdPxY5ZHKeU8f
9A7pOQSmVgHaJiRh0pu9SQ==
`protect END_PROTECTED
