`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A268ntrLhpxPekLo5+8HemZupmVcPWnrTrSwBSHHIoAJphBk/6vPesjMfYXR4rmL
yyIPR6M+RkxKBrKgM/QDXidgAMiNnAznJ0Pxf1/ECZpxH1+jAY3jDf/FNPG34YEs
ZokFmqc/1p3VLa4hwBqqg4NyphUTX5SKo0hgAReeyRHAsSLYjBaYeYdQQsjYnvuD
IEdrRKX8yT6PCXkdyQK4els4GEqZTnvMLrMdvSEKxXnLUN+2DGMlqx9lYC09W5fc
/GfeaxpE4wbemhlYbcl9yQxh+ZzV86Rdig51OuU9CmOFNSrLYxg1POfJozwWPjsB
nfQT1mVACZG0ZYZnytJRkZ38DQ1kmiSsfvo+6Kj6zGtB9a8qR30whuHPUi5llWLF
kVW865nMeAl+KJgDs0rgjFn7u/NTZxX8obug95LBVAKw30y77YF/DyCjTfqM1xqd
8iNHYvpXBhGMLw8ft40LNdDNGQFR2JjWkI084Z4/XtzM8zdL+Gc9KfHFRdX3bvCE
AJ1Q17iqWvyP3lWShSmJ6z5jznoSMNmb2P4nCiOHT0VWxvmIZ0lRAKjMYUQYXMKQ
Foto9it7ia/aGbhQBC2kWH/dfd5ll3YP5gMiunF3DsQfAS0jB1SW6fdYYrd5RZeh
J56ork/jT5bIUODrM3pi4KGbhhR7VpkGIIGjh8krutJEpexQ54H3Gsyg4b/o0TBT
pLH5WSBA+cxQc7OUyHy5rTvQBTCAH+8EBD7KHhXraPJoMvaw3BgzajusYpQuAmqL
LnvLIRiQjZ8qB+RnxgpgVGJLNdQqa4nCdS91/kW4tlSyc0uLtOWtYhydp/w34Q0O
6UZhSn3H7utNQjnPLTAM/w7c3E0bD1cvlGl/Lmo5ii+mQDvqovC3SLyP6msNZzFh
IwiqtbOtjib1RSuAx4iyno2DHtTavBP1o7qrJ/4yLmXbCiHLeQv2prKpV1dwfCWm
rax8oLNOAKmlrWJ9HYSQal5NTyCAqYHuA1C7p2qGuTOQsYjzOeFIC5I8aMXARDYm
aJ+oGyt7DZHUI3TYfOZBWTlMDCzISO9TgiRcsQsHPaswdQ8nyCj4lbsb5YBKiTHK
0QKzva99dRcpGb7VDm9ptpGaw3FSKJ3wzFn0LymmXF2ZMClFjfb5uYxv21bnXjAb
e9TTXuJVtK8j8uWOqIQAZ9A3R+1dPaMlNEGILHVmtByU3jz91dbAcWVFyyRo6Gld
OaJZBeLrTfmBGlB5Qm5Jn9g8CUHI2Qhi4HjmrwuxUXPPPhs29PooBWLteUuiXWhV
wdESfNiu12MX7NZdOKdvEkIpg58L9ELI5D493Vwd+IxWWT+Hb3RVDrJVtqt1dhXN
hxoTdfazUUxI7B47wn7WDFRl3Cth6EtL4/vcCNSZu/g+iNkHHFyPsOSZdMg9U2o4
moRYvD20tjjeuw98CybjcJRcxWqU3DnVAGAD71R/AvIuuVXmyGMQFlZDj3Kqa8bp
HcmIpk3qFiiFMfl+4NKUe26n7kbFQ+Ie50LMsz7zaOYo5faWPdirgE68R+62fdMA
1bQCe9EN27EUBS8SvjhPG2hgWK77uegYquhpDgikKFQmoxZpmCJFsdSJ2ILMYa3D
WaShzs6346vfK7401lfgaCLsX4XM+mdM6lnomqzESSNnqEoCrnqT9+i23k3j9dFV
RHgzHvBVzNNMlrB9EkQ7grO9jis/LVd1R8OsPyYqMn0cPuOqsxMcGc6QXN/EPDwk
ulX9P6NbZaKp0p1SMemmfKdmA6P6zdhN6rdgdUONYEz0lppcWib6u4wZt19YKKyF
erCGz9iZqeLnJimklBeIx3arkDw1SuHmDyAGsNq8oHsQ/Y5C59LZOIQ5xh2rEja3
EJ1CbZJ285u/iHGgiRgBV5PYBi88PQ/yf88BtKLmL0ZcUj2EM3VqAsJjsUNnOgdv
3CjnXyI+qfg2W1efo2vh7wVNE9KWOJQ2Gc4L3jLULPRlYGMrGdOHyYiO0+IoJuo+
YAQt4jOxxVjyZG5kGh867E0RWDf2PfDx9o0Md67CstL5E1fdg5aIfTqkG1YEA1ve
pw0XfzyZL7bPcoqBCHwRGAJ8FaEZ4gb/1ltG00DYWx7TZr53xHs1utpDpVwhg+8t
FDZB9ecPJ3VdjWF2V7R6oQcKjYdk40LAfryZeJCOmuoY4fgR945aBzHTB7lH4hPj
1yXcFFCkyni2QakcTg/yGaBo3tso1PWyCvUCs9uKL8dsjW1GUFkEd/6DRN0EpQZ3
CjduMgmFAXQKCUMQdKMAZQE3CR8ohsAEMejUqsRCthtHRIHcCofxkxndClBxc9e9
hGY+VjLG8WhEmBgIwvG+U+V/tmQ9u8YyE0nC1jYIfsh1+VIZLVjJwupvuOulsufV
NGgHl5D+XeGa1ys6csKkR+XEFPdNxJtBYcOuGCceb0I1j+x/E6MbhxlIKiYRTJxx
GXkYAay4ghyH3BEvvT+9e1CPuYt/aWQhE6HT9vKgyGfd35aEi/iaq3mO8Bogf0Fb
Bl12PVdqWTjqP1stygUqbUvfUVlNkq0nnGiSK62y7QRLYCY78hrz2WP1YU8OonNZ
HJwy8iOci/CH2TZYhT6UJTk9HRLQoyrUD0yEjMx9tsO7OVXCcbw6aV0eF1FNYLqa
8qJG1VhkDYnp9v7JlDaaiVEeIuTjbmH2yyWphsfYnvXy6XCEO2KMGGbbpwaxCcc1
2XknD68KMTPbtquLPmzN/OsbjsbkZBEVVg6IWlSVCsFBDRvn7xt/T4IQUbwh9OoA
Xc+0GIxAHVXL8lyQnfjuh3hsS1vQYL9IqfQmgP8JS2pAqMkbMRWjkRlwPR6bxLJ/
ElVAzW2tIZlBBSGasF10w7zCHlUH8Gs8q+AAlZ2onEkSTSp6INWzukV06Do5pQ81
tThVBi8QOuBeg30siHFaNjCRGZcv5KD+GwuAdVenUD2i/ic0knaX+N7KZF5tNCiU
S1f1mqqRF2KITlbMwTtQ+NkaeWoCVvLk7aDOMl8YAhgjWpqsfcFUsEfWb8ywyEV1
FynzXeErt7iEqQnS4fSksPLntRVA685vIaJZznL4t0nz5Pcy9UZdn7aN65IQ0SR0
cbvV0JqIBrt77oHge4/ielill04id1MDfqccIXKq/4+RMAZC/AlqHHdxMlQkZlTU
L/c8PZbDWsZ4ROHTRh63nh3Mzz34xOPUiV18Xwgdt152hzRpiDbcJGlPZXdKUuZV
w5xeZ6RIka7ze6IN4pFPbbO5hdO2UiaE4rbsLZIek3XFPIUu+FhlyPHGQ+xH1Rl7
mcVmxx+ESRLct1Ale8u8ywNsMu53FW2K9dE2mPmlvSLVRTxba+LPDwMrsNCeGt5U
oyFFqQwXV68zU9UwLsH1rCudFgSvDYGgvsvxGRiHhZZrYVr0OrCq7mTbxWi4OJWK
hTDa3EsDSYu77ci6VNXy9q44suv+8YQeo8gINbmlyXaJAQ3XZzkL4q/l6Wmm/ush
bm+5KRzeZH5Szond8n7velULcoTT+Cd7eSVgEwcaeZ4I+QjyxLZd88XXB2LpNJid
ghwwZrHq2lACWd9uHmoearK1JvH9R4molqWeTc19zHHs6pxWISKtWTZTj8esfphq
eNGZFRrzX5I0n/afqrboncWxjY7Gkqp37FO2e0FBkDpMvsARJFZ379yFG7MUajFU
wxixa+aoT5bI9Kw2LZvOPGdw1XEjOYHCN9LDBl19SRkwqtJDFEMw+OtMcnEkrac0
/dcZr0G9VQkRhs8HqGwLca3Ik87XXCACDbHVdrTk7Y5HOcRSr28nkhyNafYOd607
22LTTo6V4mfBixoyKxc6bX2bYXCMruwA2zNHZ1V6rhpDmU3itKbRR4+EXrY5xLGl
JVBlR/WVTpa94ZkSSCfihdHgBhOgerF67ag80G42MbAuw1ic78fTAuBMZgSgdK/p
hmrX0ai/TIVqBCPsouPGNSCyP31iakx3I2EP+wn39H/71qpPtI+zpYKohRaItHjr
ybk4Ze//L396G3r51YmgvsgRc8zWo/TIJSiJNxHRbsjQm1YhxplSO/cigZqzGyqM
ztDDmaGOUU0lEKkxaV6EcMAyT0eK+cy2lgdDxb4s+f48eHa17EATz+BnqIBXql6V
hZT2qXb8HAIWud0dwor3OTWzbyms8XJoJDU/6oId4eQLkScT4B+x//diFAIIFqrj
q8hMum/vq23NIs7Nwpn9JKeZ/Tn4zigbseLMlPF7K3rl55nD862Kc/aT4nt9ZHGD
ggN5reKeW7k8rvK95tHCgOsAnjTG89Aeew4O2ORL+OnJXzN0iMQKrxd8SHIE7m6c
SA7S21a4TC5E4/57LrqO1S8AeN0sUzTOka4yFmLB+NZ1RYwnjaCVIjdX+N0oaefM
xeoQm6vNo+tg3GUf89TnOWKOKALyAiUWjuGJ6CtPDYA5DAbzyU+mprKac/lc3g0/
gCExV2266IGKt4D4P/qxSqD97gy+MeIxmpnVe88dcWE4UBE10cK+O3egQdManlva
61GPnA/LJj5WPwCeQFPam1ZSVsMOzJiqmZa2e5+FB+m2uhb9uHql2iHDoVgChmDQ
pHLHIiOk+Q7S7jrJ7LO0D8DSal0GG0pO8l3mOj6lz9vK5JgHVKFyHtulrqRLULHD
gjim4GjIPoHRbbRztIkAWZSxJbkUICXGc99gBZltd9G2V0M51QN+2J21AGQ7J6sH
ffRG4V64hvX9LuPlWPdbJR8B0VXDYQhiMxr47lesuq0suwcc1ruSsNEap1z5xD0K
FVTgSr4L2y2TlV/M/yoJMjg6rGyDN9F7Ix0RD0FdW9MHEC9cOOtLNRG10YYvMFYd
U0kOFxyAkaUhj3P2tgsislpQrka0LbHEZbQN5ln2yK5Vnys/gdOhGMJZgRhpuuEt
1PfjAOwfXEDTJUvV9Q1q10cDw5dwFMIqegi9EAjwaBxxHZ3R1ku4fcMDPf5b74YW
+Ghzv2VU/mYoQEALXkViEXPCRAqo/pfPyxgOxcu9DT1an/aDpkBxsUISfNFz/ybG
6brYrw3Do8+D5zlP12Eg3p6zd7aKvRK87Xz3UzDMFxS+XWLkpOgTWwrbttFZF6Z1
f5v7040HIz1uxeEZ09Mh1R3UlaEusn8w1n04pMEVKeoCGrT8/TUKeEKAfqcWtGf7
GYUf4tKpVgUlSFVNg/TEBYcT4e5I9RTD2VAUGYj10sKspH/KO8KymY4XpRzISYx9
4an7BLibyrCBu7eNvQ6KA9pUI5EkrEghhKGxc43t2TU1oZZV9NiM/OMDvjzGUayb
R0A73c7G1UpaWKiB4FRYicZijQ1edzE6wBqEoPDy3nBG2dq8yOTmyumyerxbjmLY
KJvvRC5YnkioDsBxIV5trJMpZaMhBqUpPnIshdeNdIV+Vmf8JJhmuPNVezy8HSOE
p16kFt2sG6SgFKoC0CvXeI9d7HdosmOe9ZdkzONACnr5zuGX1OLxwX4MbYXaotnR
V5j0ShKes8UhpIgt55kgiljRO0WAbrTuAVN5/p9uuRwYbZTKuJmu91GFRtz/FDDc
33Eirl0738s7TVkMPVVLNYhT+FQTzMEYT3bQoxjobq+xpxvg3S2q2Ee7RDf8P/Iq
eGDuEwXSa0Fz9d1Mwp2QzVrnxLYYGmHO8mTHMIea1DnvxJ55k/uYGdkTJxoEpquE
+ZLs5Iw3Xi4ldQY78GfYOuQu8wc+KX60bNLHpZAtONGi1vrhXw2u0FCEwJXZ3D+a
pmV44QbNIDOfSXogWrSJ7KCutSekWHigTcaevmbK7evGPLyZPZf4cTsjBN/nHu5n
ctvnJ4Sf5FQ5mMevyGkJpN5M3LyI1zflWWeh10/kKzUo+eGREpU5oUs5SJstpDoB
R6lYaIlmjqCU9o3tEsBg9wCRqMWr/vcOZSiwLaMIrAaMrA/kGkzlP00L+Str8HlV
TjxQN9ScGdiXwucKdxXz9UphHn7O8PzTdpibqB1GkqIOAdOd89s1vkXGKi0uH6fy
4ElHVbreJvRBZRPkBBQzxsBwaCArt0KsNEf0vatP57M2P2kfXEiCaeQnRKkScGWX
vUiFQc61bu4PoSMF5HckwBKmjxWO0zXBJciyMK58PU4YKWVcqHzPdytjzpPYBjsr
gWp+5C2IldIYDLMQOx4Ijh8x4u8QlYRgLvZIqTq4SBc9UCrG3X3DHAZrPQNxwcEm
P6tngPvt+qmM0seZqIP64+d5oa8O7+ri1bRb925VvHrd3a8X9BKdXADDXIFL6rXw
JlShGra1TiFwtD+HEYrpDs1pDs2Gub4Yua4j3G9YXGxTL0MCEGw+rrqF/cgRNrxn
VxyBQOj7DmfPcsdzqqpQ5gzew2HmIR+7AO3D1/CeEt8hbC+6r8URCpYoKoTQcvVa
o3EcgYOvdeDSwVm+L+IkDr83nbO/ItF0TwlqozpL1l5+HhgSveu32V60LJz6s7to
LDm3SDU33w0ljVGUYpXcUIhiUBJilY9+Pot60yx3zWb8AVmXfq1BXtqH6xaesovl
41Apl6erpaU4YNQEx7jzwwU60+5Y45n1A2gSB6tVyESoRJTVwKXPSSnPqSGY649W
C3wEQUACi6Mz66JEGpHMmM++yfavJKsoaq4zMNfrxW8Xs8IBmO6yOkVxgsax6PJh
7TB4ReD+Q5ZmL9GYugcoaKfjm6N/pNXnzzXlLRLYmxpDUOrHAB9Y9+XgKABYni6J
u5Wi/hti4dvKRMM877e6W+kKFWVcWaOv25gX5HH+JHYexEoxdvlCMl7vcnQ7eTkv
/SJUCiuHuuF5ZANb8b5XWcBdqbdkE1wE1SH4yDrMnDtc7YHM9p5Epgtayxvk9MpN
fpIvCWRsIXfk5NsQm69NGktj5iB6fDDta5om/shSBqZGD6uPjU3nHYlYZyDD4G00
8pNwoXwGkRIyNq+CV8pQKZS/ZeMOE1u4bk013Fmv0gfNS0Szl0vu+aY+zqu2HI4N
vn+1KWyvCDIccD7vtcF97rkBSMD0/5vd+YvOuiAkykQXQd60owBp+iUBQ5UAImuF
SzgyvHEIxHlEkkvPnEspaIp7Ado+ovbEtChUCNpV/0tikHd2zU+Gmr/1FeLSTNT9
2SiIoz0X6po1yNQ88MEiB5NAoK4nP6Q0JOkKaLg+b9AHoLVxXydlw+Wb+/421Lil
n3XqC9vfjXxt77FB6LkCenL4aIN0sFKy8XSmfewb0Ub0A3WJdF2JMmIF41r/VPbb
3moT+np0OXqYm15gcxPOVZ3ZBs9ML0cGMNuomPZvtpn8sozrj4wuV3WkWTXJtWLX
oHqf9lBDkdSHRhAVWJS9XXSqGYzfBUPs5QIJrFMI4P5f1XUqkQJfqlf8473dZWyk
CcAT1/c8zN+dju+Z8SnyNNxD9UKeJjRIv9HiyGL6PJYDLk695byU9epH1H5zr1Ks
mA6CuaLv7qMySceg4EGbPrcByqhm3CTHhyxWze6AqsIuILQiopibWjrb7zj2/SFa
/9aHyMBigytZdXqYrWUm068BBXaG327OatIpN1KJ/Yrf/8m7OaUHmy/W1lMBf9Ve
/K2mbSTQK0qxvYMMRISnYzaJQTocE4x75PsduD+vWTiVRHeSIsgupfpH6U/3hNYR
BrXcI9PIP/xvfD1up+5RatP5vvjTKo4w6RMzG99ZlECSLux4vEhHanjIKoEwc3Kw
O4oHUD3WtylvjFT2HYTO3apU1MXbfafGm/kpYg9cyIrgFsmbf2jAkKYl/WGqYhhQ
LsDced0qWZ0i8idyqM3eA2phkX8WXSV9IzQXcvzSHSjOdiB3EYAoLiTTkBIG5BPe
ESuVTB65yvIUg509Hu4DCYWdWhAWxRE7ah+1Q4ru6Xw2bGm2Jjl65jd+h227bBA3
5ew+/zra2m7+UdpdMRJAxbDliimBgHnNLTKrNaTBdFO+b1CqeRtgYBtOTswPtNIh
WVytG6IoYPNud/pWV5Z/yEuu3HhCiwb7VWX858fCcPQfwTL+z1I62smyhjbRJsRa
qo6ghHi2HDRZtTPT0hyEVvATKcO4g1KFBQQ+CTIUMR40j3Hrj+aClgFi3MVZOApy
0ctRXhutk3jTHdSYidSDZqkHLUTMUGxegys9ugR+4XAjargi/iFRhe+5ZhbwdfWm
N9TvxfgkotOt0PdJPazfyMAg6YoqZNMGI4k2IZTs9Xe9ex0honFTXMgeeBjmIHBd
I2iDP54mj9s8tIz6KaZYBKaDV5mbiKRDy+hhiCui4MLcrrJz+xIo+SiXPXKxqFc8
xdTfJJOkR1iL3ZHHAtJy99q+EwvKCq0JKK2CTr2D3YKH4fO+8Cv6ylEv64v0Nk1K
bTjNqrgHaGhzHe1wL+TzidL6Ue814TE3+CY6X7BbNM0mB420T0Pyh2Luhyi+mt/M
8ZhgX5tb5jzU4lp2UmkcbtARnwdVfQpHrK8M0AWPMEGNsUumFiX5nsSU4aT2fxf2
J8JuXxyi3e4FSLycDx6YBmQTqMOehNN3paTKrUKI/RRMhBXFGm3mCUbD/4lmO/mM
rysXN2htE/u6f3j8xfA6qViFSevBhW8tjmSjco1Wq8KCo1l95YOj9Y9x3rbKNdt/
bLBc/s/ff8T3ipk9bmE2eMEADcDbCCq45Bsk8oYEHk7R0u1iS+26CY7jno8B8Bnt
yJrhQSBiWaxKFUzjSmwpV/iqau59WupqUoX44oygBEUjub8DHIIjtbEYzLkXQf+q
WvR9K8T0Wp+wPQ2361PqeH84JACjwZwCMNogSK1vOaMcw2BhUPZdnOOA5rXz9kvo
s6S7TKaYdIvPwRm5xyXeTLi6tL5xiP4qm8duqZLuc/9eRgl7AhroXZ6blSTqQKQX
yLASzGp/uLnm/2B67xZ3VtYUwrXOzM9yty9/WFIbzEtEkcaO5xB2slrhThjEDHF6
ajW1IiofBNI5Bv6Ob3SDBPH5NKeKtljGcjjAqbgIImfCIG90xTv0NO5uRtmWAhju
9b/xtOQBuB5vttA7pxw3pgNMDk2VWVcfjAnKSnj9syStgMXRf5bdNOi3LBQkXYYP
RUTaQjgp70iIPMU62wTCyi4uaPg3kWBbm5FFEsMbu4uLdv/+/oNs/bUpnZYt9/3u
H05AzqMvj6DsvQOQ5S0G7NSjzLHd8A3Jt34K3FL7qDNB3cdmDEAFqfjoIaqbm7hF
M3cvan7LTCDhEG0RRNYLHyxEzEszN0Dz9PkBSrWS5uFc5tSyTwRNwE3k2gMo7kjw
ReU9+4RJhjQ1kDriRtXBK8ksun4LFydLAp3nxRL0eIJJnCel0XCrp62O4cnMV2Ok
QtX/y2nLx5jhSRUqaVXjT5uTwNNavmtP0eiWDR/6SxubrwfUz7P/PrMr7Gn1crDy
YUjGm+VnFjHP5HQIv+mKOcsSdKu0znD/vGjil14q721FKEvKs1TxRHSW7joCU6/m
EVHyrbeUWsN+iXqqH6AUdMxQX/TQ+PodZwNpw1S2XCGCWcJuXKPLiNUMqHSnYXMT
RDRsjZEj0S2FTjXDH4/mInfQvojraXbevpH+GZjUYo4MRQurVInsBGJghhMiOU4R
AukmZokfMBQtRQ+XGxb60TvyLBt3qcZxR0iskKkp8lNJk46IHhLkrJmIIRe/41tG
URJgyV9WX3IR5vtodemGqs4fGbDe+1E1cYOPOnWu5L87vfUGXvyMLSyLmpFn96Pn
ruoiUbvosU3mWTkG0ansC5Erp2Raojqrrn23DVvVP2NhMop76VtNa2+GcHDJLqL3
`protect END_PROTECTED
