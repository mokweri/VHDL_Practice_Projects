`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+nb+sTDNjvlA88v2HDYkz5+djriQ3bo6ZWXaJRDG8Qp8vPPQM7IBWwf4pL+XC8dj
ESHfrYBuNH8Uq5PVqK7uHm4OvcL31upOTByjLAsh8lyNQGUgj0LzyqaZx6y+Hg2U
UYTJNaxzW+w/SFrkvPW09eSHqG31eOG2fqYkyHREtPY4cO9HyG8lWd8Kqt38chyT
OlKZBcuBqo6B2cpick579cRRjoFVE+yztyTUXqtQyC0QbY4eNKNxAmPbZMcvXclK
dfaFJSgTS3GdI6FpYlvvINxim1V+aLGPcWuLU68Hb45XVA0D1yXwPsn/GdQNmfdT
mKHhF9wiY4I6NjMSuiSbbKX4R8ZKtst5Y9w1rrOhJhJY/j56Cp2ZGvE2Zj9Y/y3b
dg6hm/258QcYQ0x0gmlznFbo1zgq6WLl3iefmsZUA+Lmaa+IITYBlSmfaxOuXBJT
0dEKjyqWsPGKmaDfXKYKlCThtCOTBTZyreSR9E8Yd6sEmme4eLx9G2cCtX7z4lce
uNkOXRvqRI+rD9mm6q2Hguq6bXyQviRTlVv6HDNe0iYPeddH2Whz2VEPuRAnPSWF
bLlp7w2lhHU4xaFTKauAIdTUXTMIsURjtXEqzxgAuZSkRt3+bowLqWsQ+P2XU23K
okYT542hSwEOC/VhtSpAaMgCBJI4FU3/58C3O9+JTiKybOAy9Hyko9Wuh3zcaGuk
`protect END_PROTECTED
