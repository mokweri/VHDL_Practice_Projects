`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0ajQCsIp3pT7SZJXIwpErylFbxKYfo9FknE7j/jWqQmKTNLshyVUbv0RnNq5iRd
6WVNQSt0LCO4YZiR2wp+B+GJIhifaA2iAabMA1UBC1zm6WPFayHkmkkXMPF+zENt
3tv+euRkCcRKKqVe8yONUCqWWfEvG3leQNlriI476NXbsb/tMLGF28jKCc59toQJ
EPZ0xhVtZzqgiMI0vya9DFMZ4QOblfD6aB+w6cAgifivKob/n9ZVQ/bCP3X43chS
RttTw8o2CBuEDjj1t3UZlO3RsN+pRgpA6mjjswQHR3YaV6fQVTWYVItcLjRIW1c0
wSgB0ETuMsDpR16D2ng4HSWesWuJK8zlqYPygF22jENzOUv0deP+poPJohyfSjbC
8myepbXSUntC+VIg++vw/8/ZRhxFSBVleW6Ekj5AlD4R7yJwgR7mXCx59KOK+ESD
ZxtDggoqzV9TTZAkn95KVd5anSjFtXiikfEYkcQD35iCUvnEmBreCvBzmkmfE6BG
3VxUheaGVfKd00D3BmzCPNKK0dYc8io6DVODa0synniTROXhy8Q5xyHLVmIH/mvj
oT6RLLXlIlYReLb5Iq9NPQ==
`protect END_PROTECTED
