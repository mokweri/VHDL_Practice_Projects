`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSekrA3IuVrQqCAhWTL1oz3DmKCOGYh4AeeNh7n5FlQltSw0oWrlONodnw3Y6KlE
G8O1EEY8GOWyaXm00d/uA2/eUTIZED6yYo6xQYJyVNCJVtcVCN/YxhiRlYW5IbR8
7xpeEmtkyXz2r0maGYFDkhdO3U8ypRyxCrr/X0Iy/+wnrJr4YsDI4laEwlXZF5Xh
6Ek+JL6XEaKdOyqT4ltUx+DMlXRL6s+T9cIo294F+MnbtzPlKzxkaLQnPUP3vgHR
040hfx4zf1kb8HpAfLDczPgdMvcMNrXyKfuuL3VHY0XZEjGHNSMqECwJXTVqcS05
jLDDTbkmbr59qHLZ+c2ArM7viS2m+Fq1hwzF8cVPGLxv1XCE8ibnXzTU6MjTy6L4
abl8TSjI+46JZbprQhZlpgj6/twIt74dJ+SGHxTWAmGkrjSfosif19Y/DGc/Y9FX
eo9VV6zpA6ouuUmUJPBQBKzrLo/f6RrEzSS1BbIffaR3vxJzxVwYbTVkjKUrN2P/
fenn/7joGSO3NYHG2bmaEAPpS3uuzIQOWeGhiKh+Zkp5XF4yeMJpoQJU1ZHUJoKn
lKGEtw/TrGPuAoH8MnfxAKHGuiH2Bp3bPpCWtGdXeLv9pfxw46KSmPnFMMGR1IJn
ROjw8WgQsyqQJ+HTaJFR7B3Vpcx4a06yx76Jr7h4RFlaokY6jyCf6TL8YuUOkBmt
TzfHYpoY/zICpBTU12pwxaMX9ikdwWYyW1AWv5bdC8MB+kSEr2ML9EBIOaNFnz5K
wU8yEwhO589SQLOjcoMyi0Hm7kPuQYethvHTaDQrA1gGFw4QHGlg4LpXUU8MYFjO
MOBlUeQZMvLX2wOmgGncWy/+Ese8X5/eH5SXDpUPL2+dQSl1x4HeOedM7/Eh/V0O
NgPlgSxJ0pJs3YKA9cS900oACQ3YlmdH1UiwzXPqX8CVLgh7WVu2MBoCq3O4YkAK
Pz+9RvbY0fuhZLvPmx4yDUX4nRV0GLo6wmoVKwUkVMd3zbX9ubrPs7NVlZHznwrC
goNWlYOzEf1s3grgyBuDiq3BX+ORxqZIeX5lueSYkU0AxdF0QCb2ClCzkgSs8DYz
8FRK/kFCdsJ7mvTM0fI4VVwRrOWlabzeq4BL+orKoEyNi99mhYNXswmSqk6KGHgC
oz31lbwDDGMxCgFVCNL+hijx4MA7F9DqR7O5BToiwFUVx9ht7ZoJtLPyw14+CE9W
Cq9iqAm19u+ox6/1s2pFQkaDHK5veu8uDPnZzBNMRKa8WgZSFEUVZoSRvCYl/qq4
33EXdmlgChcAwYPYJ07OHRVUxp6PYmZZ63Edp+LIcChr3MkFhLz/psX0hAMHLigm
CktW3dp3yh8ZqzDGR1IREzYjwW2VJYyp4Qb/D2XFe7FbgIAekEHZDeKWm9yZy1UM
4jqeD4//7MktRTv2chc4nqD2/JaqDXR8i3DOzEikuxFwaYa7pmaT6vSS/saRwZZx
k2iRjMxfvs2i1yiIbkgoenefOr8XynnFPiqE+VD7GlGroMNc/2Q0t8bRKoVvy/of
Ygu7qXwZaWdxugYJlwnZyzK2QV+jzdMaIjAvmqi/hPLUo7CMfXa595KA7N9q0Osj
SxCS7qqjgAc4ul9U46TwOTT1V4HahgYGLYTt7fWp9g7tP/+egAFrrx5soIX3uK1b
rZd5x9KFlTMF0O58h70Q5C6TXPwGnUMpAc763z5G+4ETNeJsQ4DpuTdjSvMhJJ5I
EGkTkVX7H5IxYKO2rKQgPRdupz5/+UEBl0KZkTBWXWFyDCwBdAwJYRMwNqbh/9kQ
Zrhtmu8wq6TwH70K5gfulSYe74izpOateq3qqgnT2V33Thj0Vs4xEanj0PfkL5wN
F+s3kiJx/qkcEW4EBYW4QohBGlT2tCl+rp7UQMuxMOPrd/o9y4CMN2X+xXBmGgZY
CFnjiHKvnDgoTmS6O9ui5GspXowU+tAacUGwZSBRxnFZTCIhdNJiSpGnFwDrmmEd
ebSCi3pnCaapT+6VKjPs5GmYvWdYlmvcWcZBeCta1+04L/Bu0IWiCnKjRIszaqVm
GJdyFUTNvT7c5iiSXAkAfTyZp255MAQKl/B333y3brueAorWHWSkHe4wlfmFTEt2
hm8Fjs7+Nx5rVgAKcHoisvu6s88iYI6Xg1mGiW4vlIUhX7kE6eodOZOd2VuBbxHn
YRjLrDbVE8AYjyN5a+Wv+dvQtWorOGP7HyjED24APWb8f/P7xO7OJpgIpUP6EAV3
i2Ll8I0uRRH9ilc9JOKhTJWqAdcqrtAzBdjHWnZiGKEG0z+nNSCekkDdGgtvjnAR
Y4iD7cWk0xFtR477DKljMnY9m/RyZPyOkNna28jTTVwW/om4vX6JtptBOzz2v7Lx
EGGXRhp/ko0E3MMlFqQq+pjXc8/gTEgzd8HM13fc6JRp8VhcyjgiT9Hdszr0SLPX
BGoOh1TL3kx3KbtkOsMWurzapCLOjGjJGdzMKdifgCwHkHGez68Q6FKJLNT/TDHd
5KdJA29goztG14BjCJ8qVofbqBaJIS/OLzRF8qrBQKonUOrcD7KaNuLXlGJcukd5
0j3gouHUpKiM4FTXi5wpemEShWUlcKuyMkzR6X2OPW2DF2HZK271uF7evxmnvItb
CdmO5GJQdKdoE9smcgpptxNu4fLvaAFXYTRYJ3tXD8wiSeK6yTluwwhjMtHMFeB5
8be6/Aj6MPr3ngBpCnCHtHjDjyfAKDH3vHiPPNbGJbQcfDqEH4Hhae+BeuLalluF
P1Nk2+CCPCVM1Nd+YhVHsv0aZXzUCKRXcDM1zT5ojBaqt5v//TJG3aD3xjAm/DJR
A5xZaQkYqI6M8HXzQh6b9hIuJ1AgXLcPoINxeIAFF1DfdH7bMs+3VNRnrBYqHeZC
EbQq2VqBMYWyn5oaiof0g71lhHmyrzVvK7k6Gm8OUWCXcfjSioAm3Sr0lLvbB8Kb
HIUWe0DnI92Pp4BZl9+xtyKmryK/r6XAmkELlbrepCkSpATYXpF44iNY/UPuUeOb
cl2hd97Cr4lL8hp9P6iPywrYwpOnqhZwyg0LmKHiBzE0vJSbPhcP5HjIySHZtelO
E398a+Aeh5tx7CD5FuY09nqhZvB931NgAZ5fGupRLoRiInMjK/zus9CcjkXS/Gma
PbB0935vNpSKvyGO2Jlao+hJ76+Vki/fJIuC4AcDi6nGAMoLKXRIdkIEA+sKhQTZ
m3W7/QKyaGXEWOG8htE+pY3rgFFJTnFxs161Q76L+MxYSv66p4KlLufHYBktbct5
9Zdban5SyZM8j5jkpV+RSeOXmhU4+c5cOXy88ysLlrlPx9sriUDHzmUvUNXf2Jm5
1pWpg69oRe4SZiQa+7cciBvRl57qpIMCGURqEHg08v/Yv81l5jfrIbEGJb8PEZ9T
BYivLLnEvzYUp1X73+aHwVXycWrVUP1x/s+Pedfwk1306PegO2MpzCGHpW/w8FEF
y9ZwrkroYQAVH3qs7zB4FgFec5C5aRKOVu5PfdWf4rqayINFvJrCFPz4DEgP6DBK
dcqNLVnn+2KgxEd9pMDsw1GIM3pUFkalyHMz2078eQlujbEVGv7GHsomL0X9CBzM
G7ijS92fGi8aSulrZi7sv4sQK/pbQTSVqDm0YH0rzFFElxpHND2REZjoi6FFVLwk
D3p+ivZLSIaOLGGx1VL66zW2yHzzJ+S4r4/0GEecAbrsB9g4WOwLJrKq0fWtWWKv
uTHhDSJ2PC8Jc9hOJ0fWj+w1ru0yX+YWR3QTqMFGYaGtk1S0+9TGTb8tf2zveCtA
tebYQVTENkM+YZSZx5VJKPM27Qul6Tu8/KyFgD5r0I+lSecb/mnut1YN50ybMWvP
XwglHXyQYum9AfkiInpYxigivbow6mdutpG8uPxaRD78E51MXBRmG7G6gr3gJrRV
1swzSN2FRPklV6kMH6/n98i4fVdf3pmNE7oTHStCnty/JsHvfIb89x1S1T5qjQRn
pmSUmKsmck67nTvr2lWF7T7t0ukBKmUHtjEHuE1sHlYtPED9fZD3BJjGyTT8Skrl
cXGfw7GTOrp6lwq4yiOl9QN/OjmSB/h1hgvrKmPZrpbuztcxYHyAbQEywBZbr8AG
veuH3CrR99QxcChymfPHqU0YZSecHr8tAoALQNzPckMEBU5wYNZ+TsyVJFAYGjBr
AMGdkvVSrB2kP75jOcXmBf+g7btAQNq8C/5UgxkHZe5l7Q/JZDxzvaNIEV42IBQR
IAzmUuvJ9ItWuAn6oYghPMCHwXP3P5FPv/wR/nIkcuPG6J8omTCVAFBN+zZbkwMh
2Xqhqp7YxJeSlcgkqb+Mst2atf2PYZP7pck/lUjDVFuV6X0sSjtCs+ciw1YhhOuO
GFoD/C33rAWIRLRa7FeEhKmiBm+T4bWdYYxXqVdev2m1fukoyVZjUVX76e0VKXa8
En5nz1hagnryboqK+j3IRj0lJYwQj9AsZtZ85BppLPjZs4jzrLdFB4XKSRAozk7v
JGpJ5pySChivk0k9XTgT0gxs2529RCUYdk9HGF7aVOdTcuu/shz/yk3r64+IUvmb
f1+Q/PT74UMGQaQsPQ8xC1XeZMRELTrUKnNWpmrQ54BhVM86uBp0Y5kZS26c59+Q
mk7OSzKP4JIbY6Pf6tx2yE0OYx9qP7stqZZeTtis4V+5fP2RQuB2gj3EtESgj4pl
S+QGpWLDNHZsdObn1L2awCg1BXqhW8FjHBIqBkxjozyX67SPue79Zs6vdn7IF5ES
FcYJQcGGGBJ352QMMoFzUntN8z0X/tFNuvkbEaU0djUX7jwcl3AO3PpjkKWaiiPg
I3h0F28tPLumipdFuPx0m9tI5oPoPf9agGSEYiR0ycHe8Xl3MR1gASEj9usbHI2A
EfmRQIrdju9ghE01jpL5oZZjjwctMhtFD9idKna2cXeIl4hMBzLunUZAqx0gYKkI
gYaVfHuq28eD0SQgDQAUCQyjoItzp2CTGib3I7ObGMireNxwGpobZ/TsDvK3jSzi
Tz9O9vSQezbjaoTVZY0b2oDhJPQy7Y9jOYHboUZbOfHuNUYNsSQhnK1vprytXBNh
FqX3F42rUGPraifLTQgMg32hkJ10CQnUzDoTz6NdohMidFNGXQj8ZZV00fqRjdWs
eg911kC2mOUt1OVhkOsWui/ebTUrYE5GEcFtgII2B+kW/5G226RcjPMrRQDzRKeO
hM7vRsMyeFtVGP51BHNvVSBEwMLEn3hVf6G4DUjTPMkC5YGDJbTK9gyUgSmfxCVL
vUTRW7rN1BTMn/nGYVK7z1Ek/0vUlOq1q1tfoqeFbFQEAIZE+OVdkPPfqTJDmQ7y
C7jGylPYN6iQYs8N/JEvd7X6mCgL4g0/P7Wnvrej3gd6OB9NSh0q/wtQwusS0/cB
9p+JUe0BKugvj+jL2BGMSOlOtDohdLWtwuM1Yw5S7/gShvYTNQcPNOF1TBlHZLCt
VSBeM5MU2Q9mhXchI6IcIlJ5njNooKqjEKhf2GOPBvXvFZe6jgc4P6In/gYWyltB
LxGB90DvFmZ9BoFKYTBjuPOEeOpMPyZwiL5yhmmUMv5R4FXkC4esWiU0KSWJ3uu7
S7R3ePhFhLF88F0jrBtQxSkn01cBKCQBm0/K2xoBZTA6+PMBfuIkdawRbHnbMRvV
8hIuZYrnXS6P5Y0czx+AuZxxK3pOkNZWo0tSLoHmr4eE+pOARvtPp+DVUhPQ3mxV
J5JhxAtc+jH/6lcEgkuK8ddknKjB0/KYv/C2gRfdw0whehD95PzVEeB2R9ELstYW
sRsWULq4stmwxwN9shbG4TtArVGU3uKlgCC4cBIHgEXIitDgEiCsBLK/ArLUT0cC
nJWDTr9n+3FOC4BuGpJ0ik2M1jZcd8rSF1HeCVg0jTeoqNjmWnw6CSz+g2CGNRc1
Svu6opNfzy1tcbIITDNHwtwW3FIIH6PueR20dKnRJ8wFEhgfxnTzIVQh7h43Mbtd
Lgsytr3fvhx4NmExvHQo+MxGnbGxDjhnrLh/lsoKzWobT+p/H+CljX0u0TE8aX3Y
4wTRm2ua+t1njhQanF/3awNCfEfMMc/4n2YcwqX/NF9hXGDnSXqWwgzpjnJwu6yz
7sBd/eoXMbFtqb/gTCUQERs5I2QWnqVOMAcGfYLw3+jY1fF0Iye89HOcK23YIspt
qZFy5ywmES+i3SVK6PGKeiHAIgRGUMNrXIP3+GC6BibsSyZ/AdM2cW5IERdLcXBZ
SJ1RGoLHiE95x3M+cPIKzv4NdES2Qa+Ba4b4LI7ulz29angRz7VsyTuvQjmzPXFx
3HQrI0VtF9TRZL8hb2PU3AN2qC75Gvwa6xvUGsOW1iLKazIQGz+bAeaENEntvYco
VRJyYm+WxhuZwJr/YZqxjw6uyDfUi4881OW5jK6Jw2ZpkfQOh6nd1EMr4AEljpwG
MoYKEOFsFsU4f5YwT4A8Uv9w0XGbMHjy2OzI2qRY6ja8sBRLcpJB6PkW4MCbbsnD
+LlI/OSyEfmpL4CmL9d0NXW78fLngCYHhPTlMEVSr9vFQ65FP2g+VPEcWFzCWgMZ
kkcAfuhYWmtY5h/WhfCVb7dHRVYcwOsd7i9kRaEeDOc47627/zLi+Df0ghESEA2F
yQbXl+v9oWmaE6sxyL3WzKJerUGDjQ2Y7KtdkECTDULhIz/4MHTqEIYZj9ItXLnc
9lXVHXpF9VCxKuGhLDjrNQTB6ecgvodSlTgyEYRabPQtKcXBpetmV+dElcM9HpON
IEUPcaDvbniX8BXLkT0syRYbNoFCyHUqjjOuHYxGtwXKJhf5VKUHOzUx7wMqTpqD
R3iAK8wAEEC/NfWJ8quCuusTEyBkXZqvD0yvtXnQhsRnFfEGI99k2lMm0AgDJ7vn
Cqo31I1schHGUgCQZmzJAkoz2Djr74w1WszTgimzhN59ujd+FTenC/N5HO9jnP0z
cyT2LOM4+lGeVR4OUSCl+5ARZ6OfHPV3TTEat3O08xg5+0x/QmAHxcFAjLppQ22g
cC/PbHjRCSSPtscEJ9B0i0OmeItQeKLaW/WhYg+GSHGW2avFwChD9veBHo5exlbp
gZh8IKfOjEcUY7dwn8ukLD0fDLGMiOQNFNyEsCaQ3m6dtR+v+dzaYMkhDHgb73ZO
tLclCEU9i3HoWi0cHMwUIWBlZuR5seiFhzp+EiXY76Rx5YTt3d/5iMpJOAFi1FUm
AcIzMmZh7p9k0ljrJAKyN/DcHrb5ZS+4wk03gu1SHjVwGOzSqM/R5zcA1qOGSpk/
BqNcaH8pHGu07rdmcD1UpDGJi3434jD6S5s6bygHDFJhMPVI9stbj9UfWzsJ1UEM
LeaKsetkzCj53+TRaqZ7lPEfraJhvvtc5LdB9EAlGADm6duWfXhhFKbvXTpJGanq
Cflh/H2SQF1rFXug/N9iI79zeA3MZoyy5/YIjtYJXRbRA03NFhFdvPt2lN68qOcC
p0EKx8AUXZ+nogFzwowlA/DJ8gTwa4+RkYZmNKGpFija7mohJ3PK7WnPWsARxyZO
RJKNgAi6pExy7XAFsfqZ79gPb7bLA7Gt4q7XECVIrIQZdyaajirbsE21usI0YA29
Ism0ae6nsP4FzJhLH5J2Ijykf33ffbKzr0Lamts2KwEsK2YyP5V7fMqo26lFC7eh
2ZCwieOIcvi6GSyw8VjZGbrGbGrTugF2pPjb3u92lD7XFIZfJszv/3eGY+D9WZgy
/1DxaDfBMLThNgtePH8iINQtnfWJx+C14aBGwFnnmNpTjrkPW4PryUEYVLG3z1bk
nKVtvwEsHkVvzZZg/6h8fAAf9L3R0GOEBfqzNy8emHznAzmc1e85eK2U9h85tVJl
2IvhWX3R3cwYtcBBbnl7b9bK5fb3TGpMV/nrgWtHbjmHhHPeLHcmF73z1xzIH7MM
7Iv7mu84w6I3kVM0wFE5Pjn2L/VWD8yG8eOuRSIfWJeayM4T9a970N6hDsGRUaGA
XzEFfYc1b5MQdqeg9bEv8pOfBUCrbcLtVA5Of4OsQ+cxoooleePl24k42anUAWJt
sgburpV5vPmQsmJEQ8VHvVmNSIhoTFaDsCo358tvFAW/c++tne4q9+o5IgObi2Yd
nEHHqP0vJd5NFHCCRvTYR0s+F5cGkwQhTpZwDrsZ461LpZ2LnOKnCKaibqjnBAQt
sr+4bZgcZZMKew9kDj0v7f40K6nyiVIfkyOq/H/HZ6Vi/XR8t/KjBYVShh3LSVnb
U4N3n746+5DcxGo+cmEDioT3ts+KUDmPpUTuKHFdk4PetrpJYsiVAR+7WYYA3MkD
nMtVY/enMEGe2dpKKr5qbNcvjukGEVooKdBnrlUVfwWGTPNlv30C6/CxYx1uLUUW
seUgb3lusNco/yWVxzcszF6Il+voLXHXRrUztP02eYME4SggTWdocUOf7zcA3PGR
8vG8opj1ia3VRUc6p9KaCEuWF4sCgx1qbZT/tci/4DNSWKZFlFwaFy9iPvLWfcqY
JvCFoXmytDPvCzWAF3iXth0NW0RMn3HGri2jyWm8laWSZhgcudIUfi5ik0R62Q7D
jj4jN0BR7wNjKiJDeYGMrRSA+L3SZvw6vf5O3nH/KajSoEI7vnCzq+z6S4KTCNAR
kPK8+PYBxC+fMye/FgdELI4yZJMzP2tPl6gvMrTEsuBg1bKmzrZKdQVgM7ZnC5Cw
GhmJOe0rRmj4NeivTqsyTCSbhvNl/w3u5lRs8Wk6isvLfe64OM7crOQraokcAJBe
S+/jSHP0kKXRSgM+khBQQpjdxlXpHH3j8UqV1FrT7ZTvhHvVvjjGgwXejbh3P5wh
bbuEoPhQ/30fVi+IOLgsTVUq+zR0QyKlETfMAVNtSpB10RaxF5IgqInlAau3mEfO
vWwypKSckBvhamKFN0Sx8hYeObBx32InynCzhoL2ZGA8papAZ8I8lyYy4IE2RU/k
xkaqrjPH6jYlJjEoskRkLVTat4I0YXlOQyCXZ8vZ0wRHn7VFKAZZbtmiNFMhB0Bu
yb5TnMsNfUqXz4X3BmKCb9AhqOFy3tp1suAyNgkcxjm4nPmCL1j4ofWHKIv2gSMh
T3O5oalLLzaEl/xBoSd7rhWZmRYTnxAfYkbeUHUzNKqm9SKXHQBacYGq835/9ZEA
3RntnVYZZJcOmu6n8iIbHehgZHWJ4Q7PtdI4HI/YT9rbD2pm5eBFEnOuFYUozVBz
pJHe7SXYnc23AXKN7or84kLVhCFYKe6Hv8LXQcFeMM6gEHSrLXfPY3Au9LEnNMhv
Evo5xX30+yJrQTgEIV17JAomnGDra9fKWN6i2ca4WLR6Tusp20D3c32nVAkrad+v
sQ+JVsG+pvhdjY1E6DEE6gqfhz5qlhYg9rdSjiENM/bDc2CtLpQqcLTqOzB1Nyw8
KHWi20DWanH1hg+agDYDBJIEl57H5AG5Eoe7Hm9E1mS4JifdaaPCfukgVSKDhmME
2fxv0UUpAK4DZnDrzLaQ9t0YWSOdY4tfETZcKaRjf226tXYBsUA+KYCd6yQ0cAMD
Nccbnmz+V9iK2NT+bQIUHbz7y59GxXA1IaVJORgzfoxfY3jEWXgvZraOW86RZtET
ozxLCqqf1GLJcC1wf90uEPXzbXSf5EFD86UrNYgzclsD3GUqM2uJ4ICHvlTpzX6i
dRL0zhgD1C/mdq3l3dkE6fkWzeqBRdx//VYgATL4CdOn3OY5mepcdEDmE/2hBWB0
L3f3bpmnB1m/OCy//Pm2tpvQkAm3bOdKHQtdl50hjSQoXhlX+eCIQHOgvcr/1HrZ
fbD3Wp2oWohkaFXSjYh3hIJ7y3y29U+wdas7b5WVOvescdfYSWfbk1Db+rtVo6Qw
W0FWGSwTmRW/O6Zy1/KDiTpxfAXRhdCxZgxbUaXvyuHxzQfZA7CI8BLKh+mlwPUA
w4AzBlXEA7Qy+LjEdy0o6lVHy2aAQR/iY1czhCE9OyvMZZid/OReHABIkiuF9Igz
TM3199EOtJqcKOW+Sd+clfgIOEyfZAgV1QE1vKvigVOa4anDY0heDObqC0HLaBt3
txlplLdXQzXlzDgYyzLEHOk5c5D6uj8H+38m0zxsk4+WZDcpohYqCCBgaEOWlZaV
hSKnYkgT1Q5VGk7a2yw4Rto99QJ/U+fYvcqna7CaW7ot+SBj8p4k3TVV2vqPdTQy
qvaXncgBcZOiuF624fXGZDVnRmV01fQFdCvTve5yRYbHocIXNw5e5Np2xdUv4JRB
MKSI1P10PQqrWAVycVJSUbR6cWv1nmsgUv/ExNt6XW5LZEB5Er5MvjcdkZzeozIa
od9u0G/HvM7YBelV7TXLV+794qI2jw5DZhEBIeasZ8ai4/TKJBB99Px0Civ7aQdg
zpun0GUtsnmh9S4fgd/vcRdjKl5vQr6wVK79kfKrH6yk1C+CaeSvkGwBfGxLi/ww
h17OGv3AdpKigUwmUBW+U6lC0DxhvF7svB1uzW9Eyqm7e4n5jtElmFdcyEEcuz1k
vUs5+RyVOQ5uY/QfXuxoMYi5n3zwtCAaabPAmMuxu605pTCH22Qw8DGl1CPqV5Lm
oA32oo/kFRrteviAfvF6VabtKR05QqSIh/u2zyVm4KTCUHdclpjzHwlRwsDTXY+A
dhrXCdiWZw3H3cqpuawvvrgn1CAd4ptAnNwXLQsUVJqpX2HhQrOMclX7ViIdvv3k
34QEhjst+HVmrIklTz8a9uSLF+0WP552v1mf28poHoR1LzCFvM9u9A7a6u5CUq3W
oLdsfjXlbfHYuBD5nlsIRLjWIAxOriP41/irBaOIjfiTSL1T1n4nLam8pkO3nIBy
9gIibjPD8y/fEjcC5l7YrDI2uCY0DnoVBHT+lZSUj2b414/QCHLZV2SzbjOa05Lc
3dUy6hfmGnsjjtLDM6BXln7+hNloOxETqpsHRARim36wktGoTUYc9LOZwBZMqts1
W+MR9J9836cC7ReYwg7QrWQavEBdC51X+exTk2BS3SSU9EzG/tqhCVEmPpr6EAxh
VesnziNHRCxGKjeUrApYEWpNZPfzTyv+d//+XRSNwFHZ0KjEi7VdPdRxl2fNP/Ds
+WmWR/u++Z7lXAxmCQuXPydEfxk7Pd3fwAx0i4mAO9wHItuIoLeVQL64K9PFC7bL
pv+oimYxNwzW0QdcBjQGtvYXq9dXCzVsjVf4EZZlmh+MOR/7Aqg2NLI6rJ+h6QoN
ShCBodqpRa1KnX/gvy1lVoGMHNSVR+99+eY3tcqs6i1KKiBL7UB9ts8Q0Q1XMXio
YXloyUyf/saHOamB+cuYWtOlLWcoJMIa6Sq78VU59cC6Zj6UZplWr+03g/77QGgd
4gLdOg0VVhNUFhtqCQUfQ81MY4+p3pgRyhtLB9MOmdnPbcm/Kr2JCQRZrUYaXr+F
kX/qn+ubvYL8mJm+OiwtjHGyrFCUZy8sNpVCDyoGTcCzoSk/2xMnOjuWQJkIxoD6
tEmeTVYoKLVs8dM+eQpmt0+FwFk7ShV7l2MReNe8sXTYiu4tdVH0fFs6fC+Vc5pv
fHqoKCs7glGatZxiCzlg5nZkG+ZWly61XruxSum/dfNcBZe/LO11FeSnwECxCyJQ
SKwMeEbhRZsOWPhbjawziXJkMlMx2JsjSo3nzGZp4EIozSu0Hix0uoAOc1a2bScf
xl9jDzjWEauTWyR6WwZwnnG9JfQGA6uvoKRjq4F+D2wwL2abyPM5tFgDALxa1wl3
8NwujlrtBVlZlBW8+hdr1rjddXuP0LMKUUaaCCvaeJjpwpBMXwLIJSE1jRFMoabG
YinYmyCFt0zLH4I5zDWv6IsFZJHHkVk7nGanbgWSRDMbwujx8/RQDZZGhSt9QFqP
r0MbpOG28wfkhncC0LB15k1uUJhrrSQoDKxco3ZV2GhLgF4F5rXvPlims1c6Wjg8
y7sX2kaVIVUSrMmXgRTZA1XBiQB63UMSfDfF6r2jCh60SR1TZl23IFpER7O2kP6t
1oBBCso3+b6ArzNlEvimUyyR2Jx9hU4YG11h7ABM3mhkshrTiub4tqUWvLeYzi0v
+w0BNo/OGfR48X+jUYmu9NBwEttzk1D46gYIbU+hwBwXCYIyupevEbrTXJbat5JN
vVMRYHpcJTdG+d5jZjSIQnxTCD/KFIFeWpWpJv9oNjDsie1c22U7Aits9xBZABlK
mKCdkRWJ/RDcEjTt2Ekfr34GEGsK7eBX6XZ72NNu91jfl1TttHfqtHG0ThLdISQe
b4zJ2PearfT+Lu3TW+2dUky0nC8IbeR6ke407Cj8aRHxo0LTakD/qfdOLrEA8YcG
SEcF2mF+K7YJ5JZlN5D116z0lsAgiJPYqnXqtSH/NJklnajg06AzPcRRzlXbyAKu
7KweZSKQ6OQ+Zy5pcEpzT5j9Jfxjb82X5Ymie55FqBE8sCyrmI1CJ7+OaDWceM5l
SR9x2nRsg9OlRn+mfxkJvu3nsBV3Cs5DShGm0o2pZAGjqaHiMeXWcIpURa/EElVr
kpBedBRvFO/90oP0KlWwYKq/lrTo+MF4cFL7phNoLhnPY0yeRQpJxnZjeWo4Sn6K
WphdukvWd7bZJEpFkqPAoD4n8XW1zYAV3dDpCAU5K3oBy/gnO8uXcIXT1hkRia9m
MBpfuUeZkNzSeaqwLV2B6mz0rAueevaBCWD0PH8qOaIUqwkTE+uYYcOqOjGpIbKo
/oxI5ya6smrTTz968v9ma/BvxUfLiSdhGJkeS5r2SbmRkHYXeEvxB6VVAiizJL23
McqT3j3+cvnaKPK4zLqAwjuLsoK4QTVRnxyBHvw159heoEbeomFYNCzj8sKsxEav
+7hTUV5+0vZwtBdU7nuTgLw2hp1CWYjDCMG6Zjm3QrjNv4kcF3FYFNuQbebNsQfv
S4/Py37+XW4dYwWtmmGul7s0cNtuhSteATi3azo2j/a3QTOwYzWVuH3Eu4PKLlve
bEi9RHZAo2Gcc2EEwczNTdIwIflYfKtLapPPzCoHFgG/KQeE0MIRYyLohqnMaHWP
PEmKbb3a/UxP63r6TKVkhKn29l6wSrPJpCjyrhiUAz4UtmIqz9jCkkuS2HspHjq6
l4ZsCuE/etWMiqa0DZAy3usWBPSIkulp2WS5lWBRQJMeJNLdeV4NGPLlAYjIQLl8
vc7brHSVLPcOUcW5hDFyVivNb+LKc8OSndPh/HPoQA0KEBiDUkfoLQof8Wis6TEo
li99nQmO209JpjdxpVFjhpt4OmTx01sHkPRBuy8o7s7blirFdhLMJUA9Jx13mF2K
abT9MV/o0fZ1CBAPp0Qx7Bzc2+cPvORuTsb/+mdJTEIG/NXSZEbH4Ab4c3FcArmN
UWy1kMW8zrPL5TfiCpb9tFkVArYcrtoPQ8NZr4eIa8W4FkDvnDcvHzHTjathlt6b
wmmbgXjK6tnZeZ7//y/lSf4RwDGRpiapRjYFqSh/eHOHqSRqLOJUdk+46LZsvrGF
PbcpVjHVuXV0M3mgUgwU05CRKqvMqAkFwyTwbJ0dnZ8UB9XxRaPES6LGxYJi23+W
KOY4XmknfjFQfjYYJc0OrBf6tBbCqjYPG3nljhKWmgonUU8nmoMHuunHhTu5DZpf
cT5uh5Kc4IZJxGFbNNMJl3mhLvDFd8X9+3UwX1fX5q33OWYU5MTyPz6SCtQ7FbRs
BlE9sZBqvQFn0Blx85yCuKr8YBa/vtXqXUIJOBTRa4JPdPvbY+sA6GO38fYjEMaW
1ORuGjpk05tzbC10wY3gzNCJ0JoCHqqTRrQncWMY3LrGpV8AYR386rlUsSC3MaC4
QcekqysDTHS1gh8t3QzmJ5gMFSbP16bMxIK8pnn5lv5QUzOBcpTFfCnUWz59L7gb
B5gOhYfYKVpiqQ3ulH58rdZmQ+1eAwYp8UObiLwG3fvTqoOnCdUyzPhgptcgGu1x
WkmXE6EErJOUxAcle7Q8u2EvaRgb7r0FOYKs0QA1EKxQrHCwdHjuFSbOXWDBdcAV
+TbMEdowoNLW7W4wY2ymHfTx/vaCG3sazMrqjtQyKCPUlgljkWMb5AR42kCRX+Sx
GR92GX4z72KwPrTh3thzw2mZPNBqzDOR0OJ53SDjlxrlnpMV8fh23/qPbgPAb+CV
9tnheRBedlFAt+Ar5V8KV3TpIL7T3/7iyB2NklIpMAU1Ja9oYClF0o6IhE6YSwbm
dRwthjSTNY4U142Sjgry7BhkaPtezLjMdh+asvA92aZDmmV9awzquhW61YtEfU8S
oWc2iBAcWkmoFEWcIety+3O+cg19jjcKApb8w7wd4QPYomrtwKKDsFW7lmCmzvfG
Ijmyi4wgZVqXlvvofeVESuRKPIKEljtOBEwG1TgJtiIUv9QWHOpiWGzDiChjj80y
vsjpMRAeu4ioSaYlMQkB9gdyoB4ZOGNL0ucL/gtw1+25J+1mnwXSwDesjaZxBL7w
nixKrV12BAcLEWZWaitKDU6TaX+OI0pPNl9yuXtd6bFiDQAGGgGmmnUgJq1Dsevy
U9cOzHfiWz94XNbab5Bih4oWbA1vGHlMuhq1y9Sb85N129RrArdj5lNwGX1LYjt3
lgR2FPUXQPwjn1EYgoRklnDVG6w+m+lI7/9hDjjdTHmEIPLdApJdrb8tYLy0DgkK
flBSAnsVpY8kYVw/aH3vhVdR2bX5FIoIdPtjMHLCQ2/t20ReX/01T7dH6hVvxBSU
Nj/YNTDpGyEoSNE8aNywWrGj/zpGDQXedqZSYYnIgNLZDn2HxS5LYdX6NkD1F5V5
j+Geckcl4dY18udu3qMfYloC5rANo6EY7TU31XWj8hkGIFVq+vmZ5IFhCkHI6G5O
h9pUaDVMY3yCO/98puEgV6d16qBw4FjFD3LpGFZrx2uKklIAAl0Eks9qd4mwOKI/
ywRqifJ2w9QucRtwfu9JHyUreZPsRss/PFb85Jzpl15cSxzliLzEjZbCYzAc4Hwm
rmwptdZMA5gFEx7qfRK0f0BWuEnzdSLwoT1zRmk0AGvU4mTR3lVm44ghd0FUQzxW
lQ/lnhIzdIrzz/JfnUpTp6L/ESdfcDyus7Z8rZNmoqbDqkvhRBxTlk2IvgIDAfoX
x5fS5fwTCcV+/9/9mdItud1kRr1h79+x9zmV6pQM2Ben92AE7DTvoGtVUDWEmjU5
v6maAqmtG5YREGQRI0fnoEllZBLosPFHMBKb/8swyGeTdgl/5yzN9vyOv9zlE/Vq
M8R5n4eaF3x5tWHsAS7xHK4tevb4W1s0U4sxrDvYPq98aPmIWFZusWeeEl7xW7JM
4LIe0g7dwPjFow/1kDW7FTNYgsvlhO4A8qbG6ftkNX2sbO18Gs7pFPzgzT6Dqfp9
SD3GArXD9S6ZGRRZ+3EIoXOamz1F2wti5nbUAnHdB5AS+JOwOkSSTg1K62szgnou
alTd7YApUhaQU4SLh7iLaaw4FRyCu7VQRUlUcfQofIi/6Wt+CSey7pFkUhcL5t9B
JqtrDH9WOJuK8puBKU6YPPYAXYESdc+fcwDkWuJ3JegIkMNlhmxJenH5R42lPkM+
IY4ml3cyvA2ak6yscxLYDokHFOR0YsNOeDaX8Lliw7D6wUstptVd0SWLiVLKCEJ5
mIRRR//DJWeEC5OYE+kmkDYUj9HNfP/wUU4itdufBKj8jeDnxJscqwDTja/52wS2
YGm/mlGa4jNMuTJyEyGYTqJH8ZSKMWs9ni1A+gFSrynKVfXiLTH9ZFU29QjAZYbh
LyU/L4/ME5NUPw+RrD9A3xT+/qFCjxQNqaZRySHZ2yf81/t61dRdQhJhPTeWJ2kU
yxAe5jwi8Weov1su3ahg2KLG28kHuPA4StTYiuECHp0VINlovjtLt4pMeCFCpcob
733FL+cm61GtooRR5E2ZfSPHjFGUJITJlThrLxNoQYD5HKIPxpmhyzvmH3pTBlwE
kIuD/0f/s45cWKZrWv9GNaWMbczMi9p3a884R8rC9PcuQwD4dTDgfw70SpSpQRAT
op7lJTcMlyfNYEn898Zx3UOz3DkQUBdChUg/ifXXxAr7dTuVxDQ17SeRBAxHMQTo
a//Xljp5NboQs3QeOJaSpAGEPq30kgcsjsAg1WYJZjjGQKaB6a+/dlgkP9zxPEgc
EubmfEHjDcpocibcM/EfFHsj0AH2Mx7TSWZ5ihfLYRMO90EPwe5KhBL8TMaChiHA
/DgopKYIK44s5KNwo9hunICRWP+8p0SegjKkBK/ddRtC6j0y/dwc5ob/iOiE+5p3
6VzJUDGr1C8u4u0LnQVRJOo08csFUWfKZiBAVteQpLAvHEPF3/KVBL5ynhWQIHvL
GP+dkv+LreJbo948XBACUTGtkfTTga8Gs07vOQiNcrFjBjU8Fh44iMf42w4GgHki
rylrOy4ZGSlAZQ2EUsi8Tm6P9Oj9Lfb0oVy8r3QWHdVWYP4u7XaMfik0ZhL9lW0J
UC1k/5DBdqfYzyE+WE/16nXdW6xQiHHQKZvvt5yvfNY+tffb5Y1X/qCgXJAjNXVi
EaO68SnHgnMs4G+DsR72hUjoFEE4H9a/zRPjoT/1tR7OYL/Ma2nPVccBX20sUO8v
58eheCoNg8QZSp1zvsmBthfj2zi7d2A7ytbWMwVwdIEb4xb7e2/CBn2jvs51KHyF
G9nj5jAHdkEF2vGBI+z2qrWceVVpmsL2seshpMaMFhaR238Ap8Rz22naHD1HA2ao
m8uHEOLs4JHeesdfQ1/I8DVosnDq8aAyC143DQH+p9YDZD9/p3BIunjEdJWaY1UW
1/0GNn5Nuz4sbrinfcvcmDSj58RKqx3pRWRHpn2oIhORw03cgBpmQVbDQLHXNVsn
9rAUM03ojYjdHIXcDr3jiZvR7TFyz7TAUHp4CPj+f6yeX5CODFfcZBI13YGjkk8K
zPtaaUOYTkl74FOWnkm9tl3SE6PGg3x5IQYzhEkGpb8Gc//bnUvgwaYT7Gw0xWcE
1MHWJUX5K95aKD2mbC+fSrkEOvhs/wPYQJq6JMDxUKaDZiCakcdPrFZA2uSnrQcS
ChI4G6dZZH9qRHJ5ndCP6wy1lnLHlJl+d0JNfcrrOKO69786e8fLL7m+0+x2+12y
8Sj5dLYq/zJQW59hz8YNJdoU2A2inxVoUPwaS9RJ2Sz0MY5VDYVWgs80//9CJAhG
DCK6X6Ir2h4rBs4ZsXjQfR99oL4N6kcWoigvQHjUgHJtJqPRrvRRL51E5eSpSwSG
S5FAvls94rr1MkNqJRWVVfh4aHhHX4XCebTZYv+iV1ufNKC9nVrLHz9sZZdpI+Sz
gAewdJF0GIleLpG/kB3ppvMxDv0kzkPf+QAIM2Ym+O5RDsv+ZA5gDAwV938YkDLR
0rM6928LoaktkYj5hzs2xr1vZbKWpxrfyqiYq6cspAai9DiEiVQyG5aJ57AarEVW
AwJAWEzFmPsc1LRm1UL4nlJB2RqE4Iuy2C1KQWaim4DhgBWy8hPip/HhYN5PWdFI
xs/Eqq/oe7vHGCQoB91pbj6T/O4f5NJsOGuyB/1IOdzbv4LXFs+3W4KNoTCks3oD
Df6lVoCxPxNRXPZoThNrDiC6WjEdCp93f5YcCPaAkFhY3BiXjH0jC/tu9cK5KFPT
lqTFSzlsC1dKFiwVZhB9etIfo3VfpSdxR5ac9Z1LrmANKVYdzjBuVIYBavtqvzHW
KpvgjWJ/qrnHp9pFDX8sxuAJ8HXo5od73fh4OUpr9Q1pV7MtrbSwyCkQKml5P6zG
akt8FQuDDOhdPNNvVzSgZuEyjfTnUqnoaRM/l961A6cKmTO3KqaGv2e5bx1QCUWG
bOElGIkEbJ/6RwH6DVBrFfhagxumhphuVM/sBNx9j/zbzcAus/dYJa60ioXVaWWi
Xh7YeGIhe/xEBTGZmDlVZcDKopajt9dWhUyVYGuyzGOYbYefceiSORc7Emwca8w9
f5VPfyT/Gy01uswRdWoh7KgwjQ4pFsXJ3DwDejOKoSVPYkIih5bw0QMvdxjBFXFU
fc4BoMIc1Ddfo2ZPdq14BnOM43zOaNHSXvbWo7J/CBHoGF21FovTtNbm2JAxwy4A
2VgW3eR+b6ZMOni5S7lMQ6KIbjxZRkWqmFxnQvJSWJEoxbrMF76swA/3oXIFBoI3
3vv4I3+IZVHamS2XK2DS3IwPJBhVYmOnoxhiHafadgk0mn65QRrYSnZa8qDgT3uO
EE68qld1Tkz8VylikozInP2qkDbB5pFTAX63GWh/HILejwSwGoYk8QZhylhELA7Y
nvUeP4yzdaq2C6ZPJ2l85BpDoaBEEuDtjzxv5Rpuq0m9LaDmsGDvwzODk3pR3rle
TSBidzsK4J79HX9fkez2egvr5+AKIo+WOrhpYJEEf9pu6TC5fs6QpNIIAkoAhVvv
iJ360mcMXqiRYeZsCVC8/rcklEkuz8FB7mrPvBwadueClEgxOq04mceacgtIVwWq
igWismDxNtiktnGaqedNSEfnkzXUzOawU/6e6xxHdos0ZLHYdf1Met8bJsmCASJH
VFf7ulfhfmNyYETP/k625nkcUqjee1IluVSxgr98bPvNTTbZL2tvK742cxi1+MLk
Y4AWm0OBMuVW9q7m5kxTpdcjz0hWWM2BkFSIHitfw4WfuldTIfa962akh051aypr
WdjavBLHJWZxjLJ6h5XPdP7Wd6h7V1ILHkXbi9RrWSnWmIBnjRWhO28DGyLNlyCj
s8xn8ZH6NczjAfeN7zQ9qcSiO1T7DMmSTnZOazJrfki9bwenIS8rkdCCt0V7iOIZ
l2z5rqYlzH2qhnCXLS071YRL0riCPeo/G/8Nhs6+2p/a5dnCV+cZqGKlSsRoOwtx
abXWO7BcypLXIwHhQ8egIQ+AWJ+10ScG/FXq+8GakGTSrceI6UEaUf5OGCCuc3IJ
M51o8m0lAkSIhn0BByUHX2zAcF3R/UZIsTUXtuAG2hCHhYR1IBOygWuWFWbbU1yU
VoMe0bmUcvsOijqOrIK50Gm0ky/0BUHCWtGAW6Uc9K0xB6YoZvoDEi6N+HCLWlQr
udz3H0j6oZMjFdhNTL3m2dUwA/f7ssu9UDATziRfJvYLZx9PvFMFd2LuUlGKCmy9
DFj03xo1vHCY2HsnGdWai59ZYshjBDhVsGhAuBbDu9EbABrPnKU9fjAdL8m+GYAe
6kBtehYk6W/HOiQ8CUIGnXHt8+ht22RrTk3W69opyi7y6gS8yL3kHDlil010G+8E
Pzpw7GFoSWaB2s7Y5hbkqCXdMjvVicKyBLZHu7nLUnthqavgr2OnIj5kNDMHYeAI
/KEtPQoX5AWcCSR4j3r8RUPhXYVJhULK3IVFr83yPbnAQAbhL7RFh5ffy8HcT1Fb
5UHUsW6TSVFhqvXE3dEairvQzkGrEScn+4cmpsxEgmpdgo513aSXgj37T4wWHEaN
Fg2S9lkBKPgNmEbIeQxbmKsRr6lFGoFmBDER5nETrgATqWCTgNG/e93W36DxGdpC
/uoH1HErjEx905YRmN59rcOBmBaClHw4P8SiH/7CC6TSPt88OxGNcTrRS/qBbBar
LLpafoBhml6cYfkvZFq6/iV7bUUxpQEKjldAEVIzGqdmg/sXvWbyaats+h79kKbL
jO5QFfr4RTFKWWHDH2PI3cYjzVGKfv6NXZBl3iWvX99yaGSUfOi+OOT645rlul7N
eBZuEsQjEo1L5jEybwcngdXVyCUIJwul68tMtJqyADEOfQWXeBDJT+V//pjN1TDO
/0UoVKAl6mcPAaVq5GIODPoHFwBYOm6gNUDGtzAFkSUGcP5W3VYKiEGFfsF0NfNC
TxeWxysLflzfdbbDvaDq3448VRa8IyK2YiaNORVM3PEDDYic3Xu41QxhM+Xx7ru6
dSGiOtk7mEbW2AC4hD6UcKfiq6O0CTlneJHQKkmydcRv5VlfaRh+blB3r9rE8DUs
cfV94NuZXR2anRCy6euq7zMcJg/Fo806FkDvIa8boJWNs5m21qVnE/52GLixHaYd
Rs6xr6OoaVtBiyAm9vTVqB0NIzn6viVEGkSWG5HUeeIYkvi5AkoG5SFDvBCyHXTj
N6jdMWs3KawQzPUH1OafApDe/5U6ex1nQ6R6LCEUmOSOAIJGjwu2C+AfKSEBBbDb
sKXTS6JxuezqjIA+DCgxNH3pv60nRHL4Xoy6xNci5b+nyWJVSjNlOyn3CI+zFlWN
TwGT+l4C4BM5+kInav9hgBbG6g1F+Z+MMMK6aFCqmDGOS4aVyzzf8QEYx3cbHDqy
t/xbC2SjS/ISTBr3sAEQlGJgLg7gE6fdLm5MqTUyyDAfd/5MbRUeM3KLxc78Zv38
bH4c6MwJukwXIl3AGkHIliP2IlV59N6V3k22qvWT3uSFJqeE4uCu3p3RuFCVd5U/
+y1/uPWGjb3HWHgbz2vJ95epuvpbM907lkUa5LVuv4/6zxwuZ1QXR7+hIU/SPYkX
ODggLBxU6iRonM3l+3lADq3L6g8Doh3XsVMGAc20FKUPb2SMpYxoDhF7GqFt+uiG
A+ifvJ+dowJ2+oYjUh9npm+FiggavDHMJiBB7ibqyOlP5MI/l91NuXjlEqCdh7Nx
EG/v82k0/qcjVjpp+XLdiIZVqWgennLpmQZxUMb9L53bd/46YXwSCGTn/Vgtlwjd
TsPK800v/itfkrZ8WaPmeK4Hacb/AowVMf0NXFHjRcqIMppityCG56U4aIewXtHU
3HWVrFVTLkFX6usChOMu4BsNtbPueVvkMnU5HyBe382FYrPXEBDewSSGD9gst9t+
8DAtoreyeGjCxZxlXcMOqmsPPLa1cw2v/jUKl+yXxmR3xfWnMHGqXSH2iyZsxIpD
URivyOYdG87HDqYRzAPOaaz+0xDnfrrDVeqdAMMuvGzB0CJ1uNQQIgK7WsLdI148
Lgb/r4DHU2aekldAAOg5FVUJwIsxsKbga8vQH9rg3vs8x+AjaX/C76NFlJTZN5g0
g8HYyI3/20eLyacrnJxKr+ZuQjZzXs9XAAhlJaPOZOUyLyCDCj6R82fYul7driBg
2ulRIl3dnMfirazo6GXsqhNdpRDCuqfXvMJU5g0ZM+pHZ9j8e1ztxYIr9i7n2C0q
n2s3cs4sTNhtU4S8URrfRvJGgG2sUx6MBWhaD9BohIeP4v3HCr2jObylRDDJ5r7m
tomex+GLNMTyf1IbewNIasCdEjmNZsbdn2YQidFt117XFQ9LpWQ+vR4+YYshVk1j
xzIBQ5deoiLWuDvXNTAqowgCSmn0I2LsPwM8HParnoSpy1zqOcV7mJuQDzg+14+y
hz6q3jsfBsX6B9Xksmr6DvLEXnj2is19QcaCXR1Y3aLPfZbdB7/LN3D5qcJURo+V
AcfI55L6PbV+6iFBASpZnt2tj4dNtDT54sJ9dHvC8YidY8gUn8RFJy7HCANNNFrp
cUcO2tCotMMOQLfji0xzBj8UGXvdVlL6XkpbwsGE72+9xCvK0CdphIV3VNS2d1vV
TZrztaYN0XxXbEv4VCucU/LntRrCOt+URtXlyMXP647JFg3uEpFsDbHHPUH01Tno
s8lxyMli/U80voMK2klo7XYukC6r/Rbx4ZZsCUNod9CPvr2Ztd1/MtCRMgkQ1X6E
B9jAr8082tngmDUdPbCjDMTTHPzni/SXwOG8SbWYXBJOk9ycQf06Yt0v2WDbGh79
J0uLlWXqbhpCXRO7u3naOMXCvyNh6Ml8zhwjXD1GsPlNdnN83t8/ISIvnbe/ia1P
7XkGTUWKnGraL4HsCnUFwsy/glehnykJVvgKtybPVd9RZrPMMFHeyO39zYnG/4pR
xz9TldDOuxe3mbFuKpxZ6pgB/qf0M6qNMEEFF/jKWXrezlqpe66tWcvJhUJIP5wc
dfQ8dqOW2UBf+HyYF7LQYuPn/uKHCF2iJr/uxmGVc7inOBS1glLNSJE7umFQSsgY
qUC/9qidfv7sVaRLiNNt7no3JFoMtErSv1OBFoTOwxxz0jQS50TyRJpZC+ODOFvO
woQzV7pXvXvxSg+UIqESTJdNRCNFfkq46jF/Bp1Ddra09tN0XSH8YMRsMA0S17R8
a+9L9AGTtyEvCYDHoBiK03rRUG4NHfEaUfKVNLXw8k/zrHQbBlhuM5MWDiSfGPSo
wzubDOeSEeocPKIvRf9ruXaZzJho50D5sF0HP6HVbG+9RLLdXPYXJE8wman27NG8
uFB12ZsKFTePxreuJdheX3QbFkOB2kh8mrTEeg5Z9HHoU6qBv7XuPBVihP2Y+qaD
Z25vFuOHDqY98/7clsrujaXz0xV3hIQGs3e/QWN/wRBR7QTX8P5JVZCEHzLQ9g5y
ye++AFMxidvDD8m2nQlwfUVYx58X+GeBcr/XjYRbL1kDYD9FLXiyRouvP1DUz8cP
L35eEMxh+BYU0zRGvMqZR6STS+lXxhpggvhYIZ0gzb/pgyDcOI/hM2XPAAw8JFOs
kabVqGJOBQ0ZqRscaLG4/bGAKN4uuykXI7WU0fBvLOBRKcUQeC8DpMeDi8EHy7mh
ABuQIOIzlFCmuEsl+isG8a67it+GPh4ywPJK9CSel4zfJOoPn7q7i1ktopHAR12W
mX/KnyHXWzQD38jkAAy3S5v5WbxmiWo50GXsopFJA1QYtu5idPkpOBsFvr8XJs/4
Ggio4nCisYBns21U83CH2Q6XxZ2nxfbQ3NIbvNJ8TlrZbOaFQixqlfkR3wQ5leEA
iMLsHty7pNiCSQ7GWvQ2Rf2KD37DoYvRgKVYEFMNTu7bNJ1BI8/anT8HhZu2gxps
30zKMcTrI5isWgX3AW/NQyZmWQo/AvkDUOC3PK72pic1ha9Zona47c5gWH7WX0wN
tKJXZ2IV8RS31Fk+DHVdWFz7ha46sN6evEk8Z3Ejr7+2dBJITJfz4wgakYrm02yC
QGyw+aVoCVTAPuaLW9Hqgh7rglssI/mFxTzFajkCaUO4vxhiqwe6TfYW3tueNHLr
9RIUVCsEs9DYOkWWyYkRbhbpRTclzARy+Z34NQXqzJ0OcdcOnBhlLvq6cKwxUJRB
oTbjfsQ9Lyr1k/m7eL4VyJY5z/LzEmMjZ3ta9bFFrBd2ihORCsIHICVbu3hjLped
fwlaJeGOAecKsbUZFyhsHy0Dx0bimBpJWObw9kql9RxyGvAMUXaoaV6OL6ZsuItB
rb5AqhzFiCxzzBhmnwwyi7ATfKlNhKe9KhKGnDl0B9kXEXj4jZjur4oACHj3YSqv
VLeg0q5OXEqP4Zo8JHbgFS/AWaErqkvRgDWyipy3/6OdVZMios0MzQ3vs7KonrPz
rAmsZjhtYuEK5fd3++mR88fY+YkZymb93nhioofYvezg4UwJaLtFW+hFTTNPLhGp
jZ7rk6+yCd2VzyeTBjpEuA6uiFD30nuKLNx6nxnbjOKxxbJHfjwPdZSGTLt2hySc
/ijuwm3jTBniv12NXlS+y9l2Cuh/s0S2oYjwsYV/EisFIqUvfYq2x9jLnbC2nbUF
ivnY5VyjLcCB3iqmXvl1PF2yOLxvdy6dJijkFFooF+mhKppggIQmbd6TeGKLiJE7
a4l4UyRKm7OQROXEdMFUksQxJUSxnEFF3fzm38Ivc/UtJqM0G2A6Unsmht/3l97y
4pozrSLCTID15D9wCAREyJDk0WMsOvrrWSz5WyiTwLDhypAVt+1mci6TvP57XvtF
ddodDJUqkfSi06lRu4FqrAHR31uoHiCOUMGCCpXQQDXy6V2B4o1W1I+wDWX/DeoY
IKa6ZZzrDMpgco6KHm07tq1hKriPK5Kyb53ZAoW3/eGVZu4wGEeVKi1bI/sZEu5c
8PAF/fvqB5Dxa2gwJeAj6CfQIWZ5msfbuYj1OF0XDMMNQAmfoFcXQqrGLCyUDTFv
mPYhvYbyhRsQ9CjJCpfCsUsOgQqbzrIIlhT4Pm/jMuymf7C78cE3MaeGK7uBpg+u
Z0XBx9w6uecjhJvsRoTwMFYvAv3mmnRlATG5A/75819Ueg2YWTn6Pg13sf5zRpL7
Z2wjy6irEHFkGrumVKpw52v6N9RApM61SN3hfDBx0OfQWJh/uD7spf+npRasSJNi
CCxFJKt+5YG9wyC4x2EQAN9j25PjitAi3T8AoapcSxVQvAOuNvX/+dbgYP9fW88A
2ZMXTKf9p582wIryt9Bhd7jJAQJYGiTYF8QnP2DWQ5wvSv9avewbARTshLEIhUJr
LuDntWiAOj9Bn+hkOxhukYrUV+khsdTUqfpQCN9yfztI0bMNrEXs1z6h+d/kcxeW
FIf+SOFu9bIiuhWKEQqGo7c9MG/X5Dn+KTijupltpVs8E5ncd9vjZXlVc6gX7Yol
IAIpjT3sW0m5hZV2uPVQK37DSf5tNj0z675A8xWh7HGNzudzchyIyCllDKVQtZMc
73C8Cga5/2PvgRDjWmnlyx9DW5QpElOcY+LqgmMveA6NXRK1F0GX4KVkNkmbqxG1
s5223UEoSEnhpxgxa+ZOVXepmGLlgo34OvNINLd5+mtzoMM0TSMWTE/iVdJ0ksBl
m3uKOxPy3aetxFqt1x8GroslntwULN86i9byJHTfnisWMGmraTsBRkMoOauRmey3
7gdA6GbvA9IAHODYjBqogt1/6YOGWNpIQRTCcirXQTMUEOlHWYZv76e6YJaMXmWO
2ryjrgvvGp1lUap0MsOT6pyrmx5tnMjoiVnAKNzeaV5kWPQ6xzqlwYDBYzIcnUek
pPWV4Y82+gMlbXQ6LhpFCYDGp6AFu+xSB9AM25PrPwXWuK+2przsgssPnnVOEG+R
RcaqApU6tYNxTfd51vcMnUUMG0ic0SGGgNn2bYVWVQDiVAUhsEp/B5k8xan2n/6q
MIvkxvdEVorxOCg6bNhsJRSAOMi6DqhuyAp9OGUaf5BxR1laKSzZ+Aj7jTRfPlEZ
P4uX/axz5j36j6ABXEfZJHl9eOHZc8KfKWdb1H82DR3en3TgVnBS343M6+qSA5I5
58yZk1WVj1SElO6tRnYiu2vX3JyyWgpyAD41ej4S6dkarKjAaD9TFgEe6calkPRF
OKYMplVDq3cmoNFn5K3BKKmdLoxX7CeTuUPeH9V9xYJ8XxZRT33nTrVbBzaMA762
6W9HyJ7k29UQUVpnmTNmxaf8Jr+PbWBtIXC9d2vmuuMpu6iTDG8W6JCXnBarvUBF
CrPwGCu4eoRVOxh5zK6xPo9B04KtuzsIAnDZAldmid8UdKxFfOlj5BF3Z5nJYEjT
daUDOFWCrhRpycm72czCncm2vMjIIeA507Gi1R1pQ0T6fLhxzUwRp40ZEAsoNczw
WtePlJNJpm5hS3HMhGd5oVMChzoSzz57hIGnnPc5LPfOb2LP0aCmVCJxO2oF621z
Cpk8Fl8WFnPW6J01NuQDndh+lblG5lsXha+s5TgWTzCxwW8HdhJUI3qt3iNfUjaz
prRlazapgOYUGlBgrBlglTZB2nesFzeGvOfVje/7uxO208FvRzglwNDzN6AkZDbu
U5X1CcVfM95qmjILSUKVt32jnOYZrjSf+xa0puZqrSAO2cjhG7T6WVFUYFIQTmWd
hVLJHfTWgnWlTcngJpVVgVqPktzx3Fee3JtJtfRzRvaJKOVKQcOKSOd7XLi9/dtN
7OGt999Dwg6bv7LJP2fii5f4SL06tv060HkFf2qRnfph54quOf9EJJvo5lg21Inh
Pp+yCDYejjI6hcvvbyjhkm3/YYUzXU7twu7WjVtaaoEJwa/WaV14pNRE9D3x55ot
SLDnnUuhzbTsTNON+eSh6kq2NXhp6XsJe2uns2IYK17RUXb+rhEZ/gPiPM7/nwGL
kttq3eXDX5/anI9OZIxd49YQnnrDEdHRRjnXdScEyLSsp8q7xG8kNYhbyiLWIzVd
7m/IjVgqzvgtAiOfLQSW+215KIXM5ojSWnunbGpOpw262p8yYo/jz6E6jnPvgDDU
/jLqNqxwjn6spHlEaY5J/m0KIENkKMQcSrExaNz7/08CC94LpJceeJamBS4HMxnh
S60jnWinVunVSspt4TnzUXwIQ2dqNpoX6O2+AW91xxM5Ghq/R2UJLlEpowvrrRnn
U6lYbcNNS93oKhdEUTI4nknCJAV5UbjE0Gs9qp3WXYpeyTbHZZXHViRusNEPVBdm
5DU2A2p9oalOuzD1CaqmYtGZ7edtgpzw6qUmomDOGMms/QrLQrGeozupmdDkEX6j
MnZGBsZgwD3EW04CG+UOw9Ghd6RpxfAe/GxunUfLNVp6OVMp1/1apCrsa4O4VEz/
weE4F5q+KrH/ka+SFQ6Djhd8/B/Rc8C/KqbTmzqTKEoU7yxEGRCaZYQiIYQ7CIcZ
OospBwuQzYNUmd8Yw9QMgBxaP0MgCtzo1Q0eQGRn4HQA0Us1sp0d5jIksSpzHKMQ
sVHZI9Xq8ZbJrdJys7MQy/a/kTWLagYLpdSGgl3GNOeYv/SXN3RS3bbzDTFaBjoA
Ps6mPIwUp6EBzOuIbskC7AUie+cYAba39qnrVGLDRPIbO8JZSCGf/+iI/h50R3LF
m9WlbRmN/Zwz3dbkM9N/dn+jz0S8k61VglNLE1o+U5oI9n9SMc/4Fry/IQKIT6jN
tRNbLTOvgt23pPlzBomyNsO3nvHOmrhJ8D3+rHQGoAihsul4eUY1Fc9+RkEIjOBi
QvXQvWorkDhzL+S5CalbglPzcDfzaL9WYFP4IvhsIVX7R1+Wo5aLT2KKoccbQ4qw
cPIhexowg8W36hlzFWa9WXqm+tHrmqQAsCv99fBvcs8spY2ucNK0aiAyC6atLQOg
G1Jn2KZaBWmRcAwHSDjoiXzgUvfgO0px38XRJrVn2PXDMFX2wU1JOVp+Uf/vZyuq
Df5LGdW5V5wVLDVDNWN6e60CCucv04sbfzCb1vwHY27KpFzr4egHfIUD//k0Qqaf
psc3TggxOdqPhsaky1Fv5WkIcvhkq164rbaMZDW2SnP4QV5MtKXDbVOPNH1eu9gP
uN8CoUQVneQ9ZKl/lF8PyQouyVn7CvIn0oTTZ7sZ1UR47J5gFhcQmWy1DJzOmIZa
kNh0thFrWarrnwDD3eXZL4gWHiG+IgymZ03GoiQ6gOCnSGGlqduC26Ca2Js/vupr
n9xdlBs3S+/Ch3c1P7i7OM+iYFeJvCexUASbr+W2x0/GROOXCGbCVQnZNBc+Imhv
QCc1j4/55H4dhgioLtXcu09YvkqnN2xZpDW1pr78VI230q/ezPo2yQfLRviPeRsA
U7UgRmCMDvccGBetRKDgC4+H60YYGyoKuY/30q3P0XUGD1QBAbpvXpyZeZo2ykQR
jSoA1ND1fPOlEi+hMaAOZT43efs3vchGJScLf7xH3X2VO9z0dUN/uZuP7YNjf4qS
xSB6dJL9qU2Jl1cztLC6rZzS6TbeTOM42xj8FGDrODV6FqN4UXHv61dv/lEfN26u
T7FZOaCtXaPC0FYfmLaXA0/VIKEPeyi/q9quetG1SBgKFd8cW7DJKb6Mdm+JDnlj
JKoR7OhSmJSFvC8vTLqEafrhRwPeESgiRuVy4kMOMYSxoY9hhLcFIDfvfquiohGw
TJnfpUoyysD29NxbGGZAJsC0IuG3i/X6METkPqanpbFL+lwcnoat10RlKV5hfXL/
u6FyfQdoNAAhubMUrjLHcZn1y45XKm3pXdSkQ40Y77Fue6nvPdo1iHYPdJp87YWD
L2oTxZ3UELYmlG+9nh6v0/tuJuwxa5nX0v9whwGUexpjY84d4OszY5KmYFh47dSc
3QR0GAo7xOxc0hhz8e0uT+LO1CjOnamBPV8EXMTprmre4k5/f+/omwl3LjPx3rkK
dAYQe5M4+rDXShi92ZvR47N+O2U327o18DToxzXXZhJiMcJKef0ei65+Lt680uOO
ktz+Oj0+M1Y33Slu8SQsFS8UFGtJNaHWBlB6OC0yqCxAnjAkKy0g0g01FUU0eNJ0
w4xdqlWY8ewdV850MSn56P72tvFTx+0hCuP/CjUrWjmpjo8BR1B0P5zmRewy3pb1
zombXWUTWrPwocnI84UQcVQn80b0yRTLrY4CYDkzFnbSqcs/RHmZGjCNJ4rl0RBJ
Hucs98jFX4fhjgxc91v0OBVhVT0ZCD0TCHM27FDaVs+Jr3FfUUUkPGqFkXrc08jb
jUoNPhwrjBQsyEpREoG5GyBdl2x1AOHOsxGeiP/9CEwMhBT+CIX0vOINCfVe4gcB
1Po/AaPgHvuQGNLftaTIqt/GTWgldb7NYdjS8SmAkvxMhmCHCozVs/UbA3+TCjTV
o0lA9ny/BfNZnW/wxsjkkd0EdSDozy0B+yvkk1wlJF1p0P9bjxfAUi1A0VVNDlC8
xw47lKeBisxmJgEjpC97Q1ZtDIKavpAt99+ew8LayBGEYgWjN2d71R7EEWnI2B7B
lZjihozUUeps5GOp8SdLxnJ+zhB6PMMTNFR7eqiYrLOri7xvSxMqDvZ6S08+FNwQ
BPZvBvmrs4OZ+7ejL9IK9NSwBixLeUGIbreZr1mPr7a8fuBxsej692TDRQWhYWPr
Tv0K7Y+pG5XxMeV6KHUVOyStvgFtASURBKmbC+Zi9Oe45B7au3WJxVchLR2Howym
teaqTKE8LP2g2erpm3uU8XcnTjzKIFoHtVj+E3EnwWyIg3vvSO89Mv+dYoFCo7LE
yspsw3Ez3f6pM8+eoUVtCzEiTO1G5e+eHAIKRpYl4WQ3ki9rT/oVAFc+00+58U/G
GLwBESzzxC3WRxt0c2k8hAqhgFVFzAXd9CV0S8uGp3cA7ul0uAUSlakN7qYPnGz6
ti6SZcRMhIiPm3G0ILr024C+ykBJrnjv4GgXsqT1v6A4f1AKuhduo9PyfyvpTiPZ
MfrnaTbdP80+tHhiO1qiHW1FA/zTBb5B7g5XsISg9AVW+H0CofvNAZcuNptdH/La
uBJ4gXMzIdh/5BNxTP6YivJZDowfZgP1DzRWUsQjPCMWsdAUq22vAvOZL2y/d8kJ
uFGLhFwH+fASWZFmO1cbcIHzpSvrx+WYsmtqPQknZY24OUDUw0sTvPfsAhnP+RsO
vb2+peCx1NjVuM1jOKcMR1oCfKfzFk1Mivy9n5WA8zzGq9u1hH4wCeoi5vNe3C1f
VzFOjr+yz0uApeJg4EL4GfzJQ0sUjr478cotRoeLddv7Eeb6Opf3QJfMJp0b12Uj
w5p2RDHL4XpSVnBJJht2DsWCX2khh1UetgbepL+a/IhDsjEkskSk979OuP+f1/9y
kJYTGo7gNUoqcCdXXIwYw8mnxoIxsM90f7MKv4Mv39swlmss1S5+kn3AH0BTtywF
98QquvvdgEf4FhgqRtya7DfFbMEzklOnuFchawLOzkcd3L6zPqWUpaVVBHm7p2Yg
/hnnx200I+NwEnMnAsn3G0E3zJV044LjDLpedJKAMi9bKRhH4cEkXGeElEFd2O3A
oCd9PbvwR84us2qM65ZBaiBbFeGkJP1d8dfDhjuN3r/gBtqq6SSwM0DIQuNyOU/G
Ev6t2tImq/WNnpCA+MWloiV6rxfURH4USg5iukqdvGB4bhMMH2+K2p0FYDJxoC9o
gYFiCHU+ieNe3cLCdBTmiXtGmIjjzlkAHU1eJXqpikcSTEh7UcLp6R9lVe2NGy1C
QBihDQ/wZHURLm9ByymVLVTstnfjh+lZgzGzxh+lpvrGuy0SVZWPZ4AQ3YnDurUI
YguAxTDukFSuDcQGBo7CSCU36lCLNHZypsU/1VXZRH732pBzTrey6CxDKa7WvJXK
7Rs7B0TxZDoJT8Wj+ntKDGLPt15R6bs0Xv3gI5On43RuYVtcmkuydiittqCMcSKP
yABRHdTQkuxtUM5py/k/BwpKI12Y28+iJX6ihPZgvQdZcx1NGZhyJaF9rcluoXnh
DYPg2vGTRGtzZ1ktyrvwHSd7JlDUwS8ItarNosiABJQSJSc5GVMB3rwlZNynkDJy
J1pqTlQ08sP1mBWY2lDSKN1TG/NziIo9xp7b7Q2Pq8MvEYuRhwujPBSk1FN3jmWB
roICl1aCW7/V13eZg3dIBrndMRiH8Iz5CUZwo+vB9k0xMw7pRiBCJ87vwSiWONDf
hCr+TKX3pa0eupyt3Sz25IODfB8qnFZKd6LOTPsZ5VKcBizcuoj6DvKOw/8BL9EA
ngx3uFLj8Zuji2hrnRAMTNvfqjK5FhZXrVNRnnKGWwSUYllo348Pc7IwV1lpTfEv
hChC2TCzoUNHOygZQ2135a0bU7lKsDQI4sAqbiWtezWRKhwdDh88z8kOAuIbWpK+
ffM5NNaqYEHX7BDsqD7JDZQz8SirtLd1qZs1cONLrnlJcs9rKQGVVNV3FNfPYZyn
5Vh04W1fkTS4cqMTKeIJfE+8XY4bGl09fjKmsjV577ezHYaHM+ByT0NFcGIkmsmv
jFGYat8XKCqOPGzrmh1JRkoTi86q3qFPiLIW49Y7FOuE9IYILVtIZqAVbWq1Al5l
K197H3LX6FgyZIvxBEza+fM0JGmNUMtGcMQotG0kYPn+udgT4sxvBNjFp18WkADI
iP5DwKIb8OXB4I+T0oa+Yt/C+dcKcGsh0+TST/ElEcGZcRl0YgiOEE4SK55idIis
gd0UD/qdEcZ3XEbbi4sJL4oV5mM6Qzv5Cg1v/tvTbrmUSAUtI3aESNzVQZeAxNXD
BfRy4mAvW2UFg5n8Fpny4Nc0tSn1UdjAryiA5mIl8cj++RmwjT61AkHQaqkkRTbJ
JADq1B/fSqKOtVv8b70SfjgkctN7a20W5Pr3/x5M2sTbMESLMVjr7VGZx5t9hX6L
hm6Q+WZu7NX0gA8dze7b/9V7blNjAWrfKBghAbSm76TxurRI5e4e8FCbGo+lAwrL
LcSCmcUap169zNNawqNjUL14lBbOBIVwP4mjYXNttWs462Yc4mREkcf2i7oj/89Z
g31OPXuTK0FOWxDYrVWx9d/S/4mY1l1+ungYqbw88NMuQk01GTmIA7v+vSkPBJbZ
b2rxU9JxZRgl6NZJHj9v2Ipbwc2rcA2rYCdKrBqHK48rDwN9KQq2pKXnV8HznXil
fnGTU4GukiDX1PxBTJvYbzePsF9oeit8H5oh1d8TvFiTsOk/SvbaJy8cgoExi0m/
Q9Z0tvUgd/2v6ddbbUo+CQJngg3i9h1Xvs7/ylHFLEUG8wxO2+bUql3nyxFEMM56
MvLb4oSg/hdpoxDGo+uKUKS8iebFGYiWCa3YNevpn4QoWEqgKtm4WbncpRyBV3Op
WPE5jLerM8VCbCleaU8bZwt/ATlQPig6Q0IsivS0BEk/bWZuchEZPy931I1TmdC7
i29vtOEQoCY/WVhzZGm/MKPEj8hkIaU/Q+Na2XaBGrOApCsbLUk1oMZybsQadmxQ
qIh1fPSLQxL6pEsbO8aCagXucMrsSjn4Vo19wYmDXeLm5cNxP0MvojjAViahQslf
b3GL/9hMMROxS0lx2DfWTv6tyQOJeWWUcoUzberhbVMnpVgr0BcUXLngIdPDOb+J
2OTpS5/HhNFzbTkCWGRNZFs/u/HHADllcRLDXTMeDSp16s9e/1DZEmBBp4iAKFVJ
mp0hm0rUhFhGJskQlJ34nGh4pswzHGsMCjmfDczjXGEFUcwBdhVdivPdVddT0Unt
j72HztmlRUlx4sOQJo3gAiTYi021HsjvAApYPPK4U2JJsBWE+JIKstjbg3DaMj/1
DvuF3OH8vdcq8YJh7xUgqHDRz5E7LjMsC5CM+4oip8/8nxwSoqQufFvcuNrIUyVv
9ZLuRu8Ei6eZnUEWJ/7MfaxBZb+aRMIcCGiYKiA6Mg/LSqfLJsK6r8odmOktB80Z
KfgxsFJ69pw8Yr17fzjoeLzApkxlOID9UWmuiqPIUipK6sQnwZMQbjZZSkYs4Bih
q5Es8k5Dn0LdlWEHwiaPX8efxcx9/VnSop5TABTh2KAni87k7vC7XzlewFY8cmPa
4Hosn3U1LmP8DeZzragdNGO7668PcgSHnn49emV0pxwA4rnd5fyMJIYJd5t70Ms1
LZFvz7EDSPPFpzWaIIZaw9VChT9KRWiKZsJz1Lqfl4XtI33N3i5x9+EnfWgjccF1
0PLnkXdg1jX7/oaw5+SSJl3jRESuEXCNOPvjM3zZ1qW1EYpWYUYA44YUatO1HHt7
/6f7UPy+HXzxNMdU7zcnt2uFkby3o0lceU5szX84SuYPZjJNeP2LsQTsiSRxEJsa
G5MDUFAxaniqUlEuvbd5SzTDPb/5P5w+07AewjBwr2mfjvHuJvo4NxZQqAtQK3gz
FHy8pTc09RYR8GXkzl3MD47UNDgFmN5qoStcomFYCGCNIwx90/cCJYyLiW+17bDC
ZbGG5iqQBDDpqH5bFdDQgVRSe081Vp2Cc2mz0tesyHW1O1Z3xQpGeLXjMIjO0pXf
mS27ebk8+t+dWjqcu9MtDAfS8pc/W7ykTsmbXbCiPIctgWrk8o1rfGFFYf/wavUd
whbUeLg7VTMNU7sRSOxWWSWjU9EWUop/fKmDutPWiomfq7EB2uzMxKvoSPr9MW8G
J/heVXSdAb27eXrC4KRJDHLrgAVUBUSAhXXPEN5jqJiFMW740POAO9TtxgG17z4+
WtHFCZCd96NbZpwRBlNi3nID2sz9tpGAm+OreOtFLgsBt46/1AHegeqH9FMfmqO7
AwJuErNNm09NZTQDNlgIQNZYnSiIDPO+Vs23YUPBlWof3UNRsO4BqecN2Yr3ylJd
Y669GEPXHSgC5/ViUww+SzXS44I2/e7KjgISon1bcxa69kyPCIn0gvP1F0zeptk9
bNfmCXm0YA7qckqp8Vjr8jk6tjaAvW7Gjs+T6/6nrANotd/Njiq2A8tTimm6h7X3
VbJCins8eu9ADFFKWL73F4mD96E68EAt10OVvo7QDNDlzP9gscWikNjUGI2WLIV7
pUHFulBFhcyPPj6IZm0osTCdOoF8CHmK4Tr4CG1f4FRQ9AQN2yXHYIGWPRgVSr7r
vR4frvZsz85EpxntgBEshW2pInIuGMQW5LqTs07uPxFMPFvyPKXsOROkeMt8M21D
6K/jxKB0L1E/H1fiBxM+DPh3/y64BjkEIX/CH3togCxrMqdoyZOCKrF35EpI/RNS
N34+Qee/x4/YcpD2Qtq4Gc+Nkh7qKqye08I87T3jFfLQmP16nORFUl7KoG0Qqt/f
OVaZ/AtJRXpu9vqFucwDcMGwZxr3iJgxqfH9ONaICdieHyRgNiVWRz7kJX7LL17H
FIGlI2TaubCOQGby9CvkE1WmifiTdNuutK7x65KzOi4rHj78jtTJcVli5jA/RmNC
Dv3ytfMdUOK9AEQh0rTZM8Q2Er7orFVXQxEKGXh4eloWBItbssMLHchoqCrqBbYV
/8nwr5AxY0LGUgu0+sHvJXBDAgQhkDIuNZ3ygx6ETrVT2hPsiJxrB6ZwanriB22K
K01u6WHBUquRMUJc+6lwuYoGfjtEnJB96392vvsZMlRY2SvV7n04Wy1Ttx2Q2U2G
qxEs3QbK7IO8QeNolxsy4L4pUqDeo+NIDn0iFRFMyPNEDSlrooK5kRZI+UM7bUge
ihjeITcYaqdJGDKEhjn2T88avxC9sATAGlE8Ljq7miP5VYoupLoz1xBDjGC5VSBJ
u+pWUyauI9+rr0wYHZszxBnRSD2jYMBp7FddvET6zppSnjTXqzrDGyu5NiZC+ofy
/4DciK8dld2txorG6Ca8Dkl0jBc4f7vLYJE3lGpsnTE3l47Ok5wfeQ5FpFuNLnBa
65ZJKBmbOrKwFbvRdpdj8n6lsyseMSbPwh2Vg9fvJgfu5etEllOH9B82coL0uJ8m
BRET1HIg7rzAEZtAGIRQB9UwSu9N0NaNDF8wB5URHBy1BLvHe63ljviruUgzv8ak
TfvVlKF9QaTC99DSuoZ8HWmRuyJ5+cfQOJoikeiuGsC3P68BT3JwleMiON3sqEZc
d4HDvzDLLHYplCrcS6ng96ZJK81fBwU8/+vdcMJAV+I7w+hG6mtaMDEEWb8INERE
kQnxjIRVJuam3hHuI83LJUmRCXXB1zFWvh48M26RpoT1s1Ny/mpmRuiVTL5EPcjw
L26lkPkk/TrAwOPFGQRtIDO4tpwWHoN6X3olZhbZT/GAnWD1/B08EUGVX9JfKxcu
RWQ76v/neB9670R7u4r1BApL2USPKftOEwcXMtemDcLff8PX4xvleXM0Go0JW6MZ
2SxsGnUoU+yLtfJ/cLZEqmusNz/32d5dJ0A7Fz2EJsbslIxJ4W/1G3QabGO13+16
XmS0B6HalljCmUEznEFDKvHDSoBf+N0nkKoDUwt+lyNEkqT7b8z7WMjndRlQ3Xwe
SxHEA4c5TqAGCJDJvAtjNdNrcBT7iuut9EAO/lI55iCEsXJ4TH7ZZbItUkqe5pJx
My90B1pZJ6EP7tZ03eY593oL66EA1fvcrtFLusx53FkVNBqbWD4hRxdnjVMJmR3T
dWn+BFzyO/79ivR4ZRPSMP8nc2Xm7GdaaKQXqjFH/4Z4sRY3SKF6KQ5DkB0Kqlgo
1F5VpSqA2NS66bPf+/W7Zqix1IHMwcW/ZqnCUFxeYgabEqUlHOsHZn8oamrbSHBm
Eu09RuSzuenB+NnyRtzCM59uFPpnkxDIbIxiGqT5AT5i2M6O08biLANvPf6vMm5u
k56r4XzCNLEVYBIcIi1jrujs7yL/no5TvBQL2ycvcrMERD+eHmfB+E82cJNDH5op
rXbIBgh7ZscBAKk6xIZs7xhYuzKtUH93LdRV1AXFk6z+StLYmEG/CBD7aLfrkbgF
D6VD5kGgRAhOZtHA4RvVOCHQyfymn3rGDRXsJkmGzPb+tlKYgE+TEGWvYwzYGtLP
pentK4ab2YZBgtt7y98oStue0lRZOJGdAaZpYfiEMSWlydKp0wwQ/aHq5YuFpNjd
BL9JLsyvSUzfqHhg6JgVuF2j+ebnJtbreDJhLOp2v1lVkkq5AvNqNEYtnTiVfEWz
0o27kge1Mo1vE9nJ3Cq6XwqGbOvPtbfnOzLoZYE0dfWf8VOdVNL1OKfonfWllWNM
wZbsokY18S851/56eqtT9CgoKBpdaEIe7y19w5iGNpyXbbTXnGoJ8EhUf2IJ8Yh5
fie7cX5eQmIA3URIurQPjGYFdwVXy3P8laY1RE9m6qcwxLr8wEogEIVJ8RZ9LoFo
MjLvw8i082YYesuBpo40UCqYCNN03rbzR8ghnxYcA+dy7ikMnF5C4ihbInUBqEuP
aE6xWmBM25EUoIoIaYFSIlgVbhQOdWRAadNrf/Rlki1QP7wMARRrym1ztKzPcEgn
DWFLEY03RMsOtgYJh2u9lypFoaMGqvtBwROji82IOTVh7DXmv6whFKeVu+tubaBc
rcgAOHplco9KZwbnz1ExYRaH3ke56GZ2BQbhW8+3vlZrGgZ9dNJOwp6mwcqOIot/
iZEcFiImWWo/7gU5tgong1OZzG01oGmZs/UG3XSVcr3YuTzB6ZRHhcXXd5AmVkY8
hVneb2b3ZBWhpCJRtxuCBP/yWZiOF0OudBTiThvKPgDJqEmRX2ZSfvCqgbKlDjIN
ovs5Iz+KzBCD/4kMGOzGq0B5tJFzlDKaQipYImCEdEMoL5HFSPZgIFMnWInILFJI
p8SF+QYXpuA7CFEAMk+9imfIeXWIpzubRkzorBzHh2Tmr1mAlBxPPvp/1ZiK+FGy
f6cBl+pxKCDJFQA5xMBw09bf873+NCS814BaUUJaUiWQsyB3RBz98WFyAV3lxUgp
1QAD/zGlDnQnwg7tabhJiew6eX6zZb12uSgOD4sRlmzWjyNpO2GuWNzuO6YuRwJ/
6rND+Zd/9Da41AziWK+Ghd71wcUG22z/x7Bn4Eu4BcldFGBCJ6VnQOSzDgFsKN3V
+W+uQIfwgYIUAG6dP8eL3H/JJyBt+DUqd+VxzHMsRgq8tyvYZ+7H3lTg/7bpGPWG
WAu6ggX7DuPC3vRth6lJcOXn1y0CBbLTxDnGDy816TAgf6LE3t6gkB8ltQRe7PEh
RKN8RPilZnpSra9E8PtCeLwrHvXbo7O4nOVzwMwLaImkzgB/sv0PHsbOosXefTNk
6ERfmKq2RVJ4T8cUfMlCuWU+edK4eK3cOvaX8ThiZdw/n5LAByZDtRjIoyAG40nt
OfqD+owXskY9htgBoOqfnUVdtJOrt9iEay2KsqpavFF+ViG467ByZMDUU3n2PhtR
dla2NH8KXJDRuxL7gMG4x0AnOq4ZCBfxegf1JPAUsNmQ+euRvrFeNcO6ILd2Ls29
FPNLNqAYxoqTqho2Yoj4FVuwcH8BF+AJCJKHyZ3wPdJjzlpBt2VDnqbV0Ao7V0qM
AdfmdfUGh6dQ/putNbPW9ISUpeevK7eXnmr1p54s/3YAskbjqF6VHguVx1Sy+c9D
LTtxpOp5nrFfVUh7FtVj1SebAp0OjhcFyH/BX/tkN++2TQBpNfDzQRA5cIyljalc
Br99TsWm5o5oc/0uRVeC3XzSiNgFZIVikFnscDN/Avwu/7Cd9GwBn3m6hwUEtb8D
yMAQFKmJCVQ6sbs628V/r3IGv93A1ZMzhzabmHW3dLYZuFZqcehhMo5F+SsEffYc
u9cP7JXf3DcuE8gVZ6Wzs9kwzsYYvZHOulfZBlTR2a1f19503Nl43GP32v9cXUrM
V9fmrw55V2T82Qo+0k9F/QyGEDMcTZHeeQpOVRl5i0kW/CaqJI5l4OHHWRoKyYHL
lNQqXQGnK0niLQ0SLaCI1sRqLi7PheY3Yhs0EJKXB3B2qdapzYghA+LrLlHPgmKr
tfLzcsjA7krs19lrH18EMMVwOTpplFU9i9VxeErtphLYQpW6Ml5yks8u/TnhTLvR
f2vTu+p5rQVaKwklW4WnF+HYjHsHZzGxK4WO0Sualb1pMBurIX9/oyDpuiBI4Rdf
H8htGxwzdijpdAw1bBtOKSviiqarrBfk4M3qkcCr2b2uzQNlB847BxhGbcC1YJyq
yLSrP27a8ng+7S6ZjG6NJFvh8qz8BI0GK2Sv5ps/iAPccr4uPJawXe+sebvb9Djl
EeKiMBzCvL44yYVGxCoNGW+nOaYT8j2WwtXVQBRE4jgrloByX0QJ+DOJtIQ+IVnU
yRMpQAP+Eg8Bhq5vKivs7fg/daNPjHtU522dMIIQjELuy9+4tWkEGv30zTMSMr86
R6AA3Pb0rhDLUu5whbwtFw6UtE3/2DG81wPuUOE0OoLgn0RmQpuilo37hvz8Y3wy
mytRf63AozND0IaEGczDukZN9Bua/Dj2/UE58RcLw+b+3iicZDt2P1CbzmmCswxb
BFg8DRN1+F1/yZEPyb/3utlp9bpRBxbBdpOEvqvHk1IMDqEoFUQOBnKcVr17CRJs
CxxQg5J7F/suwEvOaWL/cFEEOMGfsDkIUuWLFFXb+lnWagvIxZD1ZGN+UJvoXsxF
7SyUrqsXmyqsMHPLxWXzdAca0ZQLHfj3DFO2nEJVnGFpH1feUDLO2LFGNtFb6oBY
sVYtkCwH8HW9xbzR84KpjUBT63LTDov8PWLYS2IX6j7vaPbMul/YNfW6I8pupkGJ
xem74CzQXVFRdz7r0GI1qX9HzfrwYWpyDKIovniDg0q7GIRUGFYbSvoK2ZXT1+zr
YuuUQ9hf5Ut1yvnzj6r+6qdG0bRBbj1l4+SmEfzXzPTZjpFQDnKHHQBSBI2q981R
hzGMkXb/JLl7aMLVAFTV23LYCtd9Lze7wsB+kU9IEgc6ixOzCIG3J0KEaF9PQ9Hl
o59L+55Hs4bF4U9fmJ+S5/yE1KZ4Zu0oLeY7b8dXHIFjdmzkGuCXtoaivSKfx7fx
cMnoI/qGSxxUBC0BHKc1ykTxxBpmj4/xptcoesaMl3dkRwGLAw7xCqKX1775qSVx
7TXMQYCs4sJXF0FIpMPJDuV5Uf+IaaBKsKuKNmU6jD2WuTZj8Y0Rcu6zzOwLKjKV
9iTnDhnvwVpdShJ2jMobgW5MUK9JU1QbA1tDP0TkYyNFXHua3O/1NKIWPvUnctGd
VpAHjcODvGnU9tZh+TYh+Q8FH5TzxYbWSxFesUkl9s2v52wvNm2/PHz8GQB7/kKe
eSjsAYrHKgL0Z0y+uuwWIZx44j3r0OlGNyDruJbzhY01//V5XoT3TmmF3ligJu2Q
anVNTkmQUcjxuSszMfH0ZQ2AkcPHZLnMGJC4vJVcPTPJkBGweEt+PDOieQOCuC6O
Bd4vudInePSWjysC7xp/gWq6BUsTW4nIEzbGeKPCCNixGzDgJnLqn2fRec75dCi0
siJ9RPfrxs0Bm6BOUCk+9kPHO97YH6Friuw1BnTiM6kymBuZ3RSl/d3xSRo53ywQ
1RTrs9vot9yli91AtAP680t9jKKNMvf4IJpLkVUxa3MwSVkqFGRvBEp69EBMaWDm
P+1yqYVJF6xUm8TpeBUpuIPq2+fNzk41OSpBUZllhCRjnDSDmk2yhezXqxnzRxxb
WuPFRLhHlAyYkOvnMYqYjxziZlZ5WS6Ffsp8YWEHWSECj0vK57KcOyz3eXOhXYxk
CYlJNN8aqRYUzYp8naXnFKFTrwey8deLG85aERU9kA0PsRFFQreicVHYI+o0BFi4
cL+dpVyEcpsUw8pid2Q0aFAoMfKd+fnaFsOGDPcNTNuB2jAacV73X3d15ZjvlJ10
z/HWRkgmOz/AgQteTdUW9TRq0Q7ix1VdGuEGsuTJn4CaDG4JSOzE+esHSRZIs00n
Ob6Vj+AOX5zA9J/3cD8g6fcQGZZxfRrZ4RN8okacBTgFZM6SD3pp4IYmI4y7wpDW
ak1Nk9g9xmpyJlm8QXdoT8h/rlZUwTGnNSvSGpy/o/OXnEPUVxfZW7K0amSdHDe6
Zbd0uNq2aQjQXt9DLtegXvhKlNlvJ2Fz7Gv5hR/1fFwxmdyskvqkrXcy6jcnOXdr
zgdP43tHWgXqnqPY0cv26gkpoiADkExyH8Q18pv+/m9PCDFRopoNQTfXNeh5VlbG
WHvqeHH3VjFvIzn7bY20pBHaKSe76GUV15twphnZuqA1lzVwsmm09ncjUQVYGyx8
MDvQCapP16SHsMemrNWCiOvCH5BnYGe6mSWmRck4bn6RePLnL4EHFZBb7vxQh8lh
fkoNxQ0vE7eTL7AVGs4l8hI5WSUogomv7JsAsVxI1AVddNi4wc6DvaebquPivsMb
Y8eCX1o3rMytpdF1rO0ns/kZJ3mYahI+ezfapr6gYeKC7U6bsX7wWtOu3PaUrubD
XA0r17pn4ZEeCTekhoJkPKBJStnKIvYVJkkiPBLvLPZmDdbr9BsfzHpxtDi1RAHL
70Aay5G2mOe8vj4iMLSECd/nfsOTL+AU+qYKc6S5nq1MFq2wh/iv7ImyMnJNFDBI
FwjmLYcso7JhZ3J2RCer2qeFib5E+boYFKVAMjA0wQCFyehjHcML0sKCjRQ7qKIj
D0QjzivB+QpFfyE77kBdXpee15dA3gnbcCBSKhUtYzqej4849ywqsOdCtSw3qdWS
gJTIAzGO6NclkAap2Jp4mVk9z14/I4x4ka8s7SVGtNI6ChoxJNE52cyqiCnSQPjs
roGFxT2ull8UvHjA9amlP87VkJ7DVI8MIJDp7KN0vwlZRcr7ltcVC/gh7rwCuwCs
PCFhPHGze4Y177P5vFvSQ/XMU6Hsq4121oOVcq6gMxDN03zFidKF22fTxNKU7x8l
IkKeyX0EXMQWt73nfBXWIMdCL6h43YV3RLnakTgu44Qx8Lhm+clz+Wq/yUAEujul
e3QfgYauyE78PCgzlLtfeWOvFQoGnU208X5KDxJF+bnPaqyRVgRhHSJqUZmVCRa0
mK85TMYSanutWKWXg+9CsvqS/qK7ywlmZnptAlmhsb0viU51MdBow5mHq/KYHpbG
QohvDeYCipmMaLFbB2rMZCjz1zXLNv8N1s729J4QbzJsy+kk/G7aiLUdDWp09NDg
K8lH7X4SbQ4Y8wmGX/VBlNjlQTvuov6y2xHqIT5E68sM+Z+G8kMxN7E+fXbL2vCu
EybEFhmsQR7pRJc/Wx8nqXbGo6nk8XvIwayUw5pQDePgMyFDCcYHaVfpSBWPfiWo
5PFJBDWnBdQ/Jzu01dWDUhD0BwlvONJ3shFGy1MC4PGVE3Uz+kdbidI/R0Ie5YcO
ZTTke5ppYFY4v6PaK6HlK7c3p7AVDwazsz/ESJMAUggg4Mxe8exzgOYAnhkiSM0Q
BPpE9dhK2q9EjDtCRc26XvUOy5AJpccGFK8T+NqNeZ6cQ6kq/pTzJ6FObgdW87EL
tQnr+p1nqW60MK0Tgf/mx/yr2EXSXK+BYk6R8CcL+azQmZiupEeT3hEqGV0eBLIy
dDiwPMbG7WG905yM6VSxyRmUC4oQOGMyWA+O64fJjjcigUG43LgxVm9Fph2EkvKc
1OhrD/OKZ5+UkrTQOpRif6gcIxApBRVFHpPF7yxmWFe0N8E1hQGkqrKOKYq5ZXXu
7EFLGHDUrWXFZUxvaZ6jeIMrcUi+H7FvThuHqxPglTjRgjFW+863gEf3vvBEQSRm
7TFZpu/U0okt12gN+Coy+1OomkXP1eBxenlmDtkpu5Cm9KYzqhAFRbFCxVK8kWYT
WN3MXmJPPsWzsBE9sJh/NcUVUMlZnzRPFGW4zz/fQbYtYPzwfL/bj5QBMuN1Nlec
1XyE1EOhpMALcB55PoC5ysQxkQU9Gq/NgA6ijhrOJiimQ6V46i2PTxYFkiofdyx/
JaJVQmuMo++MHxPQ51ib69u9LboXJR+zXITeFbi8wdT/6H1jmOawbXcvaU/1i8ZB
3qfOlCsKrLhi8z1T28oAIA9SjybZ2KBQh/nHsDHbiEUJ7tRgovVy7jvx9kh6E9Co
LSfZ++bUE/d6pSE3Tsnqi2Tm5NDNdY4u6pinUMRoVSx63XedFwZswz75MTF7BRrE
v40HauL+uFKKBvB3wxaUT2eQxWlAMb/cRe/IVmC+1ZRUgkwyvx7IhrNqr4KHHSCn
SsbxBsbZa1cpj1bc+U6Ngs24XImokH35Hk6PyCCwofGC0lRL95UW3j3ukd3wWgIO
y1SsdjFlhbhjfSyOcpzO4SUBqMp61lZT5KDYFhBWdl2wWGg002ZZf3O7AuSloh0w
leS8WO3VuMBj3xUlRlc+oeyZRS4KZnP2hCY9fQaciUv1HveASWwiRh8T9S44av+S
f086HUtWGONJGhIYElVkAM9JhxX20N/2wLd/dOAgmYStnH0dEDJoF6ROP70HSJg2
57sNGYOzeIdJxX41WveqMoRNNo7iPfM0znFuOqxuK25BOwqzSC9y/MiN3vDxr8Mb
9EDD5vLcJNrWNuMpPQrBtgzaWrsjPxvP0NoYCOeFTPjNC2sDOGT9KQ2BZxLJg5R9
EqUJIfZqIrDptqWpSG7Pq4zIZYqd3tbNkCjBipHqZE4ZWc/PT3BUPj3KA6X9vccG
aw2QieAKjaIV0/HFY9OkkOTZHMN/tsZdPnGJZVRLYWCIoZTOpKt92mnCuf2fv6If
KMr6mBkWTFyCX3CJBSbwt98Gx3MdVQ0RzavYWA4qJrVKiYeM8E3L0wD6bsryzZMd
7n+vyjJ3ckGPSZwFoiYCjahVZc5rxLBUAOrNt74dX+GghQ7Mx/oR8Ng3ihk6lXeH
NAKwHz7ATA6vmRyYQ5yBuSAYwoabDy31E31DEUT5fUoZGXN/frG85+8vAiNuW0Dx
UNddg00pANe0o0lj8dZUqNo0zMSwiyPKLMus1j8cm9vmsv5wBgCAojT2yBY2/uKM
7tmMgizee9xTQMKOHZOy/1v/v8zBK787GJc5nHBIYK8McHN2OwTlgmzvbiUaROBa
IIIOCxN+JXm1TMd3oG4VJp/EofXqvb3Ymb38aP4QRPVT3W+seTRSHRUHCapqGsnQ
qPbHEZT3Mfn+JhbkIvn3B+ftUS5ziYquigUrzV3YysK2gcfyhAALQsRXVAB1RRAc
3lMeH6nz456w8qFhP9xIRSF5JFS+wLtiTj3yzZ3pnXp1HRQp0PDyBpaS2P4u7W4A
9kmDfHZ4dTV293/MeT1znPu3o1toJ1swH5pKHp8L1lVHl3DEo7LXLmZwUbcyCdG6
cX5bAdUdR4vcnTO2oWwccTF/dLSouD3Kd/J0THUi4mDPpwxVVEs4tu6x9J0SDHT7
O31L2m/2xwq88SglHpq61Gm4VxMxg97z4PFTdp57knde2M46+MpzndOpHsSoPbvw
g0IqiyPtX346SpWrFWATH0VfMGV95694wlG9Dl43EYIABF/k59nfLJjkQRBFEMgf
X9FzHuLvqmRnKVeoPggH27dBBFOK1YSwyt7x+N084juO/K4OAETTEOLwmFVAzJr/
ynYSZC4MfKqXB9TCflsIe5kggunkCM75iNzzYCqQ+aFYZA6lsgolOe3pt84fOeKT
rbDVk8y/V++k9+PJmc3P2xKi8cvfCBiu12DYnisc7XTWdxWQhRkSIQ6jSN4ToDdU
WA1wCR7nUQBpc0ws59ym+hxZaeLNB5WqekWZdBdB9fMmyvpRYP7iUh64FL+HxnnQ
iohhML4vEM6lLpxiF3DTN8PJkYRQ2j8uNiAgV79rtsGPgS7tyO6bDOegIicXip+X
RykyjrH7jQU/KvwAXIq0XlyDtHchFgefNr7xl2peleopNMG63odNibcVF9QAjk6x
5TvhPrzR4FCPqKifFjEEqA27ecskzPrFhhDO3hem0DzaCa3dB4cDrLVi4+jyUZbr
rEe7zRHI62+tM3LDbg3BtGUb5HKfw/G+BXQ3GHsdK1wKE869KXJ2OUcOsSCTKzEX
6DLgpO6J1nPuiDHELotAQsiMvCXzxqza1owyC+NtjhFQLc9X6Fv9g5CF1plPNCzp
TwSh2xcNMlO1HyiacXelS7dKdbW9ccFXYWp/Zas9nMIP0r1hQkC9rrbU/vZuS2U2
AajLmfTMYSeRpTeYSXOzn3OJ9b563w00sk2zq/5DdO0GUuJ0pkLfopZIKtEa1N9y
TOenaDClKiGKd5dFruwK/zym2rxsfSZRnBjCY8Zry7BTT0UtPRGl9KuKBEGsuyaF
mlihx1w7wtAiYMJqc2VkPfNFNsai/1E2Iv1Libf/mRZboYbVyLSrYb0W7XGOYKsk
BiMb+8yLgv/ATYpUAEnAQQ9Gxsdr67DK6QqSzBb5w/l34qp9AdW3QQVl760h2YdL
Tvlqle/1KXVybeteblslefFZfO3o4WPjSQe7kf5P1BeIqaSTFKZ6fUiO5MeUn0EM
8ilqnYC0OWwOCoGkuYFZlWgDYonYEZ7y032ZZu0NpnG8Qe6M8TLhRZRyvQoEcRyk
tC1E3OgoXOBv/nq0FktN67ZQNDR8tnq94AdeTa7vIrKQq1uoOp6S8x0w+zRBa7zh
1ZZ4OpMpE0qAkc0c5PnA6uKxqgKEY/tIoYyAPDGYe+/bAWhp1mR9Zr4ndc5Os/TO
KK4sQXPW9rkU6RxdvBHl8n2XevL7r4kTiVIyy3vXHfkYzlw0oLZ1gp3De9gtC/dp
gdmoNHTt7sXEL/n0Q78+EO94oly2ljfvFxJAjeLpoudyFfss6vVqju9cGiwiblFJ
iDspESSvgtwdsKtHoqGVi2oxbuunmXqeZJ0yX9EgikwsBH5UgCLJtEpACUXg+0kc
ofqPkUBee9bZsrTCP9/VMOZY6lTJ84HdZ/aPxtBITMgKgiYEhqAJPAMlCUVv8lOU
AYEpAgqkHiKh/TJFKAQEjFk1rNfxMU1XnfSpaI9TvD2h0PNLH1RGE4HYKKcVWNxr
BOMClqxU775tUT81801PX2dEJEGPKoFC7YPG4qH90uRQURs6cJ/b7LbEmOfHRpL1
ogH747RvD9qzePKGtGBgflkkyJGKcPZ9Ry2MmpelEf1YYRACYIimacg6oRORXBCK
4uvuvj+8tZra+0T8X+yVfpYXeqn5EFBGGodeARHccYY9NcLv37k40hugjIiRoEB/
jShj3ChFAGYJWazxFCnFHyE71sUNm+gMq2CSCikkrWp9vlKyHoDBECymj3tOcd35
JdF4c815vHJj7+dPrYnC1UnuGMAvPFn/T0LPbW1GfDxrvk1T6qQItv58D91cy3C+
LQHZO+vdq7riH20nqh/saQ+rwebjIW1FjyD9V0+YFvFXGdM7rCS9nZoFOsA9Icug
VP0AARCWqZkIGxhCjjO8/bZbu1pHvZW+aZ1gpJfUp9HqgF1pFPo8bHCA+ueSltI9
FdOfkpkHqucn8RKTqYWOLmZEutxrviZhv261yQhWJZ2mhqCipTSrW2ZWpmiuMN7K
YbDMk6EDyPWF7E2bPeNNh/75/pOblj+GTScuEJ/hK4ys8y5qVi6g+XJPAY6XLw9Q
86DFOBcurntV5CYJrdr0A9cVLRApl+v59Zzo3wG0B2gV0WiYL5lrNK03yp+meWej
h/NNatbrtW0VCO1mZ3pzDwzlYg1TA+/UduhFLCLhTcNHMG44KH6NHyXBPMf+6raL
6YOL2AZG/fmUvqVYy8B07yHFBic/lhpV4dQt6CHaxmDWB14tliB00lx/e1CBCqzh
1sYiP3DiY6I56wPkTx2O26++p1yP+vHvJ/xb2yLh4DRfbxHZqyeW8wpiRkemtUpv
O8sX+8Z8V51hkKDrHU+vYLqSZQ2XZiI2OQzGwaV0THfvzhkDF4wFNhtCvRPJbhBY
UxQTpUaDlwd4NE0M6RaDiqY/C39/AKsqWLjWrmo7omp0pr+zlxzSrhDIFIe9XNAQ
0Z8ihdcnUlE6YRNEwUCtsBNDCqaogoCx+avL+NjyAGcOENYvViHA9byd8WFycE7c
izpz8G/sYSg40n19y1IO15YMTmcz7zAvSuC+Kn/Is78wovSjaw8+Y8EGiF59VB8a
LodcxNtGOBXl7uQhJOnQzLet9NpvQGkn9bStQ8lIFTfevfJbwTkOkGbuwcsOSaK6
w46PL5MHOthgOhWOiG9ywInNv5SFrqICChtaKLoQyD3S5+p3lyzDbPpF9cHTqtCQ
9ZNmAA0QLqejeNdGMPCyD3qxUn8F7cUB0ZB15RotIL7auFomaFXM5J5ZDmY5PiNb
qRzEom1cHU0vnT4vn6Pv83VThA/GRW8EQ6OG1TqqnBrq6ui6hvMjG+qFwISDGfiO
Ef5Btbtv/ZSv2lyucidytRutwZDdikgXUumzfuwtuucwteW5hcrmpCfImExHcAdJ
KM00ODXEZdytOt9AzU3WRzwN0ltwkhoB6+BlSWIaSea9WGWLZqQJBAPbaD6dBnl9
K3dlF7FYatBugyD0KIrNpElZ5Z6MguFX29J+xjZLzy0fXUXKYOoOUwn+lkdQQgQq
rNvYsf2fW8vyTehbAMKjBI5nBhQ0zN2LfEdtl2qBp5VwmzMHRWUgl5DyGCzEcq/T
KLRhNGUkMPf368W87xOKpfHdzhUX+wKFeSd77rCDHLBgPj/ge9g/hi1a153xWvF1
VV155Kf4tuLKF8wa65JSxrGjYwOaWwOrh3vwVZ3lkNFZ1BhDq0XvCy02tNTW+Xp1
5Myx1SduadW/0JGl2iJaAWB1ekVC5FKdKfmGbn5SmzEb0tULF/D7XOm31MiRIm39
65POJGB7Klpqg18/76ZBlEUgwPmT+zdrXhvj5tnrXnGZnhGELHawzi34EBlZ87KC
zodh2AUgzMbN83Ox1+UgMzpMpqdn/fRwGZYNyOp5pmoBYInGKCjo8HOskRcGQM2s
4PDjjl2EBJpIXjJXLrWCWDASDr5oIpyUF39h4zYixwXWrMH7y21lFRvscdPXFGS2
qfULXHqtGrl9L9AC2g02K7C+4zkP4GQ7uo5tBHni2RXburij30RO/cNu9cWTVBOd
d60QHaHbRMUiagLdg8MXzfOp6sO1jr3lBctbPxekAyCOkSaBoXdBCzGpfOkNGgI8
Ah7Ts22bcuP88xlV0pWpg9jOb1MyQAiDMLMPJ52TRzpsGCrwWtarEWDWK0Rhd7mv
BxvpyrFVL8ttp6CFOGse9xADzxG3ADiOoGK6jbbLhnEApcvLxWYjHa6Zx/5m5J+A
lfd+h223tVyDXcyH+ouC6ifv+6Mj7TRbtTAX9Wg8wo/vreI65EVsrETfrNsH35Co
vzDtgwsmsA5CQeG0OA9cDhfNwmCdpgmZZt5lD6172sI/rb/Oot7PY20/hQX4gCef
7tk4TBVOzXFO/34m1rpKzYeMhG+O53yLdd2mnp8dxnze4TIA9QlAfDEaJVeHgEOe
UH0jnb+L1P4WDRZ5Jk3z6UNsJ1ghJZn9KOYTBzf+w7yO0Vg6QKnZrqbvqk9X/Wj5
oEY3lkxdubteBIxhHq7c+p30HBiX735eyohDS8+KGt9EwcjE4FJ8WqzNY9wNxgNc
B955ItsZjnGOG6IcABnF27wGGX0Jb9M2RFBpJti1KF5KqwnLZTrXbsy2NSHeMgaG
LngXuAgInBaqF9VPtPcTcCN/UEmX2ouGXDzvs63+ZtlGNm4khPc5BKGVnopnJH4G
oBG8GeVDER9Yt4a2AVg/QYCKaS2QcmvN0sItPCo+FjHf6cfSULj8kVD3Pa5zqcsq
xBiWxD6Xk9K9QR9Sz4QzJBWP+7U13QCRSsV5JtDDX1js1zA/0EW9ytJjV3/oFnOP
qPXA0OPEkgC7NZQf2MHVqphUhC/+O00pUc9469f8Qm4z6Idbjv8DL7eaWsFBEXk9
pDCl74PMCVw/kzhywYB+oSdVr3Vvxik7+6NtWmMC/yeFieEVPeXUuwzFHkjPc6zb
qPBkCX9h6A3abb+ee6nj0OwtwIOyW/YRpxdvVrtV5I/Wz/qj0bkX1LABM7VLRO+J
dSG0wGYSXdKNlqg0ug/0d2gfuQuKSTbJv2nre84nI5Ar6K55DAoMxM+sZFlCq4q3
4HTTV9EhpBpslW4BSOIE7khdslIq3ruOc5Xx88H+RY938+Ev9culDv0Tl2oyBw+V
9M9GQgSypituln+UhrKRElWrDHRNvbf51rDA8WTtoXNnwRN+2F+j05UxQ/q4TFef
8fagravSmmUqItT/pA2Ok7npIrHyecIPC5vehXxcHP11WqXHbwuHvqml5A4vpspW
7EZ9Z7sbCzMd9tXO38StDG4XSetzPs8AztsPZOLLp4ouC1+TWGUMJ6KYFSLyckA2
oyXGEg5GrAnObYsOAJA1wb1Q/ieZCudQdREt0Gj8fnrzjbFrzyZtWS1U8wOcUNCN
FCqtZBmzu3P1bXen8xouu8cXndPgoTbk84zO1Hnv7V1YBq2yrHnFSQEyJ8sUuHTV
QWS0R2G0OmuCYT+lVW766C+ejvkqvIahwfKq8Gwe8LggBcHwF2WfGYRVc3K+KeG7
jWagGtLGNlNxPSMLFeaa66OnsycEKJTBFpJBhe67huV+DxKi7O4OlSS7FxNhPyaT
RT5Luor4rJkJ7xR6eaUfKPqvMixZed6Dcz7QWruk1FaaE403Ee2X38UJwkg0goYn
CFC7Mxef0AFBlypaFPNuV2Ddhv1D/FJy7rGF6fp1SUtAUf55RBLtSQJ6tNXCUdBM
jJFLqVBN2H4wWnGmwC9J4fe9twHS2T6Bw7KSxwrHEaPVjVfL4Sc7f7A65Abf8MvO
cguqO7gzvfRgcec09YozXxgBg4qS3OJGG5igAEpMr4/HvsF0M56jEfIzg2tbtbzC
IrhaqhJpFZbCm7/6t6fKLdxUZoMPvckTRzr4m4RozUSwh+PoWr052TewA0GYTIDL
XeMFDmsWtqlueQDJ7S5yy0FTk+N0McfgySZjdUykJ4JahE++/pOJg0WIXtDIxPB6
Kd02wZ9Nkf2xUekT8gpnNoJGPG3pHa+FQBTrK9o2B736li0NijVOL1F7nfYd8uTZ
RVMznQEeqsT86WffdKjhKXxtIF4M/bT97UV1wBXigZKYLkm2F0v5qQKKW71yoWaq
SnK2SEpyJ16vhp1cTgwSnD2Rwv5yfPeLffQppXyCAk5dd28EwnqfntBW6DoGzBSa
c8U6PyPGiIBsOspQRRKpIbRdPun3dtqbBxuAUyQ45hA3f+ZdcYzSQtG2CdwH46YV
JUBDbK5ymtZpae8U9HWYH45D0qg226vtQ6hE6s6d5wpCH6qUPhWL8P+/Fft4tRNY
PF8grgT1AWk3eUlUBdzkr76/S0qPuPzUwn5xNxodd/Az/kUTVjuiOMuDQ8CS7YE1
Q0rOxn2ESngujjFQnb96IZ+KNrrM7ZSWU40YP4Lfx+55W7rH7Lo7MFwFNOgudu/4
Ir7zeNM+bNjS8TPXPRaO5GDXV7SJPRpb0b1jQ+0wO+6wXHVeFNakhS8T7UxwcwJS
XlXxVusqchUZqLtYRnX5468GesxJZ7foQ/W0Zpl8X4FSAJumNQCxUmIUI6vt9ttb
riWi0ieUsTpD1G8A7kduIFSXC5Opm1lZV7YGQjeUX7cejehFkZWO7NpvbztRN/KQ
kl9hIOXT0zKNni+TS+DP+hPynHBir39tfUDI0gyoG8M+vP4RbwXsDnCuXN0MykZ9
t990kUqUq5ezOO+SkD6xZ2tzuq+HZwtQ20lksofmHJ601pabyJJLMtv488yXXMDc
Zgp5KlCrMBlMO62lSY7XotrNVNcfbsrUXGlTcG731STiq5kr8v25ZrUIqysA8ke7
BhGGaNhGl74WNW0YO5Zrf0cUaT4YbYCS33McYJOjhvrDPVsyGV7cdtx3cHM2B6x4
eYd8eBl4foL/Md7BAldSeQpQBvluse2BaTAc1oH+MeBP4MO5nH+VKXG0GgpvtlL0
/bmwgLmUsvA4SvZmHYEVM2JNV6Tc1OqdwO5mMKA1rF9YmZowfiPFX7IU+/p+5Q6z
DzwdstXVdmW/li5U2HHhrrljpzsKbrldVClJRMuf+xT9d4Ezt0PcGQjW/FmKIIRJ
9mPnfY8Zv6zdJBPTnehLWwPzZblC78qKMw7tMN8egxwjrTNsHdI6ct4PftLXOV/k
fS17iMRoaKiyx3BLfkB3036nllM9cpg/HQMYC85qf2/QXgtqVHNK5x3QCIpRhQFD
IA8AmRs9Kt87iESoUorjFM6bn3U7L8mHU3I2RMh/q5vk83sJ36omfHIzu6go3ztA
rMFirNmrujK7b9JSf64iuFUPzTsvJyDUdkUfB3j6VI+oRo/XTV+fMorOm8a4540a
Jew/bYBEasRNqUdPdyxh+s069SjEF+GV3aDdQSxMaGPhjQ/Z+zcdVC3TWF5pyy35
cmGBklCRhZxMFS4/FZuL+grv1HnT2EnCwO4CGhUuzHkJ4DAXEMMFFur1E1mZXChE
jFqVOxElOOsGXAGhlB1G9Kf3YAQ8BN1j5U/er1SSsxEEh10l5S2Timossr5PJRlX
zPuv40OohVtsiSZIjHZ97Fdub7PhiOMlLClw78DZNG6xROty4hZa+vrbT3XW1JnB
LnsFZ5DQnqkGLIo9jSBA/Uwc5MnMYifPgzFgrtm9qYxidxT7tojVCKe0SE7L2b+6
0N6bpOZyEnysA0j2KQ0iwgXtoIXncVLjLDGPjSwtEGzZdxr9M78n0jFhgkT6sYkv
rAn511daNVSOrcsvvHZq/F+mcFuV1G3YU21WAjdzi5QMDB6xhL1z7xZmEggFvkpq
nVyXN5irXgTNfyoReha8gn+JG6O3d13RST4B4wPAf00pjOXkjrkY1W3ghVnGhPiB
IE+IR2QomzgI9YDDKLZen2Nd/ZPPf6X4PGY4M/JHzwmCj13u49fcuZWy2OvIWlCI
c4Ni+7s9aWkB/zQGAWad2CdVbGuFMiwnlzGKYI8GqV2T3HJKvzQAb7f2EUg/Wcgu
QMBZAG61xWXrEGTbiR/DO/ykhc5F98gRhJvGHIeNU4t3UPH9EX7lSY9BOZEubSdz
c6hVbRfxbUKM5KnzKX2vBxFUIwHn0sviG7xJjR3vSYgiA63OOco38T2b3zghYotF
I3xcF6u/H0EbKNGu0EikhJDQctGIxQNE83K1oUSoss75OFnL85scOWE3/TnYvsqQ
ysii6aNr+0kXX+RH9pbWihDxH8tUtIR76j8Jzrh7jNEAdrbJPp+cwRWxKjr61QGy
CVzY7NyYH/9Bv4vN4rVfgUO14SMyDUXR3gPQGTNk7cdYJdTa/T4k1Efk3W1a/Omy
BiY1VCbiRQqba7qwBZRaMSXjk4fZLsrn5HKcx2kFoiZ1kAq75fAV5y/OjA1orSJ/
23YSa8D9sbsvZkyyQg8714EQ30CEEECUi014tqxrog3DjXYENyPX45IPP/0BAL1z
RO889oh+ZNFYEeWxNhJ/jFAsSZ8tLbgAupP/p1bhwGEUgD1Q1ksESZ+3gXMqjb50
eTMlOLcqLDwATFvqxqRbQPLQc2vsS/lFOkZNNy9DoIPiE/jLDuihE858n86iLIG6
PZlDnXYLKq8I4yS4l54m+bEdNdKlgYInyRRUgWS6bzMHPw2Vz0wFHGA1tSP2Rw0u
lvyf6j2ehqAcdbVeJ9I1S+Gnrg1SIw7hA+4RA7xyiFEKikTGoTqbTtHR3u4Ms7C4
GQW9KMI78zKQJplRACRI7zx4Wm7y477/3deUyfFbynNxbEfho/AiBpOfpd6Fq8D6
3l86fH013SDEn/n2lsCw67CIAN+wasSjb+sV7fs1uZKB+/+57+ARDPvS/ZL0kL/W
nuKNAN4H+2sqTeqv1Qalw1y7nfU0is2gmY2PvpjxGBbzFqk5d1J2JGuCCz4WmKaz
wyeMR6NW37zV6JZ01bb2xxFHcfUGfT1FVuPC/mXbSA3rkdvavMlDFqX/Xpmu3gIX
+pNqXlHNPkNfif1bpY+AtBIlpX3CXqBoWKpvrD0CjoDLBPGDYMTIYmNr6euPtEwf
gUqRcHe96H0XaJMOM4AKGjpKyUIaFQ+Lb82Zo6JduZx2G8oUfa5MdvRm2dNEDyOO
Q44wI66jY94PuMK2T9hBwBDMactSvFFLthQF1XIC2SWe9V0vX5Ktc5aE8hOO9IHw
6IPzH5huaAkMe33o/us9LDmdLLL2NrS0fn7DPeSC6Ael/wzeLmHysVUW07M3Xcao
/xtQRq61/ZGcFazcArn5QZv2IN+VTq/VLnYdG+iVhXBBN9NfxAKuKcaJIwEADmdq
ZP9Ls8V7hqekEJ51exwIzDthdKypYb8odYALf9cYy3w0n7NIxhSuhXCwsowt2hSk
/mDtI7Pl0BcmKQSWng4TeYkYBuiQYOI07yKLJTeoY3/g05ija0NpTsyz/zpjdgpW
T15xYZCaUg7qi2TAGv/qr2SXUggDmIFalw1Y40OyoY0ZgBVJfTldUscO9muR/V15
kz8dpJGPu2/knv9FclhWpwjAtl8SZYyW3YogBr38E/0cVOD8+S1m3fuFjrbd0wuG
lzzxlRQWOUeLGWAUZ0I60cadEsspfwSwfakGa7MCSIAwk7QGgrbqpEXyNTxK0gN8
y9Fj6kApXwKkG2W/jfj8bpyibR6EkrAJJ8VmaAaC/+kmlyGjq+9p00fobXqcF26A
HXIiqomQ4S6iB4kZCKpW1zGiIyDcpcqT0tvMRAMN2jwsGWz+hRtGejZ5iqIEamTU
2S92AeTxMOV426B824ecejGKrLIVeMJeqBOAWJInKkO9AgpkVoy0+lpuQFOyX/ci
KEcQ/CsOZsa0yvSZFaVg2kv4XrZZiyVMBp8c5pod6uaZAaVOXDo2IrA7JUR9nv1D
TleQdNkMvVhdsfGUXJ0v0M3wilUVtIQOOW+gHWfwNQoRvEN1YjGoozF8yKVX1j0a
Hnq+nTymijXDyHPb9doSqe7L2uxRQP6aKWCYzjvaNGcSu+r+L71SBKa+2AV8GpsJ
GsmzuFnZNTns4nC91vRytKiFLOOQEQY0d2aRhTKkBYBLkOYZQJ4Yc+9g7uvnUOai
csmci+iObkRHB7OS5i3h3GeQ/phVAW4P2rZfguoBk/H45eUqGc0A8yIk2wX7fFHb
7SIZ819fQLtXSaf7LxTtyresseASfEQGsty0jnHRC0Gm6o8cazRlt4GJcdWRlGA7
NixV5bASML99kcgyoOeao9utJembQxFuAXW+E9KOVYYFyoohI5ERA5lgdZlhRR9H
PQfsdQtR3NSjEMnuy7foMjgQm7r1tg/kUyssEiloItBDjhPWGWUoHedtqBPL/Dz1
W6L/SCQi24gh5iOo2oCyAF0hSsoRRITjKXiqFlgVxEZFjRO4QlbR9Uyva+SUa2Ui
p+evtN6G8CCPfyTip0nDpTEnms2ilnpVEDtUPnj2AtWJDwWey0I1v8fNjFK3FVg1
Fvfe5ofdW73Z24MpgMVIhMLK4w4AAz313nD6Y69MezgNDMcF+wiA46f5qLBmTsHT
5pWEe5jnhSWaMrr3PmpZbc60765x+iXNzlHwU5GBhN1aJIjJ/XBohRXt7H1GuYih
4UmJroGwVMEP4mu9e9nrdXq+N+XsDtg/laFWwiFca5iabRC4rc3NwFDXYAdk2fIz
lnvvPlSOlB47A0GM9M3hbd6XgpFxyh2HdioenBMObU+vgtR/AMsKhnwmf9Nlwwo7
d1dTVOcskodfHRQuTCk9Uu1vfe6mi0/JEc/3txZecH+YPUwLR3+oq2CNqeTx6MyO
FxqKw/Kgy+p7nfNGI2R/cOXGiqPufdr7fdsDNGX3HtS33lHBS9ieSmMFSutI/Zeh
g6S1EXF1lzhWiwjzbvhClICau2e4mkcTOi8LNzz1PHgr9bbOxXKYnPc4egyzb9FQ
frHWsLKofl5Guep0relnpZexkX6qf22pw7Cg+pDO508L+jl1VJ/01TFzJwB0VbTO
WmKfV78kvBfKIS7QwBHtGgd2CO6FA4xV4R2Ggk50T6YuWJE6gzYwRCTtvznVb9EG
7l19UzKwHJMnXmyXLUOTg2NhmHblH8uyVNx2YmTCQDP1zSeIPzoZZBLqSpBELb4v
zgxcuOvy8QALf9JfA/88nDf1bGLgN56CPQzStjvx+v0S2WGcluT+1D1arx35oQ1B
qXoNOpuzSvrRp6apUEnWYUXxfP8UT5G3qaQ+qxfwRGd4r1z0RwIxMzGzURYuXUSa
ifxVrq+eVopmiMtHYjqltQa9RYhlKqTIPJHxNo2QBqhPvWXORspzvVRRslSTLGVn
GN/FQaREmxF9A6am4ODVM8+PNVRGwRE6XPIuzYYRNXQFOUUbm1nddgMhSunvEqPA
T2BmzWrU/NF2JtAKNuaLie+DOLzEHh+NSBUQw+AFB2SFab2ukfwx3mhA5SPhM7cR
UVmWobAJiYg70U90zhcFZBGeDZsO3ywTwCfLQSnPoMUb8t9iW82C1NYQqwM5wLmD
Lrkj+h6BoP/tLhYItGlOMx6Bdas99MUizIZ9ZyL3aNLdF1DbtjKMXf9aWM18T/cb
tMyQOprxmVKs65Ivmfmvnms8S4+J5QpZdDSpnbJYh3sbzZRXzy1v/1UTE3oVjCTX
wCKHBC0n/bHjpOZ5AH54l1fbLfwIFIwffHeHVhXx/b38IZSlnOTTVs7gC7aHQnKT
3quZfEJV/dClcGk24INXF8zCJch5nMhqsSYBqb3B/FuS/JTls3rg32g0Y2aKLa+4
6+FCK1V9vkB6VLq7BEVKDCX7BAvS73PpaS60e7ra/s0e18kP2FRcQatgOx84mfhe
tw39NE2OzDrVkZJ0UVnqav0RegSuXRF7fM5KQToGXL8PQ/ssJx6KHRtk9NZiVmn0
HXcHWUWLfnGzG9uKspK3/dvDu0rphdJxmI1n8EWnLu2jlYy9+0HisMLmUYVvuxuE
hT+Fgv5jDf46da4pZpviv5y3xoftm0iRL8f+8oI8CsYu9/qVeWZMq80gr/Nus4X3
zOLNLxx1LnR0SqhvmfWXK5BN8yrSt0F4uBvui0b11tgr0UHWQeafztpKzyA6/lxw
OxjZNLudZ0jDeaMpplrdoIuvR6fk0oP+W7G3LZI2gt3aDcSUoy5wPXcg9qMGq0UU
YorTtuDs2/K5ORu4uBj8X+jLhODS6Q8eZY2LVykLh4ALnA6ea8R4WDM2fCLKhbH1
dKS6QSZkpoCmdSwTuoyaFvqUTRyp0nSwFEEWvaS/xNcR1ghXUrQYHU8/YEQFnF/w
CecQunIbnh1uuCrSdh7T4qVlUDKgGMz4fUNlVKcGi4slZkrrRAdX4RE8+mcuPFF+
KQh0nNgCwLiKEzKrMQ+fccawcshZn/V0a8Z+YCfKqKQUjsfmiwwcy6qLW4Aioxe+
qyVSQeppusbK2VG7wtTHF4eD+DJt+DJAkb+O0sE2uUOtOJ6juxKB4VRS5T9BPFfO
VPbIYfTnwpRzswZCCUZi0flJ/b0USGnNs5O9xvzEWGLmVFriVgvXrIiy9L+hy5wP
jSrGxE2wcMfongaLLFiGC+cFcVAjD51yLeZWQkpxuDwoECn2ZR48aZFT+UrAkUSh
ow8m5EM1934I69GYwdCj37S5xh3WmfXbc3b7WllCsUhgqa8k6HrzXfpsU8mrnHUN
Kp37+WBxi86NYeOsxgNwwYSj8WyzctUhlQgSVfsgKf4bx4V26rGENYYTK/Ui+ZS9
RbmACb8n9k0Ab9/nWybpw8DCVbwL+8a7NXO09Y7f8avXJjdK6l4mchurtvMuMy4Y
NsXbmwWnc0pb1b8yWjRCzt7G5zB2zazQ/uKeIUgS7Cb1hVLzSV0+tVA7zOkQXOfA
skiBDiM+UV58rGCeSJRnZsSNKXQ+NKVgeb9GVPik/QpbRXqdQ8sMZS3iKoVXJWuA
AkWlSqSYdicUzcUT/6FLiiHBfyJVVLMejFbVwApPyWT2V9lml1TgGEX6qmP1yAwm
q4w1bIbgbAO/nTj+GeYmS6I7OrhhLH/JIaCcZqLrrqJvOfHBBheN4FpbI1eY9W6D
SSyvRzVzEqx1NAjiyMtc1ZZmJ19NNV8RKL3WLAYe2ju+ZdonYsO4Gh3cNtzKuZbv
8Vl+vQ2vcIW97t6wsrkChjdrXfOvNWvX691c8sCbNFdE9ZNu6CaQV0s5ApCE3e8R
FnUcgvAtM0z6WBDDvM6mM/ZJlyvHTMCKRds8cJ4UCHvlfv4hVgGNvZM+KAlJOIaK
A5weAkKaswewTgodw5nLZTaiLaEyRpcbQq+1N/bTvMPjsRxAQ95x6GvziTAg77L1
bwpeLoZ3nHTvDAz4RWrcO+BkDov2tS+uC9DAYUjwzWxECUx8sGQ35gItSPfBB3f2
qqsP6935Y1Y8Fa4rnJljC6w3V3BXLaSVemkU6wCjKwrPC5311S1rLdapWpg6hNdm
BOJulenZ3ZK998xasTM4TLjt2LaXBFrL//fTvxHWAiVr7+CIyHvXvbOiIuxC1beN
SiF/LtsZq56mmNhA/Ph4pi/H4bT1/lBSN6geK1xlQgBXc482Pwc59tNoRdz1wevX
E+W6SaevYxkwLpcLclFP1ilmRl+11GbdjsNJHOc0zwitL+w4HE7y+kbzyAc3VRqB
xYGfkRG3h3ie4JOsSCMQ7458Pe522XjQcUCijifedb3VhOZZlzFMMKqkfTgCSZC3
w4iUTCk02j9w32TZlZdbj2qG/UQ5j66j1XrXbVwhy0UY931s10CGkRcMPreCYHaM
UcJd0GcEVVxSczzQgbrYC1pQFpr0o+eSs9v1HDmDLqXVgeYYZnRf5NsJxNLQI83D
Ti6jNxT6lgXXrYY7UGZ9pCfvDMba+8RxFsj6nzl7M70bSDwvVHULxT4ORjT4uMpW
iLyVxMsObN1WvRJ68jv8dtvYL0dSMI5opDRNSsV8hMswhUre+iCJbkapkeKUTzff
4oSd00sDzHC0241he7Bh40tpHyOeXKkbTGC95PXfF+XQvKO9M1AlszHMvK2QtfoI
jmivHHAiOd+B6gl4OriT1xm/WJvMB5rYts/UCjRR4wWPUxUIdBAzZ6GuqVD18Ogl
VAfskRUiulSzIJRGPmXRYz0fKVsKX5qtvxqNkiAVLDm50aaQ3jEhjm+1w4Rv8eY0
YoQfG5xgXkzp0YDDSKCe+yyqBNmuj3M0OiVKvricFz+Brb84iB70SCx+4/BN3AZd
DA2hoFmKXBMRzzyW1RI9fdFV3NstlR0Y5r+M1bRbMc5tLX7lMrcazahpRR/YoPRh
Nhfzm7/PX48qT+NwqukH/oguRCHy8wA16j+eKk6OhFCxLjBgDVV+jxJxQcRAM13j
86pJrO8E93Asn5deRfRidb8V43WKrM7a0FqCM7cv8A3mphljIK//CW8nIs3jlrj7
Uszd4oUeLWYxSGFB8CWofZBTT2WtypUszt6uxrEqtiPER/AqUOAwrOq0IctagIKV
a4bpSHIyg/FjzwJ659rWc+UkQWYkFcSAyXUvaCeeXUYRyfpVSq9YEom05Pj+hmiY
d/zYzg+rYut52GAAOUiDIfiwq8qH3Wb43xEihDhpUTx106urUw1VOntFs9CUeGHi
+m3ijMLI2McCV0kRtfsItyl8JMt65rUySTD+dQpjNExHPwDx7agqmbcuK9hfuDVe
9TURsTVvyhrKf6AZAW5Py0uGAMOVX5EdVGWwvdx4HVY62hfJdifYHvINTHXmqCaS
cN/OcKBJMq0KDxJd6NVgYoLfpDfqOTYybBKjIu2+k/0f8UCBt9oKAVc33fL0CsIq
OD/OG/dRkzuxi3LNLIuHI9oD9J3Fb3R2ogzPaiHldnAeqkr04a1Bzqj68P/nZTEE
3+oITWG+U1xutW4k7ZiESk2uDFvIlkWuFyBcCjTGUd8tKEJKklVut+ZGinI4lQYO
ZivD+GdHapSkzbzrSr5mvnLTIJmkGdjQ518f804MVBy0/UsUpwd6thswhZYhlZyE
Pt309ZCG4YE1+6OBfRRmWIZ60yjC++3xL4KE+ziDJQDK0xFdiYoZtz3cCAHzDdX6
TUJ4nElr23yi2KpgT4LRGlaBd4JPJf7c8n6x4LW5cWOKkrfyt9H5NAdCDO3uFKJq
TCOMdCTx4S1/e1SDyNVcgAhGnkOpmWIJwDUY6mISsc3Uhe+XSfHQP/IqGWulDzLE
IYvLTa/CxsWHnfOL7kfD+dmrQu9Pgb2YL4aGLt3wUC+TN7SCIiSvHBodX9guJhsC
iS2mAlbwFFZnVCq44qBJ8NNgPc1MsZ5v8TcJplnB81yjukGbx7EeYlvBGuwWBiyS
uMm6/KtxWqy2qxJzCdQvGkC2jXsr58bNt2Fv/p5fvz/C1+6rfHVjfPHt63b+pUJ+
HfgrudDN0RqVBdFGb1TAluhq2XounPIkzFFKlll3wEdgkIwzlLeYqO59FA0TjPm1
U/zBCcM7cuzkDRgmuGnCMSDLItqmXIfLKb3RNdxyW5CxAlnXW93KgOa0MhMHUwDA
aMgagUxfQF7Xg+sxl//OtpsNqyPhEhEQw+1BwmqxUfsibdJRVulY+yFgKMq7DjKG
71z94w3qgV6cVco2P0YJsdVnT+zEzdIjQpyoKXMn5qTvzy9R+zbV2kLilz5xq09I
jdzrzwjFkG/3X6UlCixaS1t/pWv8M5MjNNNEpYU/DjCfOmLMdrkWHL6sKdnu/OHA
tXnhurJmyz8maHP4GBWTEg3M1rtOmwKnK9IslPtoMUHtgTS0usDb43lckVIgxJ5s
NVO2Rh3TnHidtQEMwnMVAHv1pYWyIdYe2KqT2YEDUCchIR6y+1NkfiRDhYQNO3/o
cqialClsDFJ7OR5vHnXtpXH+yLfreo+LbUOS/1glnL/lkFGKbmOjJU/4ascZmu3A
XrvLtYPPPae+GKxrrBWNg9x+iI9thBlDTeLGUA9kSXhpS9FBMKDzAC1b+Mm6HIMX
ufeORt0eS/01zsQ2tp1kRuVvVoLy+Gtq3n2ffZKQ7aeWdK0VnRmE5DyAgtnrq6WC
1Hdi1fIbCTQNpVCMv0wvF2mWR3HPe/1JQoYOEjRVzvWd1EUWIq9a7EcXHxEduaul
dG1/endwm9ELghw3YWGMhacaTdAyj/FhnAuBrT9f2Y+1RIvHXPAnDQYLel0bgDNr
lWrtYFwgpa0k5Fw2/ErH/ShFMbPC0Nc/KE0b4ylYl/UeRYvJyrjvDQ0v9QpOYApF
UPLUuo+bqLNtGefrXPw8Y9i61ZjguzoKhktCn0AEwx136kiVkE2QfRsFcjSqlLzM
TtMlxB86ewi7QsxMT9I500iRAvbYvIsjZ2iJDUWtLA3xV3yNrrU8i+lHex+u3pRI
ANFEusF6GXbgEMr2xAVib2/0bGb/UTD49OiFcMWK42tJvtjxCTAkzhHW2MyzEkHB
5LbKN0F2uoMpt94HgZuEnWUdizk9hoIyRBL+XlqfvpFhQtRiQp2EwlGH8eleWUj4
on/TrajQ8qcvFyyXRlnXnUU144ZHHSNf/1rOR/R14b0DQvhOQ8D8s5ilpYRKNzvr
SMidgFgPTLpWKhWTN1B/liqT0tOEkHnkgCvyWxeEwZ/89+qd+yL0H2kVBvtBLlq0
q71YV7onwJ3wOMobbyOo9Jl7+9T55Jyy42UyVxl4l0ts532rv4doujbIwRCpxBue
bZ2cWPlZkD6XEFX+5n0lwbSDbRLVq7aT56fWHddtoY0MWRd3P3FDqQpIrxqGywiD
fuKUyl1yrGP/MLJFX9B16KxUMYgmas49heRIYEdlW/lfay9wPUSe/a2eFIhkKwAf
lwi8bRB76Y4l0e71Rx3lNz0o11e95NhZZ3HI79qX0UEFpU2mvKo3rEl/0sH8F9x9
yN0Kgac7QGHgRWxnUpYmGY/4x7gvq8F1yEpWavdtwkHNyAh6VGecsvKjzkVCWiHC
svLzmvnxQrtctPwh/I15O96WNwpDQPaN6bB1kqBZl/abQO2Egwr9VPq99ELBXA4Z
dHDHj4zNq3AAOyt4IQlTYaxyKLq72f6Z2AQp+X8vtqsjDn3FeIuGiBJnWSUsvBhC
VV07V8Gq/yrGNMYfT02IMUm4b7yPtn3UBe6t7rnwIGOG29NwYEINuZ6sAqMN65LJ
HhoTpFlHbWNm2oX6aK9kLiowuZflE4/wx1SpEJI26DZsJQJYSt4c/jklDrbabYm6
zRHZfMWiQ0ZiOVHQo09bDPSCoHg1ptUP6o8V4S6ed2r83Fwu8oMh1tpQk4gNwsau
RoAPWfRjr8YY1QO2cDTCcycQpeWOnSJHo2UV3gRZK5zCNns7zWtsiMbx4+riMX7F
GSx3b7EaNXPhSUOCN/tOSRqwX7wAp5xIQzLJRZgdBhGg1IhaOZhyQQPYvhDskPPe
16OyOSQM5lk49gKi6sK1g8JhM2xqdZkfSthfZcGdcZzq15P9k5WVtZVqqcChUXOy
oTeGJer5GOqkqkZMFzNSK/xFhJHQjnN3rfM4ZzTfP3GLxeIKw8301po/56jCRSH9
cZ1aB5iyeCbdiDTdQRLZ+RH7ouSdWTYav3xtFrNUV4b3Y6fCfQe80fhRL265XRDp
P3e0GZcw9/MCtAoSLcIGcT4iEOnBoRWeaaaS4mlTwVnx9fa98bq3JTja0lWfjZP3
ET+GJOqMK5l974FB7TxW04jNva01PB5YNCzPpZkWt7xTy8NQiL1nIGdk+NMbU5uI
T39fTXB6welgpC3u/IvUYdiwnRQf5sx4QgLlDmzsBhORCjy+9jbpf6lYC+P8EoVo
tiJXO7f6hMr8R4DwLgFqbpleE+6F9vK52JPtZlTXCeEpwjnqUK7Szk8nY6eewQC6
KnUL09VcT5UsCX9NWUP9NMuxCbbJqvO5qXfYoTuKsFfIbZsaTIbQo2iIFDeUtWp4
exfXh/PXSBXYFzKus5qq4gOKL4dF/7kVHV15CZs/A30o1iOZMi9JINgfV0crR3qu
nz/zNLCBFq9/4HqWhO+z9o11owy9duuIdQg++/vl5VOH+Kf25qxg/iU435fzZXc8
ttM7f6YksAr9ry9Lg72qMiEtl6Ykr4sXyQPPDMl5nRNaDXBMoJjkSbhobhvpRZ7+
Mxrkq6yrXSMRjIFUcVwXoSHwwdtdYhDHndTJeje2GGBtIamez4vPfAbHXIaFUy0i
C3Yk08XBndhv7IdtLnsnPM8l10Br3xTX/5nBs0VKtri7Z/dh68tRCDe20ZV+O9xQ
tIrU9G8vZ+3yEJoiXAyPVQCPbTRpIjcIkzxMi9DvSDFESpZVUDj3KG89Q6ZFvKrU
6J7AqJgEjNboqdNrJE1YUVMreaNdT8Vv0DlFWPvEeH3ITqxYIY43K04zg1aMSgVx
gY3Fw22mDrGdDCgxSY7jl8FUw0iOp4InAr5jMWTJRlQDHE6fQKoe2oozFUoY7s16
f7dnCp1EpdcaKQHKB3rpHbjziv3auq+cEje/8JXsOmcKZ4U/uSit83z/Sb/0l4TF
lXA1VWnQyaLg6HBLfScVFF/Z7/7WWFLd04qHIhrGHfOBLz+4ELQ6VLtMhmEEjtml
AuYf0qH8TSG+Y2c/qnxRGacFY3z1ab227aNqFn49u1z6cb4GkNv5ktEktSPqGwjm
viwfTQrJrSrfJLLpBMapb+kjvAt6LqLMgnxLRiQqa15zO4Y0uPKMsC/p/FX3kSjZ
uWqyaEXavzw3F2q52QF6LkrdJk56k4sfDTjrQaJXkOIDybShBAyam+yy/jkm2+zi
hh6TqRDC01myFLtjPgKP1chJGRV/jBscg8tuQb8bCJaq2k/I/gTmPrt1VQ4d/3id
+kxqYlq67/6/SXH7PjbSrQFRVs1A/U785X1RZFq7njDRnVKuBWGULMrqjYYq8dwi
C+2PaVqlWd+kGnt1pwL0rOOWzpI7sva6+l+TqqYaKtI+nLLMG0/2ES6rPMHLyphl
lSGXtDXPqheLpcK/Ez00yKcTPA4+IXtfyRarzdxzhnKV7e5lrKyNoimWQFxdEgOD
o4+gjguU/UnK0yncBTQmS/eDPVwoAYyyUBcs/iYrPueEVRXodZVy68+JoNSnF11h
zdkeSVGtTe7LvqkK9UDC2DZ5Xmkx2slfEHRufCFef192y8MClbC7b8Q//XTEg1da
vPycsCTJH8pvdE7fV7WkioTlCWU22G1ziKqw9EPyJ6Aei2Mewq3Wcsh2TSUTEInC
foWw2aOtigHVIVSqRLx+q98fa81VU1pustKwBbzjPK9plCbq1pngLCBMbNgFNicr
qkN0uF7KLKZWukGgWPGs+2reM5hpeEDTENihiksqZWVQvko9fv4+Vd78BHeoepfF
r2zfALdoajMJarH0nV9Ya2qeAJZENVi7MI+vRRaQp8+RFapki2Mbd2sYns09zHAZ
n7R2j6GQ2Jgss+/SbemGP5kM4/1WLMnxBHNxKhUoungk/pV1epXumFpNjLuBJAyw
CY2rX30lLK88hZ4nO63Slh09qiqr1rtOl8rMbvyZTv8Ine0FEJN4drlSHr6LjnJP
BcFNnkFbm5thRVR/aAYC+8bY9IxCXKzJqOlqq9snhy/lRtJ8UKopMe05Y5mEwG62
GAwsVSc7bA/2XBrFszgIZvIbIMg7PUg4KfhsupFDdr/EW9VnJLr3itWnfFb0DGlz
5jlb1flAUYXjqo1K9mTJE6wc1M4dixly0dOMK9kP6vi9rCpI5B7MRXLDbbb/s39L
QlKhIQdHUFbFgLiVBilNJVk1ryUc/kSpHMQ/0/U7/NJlidl+bsRVYVOpQXO4v1pU
0ufhngWZcfKm+nGAKrP0OO8VPqo8Atjdb932ahihygtANvmta4mY7Ehw4irib5TZ
VyP4g3S92Cz4LVKZIyfvxuL0Zq9+FjwnlKlXXabNpbUymu76NxaX6Sgo1uNOGRhd
nQkMX9+n4h6Pyn+btLe0k182PgJlLgsdAYSC0i3f7UIVkxsGZYMP95c0TrZ5luzL
vJh89ETbp6iIf9Mo9+n4Rrbm2cjfzQu2VIovVWJOIRpbPzaMEnWIgFpM8hS59FTr
7XsArHLZ2ruP5oZm/SaPqJI/nlcr6y2vW6lOARkC1f5BsyN30PKm9+LBx2/+zf9f
Cl6eNJxv/lJNz+DVwCD981v2HNLQfuiPFHTbJGcNaG6cTk06cu0KEdHsaog+ZOaU
p1UIO57ZoIip6fI5l6Fezt0XyDrEDpWiI9ovwmQ41bSOFBtk1vpuBH+1zBJeezKv
o07+XLgLZVf5WEHzD6i5RA6tWV7oP/XxS1XhUGNAQK9MV6p6ci97PXj0rbKoBrnD
I7PucxCTM/CVT+4fHk9C7ID5jeFCHPsZrbXzWenfMukVQFSV0W8G2nSmJklVcp7S
ePbs3Bt9WlOVBB8MBCu8DcWvo3H0GStxaSotSbjkrqCh8G9CsM4wMHfUkyIPGUR9
YJPB4ZnWRxo4FqEEXJ10cK2zc4i5EUCka46OJqa4U82bE+wHolXPC2DPAvX/eaQB
UbyfXfaxCXVqFamA/H90xcXpxZ/oUZp9nR+cK19iPWJVJchsWhcwKi6B7reU2hMx
gNUaM9bamvFOkScn/+jKfuYdiFcX0n+aNvNfcio+o/J55WVWMhri9rXsXUQDwfAo
gssZDb7oTbLgR0/g9NGStIIRqZoiAnTRlwpfUY6PRzUtEZbSseXhi0SqSDQGHckI
MMjFOPd7qW+tNawYhx4srHwiojxhSwkOa4gKHDIfDJ2L5eLIMjts0G7T6YN+8Wp4
DdrgGASvOH5zk6/4UhfKDxdP78vHf3c7xwhlzUhupsU91nQrCqPGtgciRs5go4wo
hrYUWRgy+5usqLcxYoi8j9Es8b3ESADWpU4ccaerDdJl30dozOvjbvxiq/wpbNPN
2wZHvcLwOhcepsmJH9pyaQoBi3BTr84VnXHmyuoDIxjTCsBZmKJKRDI0vrxL1vP3
fAgr4+hvZOlAHS7xdttNSzAqs/vKvUnNQAiMHANecwCe8U/muUn2ppVZNRmSzvRn
cxUQdQ2TgjUMOMjDYKqLq7fqLCti6xDahVDpmm87jSY2dnp6Q66XEiVeuApg8NBi
+zbwBWGEs3F4Ky2G5Y38WabwTmK6Wu7FDqo7UNtxxIyBdG3Fa+zojjBxMDDROc4v
dQAimTQJJewXD/D/UlChK8AndRiePdkyVlXKcJyalXsC0N82JDXMnxWkhPn7hha9
wIGBaVLGJH6uxzpXXQJmJEnc3INZukKO8TttXjFN9m668SmJFe4/MlYKrEJEmV2g
rUECqST6kIyTDc5jduhmd3g6BAtW9Vr7/9K48AfqAbOCmmnXLe6Z6JWdO5rj9pVC
bnhlu6Dx2/IUwiwisF9Vxx3mryuipXW36xZ6hNjLhdA/skdhVnT3y323+zqZNxTh
95nwz1gbSD5We+iTuVoZEbpQYixqBb1Od0mTQk2IpMn4MV9pdMCUU+Y1HF3q3lzu
0OUFSM2mtg4YFK2VZyrTNMrzASV1qYa41O7NRlySpF8zxUCKEwk6iBj0mWKrGuKb
iqhIKdl5GPqCFoB/cWhokaf3m/BNeDVKjTew139Jc/yKxyzuG1XJ7fQFZgbR2vOD
AeLiMPxRnCHGnX/IH4YLdEX71rsFEVzP5VSCdNtch7n49RX/ErVnizP9OQIc3OrK
ruRolUdGgS8OaeJEpsoB8oON2iWByeGTeibtDai6PQQFFqi+bATipS9pbWTiQUdj
7IRQYI0Y6xMCMP96YS0EDQgJWiFgk3IAO+McH/Q424mYrusdygHnW6Q/LwnA6Con
8wss3w6n72B7WEeMy18JR2zCFXhvye9jldDC8uleu9d+SrfXPLATGdHNY9OlgPm/
AH8fBNuqH22TD7ky6e3WDI9R6nYyAv0JpZ6nZtrmIFIBKUW7OTvAHdgeWhHJQTfy
oAukykiy1AjlHPSiHFTypv3ZlbqQtwOru8Da0N5j359Z3i2xb90Ij2S+bomYnFxt
mcK7zxrRuMHjDF48pZr71oVUm0/ML14zn1XlO22WScXZ/gw2FSsawEvC4CpVKwwO
8K0lUWBYsIE+6qhXFlsmnT96oL5LgNOdeQbKTJdyrj7dT24FCzdTFCS/Zgo4Uklx
MHp56GRIBSbVPDHASwAV4nIknFixSN8EV4s/NQe2JgfvDohhn6fyuxSIdEe0L/EA
NsGK33PYxT5U4a7KepHTvK9KuJ63hcEg3d0j+XYVGXzBOE2GXqO+DoPk0X7msy25
4qlJTkfpVbnXxSkxzPWKDIwpwDI6MtuxeIuyRiuUqpWZeA95QxCW0At/6BCLYDld
YZLmeWi8OqqGk+kmlMFHdHNaZlBR1KfJ1exsRvD4xVCC6p6OBOsCFCELYrAPlfsv
ESZ0dufQMviScv3zFh7mpouH0injZrCb/+ArJE7qHUk6Oh6OA/Lx2RVzhCcXrAwE
K3DdsnjiKWrJEZENcIy/3boHj3ESBy25JS8pRfJYR/Fmo+BUH1OrgiWdEhxzoWFP
KEn7lfuYCuZp3DTW+75LddK2jHwA9/bOHI0w6dRTmdYYldafUFQCFWE6D66Xaawc
5thv+9vGrv9OZhVzVILCfH0DYy0Ii+ruqaW84t8FAlANt8vup+iOr8mAjgsnI8aK
Ehox2cwKpIL69V7Gug+L/2CW0Sngnd22uSEe2V2iaapnmFjsmZrqvLjcPhvy92EP
5MGNEIHJlLBfrO+zCO7ZOGg36crDh5z1WlpjQLStI+8cCCORmUAO1Gd2c2QLahY/
UKUiOQkG9LI+3Ec4992gxkTuSvVTJoXFWjjGxPqmKij1uCcHaOkLFndvtTEAWqHV
sc9HU7HSI4MHH7nEb75g/Tg1iqxkP/YwQmOhgd913cvIn0m0LDR/OlUtG6+wIjud
S+rnecELjb3L2kPTSenXSTAD4MWyrLtO3D7IOzse1FiSEph+HsKOiCnHA1VpzzP+
wy/7R3xny5F6RHqUgDxQpDyia2p0aFsYxaizh62mdrp3XCxit2rGJZnBdoW2vo5R
yQOjrSpsdpFfZs6vTDEw7s6z42lpesnXuMqXHgJjAa5MNooSSPuG/S/AMilIagMF
6RA/qxqhk+Hbhg1Au4XIg/nsl/lIPmdFhHhRHKBr5s1AYPwDWwHYtpKIEY96z38s
WBvYER0K0wwIWjUeH9nV8gCD21G/aWWcTQ2c1QjC1DnGL3CTAaDdmMjEVDLCncHA
giPhm9G2bgxAjzaEc4HVq3wxwq+Oj6yHbZo4hQY6BZX0pVoP4TBJPJP8IQYahnUO
Q04bkCYXlHcu60P215P6tOeBRAwzrymDS1ufI2KH5dsTQubn/p9Qo3BsRc+SCHCQ
jPQK7QlolmBe0CX2KGwnVFN1mfHXAJTdgdh6XzKPvlZmCN9iL/nklxxeemeRIZQS
nOXZ6WaU4b0I6nnPuNC5UGLeAd9avFOsNgf8tutBmyClPb1c8zLGIGOWTLlDS5Dy
Xt+x7cxJyDiWqzk5m4BpVRytfIJIcgl1HiAUjhYQm0isWg4iCG8vcTnV2v+I+eW/
CZwXh1aIJQ8FGaoGoFGb+Ngq3qihdKlXAIs9RhvfXaEZHdXYnLJmjRP+qwUSkXT+
9vvkLfsnAC982wPewL65KwoddKgdt0Qbhffs7usOJPe44dkd6GX7AW5VQq/zNxyp
l0mkq9IIPv31KYOAXVzwfjpfXYz8YkUpDSVP+mFtXQkwRGyJcQEzK9p6IaugBvUR
a9PRmi7mN0XE8OD50ixK2Bq7COzxiqynQun4EOqBPnyveR4y6Iq/zYegFDYjeJRq
EhFn6hcdUSQFosOAlc/HdVudjSUdqljY0tAtduj7zRPub6Spo9zhf2x5rfOP4qWo
GfgodC9ZcNpL7+09MG0s/+4jAazNRZFNW5JawlxoPhM2uHRcNk1qMKRWbr1k3JkI
rJWDMnEmgzi7ad5yHekRLaZ4oXtBC8o3L0uJuybupmz42wPdi1a0RatsbVmkQvEt
rV1L0yp/KrqE0H20IoMMBz35Rydk+Wqiopdf/Cz9/7Re+uSjTT/1bJS19nF3J+Pb
O/rCPZ1rpzAFGzUhnB/rwB7pCyK9UAaHnQYjnkWpvPrlVyavVmOp0qN5o/iSeWpq
jCv4bcH8NywjBBU5WxTfRkJCJ6oPkQjs1c4q/mBanLsBvs1EPE6aHEv6NRP0X1SQ
g1ksTuxUcZ6wJSnxxlQYCm1vdnvJ3QPDiMLPVTn6QwECu+HxmiC4XkVAgUCZbJOj
fol6l++ZDMc9FQPUfyiWcQd6o+5ZNAoG7KtVn400Nt7OY9TeVPYhQOYx2SJ9EhMH
pnbBIJU3DoEqoPlW8XX8sun5czcbt1vGIvi8AR3G6cUiH0N6+J572SsDCaq1ukME
KjwjPjCCclbMyC3q84r1M/0kloJAKGuW8QanRUmrovS/kCdgeTXFPNk+LK5SHA9Y
rq08SEs94i4aOafqa9mJd0zkm417DJng8WRmbWd0+A033QwDTz3obc88A5kSGnD9
PhTyBNTexKdGIB4VMAt3DonEus1wt7eaVkBFsHAXRrfbr08sgl7hvrwcoqgLKAw6
oQseejBx0grljCCscNvsP2Zi6eke2M7HfMW0SAyiZ4W2c7n67xwbG8B9cQ559JVN
CU3hQwqniDb8CbNtrETqiiJcHqofzoBpjPHkp0M0jFtsLObW3qcIPCoMXMB9EeNo
94KUIu3st2VSHGlLdbtXxHte+Qnr3qJofFUYEmJ91W9SJA61tW8muJNd8RqVklOv
gaUNJMAyzKgde+AaTtMXRQFzH4PyEXhXMF49koQi3QOLkQOMYOle8FN9KpnhV0RV
Z02C1LbGIdAzb4aHl5lBZSbw5SorEeVP7JrqXSnSli+Z7CiM27Bk8t4L0VLyUHNp
5bugexkiFjJGdu6ut4KzOmJYQ+7MuGViosniPcV4yQ75Ln4sFi0AmwyPQITd5Bv5
NEY48XjC+XX02v/3omzVSmCCI0cNT5Gw7AC6uiCu+gLCDIuClO8DPFVgmDVnp9wS
+62SMyeRsToPYu94FIo+fBNLApIVdR+wsNpzOnYrDHHLgqv0Ue7OMn15BqSOLnoq
AVTRbEWrIc33R85GEMA9Hn7+g4E6br0H/CD3klEvo3Hxt6rayp8oBZmUeL8aoHCU
ihCFoA1+Riq+SAUzLYCw+5oTxC0yUt8X1VEHx/EvuRltzyrv6wM4E2E2AzOKW982
E4Q2hLMSFk44YCHbc3Au6tvAgckkR2MlBFJIrNJJC5/AiCu+Q+ben7KZ2vb5B/XV
xYDJCIdBLldAwx45R3Lj+wcm/tshXujtUq1eXIxkyf8gHheYvI/7zEFXy/Bcfv2z
tlfCtJJnk5OXZA4bRqjNBO7yY3YQ4w8g18gVk0MDiG5T9vpZs8RNjDZF71sqonlz
7FIbao0PnhA68JgHyy4VdsL3kVAQWwHyiqYsOGB58bFZ323ZkVxVAfJezyWAE2jg
/p7vLjISwkwqHyCi3G7XTUYEqk56ZRMVQn1rtRh7lyiI+B+fQE2dlfc6mrUYca35
g3iYfaBQUnqIabTtE+DxTQdZuP/sZMYzbZ0r89snrNd5oy8r/9RSbjtDZdqrEkTO
e9/fGknXiWXYYmvCEGsqWafJppoDJyU6tlsJP9+eQ01xxrclFFrPDL2d/aJkA/mq
5SgH7dGe2Rs7/rIoKCMS1Vr6kgWOYc8/bab72ds28G2ddoiNo1yKD0nnVktAkg4W
TdAoOR8kzzCo6pfLq1LKBbIvIrzNXlq05ixjv+s1OK9BJkOlrQ5mtiuWISa7kQpA
WPwf96WwYkm9qv2n6l6qXFWj3L0oGkBKsPXkwZrjBUN7lg4a1qBbj87yTZaFt75t
uzrHOlcZvM46KDoHpuqT56cdkPmACRadSvEpAi5z4m4LSfVmrQ1Ig/ukeC5uRTQY
hcp1paDsMQJr6zbUusGgtqlkARAScA6Gkg/k3OoLQcvtdUzQZegJ7s+pWr/D0Cfn
aLSYOjVjEZZwiFf0ruTnvF9j0UWGeIohWRIR1dxA0F5UTSbc3jluyqnHBPjwe0qY
aNwfiGuXiWSy1Qp2uS5F6GM+I7GSfL6OAtvrf3aHZo6rXboZKsA+GecOe6wlg3uM
NzNuWjIr2vUCHCFvfq1cHasACKsd2H3XWZU/kqOm4jmnrJ6RaPchr38iOHsI4YaF
LdLKyr6/9EGLVgQ+9DJ37ybDUIzvck2AK8CyrMUlLdHgSvMem2dv5U4gIBsU8BBl
TbkVyZuYN3DgSF3049qjuenlOtuIMz79fPs99dXBoQQnZ4YSWZtcM2hLqlkmG5LC
80QmJmLOwZF1ZLU9VGd5mgs0vhMdSS7lhCEZALZOJfUjI0zJFx1vp8lfNsopVztB
v47jJPXaIMxtSdFDKvmx8epnQGymrL7ZOD8SvVcmZmjzHZHfUJQIw92rehqepFaN
kj7AVfPe8GM1NYGGqQnGoEfkRIekehpf9uPi3kbfk84vqOnTSL2U+ejukvl+EmeO
yQAnzWlFmPtzmlHX9qMOphbQ451g/Yn/USsEhy3s6HqhSAqKzoc87oRF88CLKl/9
mBlTY5isEmyx9wZYjuv62EeSTaMr+CTxtGMUtDCYJBrZ8cIKgZne+nLVdjazH5WI
p18TS8stn0s3PaCpiIBaHxCApSOqrL1iowouKLbmL8QMEhmyXsOunUJtUVHGEnmD
0X4DHygOBqqqBYRK6TlturBOi8Sju7xeAKGD/kkUdthQ+nDVNdwBU4LTazR0yPH2
7VsSDM9gGyvegnP+eOtHVjbCCNEhyx4chfiWoFFtgTl/iV1BQCKGz4eU4LxT1R0m
Uz6LqXlQabfPtFdg8cxWGdIcfbIcz903YEy2B/CcPmL95Vl3cii2KfulatBIUNXS
aYZHhWnxxMUmBicqtu2LoyMA2JIx602/nLcEyuRYpKsvqwJ6ZF/P1e0S0qy7yrQ+
Cwq0GMShNPoI4gtgdMZm9TWUGHUllFwNHHM/0V9llpLg6wEyUHB0uaJTDqyqbWwt
DaV3spEsYS0x9vQu6wa3UdfzE7pWfw6alwggg7F6Sfr1g3JNrVHONzqIKC02kOJn
l6r4KjS8CS1cp5clcyz2Ud9Y1POi77i0y/yBiFAg1dg1DSD8jroDj6jRl9xsQR8S
oM4vjciyjkUj5ivtT3vtb/J0iGyhvmZlq3mMJoWdEVG2OjkMMZimY2QWS6IfG6JO
cuZUCXrc8YoIiv7K5mbP1BGY5GcY0lgocAtLjqB3kKDmS1+Vxfq4tyuHGxykICRH
Q74f9jUqGypgpu0946TPPQ0CG8s0AAxGnqWYHA3bwNn2ZgXWG1J15hptNw0ELgSS
b2ODm8+5XD/P7l6UehaVPdzESqwNy62lZHln97o9RY1lPntordxFF0OraZ/By9Xr
6fI7iHqAU4PYf9smPwA/M9UnyMEzjzncR46T/kHOtugBFcEX2rGlfYEidp8IT2RN
UAQEJE7QvYmJTxe9MzhaEA8dhIaVYDTqOrXRGDFbjdJwXHkvQt4q/kMT1rYGj+bd
siVqo6IteWuBaiBUfHNmYYjv5f3tMRoHsp49W0hNdolRliRCqgwQcjWQgfXSSLfV
N8zfBOzJC60nKse7X9f5qoIGwMGEaf/gXr8BYs3Cx7eDOtRCILuSYaIJ34Zrxo42
S779iPk8j7Ggx0OWAUw4/3d4KZ/4a2fP7zObaf+74Sxh3A8m3JBQWaAi7DQn9OWi
QzzzfKoWllcTXSlgFKuBtyM93ti7LR6BBn6sp+dROYeSmRYhqerCS7ZQf+KDhh8O
tYCRGLhKOsq0dwqN63DTOTC2yUp0esTItl3fnLuMQw0ht7Aw9ji6SIxktEsrg4NL
wtBaR/EntGsjBa4my6yxNBUw2uhUyg4kYQQZFLsC3Gts5Vcfpsg532gJgqqLjrMj
hXYsUqkRJ0TYxNzojMW1cqwJbuy+pyjOtJwvXsFBGp7ct5W/xyoobKN6OMpTlyfk
9vN+61HnaPl4UBQlQhjRVGPHR2mlyk748VNGL4Cjx/3JdO4XabdgfwvAz9r6q3Bx
z0kp7mzY/4b620shMRi/2vd872ZXF8xcpXv9E+lu0ttE5QF0piUAoCwsE8LyybJ4
ISjN748jHLszAJ9QH99at2K9lhhhYTiEiq63+btCRbprhdfj4PsRgZ/BiERY5nqG
X+afLOvK2hQaMRY+9iZ+ElYntGN8F6tak5DqSTA65BbZfCI99q6rJn9t7Ne8zZDN
c1Uvxl3MlztJfDxv6lfs/Lo51vum5O16I9Bx1wWAb+0TYY20VkcLLJsqKxkU4EK7
XbHtL01J82pPDX+tlPmt9v6CFD2V22olaal2S6V6mZqI5fsUqNK+39KKjG4ezPJ4
TsCUql2bgGgaaBm7g+sIjXpk0cNWZUQx2NRt36ayfi9j3z5Bgw0YwAPsO/8NSXe+
/LTOLtj9kHppzzmsDrmA8CjLMwP07+ngIWvP/MhcZ4shhE4UTsz1hOUa5A7n1N8c
5xeIdxFA4I9htlt1Q62YhxjDwN5sOeR25eBXgCxW0w4zI84XAhcXiWASs0iB/QQ/
S+5dWpxtLew7wHbOWX+6RUKnbGqU6NXmGWCRgz5gY6MJtT6DdDoqKHNq2jGvVziR
uFVGsvF/ypfityf3PBq1NG0zDxZULSjV2bo/20nr7u5T4jVfcW8KGqlHtBFOX2Yt
dtIaTyCE3YTccIrbBKElnaeXij+WRrqnHgGaVSKCDd1U+zarEQsL4mNgPyH+ffR+
XjhyJtDj4AZQR2pvb6w0BjNiOBYRznwdthY+55QC6n3MvQ6syYAb9r2NvB6mASYf
+58he/3vu7pSJ7b2EX6fDawW2nTULjGmPrib4+MAPB3d1O0wqTpxr+5jWRHQRRIo
yq5vUxIoYfGjbTOZ51adk0iawxQusWQCiyNQPG7TntSA3aL9bNhwWN9giNZ6CI2h
s9gsVMIt8C6K3PMG/4PixZz7B1i5mnf31MhfZdMDY9bzpGqTo6HBvZpf18qk7JSY
jPM1yuzDwqQ/P9+pOkbdjIFXYtqRz2ZyOdq90lkgQnuqhcjBzi9Z6Yh+CitJjgjU
MKxNDL1/f7MgYL4sO50vTRL8iu1MvOii9AMfIZ/bTxjnZTwDaDFZ2duV6CbZHDTB
yLPtKTjWQOPcHEFJQyLoG2YOS+3res+JuITpiI6aia91biLhaxyCcGSceX+pX1yG
70VI2uhpJQDuAHagSCi0hxF4hVTFYaQq1uU2UpjxFBy6lMzmxibgYSATQ/0r4TH0
1HOXzgGaJBhasuyZA08IroA/cCHTk7XYB26jzmZ4YXKqtBpjljHxk3TvdOFXpMOP
eASIrbFffXKdgzJXDuUdgazg+B6QrRPh+zJts1wA2OFB2AP2CuF0MSoIEJRvCiRM
vs8e76Rw2Ii11KbTv7GsYczeucJzyR213MJmmdOt+0xfu48ZoFuMG8X5Kjc60sXZ
VLzmyYWM5HdOxQtu4wGsOk3nkFGix+TYeuWJodDiuwuUl9iLI9njaev2TFaYKuKg
9b0/rbMGhcVbbg8R7ZtAJB9DD12+TntgA+tFQP9cj6398OMUvlF6bRB8/X45vuvI
GI6jItzMKW4yEHukIPn50JVcJyH7kdVOyCNo/k8rqX6SZ0XguoI0818AJE8XfMJY
EZQA+OUs/EVIRq1KCBxHDeGJQeV5Lamy8eLck7U9a8Lx3Vie44uN25vBlFkviAEk
6Nz2iAObdRzuwdGhNTAR6H+QTIb9jnRAKJr3t/jEqZI3nH96ehDOPydFbRvi0v+B
ZkiHcIjJURCUoeAAIg0ctyA7Q5vdYJesG8jnYYmrMGMzqcMeDyG78tiVx8qNw1DO
5++naJLfPDrxC7wRafM4WHsi+jM+28wIUHCElF6sJIzxreWHvYwJVOU1p9Dm9McJ
KD190wrKA/0ltrYmZx0weoyJK6LtkYFGCXghE+SDSwNLObK6WHpnLu+jiagTivp1
sbjY2kIMS7m02PZop5SsEGliHWvX296pmIGm3o8Z2o5dYN4LscsJesr6q92aa1nb
gf4tzPlBVmKLdMRUwyaSqtTl7zArvRoA1W58EEyuvWvbBPL3Qg85+T++sZXAgmR2
6H7D8IRe/NuqSMOhDNVe6LZCje9K3FdktGcm2vNY5q1ibYmQ+sjwxrD8AZOv19d7
bW90TXu4h0pc7F1vdEZGXZZuqSPvjCxPMKbDvG/a4ntJ1KZAzzQV3RM/4m1QNriV
geFe0gB8jVDdmVtaWDabZuxoYNEzgekG8tbI1cwZ32L6z22jcOBbJdMN6YsKowHp
XognnErq91MldJpEGF+SeOnQTsGufwVwVUWfriSmo0dPDZsX8UZwA+Cg0FHmqgqv
3rIzpOJwCTTOe3aI30PcC5PD1LhXhqEtZAHSWmMRiG375ozKUrTAI+y67LK2y6BS
p23jSpMFk6jzfaDuqFitt0buAd7Qcf0D3VKxNIthwEzjfREUOVYQ+GiRq0DRLif2
Tta+HMHABC2gjPbJR35eR/vrVEY9V189dyRu8rTPPTVpQVRR+xAoh715ec0nBBHw
nOamcESSweV5hIRGy9jo8l9FbuY4jt/bwGviv+tqCoaxm9Qnb330/TZGZYCAMZyC
Zlt+bZ6Usswased614eNGFXoWrot8qHuYrLYFgrJJaS9i2+M0ce+eesgjDs0BDOd
N54Ar/26uwqGSLxu9p2czCmAOD2C3b1KsiVgjwQFYgkTH7pZtH5iAyUU6ytU1O+k
ClSMxyCb3fDHVkQNoHqWKdAysHeUd0zlvb0GuAJYDyGLW0zwmEOtJWXq1oLPxxHc
gEbfBNGoFxhQE7CzUIYNP/yi4vLStZIDKolafH3RsggYnEtGv5XjMyJ7W6nC/fp8
PHLmSCnwNMgW2+2eC0c4ksv5SNq/Gc1OIonlswAwirxMyyFoiP4VGZTBg8IDdKmZ
cZYK9m+yZyt1nf1SwAhU+Qz4zZR1muXZLh8U4fplsH5pMIn8288TpAOb75oBx9Ok
GoD+Y4xyluQwhkctimEqcBenTE5JOvWNu2FgIekM6osUBMQm7fzdTkkYVVoeSZha
q+E1bqhMdAIcrnQmCXrJMv/3z2VBkZAf0tV4G+bOsOlI+5Eo8n/mCZgjQ7YiDAOm
oPhtkKf7W+E1fRR0SxZpVAbKKIhgS6zMhAi/HgKjdgEJXtkgtlCgp7Fun9ml+TSZ
wkd42nuVVtgOLRkSe2CYEFY844ffInV7tNRlb3VLRyPmch0+hcPVc15+sgnrjFmC
TIx/ZVwPF/Z9jCu3MPMJYm6NEubKzm1WPEr2/7UpWpQ+3N8lV7U3+Eo6USG/X45b
wo47PqDQg1C089koYNw3e/U+xfFuKT63WWspPsEgUR8y+669ZblrKlZDq4rOHyQx
4ECtvAuPqeEI02Ny9DkXg91SlV+v7rc5mZRguXEWyuEfRUnPDYyfOVJYes8tQBPb
orJDeVDPIGMLKACM/FVTk+qeKvhirnppGA3DG+Zgofc32xsc9umzThT/zwOr0xb0
SmIqfOIOgH0zYCyEcNsmVtA4TIhqlsYTcfpdQJETeAnFe2RPV5wTJXQy+HBXPM4y
JFl2sTPC6MomH77bfmtzDd2RnEVh+cfpfYlYl5RfFFowMBk8Cr+4EmVHmVh7kiga
tZ0ATEXleSO+b698bZUiQeYN+AVy21CyfQdQyOkh51tZAVnFyBaTFc1Nxfx8Hwfo
2HuSxdIxaDIl35/wvNZwvpcbFZI/BnFFrc/7eXYr+k8+qhtlBRi2pYyASPpy2kv/
sL0SU43OV8v2cXrvdUDXlMbLtytmYs6GlVdu2yW5v+TVnkt/w6zqsxzxkvS6cgKz
hCym48wGk0W63yzdyVJtW2aq+JqCvPJb56J1Vzh3ahCTvB9Mw5es/aePZWfebMz7
6O/YY+YIE30FtpUCGSznmUOmJnVpXm5Y+goHag5vex5vDSLjarqtTrI+KtuFee5D
34OpL+u6OoJwM6WByw9MAD4DDqZBAHQi9JMoTdpjmMoGSBJXcVSn+n55xVGrZgsW
LEVKXtsQfmvzBbvyxYITRk+OWUkNL4JxFzyWPVKrqqFC7m65jJt8+rhbyXB6k/IP
knxH4/pRhSQHBQM8Uk4WUaZlHFYqPXsGG9i2Jw7SbB5/MciGzZWfLne/yC1L4mYZ
XXLQ4cKm3o8KKJuzZVPDA4ZlcpXpD/Wx0760HenLQRY0VSbuhzyDHIz1THbnVEKB
Y3EgpJMJht9xrTqFvithewayp/SeLSrJqazhpKFwTwa/dQLlpiwEeSWO+thlK1Sy
cV2lcJVYIfYiErIHx55BIvfksk9jQ4Gdoa8UAcA/+yehJ3mggLMENP8QiCinNJho
O9ei7pTw+neK6r845YRG7OMEPv1U30JteVKPF4zxbNQ=
`protect END_PROTECTED
