`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26HDBGUdPf1KkkDN1d6amdvcZRon+5BktLqvLRY7cJaG2OJoBo8mNC7DVhXHZEuK
n4xEC2nPWcNhYMyZm/E5AhCRedso8v7Dwd7LRyRdgb9AB+Zo288Ys4kAYxdA59l9
EwFreu9vmLcO59v1Kk4hFNdtqN/dquff4NAwk9VBBQKNnqlvZcmw6nln3b6/Rets
Z4uW1appfPYc5ICtw2uID4K+bpjPw/qDZDf0PgeLconB/IOl6bZKF9oAx4366BFO
eG30oPhxL3K7idbOl/IiTZNSBt+z56h2dRkhiTMEDNZyOBfRxlj0403WjABWEXCi
TOeGTljK2YOe71nFOZXJ05zRice19mp94Wb1AHTbd0B9No7TUZ6jSvs67YWN7Xf6
JZ8AYIhTaymSf2ssazxLQbhRDAGg5v4pZao1uozOkn99i7pqccivNwPPkV60nEqq
Lr7OW0mI63BNncgYDExK/Djphl79T+UxV3HWnjvj7sallY+SVIcyyfcmkOGBjnpr
4jpgqeCZTezS4aklA6jdKWRB+FCyZOc7S7oMX2A97axJbhrMNrIdPECj2P0vr1lk
Hs2UZOyGYrD2UxdDjfleVamhHQHh2UOZeIT/YAIeuWFPGk/ag9fh/DpNb7kOx9B8
bHirEkC7bJ+qMUYonTbHoE7k3DJpeaSYNDZ4pdMGO5U2gu6KOoktfAXmUsInSS6E
BnRE8kAxx/Du9ULn+YuKGHtugHH1Lmp5QaOOrxL8eNY=
`protect END_PROTECTED
