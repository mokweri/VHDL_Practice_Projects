`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyRSgI4DL3SHKaCDOBuyammgIPuKdoeFL3A9cW+vt0tT2dxO5cYnt5x4CJF7boPa
UdvQSvOcy35pKlPnus5jNQbOARmHebgzh+1yWhmHh589twPRNkGOpiGfTzYHqHpv
U/aNyLpdhVVa2VrnfM6Ys42r3q9s02Soo4o8P7NsESmhi8Q1d3rEUNpNNlO1u3TH
8Jc0rtonJiWziWVsGxd7bXYeSIu/ZigJOI8C8I7KdD/IERqcA+pMBJ7451fb+Z9O
XV+rO8XeWEJzxzeCkSWMeImadDGr92YNdB66DSNH7NGpK2qdAXlQh5FtHk8wLKsG
7rfd7OFEijNWMjWYf9pa3cqh21QbF1Nx0HQY68ASA/ajisWg6By4iP4gHVSt5Kin
tjPbVWolZVk9h+1Z/NVTc1ytkOAkJghWe1BpKmTx2QYMmNrD2Km0/kWLsUncwtkd
aiPOXzqoCocuRWh2/JBQg0UKYGcsF/KnuD3m5d0uhypAXSPbCj5ua+7kxfaEKpFm
vF84aGfo9OxgqcXRpdgqdKKFkyAzKg1Et5vqWDuuwcrk9DeOvSWZu30QumDVzlta
rYB24qfLznkOBEe4bEcs3xWZKdzpMdOnTSrb90fS7PJLg2gxgS7DVhP/EwM50Yny
025tkok9Q0njZ8TkblXZRjfRldYPRDfk8Ng2eJ6DyuJ3YFRQOIwlnOnnXiETfm/p
zptzGHkvH5MmjpMBfhaoO0bGEUTyIn+8WVWcA5DtbWcCM1gOJeIr7hd0QKqq1puX
gopPgnSO4I4ORS7a1iI6iMC8M14nimsVyDjYJteLgJpTADQJDuBqtYmlrepQDS/k
ncwosCZ3zNXwxBAMLieD+rqVX7paEiS1T3FD/2dgns6TlUQasAl9hImnPx72xQdS
k+hEVZaOmqIGOalzrTpyAMTMSbJeuuMftp3UBvuxHcaN8l7z1ws3qX79XS8N16If
Dmok59QeOX6WAdV4tJGsxW84EfdfhX/4/pSc3PKJeyFSgvHPIfXKH511s0ZDZBfU
6ct1N5umRDM3vB6hvsx0npd8gktip9eXI17YXbw7IPmqE+mkk0i8FGB7ROWztCxI
CpWt0AYjG6fUdopL/sAi7yw5L1TpXQkgps7VXOSVi0reMx77aECEjwsg2Ql7IZ/F
7QdZgDR53jOzoOBEVrOIrDwZgUHwivqB59drR5n7oUq9lqKndsvdh0bRYUyAZ1ht
VDFFG9GHAktiSwm2BDA5aOt/QuMKFSAhisaDCWTi5UTK+3ltjdqDOp+XpL5ikSiU
iMIpWuejvcKR3E/IO36+q6N9Gn37zk9G4dsE/FrAEbgDcWLHVHgF8oFOUar6Y4qe
hNUmcGMVmFFBh5dY4G4d2tZqT1Vy5+rAEnQIR38zGn3Mm7PaL3ktEF3dm3VH27lt
55yP/0GvOFIv2EAa/51n+7x0FSTSqsUPv3//eZxn4Tdap8B3NYndVyuWP9ZjeEsX
+16WJl/JG4pqyKq4UySzOBxwPNssEwsHE5kbwjcnwFJYFmOt2CpB7XrKX1TBLPvE
O9/WMlFJb0lO1UH9rz9x+EHDiFOLxo7e/C5FO2A+hmxjWeCbQJxq7pLuCaQz0BOB
1WhjJuWZaOcAEG6vFWzDBjEvuMDAaF6YzWkt1md2gi+0Fn+h6sx6HxgQln3XHv+C
q29wq2AMtqWyYMdqWHnO0CaNljgHBfdtXuWsYFMWEG+6jAgcRqyO4YfcI51g79Fk
DPum2UfbF/YhtLPdX+PQwoQ7KSfWJXf8cxuP1YNkgJ4mqW9WySkeyc7QoQ7iCq5w
qg8O+D83NmygCL411GnFIS5LdqD05I6CPIXUTlXv+IHS/MybXbKP40odODgp/FgP
0tLTI/BbrILCnEuYaX1TMJNZ7d2Tqjen7h6zRx3ogwV9yeg2y84vlnuq4m39xBSc
M/xv/Ay8KJmhid7oyIvunEm9LJlJeDJf4Gsh6TbiHhr0VESO3/lmhrC4PbEKqIjv
CqRmwkyTgDYJ8Q6mkIAEiyYwQeiPOAK3R7RoUcjRhXkUmafORcGfeUHGszBSOVEj
MkTCFylwrova7OrdzxES5mCV4KVLAJ/LbbjX3S7Ck9exqhOUJbeHV/pN7IJK1Tbe
pXPEP/nwASwLEFBdhhdkYKqx9KdR5mJCQ6nwb10SH3igM2Xcs6GKBpHeAN6spF2Y
vQ/wycsTr3dQ8kLQcwPVWC8WJboOhLn1Wj/Nu2FmUMIWl/YLnjTVuisrtg5qESZ4
dOGoh7tqhToRMa/01Bkf75axuzy0EnQwByhNXNqk0FR3/cXdz7Iwa/tEUeGKoF42
B2G8PyE3c+vzY8ghCWWgtuBdCQQs5dWhA7uG/bHg2Ck3vGJGZbCdyqKFw2EwbL/K
nI+yfHUAtH9xSSpqXX6RCr4Cwr2gEh25bbuweoet3qwlke0llzt155W8CKrHd6KB
FdXgj5/vVLPSt66V36mctudWp0WbpT2A87oMivgmChthK0kNZ6cq4LN1znws2k2C
i9kaT946RRVt3GAZavKuUJgvK3ugu+wpYoMNcRr1t/uI7N98JRbto7lAvyw4mf11
r5JT5eVRPrQucNjs2cJsWNVe8BlhjUJVExsRc0YTWDPc8XmgP01C4mxH+fRSoZIa
ENKa6KiYh8oI/lQWS1SkjKFKWUr/nknv8wROokshjQ+93QGR5kGyv2HlhSHFUtko
pWJgEyRB9V+aAhsvAHMSGw11pMqUMoTJ/t460OSXQlMoQlGUQ/ihmJWxnZSMvb7t
K58Ysou9W2OqShOWnqUHKX+hDAujSbDlzhkSOa6XI5pri3UoKGDkyjUL41LA2QbP
o7RzQMX0kLal/fmGrxfCBQ2xVVuKtkDGI+BnmVEKLYHsSvSMx3daP+ci27ehAAo2
OaB7+p8xj/jgGh2L8EWMXl9R+UNCCSVTAiTfEZPDtcjJvYYrJpohiUOGN31cUzzo
hJyQaTW4fvCefS62LSIzVQyYyvNoUhSSgqXvHmZJhuqJv1e49MZR4YYnMRR+4FQ2
4w2aGH2jwjatTnex7Qy6om260O8Af0ainqA/nr2C3v7tSEAYO8R1XAskuKPuj4zy
8/cj+ZxygaZbLbTWZTRHtOlQWEyiEXWvD/VIDwTqaLPIq0TkXjWTQa1weSz8kVOb
dkdjzId6xeIW4yc49jJvAp3FuOXIlMctA8gsytrHO5wqOmjVYHyGGBaClpSYobyS
p3Ci7ayJZlkvLKVOSf+zEugRpZMzZKC6cPdU1m7QhJR5lYqr0eBwlCfHXrpNIlJY
YXT1ws8hciddMlxH1289xOW3so12UYbCZW6RYVhH6Jx+Ie17WmYzJ8+YDpin1Gmx
95mvfat91O+kapEhWajCkPEseX3HSMzLlFlFAGDVmzcPo/9PZjrV5ulOoyK3fxdH
H+9KIUQi5nIlzfglUY1uZpzAM8/DyiNBVVxKzPLOTeNmHbbY4mJ2oOc1QdQjuBTw
9Zd0yyjgAwjuElm7byNYSqtFk9A2Rf3If4fhcOvTPdae/2hVvBl2TUzSOZZLiQeQ
vfLfqbwDWFYiQqJzCYyn99WbsTL9tnBw9z8ZYgVS7/nJQr4gAkKlYoNAWiDtTEmb
dRjE2ivvr1Mc7IhlF7t+7klwcUMhRMc5YcfUfimUxIaosAfVeTcllV6CF5kKWfSG
qrt+zGuwu0PyGSWH0p1ZFmFycDmlSHV/tETg8NtGjbWl/g/XRx4tjxn2G0/K7ggP
/orXWw6bg0DN3ZX8/ONdYciA8OMbRpRpSgJRoPkn1LbmUsabk0z19Oq5ddTyUfbw
L+xastFStSPFmUIbnlM2cglP97BBfYjMsqkXv/Rnh3q4k2axrQ9hg8J83UKm8HgI
TInBLyZVriTZ6oSUO2i6/rMNl1WnMIQ49OjWqSVwh5A71tIspEK6FQxxqGu6VE1y
r33oHAM8OlpOpy7oYddnUf5hiYGkdhefiN42PuiakAJWYbrUhM6kgOWBZZn8uTyj
Ej6Ykx0wW9IIMapz4AcG7zLnjjWtHY85jF1AFJU1fa1JHqHFcI5qYu009veNj5tj
+zvIzLTFhrGVEj74DMcWSvpBK1pi1BDfAR01gGRzstlHewiZO/7vQY5Wa0RpZvF9
yN39m2qzd7yrbfQTweGy0/J1bSH0fqoyDSKcBKPOpUAiOSi5oafTxfOvCDS4d+tM
GYbR+TINl8Elc+KWmrhDmTq6qHX6XwLM3K1IGZ53yTAu7fCrc8Lw8wYUPDMKug3m
FtHm0WBJcZ+fc4MtBCqOCbH+ihQqE6+b5TJBGUSFCk6G37UPQwYA9FrbTnIF1qRd
x746mNoO8FMzb0RYz4ra2BMrJyiQgokUu0z4F6Y/KLAQRJgtw5y5g6cxz9z8tatR
/GIk5aKTUWBsNTT0mEVBb4SOL6QF1pj7zpbS5jWi8+elAb0EjLYV7jmxal9J4d8i
8qzaanFzKtDLI0RR37U5uP0So0qofkzzUm3EHGLrsBrlXzE8nCa618jyN98RbycH
qqtMJMz2tAI7QfIOqA03V86pH74+PlQ95eXsFescVU+kVrSV7yJYb0zWcTHmHc0m
jjIUuEYNPi0GjI6D7ZG1lrTsXkQiZwsyXFauaNhRuodwsRgJ0aJsQUetyx2mVH5k
1LQyD40rh5WdPUQgwiBUOHw0UZLbV5wfFP3lQCA0xrzmpfd7PfzTGH2SBcw9m0Zr
vPfhNC0NcViA2qcL1yweLhqnjzCwm1veZEu9X9byCvY=
`protect END_PROTECTED
