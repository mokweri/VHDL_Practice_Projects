`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7PoF8DoDHHPrcG0/jEKnle89mH7yCm2bMMrYGB/ZHD1zgyDy4UKL+8zYpohAfuj
cSv3E4EaJGlLnOW+Iz8PCSBBuhjh8dal+C8jKeEpyiR9ZeFzCKm0SyGfIu/VPf2V
XyACcpLweCF5MYNcbcYus/vf/b0rHHIWXB+Djx2NsGc/ZmkDAhpap3Hf9+yiarQX
CGuG7KUOmhf4NfnnIorVYscxS1cYReSA1RunPwZxKIRWMQF10hCo/VzeUDHaCBE1
cgRAeT75vdXX1fXy+b72FjwXCeM2btJGlVOrlvw4JWYjK0EZxxi6zATzRO7EHc8z
hXaF7o0ofomdI8ZZH5Zkn6cJkzmsneHHi1wjIY7lUoIiLsdX+FOIKWExM6PXpxcF
NLGw50GjlERezICUybRNLhpxenFG73CDWTCrCPmNQ9MwcoBsmoWYp673/NYouaPv
btL904OZSJItO03KuqEFyTHnr0aABEsEI7lcuYs2AbY8Q1SZ2r8h48+F/vTbl1I7
BYM5uB1ir7tEPwKMl64cx/7zadEEGxO0P8m8/WRLUiE2a5BLq027J15uBEnGnK9D
dkL2Vtc9yaWoBpF8Ipf7vdnveeeewGBvFG/cLWQc0fqm05XpPWCMGFesp7rykc4l
shGHMcEhcxNY+wHS9iDMcA/iOpfdbSwMZfvacQXcqgA7yLLhnQd7H5+AdFZqjjNP
pMVySo2e6+SrK6wVFd1AB5aJRjxb38Rw1/C2q5YDOFudaKyykacVQNwgCAP9ZndJ
OwrpgKKKS4fds79mhJFXiSXhoQ4jHyeMU3tdHHmvAJFWh6yVT5XRqxKNnuaywCGs
3pT6ydNdY4rfnnRowmRacbBXwxXwO9gkYvu3QqZzui0l4ZR3QKjM9qDs+VKRHdR+
El4QdccPjx6W3CfpNcdfn2JGaOrQqzC6iPKZtYqwgHj5y3TEyf98aX43oIwlwY8P
w+axm0+GlZfxFdtAIFXI2KHw+9o69L8fnmR8Cv2qZURlj+zbm9vNLeK6JrnqGJw5
Z+p1iYwHs4DPhNhR+4PZ4/+RclVx2FKbiYQPofhroAg6NSh4QkcbMaSS07h0xR/2
CniIO/6FXoczoGl4e+7ykU74DQ/4tlcsFY42jAsaBIp7RNgBvPQ5lyKtus0Ma9ek
ECpPHa5UozDRETrIWDZgGli9Xy2DVR5VLencW06IG0YEsA6y1wyZxujiES/wAruw
IZ1JNWff5ddki8pdv6xCB2DrgwV6pHM9EtjM49fMAOeyMHon3z7bE6BK1p7Wv8db
zqaAsNL0loa1KSi09n7BmqD+pbtD+9tMwHuYel6DeEPbxFtbjQ1HSY8/Li+HtvAW
Z2ps3ky6Bv43D/yN07g+wWzGZDxRaWdgeWAJUJ9a9s4ukAA5Nu5fU+bSP1fm9FDJ
/yQbRMnPifW7vwvt9+8qBBA+yeUfLSNGljhmrwouIqCXw8Ihp45bKkA+suc5Xmy7
IcBmDUdy2g0fs2cLFH7j6GwqwILTOURWjlV6EVTeCzIDlPm1dDiRz6qiwXM0NJYz
3bHexg5/cgJcxycRK9HokdLAxdFgY3CKr3SlR6ppu4qNIMWzVeCpNf7oYIfRfx0T
UE1c2H0WRvvRFj7S7lvuTDq59+qgpQizRXwzFgidOknpyz3UJch7b59jHOfXdrcA
XhSzGpUg3uOdJc5b8ifqJ3k8ITS8fQx5kNAhRQw+28sPrAibN+0ghH7utk7ZHp44
X9i238LWk+T38j8JgcdRMTfB1t08s5KDuRbAPpnrT4Que36vc1xCuNJNIsxhQyI7
QiyTTosiy7z6J2ud3DIeIL8CP3vXcDKZlrrklQEGAKu56Ij9uEOncrhvUwl4ETLE
T4AQniMuD7HYWDWfhqU3sFz01CGYNcOSSeMpA4RPJ1fVjNY4/xssgWNk0xnMFMcH
8bGBoF7oM/IfPlEtqEhzwQdzXJ6YJ5fzeJNIqRxJFJLpDT3igZ81Jh4TwdJA9EHZ
ks0+GGx9hu2YNjb8jYIwghVkOBxqMXccc7DjzRz9v34y0zRMOEeVa6FtzdUEPgVO
S11k41xro94ACCS4by9//im1UNQQjxg+Dx/JyR3fOrQVMQmRhlX0Gp0KCc+aUWos
OsSFtyHGU/p9ExiMu5yYsIfsAaApEhFdQcPlWXLCUNHdFauwqlTvn1VtNQl+gatn
r2n96mVZEbhtl2c7/3fqwvQga++dJBwFUSKrXEePuFBZx9/LifEbKRn2xJPQ97NO
grA598/Hp4x4oTOMZ3+TBqmfvMfkGj77x8ep1Nlz9RnJX3KF8mTLDZy8VWxX69Or
q92FyDbjRs3MLrIfCNC152+4nLOAtGtzNbpvrlv4m01Uir64fCFiu3tFJZw0llHx
WYRwnTYbERxIZhfBbDnZTEQKPVpUFpHPyXkQBkaJ5E2vmNu+DKRelFADG5Z0uL9G
0ZIl3dQyziQaZcsySelXCdmwZmOPaHbGLuQte/RNXa0CG0+inVDeVh+XlkN0B0hd
iz+raKq45TCWIaIbBKtuyHvX5zprm1RFumMrAb/3CAgcrF5dbyBrAyGLWICXeVsu
33WQ6+3XHljuk/mxUAfmDCrsNthiXIohkMJd4uz+WYGb3L28cYqIN0XIjU2WaZtj
fcKvjHtmxRBN8rcxTR0VoGbvmJcXTR2CxPx6h2pF4N7MiS9/p6YoFSmMcNbU7O6z
Vrwl1iJzYhk/6jdmNEFogBrfuvztWMh4dZe6hNFhgT7Qy3vTuYv73hGlAiMuZjtC
XcTKVxhwl6FG//caKnCieKXRbC4hgJ76/+Zgx4lEOM/v1k2XIoMfCTcxvzUqjV8u
xks3GOLGK9OB9a+9j0ARRzUbSfONZ/9ijeXfnwb84k4N71Y/dp5nZ2KP8fjEZlmQ
jw2Vv9fi9540d3AZQ1UT19r8CJ204JSDQegaNVzrh8szXVRGOiAPwNaDrYRUa+F8
tv5iSGx58yjtIhOZQFEglWpgQpwRiE3EQojrHyPQg5RcV2kFa14AVWvFvMfYoOld
pOz6pTvNYWc2tJVxu+O0SCxtmDt/iEwFaS+AUC4AC9Ae+xNx6hLruQ6nYRxFf/hT
cNJboIoKyFi+NOwPTlAhvlHPFFSuo7R6QigBSmD2nVRRJUudzBYQG+84dTQ87rAS
ElmFO+UX8Pqwqoyl6W2YCnvcPEYogIKW/VoXLJ+MGNr0x3WJ6+8ioCQq0SpaZ5Q7
CJ3bOggvgTvBOGWPr+jCZz0unnuFO27Tj5+nn+8yluRWEHBVTBeMUBGMzHTLVb3K
cQl1Uxxr02JzdSp1iFYnOfd3NKoGtV9wbWceibOhpbpDb9g+4vXk2Nh8nugXvl60
GJP/KJW1dCra2c0fW/Id0RDY4tAigoL8r+qkEBGd1WfdMceo22qMbqEFBzGijxWd
K0xTfHm+g6cSyhySqiAp7eYvl7yx3IouPT6vq4L/RJCueD8gz8FplF0gyRXsbqW5
7wEuIgecCbmyZk2fz9hW9OXRz6Xg3ySNht5EaTNp054v7GYBMXXzfQ1uPq3jrEMd
vKch2BOka/nQyiW6233L8KsDbb3DhjcSvcq4In1Iby0flAY5VgWX6H13kDqSOiwp
tf12ikeJKIRK2IjCl8MzgPuCNFeHPp260pF/vYqvwC3HQTRawARr6Eo23oo/6Boc
DoWAWAlDA8VYGwV7Ho74v4Qj4kW24Z4t1Fhcdzz0VEJupl+H3RzbGyAagjz9kMyH
4ZW4578pUE6PmvT93b5OxXregWcEvrv1iVEouNTpoqUAIODand2OkNjiC9CCOTgc
63H8IeJZqCAWjUPPccHv23xjM2E3F2Xvp2bftqEQWKS0pP6/tZhOnheYawtby+Pn
rCsY8cFtk+miQTLuvCbl5IIc8J71zlF/9ET62XRGYnzP+VZZWS3Zdbbiv0+UeJd6
Gm0/7pPFT8uO/CtWBH0Y8UMWX3tVes3zmHDg0PC15YabZrDiAx6kSo8ji3EgFI4M
v8AJ6Al1sJ4JYyN2JJBPNkEXGYNaf7Za8TC2wzc4ZYIimKoy5wjy5kjhRTUGnRJc
lABsQOOMRqa+YD1X+bPGofjr0JxWue5lm6CkwAKVefp5vsMIz5YerIgLytZzyyQo
enPZu7q5Ldi8mnBHhyKtA8cNasIuRA8XeusstdFF+mmC5Ah2wnh+ftAiHHue4HZ0
2nU7DLAkfqPTUqmsHGaol9o949RzpE3NujwHfc2ZufQM2Vf2dQRiM2TPR/JEn/by
7NEzxS9+2vw9egF3FYTKmmyQ6ttnBR7snw3ncl4Qk5sY1flm2Q7aEbuEgnIDtBvB
AVRMK9dpnA85Myh+ifm2YaAlOpLy5qS6sVHmKQbAaz06QUp/fg9DwMnZgrQkDCJa
xf1F9zdCgYZdohCDz5xYv7C4nsHOgNT7DcHx9sMw4QZp3IIiWtuLud5Ez6gSKRM4
Ixve5/MNAj9CtTqXCuDMY+UIRduIaR42qbayHUNIfeb+G2TMm8MMnZBcQKoKi24m
R7cCNmB3qLjhMRupD/BvmjBPR+y43vsBHGwHp+IblPJe0V57pqTmKNzwgEgOqLvY
sryWqNUkJ0jGcCrupWvpoOA0iB6b3hV7smW5w04+/BRxLe8qYC3ySt+igRoBsN6j
+oBLbDi5UT0bsTuSOK2HvTcDZjIspr/Oj88FFo3AzL0OV8kMi1ar1CZ72eQUJC8W
t/xJF3JAukQR73PlGqpIh88GUDj/HJV/HsQOsvA+ovlfik20ylaBQQ+6SLCOagQm
nApQKuMsnmepL8VsQF1xKHLvLw6nXHhEClmaSQWCenEoE22K6iPkQeS6CpReMnlE
t+R+xg1rPjIgBvGq4p+VpbfFqOfCDZr7/q0s9kcuyJ5GGudee7Xsquy1jf7d7g6G
c9qIYZWMzM8w82/50PKnJ2SiWmH3rBde2bUJ/EziQZjQtQyqHzVzq0f7u3AGIm5p
Sd1ksZmWkc8nmgMSUwa3KQpH1Hjm+zOwbbB8HeOB0HkL8w/dFDBFSLSS89tYlOy9
7BXWON/bAlXLDTpaK8cvd0nszAFe3xB2/v6T2OROL0flftwOGpvr3UPG3CshdzB/
ga90vddkzqJG9wNhrR9zXfkGZlvfxU5FThJD+YK3raVty2BBNbRvB3suUN/uYc37
LqBJwKpv6IeXcJUlOVkEmtN+u8Amg//zS4O4FtO6kgjELxNaOl4eGa0WYtL8ni2Q
+sevPC9ovqVIBeyymJK2k6xmPfskKWAh1bQITq/lDVIsdcvDgHpZWveNC4yCbIfh
oYL3/iE+3ivjqXJQFNq/VLTgyhLCI09YPyNsYeka9s/8/qKW1itQXdzch8/rG61v
YMcVmNk7pVGOPEadMi77SvipY5rAYlnnjcBTpsHL/rMSB51IbFDDqeUOSmdp1O3n
uvUOLoITeuQRvlv2hVTTfYC4aczQwQPZV5s21gsowLVUeENaeGaASCr3dvgioPhT
iwnfsos1xXqoFKtkzKX50i2wdvse7w8LuKmH/+KQH/tjFFGB82ejEx6YmHka6AyL
9wlpKhlo2zl/p8+anHAtsdApPmxMIz2Q6Twm8qGJan6WhVv0jL/NvcKRxi0zWS+p
9uxbUwr4e/tGnah1PayweVkiaw3NaxtpoXp6yqh+OytLT32scq89WkI6pDhE5Sta
nkDi4+A2HxtW1clMlzJRJTYTh3r5to2hPTmnOygJeAhKXIsdjVkkCJNmJgVPdAxn
rMEEK9L5Mh7uJhTrC7s1doZo3JMFt3z882eaoBYw2UoVt9VsyGDTX4TgUAtlMcvE
CVsppvGHHn7DEXe1m7/uJWI9zskIjNYK3ZkmQa+CRyDC8HYTEeU5Ya+Z/CiD0UmR
0ly1gvRGW88sOq/N8c9Coo6Jm8XLNhtdgE8pKOxtTxwFOsC4JCcYi5Yc0gKn5wpG
D47ay2/AGHfaSM8EoF2bk0CxivFZ821BopzB1ulJGzd7Zmzatzt2hnLz78R6YNMp
qn2xfmXPzZYC53MkVMAdxGQNtCWFTN5oIPIhln23E7Ufc6kLKoabQdw2GNW0yzwQ
EmuTwdhhafalkDfSsN+o8Oe7h6DOhOmFgBxxeaydTLH4SMsPNz1UskDyXKKbGwZ6
TtOPs4wqxEZMbIeLkcTkHxOUdE5g46GIhCO21pz8tmaloLLdkqQ/aXJXUl1s0g6n
151ychGSkhwhE5M4C9OnGzFuaUqSjDKeExVJecYT7xtmEfUt+geZEz8bMDktIar1
GD3Kb2HdWYrbWWnsaVLrq37q2QxJudjOvZ70yscZ80IAI2QxByjiLcW71mBKF6k7
UCc9UsaEIPmFNtxmPwKVTq9mvKyUgisGxocmxw9ZWB6cmCUt2H0TsuHxuHwILsmg
UtxfbevXR/N01AQGjw4XftP+KWM3oqYue8rb97upcZxdY+vrIkfGBdiB4Ry/PRep
K6Hm0MNwcw9i++/XD8ESewu+O5MMuJkRx7hAvnxLrT4xM6pEzTdD+uxvEs1suJ9F
H08zSJRSAETK242khxlkzjVYAWrJ61BL6R9Noo5xwzEySpHiJap+cb68HizFYDkY
Ry6qEifnIUBrDQQlDvepiEYHbWo6LmAGwMkSWHc496fjsa/VriVscKAklWwi/kM7
TBHlODKGPj1+fsVdjRqWlYu8HAOVjGmqroNEKlSUNzyYE1Ll25YkWQ5uwkr6lbRF
0w14eigqjOMF+4yBoV6/nJx+XWgwDaedmyKrA9o1lygAsRSch3fKj1TzNnq8gHlT
hxFtfZlgDygktQtCOK/SzF78RwT/dPJtEfIl9h5+sQCyMTGr1eOOCyrYMCRFZZDU
n6r+b8R0f2J7rOjm4yo3vB+e4qHuMhR5OErhTwIXG5UPRXQq85KbAdNYMlv+6vpX
LDU57XXRistSY0jIIBVKFyuy3OqgE/ekJTOa4UGX+9ZFE9BUJjc/XTVRnLPpvTbH
8E9/DhUJZCZDhyP+9ghjJkUGgWE1BYisEcHyeVmV/IBXIiGhLav4OwAq2dYcPmKs
sQchA3McUBMOsObhy5jUTOXjYqSErzSk4To2JOHYe1UanQaTjmBm32vBizA4fP4X
TN9UGmF/vAqRXuvH0f5/JC4miNbToeuBWd8e78wJFj7p1XmndJaTW01all7Y4MzK
E4c6jnSfYx3qDnC3/eNiSAdY1jVuDSSjV8l4B3pPHPLZjU98uBqIdYT13tJKn4qt
gz77PQXbPZIq6wlHrKGVVGPEgPNPnsMJd+VsgsTwPwi3OH/rkgWlSrH0vGdVG3gy
TM1PggLeezCODVo0l7IGRbz/dh2dxE+7RpGEzlv9sTk=
`protect END_PROTECTED
