`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GP9G+X9WJlEtMq6clutODoeyW/kqgNxnEEH0QSNr/MtaGVomERVMARqwXE5KDSi/
bCO2iUlp5mK2xTtxTiW5RNjNyRbLBhcDb7tPbblATfJkr3O1fbbEn+I750yBPK2V
rEJfP5RfBIIbHA6fTULDPyLn/Ou1pdxgzxO5XAyHQ+M8b5nqaMEIghYLhaFGd383
Bxy+y21Ehvne7ZGaNqzWzSBavmx1f8ghJ4xetC3N9wuqUbx0RGFnGJzDeE+LJwcq
j2jkiukxgk75dQvAPIKFcqfbkG0bZ9p165knF/HC/Ptm82gSZ6NYKwhZtR06DBaY
gnWjfd5AS8Cl44HrM+ptCwTENyRyzqNTbsaoIitZAW842tYj7Gd02geAuL80Wnda
hiyHPX/Pe6VI9jT0I6f888tj4V1AIAxMLavRs6XDm64UKm/1novm1dFhrptuRtWT
qm98g/HvQWia86GTfxeE110iy7bEp39z1QvrsdBmoFN3iqAl3d2dd8pA6aWAtPnT
vC01slUL4OrwhXYShX0NmjHxLeHDTPlHcUsh9qvppIWYnDhEvMb8BlIxn7C13/T8
dBa+rr/RJbXnaCvO+7viKsg1l9OevTUOlFg4ceerSpUA707TNFE3IO8h1M20vy8Q
rXJLDXh1TbclRMIUN06XVSSToJSI7zc0vxXxp+JGHPri+RhBg9RsSGmrkk23PZVH
h4HoEC4Whs18w6Jz3xTZM71PN8gwUc69xAEa0VQJpQ9NLmA+vh138vksxeaDpaAb
rpEcdWe4fdxSyVIBFw7E/oWEzdohqJmIcepi+5sJrik9ua0m453Zfls0r977CoXj
X91mbofTpnJ0yIUZdFFoFD2lazfo2fuUljRtv0VwaseZsqIWh3WR2qUbJR4Rl79r
blSvu/+1wUX62EiwP0vdjtsFrBP333j7CpY7/ikB/6+nLceofkxoeTA7BeDuWLf+
bzJN/A5T5VOOUMWBBIbBbZCZaOPrkp7yFvdjMyXeZ+Qz/uX0FqsxLAe6Zrrr8XLd
BmQNspj8HZZP2LeuNmahc79E0QiNW8d6ky5UXCahNFamIJbsP/l7avR3q+hmLthj
uP+hcmX+Ew/OmxLs+6Q6sP9YNi/QvR+k68re0hhTd6uECt851jfvB14X3jiCeMNE
dGe1crZXONcwNkOjbYrOZleSpThuq751UXt0KQcCJRhHqH9dkWGsYHwPuiNVwa6B
PB5aji3yug9+5Q3/TvVzDmmSeHWzcttAP3m4BWMF0vehnD5LqV0BecyonBgU2BgA
m0M8f2eAfgVAD44usEEJ9Y+LjFt43WgIpsFql9lKPIvGGvg4on28M7RGk5e7OHqA
h5JTUekXKo5wwN63a37R/RovotAb5BTxAthkfL8Nnxk/ZqIx1QryxkPtCIe8QQsf
MbGirfeW/qunLnwrMzUfOtUv8lLZCj3uYcThI8940vQxzSLaXyK8tv0BXsPlokj9
bseliMCSmfzO7MglDdv0f84Hv/v3POr4oYG5Sc7nbhfgkl684Nyxexc8FqbgtYtf
xuSeZfGc47oz2cz+iHcM/KHMgrYoUTcVDF/GUDCw42nRIXliPo2INbBgzsMAyvI4
Y1kQK2+ipimjmKnjH0qdQYhL0DPKbh/hwoKPrCkMS07zoTUHKoOb/yfBRRUM3Fng
j28lwfwYyhx31t8i1wb0iASuy1y8F8XUtber7CinhzBggK0GNFRuwUMPOqC10srn
MkM8zbhttZjmgJ5DdAJLym4BmydLXHxQV1ibIVXQJIQUEydd//HfN9NakRDuMUR+
nby7R9qh948lbahwTj8WgmArUdp5dzU4W3tDB0czAVM4txMDNDKsU8gaXHaXfwBK
YVVY0xYUBbGBrBGu0uAOYlY+ou4sBY5jvbhxs6agzyZRMNHNzcEq8MmqNOYE2BM1
mqZx1IVsuOjKxog3yFtxhRx5U6NJW9Pmbjpur1/S6PgUZ040FeWYZiBzolTFC7Sd
tlfM+0wtQRZ4nm0RN+MGwkTc15wXPxJx+9m46RwAYdegw5CFuJa9ci6ZqkdCpCEQ
EpuBvv67ruZGEPlUdw6s5J3VHYfOW3a0X6asIHtuJjbZU5qd3mtirBp/Xd2aC0+j
2wcpa/1PsxZflpmWsxgqG3e1fD6X7NtC4zLjgnw2Md5K2OzKcYLy58rAkvyiuo7M
fKD1amtHLNAE7KNkglniAB9EPqzyGMTrc8jtEwa05l8oJI/tEKYy4HFYTltktExj
rDpGVVxtOz7LC+E+o8t/xssWpN6H8e88qWLWVvT5cdZwJjhsu+Svm/a/yr+V1KaR
3zM29IAtgI82DDhVxHr726TOrKxYDcCSf4IwepWksXh/gPGhIVkvB49ydF1WYQc9
QZf4CHCHU1+xe41d/o1UIgKSVQumu/d/tCdFfc5vgs1+aspI6VCBQLQmcQ39tB6O
QLyp1Rz2iyY7tWEwccSouYRbl/ba1VHF2EOSxAkrHCDywofuhVd6DmYxjsTzEZKY
SaXJErwA7khs02O7IxE9cNsAypofp7eYbfrW0DMC7BbEo8C/jre7Hb04BnBrHiKJ
rwPDQahEfz2PEHCW2oZZzxJ7uQI5FnvDucddR1tkAoCP4Q5L4gFIaoh2JgwXjRAb
247shA9LIu0kt7R0Xz5Cl3xBxM5wHaRyNLnZm8vll/DLw0A//iRUrRPPvXX8NGyr
TH9/bU68crwHfdnKzW25S82hJmH8g+Dv7JieKeZ6puKSwsixh1add12CkWLd78ZA
GNJAzOzdyk5tnz0X+jfBM+tEXJ/KhE+vnfr5DhxVam/o01md6DPiLjbt1YDhMojG
wl2qKvUggMCtxIA10GBh8HLBa2dVoH/sw5aFoxwRxntVcf0QWz4l8e6jz1k9A5lC
Q0EHBGJ0qDCdlx6TQIS5QlBeDIckmsYvfPRUBaROP3V1BEF6BZX3/aUN9FskTHIW
V4jJkQ8zmST/ILLbLup7RQPf/5/JbBgiMa9l3c1Mset8ysEa0EVxAa74rynlXksX
vuLJq/iDHD/MPY3APU+6MAM4cOL2f91JArGEoRLTrBACxyh24iwH454bkSmLf9us
P5sS96QQcU/SvQQgfeGVZYNbtHkM4wYLdt+qSBYchMdlUeqLtwUj2AYYh72ERz57
Z1B7XTYo3otQ3pVNn0WAaj4pVH3srfragFg7iDgXY0ZXgB6DlkjYs+xSGW6lVWPG
xkMlXx8LZ2PD3T++ipcMXyNSKPX/9h65YKq8P1leknqjXlmK9nswP+mp96hTTGBh
i7ivYuBqzOFyK5eNx2XNYSvz16qfDVh9BCuIyfHZgGyYIkLKhtDZwVtjMMwkZm5v
Re2tL6KQeFZfxa6OUFJn8eQdMz8dFMkn4hb2Gb99k/YGN/xqKLgCNJRZBpe0SqC6
EErS0XQQWb0zJHuqUeopmSCrvepPY+unvymerB4LVrHpLcLSw4XRcvpevL0LP/Rk
baTiEiukqzyEKn7YWrsQ03kAG2MeMAVLD7XHYqWFstVaM3ZnAoMh94v5whFqH502
JTXQC+QniWar+tmFnzh6BayMWeGAp8gbJby5GALhSSBBjK3CYAt2651JJ23byznJ
oLjKsRL2RjySlZuJRiwqZOiULgk/enF2pt7PI2mhTYcEHMB/kRP/bB+61D1EJVDC
OmshZGcO7j16kwgW9NYwprxWd2Sv1/iLoHzD7pJ4XU/bbiBiSN16vJjgsGOPKUx5
fq2ZwM3rMUFKzYNU4v3Tt+qrOHPjEnal4zAFULokiCmXemZij46R88jYKlH5NG6W
ZmzRM/b8vzsLLu0EvM1RllqEOdJTcQwAooBFQ/uAVpPqGN34HeCvAyesNHbI/IMx
4vKI6Ntb1qFuNc7i3OgsDWPBiABL3DrpCmVp9u5veR5Yjuoto/RFnTqZVoc3M2Kx
jR3jLwy4/bKz5Zg+eC22OBqBb8KwUFRaHDmTNKkm7PosPqb4CEd/yMKmYo4z30J5
u4uqmmPC+4ihXW34M0nENiz/18ts4t9iEPWJYJWrzbqw6+cIcrQv2vrAOgJuZK9M
zsXP2KTGxKzrGXs1ZO/gn3GRrzQ24cEAerIag8Ei1woluYb+ULqwyAw4mywgREMw
9VH8/P/hhhC6wLZh5oBdMfzKwdWpL/j1O6sHdU8twuzHq4zbIxiydmbnmVEQvxT4
7rzlx1e4viQLQhU4yhqwlQCLjY1xKRhhbAQWaoLHMo4YX8zIdaR5IPqIYaXShyE6
Qtc9RF1zT4Mn1e1de0NA/BD4ZOatbR9BjuYjXSSTjmNLL+rCJIKtHT6ePAdx7Gku
o/68eNZoymhokutMdBAz7XMlXuxazmZftwDNejnBQhgnsCgSl1zEKblAXgx7uYbt
S4tCi8fY6NvZYU3NLNrgHi6nMDAEpfQa6hLsNwpAQeUK/BInxscXjrL4CFKABqRW
XTXI/z5maPW+qfcR3AtmF9FCjWWe+c4N7fCQZScqPRU5j/yBuERyDSmqWwSuH6Vw
NKHvN9Vn2ldwjpW2gFDVRG8SKimprkAPmczsYonObKcU9Mt7n4IZa3jDtaSnoirL
+olMt7ahFNyt0XR8Puwa/wBj56XD7Ojv+yI2Eo+pAxgx3WoR+Uw/DBFV4zjdBQj+
Y7NJIdiCIApzmUZemgQlFuEjb3mOSAuNO6TgT0H6tD0+KHZtHm/ypyt6nMOfcft8
ZInX37Db61ODuqk+3jvbrxl4aMZ7T5alOAD1JgKIYFMOPSZdlIHEo/N+HHPe+nTM
4dcHJykm3vjTOjgWEhD2fXEbxRPQejH/E/1WnMJzVujEDyGGXeU1D7dPRC9VpZMY
ImMZYZdmjZZHAZDOLe0cF30c/3DInTVtZoWms5BnMXAxlDg4lI2pl8yOSfLMNWoI
/aEV/GWN64MSY8TGmYm8WPvBSqsF1smQKnnWSAw5l0qEx/k9liZBOAD5dZLGhndd
BtxJWtbDXWH+qDYDbzIXpPsylPgyUxdGMgIpev1Q1DI3x+1J2FKNir8qoPyPwAb3
+RP+QNBDLeWo+hArGPOZQJyDNE7Kue8kur5iPxTeaXwKLciWQJHGK5nDgH6uX+6+
DCgHDwwXUxTqQnZ+rrGvWg==
`protect END_PROTECTED
