`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8Qlw9PEBlYCdYgcqgGGuk7ut2QGZ8VDUTi++NN9cW2IxkuKoaiIB1/2hIMG1g2k
ULtBUhvuI7G2tdIiUKm/lDLzI/P2/BSpMIpEQMphvXwTwtoulmUqfYluTcWTtdVb
TVN09iaMmpjwYnCwDjkRfw6A+lb7WHJ7k1Gi+1/m3QLB2YX5nAKRiU3QxteUuKIP
5Bgc0LjP4pgi9RdTQg2FLwJGgMpAgyfjilmCvftIF1qw/hEQi5G67rR6coBn7QM0
bl+VuvR8c8LEuE2+qqe7ks5wrEhCQGyS3Ibk5jmmVAUNqUC8iHsLsEAAsvg4E1HG
H/UtedoFmqHiwEu0wqV7TrHzO4uGs6k2bEHBMOJhLda916Ca8nrZp4t0rtxkYILc
/vjBJex+8rGy3YWcVDOJgX3RAb3pV5YHfuqEb62gBny6nw04l5Ttjp0QM7JtkVkU
6gCYRkoUJCD5BTqJUeyvmXgmLlxqgLOjacPgoH+oNzJKOyV//gtntC1wOrw5WPSG
f6urOzps+C3bBiM7nysPfUM+BTtDFTtGzHQdJq8i+6UF9rVcXXEbDItE8htmYT2R
V6NPgIhARWnUy7Mwq7KDzdiNQSCWjXIGKHeURpTB86P1fxYb0fiitAkGmyixHESv
LvmYrzDz+XmWM/qKflGFh5eCE0D9fVyC/6g8K6kgdQwaBKAsFd3984ukjiNhPuEV
B8b75xA/zfSfNB+PUjMS6ukKlY/vcd4OfTj44tq5EkwWh/879lQpG6pEVoOkldNm
MrZJzJo7b73CSKeSnbj6XmaYrBtVF57ucm7PJMIgOV1SJpSTOlFvx22421gjnQYq
WPeTVth4TLdtCVgzeIVugabiz4GSjiNkK40NCZYXWPoSupmioV70jwhrIRt26dtk
ix9B8nR5yE3wQtDjiPReVNCrKEXkLHhXLARGzMb4VcEV8qAKOiZKLqY7u+UxuDJD
hEs5khaXUwSRqOKoMAwKV8cx2FKn0OMGnxa9PH8MrYJCn5AIW/nerK367mxvOgel
yE/jcpVAc30gwNxbaj4WFlpKpXLGVopC4Vvv56kTlErEXk8iKu94nhraaRPlR/9U
lk3GI0Vq8Hr9DkDPkeHL8Wq1YNuR8pI1HfuU2nbSXrpQnmFlRuOZo0/Kn7B1hxag
p7ib1764ux3Iw3iZuJA+ulYT5qySp4dmtOs/iMsLBsIF1w5gpAXfVj3GY65nYBCg
69IcKfPdZaD4BUXftRFXLgrz9MO1oaokYH8CuS/ebbDP7jpXdyTHugHEweJzcySt
MnwyzHjTdvJkhGUYt/S+gQ==
`protect END_PROTECTED
