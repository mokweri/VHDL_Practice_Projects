`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OafUjGbY8r3StHgdSXzXmDIRURzTDh7iJAqpolbude1aYZO7aZmXCqN03bdrvrIl
qvw1xxMohB1jueRq0y2jQBcH5fTuXMhyI/qYGCyM0YxwXMR+uN4gsx5fRPqX/Nv+
rMTkifl67V6w9JsPcV7vCw/kJQi1DOjkq8wLj7nknQ95jJELi1UlfzCHJYeuXNEe
ykvSxRDmeRhbZ/WOxh/AgP/ac4GDWiUuvVUAH9bEp1NI5Y9R2vjK3qS79R84NnQu
lA1UJNS6vGOSXcE+xlZkCslxCX4ZdssLuvY12fVFRjaQrUK7MLldw7stFVtPGBKz
UHLz72sn9wszl0m9nOYZ7bW2lClkhu1cqfbo4+TSsy64vXJPP7epa6ejpo/jf3bZ
oln0AWkdWJLs6JHBSLlT6P03Ie/3vRamtm9zhabD5tXH/BvsCtaKDi8Qt6XPjD5I
qdZ8jpyGAr4wl+78UPicg0M/etZfLFXlr0G0PB2qGt3P3Tk+DAsqdU+a9shaS4La
EO4QzZJATGTElZpmteRGlPQZrGu59+T7K6Y2cjbuwCUrC3mKey3VJXzKs7a5+qzo
Si39lmGeWwaTSte+pNqMhJVYKgBWsaVvL7D97WhlGQb++kNROnej/hzss7sYPT8d
Lgko0oI03982NhM328JyrkMaLFoRz396SlOld3e5sHim5QVr+dh0GBK3vbvoNt3T
+wKoCwAVFJqUvL+3MEIa09lI7/j0iMjkPmUc28boIB8MOeQ6tjQMcKJinMwh1Pz3
s40Vh4H/GA5gsNr9cyONOzJHj0i6vlJD7SecXqEu2su6RIGq9XP23MxKCHYULT4J
JNQuVHWbPMdnJOuyGWAqoX1kIeisQgwwy7v+bqkT8xGZFTWEM+LwkIztVlWhB0vS
tVLh7u0oFq5ulzMWUFGPH6A6sk79C3+/1z3OTDsIIJ8SZvfP481W2y1G8RNPMEd7
mEBd/AfgkXHJlSm6Jt6maERWbMbLJHwP9LyrLQqYsD0wZr0FG0nNegBA1flDExqp
2Wu3gY8dq/ub9yXzj71uaAc5kydKw25ENryTs7mB7MG/u5ZgEiEAikoxXQNqRXee
nx2EITRV1Vl0cK4vZaUoMxejVByPnrDI/VSyLAdYugsPzeCZjDWE6iFQERtt78yi
jGGFj4k9NAvmYOHeF3n1pmvVoeiWyWrAJzetZOTThaVHAv7t6kFQCXtC9d6aL8S7
ZZh5rYxtEid3uAWNaPuzr3b5UX5CusxW101QcHIKVPoZDrbphX6h7ocbjbyKDHTw
ECuHzyNXTeXVsDowDXPXAiuUcrxi5uy8W6IhHrxn/uRm0d9IkCnJnRQt8bZYT/3z
/umQl1L2Msynzhp+s98SbLBFJTt9WJOzITIV+khX5daSZLlk2SpN6aFIUHgxsx6k
t/3Kyo/UJRDrCHn271TijtkpowaRJ27VqXXeHmlA4qTBCBB5pGXwnmrzzlw4IBU5
RWcDw/Bd02yqSt2J9mm2oshdo+r5VFsGdzTKWr327cmNZOyKsZWEYeZaxgpvJ0nS
fEXfypdEvOVQ6jxHs1ilRrAMTwljtIeQJt/vaxFxKKX4wa5miQmSQDHK3NvoiZNy
`protect END_PROTECTED
