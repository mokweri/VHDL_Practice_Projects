`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XoSoshLnTxFqqwnv/4+PTQMxZz1oCydecjHW0yACCVK3MbpsIHY46Vh86ze1d312
o2LByyFO/w2vV0EXJCvgaSDIQ+VuTN2MwyOfef4kBV7qmNasC1gbGIHSBckP+40u
qDJh/GV/tSAJFOk6LXA9EPiYcNr0qGHe2BpSfLiC0ylivmX0sx2EKeJVkxyBfiJf
9yoDuAk6BOIJ8uQl08rG4csm2zTpgQHT7n3qCwGGy8VSOkxfbZH8m3BNBuOFXAE7
0K0ETIiiaT87Isavmb/RE3o6bHHl3fXqsolmsI26Q6D6kdjHNtS/lpUX91KaACu6
feyhXOYempjv2h3yiAncceVbmGiNb4ZsOwkHrlo0Li2S5qka1gwJgAJXNEh53ji+
QjqNvZMNBYV+syPm/6mM0ErbYlrF+5l6dWr+JOwNzDZ/ZRFNaujagNvVNJzrzCSa
Sf0CxhSVcHuLjubSgrebeQdmrJiOjPIr8iOlNMiSd4mMZzU/5saofdlEEAjNrTAF
wk9WHkPlznXmKwTwf2m3qRrwMSUg3mmBbY9Zoq1p3oyn1rhTgDaszXT0xZ6LjCDF
3e1eYKeY8nMiRZZivqx+xdZxmUM2fcWkOfflsHY9bb9m42RklLhRft8RHLy+ixbC
TQtNi3may7FxTuanctDaCuHbo9Ww9804GT4u+zikAbjlN9/6J/j7Wsx+y7kbt3kn
aasPZKXBhBcbaJvhFM+maNvaz6n4JoiBssBXfTRLJqn1MKgRY4O5ldlrCpUNkpUu
O/hMquCSI9hxrk7Pbd8Z9DsNx6RFWbr68uDg2bfBy9ENLTeJ/Tds+ANbvW7gObGl
4JdewNINxT+u1Mzt23zFaLdVdMsJIaAJQgC9S7hpQIXN9j0icrJWcjrPL7szZCJp
VypDYZlNqIWwHTTobtG7TZMJbSTfsNjdKqoWSTQGMzc1hg1F6aU/oe+YcCT4JkH4
PIbLIAP5+wLPxHzkWKDCrt3qtCnFi0qeJ6Fz6bEzU5Gi9kUjg0Mu+dnK/4pRDnrl
W4F/HumRIlxzup+zoyQptEnnCCl601L1lg/cZcBkyD2uE10UAWTrP+Vxsam50nrg
AuSiCaLHKK3DLe+mVffXD/y2/kliWV7G/tSPEMmK3LQ5z2NAK1clbdIZHQbwAYUr
+3/JZaHxPB1c9r8+qePddXW3IJIJyToQlwlVc0/4Ja+CtA7CsOFtFLuybwFMzXSp
7bzHDRzs5SQiL4NGQWaMPqvmx/MLBUfxVmlAUqjR4FG2h9ZSHubbzU+3zBxA0oBY
OKTC34asv6kfPZonBJ3k5pZVn/89ZZaEneBRX4knWG0xhif8m+HA1REz1ovtKV3R
PAO4WTmezOsftiM+PmA8+h5otDqWCkF7TEjqZRnfSg2ZPCe2XRs4vHpZt+mHnV0V
YWtI+rKb3QA/su1krNg0Em+ZPKsjk+C9jkeiTaGhltJiiQpNcVGdM2cZ7V0aNMUk
HmQIHMBkcIUsQpJT8tb3pSDQYmEgyVhLWsNfGM0m0hWqxKxP6dLO6IHqzzfg2sE6
p65vtwtNBFwvVAZrfMhPtKddLTa1zfa5OOtimvipKyX9trarPk1xQV3/gi62d9pY
MDLA9lXU9zpDD9+lyE6luJCMNHZBEgBR4U61wLSPcCRKEHSNgAkgZD7ow4xk/j0c
Q8UJ11G6URea+DMK7vte3YJ1zi3LYvydiMzoTfG5KOGuSTDGfhNu1kuImGqsTft6
4T/BvV1rKrsGZRXJ+dQIzIdZ+4k1+Mv1hXEiYvtdP1Y=
`protect END_PROTECTED
