`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CHrDiO7YHaFDgrzXUIRvlk6ItaLP1Kf7iGnW77Ku1aUUnHxR2EAww5pdr+lgTC4+
MCp6vVA2kDz+f439xdqbLJU6nufaDijV0jFhfAoiIwmhQD6LsXEv7prqhPA4Z42w
UImBMF6iSqh372ivdSHOlp6PvsNYOmb+F1ytj0HfHPv8stg2zoTuEYsttx6tB1rU
cwrBAnC0ClT4vpiS5IvY0fkChaMQHtACIwU2NtiFRJ53LrQPm2zCgZfN6oFmgQaP
WBSjpGt4z6nxLz8Xw6eedV5Y3HJfD7dMhFkqfGFZUAEvzfM77UmIOabeUVwlEv5Y
ctSkvMZ9CFiJ8R2K0MIIGQxhmwqYrsAgrEcem3LC6DHhVKU28hv650/g0+nsCw3q
WaFUPdtAcMIIDg0pA2xTnV2EjLIR3ksXaajoHCoTUtUyqx7WH0n75lIbvPvBD3Wf
nQduxX5+ksgMajrgFxNVi8KNhnuK0BsatHchHt9ClKsFRQG49DMnxUlXUnaFdf2T
X8eltWsyz0R8uApOCdKz4SZqR/oZ1ygstT6XXgE0YlsiKDZNZ/E7/XkXB5umqCE9
ffs2Hhrn3k9JaU4CEFxWtaq2jLcOibDBNkGL81nPWQMmPAzDt1OgHCo6HYU94h6l
FBE9WZi+r6r2jgTP41kSDAVwni/gy792gKiEy7+Gy9rouixoT0eWpPgGn45UgtOe
3KB3hqxdyldXU21l6jkVDQI4vrBwckVJreoGvrCJWbAJd3A8IsdMMm99wX52oUaR
V0n9wKsEWZx8ws1UzjEN8MRuGLJJa36ND5iRWd36nHjdXvBeeI7oFWKoGYjj5LSZ
l2izxc6bR0K28FJ2Y6C0J9zmSsR8rF4lj/kRTeyohd1nAlcpp6D98DEwhVG3jchW
/SrhwjqtXhk89BYUVnaqyFGlhGlVrKmirFoaE9x3oFo8+HAbI9IDLFUn09dEmOVU
MKfr8E7phqd4SMm+iHqFAy5dqfYzg+SRCzDJv2+WSxh5bh+nhfJfsjQecI91uEKw
92RNUcEyhqGmVeTSLeQ5ebTlgGI9Ry3TQ3YEqSPM+5ie0o7xg/8IbVRHx/YeA+xr
Waa8Y/XLe6MU28qLQRFQEUnMq+0sXvn4KIrIHyEgniuBMC7VmyQfu9010RvkkXw+
QDQcwlAL0YSrqDzsvHDRZjo2LzHUV0GhSud3r6rkTyBWW9A8ufVKFOQV/1gTztAY
HVPLQzw8k1tOLztFM/ARy+3ra93ygwJN7H1dgibYsTSkonjBqX/a9IaG2tPqBzSk
JaxfUKisbqgmZcNIh9qYrtccREO70WFmDIpJUgpAZEstxr9l9yLFs5fQSeK5l4t3
372lMdWlkZ5Urj5nW0jnUvXGMEGk6kfiK+A1k2FdA+IdZDBr2zW9W3OfG4nGB6UD
0E0n6zdp+fdootMqaCSZGY3UxlNqcxIegPvNVKSdWXTdOMUCc+KvPyVZv1h4K0ep
QUhqBzCmy8b9y/gBMBKu4kio62a7HQLZEDPMoucGwIYgPiU4on89JAnimU1bzCj8
oJ7lslSLgD/5PTdVdVyxCi62iznH890ZxzRJxCxlZuZ4zeItfFZhrpfCehcApqkN
0MO7ubrPQO8PDDYjW+gKvlo06l8uuJGEHS4nF/AeHknUXjJN79N11VOpevPfpKY3
V3OArW2r705RxSsraROtH/rbOjyXSn0bjudzwFgj1MbRPNGIUNrOZq1iAFIn6/et
ZTNSbrE4EXDNysJCrFHqPNYIv0DKGW7r0B56Bc2UCYNKRG51LmdH9QNFWjH7/vAg
0MzdN0F8N/mVp8BBub+BCdSraI8Gmh/Nd4ngg0jJyz5MjZ2arN1wRl1UWVsk3s3N
0FxtGKT9xwUHG1v/4eLHaBgnncPbHtUUtNKIbEUFY1U8NngXZuOg+S9dvdcWm9rk
X9kj4DCgkrqzOIAIJ53mF8IYgF/tw8a61Ssa5lbMNjacf3+sycKp6YpgRjEOzL4D
OenSn5QjDjBfrmwvP+HuTsUErjmU9RxpulczHhjXoTOhf8+XIF3SIjlfeE5zQmWB
o4QJI7PMmLDMGUIYxCcWCLv++Mq1ACVLMgLsFkQUBXhD/vX4XvHx2MQl2Uyl4QQZ
IRfsSP8gUXEN5XiGQeKIxnNK8p6ZOjBf5hISmKn9iceMmsKdxYqnBd3GgfPYLHeb
9Nyn4ny8Msw/0WvFPXpaDk8YYWQjWVuqHwIx7ltKc0GNaGXc3okIHiQEj5SuSh6C
7mtUOPHDXHXJtu7729CYcHin5AWKFhpqgakhWb7fohM5lOQ8tCJhLQ1eLF0yXVer
kYMAapYV7HoAPsMLu1COjLniyj1V/e3BiLv5//avh+ysRyZ5D9A+xkGZYgrZJJ3m
RFtbXhLkBOfWQQmJbLlMi2mx1T8mhrnMvXOWzP06UQ0M2uUpgMV4m7v45zmhwEkF
6RHQura12MXyMB+hDD3gyWHQVKdcrVPi8A1OU9i6LoScaXxqNwzfpm/dH2g1CPxg
ggldfsdV7Xa/9itMUNkeMzUEHdcEVcM+fIaf9MbY34cPYDY2cI7n7qCqmYwo5CxN
gECkxu+j70NhvtHEyK90ZDNyMcTVkjoQOHAk70NR34LhjGWq1sOSfmId1NsSuzc7
grpdv0Af32yGfZIRVI8PU2605yILueaMwFrP71+HoCeP4OpT7ghrfb6qnvc3knYe
KeVomimZglE5Al4GLRmvVoyXPNvXUDE1UixcPOaHxeWRZE3TeO6E89XYqZczReOn
7HAin9OilcSHOC6in2p630jsFSdHGTdSxnif9ea9d/S3ENV5ozGGNeyQQ75sUc7J
Ohr+vYeGRd7+YINvmeO7lgaa9RhfrrhW0LDjq/vPSiqVjWDlAvTwLXHDCeKkvBMY
b+IqKuysC06vVLDUPcdXMNEAS2MSuYKEHWIt/+vjz7CFGF0Svr9q+4FIUVkxVkm9
eaRrcY+Zm6Ixx6A55H15JTxjr9fNvCF8mMDnlR+kJ7qUSWVK1TlAatTciNuyT5+z
d5ejGZXe6RtvuWpiRucV8GFrItFcW6eF6Q/C3DjNZIcrmTCAbafF+XpB+ybpj1Za
kI0IShAxggGjpcZal7TmUKSLaORYca4SJpgNVF5E/sGhO90k0xelkn2J05Szfm28
Dc1Bv+6sX0NLmr1mhW7M5UkGwqIwM8fQxSb8egVVsfF+iGuP2pXgKPiNoHBog9Tc
MffVTm4Tu+bOMnzO4BPMpTVId2v0W6c0JsQ/qXRUuDz+H4+J+fq2iEQwQ9HXflXW
1TL7VShY4Gbyci79T4sfZkpw8hMhhCkRXHBiLHeoP1euD/q4XVULxpKQblwmgumN
1RfgAk57ocf3tGnRfNr5S/lw7sQ9QjvpaY5EiQoQeQUFT/74xImVHEbRpvK4MYdB
eXcTApYYH8qyCeB781ZKo+uPESnvwrcLhYOKMp0M8idDwpTFMog7rgQPZJVto0tR
Z8y+ENjiQ22lEnDqG1TulgRwQMiB4oO47UXHH0U8r0Aeffj0g+bAMI3DUfQ6uzRC
ZsWa8oC+6YxqEhZ/HROqK+dwqfxb5/1FmOTAuaxMBz5P7XCcoDzLEccVo+zkyTO7
U7NRuMZjF7jxM8Y7lqvBavG2mwxYlAN3N/rDi2LE1wY0ImxKX1+h4FZ/OrI0Z6GQ
K03RqOGVnph4UiGHE/dwV+R7BagzcNPmH5/Z18PTS0HZ7fQRxdhG9+oIaU72d6W6
u+daGZ+BI4haHDKPEsWS38otM42NeLglVPSV9A9FxX8XqsBIED7e+9miBGEmUfu/
qTrHTIc0daLM9GY2+kWG+6uTe9tSZV6XnjBISHTK0zb7CQVivY1hG8RIdAbPGdtT
cUojDUACFJr/lDQtS20tRQ3E9smXeqw3Gr0DEYRDX5iQ5qo1nBiJp2Ms92LVGSmx
DhKBHvxfQW4Zo8/P8dtw0jfZhoK0q9AZBxyx75rq//2pvlnoZHyQpWKUgVRwn4vp
bnT0naGEqaKsW1JJF+VqpJLTL6Dt8eeDfFtJ+lEbOOdiSxW0dlwC8Yw/pH5d0/gO
XxXpTLSP3SBR2zEjd+4/Iem9Eb/ewwXQlTGDDfDrod4t2Q4N8BWG4akUhcUw1J7G
qaknfiElbuy04WRMBdZZkLTeqqfFbo9ravJbSjPiLrDAWx7Ef4RVSL5yLLtJFs8K
yDxA3+ue7c8NGGi23zEaqMlkD8rEqDoIqZFCHzE0Sy+IR/wKJyXa0GNY+yiMAWA+
LRPqOuFika1c3trQedu1fe6yUVHDq/IUg+2wHw/GI2BUTDP+5hFky6J0KBSwhAHg
PFTLy8TczkaER2HmxkjKJGSmL1xqygA1lZ8B5cG83JR49AiCYDd1/TAfmFIepI37
pWARJpALds5pS0iaZEaUwOrwLVlqwiIoEs3gxc6/wyskYmQy1feqT3WgQsyc9sXl
h+FnQc+ayjY+kEqnoM9FiR7fNZRAGMi7DtpoO6sAQxpW31fRKibxrB0DEKedp97i
UExqusRgwUDSXulkXYBqAryvYTp0Rnu+ouLB2r3snJsaZZxHfE+qxrcK7ctRJTc5
rw5vNMxRLdKKvye8zLAaOobbYe36kR78wfjKEg7m3baWoljwdTc7eu0a0loD3Cpd
2rmNzRRcxuWTsJQG0H7Jfpa2wQbs9cUTtw3EE2NVTIrmu1puFegrBYFcaXNYJwre
24UMOG0sJrPmGl19umhc0ZmFoHpgcfoDlsAGmRyj/5aoC2ZvPGmhQywAXz3LBgMq
PkAaBa5iYZV9AXVpq5iGoRuHGyyuO4uXXlM4yAJrGSfreM7fCSz5d3B673Se8CpY
qDXnZ/uWCVg78QP9nz6euKG2IijyA+xgKvSDABFSsQXZshvw/brAA5YEdxBMwH+3
4AgGgEJq9JDVkg0EtgXRz8hd/JXeVg0c0+NuNkaZSPlb0xhtea35V/xZ74+RT+q+
0RMYWF6ZL78gOJW0l0l8BDnFYi+Q3kDwNsGD1HKpAyVtM5C4keTG3tP0ifdFFJf6
KrixIRhBA+xI1H1maRTMAclrYH+HnOv7AnIANH3txEkjuMe43GVqHl/6sW2Xlmzf
V+QdhXCMNzhhYrnW/ob9RGy2jEBOwN8xUYi4mFeTmO2C7/pCdK4jM+/oxWOrhTh7
DFCxgDtPhZt4EEh1VcRZKcHUAlcPoHj2+206CCR7caHVjctkWaPHPDY2LP8pPu12
A7K4S8rfw5KAOMsBK9xAdHaEcbuKTewL9vP+aF4RrJVxySY7WZ5jOG+m5fnWg7d/
KzjUZKz77E2c0/Ae+qbusSeni5YoGWvd49ruwIbm9nM+/jbPIP+ry8D/R7Rimqoq
dsihCvT1bKi9eIAAhnMdMb+PhcaGRZQ2BtOOZ+CqQVGATKKYcujH9uTEXilmW1Os
0UB9O28bJm4zHx/opwMpHBXfkwVRetRjs4EI4KxQz/aK/vRLklSC/lPx7EB1CVNI
Mstx/AeVrpXBNXWkPh/zZ1IwwbeozRWY0H801UiMFdr8MDkyEPL5biJlC19rz7dL
x3d3ZMDZPT3mn06uTfn1lHFydFG4MnETUT3zp2N5cWXEhrlIRBv38haRrn3BD6HY
q+pVBPDnYmpyf8zOWYKaamShpAuNtHUU6uDcIWusL/7BatYtNvgfnej69v337C0e
eS1tM3+sIe2kyH1+g4Cy1p2smfsKLHa70sfbHS2MhaN3ZFoBo75U19gkVId0nIk4
puu/65LXfX/TEnH9hVXwuMK9ZWibTe/4r75dnWolEMMP+V9ptB7arg05y+MVg8i2
+rMaNkqTD3yQoCrB/m5W2KQnDctoyTagR05bCL+qy70fuKq2SZnIdU+gtZcubH3N
3eRUJiYsnI38l4yNsgLPkjjzAGICzoHPu1AJDyRYyXqt7gfzIq8XCmBkQjXcUkTZ
OVrDAK7KnpjJH2xrdOIV0MwlAKzSI/W20N/xJB2JYhR+EXKpeU08/FZ3n2ySVo7M
9C4K/lrrVqNC6QWvFEh09fH1/IKMNwDW7RfHa+jkPFv88L2rz+qmaOc059fUbvUu
nPEmuJklaVyB5Bm0jFO2YGFKX3fS4L4B+ZXe3q+/LBhBBpRbsRWsZcE0TZyBiBsN
sduds9V6o8lBhJsC650XBcxJHMYchJQO/6Cy74d6ECh0FXNxkblwdaXj6Oa7yXng
A248CkRsUh29HAR1RwXiRkcqC8J2nY3Kgw8PHYM264MgK29PZDA9ISR0KOJ9eIpb
75S2SS4ktFYoXGQXSJ4wAntu/sXLvxFp2Dpx7amlEhfO/HN8gKxx/TNWVofh2klQ
0muivDdFU4edjaJiUfy7MhU+vWMccE2viqF3ImqlXVW37eO9dIqHrYftLjZr8oeZ
GBBufJmgwBJ/kS0DG9zO471tIiZRM/ghPBE2qdNRSWSJkPMIMLmbxexc0NphrlBr
8nmmIgaVU13BwWFwY7HHIATAF5oNjZCLPEziLRycNuBjHxPDgkpH3dGtTlJAUX1d
i2Js5blvWUW8/3QcZE6eCT5l150wSVsam5+CLElhB3isVpthrE8gdt3iJrPsVs3G
tQ9FD+70Cp3QTSdf/nwftj5515h5Q3Vl0i8RavbhQwrlqp4Uq69Q9sj4Tljm10pN
56O1HRsroB7saYaCjFUW97UNgXBg9T9xyc0TKTTKTOTM/NJnbdzfdUeo/m5JlHQv
nceIxS+7ZUPd6aYEcbUcQrpTs4hTj+biDtuzB/caxnmnuvsoVuflagS1yeBdU4Ul
yjI7istHQWh/Y+T4vJQC4KHzDq6EeR7hokRWa3wSeHPquI7lbG61XBJMzj2bIx1i
8jZs9n9KVrg49rc4hiOFh3/TQTriIlsPYfTaGSiws6JsPSAwUtkkJCDNs6ViSe5x
Rb/sJSDveiNBnBz/ueTuUsBLptbN3nvzb9ySIeg6gG58Y0N2pAGYhaWFe5P6Yc3D
7Gdu35+f/NbPm9bD77JtXIbYudsrtCi2HpEXWxze4K4xnWY/WrqRTwmVRZkIH/QU
x2xchxP8H32UX+Pi37wQULTMCyIgFbEypIX3DI2YHWNSYasM54iAlHajkiwm1vXr
KuZvXo1chHhdV71ic1sGX4Kms1siX20DiurXLcOoJ3u+xREvODNQyOp8TfPb6R2w
aDrtlJQGwmfG4b2Kkc8Wjtvlwi66gI+CwIvfPjOTdmGaLZYmmPOWmYvT+7i6KzPb
eNFRH8bvp7SwC5uJXtI7bJGZYmSy8k9CfiVpxtbBo9Z8qaGL2x4g2ZbVY5FCdW6L
IuGvRlQwNgu/+pJVR679Ey0EHGq4AKiWYubwwDFxgyubktACaHxiEtBZvKjZA2wv
BujbWMJ+X0dSvb9aZYQSS/zYBY5DkX3EnzTvvXVJzSORGvgTJggaSprvwZqZKN5N
06YB7f+orN/7S5V+MdVFi/ZkVTwnSYMOC1a7kKdbMJgNY1KRLkZuxBBi7Q5mDWNa
8bXhYGa6R8ZUx+nBicdNAdILKc9v/3QvGUzaIvhEYkClurKlDd9If9BzhkOQ6mR1
VDzDeRZAzyugDRUHu7nuef4J9NWEptG1tvHTotId/za1LK9axg7+/fUsYGB/jrre
xBnP6YrRP4//Edkrd+wvooV5PCPLcXXUDt1CvVM96WK7Q5yo3tcS6MTIWiOmNxJL
DPpILSJUYh6KDO9898PiCYVN8iAL2yrrm1+hA6DBlaVfq9J/kBAKNtuTyIYRih/g
7SC0iVUUTkcCrFygsWSm+Po8oTTeTkh3h51i0jCmNgNNlK40oclVkidM7HoGuBoF
d78FzqVbAWyhc5LNYHaP+w==
`protect END_PROTECTED
