`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQHDgRv/ch8OjLDMHQNl0gCzdI9eOKpv7eEtIKIXk1vGERadZFqF/vg+boOwJx1J
hElMaeSgT+YaLlrN15p6eJfC6F7BNcEAU0vZyqX2wpxNid0Z1ULFs/6H074yd4dC
Lk3ucts4mZoHBqCbBwYqFye1JnUnBOanqo5YQOCRnsN4j2hSzUJ81EH9NT5qj0BQ
pZ5vtotofGSeSabXdecG7LgKn54+JKKwFNslHVnVjKBvQlQvd4vRS9qJUfBAcusH
EwVZck58N4JXTJDMIbIPC73qTeG4wIMcmMUeTsLI9zjAbeQOTm/VQsSCpPvvRHQI
vfggrSHbkCAnItbcZB5T0IJQOhiGud5VmC+A3a1KONOKhjk9a+OO9ZKOzvNj5D4I
NWmA5ywXsLIN3icrKwJbWWNnhrjdXxn7vriwwV5E4lk5WVJYtdBIsfqm1DXxkAi3
/k2qvf91kEDNANelH7iHbuA6Gjz0R2IzEKaQR+xwa0a88zLmrYIyT2NrDj5nGHKD
V0Dg53E+ZWaTUTNqD+CXqryst1WaiTz/SSWtVK28CqzV7TQak2CG6+cuXoYTF5iE
zrSXuGl7YhYqGdOXjrAZq2RkanLHRQf8zJRxdGO2GKlfSWueY6lNpau9pMSlDXD7
RXtiiBYtovIbnnsNa+CcJ/C8Kbc+wESurP2a2t3FOm8HNfzOL9Fb294LqwdSmFSp
C24v3Fgyx+GFx/amLAABlRo5GsBZvE8ywoRfalGUEOln01F7sTwtrJZyKiq69Yp5
s+k+2HtDeeihhLdoKkt2WoFDe+RL8KMVwl96i++ZvwlocZLmSV4+/IhcypdCxNo8
O41J1pjJvghUTU8fBDRgVje8FGJQSu3/BfeEcAGZu3zMrXWVWUw9vYTToadzCYts
l5OI50BWYbYnSH+hGqCiCqU08OCAYg3Eaj0IftJ1AhZFLvNYp5PVHReJbmxiq9nw
FllX/AqqE4+Av7vX0X+2pt9okcMsmjDgvGjOzwp6juQIW07hPJwhotBo2oe0S84k
rKdLAnjIT6C0Spi22nA+1ofStZLF0E3XWVxoKNL8gQz8lnuNvgql7rVfwG/Fk8Qs
bsttsEGZD+1tfUopgKbg2GIjF5DAa+b6NQGWfZCnUP8dIpggTo+2gDDueAwLqF9R
WDGaIgiY7uaRfvTu8PhSuIjUiJvEGLEvQIWhGf1WFZAhw9YSFjwxA7iAEB1GRckV
Kn4aOAO2rj2kMleCC4Oe+2051z2Heo5KFB27MfdmYjx/Ifg38AmDa5An6VXc1hgc
0Ez0MKHMI9GLce2Lfci5BbP/odHOAVIjLK6m8uizbhMzhUb+5R+58w+vabKK78un
RrIghLFV4CWfLEwRBgBlV1yeB1KYBGL4tSZkHGpg2kN1VRDgxp8wdWkFPIQcM3u5
oLzfpaeFzTMf0LVJqLOLz9AzjcLxzv7Vkx50hK0BmpnUnsleoXX7i7EhP2N2nGxM
+zGzG6BshjDY6nMCWiOocVT87R2Jtfez1PcOlYctlSdExhsmh41thUWlQ0QuPo3t
anfexZdNCSH+Aq84DTfmd2fKKf+vSIqhU1d8qjztirF2dKDjsaqwb72T1kRHc7mI
/Tmmln94e26okD9pZDq37DANuWlES+4b1bkWMX8IWiQAQefGOiBMmNqti2+oSYKo
gtbvlziRR5DLP/pGhbFzMfHyuHNaUmSeGd6iebB2wudt1R9UORm5ZvRVYj64L4vl
sWJlPzm500B6/Buwr3Z+QTN5Ge5OMfG2ulcsrEO+WdcaqbrdwtlH07XxZr1FMfoV
N8Tnlt3XjpykD5vQMpME/04qt+P9UMB02YwqQ8DmCIVSFSb8WmIjrWLHw+39AC1a
V5uiyrKvCFc39VO+4uTlcYv4X1dQK8ug/n75jHAjx5UTxevpo1zIML1aeBDZMw68
CHaw749uHCaOTyvzX1L9xwQzqOhzlPhd0LUhjFyQ1dO0yW/gWyjc2RsRCjFcBxnS
VjmTnwhWqh3rDlMcHpD6nGNY8+QgfbnXAEKiY7EdL/AGMO9CUjRh0iFWvF1EDxgo
8kR4aG6Ad+7r4cNHdzdHIC9DXcbpLkCcJ8FYTtEGuUxes2POmsS7ncNroXvGH5y7
f38AGuHdEAWDFFwpCtE71hbkU1yBubEWgqbqSihin5wq/bAO8oHNX7/hTeFxxdsh
1/vpUftWAXoky7Rh6XpbyC+W92TAB6PGsmGycPEupwUL+GPZOnr5eixl+Gb/0bAF
q/x9WbIhWeWkPGKrqYv8LnfHq6h4dFEQYoWKLPZQe+9iIjrWcXnoW6c+ovXGHj1O
CkeVRsCxS3O8lMuf5e2YVTrQKIvjdDgp0aZ6C0a/bjFLTwKIxHl/gVHUN1AhJGM1
FUopd4QO/pSxCBsdcz83WbMgcHgM48Bpbfa2bkOJc7IMeKpha/nkCVbH5ru+764g
CO/N7f9AuYL3h3ambcJQwX8cdsr+Lv9/aUFUV7neEY3Rw04VbO1dmVD5nvrVIAmZ
dcJjuac6loyQFvclA2ZPROTNIxu8Pz4bXK1Xr+z/b05NqEzHp0e3lweNlmu+naVP
eIHCDR9CXWLEOA8uYoXmHsxuarKau/edjoTLqdW6bF45vOe4NteO3NN8Qwp6Q+Ls
DK11QZgiuseYW/gMdRmq4eGmm0x0uQWYFp7EtohVc1SBP2M2e3LR7oBqdWBLb81B
3Gg+zpO6QE7FjcJeIBGdH8kDZZzD7W+xEs4QujjDfpt0F2HKxmoAhhrtRSQC9tLs
inSsp5YWhethxVSxcRxT9k0Q9kL+UE1++sdyA9p1RKGjqSIdpiY8FjpuH60NqOrU
Fbh6hHc0WWjPSg3hDLoHv3vkbEivuHgpDaUwgufsoNR6mi+zswJPUK9a8IQ3J1HU
3A9Uy0wLmeDBFRzz0EpcoyX4leYVdQa9tPFJVD9cmFCUaEPg+S4ve+xcFluVjPfa
8DxwgKha8GMMZECyjGRyG1x+cA4AvdXs8FtDSPWVbRJ6QMSZo4LKp+PGwryxYr7T
j/fF+MrjdevZQ19Xg0xp+2WJFkbtF3OthT7Wyh0za3j5/iybVC1k0nVWvQTzh47X
CRpb63GpRFzY+2UFWzYqY2ZwRa6zcKANm0TZAJKHplJXWP3uA6HAhyrwAtyHDvl+
AtTE6fgzyB4SBvMwPvX0l8W3rHyr/Rq4a3ZRjec3eCf/aTxP44hkxQxMlpxBU5lp
1zkBq3ejjFqbIyhUE93moUfqP2xcVdu7+yhx5X+Pu4Pb1QYKuOiwHe+5X+lx711A
9RWYVlfq0Xp3JvNC8X6q6wtGaDGU7xM9gO4somyIQeXEKXdAjI4zpZ/F0jC+Bq2G
JeFnxtlK+rqj7xdKl1+rxktr5z0A0q/YGCUbHz4ivZ5ua9/21z8HrtLpQ1MQp0xX
fyrmsinUZG9l0xI7Mf8Rf60bgbQjGu2zjAwTPJvQqhrSf+5ye26IMutXAsxQDIT8
3SVTgPxbjOXMxRqpPggVX6GERD376VkjVLWJqY0CqVusYNzC199rtX4vA4dZnE35
W4207QMFr1Os5MmwmCLThJMmjbBiIxzdzjnuOrLgBZLiOKFpNpPrpDX8/+uHhmf/
4YeudIGLieV/Bv8hxahMwUlGvRZBNRHtqKp0310Sgg9bb+gb1SDQf1+EoGd+4GOr
5FJ1TxT/eKhsJmvEPefGrkNFZLspoHE35wtjfLEV2IA+Zkc8CMUM2ctc0O9vKXfG
5alvB+cxng0LpgJseWC6OR445ad8aqbT02ONKnbjtRbzoEtEGTytFWHWQBQw76aM
eKxl6W04Pedb1I8A0ozL4/q17KufEuIg7/uvFXX2IR/iRSTkBl+FrqLuZiszKnTE
Wj9b4wcj0b/kDFQ51Rsyu7xZXAAe8XOIcY5d3xv8bXrSOngtL00mLhrtJXP0i24J
U3DDEPfhHu6AsDPc3jvycStJ6y1h5KrO+tUziPL5ADvSF04YxT2GhWN7U0zSOAUn
8P8DgJ8TIFq6auutWyNlVq4t9FPot4v8soaYPAm17z3pWcYDuwxRGw8rJHFGWY3n
DxFC2luHA377PffzV1fQ8RGarOHqbTZlwYUysbEzUUEuaPckUnCBzZiW9vnwSHpL
hwa0oaBGeVk8SLaGQRQAiHrddB/76iui9b+UhKFFvkho0CwokWVFeJR2UpsTUM89
aVKSu7ahR54sWGuiuJ/VIOYHHRdQRlxmFsiquxwx734sltR0hi6ojmfGCWpqI23B
1UUWXk23PP8B7eJUL+lXnivPXH6bpEEC0dKwfFne9hLOWNaTrCA87uN1W9JWBDYE
jLL3xFfEOQnazXMCpmV+k8r/e8LgRoZf7nj+DF3xDK9J7JO2rYmFGAlKWQm2A/MX
LMdDkPeM2T35YTzf1DzCSnK5VnVud59GNcY9sRuuT6b8hgtZmb9GbjnXUQE5nXRi
yeomqQUL7iL1luCYNW4hK4pMbI/7nztlKefbDhWcYabAwtNvK2ebpuml+vPGIZCt
0daSjjC+/RUHQEEJhn7Veir4zOaF2W6Y5ydBezkcBIPX2QPZ1eeLiW78ZoCSoCKe
0kRBtj3Q/5F6UgNNb3c3ULcizHN88Xjh65EsVf7LPxkVA1G/OYrlxCfpjvHBI5UL
DCqCfjJx7OtaT2aBJycqc3G3hHwZ67mZGrMAw5GOpN5rsT8R0WsQVgaCfC861meX
mS1JMyLjsTD/cLxq7o3VTi62Ib2pQRQ1IGfp0FlpQppaQhPldxuh9ggijluVHI5v
jD/lMeRUT/HLMOslUfGtgGIMhPzf7lUvEHjTdfTQ4BG6/WlXn5nDBNhebFt8KtDE
RYKEIOH0Ms6mvmhq4sd4Sa0rtJknFcROfUwEV1kv2JfR67a3axcfN8fjBBHakFdB
ikFywVeTDxWrxr5dSVzvq8c1LVXfldVzvKYpCXSPHEyLXacGzscB5Neut39IfoLT
0NEXNAn9zJZHNWuMcAruUh4xlo2/sjiOu3yJ+eY4O4gMr05HhSrVzvVPmPuOdxfJ
muUs6fgUw7Qw/B5wtQAoQCfyvfTMyRWX7JzYPfxqsbYMFIC0uvD7ddtJ+2oUjoTv
be/RVjsXWxX8XncaoSoHLoecvVGLpP3BnOoxFj+u4G0DucoQ5SMVE9lFHTBDj850
5FwyLIMRo/G6kFxmSH7wp1ELhX0a7Z+kWl4jTQp69onseGWkdpEn36EqO2N1bnez
9nV8m8vY+uCX4UmKpiTlZimmf5XBXQ4tUH3F5jg/lqMU9HXrUHOtE12fhXBDDkCr
9VaWZ27bRrnFJciu7270u8XPd7SCuOijZuKBWDp9HwX15AJFg2RD6MGqgGSR5IEg
3zRdwH0kKI+qWwq88MMEwSXuasQVc8d2tQ6XuiIDehD6lOaH1NfRfKyZz/N1XojL
r/hulhzlTgYNYYjDr4R31rOU+kUuXMOj5DMbyknGOCUN9G3SJ1quB+SE/OJTQk33
7HpnS74b/Rf1O0dCysOGr9FF0wWhlx0bmpc2l+J0X8Pnfce/P6OS+fUDef5Fzt9w
sAdIiQnGXw2Ot+4AC0N72X7om0A8YBMIeOeO2NVLcC9tzTl7dzhsZhw+r1nq16+m
++lPhn4ObjGTIGIdLKjqciX1G+iVmVtREJYnqY4ngtZbUOS/oZuuAuKWYUrh+gus
YU5bzH8ndOChdEQ5o+Ay/uQ26qPdRezRhh2CLUJi3+lsKWKUFkRJ7Hj8RJ+gNAvs
pB/hixc8hBBdeKmfwf9Qt454qRpmY8Dt4qwVgjVp0N8S7VAa247Pgkg9TwEIR1Ug
tFQL6St4b06yTNNzOUTrjNKVl5c4jVyuSPy1N6vKJ3gncwIRhmUr2NK3rMpRsSJ/
pLmM84hssHD2WLWq4diLhIDoPTNDyRIdq3KS1l9UhuS7fP2IaOfggVvj8WGP3LeS
Pi/5yavNXEXiCFbWlzJSSDhsqGMpN3E8I5jHSsX877aV6RPuVMG1s8ki5sW/ix9i
V8TSIssdO7XkkTe9Df1p9wXbfpkQuVnsAPpYPH6SZdCKT27SfkikvCI7j4+0BWFz
PPlQVTzEmnUjgwfACZjs2kE6xwzQblzZAg9wbUSdBZWq5SxwqW5yEw46elGOxB71
QNNy3yKWJa6HRvwTko1bo4kKzkGCEP82inNF4JxzYTYa5kCP2axED1HKBFU9sCxf
s4EypJw4ONE/ZbEqH4LPiXQD7aJlOn3HL10QN1crft212TfOSJgakXv7sieWduaH
88Mw7yzw0DP9vbDfuWyhMIqwZ9DXzabZWQet3Z3lsxSpvVBeIHuSfweth/Ml+hje
EuUD88oCgLR5Jt7Fb51Tzvk8+lHiQ1DbVUvmUQO8LSK7azYoMsdD30Nf35hPnyLO
e7WEJwgctJ4XL70d9bxXNWUXqJyr4CxUqr0JV48GNiEFvaRXqXs0TQSBCJovenRP
qvAUI0BPhp72fQWR0IBBlKzZtUBoOaKoOG+gzZH1R/Vl2CK1aLmMei6JOBy3+Ssr
bWtJIw//A13ZYNxA9ssbmT+DfbA4etsXLb1zByYtDQkFkYHNXV/ZvuP3ttQpNDuh
79scx1c7MDEg30G3KZjerYeOAMJVeuoTv6c+lQeiP7quLs0Bae0Jv2Ob88P/y6Vl
hPh+K2LKjGZ1pyndz2UW7tqG9IuQGPvNs2ynYeOH43AiTrQijmy9JW39TJIHrk7n
pAfEvHjEFX+Rg3Xi01yrWGsCd7Oe0noTGbauZusinPDBPleTbdHszTMalJAMgAe2
hwE/ElVKSR+e46XA7zNiNQ==
`protect END_PROTECTED
