`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5x2kAn7GQ3wDyS6TRaS7FqyVYcCPjWD/rYQVFz6cfUuLNAPkxeNXpvH29gmNFTJo
W8z7vScHiBxrbAea5Nhi+hNgGMl7lQ19aEMjnWox3huI8++weBJ5VEF6pyZhv4RY
dmLQ8YZ/JtBNXCcMruoLSKbDOKl/2lvHHj35sGA4ZSEmBZzg1/5vOgzt1ErkF2cn
hvRWB6c1AyKLfgKwBl58i4OO55qxjEP2c1/Sut9bw3h7wmUP2yiA0fRFB00kpopg
ruNSzjGFoByRj+EnFE017QB/qckDmrL4ZSp7+7pMS5rkWsSKQEE8w0NrCtlihizr
KaZaKopdRRjuevgiB1xiPHX4NvS38Vz5+/CiJneMshj0Ce6/0Raqqgrydsd63P/T
MZz+Chzh8XKaSaIJx1o2SUcWft+Dwguwp1pE5mKynWvsLoHd3dJBf2vaD3f/fSgg
iTMDrVKZTPddSxKdyR4TvvwRVeZOjHSefE++8s/meE5gsuZztOnPWQoPWboHscyT
Sm9wUqiTXcHQhtcN9GgXuQ==
`protect END_PROTECTED
