`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7vh2Ff4VvFhmwcBSldIFPkSga0OQv5ob66Zh9IgEudT2cyM9C+y5JvJ4/zy21IC
I33+OJhD2IFeP0jJk4tq+cImvzW+DQcANjBlBmMKqReQynZCPFuzla5/FeobKIel
nyKX8iXxAzOjOLyNpFMTGt7fLRsd7Dl/rMvAyZcCmnQNpWlce1z7o2lJO3exXF9x
U8MXTJrUkTo6lzg1hOFws5N2HJ4wpwrsb5hpdG2ljZerpppTfzurvxbaqgwS+ROG
f7PCan4hpHbkWuo3w06okdFBr/rGpITcEJGI866jx5AwyJ32H8UXrzFZlGxJGLRW
tM7U2DOxLnGAWIZKTMEn+khijMrJNIFxFTvAh7BkBz9Ezx/ufFHM/R30DImBBL3w
bpGchwebO4IYig9UBoEQPhuGVq+Q3VcJLeKf7pYoTgAgJH5E+EbA2B+bWN+cKgzX
61BaKUZusO11D5/jJ0Oul86LDWo7pdd3Vp5DDTFjER1ljD9gnHMcRjGEZ/blE+Bj
I3wRXRuLQy7xrl1gUN/VlCIk1zjifRsHKFvBa1XPMqbTRlQIegu5ZA0AgYFFKbCG
o/wKWICq4V8o18IeX/oOBjHcuWRTnwC8CWBZf+Y98e4qzpt8D4OQVwTIpXFL93bB
Zc7ir/ipPhIhJh9Fqt9BgcHu610OEQIWgaD7y0n4bLpZLyJXki5bKSuTqVSuVOQj
T0MeAF6texqJaOuJjYnMvY8HPK3EGKdQI7HrXQqo0r2zYY6DmZXNa7pvWyfRsOMN
fD6Ts2b/5Q18AfZKmT2l5VM/NK5Luq/B3xf4kLw9TtwhuuwUKtFWdtuGCGPEdryG
gZqDAye1cw/l59Gn0yMAjKvQcTH6F2pP+ATzHzZSRTyqTDlmsTbx6pMZzAtUtMAT
u4m0sQd13n971+nmqeNWz/uKauviI17pCxEL05D5HrNIvV8g61YnU7s4JUMT3+d6
S7a1/b6xztrokUAYV4bAbTYw60eo0wtjaXtLA/E07QhE6L/qxLZ2At26q2pciaFU
y96v/cv5RzDwpi10AKGr9j1Mm1b00/OWI5H0xctoQB8biDmtbKsbWgxKrVGRiIlR
iRZZUKweQSyQVlYQH43BI83lu4MuTKcla96abtJExGoIijVJM24Pdzwu03GmUoAG
DE39CZPghGEvyd7cup8LIvQjf702DI9DOMlLOZGmeEQH/NJ4xmH9iuzjomrIK7mh
sP3aEVSnU/nhAtP4nMohBkCEKXwuY7Tnu/7B8uQSv8sFy7mZv5GkT4u2vd3FoyDX
7NgKXzyfvt1PpfvSkTdiOhDPKqHjq6VX+zywgS782qSCRL4RMoa3TsrH8wZIZcM3
5A23d8z+RJOCm3shipNNTfdktEr33ng4lMfbsIRM8p1R/+RFUTVyg86uQyLrycyP
q27+IuWay0m7Umw5zx1Cd7JqU7NBmgiebygZJ9Xo1Isv4SwsKi+J23VifXAaJ0g8
hxm6KmHgcPFR5TJ53E6eliKkyYUYnPQYmapZmARCZJo=
`protect END_PROTECTED
