`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dvqDEf3OwAkCcd4zb51NVvZrS0YYysqQvDBP3jH6CG0n4KwxW0u+5OhO35f09UPR
6Cvxyg5/qvc1v2ZK/PL3F82VBp92Qec2m2NwZfuvYWpmIYSfQa5d1ZW0KZ3GV1nQ
dNI4nyAc0FpcOe4zeIeZ7W0Fpe0jwhcMF0hM7F0c/VwtvNDY7ChHqB02agt0MSfy
VkCAF1WpT+NfuKu+qPmNt4pHQSqfgFiOWJqE702iGAPw0JFma1dI5VFgArrzUgZj
Og/DAANl14qdCgCea8ntTGFF08gl/5MJ0eUCu8/SNMQX8HV8wdv4efD1pFSjS/5l
y/XfXFF4V2dhQcCMtVnL1ZIpzde/MYlrYQTTUeVKOjBNllDFXFVcsjmwGrSPkAU8
WkE9Bo8U87eg7GnzeH9yuPBuDKkPzQX3510WhC1bsBls7Yg4J6NiHAfu/3HN4JR7
lZ6D1Wef67tpnq7iGb0VzEyOG47pY+mVvOlKY9vRSKXf9v1VA2EPMZOCq5NuE0oD
ws9LRF61WYZUjK3vLq12tTJQloq/vdfvcMFTAnncwFTTG1KRxJXonyFfSV0CVlBJ
ua4VnJA3V529gjdjV2MEINH4A6mZARNWzP166yMHdqkh1nM00q0gbrICsJf8vIB1
yrhmeY6iXJxCvMcDzZp1ooJ255TMOMyTMK7Rd2VcUSdroejqwFkTGZ63myrtRsz5
i9KVeSBGcVyS74AOofEFZtuoaoEHoV5Pu4NyQZDRCrOYx5Y+HEZxn1QGOMeuQ89O
+sFiC1FK0MyMqyU/MdRBOOp1xSGZr0cdMqezVkZD0pXGqqyQrXeiWSDmVPaiOtoV
9xz6/+ICiSEufuMFF+v4oX9A9VxWxisSjBcu67XB287vOrt9OURGVSFV+CbXZnO7
sObPXl6AKECJ9TMqNxGBrKQRW5HIuZcpnj1rbqUV+QiLlt+PuDQn/22/paZ+3PMR
vWPdIJlRCjOYM9spBQO1x3PE0kdR54YIgWYIcUIG5zYn8g5nY3M82wKcSCgAzSmU
XcV+oGp5m4KO6hHhHdA229KkDP+6EQSkMzpUm5FyoQ6J8TJ00Y0WqjA6ZtMEHKGh
VnQZBCRLFl6hWcclSJC4F2ZYzgj8aJ39U3Q7m4C+DWnoO2NmPQu9CKA2tZTAlCVk
Mk7HshXUn91R/xcgUtLEWE74SQbqqL74GmEdcraMR/PxW1WkJ1H+E+xLK0ORD/5H
ux1BZoln5tmAQS1nQlyO8pgQ4xxhSJD2bLCNxv55YRtdBNYtpWlen5BAairhHADC
bR2KfUNpUtlyoOOEhDjGJyADuj80WdLW3XbWs01p51r97VAISyNqj0hNQgbpQqg1
kqtCO/c6P4oA13VpOPkcVGtead530hYSC+YdhpeqkcWmP7/euL9X8h8Qp97ccrxy
/PU+22m3XZpgGtqc774bUMhyVCA7KngBay6BqaFmWoHrRreA4y0g5V+YoYlmU0YI
XbneZYkAgd0I0bkXWCn4p93MGrv/n1j6wRhz9TPorTLltoIFbqXN48HRiOJOaWne
2X0c6n7G7T/ZFX1MvrAMeqFS9DANC/cdw/wqwTNjvmE1qm0MLjm+u1IzkmITebXv
RBr66riMBBpK1zTbrqqNY40o9X5EnXXL894ZUCgTtsWZab6cm+QnU5e8RbkGbIRX
6utbTVNJzuyZ2aPHmn7+jAGQ36+ED2pzm6UOqOOICt/DhsgcFoiny6kY4ZjRym2v
P6Z5mM+tXajiKi34/IPRl9ENUGPzFg94+73g5+ntGPl+31x/8sWDED5MqmKcQr/i
nW4LyyhUKkG5udGNSmK4gfGtFcanwJsXOCeLNYwjYv2+8KhckJA2cir8Zg8LmHp/
wu/9wnZsnCnYqYTgtWGeAFqIPVMMuC8g0wGlnZhJfsd2te3v3qsPb6e3sYVXTdCM
m7APW7tf//J9r4AhEbZTL/QXF6frUfjp5BKrhJbNmlDjnXHsmELyzl3UrUOf6r86
oXGNA9U3Z7e4jEPFyA+fh63rZQxm2lhWuZOIou0J4q0Bplk/UhzPo9Dv56X+P+x4
NC2chaTnkSrDOe8h6QhjN8MpKj4NKILRimFGsr27bUnZWKg9ur7ZFLzMQhjEwz2w
5pBrgJQ/8NQCu22WBDYcKzJisGM7wy7C30OtOsTm+h/tXFXUsfaVzBwC5tWT3617
3tz/HcSa2Xn/PALuFuCBXLKUmEB77Xq224H1X9CDY1uhEA5lFHSydOtibGzsWA4n
RXtfD1r0UYQ+1wRGPNOEp74h1WlKdu9OCLjlw3HqhG+Wd0aV1kMb9/nLTAeIKwGz
cSOGuPpf6OqRck4Ay2/gvdy5J9vDxxl+ohMe4hg2jD/K/rwadyINQTLtad8wsH45
VdM3NA0qz0a7aSz6CxoxeeQAYV+IzTjBXg3ADF3tBfmCW5ndhaEkKJ2pAP9TF1Rw
5J8pGeAbOhzuf5TaSq31DQWZKfyh32luk/VHJHxXmZizBzsx9sWV1kg3FfJEmWoX
OamVeokUymsFczr517BNH3HXh4sTV1VMD1gE7xKIGuc8mdLJOcfDsi9EKo0zMiHv
A/Mq6eoby1KNxdRWRuVhZAeHOLxZkFtnHBB3PI4DIekxiNE9EELYVD3521e+AT9U
LBLPHt+00CEXCfAGlq6s4ciSpTFFKcMOxbNeSxbJ3SNKeLJ9Uo30hovDvMxbBqPy
D1ODcdZ6xRGjwpvwrDKinOyNuHC9eS018H/ToSDAEuynmOtuAbHg1+7jUjWRI9F+
AVhbtRZorHfLq5gKDa5/3euM9RZU83vgr38LrJ7I/PzDw8le6vrOnnAC81v3ZVh/
YOH7W1AtLz9hA/nPFT3eZpBOdYryxxfuByyLoAsKQfnwa2XxEWrRi1E8QaUlSeeg
PRxZFpQVn6coaQDW4IKo7gKzi0Axz0pb7AjuIAYwGcguWlvvZGXKojxkWlXGVFQr
1NSY7oRg68JFIemlIFwb/asynTmZf9JwLHWnROlyDwmpqlHdSG07ab0sSP7UMcQf
kkrUgEJ8pH6+hHSUO0CqTx9Xwm++ZjmaIOF/3w6I1G/TRQ2XaJz2vutdcBTr7uxP
5QYZO+B7RdYSNQzonLCg+0shhNFOQOgzh8ZwMEyEaaya/U3FY1LDbz8WA7nmJce0
Pz+LcG0THhZSBUPp3rHvPRPBsTTqHm88Vw4i5AeuB8RTZU5pPZgUEZBMyzNxshA9
ek1Lj4lfk7kWr1Ll+a5iq2sf670muZLhqIMN4lLso/7bA+F+Z68qypVbuUaePfcy
yKOL3Gt709b/1oSErxqkBIRNW0HJ+zfpYbBhwyA0m2CQZ14v85OMuIvGF31Sd2aJ
sZXgrTkHYeZ2L8N/R64pwIVr5uZBmNykJaClSS52nXjqhOm55XGwagAepNhH9ruM
cvMVkeJWHBbXrrUeaxaXpMCUqNkNIZMT/f4V0IHdBz1UgRVVsVm9FOecjP+PnZOO
NVWEZ2khXY1ZLCgQaPngXksuRwTkIPw4g0iRft6wUjr75jQbkIQmdsA1AsVeMo/P
OIWuY3nXtPmU14FFkkFDsNEfkgeYmhV+7nTp6jSc/Ti6jlJ4MvvPWY/WHsTEsM3T
TXlqGgrVn9e/aME3m+dIvcbjJLsxMi8SHEQfaJ0ypTQ5tuJUysUIrj1vi24k/X+1
wR9IrmnR9/DSaxtNwrRZU+Czrj5H24gkOFm6VE1JAFC+S115zPBVcdyMca8LlA4L
AVC1y1Zn2XWdTbzEcF5Kt5jQVSea6FjKruqbA57aW4T/KgJzNzDRHzAgilfEQYHz
rd8w0K80VaffxgP/RUNkHGNNbl5CnFfhEHiEDXZVroX4dQSXhtjMwR/S3AN719jW
5uYVeew1TQAgwBflYZU0x2hmSC727LsnmRjwLsCLrKhfa0XzQIfpVyqK9f9eDm1q
20IYvGLUbqyQ5+OyxJfxzawNJwmjEmkHucWIk1HupOwsiRX7qGna5cs2MX1lS9PN
Kjx1B9AO639J88HXetUUmV9n0r4VMy2QC4Xj7BfQLZs9TqqDPO9rBPRwYEXMf/5k
ZAr3LRrC5K9sTkwLNHDBJHakExeObamExkczdm3Y94u9bX9r7luNWL5mzbhCWaZ2
vg9lNsscPUyf8qgcIGlumehjHK41hOBjV+sMDU30sXws2y59BrB8QKdcVgQsgSHh
n65C3DSHs5OM21WMjAQuVCsw1st2jFi3SdjahaqgTnfAaJz200QHz8S9isz5rE/q
12KHdC7+pxnkyLvDLQa7rCdbeO4HM53WYPnjLp385Cl+Busv4qy1WJnEkCnPy/G5
XdhoMYSorzF3m8yi9tLtTaEo23wbCiRfTZJb5puBYcnKkiGFvCvJcjXFVYmmZ1FK
GB6jEzs42Dl3YLnrJdTzFX91wd1qJm+j6QUSpTe1P9jf7MiKDv4Q2X2BSoij1q7e
jfMb8Lk6Q7cELhGYJFvGBNwpUFyjYCsPo8jSPX3C7Xbxss+s13n6si6XYfP/sWm8
GRkGIZoza4TO3nKTZTeTcslUMtPNWcdJMyWHHg2Y9kU4R3WTxJZKF6uc2SEkrfOF
+g5TlwFNwV09sSOJGWEQOseivKNiAAQhvIB7Seyr38uxonhL3kfxSQhtmhBVCo6n
XBjlpn8MMSrlQxPtRvJK1qpdeX/M2VUVgEhIQdAMlvsHlO4YXQYjsL/5c17eiTwV
0S5yuUG6RvcQDlAtxwSUFjAauH/+89xb7is2xUf51NJXA+Fc50YHhui/Z1jHq/8O
dVpj5oC4wjvuoonNVq1PsPxBEM23vY/BtabgawvzIEO9F0SCAtxFh14W2QwOJv1M
QB1ZHKYiwbTO+klUouFCS8gLbsiBGb5vX5qai63kxiELhOWAZuqijiYSDOQ7v0HC
tpgp3Hi18yWBeebhfPOiNjy/APWMMjYhajkjJsoWN0Nj9lFffzTnEFEeD5FZ4cLZ
8Rpj5KQkKpaRhg2NZH7zUZuhfXmC03jbk9qcXXnttnbSP956S3Q8QmP9PZYTIWnh
K4LLHu7qm9To1W+jjZv6sOeFCeuh5zkt92qXKynPuGVxNWd4RQ8lY1xbNoCVbmh6
fYOiVDFaF5ZMTTSCeI01KvudIu5IT9/SqHjFTTI7wUcf0b6JhMyAsLwbmI99Etdu
0N0EwT5ZLTNYf0V3xlRHQWUROChg3yXtZetPKS/6As9cLK40sqjNtitHlkKKcp7a
HNM9xXEohYyVl6uUiHs/pcqCSospVwwJmqHzbIITzni7h/4kgWwV1Hiq6rdmbhg8
vzKTT3jvCSDy6ZyoQD4hQGG8QmihtnRZ3tUrA5qRDGlrabkd6mdu+iRAXqkfnmiQ
cZN5+JYlt5Nbqjx4g1vpXMH2bXLmSTCJ4gcBAyyjBv6SljsKp49hY4NY/Vcnc6ve
mlnoJjzWD5T9p/8icyHs/3mo3jaDDPAI8qdOAPXYGUNBBo0PLSdTdgvsYTlwNjm8
aER/F9tI9xNevwvN6BOMJ8xqhStgd546+vnn+suErUfMSkVMXlOw3lXcGGGWUpXx
IV3+QZx6DhmZHCDfjab1v0s0v9JPL9khAsZy09cJf0ue46pbXoaQQ+2hPLSXei8x
ZoNUOEFqX6ooEn9mobxwFvlViG/EZA/HQjYH/034kbEvHwkGwfNycvckFqPX5ACM
+qFO1dsG80COD+SI/J0tIyVayYC7whS4v7qmVrjnb90xIs2anQo1KRX12kVttGIR
FVRhbwqddxh1j9DBqTgERjZe7w2qRjC108PQflFv9U5hJe8wZZZeNrd7U9uW2apP
vgEq1WnH/s9v4z+kVAEFTdteVSY3VYAi/O8XdaX3HEOqHL9jU8CoD+mrkiuLtvS/
VnXb2AUI6gqGb55TtUbfLYn2lhGOKSBwpBaN/3QBmmgJN/krtkpECKgpAEJL4EIw
WNn3tOYI5hbh+DqGZb9QpzO17PkzpJgUt4aN7Q7mFSacoU9mEc2TEr31DQSwUKXz
FKAzLUBeO0ssuHvX7DagITXX6QaR0EIL1K67p5VLpU0JgLqUVwmuyNs6oN5vVt3J
ddCpI0ceG2eOPjLp8Yi6D4MFOzJn+Du0WdPla3Hv1FYcoEe3K8ePBwybeHI3xoIc
831M5X3J91hOWBWbVN0kGZHXOqlBFwjcdxNcRxuX3wTW2F2ZxLv4hFVeQ1zDkNie
Mdl6Tu2rj7fyzy+JzGYgU34bVmC98ASCiUgtvuaSfG4m5/IdqpSbGiASLsMMKFl/
hzq4evA3p+8o6XhUZreRAzHzU2qsO5+Kf+oYJlEWObNxDr+mCnZawNswM7MHQkSe
bWwIMZhBfXnpU33ZNOvhHn9pqqYWrQ7nV0uZ+xXwOzvAKtT6aCgPEkQA9vH8Af06
wnsJ1/RMMWFdUdv/g59As7jNK4mK/lU16eV4pknA4aPaidvy4KqifN73ZigthP4u
o+9GcE43VzbbwTAcX4yfW5QJwtSvJ0ZosaUxbmOBfCVwjWyrvHara89dvMBkEk8W
rNcB6/r9j+8IgHj1C0H9x9Fo6dbKNW1s3xKSptoHY7+LEiL4lEwyrF0sh2RJlitS
Rlx1IuIYpu43mRnV9Rs1TelZRcM0TDx6P8PBrXf8VW92T92lpMoqoHP9KGPkWAW6
YEEBZ6dZ8Lt2lvyoP9Iot/6u1pvOKwUi2hSD7dxjqr1TMW21dZrVwnxdFEL+DJcE
I3Eykj8ZX3cjWmqSUR47PAUgdsUaL+hTYUX0ki0j+Nov1QB2HPiXNusiklJ9eFSH
WPPT7oOjUDWj4sxL7mgZEAuejLe/zIoxQUnwkUoGFWGMbMeXZ6K3WiMN2TIF7p7M
RsXAXzmSicMj3RPUMJYOHOsqpEIh2FDP0YMcMAOCHtx8RDozVf6UHs3S75DP/uTE
`protect END_PROTECTED
