`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+jj5M+6TK/nrF55D6v9Yn5I9U6Z+Kd4AIMZpohqtPmVj42gi2uqDCSp7pXEHMgo
WDA3XmiAmBREBUPr+raTP47raRMGPk/RitYlIaPGqU+3/QD1Oj7nvByC0qXTxmyM
l5LloNv1Gylu1AbQZ2z+snlF2UMlw1PhNf3DC7ExDU6qU197FGCilQzSw45Wt7SZ
gjicY7ERik7NsxlRlYpV5QgnNNJ70a6aR9yX2xLiIrdQlDrAnnZcnyroUS0n3LF1
jP53jrCy6ZErNF1b7No7ryepwI1TJJOLJ12KSLFO0+swfq+/n7tBeDWtAHqh18Wj
SZavpZYT4o8FBfr64Uq9PRKnkmCaHev6I2wGz9uQyVLJ1dCZdVuuRKWXzpMJPBHD
w47ZKMrrsi+II3KhOEhh3Ua2B2FuxkrWEje5e2Idwhd2MvsLdYwJNskDliKSc8hB
S26Cnu3PxXHCEKO2vQ1AnppZuCe5nX6AvUIeKdHnskuZnlYdF7nnsm6MUh64PvXQ
mDlaY9teU6sww4Q9UACfR80P3f+GOwt45vCTlBHN0agxgd1ooUO8UVQ6+UDVgJgp
5b580551wjhcnn0eaNhaLN7WyR92vASDeCDWCKzQlQjFWLNldBK+32pwKL4sMyzD
alMJDWZv9jKM4lxUxtGlMWLtuVhv/NdSOqfWpa3DFLWixAFLoAx5BuB58l+S5N/5
+KCMKtKXoVt+26TMSH62MNgc8lKJdAi3VMVDhjI7w+oDouDWY3FipQtodN4M8B9Q
JpoBTpFzV/c1+CA+QD/AWFJg8dzAfORmLqIjZapimMCBQtN652PG3DYIfDcPr3du
9yGp6Ouasi7oGkzefggWlHYAucuzxY+Wp/VkenlfRCkxIJcjqPZLpQ6Zlesmc0Bs
n3PkrKCwJzoIieIb7hjWujOKOqL7IDxeVM9UWdPMYcfOUkSPNlVhhSgL7OJjBvaa
LEoaq/uSsc9BnoDyQCsiDB+OHDdFGBjiA8iKUEgIOiVC+hu/VZ9mN4Kz9+cOw768
ZeFLAHn14sbZCuVdeqrDFnOjS962L9Vzfy25lemmLDGhjgLQcKahQrdO5QUbhj8s
Xtek2F8aLfyycVHh1uzxHNEHc+UdPsvcHTXGvbZ7KDjBhba/x0FbOxv2H8ubjJYv
S7Z5avBHTMJiXvrj+o1DbBKi+71xw0bFoSjZNE0CcInoDJg95KORQFtor2nXu5Wr
+r8cCVrb+Wjp05ZRJsXeS6xL/lUv8ZCaP6R3e8hFLvdH4YSGzrvV0dsiq1j7V7U5
YPthI5Es/v3M9j99kRZrQnDKwpLkVOEg9YKoxj5/yD/plvQKWHsz31lFj70b0EZt
RrOGXBJQhvaSrOWWTNReVjTsN+RyyK5mW1OBGoCw7G8N9kJ0HhM+OzLszC9X22Rr
tsHG0RfCo2NnSOOVxuM7MJ/aLUhyHuCRsJjtAznMIqDl+MG6HQ6+d/9T5tsyhPhy
F9mNIcvh0INvYce+n9T9W1uJCcqHL4RVXhpxDZph5b57w8piLM9EfI8BLfPPkHvs
8fP1wngz0/QDS+tMrMUUzTFWh6WqQN3DF19T8zp3H1fzRv16dR5k6qrWTkUjilLP
fUSECK9p6rrqbRSnipzrgBrU+bMz97CYnTpookk8gFhcvJiCd2qHXbNghrgs5Xtg
krTqnBB6ni2q/1eebtjcsWaFyTa9eKN7w7/0j4EDY/rHfNzssD6+Lh+LMbyrGErA
BiB9dheZO3VZRT+8muLcEd1VecyutX81QRypwA4W6XGrjSkW9mDr0OTw/DS+zO/6
B0Hj2DOm/Eiibv7GGtUlNTDx6MeUi1H9FjzCoZxlJi+l4ZCn+bKrAh1nQpnY7DuE
Q/QoDP+Dqe0ctI5L4yXx/+2Pl1YZ6MMavzwdKVD2FKQYeUf9DlMXfhAeaLaKAkce
lB+smUukw82lI3K5ghoa/CdOKGq37bhYRLXHogLUOSBG4cwq+XuPkySHbgBU6JPR
WZIhsUyqLvLw2pZd9NBO8O7YvBpcPXF/wQSAd+QI949K1ZiqZ0UUM4BP0Y/olZp4
LhcSWCFckyTQkgQxa0a/K9UnJVOVK405gwbuwLw9t0KN4uV9GfWY/3Wqk04NO222
BFPtMVtFICj4L9eoIOUuMw4T/EnA2zw02EFjz4ERfkpzpzoh/FGKfHTA36CGK+bx
za3C0F/NgzBCC/i0FokZn+eo+1iCmFm0xR8KiSj+OADI6qRLV/SY1+3waFfxaDdr
6Pps+G50svzplK7CLjJL6ntST4xfDobqULi4ecijYSskp4b+wq/Rudh5/zGV5Byk
DdeE8ma7CmV1f+j1nrbMqQZgRCkaUYWqA0mdEWbx8vl57m4AnOSwiiJxh0AKluD0
g/yychtMaEwIef+sgL4WuiFvneMoOrzC0qC0Ao2H2UwSKc2QIW5pOJUVChMH02PN
UxxhIFY8U/aIyWn9QchXr/9X7gY5huFFjWw1wIK2r1wDv+pRgfti6G8Rn1uWBYFM
29btneddsk92XIPT9csxpqhtQiXB+3yHxvRQDjFBX7kkF2yN5RsdyCUof/AOUaa3
97d8B9Gz/idq/QPIFPbN5lwl2GnW0KxDXMIels/+ENGCJL1wmrGgO/bQ4ouJGGdK
zlIwyKkS0kz27PFWBGgZc3ZT0QN53rvq7VSRqLb2uLY=
`protect END_PROTECTED
