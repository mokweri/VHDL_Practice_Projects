`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HRs5wOFrK9HQ2+5qOjGZTV27h1CWkdIfu2lkFZb2fclCZMaAfVA8K/c98hfW9tJe
us/WXSsa9MZOONnFMGunxxX5M/lFjpiBszlLiyus4qzYM/olcFKwVZft4+46MAjU
X5kPa5jh/vR7nd+LQnnA4vWjZQxY2XIwEO/bUbgpOf3E8EMOAlqSwrRW6wnYv1Vx
kUxXr7xCDnVlR2JQpJq4P5OqaYFrP3jD+beiTfQsyuXOPDxtgiE7fy6LMlAeVMR5
2lQkJpUuTNf07ulH1OsVU/YhDbOAIa4UVldyugYZWuW7PcAyr6tdQ501l40LNCsH
B9vuZVCUeusSVRyKBCzvFdbmEg/amisjQl/Sj/J3+nby4//utaQG8TDtVF2KsKZn
ha3H4AJoFAlhHIGqeZ3mKM6rPJQZVTUPk30+nVRpb0lwz+nn4qFKXUPZoPe6Ki6x
DWMsaKxYjvJOvd0R4aEXHZtYJGgXaLEDMvAPpQHDRIQy7vs60dA5PdL0cwIBc7vQ
I6agY9lamgn9elC//unPz1ypdc2ykRQTsr8iq8R2sUyiDELqu0Xrd2YQR9a6FeCz
0qPrqude26di+otW8ZGutOibEEkHrv14m6Lx6gGamc2iTmvYl6oriVjis7XPfyQw
TmXujeceX/xrAtJDzv0UCAf1373N5q5thHiumKIaa7d7b8r3to4R2tyfaqsnwKw6
wmW8rhxtCd4edKAO+5mN+Zp5T/YiQ8owX9BOJW0rFBsKHTWXM+pBYEbt+sczWKoJ
`protect END_PROTECTED
