`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0XKwqxTgHRJ2V5bH6c2kprgmTHQafIDHPvSVWkDnemsoW2SUOwpm/cuBZXym+ub
aBxYG7BdnGaxThTEV0Ivq7srU5lUlvJ076UGwpw9b+ArRiBKDRmc8AYp/uJ67LsL
WlO2Wpz2jBuV0eN5+gE7WWOytn3rMnIk//+lkq6fF4YESaLI1hCkhSVBNiIsZf7j
UjhUvTfNiXvSR2UBuvQNwSLU6Sb0HgL0DH81/v3oiAwkIfz6IscS9v8SECcmh8cD
ZWb0242E0oV/VP+59m5diAeud38Y3PqXXrbpm1hg0wz3gJncXoM2IS3x7vBo7mPC
gJC65uAzaiZzXGyCCE+Q/u3AnFwrxUaSIg8tLONpsbjHQnlkKJGvfRlQjc4hOcJT
WxOobDD/MU4K9CJdzIRjMaHHMiWJucWV6y9A/oZ4T/tVlJRYXdfpYMIMooz3NS2G
gz/zie1yxG4vCB49GGx9vMGVkmalch+rRzjE+Wl2xEX83d+9D20ZPEwpOLFIP96n
gkNdK2Qw7NAuWQO/QCLi3GbP9N5XF7ZQrTXfX0Y9070xhii0UhoO+85g1NvOANFn
0OqnBY5k4DYDIaEw8ygp11757smbitpYXHVUcHfxvgE8ILn74vNkRyk5THs4mG0G
ih/tHq6ISpoGc3YV1XRFmLdhgwx1aNAcCDvgT7LZwLlbAt0bP98l3OkfDUuZKYWH
fNmoi6j1Sp0NdfFMwGS485jkuKBv9/R6qGqA8FFcP2T1MbjYK5kv91k4uxfKoAuj
dQnajCzeHecsFoYrrwcgNuFRA07U+lhQfFxHmTS1pov9ciXBHSbbKMFgWExYoXb5
Aep16ulcmmg1kdnv0p4QPdWDJj0lUEHcnjf4kfzuKpCPF79UDNo0ZsYPQdDDtGCE
kD6U0TK9TqdbOvuzCCxFzor0FClg4/9fJT8Sf5aWFmulZz7ZjWvCE+847/I/43ZR
mbH1OtMbEVdEGmGNXkPBRFSvFzTf+EX+lXl06rBbm94FcNh3YRlmNQSMWGdih74V
MCgTqj2LqPJ2Nl+mtbs86fQGan0sHkxZKoDq7LDUeEHDGWJwUZrrRmfCZeb+U23s
V2rpKPHDKBljhwjgYnFtKCxpMwW0ib0IW30JfUDEOJNq0YgNt539cFvtkMlf5T4W
`protect END_PROTECTED
