`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAz+4hXL66mBnS5jD4ZQu5oXIbjFuDUqQmmMz6jerwNP6HQFZJvrOuMwmd1dPPq4
EyFT5LOwfblqhxb5iCIhbwsLjCE1Zt2zsbjkFwVDZgwPkJDhK6xX84mDPS+9FYvZ
DF9YFOW+zcJHeorlNpcNNoQcgnVLFFXAg7LtwuOePIJd26xqaRz4id/zlLvduuT2
Vz1zTgLMjKrsFI4N06JQZenLA4DhAXOewymBMQ15z/25aFLL1Xg5Em/NOApPcTKe
kVBgn/+YUdo8mJLHtIl2jB6EHOeQ9mrz9cZ2aPv9GCX6sKxwrGY90wgiN9enOnPM
kTPcjX+KO0cD3GAOFUp3zb942crtqEGSr8FOAQUQeaMnSHcAYFgLFvsXdUThDB9W
l4Erdp80lplfgDWaBtbLNWOlZLnP8XCLYWhWc8slaIqcPS0I6ham7wc/EWy4ui7y
NTO11stKD0RxMUTjRu3MteJHWs3z4th7p0NnwmbPLCc5DkJSZdRLnY2YifYu/tZL
BxjDSUCxptfDwvGJGvBSi4REgcUfXxDSSjegT9W1TssUDl25YARexKfFwhPlOQYq
pyRvKAlk1IfM1KDNEmZYnEZqmzeCHIU8vCN7GmXIJXWzwqJ8AkPU/Y3q6R65mVAM
4Qb3HGhwGUlLfqAOkikewT9V1LpndAIo+I81kyg6tovgbUqESK8U58ourFqIBwOs
1FBz78bRuMZDS54CssZM+TY9x9kGySZq0zz/sro4Au1iNjwpFfr+cEUKdcgQs+71
4Yqw0/JFVA7I3OqqE+TiwxBBTzwEtub8nl0IVJQe8uue4RTHdh7R2Rn6SJrjMXxY
4kr5xNTc/zsJ6Fuk8SUQnBDJ9AUysy308+87QlOLMoK8rqlP1GHdhvE7smdQIUfc
71REux90RYjvmaNnXjabZ3k32b423s1T+QQNtIwG2hPZSoudFwkFRDBI5CRzgSuX
nNCFkG7xlrde1ZNOYvBqLQ+TnELaFY9zNM5SH2Jox1Fpog6ptl5cliXTsIENqf/T
XwFKzUPnCdFoVe/vVz5Crd2kaWKI0Jgjjk6AXYEgYh22mxZ5wTlXRhQI/QPvL5gm
9aRs0yN9ONqbhm22J8f5o8fBtcWlIvhxUMwf6NCTlv2qjznRJdtE01CrE5hyrZwL
HGU26H0r4K5/kiSIwjaM71nvXsVLTwvU5qvWe2/hk9I+5/qVauxXIt2ccDVr7ZQ2
m2WZSwQIzf+CFr3YShxSsA7GsexBTsUQwjIC5zRLloHfNdLwZQvn+mDyWgLc6StT
PGgF4KGAQVm/BwDHpdODVDgZ0C9hEnN7mEvCYmai4dYvc70hHvgopBS5lySCqo1B
XiYNaVI3rmqmhsWlmDrf+Xvi0A24oUR9BxKv4Ig/uNytyKEWasiZ6su6cPssnpcp
4ZhVKUNFfkHlxLIZJLL4quFdivi9vz2NRhBwJCtdxywylVJyEF8e+cT4rxLJ7Wzj
oZCxSvrXFLzJHQqJtrGlYtDuk9Sv4vNwwsRaOgUS1AFwXee/53QfOOhuNPEet8Nx
BwrrNXegmtJSjvV5ru1uCklA99owW2h/634rorlrjVwsNqL/CgoeE6FFwBtVdng7
i+VA2AOQP1+HTl33c/EeqmhIjTLffmJ3SuJuF/j3+5zicRjWPX/+FFQIDKIqBcah
Xb8F0uwyR+LLgVei3WhQhYIiGbvfffEuQULUBFpNN27cz16abSjYtkMEUiGUKx6c
0z9e2/HG5asNpUiftCuRGltbIPQakpaHDui9YOZl7h0gyx4/gn+BSvYfSrlDrBKa
ch1scV5liS8jI0GxU+hxpcks4aHKRBo7dQCpoZQEQ0bAYhR3OF3L7dnMSzwGUR5a
ACK32t4fbv3KryjnxON2H3JXo21H6sdkxI2wsNLAQds1i2+9+UfKyGdGxfG9pDn7
MqVSAafQtVFPBK4peMfsgcnaH7FdGENQf/tHwsOPiP0rwbHo5unebd1ZD4vCjHXe
OeUXUhgm3m5UFOfmhOdAsUi6SUPTdmvZk+lj6dwWYAa8cOO+PROALXLu+ft4L311
8aAxtek/lBcUrlOxcu92lAdmNCzDdHxSQ47kwhae7tGQR6zj1on2D37/JxKAtPji
UB0xmi93BQJEkhZVo5s97t9K4fKstRiE72Ro6PWuieyt3Z4ED/9C8QwrVhCKSraw
MGYGisln3EDa1g6mHvhx3nHa1l1bQK9aGmV9cVLdS1f/RlI/Qm+858jm7kYTFfn9
3YhNMmF8+TDH0CGhab7AfF6tnOabQ5qRnJRMCJsZfHKeCtv/tRrV2BUyak7JYm96
Qdo5tryBm2XRYEGgvc496HCLB/EmRzGjpyp+AMsk9FA8jvVPftdda6t6WUyZxr/b
2UX/zi4divM94bZgqoQgIA==
`protect END_PROTECTED
