`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hH4rl+KKmhrkeH38GseACotHcwkfYmx52fVLFKf0OAhcTNl2iNhWQCh1LjfdBHk
vfrdP8/n3FD3uq4BRs2BqLm9AwWmO7AQb40X3ltdtEsVc/CzzxJYDBrZa3/55kZC
pt/Uy7gSJFHQ4n2zhNQlmgp82hdQwPe0Z9pLtyht9bOCUHVOjpDfqBhsZSAMOUi+
MYbEZxXHUvhap6wIMi9MLSvSR/t3l+NHrAonGpUmLp+OWH/DCeRQZHVUJ1ZTmKGF
kvBTPxuJuAshklUYukJRbeJ+ho7OJTcwHqAJyoeAYFh8m+eZKgIhARC+bgqEy9tg
gUPfx4AlXhpO4lRc+cLeNquRWSEuQk3R+3iJwYHZ2Sgv8J11ATQUBqJNb032UoJ/
2jcsiAG4N1CASZW2dRhj4dMcGESnUbXkaFk2Czsd2xHSff8gS68EGJvztBniO96K
UgU7lzpFQOZka6wJmY1wWMKnDdYxCVFDYAS9QvnpQ9Wra4NUCOPdz+lGmxnCuCi6
+xUnHURHl6rPO2BtLRiLEQ==
`protect END_PROTECTED
