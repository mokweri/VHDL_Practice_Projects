`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z5KhvOEK4CbKW3Dp7WcBzfljUk3aZxkSPDGmhwG4htxUavLLWcMrd63sWhEE0EKP
ZfY94Uch7hhBXpcQEC96cJDFejc7V5tFJq/RaQ756b9J1peY2bKU2qHvnJjJOSrp
dQ2dkoP4lomJkTqbrwWcYP46WZA41RU/Xjp9oxNtsXsxYEpqORU+iZa9gS5DqRyI
jITgcLFgnjnDjmQa1nV0MkGPjfjQBU/u3sH9nVyAdNviGtcoD/o2DlFAyR9YfirH
ptWdnJH8pkdiFrwLNxrtVxjjdNscZ6dYRNI9QqFRaupDKgiO08dYz7HNy8mkDH+k
R7P6oIWN0i1uU19AYcjrAGvHTiZZVvgkXv8rXkhn+UcCGcNPW6gkdb+jzeDjHQbi
jif+BQcfitdwV+9awZo+1MUWJWS5NUP90el/QoQ1Ydfp2zQJyujcX/41bTW9diI8
DxT4VKHCTfniWzR7o+THIb6F/Bz9AcClzx0YdUO+QoQrqhrufTL8Cysquieohtjh
cseORM2AtrEkwoZHDo8/opRZHtDGicPb4+TTm1lD7YY0SZfG60YL9IJ0FEAzn8st
gDR4zK22f2kFaXBh7MxXDkWnwqDidLshhknc23hVOC1nopNEb4Qd/SGND3U2LmAZ
0KUBPkgPNQjwn6GXc4f1w++Vn1zzo4HCD/+AUvm0GfF5XeXGEepgDOKfhuqRrh4E
tsj5AxwnbKs9qNy3tmo4Ysat6AXEmtMYMFlPjYoutbr6MbNBoLphrY4ige5gpsAj
yiRDkuTU7eHDgzBXLs1XyJAsCmr4+PvubJ1Y7bCbSBkEgjEg/+bCtbB9f1m/EpDl
kAcloDm76YeDYzkYvqN+9xhpOPZgNhR73rl7hy6oqOWIcQUvqdOQIMCj5erpMFt4
HaR6UMeNhqNHo+gO9Rmy/Mv1elEHsCNSffrhbybf952lWqMBFF0ztKRqXMemEYv6
ZGIxj2X8/nHC/hlwXBesw+QAsrBlaSnyof+xNqRChfe/rKpn0seyvisbF6XvGIsk
gLFOkbpt8XuNdLFCOlMmnExcEFLjuhkbbzs6DgKX/o+JlZMYogu5nou69k7Af9/A
1wKp83XiHJSNw4iKN+Vcuvl80jDVSJ6zMvtgnp4hTosEKYozvjuGLUlM6kUQKa4/
WsUko63eTRpX2b2iRLlgfTkKN+NBnmRUpRJOT3B3u5Lx0dOnB5sA8szDg8Y52zo6
Xn7C4zoC0yxlUJtdqaqMZ5cRHC4sDbbRzmyHY94eo8Zm73C9NBJgPgL1v+9meKXs
wIrZWZbRAdnMfyWAzrbNtNSJQTV55XW8ge2WikAxy0jeRsAWP2yDLeJHGxgToL4s
9T77DvjmPPMvlBxW7R5pa4PdgwUv6S35/eQ2J/7hva5ObflIkp0Jct6ZB/UC0Qop
1qV6HKFfWgZd4xtMAmJU011e8u1WXaEmYxfsMT+V9JvAVWWb6J4URbJET1QnVeJP
/FDkythTtanwdyrkFOGagB2qlS+lsEWDRDkmxfrHyEDoJ1FDWMtj9gW/WyWxBfQE
AAI0Z0bZr8yQLXKow4oMyY+2+iD9Wa2YPkQkjBqXPAHF49z4DCD+WRQY0ybS35FN
97w++X4kSLBU7vU0XufpMBZEmKs/qiduX9LfAPosxaucFTTEYHqu7JSJYNHFepwN
BXjM17DAsDgT3UYKu+X8vjd2B7W2MZImmV2j1vEnuMl5N5rX/1w9u96acG52U4/N
fYHv7kURAp1HxGZHhiWA1YkRdIBJ4FYNld6rgfuDrnonEvKTkHCWcQZTMuL67Tf4
bOU9OEfKNyMgnchgStffu7fFkZsf9i1h0LcOmQkU3e+AF5SdnzDFtMavuYfLeRVn
ui6kRG4JvOWnc/V7j8qHIzIUrGlrSiYRcCHO21cKJ/R84hrN3xqKrxVrZyOkf1kx
7OFQIybpt6D6wFxwmDymQkWdfFo99qRvByRcOBYJOybP1tXYEqO0Nd8kzew1yWXA
3htRyMJt3N//+0KcFGcwi3SNmqjf4isUICLQ9DHNW7IVgtLAhwzcLLag9NkpzVzy
xWgBhwEU2dF9IoyMJqvxPafkV2MV5++UanUVZ1hCoirnw2nPMyTT7q1I/+X7ln1Z
xR7P6qaP+SiVKng3K2f39xQq6gSzAm1E/36HsgZX1zvBXYcTfDEBAsGgRhBOLr2u
rIAI+SabwgTr6MR1+dZT1S7bU3cAFlF5T1gA8YsUKVL+r332lkr8L9wPb1u7dVXS
eycnHQHemzbw62/hz4awdwC2XglXuGMp7lm0DcmBwJr8XL/Z+w3lRkfeNL4F5tYW
oCnqKJesKXtO3dCnP1cFuz+yiohYeuDTlE1c6T9hkqRIMn4GDnP/3Blr3c8v7GUo
eLhxs9eqdYXvF6kbWhlPSHoVpTEkJoxlTg8HinwHYZglDEQQzXBgJBH+CNRo/G+2
rN15Bwt0Bn6RfsJN1w1e61gH/3HM3dPnL5mDX+MSA2w9GhuRDWyKnB776M23FdYp
cGRSpK2E+jOEoyQXrLX/MHLXLrggSxJo7JlENCDcT+xdkpVi1O9BF8Yfe0iJOZTO
bO15ldxv2x8acuJsvQMnRGv5/yFVGBpUl0Vkx3kjzmLG2CCmYC82cgCLCZqRGklI
8VwCDtwrclB7j1IxAacUH1TFJ+tpkuN1UP3TjSMdDO6UAXXuItiOhHT1W8vLURuO
mex0PsL9c94gJEsF3NgDTPQjiKp/zAtpWoet5/+NK6/DzfvSO8RtTIxYxIFvB7zg
OYAClLM6Er2oXr9McN35iBfqtalaVgCdZAUtwiPTsMxqpQ6Hi0UyQ/QI7btIT7NG
5RavpmFjKHMhO/JI/ccQus9chu+lsSXCWoyLZoaKfXtjVxIOob8Q3qs0WLB1yAGN
DgwGgUtcbw/8B385hQ2IbYGQge/pVLsahAf/X49yppUUwvHGLAZ+77MTQtmsAK0I
GS0hwSV8xeBZQkxiQ2FiCryKPknYzHnvz4pFFeml8e6gh6fXycoYkN6IZtggESPL
sZvO4CcrWbrwn7gOSfhPfIt4dy4Icirutlq1ax9Hz5JRPtX0wqgZ55/zzfRy8+OL
CydHPvqlWiLGg/sVv3Bsbg2QWCkNUPtnPXm4LJFSAuUVstPwxAZzRbXfw23MGxld
9u2nsFqIbgScZQoVQ3TthSVXcl6l6pZ0Lo9VZ9SIqqd356mT7okjZ7xDf77+PkRe
AWKlpoXnkOzs/LkldBfyaG0FxRuUAMMM1zYP/m0f5lr8I+nWpUvLCWIgyUYk9Dp3
vBM9WxohCLj4hWK6CTXOITPF9fbpqfk8AUCB0jI1zgLxqvKPgzrCGck20ydpq70c
e3Vd3Iqrigv2yrBGIBbJTmduO7f58nH5fX1sjcge9Vote8+wIXoX2zFYCr1rNbOI
I7Xn1cQtcX2jL3htek2hQBMe665V3boMwNv/TBHEpjeFv8rbhcrhoky1pTtBiPjn
qQi460aafy6HS+hOiRmc1GGWG42vV8D86mvbDLAfC9CN2ndyPO8d23UeeHaTvpXd
W4eglJpjTWR/xrkCx2RdsOx4JuPisDGTcBjJkV+XRrcHmBv91pnUeDRr03KbkmK0
aZJ31KNLHkJe8RcWSivRM3IURgPbpk1S4OJJe/VIcjWsqgqVOUm8zoKxAiE4Mo1+
I3KoSowKA7HW1xm5GwhrYKp+KeANGcjZxTPcRhw0cMwrPKZ73IXklIbxIndX8v3a
uOwfhFboM6YsgRMNzadKlG8DIWAGNDCq3HKOHoL0LKaksuO7rrqOfc+zOJwCZ2+e
da7SOIEBWZBHC/UcHRMFt2yymhmFHbQLOvsOmTIPXI6edfpBK6ru80wjzR449b1W
qQT57bES2LfyaFDqDBflMba8qhTY7NncWy94n8Wya04pYg9StI6yEDCtypvOGkIs
9eCrtJWApFQx1C29YbeHOh239v+Ce7qIRdnAfuOreTxlkvJMTqnPiZXoCGXWlRTi
Uscip2/GUyLapmCc0ZOvpZuFvnTwuq5lrIONnwko3EHAM4yY7C1fpdYpKTOd+b4b
4PoE7/FBbAuKMYBlKgVW/Q4MLDHo0s/pM//Oub4uES6m6EcXGfwfuvMPx8yCStGs
EpC8ilBbhjd1qYyEaEEXkFtDbpjhVWffTNRoy4nBWCC55vu6ePsIL9ZbLCaOsCLI
J+6KDxLGnD4p1RMyuV4NlFipeLY3nSTYA7+P5oEmCuVwSNr5zTm+QRgG5oWdAYEi
UCbBgd7ifn8eDx7CCTE5rAcWCTXrX/yQ7RR3RHZ/IoAfvKeGdqHqxyAcFXdRGTKL
bipmdfe6tIWVUescnEu+xeEp77vKOnvcbOWmuQRRtTfdTAobx17aCgptnIL41AKk
6xSK48ko6lzFj28RyBl/5yw6ZhdK43NvI8TPyqhvf2Lp286us6CoEKfSfpH13AmH
Mq+7fTvGoyOMGT+E45vIAl1/M3PcX8Rlw+B3MhWqPHXXpXrzhmak51NyTAKPauE9
s1Wc3PPlLocrsxvrPNBXMmSnXO8jYuPsc0QxneODaaGnSjr6ppYSvO0KVCLSKvKc
fd3guB9tzPwtNPC15idwj5vSRJv5GauKF6cugJ6wK8BBBbPcf/+0cfMeUuhxxPnA
`protect END_PROTECTED
