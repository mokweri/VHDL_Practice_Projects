`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
soOYI4jgWTM0OCa/PXngzbIYOLJFnFXWELloVTdZVhUU3QYzWfNYl5jXX6ozlnkI
DeQjx4szOmwvce579ppL0GAGlGlpbn03QAPdn5nLkLUGJfdZK7O1Docu2asR4vkZ
wmJxFFC9x1gBq5+reriUaNF3hF7zHKlwSomAJDQHOQ3ivrPtF5EyOrIPwMz2MPDi
puwiOUS1PC2X7IQ8WxPrzphDZ9HkdKn1IC2AmXD3EHQ2N4zqJQ+nR7l3eePj+ygS
XqUJWruLQg+b0iFbS1ZxD9tijQ2kpruHyEuba7EZfsX0Kzt7syXl1//Hju3OctfW
gpGFOs2UkYEt8wVi64svIzYg8i0i8d0MhwZgFbfr5EY+NdoxEM3IbITgpu3kph41
L+zVmvdsjVDx2W8qMlP4vQRKB4IhCCYS5FlgCNmps7Abgj9tuj0ZMlNoLCZ71Vgx
/VSQn5sLAxR9nd+yXt9l1RYi2MFUL+OoZeYQvSByIe5B1XWvAlkLvyDW+oFRYCf6
YhdjVDavtQg43UvgU//pFeNA6nBPEkAvzxnJmhpEb68A5YOCtQn00JCH/SaURyJO
ET/Ku+n16ymEkNxH6RxiagzplIKU1SmaL5Kl6+JFlPnAtOZcok1Yhv0V1CHHFvBK
sjDTFS7K4P6aOhE27ViwdvtqfJ1bX2EH4jYOeJOY8PZyhYWqR2v77QZ39R65xPtV
1IDdaZVD9V2EEyBdINbs16KutwTjtMMugLBrJcnxcByyqPXuAfS8FRErLEpNn3oS
`protect END_PROTECTED
