`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqpNaMv7ZVLA8bxvQVk3SpMrck8c15eGeUIDCk9JDhp3BTNLLP7Ph0TMeE+adnk2
KrbL+7kTUh4brrxtTwK0esuP59DKb8QUtsaZTVTf4GoBlFR1GJowk5s8BzDhpgWB
cnyBx5kypC68VMbCiiP3E559XfAztur6XbbToc+xb/ZaGJmmrihhY4NHBtTmVqXn
5HJP58eepoR5bIDBI6MQlVZLQYLzNtNbFVJ0zzfkM2VW0JAgYxvtoUd31cfiqg6X
TQ0RUgBXWRzY+7V7v9M1oIPomLTIC3v0xdt9NrRcM3stpvnWo+K5fLBGFd/c0f4S
1XWfzPGWqsiNdiEOvNXbxYuChmgXmhnxPBcBKI2OCPW+rwDY71+ErmQMQYfd0DUY
CgAGxLhlnwxpZQ3X7gq2reMbNJMWGfEoPaaD9zid36buBcenoz+PcWVE7yJ5I15S
sUlgbArSrl1+5PYYW8bA77QmJAEucwD2QSv6T96KGHG9zotEaWp6fV6dtURkUh3M
HXvNfCeE6HiewR/tBJDgj3ZgblPlnyd+85OQiRiTIsCFPdZamafGaRUMB6y8eJK1
wXc6mczvtu0mUjpG+gg9UgkVmVduJjmfgYy9WhwCO2zxDLY2B6+a/I/niBg8oRgV
gT5XJjVf9ofeJVT/wHem+snyYiEQsw24JDvTJ3BGoVpmhWQPdZemecnPyW6yWRCG
DscpC/tWbZ9lQU/T2rbqRa1iJ+5zxPphnT9KBGXRr1YuP7jpx/re5iigauJvWCUV
u4bQKYij4ztzIHFMUVB9Twiog6rT6qqt+TN68ELQryjKnUmxYdCSFMXxiH3c08Pq
HCV63xPBgthtrbJUPFcdhZbpSYPfPZmALDfl9v/5CduVoJYdb25nylBCDWgAMfPy
5pV62VjJjrGIfhuzaG/epI1wzmkpS4KyfNleBgIECdJNcCCJrz+n66ifA/1mv17V
yNEj/qSCS8NurLoH2+Sm283zoZQNp0BrRrWDqxoOr06zpWI+eeZAmx9KhNb4AOQw
Kepx2C0rbQKwPQliFlYPdlQwXmjQ5IOlegwD0cKV9PPseHteYgdvqTUOyVGjvX1q
pyuIlWiaDkjUcmQuVPR4KT8a9Fn14ezF3b+wPhF1Du6lZEZbl6p6TC5bjWckH8NR
95nV+goGsQq7ATbzoO5J1pgPE0T1h56+vbPujBhiz3X6v1LcxJy6gTdlhV8rA/9K
oZUtfX5ZpJYMWWlyEgmCR/Mkjhk+zpXE0hc4cDWjIWVifAOJsshILceI7hJmIATb
eUnwPrHajfaDPybdfCQD2ZPTmCmWQ856bWFkLe1ZAkQTwmozoCH0Olc1O5T1iGRl
HONxtr3sN3qs5+tAMFbyKkryrS3kNq1OddFZ7LoDgUG2N6z7cmAHzvlAVlQznKDv
tiihle54OmigcCnCRzJr3Vj8vt+uiJz4c8/mq+Lb/zUhJ130RmtHGLb6T4gI6Nbp
17qNr4fk/AHmcDjQ3uVPRhpnM35uxcn8r8fuRiAOcnwIUFFIDzASav0b3GsKU1Xw
navm9ghHqofRj4LrSXAT2oDf/F2Bcs8NUs6OWmVnQCDdzTXlTEHbabPQd2z9ey8u
v9La3RWBF1C3oysbqT85hK28PpN85E2bWfxrJFrRFV81E2XQFF4a7Ip65nLRkLy4
T3CFg3DVJ3jgp6+dw/5fJ32QkmmsgHDfgRFsq2typTdU2SwK+nNchwJLZgRL+YIQ
Qg2c1dlJHitXM+lZQdOhF28zvhm79ymEta9MmCBvaBXNBe3N+wXaw8z/U0U0smEv
`protect END_PROTECTED
