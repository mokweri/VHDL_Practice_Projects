`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65uRGMlQf0B5IFRLO7jr6Vi18p/aPSLagn1li6rithLwMXQZcaC3gFSe8g41MSlY
qVnybjEM1BDWFhQpXmPrmy0+MN6X1TFJdgFlajgnBSSP3Hcq/LR47XSfxRkxn4uK
hzuLjZFhRJD7EDR+9JNbbXM3CUc786scPGe4vDIdOxOO4fzrV6rmhnCF361ulE1/
VLh0lS4yBcIFjPNhbaM5zedgOHgYlIdI+lztWTzIkSyztprxLbpKyBCDQHXt6t5P
eZZCYEyR6oy4ShVvG26D9mzRSjwX/LEAyFS7z6krvMfWiByq2yGwWvNuGJaWod4W
SVSyWnJpL8wUuTNqDY+L7smos4Hs6dwdWnMukcP5l+eMDp/0knZ2dz1EhguvE4o+
4CLT726QI8yesC4ozmBzlb37OMQ9gZMwRC1f7uGF53j8+AU3Z6qBsVWs3jKlRm59
Q7UA48qDam7/p38jKPXSuFddv4827RfQ6kt6zC+gyx8qF8GpKCqIDfuZOVoyY0u3
/A7gfYXfYNh1YsnA9dI2e39hSgWLpSfqgJyMUQo6VNU4Q7r/NkpyFIGAH+whF/yb
oI5JoK/sjgJTb3G5R4Ull3f3Cw7nAfhS9FFxWnPfRu/FAJsUdeppT1+SKFDv8q7z
Sz/YW2K/u+RYmX+8IM8gQ3AYW0ag5uZ7jQax6oiXle0TSe9R0WIEK+26vahvXrsH
`protect END_PROTECTED
