`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XurPZB4pdozT4W817Luew+b5BIFCcW/FNBVVFVYBB7P7ao8MC0R17+2pLQOANtMZ
aiS1tpc5rYEsvJ+Ebh4hLKMKfg5381vfC5/EXfbrQVzSDiIuOM3BDYUDDzLE9HLb
jmAPXdF/c1I7qhLLd/8OKtQ8pQaYovdJmT9T5nxgNMnN9S0DrHQS7WtI4c3rYOiy
ugpWBElIiAhJDFqGphF5jFCrV8oGd9ocYJAiR8Juh7aKtq9M6DK96RCjdCV8dENJ
vI6FCT8mJkJJVQEeLSlyP9ZC9u5k6D0W3gIlATsh5DQg5ZDsLf6QF+VrbeUgcyZ0
ODdfdpBZXFzMp9Ty4yqAIxY0IKdoPW9rt3GhqN/2B2TeTT1n7G46iqx2IBNT9Zed
4TA5E3lwEg4DhOqxEM9TovP62Rmf1AvGJ1DRGVTJATZWX7BdxrRiL7bN+FhMoGuH
G+LMxseOSR4VGNRNNDuYYnn5s3jye8sX04kClyC/p0ttrY8rxtvo6XirJfwdGRdh
1qxv0AJv4XFgdnT+DZgZmHrlsUujXsl+u6ULvhiVB//fmBqcRwWD789ezneVhoe9
ufwbI8HyXYBA2c4LSwKpN3ohbepUjYQcsbrKw4kvUaRSs12e56yU/GCA22PNSLs3
A4WFs/GRYMn2gjjVMtLHSlAAMKAulTrEI1yBZinZxRtuwM1Kui3dQDoduZzBlCrx
rUf7vM89J7W5cjnHVxHashYIIK6fe3mhaEdhRO5AIliBUfRaECEPnv4OzIKgvsaf
vUjxIBygkCVSZNJFGXF7nAWAT2zRDWnTy5YeA8MV6sIcQsNbfIY0HTkPqqQPtNnR
CTl4/jEQZIA9uOxLX2fMhmIgP0UZKGvTb99VS58fOUDKuW8X9YPoySyidXAYrDvL
Iosx6cnXacOcTSL7SiUy6aX34PrBgGLkvqnPMhoPJfI=
`protect END_PROTECTED
