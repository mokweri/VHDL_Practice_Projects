`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YAX7aEiMDOmB+yrn5idQrNwK6iHnpNHMJlRpTmtUmi5OLVv8uNAVy21937hNV94m
MLURNA7WQhNJ6YejAJQViz14ttftdsnu9jogHSZpJnpb2rB3wFvF0o4JCnBWtl5L
lm9JDdzKPRoK2szILFUQtBgNDIuIXXkxYsHg4uQUt0Gi2FNpKfL2/hVBq442Z9bk
r9bGFSha9trXfS0lVyFNjN2qPY1acLRBWRhhsYEWkZb84Ef5FZTsm1NFq+sD+3FA
Wa9LxGK5MUax2DIswbzH9buIUMb+VpEX83n5ddiz7azGswbtkywKHcqaBSSbVaQR
7KUBaB8SJGH3rMPscvh8x5bsrCp1RSb3E14hbZjrOSe7wdgx3e3/MZinHP96sC9W
bhbhID+qNSimruPN5Opeak94rqsB4fLV1so+0jmir1JbjJ1PGrv41E6MShhaS5p5
G32pSz6h4GO8bTld0BtdyRgSvC8J2nKV17JOQL31yvhy/QAdAoWZmMC/YA+5gFQr
Y4xD37458IJVyfFz4X2cknruzofGWuPNN+O7SoE8bK6IDPGaM70gFv/ZSr8AELZv
nFqe65OIkiKPCmu4J0v2GVC08ZWYN4ByeG0oCHexH7wYus5EPsvQoFtR5lVy2jJN
hL3Cm1qjnV0MUVjLzKa8mpRiMm+rMWIt2f4OUJRZS6035aSG3aFB9IebROvnir6Z
VeTGjGVXSOiAeJdOyXRCRYrNNt3H4AOZ37k23DY7mOnhh9tD+tlIc0jSKOu5kbZQ
Qdk1npcBHYH1Z2ZK/CSSoa2ktncd58u7uSOfAPkX2y5LR6Fyt7Iyd3xfBfiEyklO
6FwPn5287A8dXDp5qEDc5Sw1f5v3ZwdQJP0MvoSQwUdW5/YQx1PnhA9gHDuJFH5j
Yz5JXZBIiSGSwuthOwq7E3XECDtrIVhv0w62HicNQwdZL2PfqbuhNGNvRMJSINsr
j5QBMMbHsXAJc6covfQWP5OMisGR42gselb4WRBgnP0RmWeknGfK0g3Tw4Tg6RWG
npOhUUPOxbzXVpRJCjIt4zUqntdU9Z00V259S0F1BDInMcHTHFJcooIH1M9uelt7
GdkMhgom8FQ8Bax6LEmPBswF4oNsrthbqddvA6OAkHa25zVZDk/nFctzaOpLrBsr
F7h8H9WrB7cvx3zHcFB6PdlSOdg26/KmRgyKhZ+7Ac1wwzQkF14lAvnE7tf9+wet
nGh2A7Al09GzWXDFDwSv3lYpjdzzupv4tcztK1eSLK26mP7303ieaeHOCAWXC3SV
j7rAUSyYTnSHqU0TJch1LjxNHsY5f+aV8pS4KOfGOnyvYgzveEimrd8jKGsGkrw3
kD3lkct/hnzmj0BaATS1mmVYf9hhb5rXjm0N13v3eU5sRXaZBEeVOeSQwXcFRg3H
buLtyL2XMeCeLt6mCkeBvX1mBV47PEoBInmjqF1mLK2L06QHV3l8LBe1TIrJ4lU2
RQFVG85xGqGAhLyd1jxsBl/m7HpoUrONG+rxWiJ5GeqlMs2KWckT8WP8+nXNqqbn
BqfjsiW3v3rEjP4FM7jtspgO1fb1MxCt3nGvlhzmrgXjfhMGQx2H+xgRIl3gZ9uW
vQsWWYiHaPLCAN+lCloLGIYhLm0H01nAjj6GxiJXivsS8u9F9hCKQKjKh5qFKZDL
7IlOKYD963dcxRivifmlk9r8nOckBYQplMVUHSIq/Rdm0mWQmxDyUsIeDZH1zuxv
V8O0MntjDflu8it9U/XJ2BlaFrjfDfqRGnMmqhZ9qutCBAOt2pel5gmF6z1fnY0E
7ZyPb00V/HMCLld2FUsmry4qz6AgZcs0w9UcskDXJC/3EzC/naS7N8eA99WkN19/
OVum20l262XXO8MlIzDwDIy7qIqWNZ+XMc+l+8k/640VTwMNUMYbMTzq4aWDOXwr
oJEyPKz9FZDq44QHW8s7f2FWwiw4jUDFoXMmzsWJlQ2GjgXQBmmiXVekzZ9dUYD1
J3Kj3/k0cFFsfXUyuRY5EPHd2ZHwNxQLxJQ+f53k6oqCJZpp3Q+f+XTJlupqt35H
OdFzLVuEMe10ifRi4gla/L/NwMXaEfutqyJN4tH+NDq/6izav02PZQOCitJeVrrb
H7M9v6lrjxJ085MGkWAjlXxX07zfcDoMwXkDQpV2FdKdGr4QV56NaMPb7nczbPpo
dxN4W7KHZo+/7hBW3BOl/vWZHMdtOSlUEuUO604Q7lUTreaVx7rympM7hCCdAlTY
nfg9i8cVhQkqntZwwckYYKQ8WJNuf8QqzYrZ0uOMZr430TrbPliBgngCJ0F764GI
YUyiTq6ZH4HmSNfo9F8njZ9+eFB3AMd6U6+4a31zN7wYd7MzX99aNG7mF4mongVl
cvI5MNpzNuF40Vlt3U+P6oy3ZuvBPzEyaq0sFRXSLFtPW1ABp7vZNNKFDjOHe7dy
WQNWoDa0iqhx2d27URYF5Qe1grHrGdF3fsarccS78v2v4FfbTjT4tmIdrQb76ECq
iyuLxeis1peSKwB0ewP14KbhKyJj0uDf5J84+adektKGautNN2SaXQpxoe9MPknn
4hRxb7d2VcDaOSvF2z6ep2UBf0qwYFgj6tVfFufrWsGJgjF+n4ORC0idliUlhcOP
ijBi6sTrOWVHKT3HBtu2QGJ/UQ1mIHnmbRteyBVaR8FDJvLYcWNx0BVEzncMTxiT
UijVPHNTtO57zlQCvbt0wkTw3qVm0HL8f2ulQz/g3b/a02ok/5SGWZzOJhb5bd0+
01SrQqvkJWwbkfDitCWQa/Z3PQonusIB5RAMa4M3oMFHe0hnZMHeB2TQa0w6V9P5
MFMHGVRlmNIEAjKUzNtT4g3Z78/UhBBMVUmk93GSDHDOoLOVROVplT3hy59c7jdE
vK5Xr0xet3x1CzSfMDw0ZqlJVuqI/lVC4X5LOK8l7nmlDUQWS8Fwca1Fgrd8sZOD
emmrRHB+E9d9C6b6Z+uvxhhWg5yEp2oUxMxo6opEaNlMqIAnotObcDRkAoRqBfmO
vZcNB1T7/az5GPnJj32PyKwe/wt+VhCuWETc/KFhVzJHdk3ymisZk33xHm4iCxVB
KpT6HhBYzTrmTyIQDbdVPA71Z82v6H9OP65F2s0cmuIoipVFnuFmP+hg/oPEEfUS
8Vy8ydJRvwmkhKdhPuqOd5XkNkTw1aztjeVqtt6PrGMhExSfGvs1FDim7df2JjQI
u2XJ0/sRqiowXWq3GvnrwWh1xeEZDk36oAFXk6woa0UU47skqJ4Jgdm7oonEbXMR
H5WMdnIyB2D6S/mPOGDjK3kfqlbBhQ5I23Cbp7DjLNNUViQqT2gCSQzCPpjVeItx
8mAfXLCT1C0d0AsJHeFWVuEG8TEnUfYGrY5SFxjWzi+kE8WduOoJYLJLp7rXyz8U
TT/T9tCLoXb9Iy6UbZAiog04fniEL4WQtVuOf6Z7fkXAsq1D9NZbLd8mh5DEvV7o
COY69uuH/gmenj0Jz1vaWimvsffcG7AP60+pyTtJC91BiOmN9TonbJy2Gu/ygSwr
mYLVKHY3I7JdFEOly0p4HsbHRIVMaHMyJHo4eNrwpgNRHsn/RYr7zDMmNUmft5oi
RU6emZsU6M+ohHSOCuAfXH3/CnGWjebd3yPs3OdL3EaEVczf4a6Ywmk9+C7W2bMT
`protect END_PROTECTED
