`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wyiZjJvfqV6ePcgWb6stsVyxhcKvKAZwUbOjerTbNDRFnNbZyAxLZvhd6oUq1iYH
TG/+k6IdxYeZXf9TwH2ANQ2oxl51qj/eF3cAntjZoxn00V3tAbrU6Wo2u64wSLbI
jEp59/HmYuH+c1kXQUjKs/11j+h38qYPb69D1j92yT3BbbxNM//gh0kgP0nHsDb0
`protect END_PROTECTED
