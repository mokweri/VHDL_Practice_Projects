`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egCnRz6nw9/DgY6/bH9ufInRySdr7agKHx/qSEwx8IR1PfY3mQroat9RXQbN7DIr
O9+dR3eIU1bME/0QOS0xrd6WwHnMhYwBTeEs6uClyQdvOKCyOlrRhQ7jVH6+SuUc
+pbFbJItued77JIw9VK/DX12DEHX0Xmi1T7DyIPirZmzCGPlsNQBt2PLvXwczufP
h5Nfw2n0Bzra6MSu4eEDQh3He9chauEGY8ZiYhZMvwaNzXF+66REO9e9EXtj8DpK
PLPhLSCUL4TRaIb3sd5rtxRg+LVikEXlo6nrD7bOXOUUSVbA0P9nJynAhsGTShmx
FcJk66BFKTT59wIYZgaC8oapfMbSzEny+UzVZEOyo5fWOjLHfmY+UQIIbL/mRJsB
4Cyf7hetQsFKeBf/00PEsQttnSMdaXEXcBjU15AClABcUfJ9tapbgBKLWVk75Z6p
uP8vA+lGkOPNKQzeorb4fM9qRxljt/HenF05dU0UEAcN3RwhaIFsfDRqYWut+A2N
mGWwWKFBInhdNMPXHhP+sG8nLrSzdncvUbcCacZBcrLa1NiGOj4JPouoTXFvW/We
n/XZDdK2cE+LNeLaECzsB0chYF1XVgi8Hm3oKAuyb988P12bGYBpMVRwTsVvxS98
Ecz2MIFc50HINI3N0aIvQ9nA13E3XlJ+huTy93jylrRiVZL89UfL6NzlB9T5w4an
enryozIcBEngPvOITN6qeLDgGvlGf57uDNJelim7R63h6eBYvdkWBR4GEgA+WY2d
R9W7R1MkwWfS+RmNceHpDA5Ns+crhS5HMeDOisPEjSe4axZbVuHnjPGLejYXjNZs
th8MjMRtCLkFLzPlj/37kBZxCM38OMe6GV5iPxTatadsDoz2RYYtVvjUR4rkcaV4
CY65zcLolx/NdPdOrT+6DW9WXQgdcYFmFHHsmNpyqyP9juby6lxAIr6LvZsrZfsA
G+ElZw8HldGcfJePxnKLf9g2tNp6ffDdGdJsotEpQNBsY7RO50uPpDk8wa2l3/ji
VtfIV+4J1E94ywNNmqGWCG+2DLds6iupuWPhRGoFt86AqSb2ekRHBQbfEVrIi3+c
lKsysBHW6UM+ZTe6xZLNU878KcSNoS+gN04Zo+cc6H80bmwcY9xZi/7r1ainwHey
+vEVEtricIaSh3pXFTZ00zy4NldTQ2UUxR1jZOiI2A5RQLtN565L/GNsyBCC0z4m
eZY77a4bQ0hGwLdzgIp+qqnjQ7uhBeUAchy254vjVSo+JfwokhWJkER71JkspRKS
D3BpDGAqz2pFqQ2WGDJUQ5zZ5JPFEshRqRRlTEj9Iumcwmy5/Wnl0iemSQ2xFLAf
/HRJqpYxc4dzQWfrg956DckJEKb4cNQdzTzpj4dHJmZen5qRVYqPCK5YFk5zaqQJ
Gay29fw6vwIu9snrtYfoa7k/0h6e3nTRT7y3pumEzB0MFsLCPCDvfBG2ogScIDpH
6zYbmWSrYLlWfrvYOdZ2fV86SlMYNhEtFmMbtxFusHpt5CWd1gAes7N/BBGjfyWM
N7+IFgkSivEEPwH5RAkWof44uekH22WN+d0g6ASfAPeH9d7m4Px9qM+WsUs1NJrL
1LY1/UFqQ8ioao7WeRSCi5/K7qEkTynyZgwKq1sQzGBrFjyRfEKmn6H7esWU8fsA
2eZI4YUM0226/UZPpuQcpRIdKnjJe2+1su8uxQDpVqq5kM5oBK83ZWuUqb7wniII
0dWswMyT6pX1TryEaZhaX3Mew9RDCr7OkpJXwgBP5petlfulEZEGvpCeis4qnBJ9
sfrXQHIWK9yPBzspJ5PxJYa02Y92AKr1GvBCBLJQT6ZHRTlT+vm2VCQmxNAzG+RD
Qwowj9lHAwwXKlFZB6/hgpLEZqTtzxaCE5Xf7Vg1vy3In508BeBLrUKEyqjFWQD3
YfeaZMT9dsz8GqewqLR8dXERdP6/30/OWlAtbQKiSWk3irzfkkhJt5SoU1wchbVP
R7gUn0fbuGrm3PR81pt7TXAjWIjNG60BADrGPp9Il+t+lOfFZlNRfcmFPog662QQ
`protect END_PROTECTED
