`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kxPdDo/CJLBPRpxpiIwkni4qkFHEg/LXvfIO/nCFQ/zrl5Kg3ui8rIe+PeJNHZL
MPLwMQfME3VD48i7VTPmxADiUvKIbfgqW8k3ywQyIUETdIyVLVobdq31SZDzMf45
4NrJju4mVXYIiLg4tB6aAuMjMwabYYQGPw6JfrF3SQ82addBtgMtyrDCBqHcAmZj
ionC2tj2evwD8SuJMBiES27yDuD0A/Bf7lYGkJ23ZQPr0GFnT8eH+ODNhcpL+6sS
4W0K1ybs6khi1UMR7U1JPQ/UMsnUOCwBF3fJ9wUOmUloFjWqYSe1I0JiaNT8TzbE
EjdMGshFKgWyR06ViiNvR8uiX2eDRZ+MKNFj6qZiQ8ttCQsZlZ/lN0qAXFcSRoe0
Z8D2e9Go1y24TN16ePiWG8NIavLI1g1qMwTz4JBGcHRV+Og5bAYoMw6PrQZQtYmR
C4X6zifcapjna7iYQDqRYkOV5Uw6A6q1B8JBInPsh7WDUFdlrlb98+1+1RhqY5ZM
v01wXyqvL+iBme5yABx5eurju5xB4kOEGpLYJ8w3kYB7KOKpDEUIxdwe2gRScZiG
jOya89yVh166G5n8OX7tJzRi2vqm4k/L5AOi9rzXqRBoqC1WtsYU7x6EVHT1FLrX
Pj1Wqmk4BpmzGK30Rbs0FqTGDrgtixPv0UVb5dN2xpKuJCkQjvjXDAa+YbBNSlE8
Lv143ld0Yt2fyeVqulxyQk4UQWzFmemHWM2M3Wn7UU4JC0nbBl8M5mJcSH8y0CHr
wc5d0Gr/ANLRP7qJRI0wjY74IOq7h+r+mjYgIxwgJWW40k5R0X2WiHCe/qtNMX0T
n3D8tlYUj69jzx39azRXB4sWOSqkA/QjDDN7bflEpo3BG2W/MCfr26O0UN+xAuhr
ZuwOQopNKvQbe8En3HVv7NEKGemEWtkuHoBpY2UDXGsIvA5FqfIvrc3afflyMfLx
HqZnBx7+ZPuER3SWyeIFfVkfXwcUbrO//wU3Z+FHMe4qMJu9eXpn4Ck+V/40lac3
DvvTMUIBNZDFw53WAnabFlOkAfgQvsmXCFnM4c5GQ4ZPNJw9wxSRDx/3iw4rNywp
JcaU741ins9XppDEaeSm5hTnazZr8sqZDCdLxiId+SJFMa3xdDjpQRz4AeOPvJnF
Jrs8XGqOfi9ncnA0QlSXMulaEdEQXDLtrGX4MkgziWZLTqIlfhu8lt+w3z8Fb43E
Ip2a4HqoC08W/k7Jpx38mFi/RTSYSMK2yVwVsAO/OKe3BKmjnmToLSzIg8Gvfbfj
fWXrRoOEz+llkMi11LnjMze0xOB8deKk7RVfxR5gm+lNXBxRygn/77L7C1iD5a9R
+PeqsJY/OldgedxeD/aB9YKHKlG1YpWum8vg1ORXpjRZVGxHtWWeD3tD5W742qrY
Ra27yREQurYqiha16UA6k/t+VzURz4pHqjI/bBNKaZfOZRDcQDuKxg4x+1OCdq6T
9b1qhtkuy0Fkc4VgYKOfeVhVESz0ayAoHMKG6BjehEk=
`protect END_PROTECTED
