`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
io6f5Cg75uYLbtZ521ZqO25MzqJXyNYUyprs5dVAKC9Q30kQqd+w4+lUwdvr1znk
USInIVPnN397ktqkzGAD38lkEWl3gwKMPcYprtawlsf/f1yH6V+b07YfCRd4DQWS
NNOcyS0ZNEgm2VLqqEFmQrdP81vStpxM5whdYTjI9zWQxaFG8QsEPVVFHmRaDacy
CUHUdrCuZTl1aFeyGwFmthBm5/wq3uj/VPwI7WKNL5G4HjS0Hq3KZmxtUd0JBIPW
lNdbGVN3yXGTI6xvyH6sLHKi9hHIkZoZUi7G+1EoXoeUnJZMeCnaaOibXmkOzNLe
fgFze7cZDwuFV+9TpBs7oZ4kQ85OzqrmmbF6j5pg5VEoeaubqnWnm59h4PRvoFNM
dEY0Vz92D4xaxEZ+Q0UlbBD0PlqRE6enCv1Vsavg/BUJRbHTtIneyw3/MC7lxORW
8BA/AOkt3I5i1AWPy/eonb3hvpPlFwg2S0CTLtLPTRm9PsW8/z14BcW0ICO1YwLR
W18d0kL8H3n2mnC9ISERXd+82VVA3km4+nNIdBC5iOFxKNOfGYigcitWpUcduX8j
FTNbjUpyv/fXBiJx2QQd9AKAhFcwY9uDfKGU3y4JqHcZ+FWJ1M7gBb9+C9VEBsrW
l7NA5tlsy4XrScWLcbztGc3zbmr9k+7IlYNUGLcixeUswIGtTZ9sXbslE0GkQkeB
F0yObaZKKAsuJ/2TNDhSUyrmLiKK0MmkXHLPqW8HNTBNXgrQybXo3gsKVNJN7TQa
MSLHDG0XXagIGZfe/jCE+5oa+m9OzMhnPCllvEVaM5XC2396qZIWvSKkuoG3GcpH
FK8g+8jUYbro/XL53XsHjN5461Inrg6LUOUBfma2+/M/J1DrkrJByAyfYtdDYEVw
mu7Ysw4xFV6pQ5U07r3QiVSzf1m6g/fpLU0hUjH4oukcyFgDVWK022bnhyej9/4U
n59m78YGooqsizm2SbHGonbY8m6/514Njy8NOo10RM/efmK4UyJI7M4KvpAHuZNt
WzngXomV4Qr/H+ACGfSdzZ6ZXz/DDxjTfR91hbjOgHLLtDM1pJ8sp2H2bJC9RydR
Jx7QHsorS0NlEj00htAc61x9oW4l8t8MlVTIIC6/GzboC6hfdW/8jB4mhgI4BT1W
7xw9sYyEbN3ZhitrL+VwAkfv+h1a3zeO3AMZ1ZPCamEQoyV4Ke22GqdDSq27BmQu
iYItenzsoPw2LyrLxkzkL0NJsacugvW1pAbVt29SkCWkDO29mntdDquI2JEWYPcQ
gN2outwaoikZfs/4ArCWzVkqec1/NzMczunY4A7yZZA5sopRWTf1IKphzzolTiA3
iQE4HoV7mOFgVm41w7doMzyFZNDdPAd+OrSUGwvekSyO93oX9tzBbAz9xU+UM5GP
KAuVPDIIm0fDRluF7lyHcoaXovmHl8kJjcCsKuHf0JcdDYdFR57pK+DnQ3rZRRkf
dnj/mAWKRrfJpSoEKn8JhfHf9/3keRaNxInkfrNjPLbb7t/tqYm2ihyYmeY2/FQt
vVMOrqYTIn0YmoUKy7xw6uZBEhtY5jmWkk2StrSBLyllXCTcMIEFlsPZtO7q8CVW
NPdfDX+M6T0bTGEjpJDBiZhqnN7X92dKnrB27u73FueIQpCZk/eQ7KySaKhgVF08
vfiQ3UieD/YQnBiCloAjAFBtddRMf0ZfUSpPaeJQf8VxJURDUxyN9LrJa/alPKGw
tV0cVJM80rgvHGjaOoL4bD4wtoldmucyw3cKbyy76NDtakFvwWWM9L28/KIqfns1
28FKyktASRNHOyEP0PwHszkn4eCyJ6H2x8lrhdGmEzMYkIpl6JXHIed+YpAbvEzk
W9fL7lelFW7S1FQsbPUU+z0L5wAl7BiqDEVt9LY/LA9ZTf5OQDLbwWuxLjmIgNlJ
fmI/F70np42g64Dl87Zs+VeeNdfTdyFPUeiFvbi2LpIE8SbOZq5O1P7AAKhWNXxo
Ayl3WNYXw8ur6EtezloBJVJThGHg2MHF42pW42E9h7c0Tpf+eUZrUEZje87gu9qW
AEhELkLQsGT/3DttjQoga1UtuJRxEKvejcKc6j0dUFKUs585BXUAd8tve/6RpqE4
t5eQbw+FzyUYbFq6/N9Or5ooUxdUBFeH/ynpCqAZFN1gFLelRU0KPFIIo8h0oI4L
HhthuJ3RYZ4C1sonLy8XZPU6e8oZyq4OOTIR0vbcrqUqUrtknrmz0YEaNdSHFd56
OlBp2lzcmjdxc2yC4EUDvCokFBrlYWToaZGZLdsxWW4Dhcwf5q90rZ53RTpEJyRJ
4dv3QYwNYkh5Rwp1fPL/906zBXN+AM2RXfCZbAGBNDU02xVIJDu9xn9ww4SL3RFx
sMlojt/6VuxIL25aVgSPb0dLCJ6oCBsz6oyac8N2yELDeUhHT01U0aKwveWoRtVR
szxHfXE+4ugRO7mVIG0L1gzlXmVosWiFNlbql2199LQr4OKEpcw+YoJMg+GxrDZA
hEYLjbPVidYRdURkQCtjLBpdgMqUJTCGW8//IfLJ33xfnIc08xiLazyxAfZVj3rj
oWvizSSd4TYUO0RA2m2dOeYR4qB1iakJJd4O5bbzKaXgy/ZhFCvD8F40aa9C8n05
A1SlynW1uWN+J49tE2X01DWC30zXVxK817dV01oYFtPYp4yCDOFz8l77DjJPg8hN
qkNRMpPpGe1UDX2nreuCS++vpvSeBaxHAksoxqjpEOLoVkIGZWMN9emuFEkv4tps
fnkXQ2oFXzyga51xDbQv2mVIs74o2JB8X5HQxLqEvnWCeBnvHAl25x32c222YVkN
t2PeXT+YMKzONl3ZXPXwzwEEbndJcvdyoqD4g4SnkomrPlhEAodDlm4z1ieslWOK
BIbPtqR1nx1ZpIy4vrpnYG+yKVN+KBB5YdVTr4/YPRLt03yCA7yBPl7ABTIF4CVE
ZCm1N8Cc+huwPgVFCyJXmBJ3des7cNn8KwOHioWltP6Bsg8AhRFOKmEatEHfAUkP
kb8IaDgAI0CkXH0Pwk4XnGjAbTrAJ2a9Ftp/O6pqJegEVzBHNLF08lpaI148QYT3
cV4lP7Y7QPajMxW7fay8o8PZEgYKXQ92+IDA6MKutn7P69RyV+nl34uPd5XezLa7
T4KjgdHbKasK2cIKaqOOF7DYGLN0rvJugCpbU6C4dydXxozF38CBIfb/8ILNKb8Z
BMhi64ToHSOX19YFq3zT5kxSZcNucx7H+XA8X1tVBEzY5SCvviiyvq5VDO8ohRr0
nQ505/llP7BKtJFkpp2yQ120tcGfT96eGUGPEZceyN+kVBmjidpqmllPyDTju1QF
tSETtatCDbkDw4YuVbCudPd7fPDSzFDcCg8juPdeMrGk5320BT4WhMcaVw8nQpbF
lbmCGT67ek4uPQoXeiR5FpoQ3tsINtyJABjwI65P6vGYA//4AZbA0lNBSW6pRyRC
DVOD3W2EsJRu9LaT40DjeNGcvkFSkMh+X0aUL3pZv6h4Nl07DpdhAHvU9E3/Y4YL
PX3d2dygGrhPEQEWq4vRPZ5hzm8TWIbKd49TRHopNDZCeVsnQUkq8oG+798G3LwJ
tU/yF0naLgYr8M3NS/AKCmKE3nTdAxX1rUibjau8n4XE8/VXQ3nz4JzYszW+s+HO
ReqDn4QgyAo1xUTTRh2nAxKWspfeuu6+bpefGvlcqvke7IHnDHUYx+fTesVGRs2U
bBAmU1Tuk7TyQJhCdjgHRlrQUxxuoTV6OopmRB+gW6SditU237huP+6mAZEW2+oh
J7s0hF9zJa7xNQnumLbfSPHHQPLUw9oD9o5f6S/wi1KR/YDtNdHcB+hKwglV7w7v
gIgA//pHzs8pv24gSUva0cKHRko7EuTVbfiUfE3ZAm5Bwg+oXFFETy7slB4h1cj9
aXOF4JLcEGtlOERcp1B9g8iRrsWFeS6RUv+60bbkJ0qsvYaNCAdYMRalh6loaV4P
`protect END_PROTECTED
