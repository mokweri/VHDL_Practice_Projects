`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mz5s6HchbSRISj2tTWTbyb9cX/Q4nQ7b5+qdCSk2Yvyn+OKgsR4s+U9NhJk5gPHH
5qSOBeE1Vf6Dqr4KP2+VRt0G01XfNV91Fmok9l5uglOQs6m8cqLmHC4swcvMyKk4
i+eCeZRLNB95nJ+tE8vuwD1LvPXiswKU0aQUeWWYgds6TWosi0RTym63Zi5T7/ie
2/mX4pupTZqquwgFziJHDGRMKXPlj8M08IGBh8nDkjO3xFtJH8/tXfmpb86E3fGw
04unOSH3U6X3WF7jaH0ZvRUGaNpesqTobIe1FTolIPOCkOAO+1NQoHIOoUnbu8Rh
T4dzU+B5JKaRawtVk0I+g8LwWJqdCd5LlnpG+2nDn7xRb43EvxW7KlAtsCPhAwpP
YF0oxxGMiykcyFdQ/26oEJWivw8qh7lkeYPwJ9sgmpL5cbmyNIU9GqPPv+SsvBdh
pnV6aokAQG0Z0JxRYPFxdOe8LT8PgswoXOf3QDUdvJQd0p4IRT5IGhytMOu8NQ2F
aRv2rH7Kme1L5VVjdWYXVFrZ2ixbrC0Q5RxP7ECofqw7q5l5y7PKCVXTReR6eVnB
ANL1zJ4BibMgAZnvHZ5O7LtK5pPlupDFp9/99t2v07SIpRliSmgzNFLFQWSh1Wsu
yaucb2yaq0Lt+1IP5tQ/MV0vOLFHHcxGVJHBTLElXWbDnVOSdwwY6bBUM+s6qNk4
ccznK0qd4BufHH7boGOT6U6y7hU6STw0bUviQ0uczAOYmiEeoRP3VT2RWiqNHujF
zE9DOkcftVTEM3QZhAgDOI6eAarxB7nBZgD7fwanwwjzg3FlfH2NQLZzchNGNDwo
s2uSD4yHwkfobzQONixh1FHLDANk5JECCIfHQ3G8rX7DR2oZ0Jd+H6JsOvh7zSkA
n+XTrqGuqs/jayYvR/Gw2jY5p/qLdq+nzgonDIa4zvwqmTkSUdf5cTvVthaP3faA
UaKflYH3bRNNOq/Khht8LsHQ7ShFMn6KqnDmbbhmsm/JLYn2ld5upxPiI+XlTycU
UNxerGVBMmm3EeWm5Kdqqd6/gGhTmnsd/qSxRASaIq4AtN5MUXYj9DrUzMCtWLxb
o1FNG6/LGq+htJJEhqnLTzftA3Ed6LJEhMBiSxJNrFit6UDs4SnIccRr3BAzIIW3
yYSNeldZK71KieV23iZdnb8AChKgKDMC8J9VV7SvaTeA0XRgXzBgshlmo7hOInDf
qVb7idzA0vphkfxRf1BP16fKpw7mg5QaStcRu312u1zhcyDDeuP2/mM+YZ3TZYce
YjSBWjk6XwmSGfp6FP1zPU1zKivjjpxjsvjkfWRIyxjwJWqZGkWrOesfMHPLga0k
xERhFmzI6iQojzcuXGHjvpIbBGoineEQ3mfqjWgyOfaJrozl7xMQW7M7YR3SBeDg
6riuz1L2W0s2Sc6QKHlkcKAF5LC3CSvSNND5yY35x1tUNQwS4sd6lqIQ8RAgsEA8
ARLXfRi3upKkoow8x6+LtMYv4yVL6K+rlP7uxKpntBOIG+CFz9dlNpDU/DIdvUdq
mvyJB8503hHJrBlTEXb7H6fm0tD2g0Kecq/bTBfBKjSUjtMskHJnVQKktu0CfPf+
Wm6aJBPHX1dzZf5eIIZ3yRImvJyiftqRJgwRgklUWgUFISZglr3GY6H4tOZesghk
c21OsjCPzTwCe45YlyyfYux26HO1Z8C5INjv8Jd+KOsCT1ROFshU6fmQpYIiWASf
HVV2QPID2rrS5RrN4U28yHWHm/HdplEVo6BMAAeUsl/BExfJd9i5anXV99DTZpuJ
Ay9OLGexEpoYPiCBFDpAdJ8C9R3p7dIwiMOw98mhT2K6dg54kqN+f+PIZHyGiO7e
DxoAbzs083Gsnbdcq3j6nDrQkd5vQuYv7NkehgAE3loi9avA9Vgz5FGpSvMTKdRa
I6sJdJ3llD27r2VZaKrRmtK9ixkTCoRXov8M3LDVts31xfukAxNxEmcIJOv1DxVt
6qmLD5Ue5oPTGUEXlnstqD1/vi5sRAbe19v0j6cqPZFn3qi+V0C+ObdkpQy7zTxx
Q+jyBrtz8l13Zr4r7HFiHANZq+yuXeZqXmNwszIV6h6PluSO4UNvWIztGwZRCLvR
55oxeUdw9JgsZRElbe3GvLDBrUU4ig7Yz6r9A8uSQRHrNdMJj5RdE10ILHfbpa+p
sqQV/bZ+ajIQ66rSR0kGgJ75dtXS4MjOGDhV/aQqUg+/tUXmVATadyJuES0JD/A3
jIUXucn4JCaxb7h/1yMmALYlMButHhlOdn+hTN+RnwhL8eD3w1IOg2RTlCETQQ28
Dazvsp/1pD4Pwia560t1Zhta2KPMniJabi7WJqC4Yf9BFEoeDJhOZO+k27YQCRUT
pnWfzteS0P37fKSGm4UCgIYTgO6r7B8P9MARQdcfe6Vow1zi+eS2XBPNASKJOQSZ
IjNkncBWvmV+RPo/2Zsg5wTnF0Swpio1hlYmly3+z9ZUsjmF1ZexDVsPOTRduCTC
E2yV3OMAt2xiA+EHFiC45tPS8oGlJKDUrZsKP9SOtOtm/cLvhSywme3Fg+756S8X
zbPKfHspNfKCnPAP/87jLill5d7OatNeaHNAF4kNc2dDeRrEUwndQV7N1LITnvSG
rBGDhtOFfL+2TqRWHHsJRO8P82J9js191o2gbCjEXLMHAqBXRBGCTIjy50QKoSeq
+Q7Madk7S+NZ5b2cTozrhXaE+B9iaoaZOq5l8i0Bj3b31E1/Bek4Jpa/ff4/cd/w
rzSYSc4SJYcGpzihsW7/1Wysdhoc+8zBQPyq+3c68iwlt3XiLhK01MwHGLx0Zb9C
oAdFnqlks2eD1polnoy4ov/kjdjIYa0RmF+7ELHFVG0MT7Fe4fs3/nQKpSxaWA99
UmvKrXwejrjRSCcDfsT5nn+BcsAMIVffMMbHZ1oXEbtJyeX6WMVLnl2J6nNLaXP0
nGplyqFZzobCEXyba7S6eJ6WSJFXVnXMo6zCkNBj/85mydIb/g/l7qlgWcqIOhDF
J3Z3oVQ8aDyWvtfZunxkfEStA5zT3r3z3edBXvH5a2IehQ2qcsjN2Z9Lp47hBaSp
IsLBhsfFHkbaflJlamBEMBoizGMCP/w0ovmBBAzslmVAmGRVdaH/zbdx6d6RfPtX
ZvQtS3Y4uElza7y14S0WRIQdFUEWHWE3S+2reqR2P/ldtNsfQmX5ZniRH4SDEkO1
6X2LflBOHhfltvgJjGmNoZUbXcJol3gllKrioNnmKSSrWo7ikxrmaMly5r0ve3TN
Xc8i/hxqMQ3IBGvDUFKxQAFemCT+ZqB6Op3yYDlwPhlJ9ifQenFJ3HlcTfFbyoyT
IsRiexo2RIUptYT0fvMrtUUhk5jcMwx1gy52dZeRrbesVdQNsNYIX205VYjsNEqw
dhTxlngXzNLKwMQDPaI1mznihI3jqXuWS3tvqEPZ6z3lLOGPfy17xf+AbvYtBnJm
DGy2WAsB21DUVpJ01hMhFhWmj2y+9vRk3pia/9rw1+abVYHxZVal3AQrD7Cw+8P5
iBncvO8K/p3iBHLIG0MVPT+zHofpoZV9b+QFYYzHDUDIG/6RUvMkW4XNb7j/Xcus
UBcyglCKBiZHIX4/MY0hHIW9m6Irxj7y2bRv3V9Ox01V8+/dIolIg5cwX8BsbRsd
0YKhWk4ukx3tCYKWRm1B25y9YN3EZtShulv1IgllXrrznAlPFOl9kNPOMQw48HnT
fsg2xqrL/1D9egizR7jw7f3p2maX4ONigmsL1iTTeec9juwwOoKz2NzsUmMSKqvP
CWwQs9tOBcoqqp3HLB2pbbszziVzYu3tHt3Nr+m0oxYxT+TCcXpY8OIAYpqkS39q
mr6MbJlZaLjJq2ex5TkjpkQpl9UIOZlxqpO4k2lQUvNbJRCNHRpmVtMcG6vQjbp1
7Ctwojg+BA0ACA1+9wsUt6ilX/17kRj2oT47cJjN8w0V9kbRD9feo4d0S09t3+Yx
rXy2q5JIxG24VHryaKgzriRTHMU/Q0ZmfnJFjzqyZvPgxbeiA8wpMQa6dOFEDwn0
v8w8zS6ukMgKUCid081SQVA1dZCqFlb4lt/iuKHM58gscCz3rjcq2W/jlZq801YN
4woL9eH6h93auI7oW/dc/ZNpjEUpLM/EvQFm+falw+7ddRQy/BPs7qG7lNC/9MHD
9ilV0xwEIGxWAbu5gBuXVzpukfMk/TmqBVv1D3qmJbVKLdjH3xRLQu8EGj985h/x
FuBBudLMP3LZA1OdDdx22swY9NypUVEU/rbkOUspVk7P/7s4Y+VITCl3vl9CnLkg
LOOjF2v1J1Ez7P9JaEcAPgWkx1BfCoZOXlcg+6IYpJrgGq5mWkltJO+8hxyDTtmc
XV+W+54249iZL10a3zk85EUZEhSO/XYj+GmCulTT42r8y2g6nGuWFx2Ky2sNnn43
zzjMDN3M3uIT0BUAMyN0mKmYl1VLs0TKIA3B+GIRZGNx/ZOBt2MrhBQDkfHTGr9k
Epg1tG09CT4HZ/cHNGKenI8AU2kc7BSXOZhVU5KSedPNcbt2NkKFJHZBQuFkliIH
yYKburdh3t3NQC9dQAgOp3isKKiuHLAiNVWVvF+YBMOVffWHz7LgXhriHoLact22
o9mebyZLnTzpQWPnInKcXKd9e2IUOKcYao+EWHcTekbn9y9A4tsKwBDF5CpN9kZw
03NTxPSdpOekrogYURiqSwCjrsd21DDbJsVimDZCOEOQ58Xp6GomhuEIqmKSkWvw
na9grZdjWz/C9zb4FivZie3nnAH4xo7/HiCp2vauOffqemcEW12O8xEu6RKQ3Kh3
oed/8cpvIWv+vgE6upayu1ApBZtvRft2cAzLhDyoY461cSm6Rsz2IHpSVVpJ0Ixj
bXNcrjpHSy5ixuHvkgEti4OOckZEa1V/rUVffpmAXIkTNylWxfaoMn3VPJq6A7SX
YMK5fVM9A0q2fs8Nc4JEGIueA0aiFsyPAiE39kRmk4E=
`protect END_PROTECTED
