`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CO2jFerwjZK6HpxU0aPuGPArOpHTa5jQfhI+g2CuiaA2fGGPK4z4LCr5igkOkb6v
/mi770CmcJAFDDj2VJJf9XaOF5rY92ISHTasiKv8wZajRRybtkfC4tf77NwV0pNa
cq8UElunYhgDtOyn0KiWcAZtDbEiO+TFtDVIkRZVn0ZDSw+vJBUw6o0Biz89hBjl
TXc9fPMw/YBdpHMZpBf7wHBnrIFGeK+qOVh/gSLVIaALEOTUUk/FAhENO6WTUowF
Os7bPY4O9G5DKDW2Dp6VeAn5nA/NnfsX3p6vFvrJ4IAuI3LdsBb+9R+WfJsG9I/G
/8hi7nW62KNGVd62Aam75pG50K5ldYhTsEUDgqHMV7DllkWWMdxa1A6HNzKmea8k
zEY+qV16J5yxV7Y6pC1gNcbcE2aUjEqv0jenFyAcQt3tECPPHqwtj1AjsHWWFnOF
gGcSrjuRRhQfFUFdTSjvwYW5j+Lx/uMvQu/m56DZSgVvbmnE7/AX1huKyyJvP3iS
SHWJ3CL9xGL9pTTfA6UQ0Ahu0J2G3jeaMSP1cUWBBz82UlzlV+0nKOMNS1uRiQyO
87dXlS0ZqvTAdcsQHkVcaAoXBY1u0Woql0Z2TbcqkmpneJkN1RHHdGlep1xvX7FV
BQf3du/GxeU11sg4sv4DtueLD/lwd0EK3GHPhtXnraZiyI4vqzPRUT2YxRRz1ofd
QSdaci3aS7pc29xJZ4LOI5/O8zSF1+dF1wfWdgtSq7gK37i9Q6yvAS9HnxCXYBkv
WNrBq+RCFIoUSlibbO6CPrg2NJZvSgjwhX3SfQsa4Ns2shl28Zi4jT/rJUB3gG8Z
DsWRubmK1ej7UWTgOVZynDcm2Gus9gdKTbq5vobkzMZ83FG3oSObCqz+PQKh3ez6
65IlEGPvqC49Z2ks+wIJB2qO0NIE/S4KUT0scPPM7181Z+4+jCnx16ieTL+NvHcw
+zK3HAr3RsUnaaAqbRvqP8ZgqRSTndW9nKKNnao9QLesnTK2IvdGzf7W5fIUsC5V
B6F+RRwUaqUoSCqiknDeDg/8Ixg9QTQa/rLROkZ0j+frSBLeiDslCrTk1R20Kdoy
4VpsGISOsGwGI+jQ3/OfcjIxiXKtDiS+nWBoe1JQ+LY3ogzukpEf97frsMZHnFiE
RUt25TjLBGBuNIwUrFJ5w2X55SzlugxP3xVYAFDDQJ55fnx9Mdbs87r86TJwffjr
46STAM950Kugj1TNfdf04yNiWQ/Pr4Z9+/3S46DulhgO4ss/gECatlHm8/BZY0GU
Kng3A49T1GSvhLdiomnI7dRsmL5ck4Vfnf7dwdDxX+7Gt8Gj4olExIIJ8x5tSxyj
9FKcchDVwDRV5dp5pX7U4YDIFyLd+aTPM5Gb65Hkx6zEvCJ2jJMo0IYpJHorDHxV
6iPUB7ZoE0u4em0PccXBElozEVtCtJCrrSuhlnRVTD3qr0OSk+51ZSbSApJefevV
3TL2mixQ9b2FcIL24UZ3yGNkkN3fPs0Y48c2w8+9byCWoEdclRFWX7Meo95i2BGo
TciNtkYYJOjIEfHNBYAldei9Fn3AXEyv8aC7mrkN1VQvkHOIaF8ia/um15hNzPMU
Fh6uWp6tckiCPtjZUGdyQfrsQ4YxhVk2z+jPD5Dg4uGU43pAPNEmlwk9CWEob1uI
+q0vV9BOT1pTv1zz7ZLwscCYaPvqc2MebSF+950WYjtDtJ1kHyeEha06e6j/yl+b
69xuyVKuF6zS6S8oIN1wLlw+F8EdsqMLJLKdDv8CFZ0yiQKqNo+tna2RKQHEviip
YSr8XWjGPL62GMw/zeOmt286eX1+bOxK5RFqoUblIiaumjqx5j4IsQFE7cz6fswX
LTjvbegIARJvnK8G4w0V9S4+2j9xrchqILnFFw1MF61cxe0SJ2nQAmsFAQhxi4y7
hq2Iv1aV3ia38XK88eayaeqKtkP4HnLx4zXgII9MB9t9DrZ9HF9br6j9HHG4NzZq
zYAKkjgM6TzPd6NMAYHTKtVebZaeWtqnG78tj1liAP023C3FavrAHXisnSNQIsgi
NZW0adEiVbEUhsd/fREf4Zh02nBvgyjSe8EnV9u76hISjDiCRIZ1jbXkXpPySDSa
orkHg286v6n0pANJvA2bkfiGO811C/pmsXZklSxsect/xybSmbodEEqiKE+Iju86
yM6VGVuCJFNGOFkSlPaQlrDDSLy/nKNNm0tmUjmFnQgVO+6sal6+4xGVTrrOz4MI
CqcuaAPPxl2nPaUY6e2qH2VuLXqThl2+nO64BIWjRDbSRwi1VaPtbhPJnOsoF6y+
72OE5q0l3NMpiFc8hrg83nzsR2doy9UoPMey1fOOys1qamud/olarbmW0d2MZb5X
+uTD6xuiOwUIOn7LZgJNp3DpjmVqOMttDVSYp/6SxZHEoZyCd8DfCVQy8nMPtYUw
9F8nWz41Ka1FoGWk7Qumzl2slI+uYsKrJJ6OEQSnj0vGe5OwrT3uwUHETjVLf5b2
9FRWeRXP0FZM9wNWUX/T9A==
`protect END_PROTECTED
