`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6iVA5L4I39wL9e2ys/CmbZQPlvyvMRI1Bpr+4Ao+7hRHTi6OMjY1RwsA1w8pnLCb
sqrZi9sXXaXh4KDGAhr2cqsfUpJdflsPLUjPoWMsuimyQ2zIm+Irj1Zx9NXYDeER
5RpWBfY7jmE+KBQOCimzMex9DdrPpJ07bylIuUSPNrKz9lsmvXRzOAnT0fOj/cpr
3coYXUzMvHxkvnwK/cIiuLiscV4tuV3lbWBIf0Sw6j+BOSiOPBlAXI3iPb/jS0GF
HluQVFThtyPsKQiqtJyGRVLyAsjA9eN8wrRbNQCdXj+XKHOIueFmHUZZZCLI90p3
sOkGLcwFGCsrHq9ovdV0CK1hYuQxbP5RSx9ACoEweyZpmmBQUj7ZZOl8tQegDikC
DKsxfCCwoDAHf8FEZlJ9eKpqieXL6edzf5pYqtyADRHFFwa0ejmXuZhCAXt5bb7K
n9iccstiRnt3PSBG/LiTMOgkasCpOnNBqgjHrpWIm8mLPfCWSEhW5E+nsFoufL8c
qaAYzl9TcMo2UvyPeUbaF/upxLdu92Lq10Z3swrEnkHTUPV8ZG8c/GG5Uewlmpwd
AA8b5a2b1MbYk12BkUvHhH4y8Ib1UWMkEYpQ7p0qACDy5axeP6k2g8ti47fmiohS
157ffju8D2NChX5BmCEtGPjt2cfB/PG1o8JLmFuaC7msK0FatKA18To7aYWEwqej
ZRabgaLPFKB7LQOcpyGsAQ5fvCB+3Cx5sDsIJ8Yr7x2kacy37M+IwoRV4GgMnTl2
RZ4baaJJu6psqNUS9xF5qgadHpFFx5tcCIZmvBuNm5UgRHfKlZKnW1j73fWdiFfD
yIhKjbR1Q1JMFGd1XOXvVVLsHPRq92/syK342kyGbl9yITMu74GJU39FPWfFBwIv
jkXjv6ICMHOXjL4lmZMLuQq8g297/9bFxxK9iPnNgn770paXZ1D/3W5yIQnlsDnE
Wo7kDgfSbP33/hkcRp9vQBPlAHJJ72jMa67AV2gp1xgYAXM4jufU+wIdt356Z26P
1Pa+MAnxeJNtVir/Y2XWQ9sK4TAKYgADcLlRY0m39d3E+gi493Xm4H0vT318QkKe
EGIxPtumOPu81B15C1Q8Hdosz/bf9ibwP0lKSnHsdgAj2tkYYyRVk5jFa+dYxTFd
RcOZzg0nLmJ9BAmK9vFslDaWxKmiY81iQb+Z03uCy6Eit29Pkz8G15/hGHzKRgct
8f4O68xju5uozplwSUMspGmpshZ2GyScEnp9rK8QzxnwjeI4gS64VCIwtUgz0ixL
`protect END_PROTECTED
