`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbRnzXo0oX7VhPYP/EbGm+oBzynRys6e+0t49wd0uN6IVED2Orq98oeyvqgraSJa
hn/qvpgMl7R5Ke0O/AwCe/x1xoyhgOla0AuQnD2aRo+wCVqtN4mI7VCSJ1dNIif2
u7ZgjT3o/qLlNHoY9Ut+DhyA7h2z7KaDQBaat+bIsmxXQHVpYa3aao5nRS2oSRdr
/i3+LSaARstNRAorscRsRA+qQVHpOc2bP0I7xYXwxUjdTRkBIUJIodIQVv8hKI3g
/E1nQbdTJj46DC/S+Fg6/kB1aGO354BGaCIrEF4T5X0k22PG4BPoUEcsc3fWT9m9
C3grue2CtMJ1f5RTmfZALJBDzLNIm+W0Af0bx48ywrtId7N/wDa7/UkJh3FSjwVx
L6scovCPEkgbenPc27QPQZRp0kOiQ/K+70PjeyjP3Dy1yUBx5g/ssoXHZ9QsapBo
EXXZotTjr+bG12ORaTBUt0JpO/QFWcKn+Ws5J9zJdYkuXCKcjFYS1Dy3ucVCWHq+
x2LX6ehKzm/B1+XhNWYj0rEMA/8pUo+tKB3Oc+bj11jb/Rx9dC6sbYiT+HZcB1ca
l3PJlwS+eisaIGL1Vy9/Nt8CWrqj2YqcsLpo1iYerEzb57bNG/yagLctpX6GTL1S
w+vzrhCz5ArT3laYn91H3Ik2bR2bKLnNRhDqHzMyURUlHB/7IKeYAyJG9DEPtfRP
gtDeggUcuckv7tG0+a6+Fyi7cbvG04dJ+Jmi7oLVNe+0qrCwJp9MOPtnUI/vFvbR
lcH7f+Y4vwjRjnqXEZe6k8Jii29RkGGJIUsjbmwK2sw=
`protect END_PROTECTED
