`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXO+2poR7LZY0jn0Pt4l37Il3MajqXhVcNWl4zdjAtHa0skGdoEpNy4eS7O0xFNo
gHKnw4tu768eTd0bh7X0/iKv89luFHS1yrogg1vn40Nz6V/t9pgeHmxS2BluzDl3
lHfX4OCFaBgnH1qAo1zn2VN0yIMIGn2G3WXP0HAHe/Lv5B415bWce0lgJRq+VFhR
cJ7G7EyCmhyEVOksbXS9cViZfL+hcOA5xEwUfUD8HkWuYfN86FwIIHwWJXc9IWJQ
UZQgV2qr4BypQIpf/5tsTgPH3mdKI2m6+ejbFYiWH09a0h5Ln0yWj+l+KD0Wv8sT
ojeOHt6ygenTR7ufa74mEjdrLmxSV5sntnMwIJTyi35RSH7KfdqMknThZ0sp+lKY
ujaP8RMzkWhiq91417AImi8FmbJZqYU61i7bsS/HTo5e0GjGFQaI+SHNUbnkRlPC
/5R4L906Sje5QTsX//veexvOu4iU6Saf+AICpqdtGmvJvOGbMYRxKZVRwSG5O3dw
AbL412g76l5zq3O+BIz/UKvac1y2MzqIfgtenD9kHv+iwHSELUa0nAmfQGnQNeJQ
hBrZsKIU4Lj8MZVpbgGwNe+xjexNlRTNZuXks3Ro0DGiiXetYuP/sR78wKTGyiE9
5ZV3fKZLdZh7as5kvnYVoHDyaWkAfwp+WNZqWZA9C6QbcFIp843FKzM0tCuh+3ni
3gPlqySnlU1KFr+GED6xFRKIZX3aoY+MVChB0GlrxrOTwsxnGfvPJQD3L+XsF9M/
+P1DUk0qEzUellAIkw5YFTdQhGXpQCh3Nl/5GsvLr2W5gXrr9UifhnmxjjF3j8vg
y2cfAYYT05JU32xAPEReh9ZqL3b+FUtrmU3IrQ5CNwgaPgt0zkiCjJ+vf7kWvwUQ
BsXikwT5rIE00igsuGhiC6V7ktcumne/I9khjHrNQtiJUCVruTif+POnvw7cArL/
r3BkhBkBQTWifJ7GoldAsHbP/JW6WMuOAAUSBQxhAXIRw8WKCWNm7p8ckGt88dsk
1JxLKxiDJVvVI4w/vBR6IkwmdzdcFIVmZ7qUtIXSvMAZ8uOyhxf26TFwMYQ96Nqv
LuLzBeCFlhbdxbu/jBeqXPuUnVdGQF7YdRHDK+h1Axdb49m0WsAsJOwlzj/LdHWG
q9HSUDSAKTULPr3akxrZaxtMHrEL9Z+Qh1hzTsR4p0A6gVU15MFRyn/pDJ6Yvf89
qqwDuioTjFP4bwJKTpNkSv1KmDS6h7p8VUgccV0iONA=
`protect END_PROTECTED
