`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iLNmXai7+/hljdaVnP5Cpjm/ZClan22Y5fWVgCTItsPQ/aFP28cj3i2KYC6UNJx
nbrfgqF0Er+GrRPTeogLVCumQAzQebnGj/LhFWeBepPvKDfNbFpGZhng/al7s7Z4
kCl0t0kdHw51Ysbnd+o5BPtROxaavqY0ZEx+bCM7wUze3bwIIoV/3pSbOfvOrXbP
0q+pnEEH+MYX8hqqZoFmYuz1KlLEYbk11RE0ty0vsoBLLW49iXAc9s8Dm5ilpbI1
FtK7T6o9cvvmLrNRnjG+ABGfONCiahkERw6yrnw6dxyCYyar1XI++BW20krl5TaQ
B7c/+zaAAegPb4TT0G7mp2B9LQ6s2uAtlEEtVkit/tH7JN1iYcqdsZIPf7I+iY6J
aXiNEP4Ybgugq3/Kt5Jq40+e1HvT5jeMwk3zHXoiyGaBEnRiIDKfMTnl/2GYYLxq
BRGm2NbIkjYXGXq9Y6dI0l3VaqfcohHrR15tRefF2Yh9cPGrUwaTDU1M/iWE8e2i
6JTRkc/LfUJKbcotxjIAV92b6KT3XGjs38bI/bv/qYoS47Arkd5pD8+nZ2/qOeHF
C88ND7mN5n74/EiQ8dE1uTTWe74PxE4cm9hzGnbQjDU4qwFYk6uLVuZ7m0vxWpuR
YKAXZ2ThMfdKtjeeAYQeQJl8Ia2HJeyQiqcKclsCn5ON51HHcaTrvZ9tpKQmrXUL
CIP//LFENc70LcpfB5Zuh/8ULHO02ESkNh5q+rnm9f3RLMYwuaGspUgcNCMujfPx
T7jXe0A1Euzd2OLepfZEtHuec+QBPamRqO9zdqmv6EzJbWv+B23dSKpsGT+33giv
3Asj3PQ8+0XwVWSKdTsjwJAhWAfeSUrFCzdgbdixNj6JrKZU+z+bb4lKUSQ7DV1q
n36omhZp82P2vVRaGXdJgEJfOPQc1AGsoyWiuo1TPV5r1dFcMP6qRMd8c1MpjlhJ
ufMEZlUz5Xvq52XiknX/jO4orZGb4F9TrjJ7kkZ7cqQ6joFCMyd19tF+jfH14soh
WojXN/D4c23+IS3qUNIkXgBYcji36guUJUoJyxxUOj22J9hsfJ8Ix9Cw1hkwWBbm
7PI/i+oc+T8iYjoX4C39duJTFzCFvaQoII9Vuosaqrp5EZRTGnL+dXkemYQ55/6M
Iax/TdDmo/VbY3lCm/l5UnXhXTebaF0UEUnvlMT4nFsCcWzzQAtk0dl0ruqodFXk
cmFy+uYlApqFST1kQJyW7+GNDfXODHrvyEhmGhK1KI4Ha3r2votSTwgMG/El1lGL
4WNrSuqQm7o75WStzYJF9Z5dQTqYEkMl2vmd13fxePLzmbeVEgp3LPhwSng4O5M1
QGH+lHcnZYfs97Gg6zlIn12Ug1YWl7XxHWy15gYIiQWkVK2nRK8ftsWZy9cVVJBH
OsxLr+grpU008W2Qm8kBeNJIfskMJbR0Jzyc5Cp43D4dF6nIIQcTiwsHQDcFfPTh
xRj26HpJjyphVG12xHMtbYz25sHAmpkhFnpTZZYwSMUK0aCOe/yG/tKmUR83TLi8
IjjfqTVp8NCpYPwKoqmyGAicq26e+VFDhm9AUi0U5eD+3jyUEoMe2WgdenPqfnGH
bup2xDzyaNNDCm1CKpyDN5lHOIimrrCp+2OQ1cWtN8i8urL2IMIJuYCNFPXIpMb0
DiRRMV/rbHtbylmzFdd8vDhtnGjNeBum4K7ES6Z7TheF/islHXMA55t+G1J4tGFy
xN5uOZ9uTOcl7WMxoYwJTUAQN0TYp/1slnRd2H9fxjY37crz2Kp+J9csW+3ncVPf
j65YDOVlWc+ZOE1SbIGZnjK9mIXk6hkmz6mQGGYR1cKiPM1yd30XTWZkjnwtnsov
hz+rg9EoQ2RF6k4FIfxQ4In4bjUpP6GwV6s1UDGwjvpWdsvVtAh6AL41PoNhxIT0
A8/3pbELxgRLyUtzUlkw6wktvM4V9jqevQGw/G+C32xy4MmcHScjfo+PIQcAi7Jc
GpAzy3MFfAgZk+EtHUqbw289umji85lhLeZMxpbEsujI/s+ga13ndssg6uQY+L5X
12NWmWG5qvGWY3/DdT4cgU6hLyfo02YcbKnoLE7s0bkKU5MW7QCAIAen6DNTxH85
mR7lCmr3o/YyJ1EjH8N25PtazMuL5dtcCE+xliK/Y+lhqzwnNkoz7Cnt0t70O0yk
KyNEY98FtTdcmxjdWUGNZqGyOTYgAnGk/xpY5fUgHz8=
`protect END_PROTECTED
