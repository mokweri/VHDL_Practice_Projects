`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hb8Qhb1i+3vcKuL9ymYfXFrRYoCkKlZt6XDtJf4kejN9glac+VAfu+8IO2KO8eyf
IBmFmWf3WMZvGjy3jMfe8ox1TqgklMefWK/lHaZTeMg1+vyUCqprj6bsruavmREp
8iqmbjLsqsqhgODdRDsIq670k6onG/iEohK+v4UuM089cnQ/6mTVda5SW1Ozb0z0
ZVTrZ26XsJ5/eWAJXdyrj+lNDJlgoMxGpFZbnrsYI19N06po9RJQguHkFTwFlyro
ZW1GXfe+M+He8k/jWDrsrueIxVrDy3XKXASiUvJGPcrOtPRTXcrTquas3lTyLAK8
eWpqrAwrPjF1XqkdbZR5GbASM2bAK2SHaysY76ORIexW02dJBPMyskI72a5Kqsee
hz7l2Ca7o5bKOsuRw2Twf41CbQL4GK5le3jzM6yUhEpepZyMRCHx89jgVTNNz6s/
itxLAqb6Pb8r+gRRhgWBWk/zJz3U+uNredtKn0lxMGhKWzeg6yCM1xZ5H4gEX0xH
jvBiLk4doWebTnN3a5np9KbwFnaasYY1JpOABVWe9DeO4zlL4v3iqWmxJ2LS6M8L
dtvTdeg6NykeWzMp+qQwTZaRSnfkLa865Z2NS8teq8ZrtvCix2BYpp+qlBbQLU7o
2W3qc+8qPkHyCIqSDxjWHGJbFtbUoeOSmfebi6ZPuXdouR79TTIORQ6BNqRD75+X
rrQm1TjeRWNsvcj9AlMFiRCRq9/xm/Cxf8G+crw+8kjzBKvuToovX2k3KpcdVvGL
qVHBY5RUmcN2DbOVOJvxVJb9wdMm+jM/lkXGxqHZKdF8zrUllqPLzCxOdUB8nU0e
4Q1wWaTEK0J2k4tCeAYDJe3THUbS9IUBKHdQtBlSb7A34Bw/rS/ll05qC0r4GmlB
urkOrEB4BWPOmV2/AgxYoq/QMiEEEfKvuPLHDIcX0l0mz2rj87lu48LxlZn5QnR2
zOJd21d1W8GllXar0nkF1ePKo8D0i2UEBPD3XFqZszJCw/Ov1qTQ2ycBL/hEF4pG
Pqsk4MlBC8sYTWGWuDIqZBU4+zgZyHPktPmBLtnzKe3J7K6+MvT317F6DcdJp6o5
ThIDtJrkni+hGg6C4QdlGYI4lk9ywuOpEqAh0h5tDdEDhxFq5xK75+JwEjrfTfZ0
mYkHELjDJfVYu8/Db4epE6MJKkmVXZJHw30K0rVqN2nULLbEUI1WQXW7auAKUREI
HO+vhCYgbduSC0DZ7VPlq5DRCx977HGDI+yPaEeBufpvm/gTetSMvQueobfmBu4c
l9DTkm1DQhsC3XtQt3ihKuRIO1NQ/T9m/pchjdJP9LxjZvNU3lurZc2Tca10aU9n
V1/3SSufm3rKUZ2N8GBXZtKi+A7xHmblnRiEWVFpkTXkOr5hkMqh+fv+jt93hNAV
LxYxLGWGS99pTlnc19Gd76IbnBEv6Dd7t23td6mFAmqmaqIpEjgOLz2tGKNDQ+P/
9MTcP7NqF3k48+LTyfib2H7xxt4GSkrKz2NfZ0Aehus=
`protect END_PROTECTED
