`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QMA2mY9dsksOQUiVrxFX4Bjgwt9+M59lFQpb30d2pd+xOxaYltNhXKJcmOPATJxL
ZCN1yj1v0IAJMTytQPZ/8ABk8J8ElnXQPC6myJVB/IlFxG1GJ1QpxDPFbJ6FrC5E
jQbYQ3ed2eVQJNd3d7Dlw87CrNNQrJLWnY9Li4ARETFJkunGmijwXC5VYpcAkPjL
aqSOW+ZOwCHAhO5ScXLR6ocOis9YZQSMzVklTNCCyI+oJ42vVYOImKynhmgJsE1+
oEcDyiZZ4KM5KPJ5PGvtcPMLEkpUwA/rpY2iMH4t1Qipano9RBfEvGp8UKg4jQA1
1rkI1RdLTCCu9Cw9x5+ckq2e/5qomy5zOJ0t+dsLXQRGZ2EWPWdbAOKoImFpV6Au
4/GJIHzxepbm5md8SLKCtT4KK4wNtjmgRk560DMinKkOQnTizit4JZQ8bPEI9Q+G
GNnXSht8MO7lsPCEOO/fCyAcEyAoKmuCI4KsAq6f26A00LyGakXSNpZUNcd3q7Ts
EZoiWZ3ulvWf+5FnocfBfnbwQH2/ij57++JjzrGA9mu9hnS8n613J78S/ioiivLp
mejm/5R9erPrpzXuzJfrntxWj2F46blGL7tm29UmZwPOe4wBRgWUI27IQPHDvJLo
z06ydBtISO8rL0Xy47a1S/l3JF6lmWtMFEeqlVAY0xA7jDHOrrcnHeZokJQTEkrt
zJsPPblpwxXiTy6F5nDmlop7Fldk81/o8M+pqFxhiwk1Jl762WcCvtcMzMAJX6md
gPyCmVj0dmz97Xx1cacFtGKjwSej8JYWF82toV5dHM0NK8FZZc7jg0tKs8pzwZKK
2ZiTgAOd4vnbxruxkqzDDxCizLTXAL0ucC3jNy+b95EcOTNe4WhVUiBYvTTQTdfd
bKFxIguMU9JgQeuANJq/AjqlXRB1/4iEDEAQ+NnvzFc90uJOJYaJnP8kO6s2MFYN
IxqNV9oQ/r1gg0OhaQM8X5Rztba9Dhe7utvrgYBSu3Cc7I3aSP37AC+q3L2H1BJD
ealPNWiwtad/z2TVwvQ3MatOc7laI/EWdu0nY2yDw35vO2AVV2OXIeL8JpMCMhos
YFFN7pPL8cOclh6JDUCpneopvVwjvZlVzs6CuXqV8Yd6pN0WrTitJa3l/zcc8X9R
9gRfjS30Hvoua2mauHd7e1/OsEjO96t9rPFelHQ1gDpnWFR7bARlY6u1YKYvwxy8
rDeFdpqAc72Dea94Kzj66tmBTZRcUCse+Eq49pXJIX6B+OQwi0yBlMl2QJhBGsif
QyZO50h23AM824R4QsQz0eFYD9+JYQ4tHCg/SVoldM7hl7H6q8meAnOG5iEU1JdT
zgHA6vF1+LhhjiwIo58FgZcTJcuYhR6Kl+mcthEcYC9HtlHBVV/hBw5yCt35oZbC
5X1UZ33NmHXhjQAVBqsH0o89uMqjjXZuCCR9Nf5nTej3A4obhNS+2kMAZuY+/uZF
iE8IT/03hsOAsTrIgCBEzTF2WQEmzGRWh2QooHWN5lS/IuIuC/goR3OH1xdR5R3b
VytEe4JdXorHc5FG8RipIBcS2wT7V7BMbz9aMafwadt/Vsto853dvpJk2U+qOhoY
vBnLpN6cPvJu2D1Qkat7ZAx/Kn7nQ9TJeuT1zHQvlmspQsnH2ygQnQTZP4WgcreL
Vquu0gEYLDIskWDIametKETPrydyzWoi8ClQYNsEVQRf70dSkYamvamRPtuEgToW
bPrCvcXcx94hfpqSRXP5zFe/6vLLwNGI2mcjRM3Ru+G0VMPUZhPDJ443FrM/ebFu
K/Bt0qZGh2DpDz8khK2xI2o8jVewY4HZH2N8MyMe+tYuZZ7QxOGiGgOMWYXAGH6T
vZLk5n1Gq9Fdb/XeLq+yTKEOppY2jjQLlVq3PAq+aOkABCFeFYr2fMJx4xPs8ChV
FDLd989HI6zcWIIMQKR0GcX0UhueQWcsTdTyqC6WHJDDfSs/crIL4jP/TluFcLYu
xTVCah14NjASjuKEYn16MfqfzMNHc72N0UULf3R2z1w+N9qlAOLBUFNSkkCwveDI
OflFRZYmw13NFyLsiBpwTbvCmrxN8F5FXpn8FwBvmgktklVrclUus39H0uFLG5nJ
OoopgpLh3fKXlIox+O9k3ODOTFz10TqkwBsAYEdSm7VB15nHQC5NNHMQVVKSdNfo
uj77t2JReklddoO9aYp9YPaOvLicb4JF7+UynR9nljafEhwAyZVhT8tr0znejp4f
c1NqPSSjZZeqiV4fJKeQbyC+FaKRrwijnBF+tlkhzqkcps4neze7qBp7LvizeH18
NRuu4DHNg65s+tLN5HNQ0Pn3o9K4jsCfmoahHgxGgBovj9+2iw8E8ucPPZRFhFCt
S3BrXfyycpHS7I6joeBq9HR/De+rOUK64cIgCUaYYoczfUksdQflPKarIl7O78Kz
BY5hBtCZw+KXU162qk5QcXX/Ucn9yx9Wg1JpATgmCb1TJR6ZKTJtQPDKe5AIwBGk
mLbDMwl0zLV/K7W4qQtfz5FxKv0M4oisX5nvD5Bf5lYswqlxV1z+BWZVvghQZVC6
flbaIu9l2mTfEcyrJFG3yCD1pkUjU8EkAPyn/ihaonk=
`protect END_PROTECTED
