`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjahgxYy+l8LIiOcC/F8yov2CbNTpGTmA3PAjDbsBvUEfhBdW73dPGuwfpvcz9vT
RlivmYXor1pwWUV4CLMWJxEladHpmgt3bXgG0c8Xsjw2VCr9Uoh6dMmYLTNuWRB/
HLqHzsfBbh+t0LK32O3Z0D78DDToyhrwVg23avGLhmRhgwLL00BrZyFbOZMo5zEG
VKg39rTQfcuzTSc0ZpOOtwDdVvZMmUMDzgtioeqfIJBt08kl6qBAKW7ZMquLQO8W
SAYRiTXiEfoR4aFvwuU1cCCcdHRy84s3n4lh+HcxqeMY0TOyXkLdAexBEElWB6eO
pUTSaNsDEzOQFeqjtQxEgyaDHxwbIunbHA20J3/i5Jc/CUqBDvqZyh4RoZLojIRY
OXWMTFC4AmfO8vP7a70PGMG2h9RBrnRWtJ9wAF0uSqlMRf8cOKSK0mp4BCzGvqna
grshOjKb24RKGgTNpW6d8TR7D3g5dZFCvP5jw/bVcZOE2e7cXHVwzuQR1R1Z/+9F
KCzseTX/E2Dv5mmoeVhO3Tk4dLKVxDNsqUtRasupU0o23wHt9slXUcOqGZhHCOxs
U4skF5lT8e/aMHqH0JUbiVsXKa/7av7k7G1jU9SbvcjecTr/GO6cUvrct7LQJuc9
AYmiP/ztbPrce9ln6k7MQpAkMVvpDgqGGmjCAaEVoXQc0JFhAh/1iSe0LG7nU7bo
/pdLg2qdwxHwl1mGMQwZ8hLM9V3p+E2XrkX+eCE4yStUwnKFO+jHpuZYzuzVIaJ8
PlP2yN2MLhUi9xt75nN3HOYxdWRh/UYsklEKpXyJxorTCsCU1pMphqeOhAQSLXKY
0+yAoQhoKFiexFari4QqHDAJd1O0cz/rhigk+eFigMcS5iJa9RI7ysIjvxrb4sGe
rKwVneLki9Ym5kEO3RA5fA6KH8eTiSbvevcDPVcKNSGMawwxNfw05u/x/sfNfMWQ
1N3sW1f3WpnR2VBNOWIbTHH9C/Qu8Hp0bkyTAk8bwso/PHmGTiu2mquoEXMDks1q
ePuyvOGvqoXIdLQv1qTYN7+WQdm4NyPjwMyqcC5lm6e7o6edJVZostUVtVmnrqDs
WoDMpWNKYCyQkvnoy3yVOv/ym7btmCaZVj6TeeN9ixiwnkbCOaUWX+nslQIhlUUc
XC+Lgn6g+TebR7HznPygGuXPXI6xWNyj6ALGObxrGBVqqmL6n2VIvz17IZ1emY87
QkECha41Jp1uUI+2+lSeFmvo/tcGLPihCq4v2/MuLsx150BLpsMPeNw0K+Rr2paF
hZhmmGJt4lOPW4Z0oKUfeFYdKGOcTyEsjKTd00RX9RgD/ZcH+BSfx1K8VM/xlfWl
58j42jc927AST1ZmJjYefemYzNF79vDNBJf3Fy9kh6DEEHYEMsspIc+ZzbUin+AD
cQgojrartaqVwmX7SjM1WY9nuCsZ1ChpE18U3THSwWoJUmOf3eru0HRy298TH3hx
LdQdfdfccGZsht83U6s5gAqZUuHxylBhRv7OBaSUfdq+dfcO9roVA1jrOZ+l7Iba
F+j1YKLvyJGlfTVLTj7S+s+VdnVKgDiocg3ViWG4y7L+wx4LGH8lSOQzp5CyqFVd
FsyV0OpHnqbwplNAWUsU877hJLIC8+V3NGj4cWpTQGIjl83LBEGkCijQb3ckZKxf
u91sVN8XnW125HCq0G70fqGC8HkwiCEp2g4EYKN0/FCulA8cTuAO9Af2PUQaWhI+
kSEHDj2dAoOrcvwYMV46jO7GePtLHPwbOY4UorIfmr7sHxh1FB0VGCYrkGkuMiSE
6R9L9eHzAwczvLXC8c462n5vrNoTTqS44aLTXBRwy9z1EJwxgvxolLv0nWbEIHzl
1tEiYbVMM72BvDQxArABRtAy8SoadTP73L74yptkQZ9vQ/6LUPD0p/KbS6hlorqE
+S48C40mPi8c1ZRW9vsvVaF+JB7WqwUuwuEGlkoQaA4k2gXuhy+IAN0pmaoqpV/e
qd3cGMCly+dEOSLSNxYQrpIpRHxvH77ZGZ5TAqlbs2h8lQkl6FT69+Y+u7lTmceY
ZO1yKsFGXLVMnzTkKDT2S7tZ5nfZ5v2ryhO84eCun+/pfvPq2lmBgRAnRCoDIrI5
aRi12WZicmGWYeBhngSriyQj+J4xOVNP/Ba5+aAmANsU/mPSoYd7kbq/e9Uaassp
sGHcLtAPvI/eiJsDaKzn90PBdwdKiecoe416CYZBl87kd5JLsdjGdXE178Ft0bct
kBVVY/CV7SjkKqxjaVQNcZQoMecZNjbUJmzAREee1jCLEYkMwwTQkdEHnle1T70p
tJMwQLfkqI0fF58pQl2b9l4RN7hqNIyR/Uoqkeqshp9BccimhOdzhHlI4Wn4qlg9
bIBy6k9KSLhpkJHLkBldiyFv/7XqyK0XaVJY7KFvHW+L4RWaLPa4822rBl+CR2en
oq3de9Cg5AVg6+XVWC2lP6TWR6p7Rl0x9kAGB9OpSSo9iGkSoJCd3AQ/hDb93TVB
nJFsF7AZ9yZjN+n0c78+3Ec8Tfp3Ei4o0tspUMB0JmNKB9h5E0FCyF4E/eHaODkq
KgxKgW66NgLhKK7VgEbRIpU1hJNtv+wVSRNrmWJitQPHw4/8RnsA4E+ymtQDtqg4
kaTNoHThdZA6JfQOIZDRiZIGRBdMgpKVSlA677wd63m8lmYCQYuGd8VA2G95Qgqx
biN+eHekHTuD9kN1Ev6Y9QVPH848tTJmtpYf7RM8mKGCMBew+L6RKuj5ffvG2Rr+
2lCfi5d0KiMefVbjzaVBWoVQrjft99DZMjTOULhCMBMLp5gtLjA5k2kWf5vJqOwK
n888nBBZF8E5Tna4n61bWGjBhoexkj+FVM2wj2BylW8yN3pOSUjAJ6pqxbOM8nnY
Alp19If7ssXC4D7PI/0OtsGFTaS+zfp5TFvoYUPw0m7QzmCcPA++V1G4Fw/PFVKJ
ig4XOeezBx3SbPwkizl7IypzoqITEvaFVOf/32v3HECO3SuzU97Ecc9f0TJleYkE
7By3stD2aac5hOoy3I/9f67rXvv9CJxeCMPU411Wmo81JWDGLhWFSjjbZDRAfpiz
dQKtB8v3GsDTy7CVA5sh/+C8xcnFgWEEJqUnte4FUPTtVMvntg1H3qWdSbnq8gax
glF3Gy+w74BvcwdqWy4gvhgXxC/llLNKzRxaFmuqtR82VrztK472PzZRtjl60Lu+
1c4S8ZIsfYIJFNTh0NNOETKPwWCwv4NELiEP5OB8dxPBR2H7aRQx0rTg7udmNmna
3a5+As1x448dWSfJb7OpHizn+w1qqNUPlWYIc45Tnfx1bSSitE8CtJq/TL+x563Y
rec/aefinMWBXymbMf9RvYe59LyjXpkzr5A3yTsXNlk2w9L0gXi91FR6nlP4zsOC
jOluYZ7S5uqGaMY0qPCxVoqA1IfiIzkUQdNBJFvBoRSftuhq8dx8Kfskn+gEJx30
N/sEbjREZkTW/1cpO/BGHKkS0932KVzp6m2Cimuxo7+Ci4vLE4b+pfUHENl2/WzO
Ph3RInWGqsLAhCktO4t8scAUgaITm+F7n1IRdJL6X95n2qqttihn23oX5T7+YguF
mDKz5maodj/SMkZp0GeKr10C1r5t9VwujLB3iQffm2cnmKanOEoaM/dENw3tjHLg
Ph/QnAgxGLDheVaxWcOS+2gI5Whxv0ucNe3FSEVAXD2zPoBjjpNQZS3jS1eCdh0G
ZvTXTxbVnY/dPwN7VutQ6UlXAds/zb0ndOZdutNd9AhaqR9yS15QjXf3+7kgAjBx
pVwo9y0Bui0eU8r5zR25jcENJiwWwag5vhxmdzoKCRTLdjFmCEo8p65Ot33uPgkc
MGQ4srHlMAVDl4WoHM53WG3Om44jIpFSlPVfFTeZLBc5A9eFHvxUiijUTAUKb/GO
odhIAIvc9Ot69ZxkETd25R4KhnS+JNGUudR+XI3i1EVNAOT4lHd2ZIrFVMm/cUTe
SoGjHPn7nK2vd9NcJuspFNERutxQl4Qs4+4seRx7iwFvDKdZdsINtwBSDAhBHS/l
UMDB++Gz+haj5XuhWiaZedYUvgblp/sXB0Wl88bDEJm4cFsRzpRzJzIHOb8leuBq
kZNWLpfRtzzNHQu3u8D5QaUVFuGTiv9N012LTDlwAHu9RgQymvGvUWEITS2LwdxW
1EmFUVC9RcSxLA9NExfci4AhcIgVF4uAoYuw+2e1Teewbcz6jy03simTZODzHL96
yGtCiGfLa7xS5EQfh+YrFMeZykviwXBf8aTIy1E8Ou+SFaqugi/Tw5sEyuSmiJd3
v7zKeSbeUx78sPE/PnItR0m78clayC9RE4ewA0xvYTv41HKNtVcAUiW8pdI7sP+I
ptyWJo8yPEoDyumPjNKxWk74oU1a//a9mMskP2H2O7HCrvJmfyVC3gF45Q6/ceOo
yOj/xN5fd13qc5id06aZ4xd2p1ngvxenscFmzzhVFvGVspisT85qP6sgMRzZ8z6E
BsnrCDtBnS13+YvKsub00yxMiIfzQPa+TncmfY3W8aplWJh34chwjXFYGJMkG+Qy
zOgzlljigid1A6EQ2aCigOOcbDXvsug3FSz9sLi3c2ubtKjIY6oDdAPKNd9RdQe3
OwQ7Nh9atqAQmBMqGry7v0TGYB4xB9C8bdjF2m9HTYfiKhDgWslUVHhvoLfjSj6i
L4ug2qpyLfy22kagkPUvApEPvEujLZth4Wi4TmRjKvauf3xgLa5qnsKj8Um4Od7k
3S/rrr8kXcJv/HkzVpnTyUnQwVioxYDc+qXw3LPjBYv0a9xw+H6nfokLbtwMzPtZ
5mPeuwn8WvF6rjQdAZxH/zcN9/slnuA6uu8r2HlNrar/xO68wPA0aJy29PTW1MMb
nAMrtiikvCtmt1MAaop76GhkZz1sfmQd9H2aBhXfz9BKtpNHvyLK0PTj+B74alVN
hRDxMTvtdVMqV7mhdYsEtB2eXr7o1B+V/n7VKdEYp0/SY0YbFOjkkwMjwwCv8d4p
Yag8fP0Dtjgvmkj1xjrMXt0hFFwlNmWeMBNN6kEPTfgted2ovWpYePSWs2dcceBJ
NFSgm5xWLJwESite82NAQRhbUT6ScFawEjZvcvCR+gqsg7jXMo9+uTBRRFYQs/jj
oKhas3oyXegtL3svOWZ5vn71mC4fTfSxrB7zIqxnviPkufAWGIynZRjO1p+3hUiY
PQnNlcI93e9C0mQsCpmXqfnQz3/IBOmzVCOJvpTxNuKKbA0TYdWRNaXHcfrRkR3g
Rwl3JII7RY3GN1+8zJShY3Exe2AMuBe8VyqvdC+PrAbXoOQM6CE4Jo4YlsWzqA9s
ecC8qMD0a83iiIW9q475dXi4g2NYCJ1Sne6KWuC2bOwtJp0GkZoOb+92Sl7UjUq0
Peesx+TSiiOeFXUKcHLfvY+pA9t2xENC84dfiSQwlOEGt32J6JYUlhGhPp8qdBfJ
6i4BhTjKn/pAXGogSEDCDeAMrALTsbNnjia5nM6WzziZLhgKBL7PS/yl0GCp0mzz
uZXhpwIreGHiCsolm5Fb71ACiMbT+rwvHfvr3q9KZRyeax2VaBasRGG1JIiZs7Km
iH4BKXV4fzBQYYD4wQ/0io5JsTTaRmHNVe9jaEgSzFmGsmeVQvq8u/Do+Nvc2PKu
tvQ0sNnL/pngq6Io7X+qfN0ue+aUdvHItZ1PVSC3P4Wisfpx3GFnj7VCXgaMXBRX
06KV1fCmL6mlGHWvvCIb8HHVq91rNLjt9V4P5UtIviQVG+Ukgabb+EwonPW8gZMR
O7fYLG5LLIZXiZ4z7su3i64jbOGRA0S85sP3GoOYJAfXIRK74SuTdG1oZXJ6kvl4
HEjRQDK38VgJTlmi4r/zDpuyWn02H4utwAkD4+t4wFC7xxkw4yGP4/1bZ7fmTDM+
mEmInOVCcwerN5Q1ShvTSEyUpVWZftuCoV28KVeoPxVrBKuZPgmLitPARuVn7FB4
JQD4Pex0YQa96de+LDrcydelT7IpZC7ifyYzwcVaCatmJtI87NGjTAgkutgI1WW9
YB2tt72jpCK/XFOx3L+MNPqYYwf6ibZFsIgDIDBLgNUipAe6lDxw2nY1uxymVSVO
3HnA9kFWoxQuVhUybR8Jx1F0Mfu5w4Rygzwjj8w8Agul05gViCTEwYnOCB+kfAam
NDSso2x9waSrG4SILz4FlFm0mHoMTsXfyRshsWVUxqGkhJGDZKp8jUUql1GtOCtW
oyc2hOHaysMGFY2NQKJ4Cw51x8jAmAMcX/wNChWIPL4ESfvzPAsiHXG8hr8IT5OI
8lrWNdukxzuOrRveY/sGWam4h7iaL8WSvMaMb6TD97vk+ozSQcUFwj7KGS+CZIPU
9TrfZ1LbOuZ1PyaZ8FK0PlsWIMg93C4BYwRNq6TjZ2HfpCZEXJfYm315xwKe4vCh
O6PM2sSjtkNHvrEWVvEPeThtPxu8pp289poeOOMzYn9E1yDLPq5zL7+epXJFt+Be
gpBAldeiuOZZBGKMqs/huxqwyUmlJrUFb/5ImFiY8Y7NKfj+XGyAFDNU65r1JC0g
PaKCsRS1CjsYLDpFP1XW6MxcxAbD0iIAKVACWEJcFOciDS1F/wRglMUBn+WDbZL0
ML/GCx1p8wL1KgVpsx71CU6g8axIdMiyQNcy5gwASzNfikx2H/tB7I7wcZO3QUAc
H1OsMZ68CbGP5SGXQh79ZtU1jKqCYONvyRrtNdC0Dsa2q3YDqqNp6eQ8hYtt9lQm
CwpNCBMWs74klPIfAespLdKM+rh+n1UneLKODy+v68AqQO3vlRgoTd13wrvtjHs5
pvGWBu00+Gq4WlCZzgdTT1Gjx47QcywHYgCy3QSJL00ZYmyap5JHCiq2dc9F7oZH
bs9y+vjBI7fl880of3OicHZsFyIUJ7M2TBkHG8ibP7oXXzbRZNRr2o5WojmPruAI
LAutm1O3QUW9HamWpY62vJBG0Ztl5UbsV72Y3QP5NZt0ehiwJsnII2+w/X/llxpd
YGlAcUtQYN8VsU8A7zvEvSj7psnHuvWiYT7cWQZbh262jBQ8J/X2YF5704zLP0iv
JBJGyn5anMvt3fVCLFRIn28PpqQ47nAQsxKoX8Y2JoccTrBalk0dyfQ8/TlAbhRj
KHd35vjwJZztJPXLwf6cgQfyibQy7P5g/ewoQnc0w4xnU1pVfKCxViBgGFETLLi5
rvFcAgYJ+0+5fhUseA+aAHxbq1jRcLXuVTIfANgoMbR82HnXZgIoZbkS6pZwGhCT
mUIn3uV533FtQEacnSa07E/k81Yh70BXbUF3notzkboio1lx61fLQqHGFZing35d
O+kRW1c8qWMbdfZ800jsRw==
`protect END_PROTECTED
