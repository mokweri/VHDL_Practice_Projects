`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/YUpQOk7YYbYr86qLtpHj7bd+AnWE0Ij6WHEU938GgxrHIfMPHMV8udxXNCzqce
qcvCxkm8B5eJaSeUEOA8V+dfWgOL3Llyibu4mrxmvoeDNUh3jc/j1UrWmD4OgwHg
fw/sO5hGtnC+PDG0/ScHeTB2Ej7L+IbyWoImWtJ3CovW8+c9TmVqoMDXkm9UKbSP
UsVwhong/gpdHEWR2SMGdhOjIX6RJwnSV5hMxbk7MWHriLb9gC4G3P9rknQ7GT75
CYw4aUuB+YISGlMKUZI2HCSVDENH69rr7LguQ8l6ppddQTwpXXyAV+X+vwQG6rcI
WJZcjNFXnGsxQSkV6eLCHUvgo4/P3ZmnllixNzF1FcU4+i8tHr29UUangiZ/SxsC
7A9wqzLF15y2fHgpZlxgYRozHZccdvulSKAALj+IlO09mrGFugi+kCmiSyVzCqBn
mN4bAmiSy9O+LvfmdSLEGn3sN+xgCHbIxbMDdEkmv3sqneOFjjTGMhuMVYG4zKxk
5JyqmLee/LH1ITA07rAJs4zoWiLsdwBwWoZ7yV/vGIBHp3wWHphYhAHPVOWQOy3Y
ymTPJZeF6SnnUf4zzMM0PAYKXukevW9r6LUZ+1a+5mTVuk8xfjwjmSDsOFo/3spW
69iKMczO4Jiwlk3XczK3Z/RVzYwGa3zZz6VyEBrYd4pgSZYP8Y5lCBJGWsKOq4AD
oJs3pu5g14rLV8bU1HBz4YM9KJTmm+hWfVIULBJdJPHWbD2YtIUsyhMiHByDVUoJ
6jN7feTyggiXaUwM6xXBgWfU2IXQ9ckqP2tMJlV9ZAcr0M9iZgqKbgThSo8KRgw+
PTkqP4YP3QsDR6XgCAb4DR308e9BaNpko2Zq7HoBMFmT+UriUASBaFLAf3tkoeWc
duL5RrEFzUtRupMpWpCDuoEeOsHYNhl+8UPfvSNnB1KqqK+jmwhjxcyvj/TVP0Tm
g8EzQw1+FWH4CWhVnJY+SlbnViNwZA7o9bLX/UfR1ETt2tWHQLFk1m71O/+hlBKG
yBNtEIOAA3dpdnFJJTa9f0Y6Ts1i3WxJ+VKfVqiWAU0a0dcbwas7/TUF0BTBPk0X
ZCyulooJ3fZYh+Vapq5O05RHsRPjmqIDkVKfza57GAHwP93h5NWlUFVnD6GXWoyH
q0DmNPelO6J6jamcZwYxAnFPVWnfBmKaoBr1kLNZuR1Vl8gaz9UEiJfpbuMWdnah
SHgdsCAzxhzQeUAAnNj0pOfMjYcd8YMuF4A+0iPY+m+zbvme+HWR7ZlZ8B3Cs+jo
kOoW9pjhYy2juwxZkG4r0YgdB3pPJczjNW2SEQW8JsOzBoDAMqcT3/nFQqrxkJ9a
VNRcMEn2pKL+g8LIi+TRlGPtLgXv5UtfDxMWi1cz/lsANytOGJWmB0HdDSpyi7q+
2DtMTAaT/8p3nXCZ18RQZU1qxtQRTSbjl2YbQwTeylWNmbcZbb7ni/weTo8GzrJe
wVsmsjYSus5VqRGrX85uvv2j0y0IshcEAvaOp37jwB/GFTmkpDGliMNRJHjAbagy
3RWV3sAi0VxC7BVtKy6X9/wWeLQFlADHxlUwYAECskK2SKxHMDLDqA2w1z6EYohv
slJmJ+hYxgD7okF8SBPncqpCMku0Ui0ga5c2+/RI88Vb6oidZtGZrXbbD2WN4hUU
j/vw1QdAzMLlsZOSjfvRawmvEqjdEkIPNnkho25Nl7zz61e6Yltil/n3MRqtTGLy
Tz1OXZIyEh7r1j+UC7f/rrH4Pwiz8q59R2O8MCSKvsf/lCC0r3RrdNmSCMVazQLD
lCFx885hoa+YTqVPa50WUlRxFgW6Of6XgMbdp5hqueNFuyOi1sDdndObZ8XU/eTW
3ox5M4FdGHXrM/CxW4uVsayPqzo5hg/gpFAfgqewxBDaCjYhNpHFbWSXIV5pX8We
l8GjWypkBC7cWF697nuFkzyqCfTcUwpKArmXBVw+wwo=
`protect END_PROTECTED
