`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGabBqUqkZ2jl6wCh63E4kIYPK3DLrDWcnYc08achc2xjk+qYfzrsNMS7EXauGwx
TaHKoH2D1uHqIyDU2JR4Ejh8k/6YuGgexichpRHKEKnuZtAT/9RbAxsiEV7LeD0Y
rnbekmKRsTD2G69bGAAnCTcD/YtSWgKeZYDAEwiO2kbebg28e4VnJ0VeXrV7dXv6
vHH9cxiMMxn92r0Wo38wmukF1GabsMlFkb0aWI374ajfP+lTWqS5tNCHbmBtRnjc
ng+EOK0SvGLfAMlVS+I8KcAOU/nm+mOg/1cPF05UmfTZsdKbfWfEnx8DWgeJ0q16
1+vyoPacjzvMKu6o5bBKhQr37/tm3qIygzeLJz8XiV5kKUYBrB2Bfb9AJeUZBmRG
4yLE5cCr8/LWIo9a0EIC8fSsmR8dqu1j9yWszex6LNzHSeM/wuDbmRVjtzAAkA+h
B1SV62PpAfxS9IastM/jJbEcUF7IRTS8wgEdAz+e8wNRnCW59wxS7PvWu0+ds6cx
60t9zLwIAl50LsG8KUoNWfbJpeBoQgncyStIs6cuMhX975DJRDakSp9QgpaRxGp7
2zOvatIAVRr9FyVBf7FvfnukTjzUzLktZLt/40GH0Bdv97gfJFGZwpbYeikAYoI9
Do38XD6KJFUok1ybqL8xu5yeK/2gJA6oryNWdGSXj2IXj+5AQnh31LgZ9lCKKSI2
ED7y4Za5jIAZSXvbi4FMzX9OcGZyW2BCbB8UqY0AAeFKu9ZZ08aGs+FsBTzteqiY
eQKcyX8vRcW1ZJoqeNtHFuMtAIHmx9CUH/7G/khFJqsKZtq/ZLMrFx/kegQtVbQU
fAqu0WQDhXDIbiZzCTGBQXGFrku1vCsFJ8w5UkMNajtaJili9swlu/GWFOVUJkhg
jtQsci3nEjFNBiaeIRtMDM55QviU40guUVs/RSnACJTr7HX83NLiQtHVLKtioxn1
3ljklqNuUofhoYI21N/obY4Jx9/teB9IF5h3tbdvNyOE7SCxxaPMWnHSSAyjGZ4w
r66mcDN+aHiVs1Hjx1g/ctulHXDEqsi7ghQ3NM8Hy3VKKfSNr57m1NZ5C4H0Kelx
qR9fPIHYNQ2TspHBmW4PClNTeHODiGA6U3WjexmQJcHuJFaOWAnXkRnyTBOclfXe
9L8DBd/RRlBCjQ6v3f/VlTkSHoozl7nNBAfdtUnkczmvEW4w3DnhLTnkOqVDLQWs
CJc2EYS5R7c6KpcW/RB8JfNnqZUQlzHd9BIt+R1FMksCLZ4u94R4JEAGE73Xq6t/
Haq0oLD1UfjfB1/GbIBftjKZiikBnmMmTEyGVwL0JVN5jEONEJVXrnFJKXugtvD6
uoWCKDC44Kav6SDrRge/NV3kaqmOfqX6t/wHxOUejc/SDvSvOgAbSNuvFXSPGM4X
ci1cRy9Sq+3e5LUGrWzJtD/E6tm03oiqNWhV62g/kgw+D3yh/RvinyCQOqviE4CV
C5IhdYinA2z1S5o4wSM1v8iAElrNYnJ1Dfp4uXwT6whF/krnmXz+yL6U0ltxI/q7
RuSjAaA4phKyqZ1Mn15L2U7TLaoSTy0pGBLDv0ZegVyrkGEOciodDZ8ZKIdBKbFg
slZFVIVHxgWpaDFVX5LJX8EGDRTBbY1asFHZ+iLBnYzv/f05QdHcWLgMMqGVnZB/
ifurmO+8YV4RwppPl7m/QVK+UC1npFFo3twxqoGgS+01hwaCnu1/ToZ1Ad4BgzDh
S0gIsxfPULaVX9RGQluOjc7DsmBN5igyVO60uFi3bfB5MZBvbcdz/5dFmAF3PpF+
B8VL3X6JtAFKVR0t+GBKeFEIebfdgzkXns0/c5EL77j7193UwIFNAubh7Qt5DI+x
GbKcTrSa6TqGPgSuOFK5O4HPIjJ4BjCnvi8Mf03uUGyKniOSXLaSB/Qq7jutny7D
82kBrzKOCaaIZu8kQ/QoTscYNEZvEq4zRddGEl4bNXQxj913obNNSu8zNUcVvwyz
7Hh/XohungzNe74T0OxgQjWW6BJVbvPjp8tflQSNsj7bCVw7XBO2seCuFEqUL9yE
mQQixTiTK+FJuRej3VQXn5K+TON/avNq1KEMTKZm+PmZ+kjtgfqfvjjdY7ViQdfu
IY5GR4uKA50A5iYzlG+CkxTyrMIZdvc5sExwcphtLagOdTK0B1++tOZ+zE9ncpD1
wdRqz9xkDTmrPqd4/akrVCZVd5kAXPwVoHgMpF24OTef6R7LakMwVrVvAjswjciO
AWGG6jLT6VGurA6v/n3fXVrBVZBq4j7EIm3BG+BFFxajpP4jVagiDTRRW8jALXCK
42QLerFalU5wJ9ge54gzHiQz3GfC1NWLzUvu1b8wOJdg2d0ktZXWolUSzxLW06c+
YTm/v/ydfZn9i18SeBWEYzbI7YpayiI6NbqbN+LKMfPeUp6dAFWvsLpYn7QHiaUx
DwIoPtSmfBpV4Fg8vu4rjOR+y3i4nLGoEOpTDN2VtYP09FCPWZoSWvPDweZ/vl96
SLa4B6KLkgKuv2In0dj6LwZYxQhgmiO9jjkBloDNzeg=
`protect END_PROTECTED
