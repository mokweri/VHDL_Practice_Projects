`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NADbbz5srUFq2xwikeJ4UV28lQDLgqsSKMSD184TfHLmNWqy4DhdTBZTvEkVqmFf
/hLRXF4DVpI95KNMId2nDjtPSMQtWu45kATx4hq8GSlXkBxbCuNQBRGXEQCvrPBJ
O5VZwVycBUNCsQ3/L2UCLdTchiyc8thhgymIVME4Zi+H1lZfeJTKYSJDbuYa6w41
Rb8oefdFCrk/YLbiB+/iaicXYWOiJUNPs2chvg1KC8jP1hUoQVYPCQvr63IekK9w
sV6PTN3VhdZ+DviOny1gRch+XArb96bokWBsmlyDyahN6aXQ0o16lGJy7NzNqCN1
uwKlcfVYJNxwsqKwJCphItWsRVaGM5+zBYTzPwMPHX/bI/zLOwQ+31K+yeepG9HB
fsBf78jH+lqzIv1DiTfLhYXktXQ5FX9RrD2+qV0l0VzlKklCIssEPBNTq4vOuvmR
B0Kue2wUaYSloNf7g7Duu7pgtgSa/+iyaDqX1e+NFTWkXxIj3NrvDGJ5TgMwb/Cn
GOibLmdnvcBLOOklTmFK5GEfCAEIOGlYdcBaxw2ITEBkDJutSpeS1jn3v5h3+SM7
L0xc3jsEX4o/KY+PbBndnQ==
`protect END_PROTECTED
