`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTLVByv+4uscxzQ6xP6QiEg7JaLnrrEm6QQ1ZeHS+l9swvka8IOlhtgPXyfhQNL3
Kr0C5YZD9+lkIGyf7jieRrfYqekYcPpaN7MmuCA8gq1dxf118bX+8N4Mzgo7rqW0
qcuxwxLHZpQpHD6BXbFUV8Tuf3ocma8ue0jk/au4U+1Hsqi47741cJxEpEBgqYaV
Gg/l+3vVWad/92hBo8WnD+eDn4OKQvGCIrRLTJD+gU4ZOmLWvhQn4jJFaDzk6bTW
sevctmZyAk6wq5QNp0YiLP9h3SX5SSApxkBj0K9qMOi7K0hao+2slPZRii8fcMr8
Z8i3tgktiMJ9xf7XF7xscpo8K/UwLzXthvhvSjC2nEmnjtPQwzggCaarJbZ1fbAQ
/xIU7zzVzMV1DEaOCltlGRkBxndrrcFptNfke34MA78A4AavA4qk2g8CikciLDHc
fAUA+CLujHOWAcz3fo1HeQLba2RFD0PhUwuvlHqbWnPEEuXsflSpzSscEZfDctQ6
brxUOUm+H7hkuqrY2t5K+JtDwjmWaZ8IWndSGVbrBZvzsllpVxPGLwX0WF5A1nPF
k9rXnl5XncwrM9dRa9R9M78Ax7ryX1C2DPZ8WDOJCn/cHoQ7ELBfm4qbjPVWP5yx
q5n0zgebUhDOYyJuKlKwFFTDOe3x7pWYiA5KhkDdOYsM06cVBPMYBTXA01JSdflL
B1N4S5IMjNNbTVzYh9IiIme/e6rU1+DqBx8Q2MkZgeb3szxX9hPa/NbhSOwq0dx0
5OSsa2j11rghyo0kagLCmpoU9zRuIX7m5OhxpZTadgo5/ZZoXN3+wnps4c4DP+mb
8exQRslGH0jdVUUcglojxxNKsR2ETykOHs9l5NxMOE0a+aivXEdrxffLtiblZqrL
+AYjOL1LPBOK/z1BO/2IrGFmRJ1ScjqgX4OtwB3DaI3GBiw2NGM+PLq9pdwf17x0
9Dqe6bzbmSrtoC65s2G+4ersReBk0bDpqZucwrbuQzSQ0ZKxBDkxvpXlNOzc4Wwd
2kAarYNZYvBc0N/NP/dB5K9d/s3PAvLmqGUNra7t0z+Pls9XeT5TsiPR5ifAqF/I
kxRKgf5sYoBcyW5Htw9A16D58B6KwqOm1SOlj0vo9B6N6/cb+fdfHmw0/E29cBxJ
YYEWfkq+TN0Kpic9m1/M4FEum6lkHu3X/38q9C4poeucWjzuXS7Lxjx8LU/n/9sJ
ADSvPdf/G8Yr6FE5mtm5nDTZQW809ZFOu38kDpCTChViPOZ0EVlI+WofwgYfNA9D
HSQbEBb//1B9SWqTH2erLHBDBRRY0Q5+mhvE/yArUZUkXMVJhTn3SJdNrJUhzUH2
IzJWBwBEWVzi4n3dZFqTilx1AZgV7hbl3WraEeCCyG/EGezLnRGhQ6gTHzxqD2xZ
hT68FmS56xvJYRDqnNKd83ziWS96OKf0e9x/5e75FyJCZw98PCzb85x7Rx/8fA1V
X264gFxILtVkRRk9avZ4q18VAMkemK3T8FGqYpAD0gPfy2GOowWvDR6af5ycBFZ/
2hijkUb4u2cRvM7ewgyZ10ZIYQJFuuMME4KQZF/2RYQYqtz0iG6yofwSJKRdZ9Dt
pxgkNXi0fo9mV2vmWLfsu0imk1rOTQsliUqeTv6BNUJ/YfLLyocxuiE825kJJU23
8YjtJUZc3EJspRCKwmF8PVxMUcY7mSkOCMl210SzYeivCU7pQ/M0ZyhiUEwCkc4B
P+nGgKY6gd+eA/+zWhyrzOWZTI+fxor53Bq8xhdyVIyTMlwDC/rUJ/2NobJJ1op7
1UOSqnLkLywHejpng98Z1rOypCBAYGgG9RmtzZ5M2pnCXVW8Fj6IQOO3lka1Lxq6
aG0MfS8GdRDB5pcBgmzJmG6MSE7rl2du6Ry34o0q0+yWLjBxMmHG6JczFldNQgQT
SQutOS2CHHhUK6vZ3dhcv3I6PVyTO6JYkHLsxnjciwLKSilFE+rO0ukxpRRDrOT1
wxdYRT3B8BGqXM0uaSp5F/LgjfeMcZZXOxtXJJWbIk3WD1Sqkin3lsm2McRi0lvH
PET8vwss4JmUmGnd/0okDcp09eXhaxFAA0peMR4tWAY0h8DucPibPZUv8d7YdJeB
1wb4bzm9xsR2PHVzr/NdYLvv4/6oXwoRT4dQcM00bwknW38vcmnMBzMj0VARHdpj
ofSXz59EGoLsZ16dkTbjosSgZi43NHGZQQnV3key3wtx6gBX8QdSwG7kTswS3s92
x+5XjWQ283u8esfCpf9fNP5QagpTtEL5PUn5KoyRcOFIxM8qfeCtwhd6iRm6oEBR
7a/Ank4ZEhFsGNj7Vdf+YS1V/rvC9TgXdFjIdj2Lfnt5vNlUA446h0m7hoGQWFJx
kNb4iTBE8fTp22CDFDxcEjWbxw/Spq4wcB2vBd7zxqBIO4rlFiv8iBZrli6+BKH7
ZYm5qTAvKUFLZFX/y7WXmozQhqULGN1UKAih3v2A+avxCyZuVuR8zET2ktHjNdHE
jub+XERrBqheAzIPL5tnX2yKLjq8+LxuBBJZbCjiER1CAumNEFd/p+3xFNz9knsq
KBSxUbpEKS+e3yjDoHm3/uJzgzsuFCqzvbwu7u/fvrhMPyGzi1R5jwqFZRF7JQ7J
QxFrX953zYtAMXQN9xbI2woulF0jlw2WtAkk523Ullw5pu5llOdpbJnRn5w4nYIY
urYWVQDTcPychwVeuYgGpVIzu9cD16Yo4Em/zLfkqeFmqFOBkcnIY6PninlHJolu
aJv3UQ5y/J+sOXSsRH96r0UqJb/ExNo85C9n1kt5p5XU1TXxVA9CFD2cSIatPJca
6VskJjjSBW/JV265lkOEF5Jo+iOGwmGtElj9+FeadHr2kzMwXuBxUX2gHp0eQVP0
jVH2dq9sHtWj091bYEKOL70tTIyEcD5crzwSRF0Xujp+S2L3zFYfZtKkos5D2ACe
18fo31oec2PxItpXeokSFYIJWrJxzWSgUG2e6BQu8aw5G7k2sXcXuf1ieg70HFRT
3MaBKfd+YCvFE3uKCnSEVnODJS6g45jnJl91/I/O13f/98kQzAOr41PsDCEQGbcN
EMekKOA2W9lGrtiHd75jXjr24M6qYnIVlEAaig1szMm1EO7bfG5+svuq1wqA6YWf
Wk6Ex+w8arUwVoWQ2SkJxIv4Qf1PWrafq7e11nvOXNo0CY4RYbl2yQACrH0SBQdp
DjI0FdL6Q6DjXyc43F7bZHqb65O7bdk3yunHsjvn14p0tbw11ElWgtTzH6tX7bcO
nR2V+m+SiHuGR0pATVNYti8R2b7hSW4ok3aBxs2smqM5q8L1AwXcRxl+qGWSlEus
QbZ7fe7RLV9GQgFXE7DAit7u9GIcP+o9mV0iEvVggl7tU7vsluudTh1zVcIJeXV8
8VU2SqhUM6F+U5WaVkKGkZfmvXNzco9xXAfI9TG9ZPHm3Rrqok9D4gZdBp6F3nOS
SZhZSdfX+6msBGy057nn2AE8INseeMi0Zu53liPXnee9nrTVSy+N4DLPlYto+V5H
IzQ4qiu5tEFnqBd/m/lT/A0lItX++JTq3KjobCa8rCFNSJVzzGpD6WwlgVNnt1t/
ivWEPzcnn0bBeYFUQwS18Xy18YVmyJLqK0tYFHtLBttwWnujQLmpHnRfhL+5cCPC
iVNVfeGDpsmCkcFUfpFF5VLqxftTsRQC37k++qoq7FOi3dFcB4IqN3juESZwHnMn
mWv4OCu1Z9QExMGyHxHUvv9h7IHdzR02glmKm0daOHWQKRLHtAX9S65KXlsAws1b
PhDCjrdLCBEiT9Zeyi0FUw1Bpi3X8G5Dd9ta7NshH1YLMMCnjcYGrP2XFuDnDwUY
1Ee0HTGqGszblm0ugTHib8pgdAhyRIFdKQLtgQjv0l3VuF0tUiux1hIgs8y2SCVF
NCu4hb34bR53fJshZZT3Om6bZg1ro6MqN2GQZg2w1i1Tx0yk/+da83rTU0qCDfPd
9/LRXAe4utpNKIDGE/j4NNxnai40bDq9q1JZ4VGuvdqIa5sJgdT3gCrNRSIvatbX
t10vGPvI7hXNj1S9+TzEl88jvQ/ZV7/bbt9fhBsuKahP9qmYp9EsliJAb4eMs192
NwR4EblI51OHQQMvVKctElG49ab2F6TaHnCjKxKksdat650EQRd/C8FUtfFm5/A0
QDNGWaV2nf2lA6ln4blpEfSy+I8W9PKv3z7LFhVPV2CKx8lPmPYREX/GoKMy49LC
jh/ENaOcQFpXUrOsF/Fc2izdtmwlsEKQHTYghM9O6hcoIuowsY0kbRz7KrRkqivf
ngiixYn3bxQzVIyijGSbIv2nCPmst6pYQ6lqJSgMTtWvaWin5e6U4KEJ8wWNdDTt
i+HmQyLYVDi9AUoONxuXuOUpGRdp+Fdcik58eXrsjWENP2B3cUphVCqAnJlGry/V
2CP2WQNf+ThB7MHyiruHkIafd3ILzgZkpubqmDD5h/eXQAp5cUM5a4bvlh2KMXxd
bGdO8hDr8S9VJ9gF3A8huMyZKLzHVYUZUcAO2GD6He7iegHlORWSrZ3Z7PlbicEE
P9PdNHfe+Dz4PwpvTWd9C+9hVh2Wfuc6S927YIRSCDLWdUOrqc4N9Fs4IcleCgqu
m9FVI2F93Sqp3VWL15rkr550SOMmx5pGTKvh/1veiC5O3pBWKcVzQXE0lpgo+V22
OLiOWPObgl51RRI3fGXuSwtrg/hI1tchCcNhvdnlVpPsgE9tD3M6XS6c96s9SIP0
tM8+0c6gMqvv9KFgHT+eF0Ko2l0TRZHEsEqi9WGX6BjReYGHOdAuohFIjAuOI7q4
P/Pi9VQmCL8KacdoGUty+viK7kUD7YOaTPn5wKruYVNfhKbMCOFzNaxMqINVEz8G
F1PeEBzJaqPcWvFQ1tbExnWKdEUXHeX1LdP0Eegi4gGeHDdPm6aG2w6MtxAPyFK4
8XLMwrlFP3OxCo82/fOQIGeWWxuywk28JgTmjn2nB2KC+lExnHxb54b1EYnCof1C
TetcjJm2JqasqFa33NkakKPy9OhMJCrK8Cfaq593LTDxUtiW4VLtCKrCyRPlUKL5
I7yeY47AnQexCEhT9oHYSWxv5IDYyq6ymNAJPaZa0DtVl21LEjgK4A/ysveBlHgo
Yo95+uAPOvZoXKOnXxxFKSCnjNlGbfSpvgduBrjbUt5mUURFOMfof0psl+//b3VX
r/K8Bto9Ofn0IE/Er6OdUPqjadZqwfAqf8J52EjKnLg5oi7IBp4IZqUwfFuWUHch
kdyfm6SAdeByADyJhDMZx33mKpYMH1IVbgGzCsWq+zHJVRlSxyBpKwPOXCHRdUTI
V2U+heefOLRDhZYcOWPrTrSG61daqHciKUeaQVU4ewbnkSRjaoZQotJ3daxieTZR
8sxT+6jMUaoOb9Rt+4OFig/g/RiiIJdBapbsQLu/I+NKvfcUoAfXEsLXbE+WM5/m
jL8xqGQ+LxleVbmlhGIHKennPX9eVcNHOIqQCEIrlVpBJlMZuXG50/jKniZbquX1
0O3GX4N4rJMOn0AbF/c8UnKJHNLDLX09NRVRVN5CfZsnKV7XzYWjgo1K/MQGuxxC
V4JGH+h5OdfqiT+Tielp5d+E/HJIRCIbZmuYj55HkoZp9bVpa/dAFHt1Zp8skYx0
ZCN+eclj0lhzvL3K4D02srg2r4E1VuXk5a0t3JSCvm2HDYDB2KjOkiqlnZmxhMKr
fkiOCZCrDQSzwt1x5kcDgrC0f1TccMUQAsoh6ZwWGikAea4KNQxLiiB15U11oYWQ
K8FVdHoPvLEiAkfKspLPJK+UCIM5+Emy1u09HQ+b1z4ah9TJthqZ2PfDNPAuqaaM
f0WhA4w2wlIzgSSzzXVZ4CHvKi/vvTyORP5tOAWYilhymQLSqCd335Ock04WU4if
JubJDUUSGlN/+RshMpPftDzkB6S/hvz/xiiCmqrXBboV0qDcjuKmR89ZnPQ8UvRI
sPdRdB8MnHBx4PGruDBAD6QRAD7naebXZHmdsiNju5fbHCQ8GIRlWFAJu+UscUwr
Me9uU3aXMQ9Y3h3GVgB+7mmYDZNFXdqzJNInz5Mo0O8Fx0L8xjDrMm00Eu+HwBe9
6MlmsyzY23WP5njqy0p6VQn/ljdkljATJZdDHdtW5E6fkP8inPZq6TxBzgK8NKQX
OqsyQBUzACxBPHjUUitQ0IHA2Xc4aSVQmI71HohiMhLvgNf5F6azKg5sNbY2wJb0
WQ24jroQ8O+3Mdb8RHU5AAmWBHg5+TKxA3zBM/N1Stcgl2eerTHVj4kT0+Po8evv
Wo8QaKWL3XvUuwVRdbGkilNeoRDsV4InCJ0IFmA6gVQBWelvPfOCw9IGIMSP0sTD
7LX3lJdEEMgNijx0CQIBd7fMawkZayvhMlKL9lK6ZpQfVAISC2vp5V4zs9c8+Gzd
N0AbcAHE8EgIXEJQdWw9Ua2nNyXaUMFjP1KxRPkuXGeXT6hg+jOf0aDk5lHLRoG9
nXdGq5te5QiMBU0uLOr2Vby5TKiaqaYEZIjUw64pKuGThZJ5QzwBnsG34IcXAw5M
PQH4JUIv57jQSIr61epEdXFCav9MtxaHqasUuG6286WmFLE0pKJ5ANGvoSi1pvIO
SLx/qdv+pt8XT8RVihqd1gQBM9rFTP9S098sG7OMh3z04MOCY6HvzrrPKH6Da4b7
MhImtHkP3RzLfKy437XhTbdJNjvKoYrLv6h1h6fVX1Ti9UrrDMaxMYjMRnTxABUL
+FrxrTTiD1AlhOVmRPs1LObLMUGE+6G50CLEdTDAVSL8kFuUg5lIcg/VYr+d8bhm
WSjqN9/nG95d16rxB93L0GawLYUZ5wQ6l4VOFaCyKcuF7VBbaktARxHax25rXzAF
1TH9cC5FrwNwbvqopxAgTVdmfwKGdNcJHeg1ZpBr5tobz9YZMR5YVXPav+qSfnfe
LGTmMmMHA16oxOcbffJvzQbAruOT4vVkbmNxJ1XE1+S17RG8p+2+IkIaRO6RVggd
qG2XDmBr/1z8D/Dap4niFQN53xZeu6EeSIq+cZHLU5HExuthmK5LXEEt5zoqRNBe
uoZfN1fiZNUOHT0ZeK3BRGb+KwXlwidP82fhpNVsHKtwfDThhvXY/JNrkkT3aATI
w8JtfaAtaGxNVvlr6dWWx9MQz873JQEZ5FNVM7T0UzzLrCwYpkQi2ryW4hm2S3gz
O5mjodiski2+vKH4+I83FFNRSwlFeYjY6yd6MlP/Hta5PHRby5Qa1XypSQ1dxfBT
ghcCzL+REWgABM5O6cfYAx9BKn6RE7b/5VIayzthmuNEWKeP7KPOkRlv+NjsQ8GX
RWG7rpXJH2uzp//8FNdGT3ojIqryaIG2YD5om7Xmzbmkh2YYcahrYa6zCXHrRIGK
m+OQz4n5lFkNK+/mG16uQhFm/ExEoxDaUjyTrb/wViZg8AwzAVgm5oXM2vbQUUYj
lMGKRiMjqIqZ3cbIE7d98Gs+5ROu+B+LeBg1P5LW+l3n0PQWML3JbDTZkVUTB161
6GIkE5zWK7CKoUAwCayhN+1J58E8q6A35BcvbAM4yZuhXF0eQS+rhxMh0KRcbelA
FZAmFN4pWYQzz5zg/vVIsChHu6xNp74QwEvapMU48chZGrGNxty5D1YDpOLwmJBt
sNV6b/miBciGnDV9LG+ltdhrKjNpMeQuL4N8QvjjL6G//WdJ2/ZbS7s3LJjtH+kr
D8Jw5jO9TljhB9G0CJdSK2jldCd3o0Zf1dEX7hkgPT4aclyXlyPg5CXvv/VYNp9f
6snFI+rAyFU5NN3NhBPxPw6+HPbdvAEkxZyxkHcBjuXtQZ51ZrCWpbDqNnQ+Gu/T
UTRDDADnTjHLrka7NrDuA9lx0ytgIYvVnLSbVKnkCreaiZ72DDvfG0b4NtvnSD8+
L09alMnoy6e597iAGXR/RHB347nlhkA012aa2vnfnM2TovW0QjxgVMa/U+dpktv+
t+QQ6doSPFIvVoaoTMxJTj2uUA/dsErDYy6lkce8tG2DCkYl1Zrqmq55OjV0cM9s
MTNO03QhEY6M2qPAhblUzb8z2Wqu8wyDoT2Hw5SSfaapRJDtKTrLANCRYUoRPooh
z672qmWrEENQgDLyYWWCgJreJad8Y4BULfoiJRnMkSxcC21dism2imxzgPFklsfM
niHTiq2dk5eTPq0KpWm8+UgjJdRSeA+An/9fQe4JGQdPcWjY8CdyLj1nc6zFc09g
GcFBbZGSS73IXFr8A9R+13X6hMSwTHbiF/sAPzDXQx1XO5PTP5/PdR1l1k13Q5f6
jsePTgztjrYhUzKWnrXgE5g9NcrUywMoToVLPILZj5MC1tPxxidpS1P6RvlmWXN5
914KpwMSO+czdBvsnZT+JIqc0Ywg3rPSEjPcPnx7DOEv5oGIec82SEatBA8/Avvg
yzpF3+prhrASFBHDJQqt7DsMUdjI82HB/ZJmJfOUQmmFhuIm1IqglBEZFy2riVNT
vYLOOx7V9MXq5K44wkNaDdRF0u9tLqeZ0saS29S7DNLkB53xIAy15LoFfDe+qgmu
MTU8hhYiyD1ZelwRINdGLnjof68FUFOa4Oil8Jox02EZTrsqNFkOYbbnJ75pQzLw
hqaeub0rR/V/iDc2IYwUQSeJLZ8yaA3S0l4jx39mMdDQBvaDCwGB+02iBRT7SZNT
er26QHwO/LkMsu/nfLYMbmUSCfmh8ct6gt42Z7qGqq9/jSpSbfV5i3+5eNKWkvoK
CgYzVKaPKei3Yy9Ob8khSCqSZPawvPe754xaHcOKzQl8zAkbarOfGUJ9gj3SkuXU
YhlTLyMS3x95/R3g2Mzhsr8qQh0JNeM5vrJRxspMgAmKl4WdsDci4fY2nUtQM90M
OWbk/wmaeB7JHIjOSX8p54ilzKkGRkNxarsF7W26Exmx006h5Ro4Qxvik4gArli/
zYL4RQxBse0CX0eaeLI2t7RPVoAxOeeLcKpQz/wNA8i+Zk1o3cWAoqzlJmsGYKkD
IWIwKKOEf4FJH74FDb4ft2G4kq1lCqho1IkWtZH0FnHBAstfAPPDfOgQ9De414B5
NKTBj9CCQ2v7qpNF+oDOpk13erj0JXOPm+9P5M1X72l3F0kr+xRFCOErxnHyxskV
62FXT3BDZYLYZC5pVn3Ct9AJDacYhwxJbrKe3u+F+x9l9tblTk6OtQUwtd7jexti
E0DmnzLdjrBfJgfcbvCd3vgQx2FJWm8TwOMzdDVWvr1P62+OInj3aVGfKQ1S5jtL
K03lB7SwUNCs91URTrAV23geR+ORETMOMuyi3iBRIIfTA2BWaUcRBgd/eDi/NptW
Mtg4SP6n7kkuKCJ5F66JS4xAiWkAKWPDIFTFIAOMP0hf1bDg/yJNNN0mOHH1Puj8
YMQKtonIAA2E+UwAMcoKo+Y3pbbTSoCpLzuKqDcANTlmsxlNfWNKob5w4QPQjC06
+7iLxWC9btUx4Gh9cBG5p2Cf2M9VWDaD/JA4JuS1dhHW/I1VOe3kAUwQEKyLbkMs
niklVvO5OwnkJuWiTX4Quj2mFz91IhynOug0fAC29MZKfuhB1HGgBXA71znAfJty
/+WqyUfkcaGEtBOq3u9/d2kmuQhhJhPQJrvVlTEff9AFPE9zWTanFdpBraSSFG70
4fBQEjZo058dpCIbfIs+2VL1/LgMHCGZSxu16M5j+i5vtItfgIGuLT+cQFMzAnQn
VTOz0BILhhP442bN6ue/7Dup8EzCmWI9BvptP+QE6Bg2oBx1gE0cPgPyoMK1nLCD
Wnhz5uVdfFmPq73tMEYmS5095YqGuyL8HQXWXRwFuoYild5BI5iZkau5uFxzExzX
FVFldZMcLId6Yihblzm0VvwBrRbHAXRMRcZOt4ioAlbxohQI6ZgBQWz29HRVZIru
sfOdkssDqS9RqjMBcbAvTm7hETSWuRz59y8ushbGAgHTkWSRXhWIX/m+KGheAyjH
kY+YoEiQqkC6XgkV2WRV/bAK82zh941M6ubXKm+djJig48XnMIzq7odkY/m0u6VC
uyE9CKGzkPwEoSkNtfgMYYKWR9q0ynOlFF3MFQl+yRPhxAUNl7kZis8s1VK+DTE0
fzuagC/gzCmJKxvk/NvulViJghYvWZK0pLMi5XKGBmgJmrbsgkMuf+DIbwbWuUqh
yPxfaIEitBAjHH/Rv+zcHX5dSSswMPJVHRLLmXPLrJsKh0O3ZKOfugS8ofE4Ec0M
Lb9n9O1TGuS0JnqMZJrPefNf01dfQQlxyCfkfehXqqBaWhfVYsyLVMBI16MpZxX4
E4+TdWuI+WKERDwGvx3NMNxud/8mJCJjJLLJgudiR/joNQejzd7sBx4zMDJGc0g9
ycbklAXNedWEr22aOG5/HylhyUS1oubrBVW5DcphQv453EAYjdYHY9ECI0tZ90uO
RUyDR3Yfmcmh1sFNpA2OcIVchUahoxhvYCAkl9u0OHLsNP8GGbuqCM44J/cW8zgy
2hIhJiuH+ywUvgBbyFV8JC4ZOq7lHXKiBC7xLQXGChCSXmpMscleNrJ3Jqz2RXhg
3zEb+AAbuGt9BMJXIwD8QECHDLR3Ha1Os0gFVQRrr6F0HWcAc4UGVrBriPtR4RAu
9NOF0qVd741hxuA22ZVQosT1NkIJK8m+/Wp/yOOLbi3rL8CLj1KWGp1win2f9yje
B+23zfI9k5WrnaWOwaAm6mAZkeX/I35fzOp4knKcKE+O+uAbbNA59ieRK3wzFxqM
BP7Zio4cUpGafHlxgIYLKuGZXY5Mwpe+PDjpR5G16zGi6SwPjubYFxA+m8qxvBmp
ST+dSC7Tw7Y33I+abuSf2Gr8+oTz6hvMIVnikINyRmOMTK7DmbdpuksBpDKDouVX
QBXXGJZnxqZVz9MUhsCkY5u0G/PQAYxHxBBUkj7OlnrnCxJsXXpopG691zkyAtT1
KSje0RRdcDnke6OqxkmzwuF4jrigxk8sZhPkaVi5iOoshqY9HvghG1XSxRFoaFfX
wThO4v7NVv9F1Z/viiMe4qJfb3YpY7mlgvIb1m3ZWUZLtYRqZhjZISHsT/w/cFlq
o+lSPfj3BjZNYKCmU157iLxkTx76gXUZya1/zwmK4B7+SrR79YIvkU089vPA2DT+
BUGEp7sMp2T0eFt1YdL0y/N1PO+D/097LqTNFNIgR1xAN5+7qOSLFqB3uaJP22WO
6+obPmH4ESSk9Nn8mCpDcbDvhiEyiqBwNtnVAX4++PoXfudsLo8veX9kHAdZjy/C
r2xMc26C5L6K2hyOl/aYDQDykTPEpfHw1zNgQvg6hE/5dlCGELjBPjD2gDjI5Ckb
cojx31jCB2u/XrlX4gzSMdgwJ6o5efXR22poSHeFZdvSL9Db2f9jZ3Bx7zgEReJm
kDr1n7cbSOSXDgWwApFFmW/VKAxdw35jFOaYcu/2t+EeYbadVSR9cG3Kkle682SM
wAus+nsoRCWWHMd5iz6Xi02GDlVKCTvGhqCC6chNAE5TIIZJHb48hs+Yw+uDsG26
Pcc4KZhAnQd2FSvkP6/H8Q0cbRpXKdQ18bd3Gp6Ek0a25GQ1e8Lma0bjG6FxqYWw
V86gHA34iZKIgxDbK47s/Kvuh8WYd83fNYsXUst69loDAMxRMUDwKQ2LwUoptAk3
WirXisjQiWM5bQN0zKhL7MElHLd25rWSLFV4/87ol0KeKtpBVJStkP6sqfLEMDkY
WtnjS4gM0XC5RY7WBN5piLmJNDdMl1cjmw8Ipms9Xm9wG5yx24wiO7m3blvtYWTV
woMDdM7XITECTUXHeBxdGYzABZHO66z3X963zDVel4Qtq3PZw6h7ayS3T40sNzlJ
wXzBn/E8gi4jsxdDYsWKWojlaygX2EUZYmqdHwDceXvKoGqq/7CXO0+wZrOV6I88
TBUj7agaNJ7LiArSQIGW7OL/f/PmWdU0C1yEWkk2Heg8HzngzYBLh7lIvMtCcwFD
+yNVx1xKLyAGnWhP6Z4rWWm5QQAOdQmuhNKWIinEwGpMHIfnR9xEgS6dpzTwWXj6
05SZJKzuD5BGLiX8lxMl+xScVQo2TfYU42LkL5yoxLFXdUnJSgKIKB9zsjQ3tXtV
X5UJ7SpY0bf5bVRQs+iBXBKDeLzjbZsdOQ4euRptkBwcWg2c8ay9EACZVsLQremG
mHCG++zNhpM6LqB68fhQIeiqGdRsFRtXWt0bG8yrvVNvR8uiGsEd5AyjCTy71qcy
GA1aGTAD7SJV+Ei7NSw+HjaI9/rXzgC92IB5f7p9Yh/zQxA8F8g/gGXq9M408WdV
ARyRixTjknue9gLSfC5x7wTvlhm/B1y9sCZZaoNBrUwdMiAIDiyYRKM4gaSLtaFR
LEZDV0KcahM70tLKkQJwqOdobvgFa4jb6b+vtD5JEspNRm05FS9Rq4JnM2tLc2mQ
VpXn7eZ0zO+AVfEeXlPJ9JmFymlh2Tx3V7o2NoF790C0zGxe9HY90rJxT87W7QeQ
r+oBZ96ptJMZkmOYXvohB1k5SmIvZ13s0gnNJ/LZeJUSOIN0bz+jJKia9GQaONLN
4V7Ytzh5PywSybPX2KaRTtnG6u4kLxSwTEnBvnZbIrdD9ouhEKMXN2NbvmCa1rYn
IUc8xEuDl+dgXfWT+W6fLfWRjH6hFSpTH3QxEzblUQ4JQqnmn5+PbLPc0SP1rGZX
+RuxtQxrmSfU22QwxSvLcF6mlVxhw47SZhTSfRZoTQtn3u854TaZ+/8rAvM7ouh0
BgpNOjJ6CkCMa+XO8eI268FbUAnUjJx8XmFyIPys+0LCaLkKDd7wvZjf6UaavJOR
t0q3bcUhZfHtJluqPLQeHp6scmTPqCWkQeZR4tjtKJ10hhE6fODXT+HzitIe/mbd
K4YjQ/kDogi9wDVAapYFamTyfBlYQpiS1AchIneleJMte6zQMv4k1BfM2F9Sc8mQ
j6pFOGvuOKrt/0r24lUxUJyVYjuXxd7wnWTtwlN63vwWM7kKuCN2kpTFSEX3dnXy
5gUqSLfLj9F9984j7QGbmp3M2CWKdm0786ikAtUjw6BymxgxHok3h8YoNJ4tXw+Z
fh1Kjd756YhPE3hhYeeQgbufBs1QVOMwhlfk+BwUkyF/H83fvHit/VxuPw6ATOjf
xRSbVCgtURwPa1Ieo4Vgx7u8bn3NGQxken2onSTUJeXZkHwhQ8QGnh17fBC5SLLb
/VJrlu3sYGG71JTuko8DhrL61+oskY8mz+x2W2A4YY5vU8RipyA4tmx5zmiEhNIn
BuZtUG2Var+rZImEzVHPKlyog2HpFB7pFWD1Uc2vFtennNFlWs2Ia0xcMDR/H+C6
cAMDK/Pp3tzYFVhbxAuTxpgwzzGQ8heif5FfRP1S2Qwgwi6uIqy+ISxdGgwJ/H9E
KVyDDy9Ntm6Sj3Zp2sYUn7angZ1rjH5dm+7bmb0erzb/Swl/EuxuytI8LlYs+Xvy
i5ZpkkN+I2DNoz/rlmVx6OLI8OHXf7fvRv0ZPC3lwXE6mjGy4sDDN6N/oxpzABPc
PBj3s2OBMcJRH8aNgnuJUTefGPkPcCr/o2vb5udp5EuYIMvDXkORsNUS75HhQz8+
Rj/Sn9CgCcVQ2wakPoSoHsgHVOMKV/VLCr3/4DytgigBaq2q2ZVPy9E58RonegFB
5miXhYcwuay40dUofjRn1viPblFdsEG/btcsXqWQoZNCQlKwWEn52CiAwNIIcLXz
ayD8rgw5RDkHb8pStg3vL9eanz2TgF+ky6CoseCUo8v5D6ElFomzA2Cd3tC4K/TR
Zqn/ZaZ9JoZHezcacFxl+g2xnNfHcmHUASOVHlzWllObA8dU13dKXTFTXcAcbDa3
r1sGBnGS8QxowL/5KxYjqmEgacbb9VwhiXcgiRGcZZh+jJcjXh+shqNDfHYPPQBP
8VlAY/d5InZcAzzVA7p7Fln68gmi/OybD2NnMUYX47zOgMoPrzQjm0cZ0vLtZRNO
neXUMBjnC171LDBxRNwvtLm2E9XNATyK7ECRWFN6o54y4EssMKV7ACW+xlO9sDPq
N2DLuu9QCbZHOvqjwAdqUoYDzty188zT3UESh8VPtn/HblB2DvnEvaI+4K3Ul5jf
fAcAz8tZJyAgNjiqmBcv+6WPtx0A6IeacGc2p4Q3Ery9wxUIky3ZlCkm3jLsGltn
TB37muDL1bKWdQX7xWgsQ+Ox34Jrrx0lbjBRlyIRVOwBhgcKEYvvaKyjhBoPOYCm
cJ2qornD4uEf9qrzd7toqC70P1W8UHEE2pzfZHcMD+htjmqbEi8YATtszgi6t1ZL
3ebQuC2jOSrKMKn9Z+ZIYj3kI/wlyJqL+Wn0Cdupln+ExNoJu41+n7yGkqWFTL2t
wbYvK1p/Zc9i4PJFsBMhNWuwjrYhbnKgs72vNIKJsJ9h1rgm7FuN+SeWWfUohzwS
SmZkNYLx6bgwaCMQBTlT2T/O83XiZ68lFU0HZzFt3MM6hmR6bExq2MBSffakjz+x
kYWXDZZsL6LNZM7veIA/oW6YUhVEdV5CBv6URRwJ7AshGgyAIfula41KrxKvss2o
4Hs+SMWl4Sgd99FZ8AJ3pPFZIYF8vpMY8Wmdn9QzN9JnZzkD/uhI2W4wkThLZIgc
hZ75p2+DSBhr1w0wuSDxIkfp2vGVuW7hOWchfkqU4PkF0FHpLw4SmNgcb8rLAknR
ph75zuRDGczVmX0dcVZVjN08PN76vTEaO8+P82HbUhZAUahjHM4m9jkeXeuF5Yu6
XAGiNwvrNw43SMW9YiG5c61jZhLvyV2weccIEImonEl6z96wmQIaWjZGlUsKOFY6
JuelYYZeid06v4EEtJnSOK2k6/yp3WvXqC7kpfV2UqwKFd/mJBNCyQpeDnwtk1xm
jZKdkCqdo1lrEzblcGYSVpZD/6DSOt79f7vQTOgi9UI9crrGI759c3py2SrUUw31
o8xb0jpyycvn0+KfWcpCXbwD+mC8c6pKbcx7PeW62XbOp3y6FD5oX8aESrQ2P13u
o1b4SvSD6/bc1EXTIK+Rx+aSktb11rIJ58w14zFGC3DPHNy/BstBfq0WIrby12fj
BAiypMswL1N6xq1dEETMN36Jqs68f+TcsKK45ehQEZuS9SJUu3UND9kuNsokBdsu
vb1WyVYxx9Gww2ZFMrm2vJZpDxZ4afxGiOj8NpVqioJ1SPjxvZisWLNtLQOVbhow
VabYykaV2nQ0EFOsVO4Bgw+nQ5yw3siMe7rFjhGvQptAyEP6ZQ099VKeOpp0Ctem
QoZMo1Rn420OKnYhZ2R498bVNu+kAldIDfpa67dM1TzbGWqLL5JDnkj64F2X/JcX
sa0ZJ5tmFljVIzUYvVbYtukMelpuvQWW6Sb2Xe4llT1i//xxXoNYMpWs5ldWLofP
9ogLFK8bnYnGSoBzgapc27oZXXl0TLFA9k78Jr1bbsJ53xfyyHEVk/KAnKdVxmo5
XkoqHbaLslhtocjgigZo9PteYqeLiso2XIcdwmzpe2eamRgAyCLUtI1Zikt0MCii
CGYofZv0POGq0diCUkKk3uh6Xdn2+sEY1jf1+NwWbWcr1+PGs3e2DqEPRVikVArZ
CMPEEKTSj5+GzhREcTI8Q8woXAGz/YkBScqaSkjLPILM6cVdbEp2i08QYReEWg2n
1E25zWSXmgu7Wj81TVOiBLyi0OSRihj7hbxnmD86mGo8oEXzX98M2dBSwwUGGKE+
yjOnizKsF4VhaQizHduKcFey3eGYyiDi/8ukDsdWDLjf9xsjQ6EiEujofwHvjYe8
1Au4xz4tyyxuEXAIkQ+LcKorau8pe1zBLEWufNiZbqUy8ovA7jEO/QGZmOatC7RV
xkiDE7WkCPSGqlZ1OGaKqTqeNlngaF8u66IOxzQfEuf33gFtquVCsy0uRONHy9qo
XxYgJ0QmvBjiBvPiTYKPSbcoPlmcDRGFxYQJYiTC0W2k3WCe2f0JQaR0Ac8BDv6Z
6aiz0UiPm5cWu6IRdCTO3JYCV2FatKEAnOURN6bAk+FJM0lBeKVW4gC7Qo/hbqk0
K6PNlRqeBB3hxQj0XWSmrX6s9/8FCfMHs6w/m4ktp7ypVLLIxQshWLh1hMbvm+/L
1HvPSEL2b/IGloTsuMnsKK9AgrKhRCOPS7in/PePmEB2WBrgweXyzoh/xWGzYr6U
U47B+LNAowricx7jY2tUPXhYo7E2AmD8RUt0Kn2sVrNattLtb9PivinfXlJR2Ik8
AwvHs9MlF6jCgVayIEH1h75KyWRO2n5B7lQHplrJJgKj4NazjRxg9UwGx1bcJ77o
aT+Z9MZ6L0rCRwCOrzsMVNlgONYnrOQHCZ+iUyW/iHXAz95GmiKyNWRO7eWyARhp
qTRI76wG5qsk1J9BzFTBA0muazA13isY909Q5LzI0gYNctxy6Qg9qAeGHljCPNa9
bcHz9HjPuEkVvrpGuxyCPkx56sZhMS1ckmRKwj9XlDigUkzqTTHXIUB0Un9q3nXx
D1aI6jWPs5V/EEJfIjeJHoITwuac1bWMz6Ap0P5d3735PlqpBr8Ah5uIFdWX1dTY
+buCiawKL40+nmXOY8wDb/TFkMGPU74uVYA53ar0kqs1h4S6pR9+5Rz/p+ktru++
v+0AZ8dF5DpMV3v3C6UrvQf9kjeBVbwMQ0UK9/2FZIINVvV9OEFGTiEq/FwAk0Wv
4g07yBbajwD2JJJtKtOr67E6HSfY/GJaKeKEl0k8oE5Vh+C1lr6sf7VOCkDgN2lR
aJs0Lj71a/PyQmhhjVT84ZhiTAYUvthMu78+onJCmmW7ZKPW9hUsjSHmcRGbLDCI
TEmSNv54TynF3kUbsdeIO0IMLIYZNWNhDwtdA8N/QS9S+X1B4WMCva4KsW3MZGri
O37DxfXvDzAW7cU91xXwLmZeozKVMO44i3bX+zAbh/wSPtdDvLRYQy35BaWipk5t
BWgc2uIFdPGQdh/vYkjYCVuNnVE0k34KzMUf5dgmNpXw607PgU1woHmb3dIX7Oq9
6ezi+dldGCrdj1fOGgA+d8h8rnbcM3WctKLmqzULmyBrX+MwbKAdEIo1j0N0p7Mp
GDaD8xgi26QelNAbQJ8eOhONLbfTX3CC1+JGvaF/++i2kijW90UG6lsNtU3H7cKB
uFP/UlrWIX7GT+gpSQpE71zV6a9jlWH+Ft2dDN1L+YOBKgvSCD58T/SJxXBomoDY
HhA5OdusmcX/HVlSuYEl7kQoWNhUSIGj16Ztp/hix+xvPjEQvIjqF+/8bs/EDzRp
DSVto0Fo9vjOi2uPsEK6mMfLQeC6BXxQwZw8gGv3pXrBy4+kXcIS/xyNHOWjOYTi
OiPg+OqH+XV4OVDQOK2tSNO5P3EgeE1//I5ZgVXxWPvOYLeN7VnIPv1nImGTOjo5
jNZPeSQ74P1xuoEKb9+6nYQpx+oE9kThvokiCta2ZybGxjWwNcC6x6jCzwosJt8+
O8jNgc71wjaMLm4hzwiu4sQc8sgu69IrHoxg55bK2mKtMIHpZe5/Xz+jdk/3gvqE
xfKR9/tg9gRlE6BUOIyfQZu7UJzFLsH4B8Q1dyNbOaMuriAE4zLKEidZXZvAE4sy
hyJVH7oJmi02BSR9dap/Rbmj/cwyk7RBtWchaT3YW2i9/cw2Jj/lcd1Zk60W3usT
TjsapipkOQl2wvnFJSg+5bT1v+MSmqQklgangY8ZUblrL6TLRaIHUthO9+r4X0BZ
EQHHkYu8aAccobZOx0LJbeZzUDhjes4gBIoe7MnZUOX9Ev25wws/cqLylrtVmO2T
7rXRu2yBUl0TpTc5sO5e52ay1JoeMiM7nNcdnWB3jQ7tm0N+27ncU5HfHrcW9SGU
/GN6z4XeqJdhVPuvsd92wpTkPnsi5LhxiSuctnr2H6pcIJX5LUrRVo0VKfc8f7r6
u7VlRtx5rjge5IRuqVGloKWcCphKIySCx2+KJA/AWLoUTRthgYo/8ern8rOwYck4
x5YsHK7808jbEjw48z22KsDRgPVBSU5Qt7Js3Gv4s/GLZhpSXy8wYkiYchDPKzrh
9OHj9yVfOa2txGkA4eBILqasveHqFKLC9fXOBTwjsDu3cOizvKh9XS5q8SUJzHDO
nINHH/n4Axc+8OPCQ0egWXhjKQDGIc5YhejPY15lXXOeoUOOP9p7hqQ0vIur/r5w
4oMMEd07XpRXYZ82qxtxIh1ujUWnBuatwv2s6TToYbTJBqwLJVjW2zkmK2VM+8DE
FqZ+DckVKqlre+tvIgDwYoLYj8gIMNVU6S/wKPKFZBHcfuPH5IspNMmMuRsPUqC0
vHoDBE+taQCAvCu3dDNu1MUQqwH+fPmEIyj9MMJU0tQHDv+36tS6EHBjLmKVT1zP
QIc9OcPrS8eiTYAcsM3sNSuqlyHOAcZfXS1UVV2RsWrjXf4/UPSsb6SgvnfZFUZO
1x2ValelbvlCuxecmLjEs9SUMUUp5A5csdxLnXJd5gE3GJT5eGlGiwtBidfaxhfY
Ydo0eiPWr6hgJgu5JNA/iK7EG3Q/4aDcOTSyM121tybXi9c7JYc1VZ1/t807hKSq
ydJvl0K+CftnW3CdGgm9vK8ob8q6+5i7li/C/nBLeDeScAQWDsRPVTAwql7C7Lj7
Da8HIy5x4YgzX+fkKEhhki9vCQLeMUcuM64ejPmomltdJwlyFNXl6zZYPLHcYe+i
bkW/FWNb4RhMJvwyA/qL1q1qWJtWY38KaGoNZmvnBnqN4YNTAMIBSS3v2mqUk03S
wTFHydRc1DJCo3tNXrBxTyU5pSgoGcXs6/P5lHv1MAdtG0KwyjAyD7F8uDajVgks
RPG+VL8YbHNbCAJynTXs0Kw1Ygj0U0KSQxYnb+uwiggm6n3Yv4rI57r4ZsBYCVW2
8+u44eI/LZYOjZ0cs33dUzxUwDE/FBqP+kLBUwz/x8wE2o9BA0SuM1WmVQufLB6x
jX7turrOTzu79j0oRY/9q01LUTkBMXbqcpcybQOaieRvQ8TnQ0lJdFgBRXx1TFGI
WdbPy9TPVleExr5EqjgYtvjiRSh2bLmQd6alq4jzzwh86ln1Rt0R/q0wFwKqnZq0
bzEMKz7RukEPFLxsRsxHlGbQBfDVeKpzbPoBn+DiPWgB0Ql3g29OJxVDtBCnK1Jj
+xnCnFjf9oLtt6btSD4ey1eeZrwcT8+yLL+b2O3HBaQeBWI4tD/03FhFdj8dhdnQ
0QXjaFOwUP9QxwEifjCiMAlfcNa3/NBp3PKyRR+bF35x2hcKndAcoLJQB7bA6EJX
8MqSUcVjbcp9qTe10T8E84NWA0Peft/ru6PGJoW/uDFx/M8hYIiRZove8zq7zW40
tIyNEnG3Lq0kPfp2mN4S1Yai98q3jLxDmWPSFGMpuYcuwT4tYZGuous8VFWo0RoR
9aEP0xv3huKEcIkw6jZqxvNwQFu6TXxz0BHFe67wzyAc3iVXuPjKhYkQOFMXrj9a
6N9Nc8Je9p9wsAvSyMzYETwvQMDV90LhfFdVTOH6VTZZ5TIYIpY2HxywB4BgcfIh
cu6BXaJ4ipy6sdUSQTw/O5utvef6UH+xM2X7ft6EGpZUdnbhxpjovJen5bT3Nqmd
fqFpAWzx3x/b8te+VoZG9lg0tIjer/gyLvREfmvQRVStSV+6pQow4hA92RFSZER9
YGpOtBVDUlNFKIhe8kyL3IkD425eXoRZHXQ/SrYriSZSJ3UN1PX7RkQXaTJclmjY
8xo3jM+fgxzDDBfSLp5SQdFMMhrisY1qAOE0QK4aYNIlsfzl3f7vcNvZYUM0ZYox
EXxv62ptssYBw9OefcNKGJFaeY1r5ckCJUIdo2XoK2YUBymGrgfL1MYQ4JHtn76d
y+/3cKTBGBswqogNjqLKxF8tSuEtxWhVQ/lVeMjdvETAW5Gbf9THADmGVWFC2P/h
leienIO6x+NmG17sQLsfFxF6us6YdQRzrd0YwMi1F3XxDH6U945SRLgE6fOrLZIg
vxXzAD7K/euqaAUZshFH2ryFSG3fVUz6YIpvVl/8uTtO2MGudrq0rddrYj43ZkoW
CbV9f79jSDjfHuSI78NJ3pEZhm+XjB67SaeG9DoxFU7h+iHMCEIDEpYpnwf8C4ok
TazD2d291XpalPYb5lwONIRT0R3m7Vty0nBq4lmO1GO9ZvyGhXGwIoO2NW0tyP6P
wKOb9DvvO8MBy7/to8O/P52RU7X+LuTcq+MfSR8HRjsGvco6PZwroddF7ZTR1yl5
+hATvhSZoNSR60x6DEmuyzkOatrg1F6W4w87TIcL/Y0TzImbtbLK0BDZfRBfk4RW
+oy1egSvx1g68CIsSpNvGo0VarF14vxG6fjyy5KkUrxLxSPbXQk43u9wEG5gBUIs
49Ri2dL9o7mjgtqqRawF8CFm3BfO0fnQwsZbTPG7C11wRIdyLz7xD0Vr8c0RZTGk
m7HOEqwFxO5T7FNUQ0YysDdebb+o6LjSwjZ1LpnhJLqeXbyTsr4xzY8UYoNBkRM6
tvFhK3O5Nj3eLJEKSQx5XwlZFfCneIRlWlkEV9xi75738v6ukDM7tjWNvX85C37y
Y06A9WuaCijxssNebQd9d4jPaJS0xZRef/PZJ5dWTsOz95ohtebOw2PY8+2J8dOv
w6HGAOMxz/O6RoZjInN1KSbRIIDh0Iu+1ZZkgtlX4RaqZDKWNxhYuDIl5YBN7MLF
fWh6uFmW48+IuyPHiiLzaE2KvuwLv1zntkaj2BdX48qPQkLgpR8o21bVqU4HdTVa
5ukTEdKNYo9LAAzyg5HC07YNoS+B6kOFmta36DhBZWqY+LEw0kYK8iuaepfPwZrk
7G326iy3Gpg2WTVSwaGRSi6IHGWjh4ddkbIwIGQDrD2vp1w+GtjkKNnG0VLneOiE
cyIVpQf3BgHMRplj5U/tBfMe6U15Y3Ds6G0rRxs9eWLA+AL8DacVddG3IMPRiE2G
8s0EJI1/zMHS3C3tzUPn3xhQGl3gvOtICKKMbgpFhWSUxnE0E8HrBaeoAKfENJFv
xFYZAEw82QHguZvq429ZbEwPknf5trib7X1SoohwIqSfRaPmsVhi2h9s6SEEUK7H
1jm48bTDFP8oaigThJkDpydXyLX6pB/Y0uYfB4bsNXicbPsSWuiLxXWB8LnlV6gb
gvssnr7C1LWYqErRUM5xuqMRZANHwMepd4hKlfZqtMeJjDKfI6QLdv3WWs1z8pzB
NwTLzUKOubrRNQyTPG2MdWa2ujdNYfp8i+It1unbVRMzVAJPqIa3tuNlizEQnv44
bhF/GxpwzhwcCvwKp3+PYF1JcUkQ8JiaYeKnRuYGQ+hKG0Vf1Ky6qC+Jcae/HKUW
K7lTTCXZtD4w1DHqE2Agk4Pu1wYwcPe3ILwV3oSLluJx1v31C7TdjX6QcQyQJ8DS
NJ1atnHke/usbKKWPYLF1impTWkRTPzz1RuI9eV1Sr7ZkAhNuZiWQrxnaYul0ylW
FHvJ4LnB5MPyxjyZfGyZyJPpPWo4JanLfH1ZAZGzmUr4/3Qqz4wQuKiQ0KChtxNL
oA1YOFTdv3ymPZzzNI+tqgGzqbQx1odVuCGsYUp44PfGnDXXeWE2gQbLSDGjoEwI
FmlqfBNEt/Q7xtobZ3vKks15JTYiWXTeWwMABsqE/sluMR3XQl2AMjWLaPvgzu7E
kE3clwtugmGLrhhzM4zFZQ6Cqogw19Vt8ie+iMumuJoK2iyiSdiWlT8zn9Eiwq5X
wmZ9F3NItfrGEFX+NF9g8NPD0ZcnfSVN7fq4ZeW5sMNYpcyc88Bg1Jzf5KAe6PA7
76SulhOSvPRlsSCI8IYcxzcjPezzZjSawgBRNZCVsRjpOSL/etSjifPxv6Z35yNh
42Q+AV1T+z0nadCl5p+rbubgnok0SdbDXs1SXosTaKtMsKmD9SyxUjbXbqNLjEyB
uYJq3YD1rExo8S3fTXPlKV69G66JTXLu5neHUVQXfjcKJevDTd/i+nm3FGCnxNuU
Rv0yYxe3kgs45HeE+0XX94L0BbgDFCsbLpMK4YifS/GCti915tH/0+jKiaCSEuTO
ZJ6+A2X0XNX//fR3Cu9s6rk2/+98flBTqG8BSodF71MSeFwgruv76ewJ8nsMrJth
0PCRncmTOVW8m/4rQnyGtCTsGo4j1tcewE6RS7TmAV02sE8Q4nPPNV+gXaq0bvxy
aw7V87/T1pgRh8oEZGhNObAochn6BNQhqklVu5oYZBngyfEWP8+Pwij/UchMzHke
nuabEF60S2lN+fhqMMrZ6HMU+jqN3M5DtgnxYQ+NATE2Xb/37pKbaVeefN/8Z+HZ
iZOv11Z5cII19tfAxMutjwbKDC6fGZgFXkljdEVmIjmsPVnp8mF8+F8U4L3F1ePB
s1PiFXKfwBsWr3l7IK3jP0H5Sb0GPLsth67kBcooH5jxd/Bn6fYO8r/I1dWhOo/H
pq6GEYMM1qDDFqRParTXwAtKRkBEdDvEw99tMRW94qyzLEEeRp0EeotH/P0GA5+p
TRqLhVJk4up/Xf7yB6bpx3Sm+hSaMjA4Kn3Ee0xCS+cL7K/l2oCNUVp2YkACma5S
InQ+LfYnkMvrENz+Eg6JLNHYY+d9WrDlrtMcr42w4KrrbULX2Ag7aP1yoqnc4aut
K09M4kiRmv2kFlpjeHB1mXHG1pRxSGdt8JpKXKJM3F5/zjmoIEyJ6yv6ek0XTcgJ
GDZGBUfL5V7mEYEy37oPwsZBb9sJBWsnkUvJu1IeFhAGq37Kom9ZmRwjdpXBcZQv
iCfUReyACL9zMVKet9mZbKHddprRyel52+mty0VEmTOnyOOggSgpqq1Jrnul1S2N
IA2LsWooE2C0jebXQY6H//yGO/n6QA9rAOxD5cLHm1u6HcEPn/Jw7q1jiFot4v9u
a3ObrNHIMXL8BhfNL711zMfDQXwG2JmPfiVUpiAcvI3tLLhbXdJ70sTNMpKUu3OC
bWIv9HCcLrkqRO6YPWiHnywF07CbgLXPJ9SgdCjOUwCB0OJOlbiejfXmqjlwa6tj
kYEKMbGA1mc3vvL2lZSsjxj82/iyaf7bdvGjqt91lAWH+Imqq4dpTNTGQFt00XhZ
45cqjcz0qeQZIcB9ldnyDixBcZCROHWym+Nr8Sx8ooZ7eIPYZIhalO/2hk+Jw7QZ
QLD01IqjaXM3bDbvLEAlauBWeHwrSL187fNDCR6al4U6M2q4cryOenS2aRNk1qrM
244wMwK/8BpTYGEBrlwhV6IyVEWzdfL0rqU0vZmgokHOOUnSydqCmymmUWihWGmS
ddemRoNf0seXXUuIizqVTI9Io6g+s7v+U6KnrqeRxfSP/r3kQKfcY9eqnTfQRm2G
DmrTuigea/MF6oVZJx8nTvhvnrFRbRqsh0AExmwu0nIVuVWG759ZUDp7v6+ey7Iz
0mO0QJSX97mfiaHe3yC8wnMKEWnPld7F8xGCNf6yz80x84+BekhWquDkP8XYINmQ
NiNvbj/mSOd3cPThYF7ED+t0+ubcloD8FIShNIvA0ILTty9i4Ckm3UcMuXHEbFoE
FYoH600ZSszD8wwqTU269Oim/T2RScBCybOuLfHxoNn044vZ9R+OYo6+GmV+y5pb
8zKaZBazGcTez5+OM5/sWov6+12HLiM87SvwJa0+UrRe1oMop8xsIcewRY0xvoRA
2KH41neUrnvTy0hlHLX3dvPuM6xjDytLQNQGHcfy9m2jFACTkX8tFcj6EB8IlZRn
nmBFG1L5hIy3tvYIS7fuZNOYy7Fh+w9KaSyFttGbzSfVdiu1QHcTPLlyvboMdXTA
3WgNe45gyFl70V+9FXyY+WjqpS0Bhd8MWItMFTmfFdg4HjKutqe/pNJth1SZgiO4
XSFMpZUPX5dtlGihrMltFE4L0K4vEcqiziBuEs3MadDTeKTWAsBPr3TcOJgNMCyq
GosDfd0bZhfg8rWrhD/Wz0st5gdV5uX28X81vMh1jiT/4IsQPk8sz91v+McND+Nx
KTbz/Vy0HDb51y63Jax3S5mGNjkNjCfyViphMibsXotvKu9dInTvtAn87EIspOZ7
AA8nHT2/PNGntkkgKOsiRUEJhaHT7wg0+D9hiakERLFTH9QeIiCyXK33HlDgd1/P
W6BRV37ExIjdpdwyf+CLHJb1IoH213nAL/bawb3UU57cqVd7EomTP0r+18mZh8OJ
z+DJPPOcQzPMs6zetFCMGk+D7rgumXWvigxDjAl71nffKJizYXZCW2ZbRzBBcFQU
/U9Mkyk6SVReoL/xDSc8TfQNtxCOKqJP6QvJfE+x+iS3xbmk/wN57F/gqhr74/+n
ZDTTu3KJ9j7szZ171+aZVRCZFCC15OLmm2cYKtz1Cfo15uJuxGjALYHnqUCOgIiX
pbhGrxWaOKIqTKoiSc1ss4oVSLbmdRrERoNV7kMBhjksCwKO03j68bqyiBBiPQhr
SP8WreV4NvS1LulnjypBV19kh2p2I9Czg69pPJg+qlGS/tYmtPBEf0LDxMEPPf6r
GL+G1OnsnxwdBCAmqCyQ+gwm+M+GHKor3Wo43j+fm9Z6eBhhrqW0xRzjNijEKs1E
M4UnfamoELIZPIufCHNXd89xMeTjVEmrhGNiUXNjUa3SuZwAFFUZ0drtj1XcGdHj
joGXPFFIBWbZmDiCsl33S06nIo6KCAkqpVo8XPmW3GaDv2uO7g6mkeLbQXyowTeJ
LegJoeuY/jfWfrMvH0rjMek4WcE0shnORpvV08S7PjzrIMWq0DgZSrWBwI2ZhJvd
vpV9/iuGf0/N0lKTjqAKwvtx7KVUvdmS5mxsSLJkCHg+y1G6VPs966FnlA2VLccc
oxWPpJe9rjzC5qG3gytMTlR70nIyfFG+NJ2xaZlw56aRKhh874Plczy+dOfQmtao
6QRTmWhlmUe1w0itszlFDPqCFaoKAY/n20pdAZZUvGbmLVa7G8kiy6SuuLnkRT/D
m04ndekCXROgDm4odb8UV0VCbiRbE8RSCgWlF07Xp8SsNQ2amOzwGH+5VQCt+1HJ
B+/pJxjccj74KLYP48QuYvNaCdjPxeymhD4oXBwWpKp7DczhS5SDSulPrwEbfqSJ
uQlFO6qVMvTCp5dt8w42lqAlQcgOhLnufm4jq3WE5nd0uikqfZ8iZfVkGlPk1tMs
F9NHCjwfyj/lxxxz/Z/hEOMQcOmh0cV954mdggUTEcn060E60ZDMLtWfevf49DhE
koXIdN2G6dxHgAUGkzuuT6tPyDpkWFQrPM36j4Na4llxm3vSNuCan3L9FN8/viUb
klGyVtQOvNTiaw1tB60xXtNJzZO2+Jc05OuvtvXdfVzBur8cnCOByWf1Rg1aOW5S
BaqSlSZVcXxr4nToqEMlKZKxN08n0VF6qBRylWX0YPm0oQYz3tRDq0aJv/sPdCCq
iliPY3YGH0ENepx9Bmt+Wm/aLiDMhP4jkScHZ1rUXAoJtm5EKG0XF33tQqzNePFH
+wi9oQ8zalEEUSKufQSk8Znb2sS/Oy7PtEPW82xYsqqfMf+HyQedoDKOI97vGyVv
Y+3wG/2ZxyQSryRS2gmUfTjxC2/vM0arwnLfQJL7QBAPIBXWdW1/E7kFIjgbL0YW
/C1AU1pqnHm3Ex9n3LCdTzRYwBUdq8F6+g1blPd4soEVilz6lQ7M4LJsEjdnHoIq
0J7aCODT/mGat5SXhJMdJ5EvAzRIS0VPpzL//gL3UkcHBWWZYTZHnaP5X2XoFIOq
l6z+M4QpqxOdDOlBeqjNLQKmMgyKoKj8FXVOHTbMc0XZKN26lbUM/xJ5WeOgYQBU
kTHpa+IWThjGgEfNzp8vtIkaybeVCkSZ3v6u4TmEeUkblPUs6AYtsAUOUqrTw0kO
ZWsGNn0qRP/7wgqK6Gdj2BqfisaQmteM4nMDmA9P0RKH53KIneNr7d5Z362Tif+1
18rzJMOS5jQn1R/MifieQrHfJasOjMtDFC+LfaN2sxyGe2a0sAVs6kCUg+8u2bsg
qXC/wnBvzkd8DdUPT8+YKoai5Skc66COxvU5ywZ1O0wzk0ewSxkGRDUXm+RVkoIt
5jCTHH3UQTJdCoj8LZZ5KfuBr7phU8eGRSNqFjWKfwlVxrBHEp8sNpi5Ib3iVo0G
ZFIRULrY4g3loTO7izjreuuelLDcV2uroK5DFhP9k9ICrTbmueGFx9ji3x59zLlo
XJKNi1mD41RnNtpqNGGxAEbu7dQaTkcJrBG5ce9fmVjUhQ1tfICeHpd0zF1tRI4a
lbuu6uH0RlHO5EURpStf3+XzPogTr1PHLSixVSbQH/InlBEZJDZD/B24mgpl1QMq
sgd9UR+grljDygeMXQsTmQ+DTJmYadBVqsDfVPxw4DO1TmIpdj+9HsgApMi+Q65f
vSMMRKLbAeZMqudpmCUmHCZcdNypSw45Qv71Uj7ejMfJ62fcsgUr2MXIGCwhAUu2
nxwMxPu1EO9ZQT/gypxQBO9M6oCG7DHRzUnIXc/SvCeqggpNe4t1wRNSEfaMoIV7
T/AHu+eMXs5wGy1vfXnJtyHyRw2fERdCujFWiISZA345ZM3FcZ51fV0SVmQRWBJ5
iImFxenG4+8B3blbC9VIRa1wehdaZAlQummTx7t5aVTMIlQJxmEgTk2fB+AJg1aO
46hh9ToF/8dOCKkNeQnrz95xQVWlVpuU/nkA27eqcmfzT38WPkZ9zM8y/BliFYCq
Hc1CreAxaEUcwBNZeCMfvTO+ErVMAEFPHhxu4vWPRz2KmusOW6JwhizhYePA1Z/i
LUDc6N2ySdUXnYgzeD5bPSbSAD3tfkTYizaF0LI9l4E8rrqu9X3aEoK8JSH20jjj
j5QZiQuPE93lLv+6WBBYdK3uT6wlyzOUOrysYj5SqVzgMQzMlJctIip6ZtTRssQA
O8oc/Tl0MUQjxN8oiGQdV89yEbA6Xw1xwqv/sS/8BdiMdeBq934fMrgCPMKCHA8/
NKdWoAc0QYecXUuxwJolLkZlo0IVHlDUOXWXPV8Adm0C7++isi2kd3fGb5PS58is
+2ACWlfhGsCjnQ160DBCM2mnWe7leo/cz5wXCiqXQ8+vhlSVTQgvHPnqZV9MYDoc
r1QmxwlNWrvsO9s6mgorpb+NI6AIusubte59ikkvF+TjbsttH2OZz4Qiy6Fhgzxz
NTyETdaVXwoLnQ1H74AyDpg18Gc5jIIa3jlS+TADXAhR6RCeG4qtBXKsy1/JNKHz
e5qTZonLGQfypwdBw5BHP96JoMYj7+s+AcrXS3BJJ1jf3z58M0spVjEJeNM4Jft0
8TX69K/11abG8dfDTV4YGdrwzlcmLhgjZRKYpkglZlmA5/hyafb8XxxhZh0d5vLk
iGKLuEAA1QnsmQ+7iUlIx8yXUC5f0Z8fD1d8eZ4CidblmoRjxD+2LS+EUixiMja6
AUAJzpGOzAWwsSHetvzvxA0Ydm4291qUAkQen1RDGc+92AzQ+LLoYc1L3YpHKHYd
URGeRTAUGbJhkuCzUDZBMEHU6+1atRnkmF+j/J7eAacrm/mH1TxbHIzqLbYthYD/
GUz0VA0pGtStBwurGIYppQvYCgKIg4xpqUX6236FSW2PXqIymhySFUeDu+yKLodh
iD682rUgQEEAAUByOZGDSPp4kg8vDpZJANIUnYw8JU6ZRn8zEytdG3SOaBtaPVoH
HMFbV353FL16p9nFTPqsnOEyd2FlvlH1r7sEMbrVWYwm12qU3HTpsP9C6Gx3SBZb
aRPIwJKPZkDvMc2qpyYeS3srcypE2PE+nLHcnAOvl7SmX3Y5cjh2YNXiYnBCEoTK
hISZrPW0x0BEI83Q3LXIyVLOUKU1YPMgFS2gJC/Zue4aB6oVnTkXQEllEBzHnsjq
OwCghzd8U62+hFRV8Tj7Pe03sf3KEpiEuPfPK10oJ6aOHJDNiINljMYIfvLcTWMa
gIdVBT/bBjI3/aDvnmMZk5Er/f6Lfj5oLhtlU47zRLXXkpAOUXSRnG4mRZEIwn+m
HRObbZDMUkFIjOolbAXMhGsZVFfjSi+cgUyBbSfmM8J2z+VFcwoLF14WKwzFFLRs
Q6uDAM8LIBAZ4a8suL1+b11v617p89GYaQoMXZVBw+5QcjMzBuERPXNbp5poPt4D
9g5bYXb2lI4YQU7T/KdfC0P3BjcRAiLG074/02J2OkEcrQCuQYI7IwVm8gi1a+6o
EW4iULjzLSI6Ah2SIL7oIEk5ZCHCCedRVxHjvmKMyfW1BRmY0T5/mBSBnBg7wys+
6a10WyyTJPcJcjbVP915J7d9lHkVVuTdswqRR3uMNRsmGIzYpNK+x4PrN8Rj/2FA
/dQYi192SG7GpNnqR1UoCPMqN5m7ykLYWa0JRWEPbJswy73ksUhoqaed+eXGIZEM
2dabMbSBay47UaMgTANuW7k0wCpk4qI3YzL2z7wCVkicX3K1ENEE4/FF7ji8ymip
+NpI2vvPFMRCGyJJbpDFh5GU8CeekRQZUa5IGPBA2a1T61EFXd69HToi4sZGWOaw
3ioGsVH23uvHRkqC5TDOEAiF0ZNUyG9M41Q3xpi2vwfs8oANj5O5dJ1Ndah3WZoB
MK1Xgrx8zaocNDNMcDqzmQeKQnM3qZtCZAhCf/Px13ohG8kvfusGf0RTLwGcS8rq
rhNnu5sRYs9rejhc6fANkh4Ib+7oj9VtWna2sFhGNXkB08n/q8efS4U5KUz7X7Y9
HHUhn4mg9zHJXND/KYKEo9qHrhBs3mg+NYLWjH4i62kr4iuiUkVhkbO0Y7jl5p7j
org0GEzF4U2Ot0R4qDj11j+fmk4PEF0dxgmpTbLyFI0YmFE+YFb727ekhyJ95wjF
d+daACiMZuU2Wth8BqeUEt+t8ownZkANXCFq3avrKk2W48z2wTyCTfP2/3R9yki6
RjYDV8sYIa+C+v+kXIDI2PDxfR5GwsvLGREd7Sj8rxYCyeocFwnYsolFzOqWgcI1
taeH2J25aq2JV0jFXHNcVSP8WoIitdDLK759FFzQecfD+ikavILJmsQ4ZQnWSMrA
edQE/1OOtrcq5Cbjl0OzcT+1KW7hUgiqMOmFFxTW6RZOXWtYsrul+LCKi0NBaLhI
bStzbj8z8bLkMRojNlcBIsTvLqUrqir1vLONRDUG7/V1H/TPaSC/VfG+FumCrCu9
FjP6xTSGTVatbc7u/Wlhr/H7uWXQ4CX4AApxVZLUJe3Ht1U3pgq5v4Rx8vpzcVz7
nftWrUXOoNTgjXyZL1Hn86sKZqFfXxuZBD6IQut/D8Q5uLT2AyVUlXmQADzhTOPa
k0lSkJAPayucTN6tXDcTGaXa/c5zAhTdhmyKLYWOnTv8/6mFzIsR+0yOUsE0hMWC
8Y5a9Ek35522c/rGRXqf3w0eZu83fqViqKyUfIFThoq+k01QzE8JCsIm+3dg3EaG
hHNYmu76k6pQD5ZKJaYLVLQe7RHSTuI7pjiBPUr7UnkHbwAFrO673VOLfP3PIJmj
g6VOCBa2fdAn15tkfYUwLJc65UNYia5ZZvqvt5c4b82rLebvMEC1OwVfx7ypdRud
yReV1Yavo7eJ2y+XRFtuggVdEbsG7KRM9ZVNhfsEoHqNdW1xead2A4or4DMa2x4Z
Vh6AWd3ZHqCplyZPJ5VFsFygeL/uGBxcGo1h8FNa9q20IRcq9rO/m6OnyKzc1Cm0
Irjfe82+hYCaGvkDE+UhFRLQTtJLpq25C6CJBSiKjv+p6g58s7JnCBQ/Fg5vt+It
vHFtJFUxERrFfAFR8SOTPrvBz4WDsDsL4dExrUnZF8BumjZicgmYMx/80+Y1KWJl
t7nqwkySpZkr09sAYnHxcMp7mv/55vkA5WdAOdsqx5B2MnSHGiheUpD0M08biv8n
rHKHO9IncP2nyA2ttny3XEsf0XKxvzwNu9HOfAF56ls1OVCFHuu7/42vs/47XO+U
1kOTLJyigvoQ4Ptuomdwcmd7Tr/REbaNcQyZJlnEnq0nMUGbQeYWsbfc2M6cKS79
O4CNVVaoY/dE1dUvKC3sYiSbYqw+g8fL7w6Oz9BQGF4uJBbze9PZRE2bC8M9L3Rk
zKnvHyRQZHf5cxBcmAMS/T7tv7qCpMNvNVVEJhBZGpUmgqWEG6uCNgkiQPThUkNh
TckX7X2pb5yQ4QDYzxxmpjAqSJ/fc75PjumyrjM7a/eupuy7bocJ+ZsfudEz0NhQ
GVmOkdXjt9RdIHj+An6fXao/kBD+7ptpoA5o/kftLGH8Q4HrJ1c6pYIsgvqoSHOq
gDL/ZWDLPvRK8y4fpE8cS6A6DggakG7xBF6tiIRwYOvWHkv1zacG0JrM9CRCc0AS
CDWvjdBFVWfKupiVMwHKrg2NKclC8CYpb5TNMXrSu4SSD9sidU4WXjj33XSjQv+p
iXTWy+FN+HaDBoaTAL6ix2v1dIQkfuiBHEeBSDzINGm0WfcgpfTm6DtMvi5UH7Gw
PRJBqTfgQy8tBqYFpcrLr8V44hJoOjo6R3WxzRjz4vr1xY6PN7Hd/B400/sS07aT
diDQfLHnmFA9zkKs0xKKc0UqzvzBsf8wfp1zf6h4vne7r3IudHpMCeNLa1IhADhA
YTLTOo20dyRVSub3v8cHaKLlP8BXb1JVPhtKv2pP3wR6el8OUg+ISemInT53kVJ4
byYYqB9MUlPHLjPUvXiX8qKdnKLQMODi/2NvqL+eJNFObKgwh0ZI2U6z0l7mAe0x
xO5mZgwNR/2MTD/Bn1VL2ky83YU5Y0OYxOw1kdMo4S7f7EVBPlNT85jXExQUjXYH
kBfb2qa3Ie2FxhZLZpnw4/4gMnXY3e4yALAzxOOcUOHq6eSBoBfctGw5p7nZA1LL
P1Oo1olMscGx9miwjY0sQDrvu89Z3JVgaH8zEVTcxfvBF4X2+MpQdofIWvaX6x4i
sHA2wCaEJLV7LuH5K4abnWjbkNvHZ9ejXEkEH58g6Hapsg7Ub6At9l/O3h/tJp0i
DI6vLms6kIENL+uyJQhx5kIytwUFzqBqQSIIpUSrKvhFih+kaZ25ZPrn8iBeTW90
QHZ4P03THuHv71MSGBEmQRVjgqNCs3yt8BqMi68jgQBcr8BqFAQrqWj/6KHNPi1H
YrM7itIIIl5wfJ85xbkUienM9pmBKI+f/S86xePWhdihxJbLE31PRoQlMh5Ib2mS
YlQUXt0VV4nyD9HG2tpAHCqC75F+i1f/iem4lYwI4kjJ8ijeh3WDd6rnL5kxNQKu
QGeiJI8S3RsTHbwgRjhRRZ45vgC/6iGYiAz+nNjeXTYEcS9vYJOyJC70SBE36WFU
NCjLg2SOgScFAwOBp2H1/83bcNy+hZVeSrf5KkJKMGOuwjTGNP6XLi5/NNTOBBQm
WW8MHp65stBA9Mrp/SAgD98ewTcgIwnfAZ4yzcgsrkqUIxaTpeBYqoGFzIsIuxP2
QloQHnaVTli4265SlIhkm/7crrARHOaysqeo+vVV+Y2lpUxL2cRDuAox+LQ6E3Q0
VncmZGA6HZLS2ZihVROy0ZcY1pxqW37JDwRxskl4yvdWszhhcGcqNU9rTU491doW
LclsiXyamuzTa0rlDFbzk4vb074GNsA0+lFfaz6F6auu6AcQQMIK6QoB8At195wg
g9eQWxcbUMHkBSpC4muiWMfvDUKmUUd53V4gT4V7pd0N0RtZowMcEAtpVN0lBwha
3Lkgd5gMg3rkzRyUoQT7kpBBcPJfs/U35+3227uPMCjPJnekW6LdiP+aeI44FSgd
qZ3piTU2GuP3NVNEkR4jlzt44i1M6LCP0nxgzJRJLBPcrhiFsP7tVeFydRQtzaLz
Z2yXvjvR2ILmleGK+ygnE86tvhJrqtCSeIydZWH5uCbkJUbLO6jRRx7P9V5jspac
rMYR/gqDGTGYqWO5mOZ+fD7kojmlwbhgL6LqOTTLU6J+shqMGidx2bHDp16+9oe1
zfZdQJ84jeCCVnXoaRG071SaX+uVKmpHhQR07ULvtK9nhsj10egZ9T87bhjV/u/G
ncG6rwg9SgxfEa4uvPExQ/2stGnS8Jfaq9d9wLbfDbgnz6xPiWlx/xew7rDCgXvS
eHvnGrcV8aHoI+0YvIUVp6nduE/0bj9S/khiHwJakDnme5BMzdYNBaj6IOYEOtCu
uGztEXohbg2kI1a/7GgbQBZolly4msOA52oWMDtTixH2GhksG510scYnObY0JanW
FY/6lCuCkXPpl5xFhZMKcpXb8vxQI1wgMeuJ7J2DYwIrNHnfC/AvLM9dSgG9BruG
R9UyrJ8dXjaAMA3GkV7vP1ibcWEbd6K7az/gnfUQOHkwpWQ4fuGTfq7qcMhFuHqH
Un3G3VNjz2TYq9Qz2hjXLN16rzTzeETTpaZFfhyM9fSGOih19M6DkilrVsTIvrQd
FJ5Mu79mk7BDOsBF7O9FAvW1TYKJDvDTf70ZFGG0bgGOTuEKntK1sFP5IqzWQCog
Ax+bczjH7kmMGU1BRjUzafMmgtfydPNJybGH1YJo8LQH0FJsC0yn3neMG9L56RZB
j35ZCzVTWC/7n2CTmLWtHFqTyjNIUz5aigebKBGkWaNwGGg94iqjHZN9ss/+UTep
ehWK30LDfN6hfRfLVOZEg4Mt9FeNSAzYGeSMI9c9yqOmYWersRwu60x15/tukQH0
gT4VHII2utLFwyZQS9VB3ytPW3YFLI8+8qfRn+uHgPfgpv8AmtiaA6jxJIPa2MS6
ZfAbScUtM/CrFIGRItgkeRg+LWZMfX56H01e17G+/kT4UhNse5H52PWmQrMJG0/t
Jgc3WZHSGSukaFllo1ZylhsDJuCc7Sb6n4E5Loe0BKosy3DjKxHWoPdWBEhwg2yA
n+YSMPY/fSxpbN6fALTxd9sHB/XhcUEB4IwrlYbZfAv6adUDcrk0DBh91EWepkDT
OoeJt7bFYiTcA50feS6Qy/HEsxBLIf1LOCggogA944GeFe2GQxI5vKE6gl+PK7Aa
NK2mkMHMC+J6+VM8bMFTrIe2QL4oZmw6hncYNkQu6Gf4XUuOVAtPnf25/i0lKwoz
DFojXgbcwZIOcDgQC1QR8HTviKSntJ4CJipVLtY2t8L6TgiTpHouMgWA0Gf+AE2M
50+5KTuqL0WkMJjZAQAyVRTkpJbWASz8tzQjHlfXRr4+MpMtYiUcVAdJJQySLqK9
ZoQ1J1PDWD//7MS5dODYjjvi5Ykh+NHjja5dSAQ9GDtJz5QZUglNdgsYFGEjoLcO
InO4WGXXUvTUmQ1xMJV4qDoEV4d7ThXUimvy/tRU+b29prrd9rKdLy/YVQ4FcMt7
Z4l875M4ZhXA7VhKmgdLcvwtcM+yhwtYhzuYNjaV8euyShIkE2tHO4LdkoYRWP8D
ugM3BjIYvSG15k7pL2m6dY35hkrGX+6uTL31jnBMg3SNmQvT3Tb+UnknR2ERBvHD
wAZLUVpGEufQ28FcJCN22KwrgRsBBZckfhwzHI+pDKzpPbGw6lwaDuFp56Dt8BpX
62NBRRaRFF4z41o8EI0ikvgNcbVVljxogi7PnkQCWEGR15RkoWUu9ysaQPQICjNp
VkwJBv25nfS3io29TgK6CUoKB4qKnzLenb7cP48DoI6cBGPCOVAs5TIUIBYIGrCK
aHsYWHd9Tch9h1zWAl7lDTLEKMKJR+t2Zkwgrr3LLgqKp5T5HLnQsX9kmTZndpeY
OMVFvUPm0JOmegHc7HeNKXrNFyrT88jzFm9vOqlwyAqK/Njggh3JvjSQmyIcmMqW
Ta0Y5p2vOtpL6+3dIO933JNkc9WWvoSV7WLnSJnYCLa27l1c1YLnLn7OIWPeDd9h
fpEe6x7Jv9hTmW5nGbTS2E9E90tlgTHF8ITZJqlB9FZXc3YwtlNwTftiBauBM9KA
vM2IIstXcSS4ugwJ4QcpCjFILHOuZGFRjscc7IQahjFdTxr/syuXBszY/2hI3fJM
XnGkYyljpl+Mz3TkSM5pWqv7uAG3MRRwEJYgC/Nq/BJLdIM+fkp/xHU+0/yScFp9
JTWRNOkAtDksmTTvFiCYvtVPGeZqNoHRIs5hyx96kW0T6lvk1hEwzZ7t0BziKATd
Ldd4i/wu+ehxVjrdEPAPDXdWB4b1RS36cDAlxPOhkcBRhTMZKC3zC+SrdWsQgxJC
5orRPWxaWdDyXAr625f4ZZpGVdZcGSxFFR0XmvugRiN7Ci6RPOs+RS3obXbgga+0
agGjZJoPb3zXKO1/QkOroHsRe5nb1fKahmS6gwtudzNxg3h7D8DrUp0OGjEZMDn4
U6+fdj1panjjMlCAaOBIeO2lH6hOjFJlZrFhhICTKG4YLlhcT8mEas8K7pFw3XNY
Vl85sPQwXcupMEGguad0mmET48sLrTxzESNggIymGw2HOfhQa6lVOv4mz/A7NBjG
45wanD7cIBhiFhYL9hPDwxFb2PFMd3XSg8Mg2J/x18Iby+bc4ahudIqaa+gFXlR7
Waun9PYOLc9W4Ktn6ZGwTB2FASvxXbOCx4uzXpV/tbZ6BfWs7pEyNKcUzZctRrDg
8rdSm02UJ24b3Ox0RSPbRKFD8/pJy7XVAfHO11rv9/qaGPtJxuQ/Dn5DJ/IVP1J9
0Te3XcRKappe7VnZQUqXwCVoAbbjXzANwVDCzzUX3CxROXpokIYfMwktCnEowfjN
+dW1PigDvHEAO4nGlfVjrUdzhDzR90r+c/B1Qz8FQQORhe3+W/FKTGRTfVafLWeg
72iaiTaIYNVRJLZWIYONGGmPNvidi2xkNM47R8aretyhDuEcfjC8bj4eFXhg31Hd
wNJu0rqbbOW0ZtUIzhc1cst2bI1EsaRKkMQrBy2LEaYVJh6xricrmioh31EiaCe6
AQIengI33+dgHUJLlTkU0i5UBbvkdB0Z+tpx08Knjoo+jhwHq19/PwSj3hDZim81
K6Sb4o8/lcU2dx8i+/MmwMy6Uq8+sx8ny2HEsN34RBtDd+FlgGCP4aGgQb2YwKS3
ZE3dGVbHRDk2VXOmrIve2ryblTyRi0HO9iHhxP66vtlFhXSOSiIsnm94RVdjvieQ
x+5gLe6Ce9cg/OvZHZoPT4JPsvYrTrgW5ClgQaMqk6hZn9b15by+2UOecu0zgzR7
QDNBpo9sgLmbfRc4yFMn2AarE9v8mz/39LnVUGc5STp0ynmqV4OdhwUED8xRE8qk
Jyg9mJp0581ogNR/CKVoftoO9cFz4f8au9KGHoHOG+YsVKka+4WvBhz7Us6HFPnV
lIJjINS+TpSmhYJ3f07ouJ8KDXhRzBO2UiCJ/GJPE1155aqhLV6IyX3g+XoIBVIU
7v4GMAUe/C4DXVMMtQAnmLrT/5Vx40dLcSW61DuURr/ieM5rBsWfVLl/llofkgEf
pN8kOLMaVNKxj9LqiVdbXpCXoCdekwA2Qh+xjCxO4eqM1O68pwwwsEoarWGpbJ+p
gCnEbjZbEQ3ql8Y91wmxM2le+iuaDupzP25uulOLx/KCK/kcfoQ2WYEZAgzUEIR1
m0hRYPxPYg/3MS1Vue0IwstOVNISMgw5NpflsUbzscFiHCgFXl/QrL/m16Lo6fPd
F/HMnBFEy34mwutj7gDHA3jKu9S4jEKxuOv+f05m6ZSPV08UePQNOpmBL13VXRW+
3SVx+6wBE5HMKEJ51I0zAY/Z80R02thEdWLb5nz0p+g41VA+AaYiVXhCKk92P6CK
ZiKEKN2FuYfpCyNtEJHRUKPL8iGXIVqX6c4sQT52YI7l7hJJHCePCcEm17bfHjry
VbueyKd5TUPTFEO159JYiB4kma908ZgqQ/EcobUYXf3FtGAX6+s3T3PJBCH0LofV
F+mIXqM/mWF9vOCG1RrQVfVeK8Krkz1fUy0b9zH7oQ5RXdQ/ydIOLa9QUEtKrQYO
PxNxU7P1bduFKkOybx3lF2kEt+r+Ymt6k7rDWL3YN0Qyg1Y147zdLq3wvsVQLXRQ
EYfreG+xXD/IRspTjR/TvF/73yJNSxfMPyIr7CP5y4XcwA/4ONgyqAQRmxjFd9CT
KKF/Se8xLaHXLETRholtH2gSJ8lGBScdYUcI1Mqe2AWiZmuu4uYRsMUkQBPokWwv
dFZUJD5m0rsjxQq6GC/6oRzsoejiNzho2x8Hhl8RC5S2E6JZ0HqoYb/TXScc+Yaj
qZLrnBzloE/5vG8YYrIj2GSTtsONmo2LYvrHfLEr8c5Yr71BT6zGMN+P9cr8lfVh
siosCdofR5Nbp1iyjYNeaMBtGHX3N8FyN8McTWJctLU6Jg0VRm40onupWcEdbRsL
M0n1kyBrh7s5aXNaJDBvbATPnFaAAw4d3uSMJdIkcBLWE1WTWNDYoJMxdiwO1RyW
rfbnN8pZLMX28I8hPoLip9NlMTaAag1lJSKAOCtGxcblHOhnqXWEHO+8Bod8Hy9o
3851+GdLe7OC+F+fOQiSGzRDG3g/FQJR/0FO6ug+HubU8ttd9ENoGvIH+c4ZOEK7
KheHY17bPPsKovODCSRfjzy6jJZ5iKKOGokoRDPLjy4fGCa8OrJ8Fq2UJo7OGO9B
njeJnIDr/3WbPTP3QiZ5/4K9hEsLn78mR1CYhPks+zEUMpHYcHSeqZLHseJWQ+tM
UndnWJx5v64c/GSm2amhGk3MT2DnFj/gMTZxjNJ2GtY2NSU1NGWnkXdDoqZpoG7+
2raCW2phRAj+NrUKcGNfZuT9VuAftsKkUoUeeG9eYHx8VAe6lNYDvudwesaFs7u3
09c2dqPkBN/qkboOcxp+QDoHlFQnNSiZ1It0wVMqWSV81QuB94wGVPNh/OGe2rxm
rTrIIKKiUZ68JvCPvDVhzuLibflC0GyN5RfA0u9QcB2BoWob6quz8qp3hfwH9cSR
MELynn3GZHeLMQeZr5E4nM2ddfOkKFYL/OYTmswz+4biQhncyiKBRjX6B0yesiEK
SHBBsEE+RLeoxaKv8/MqyP3ymLdmgBuYxMRybfOB0FLhihMIV51lOPu/l913So/y
x08+SMpgsxZr+xnaUNUjMoBAXEKy9Y7L71r71c14pkmG/Vp4lVzr+I9OJ88YR+oT
Bo5+gc3W4MTII4yGBC6H6UnbeX8s68le+FngR6WTY1NG5P32zqUEjGZwcCGd0PIS
UjHuyT5Z6YGMQfR9kmfVdkI5B0DA+Pz7WDSBOWvFmYfoLeX47mzy1m+boYly57Q4
P6HRLL+4EOuWcITIeRW6Bu8WsH3x3It5EE1gg4ovhg67XHOgdWPVXE4oySB2lPB1
6L9bUyivCZ114PkqedLCCJGr/ZChHnDGyJsRy9ylCYh0F+gXi9+5YVbEsKRzW5H6
/nvLTdII13aX0mw/PdlOtJxVV8DAul8u9RHKo9G9RnJklK5sodQ/KORHFor3n7ZP
k3gyj8VeUfmZfnvpvSYp29Dn8tuT1o0ubweJoFJTTb6DcxvNonmQCGquYxJXztwV
myiLPC7+2D9Rluycb/hj2iC+BFPa5kxOTDI+Ede4VYVg2UPaHAQDtYsN/iHlsls8
XmT4c+1vpAYllL5MdEOEBfD9fcGlu/w7tbE7SJjFlL/7UHY0IISOomsnRfKhx0jL
ONsHDEMiV4i1xj0W/fn2tr3EHoITdXQTJX9qHulgCj0dxCly2YPBOcuP1khCKtBb
zoLGQIOwBJWcsDttBiWCY7nj6uBveXfx6F9fp9RnPpaIPWrIuGVBrejTTUVKyf17
BDthkPdCdQFlvexcV8shlY0NnUS39XYXHFUv2BubW5YKkilMp3tws0F1L5sQLglF
lblviw5lBYquTzflXMHXWfIue7CSd7ZZufBc3lpOArIKIWn2xZubdJxjwjE2ZXkn
Z0mJkgOLTv8vrVngQn1kpZOyMCmcyL2tUm/oN3yAasakS5pTdTeyUHBMvdFpYrpO
5YgXLdTf0rSA1+WYWv9+Zqm+h3rw/wXvrp8/49Xrs3M1J3SLWRiyOKTAOXJkScpt
bo3MfuRsU6YBI2om90rrinfn8XTRy0U5IRA4qo9T90NAmLSY7SeAbqnibX+cJW/3
YATEJUXMLaCC+zDttKgHUBIR+s6tlUtN8pmonaDGNOeiwQxWimDIToWoPCsoAMaU
7U7GcdrOo4Ty1L+rSemm0G8kcrKZe5FbEWgLK5MpxBGFVPnLWBXyy5Vxg/+JVQ50
oewSd93eIg1iGNiMjlQbgxhwAG7HzLph0VNHEY8fLK/YOtZRfZCiuknd9nGp0wBJ
DVzIcxGuJAPKcD69LIkcNresy1aFhPrsYwhlsfL3Xw8e2rXTs/ogY36inMhg9CWh
bz0b4uhXIyasnAZBrGu77nnit70OMO13sIfq/2QfmFmxK4Y1UuZR+IAo1lBLQJoe
+fjWxv09NzrqbnUvehECD2Sz436umXELGGBAn3ZAz9W6y4xpB27j15dOAhBw+UKh
pLkrayPeTwVt6azob2bVX5muL41jSzrMaX+LBpCQKCyG4QZruBRRtp84VHsU14AM
oKIuFzQiyjKYXnr2sjToJLs+/g5Yu6YvqueE4oUOjBtvnUtE2asLJmZk1+51leCE
uHVyqB6x/oBO2UzCF2Gu0wmKwbepxOhbzTkAO+2N1plXl9Q7W9VjXlUN97baVMgz
7HLxO51ub7WI6pMH18krAdu/PK3ZsqYHEY37X/PGQPNyoi65Ks+mVRyRg58znbdQ
8kJW33eKmiuQTs4GqvKvflQQ8ZdsSqr5VQiJ+zzwt8q+j8yK+4+WOFEG2DnBwUYd
n+NvUzg0dSFrrSnXlju+cy4DB//9CKojZbRLW8mJb1nYyQIPZLlhoz0V9fiQkSDE
MtpPHp2eB3/u0HEIq8maXyj8skWR1zbVKinRvLL8JdlnL8EozHASKuFWO6zGLULf
yBfrqQ2oMo9JqWlK5iW/oduJzGsr5hv2TQLSZtvCeHM0L1MFtPd9c13hG+MOnVBj
q2d6Yf8SKS1xpoT1p1g/0WJOKeTrh2AMSClX0Z/doCeBSJ3R+0n7oXHTvfZAmPi+
zGWW5IA8Mx1SlQdqmGP5MaJqmJu8mWCV9dxhoNFNZEeueyTyifDc2IP83PdCgnfK
hvwuG3VC4dJVIxRXNoM9p9aA15ItOlcmr3Kg4viSvJ6lHncHhFgbne1YiGcGcv9h
UECMLLIj72eBeJWDcKZXI2HP1RPgAFCwMci5FfAE59MV6P1TKZvf/EFzd1hCUEqn
wDnJFnJsKdpxXuhVnfOaYYQX7Et3Lfdfut5WAH2Pc0DfVJRoAx1ERM41faCma59F
YlfXFLHII7NOr/lSbA3ZIePgVI9fy1LQcQU80EIIYbkz0Xtb62A3cNIiPE5IoYd8
mnR0tfzO4lI8+lxSJqniE66XmciF6XJdnt3LiOQUoeVlB2IujdnTgGEiyq8b1jDr
CabO/N2RkCMSqWvovfBh8QQgFoeoq6hCgVZHhjkMCHzF4x9/cZCCH17jGAzSIPBt
+IBOjxx7/SxwSbKjXj95HRlN/HdIje8Fyftg6ISvIQ9XSXP3OzQ7N4TmTo4h+CU9
syTqJcVLgMmZozUiX9ue+3MTszgwKj7qtSX+9Jv7LFKSsaHHAdFZuWu2FyeEX54d
qmZ22Z3DuKUPPs3WCjbPPTWwzWEOPbtgzOr0jvWbm7XAOlpR/3kf57L0zPOmByIQ
4zrllCL84ZV48BpdykfsTpOLrX78WFJGDjB8kt4gzlmy9mxDWTwWvIwCpZvh6dEx
eo5toMq4aNvV2BO8BJwyglGj3XpTst59CnFka5PwkkUfGJ39CqitY8izQTFNdzeR
o18GyUn5zRiCUIn7F5fkNkxd5zD3ewKC+dTe8PEe44k8e+mHC6L/KIGr7iOWElnH
dcMBcN/ZciQiijDB+69x6jmEwPzKt4cZbR6rocvzZoDwrr2hTXCZxW0SkK1FTdj/
8JBBjpoASOMHApx8IVqlGkATShh956KzCYZ9Oms+aHMA+3DfLfHTARuHI83e1Ws3
txbegVhSWutzsjr3ugKhXvnRwUwcRDaV815zqUhfo+SsV9HgIVhBBTS/L+AGPv/6
fpCtYmKQMHcVRFLs/95rxFXt5owXPxgxeCuCdB482885ndckLBXSPix73AGvDolH
8/kqIqZXon+kHQ+oFETjQJQCFtIiOCHSzFyBh/H1017nxkD2leANjCw/BN0REmOk
4J6//c6CHZoIUxspC5i6K9qmXuVHN0QXEsaJxV0XULOwIS8CQgAT1X8cqUf+GZ6z
gnzpIdTRynJ7T9RbzkqGSyf4suhfdvhTaEJp8JiIcxrt6aq8oYUZkQXC60wEaWTh
DZecRit+1DVeceskUBr99skxjXKY5EzfUxbOARYC2kRDz5hg7AHwxFxqNYHhW6GV
meN/wvlVXutmCJ9qaFGju1Zdvdt9ffs757OMsM4K51x9OdkMd06kHianyeitS6Ek
h5G2QohAo+CxUgjPGUwOpQ9a1jyDv76dbbykF1U7OpxNjjLbdv2XFMsPT0QfJBck
mXW6bhgS8hchMFxz7wDKreLITw4ZHBQ/R8X23w2lSlGKTQbL5zEfeorFme3aaiZc
U9eQURZGXcp5Hf93Mo2JI3+aj9nkL+OwKoDPQXvyX/3XAt+MLvyFNFwCeSkjdyX2
lbBDdk3fCT95ydz+cMJPmjgrY2txaF85vznwlxQDGUL3hCNknZo9aNZGKF2ibEKd
t6rOL4XypguZGUOrrI6N7YALF4wWHTN2seAkxAt2T2cjdhNLjuvSh9vgZwls3lNq
uizmx3oml8ypKNyU+Jb3d2BZTSLKUQkcwjO1/uzneguizAbV7MZV23oyOeJy2Hhd
3CnvGOplOZLwlNRkT9xw55GlRKHMzUY1yCFd8PQuuuhvTeDLfDh0sfyFBYccpxZL
PDYQ4WFqhEarNvGWWH6FPMvcdjLkBOSXvsmuIXSFqmG6i57kHodUn4eryIRhrNOZ
/jwC8Wly9bRpK25i/MrK41Qjdyr7wuJ4lpA6Ajnf/Bp7ZJyScXUVAw8GBNaiMgN4
dJsDb5szULzy6SBflnbHxtsTBf/NDIAvYKjEtRqyYL/mZFzsmKeDxJegnNzQHxUx
EgqwgHge+kWfzCoowvZRmr6tf4O5O84ukrUfZ6rPzjA0y5jHU50EGfgOhwvkIHl7
TVW8U3aGTqsApzOQ2fyxYVftPAUfuBbAXQPGiZ5eVRnGA0cYIbH8VHgreVvJichZ
oiSquqk6EDLxcV2gEjRDbATW5eWNooJDsG1YnpbNCogbaMEEyrCmDd/OrVasNCgU
o1RiF0GNqZcfhxT9tGV4fTOzk85zbxA7ZHmjtW/rkdkjosGvJFBz7FuXR4DPYFP+
PImHjMtgbCSzGIqADNd/pFvvaI4rnOnZS30bCTMiy18HJP+KRb83WCiKM53jEpyZ
8jE7QRtcO3S58wSQUUlfOzToIFJM+xmu2+MYXE+4h+kv+xzIxCAFZY2NqOeGQMZE
6iuEHdsjK7aRdid3FLTmDYlbxrcrXReWJZmr5SnD5eXv7q3SJaI5YwjA2qMsMCcn
QymRjecCmyzgLTONhD/o+LBddOWzEktDo9kxM6UHku7N34x7FvK6HtFKe8Wvi5K0
YiOHjaUbs81ZQ9GIErDkr1pPLG64FiGQASLYNIrw5UNXINLleepqQjNeOb7PhrmT
itqTXPSkQX1JLPP5OsMh2NXFUWP2cs7Qm4QGDe2kkIzmC0sBxh65/o0P4vOP6a2q
HJI+gxM4sxZP8VJzw7UCB5Zy5MqqXWqEv0Tas9ce6+ZybzGavrsVNfEG9NR++6bi
weSAM6ia7/fNt6p34FIG+lMgMMWRYYiwIwEYnC2bJyMwRljtUxYqs2lPBh1xHzUF
DeiMiaXVZxhP0JS+2/dfM2C42c2/f5bcM/C9w2zdKMZWk8UlXyJv+HnjlqCodEqw
v+WXXEmv10/dQP0zTmB4gMNsz7L5SZvjEHDrXLBcfXYMb5S7Sdl5C725U3AhQRWO
ukDvCqr5kIcrekMzSRMvaiFlpHwZuZGdbq/OglLHvXzUqs84JBTbc6d014VfXIdu
2ESDzcR+AHjd6qveZZamubbY+Jlzr1yBZa2iUTb19T9YOasFZephwvVuKxkQ5voG
3+MzHcsnJ3KybIqDFSjfuXL05bKKsewgc+RYuTUrrTUHzGLR2fnecSFbelt9LgWU
YJCxfUOzGvC3+DTks+inYZgGBF5cYJAIFpPhsf4yqmnA7OSGwSlzUWOMekOuLhU8
dMwXYNmhZ+mRd4GSAomqkKyOEExbzzLFTRF52zeSesh7l3kGVZI8KANad/RRoEbL
mC9Dcd91F/h7rZKvde+72ob8LDc2MznZa3XMjZnX39mlA1/tbWGuK/BMoqz2j6q4
85PEc8jDCU4+ZKlcjQ2tcbu+v6whysqdZ135dOEm07jAOGt7AdHfb3A70hws1ic0
4ldeTXlE/TfwoKwQkpQETQNFh+zdQuaQnt41eledfeGFGCoGLGNt7OL7yE7STy24
s+0nRhwwgPedUR7qK93jwYvX5wgdtXqkhp5dnRBtXvBVmzMjcNQzTnRvgEvYFsUT
WineC/OA9HuE1oHwe0YE8cc3oWDPgOr34On+mQWKfhEa2JT0wfvoDzacXn/KBIHx
9nKGj99VTNIsts3cO22saUW69mSJ+XHbHFQ7KaG0vuGDZef5lxEqzrHaUC2Lppy9
petEIauLzmn1ZkJW2QbprktozHy/xhqU2+Dupzjj7xKO5EPuZOLdfPIp4ZGFA1HA
9yYc27WyQImzIPrCAySG0UXk/uLxxwBMyvIG/98oxJQDo8Nf0gu6OG2W2aq5J9oK
L/i10sHYqEnQPdFzIaVdcT70e/igk8YuYy3TDf6JBtc7wcvFFL3ZCnpllnydv7YY
ca9zpjVG8D9DFlJeGYYCHHho2vZjrulPiv33GcPOMzjLRLYUtprd45DvaasCnWk/
jFQ2AfYOmKDkixgNNJAFGq7H4Q+YJRO5GuzHKii5BL8+TQGWGUUqmXO55owmK8OE
eRw+hXro8gWP733Por8qXYb9oSMXUrF64S6W/FcoXDoJQnqn/4Mh8Tz+2cBE9RCa
JINDN68sk96b9snSg/dGTLPGaf2epqyU8g4aql2gaXW51VQCR6c85tkOq2JbjTmt
yc4Ibas6T0an2WGdRjxPBPOWmd+v3GcV5XWGVfefPab/xoxrj9OTJ16AQX/B5UHg
UhGsBIdLUwGnBCWNyOME272WfZZdLV+BUb/i8Ml6AAx5CBNRKoxecUAEpjki/hmG
B0rpfcopTQpmUZ+zP+hlTpRy9Bl49iEMa7FzuKaOjqPHYCYA0aRnq4NM5sEf3TA2
Kn7nqeqhsxvLstSip792tOA1xJxN/7D7dNOP7qHmhO58tw7DagRW6nb+I+58zQbw
JPbZwVWP+mapKCRQO+m5AOyr4dzvV8Mdb/mpHrVDlw8NOmSvoyyMVe/wrkw5ij8B
9x7R85iZASjdUBtn1qBY/Gm5D+QaOJIed4uShvHo40+zJMEKzyr6QFwANa/oOvwf
7P5tJ6fFhDUIPMT00Hkx5bw7J756xPA8EPpmTPTkm88F8wNHMidRSo2FCB928mVr
pFgcmVQd7NEACfTiVuAsru4uRkOu+HYz6RF3cnUHiIV1hbZe8D0tLiOFZVdVx4WD
BlughzGdbWN7cfbuCz4dq3KY3KnB1JClTUClVPu61LaYcd+56jMUTR5NCHmEVXuw
EHPr3FPl+l0KZlKhHtuun5OkYQkByvey2GJTYSjog09ouNu6bwQJqjvxq6embYeY
Az77UGwIe00JJBdKId3paXU3JqqAcqtUWGv3AKmeaUF/fjrNFvk8L4M6fFffOld5
rfalmfbQzR75ozxes690eUIV+S5Jg+eaHJAyNfNGobLUDjH6ploWScpLlS+Fqtim
KH8IgXm+fbGYZ4OoS38YAcqhwyT4KfA/S5WAxDZWTv3WswYZCRQjI5MquxJlqcJB
7EFVrjs2b87CavfUYev07+cLZLSsR+B5F1UY/pnvR/dP/Ux7YiskB/HGZRdSUAy7
ezYrCSeiMHnXaXKpHAYvF1Kx6Xgz9fyG2X+ePdIO0KLhTDSqbTnY1TRfA9snUcPT
V9yNFMRH+zyaDcrrq3oJeZ6qZzsLAFhY0cQxbtcVOijVAGBhgjL6ANWBdsQvZT0y
8VW8WeY6aO/YSxINdBSx3b2MkqyB+GYOb8ba9Cwh41101Ovb8fGbdJucjH2qpwrU
a+Lak1jDQGij7Z7JRgNJPYwIx7Jj/tf+OhKUZU1A5DNlvGTGHbvqlGFCb3cQn8y4
NsZvlOxRxmvFjZPwaj2fZN9gJ8H7CxBYKCFghEdEJqZHDKOdKNmFrt5Z3sReeUpG
/A30U82l8j5XKVbf2h+9oEmD+MbDGlOoXAW8Zi5XXCzW9S8Ss6akb/g4MhnzCSYR
v29Mg53zpmszRVItBPLgeYRK3vqoBRUfR3Sh6/E1oIr7Iv2Qm4uUYkb1Z6UzUmQR
LPvS+6YMeVQErvF0EOTZzXIHLZcSdCLW66n2+0SoOLSv6wjcvHz60jLkH/FN+gmx
TsjOXWZp3dUVM9nYfQ+Mi6DDEqy2jFrv2LDYx8VWS32UYxfIUwWH0kOmKFLPsRr0
4gfExR3sm6lQRZBNfH1N1PRJxji0X3mxMkKsjGdNap9TMZDX/i+R4vX9BIBDttFu
Kwh25+3W3Nr7keL6qOdHzMhAC9UXwb2U4YnqKbcrt8k7AMkHewwTl06rwZMCAIy2
ZpOQN80ExwXPxXYDihiwMEqvvvn0NIkY+omQXWaGEef1hYnkwMNeSDzChdJkFCKP
eG+UBMWeASPGWSunzwOJA867pTDb7xX31rQ8xcjean99PstOTHJMvGJUAOU5dVbC
TpdHkrheER0HvfTL3SiFni07D8eV0Lh1uv8PnCtOkcOZAYO5O5j19xvIALuHuvS7
JpItEJayaVAnhURM/6Ejf+9VFx2ROTJxe7krXA2oceI1uMTvp35pghyPnoAVBktJ
kfK3kQM4sMszSKWCiPdVFhRIb0gpysEWaNMRMTHDfSe2KPEuCvQiFvU+XpRKeDxB
6tioEVVzpIxEMc+Tp3Dt9Vi2w8KJkpHMxnLC18oq1RjQpGNzzvqtjc7TMetAIbVy
hHVM/mI2TdukBklwj88BfnIMvzxPuz4tWJ8tF/+SzKMmqUCvmXD/XKn/AXTsaTgu
xLhBGz1oInhSi4ouyMkZ3dQRjjdZYJpDGc4+t1xOvhJL6MZ6PEQUPwy1sQvwcj3n
xFsfYMtYk4NcAdIiGIy693KFKDJJVYHRdtDQt9AwqT/Jo/QmvqDZTUST7bA1SKl/
4RL8Izr20GTvv1OoHLqvixL9CkfL37F+85C+ofLdJWaxUZeO6uNVobeNAPvt0w8W
hlOhh/GyWVZ7q39sqY4YxYPUn8A259xv+HPhHNnxe2gHLCTkDScySWGZogvZewr3
JKkHSCER68Qh5m2l04kxzm2GQXV+Gs5EFcecKTpPiJGMoFWuqqHEMEmvH6+A1nYt
Yf84xgW2/ftFL6H1YgIGI0e3766XNc4u83bIZiouOJ4t218HdJkxKVVtacpOQCSu
PBUDSbpY8PoM17tI85gTNteyZBoOxHaYZTOH9DmovK+LSb0vS5Zt/Q4WO6BYq1ih
unUAe6IS/Mee49i91GT8uQKMF4pKysHQF/N55eFsK55ylNJm7H5SALm1JF8BCCT+
pVaPYRbC6upAWIi6X7DxNoFk3JsG/mO8p5ZAZBfBMJZo5Mxcx4TuF/I4NBa2YYqt
aMnqWz8dlOeAPTE2xMyove1rLoaIWc70yOCAm6KFEXsID01uAK7/59CNOSw6kfSR
dTpg2xyJXXFPy6ODOR380KFMvbfgiXjOgkUu9Gz3ETcMaUkZqVJq8WxcECNEcSSu
rLBDAinOEGkrw6hWXZdpcXWk136ACj6eqiPhJBklbtqGI/TC1kNtMpZsAMci/jxb
HsAwUN1CZamDkoP3YQpa9svIRsyCnkdx469+eXbOv0Xouu+sX1ayHqru7218JWFj
1meI2mYQs/MC1Ghe8VCUAn9gW5J7ChEVCtJNXZo5hb6c8DNq+qjtFWCOh9HrgOXl
BWiTh5N96CT5r9x/UYHP6/we2Sk5/kGCU6SDHfP6AQXOJPHiHB/LWddSRh/J9XST
gI5yzytUvq239698bsAvXlVZRYVc+IWoRyVuLOMtpQI/WnI5FTGA+fFdvvYDNPdz
JKzHbh7wHSSA1ni4xellS9h0K6o5Hsq0Edm5Ksp/gMceXlvT01lFuK8Dub2Yv38V
3Cao24Su2gNf+7lMEU+XlU/sY9XSvhHfZ3HQMrBXIvOZsxuyFfE4FppIbd6skONF
Y4jeEg/dvvRmrpHe4SMbnf5yXviZJ++4LfQ6N+g/XhM60/Y4c/7FUX6jUD4LxTjn
9CjN1uffjLYVL7Q8JbEeUFq1V43zSen/9NqDuqyVSiAt5RA0oN6UuCYv5Vab9P+6
4FQAtXR1gVJJGdTAEGJ6D1gdE62aXY+Hq0Bp4aLaqxnAyrKOyVRuPC5OMsltOV4N
c5kth9r8zxSyirNRLymBCPrx6XNo5ABtjnKbtA3giuRG0QQ4fVHSgtZmi+ql/oxh
pFi1s+Pz5oXd1oiFkerjo0zlvSf61hWtUII0J53trbeRexlQSbkYrtNAXyzNPKQb
7BaREOSGXjMWKAy+4NImueNi2+BZCYQYs8luwsyXtep+K9AjV38bLaI+6beFmKDW
Bt8UOC2d/iM4XW21dNatspeWKNCjI9ygMh4Nj5yrI1VaNgMMHFzuMfrbTYVTtWGp
AyQGCfge6cK4B4X6r2b3/ZHTr6yj+UqfszPQLAz8xrc5FM9A7eg3WhchZpSW0REc
2L5RKnUW2akVzDQxl9/xS/w46CiXisQu+YEnPS8eHqlqsnn9Xw62pKpsh13wK/Hl
dGjlmGGDj0wRYVF898ZXG6WcgMhr7H8uWMG6lXKz5OAnZb1V+LIj5mKNR8qcdRQG
qo7nZwoanvLO2IbBu/JfTO5icTnxjQ8ev+KltCzgFYm5O+Rta8v9OgREV3y0jWIi
5rQOOK1n4DNvJOp2KjVogFWZwNXIdrqeZAZ3mjyYht3iiCRBvgJ6dAqMgrmIJELu
ntNkkOczdNBbTgNzxhVe9SNyzyDkrdN6obldjYrvK7Ln21nYyk89UH2qyYJRxLeN
akb79j0id6OTW8kxqg0FcI7laV+dvyWPt9nJlufl6SbAuj2DmzcailwYfqHV+Smw
8Yl4zoLFadROr+X7n9DWS0vFzyP/W46ZljY+C+fUfcn6HRZnC1vXAe180J0PmNrz
5Z15tnjmIg7O8avpbNQ+RK1zJf4y9RwFqgyhLCHTh/tSj/jF7veYXGk6ZYRCDoz2
9tEVYarXT/X4DYin/8iyWtvEWzuGwKTr8dtGH7jemJw77qv9KsK4arYBzHrU+Gk3
LRNirhsYtMZuYEONO83BRQFz3mYsjievLInCeigZqjOznnwATFp6JiYnjzFYh2mv
DPQfb2Xg6fsRRQk5gfQR+U29Bbb4b6TX8QI054EPIR+Z0VAwmeIbyU37ATwbGi+/
pvtW9i2TxCMTUWm8x/zouVkge7Yqvi77KrbqnBVvrPQh3RzgZh5MWFtqzJaF1+0H
k0wEoVHm9gR97vwFDpp/P+G5y7JO3N6qYnWZO0yUk797nLRLNlToUiNZbjiXdEj1
xCdGSk6erM+5j4UXD7Ny1rCVK0nx9wYEXiaMjntv8bWLXnbUZXjzAc2rT1Yd/I2i
IepidA2Hlw28MvoTR01EH3X1DIoM1gm8KhbTlQYtS7zyE1+nuJk60jFiPWV+wRf1
lEujwvOkAVy4OKrBtMbL9XjPQnJJobDMEnW8GulPQLojdpUGfCc4nX0mE8/XALsq
fkurU6Eteq59vj5rLgl1HeZpn/jGCynpi2RQykg75Zvvsu0xQtrs7QzlL+HPhihI
IMKt6+b+6qT/CSvZcK/zQBaGlocKM133aUzHCWGiZ3/XDMQpEh1FtEEDtuQ2hLz7
V7+NZLIAQgzwcRB24evzKoVlbAqv6NbTusV7Ab4SRQlcSFrqIo6HLbETkYx0HOxG
8sgob7ocr2WyCF9xeRg4KRx3wOzqty27C4VlEPbidzlWH73CEyuaMunYgz/whQoy
bT9BCN5gOXvKXlxfDoOHJbxADJXCIRfSsTU189E9vlOgwTSs6c5YIAgLkfX+77M7
cVNdtGvMBbHmqmuT4I3d/GKvWG9uWtG3lmiwLS4fIDgEtLnbvEysnFtVKIBGPkBZ
DCPqQ8iFwXEAoCHCHJlUQjBZN3ffe0xOVMnrrSxqPCgFS11DyVnNUrBQiaJ8N/Um
pDXnmmmDVgFBJsVyQ3nB4swiq5RLxvyBlZBcgQdfLbdvw2/TTWyzhq2Qi33ubwv8
eY7WJpHlrc76iTMw8rw6iNg8FFeXqQHMMmejaly11hjQj4QccT9Et1lKnwBYO64z
+gI0kJ2epPVWpMIaW5EnHe68I9gi3QKI+fShC1W+XvB+EKKaIauK2JWaZCvme6Pi
gmQ3r4YMM0yV3mX99UYXUQWZGqKh6MenN6j0XG1WpZSlLRmTWZUwHTQmlytH9jaE
xCN+Pvo8os1YeEBvyC7FRSOzx4mzSowKBV1ebaLCLYTjr6nWuaZYkXDBTwswP1EP
ei1GKQpRTha8/YJUMJQL4SFDYC7ajEF+WYyoQZb4qeJTwuZ9z6PayTSYBdZG1Zsd
KykUZP62o+cUyWVo4WxSn7TDamiEXlP4ghOLURi42bvHx+Z2IA0WbkxVsdomGTYU
KUK0GN3hrmTS20wi83KkMOk5G077zpcJ4n4/3u8fsNL2UPwbGdOaUSmFtZdQYjQu
n64tf/1/Hiwunq4iJWvE6nUpj4KsPBKf3T5vQJBEMx6VrXxLHJGjojNfxLOyPLxP
AQ9U3JL7rHVCG7VsejxpTAO0i/Bpq7fsqF/rJ73MQ+ebWUt8tdtIAUm5Umx0/I3b
35sK/5pj6gxpKE92+0hS+qAHfhUJuC4oTRBxAjH1X4i5MUsy9Q/au2EQAGL4AwPM
B/N7n5jG21ku33HeAI4iUcZ/E/ALiEknAZhnnjgSOPi0hg90zUWxvC4DdEz9IT9n
Njdbxe5MAU/LDOSu1Abge4bjQ3Pg4FwVMI7S5z5vg3aFhuSmF5r5XbKFmdfOAGb6
/SdyLenDsoxG4h+RVx5kloNHKmpTFNSi7N5tKM2wo8BLIitjOjAqAGUjmcdyw/xD
Ky2sOKYYmH5jw42m7XknHDPUwbEsUrTHrzzNnFpoFcPHaf0BCXD4U+I/PhmJ91mS
a3eXxUvLEMWzvPOyqVxQUgn+7rFnoVENMjT7cyBGmbeFE9VjZgWbe1/hYBxQo7vF
yVoQSfCzMVilQGxV1mHOde+F3Xze55te3ohsGJ+duGizwZ6Wmj53XETrGJeiFuS1
b1iRyZDfo/uMB95s0gcHHy6cgn+RjLhLdxHUYhMaiB7GAK5t9EXhE7G0IqGokHaW
av03Wyl5JwXyWDdtcJ8dyYXPQNpVFYYXpHaOHWeGjEuB4liqDTy8nMeXK1j0CeqV
72uAjrEOCDLOX5h23kBFNi3VXqt5w1krImB4decLnyke6jU+NwdqQYs1pT/R3lyt
Hio+/vykeYRjhl/xAuWIJOjBxphENjuYeNxAeWV3eGO3ICpBM+uKseBe/U7Vn5+q
2baFPPxB6Lo0OShlZO/tcYPIDyXRsUa2kRtKsy7SV/jFcXBbYaMrrx2Wfe328fXM
4RrRkFG8MBn9XMyKiGq6eOHeO/aNlPIzdfJ3EzHZcplGRbObL7ui6sbbDlNL2h9H
o/2cI5zqk63w/oDVs/cv1OT4QCFKvI5zp9+tsHS6U0CalM4VDvX9ix4lGORbDz5r
VuPP5VgHa+bQ2ZnD7iCCmKd8EarXK7bJtugvbyVL2C9HNgZpl+T5bIMq9cF7Fbcm
LAJnvUrv+x6KPIK3ep+eIQQTHazqfPP3lz0tt7Wvwbg8QGIWcfwK13N12w8mDSVE
OnMzcbH+0zm+WWr56bfbOt4gM83BqgEn4XQxl88Jn7KR75owDlWFpdQ4GE6H88oB
SowKNJmyr6K4JGgO8dZgew+sHQXdqSE4pvcTkzeofXURufNzP036zlsHMVR+tm2c
LoWq8xZtnauF3+Ucp1ZIQTCsOWrcwtV1Xsv2lUoK0TiY6hb8hBG0Rd1LWRTlEGMi
rBQJhKQagjl/slUtmM1kpK0oCNfjxHovmRiv4Jd3s/nfJk+L6a/cJ2kL6SJQ2azn
Mo78y8IjhcVyQk8CoiZzSlpfTu+4XeJjZxQT9T+Ot3XpV7fXLmmgGMgmU+EmyD39
bJbXBJyocnpphoc0t/Kti3o8PqpRoam65z2Skgvmz1drD7F/72TZ60g1qwbg5gFV
u5UYmoE8B7frG/Lrn/50EzB4gSvUf+RLoA/I+gW63D/M7XMYLjOT1ap19S+oumhT
toOniWVinb2oScsW9D+T8xaMrc3KQ/ZiNYDADPnC6MAYGEu5I7LR4rkTM/yenLM9
Lsu8Gt2fGMQAEdfhJMDuQfZWEH5lxmOaET1R1Uc8nrfTH2SZUXEn7aqTfFLtdoe5
HS4FRki0T5yNtdlVD6snqt3UQYsINUppdazwuLbv0E/n5+Uhtx6K4Ip6ie2no3IK
RM+le4QOLhrIBoRtsQ2x1bReOC9odvtZFtBvCSoIcSwsyGx/qkEojvt8EfTMTZ5M
gPionWP1m/niaHDuqykUzcdSL2Z2dybCz5tjv9OkC8H6Rv5AcQSePeQb5b5w/RZS
rJ+k9ex/RXZSx0y1rg8N9uu/JwAGmOciuK6BkZxxarpINvVFw/7xvalE7XN+vL1P
dnlAByD7rC0dAm5s0bKxxSO2hp/fvBhf/4+eYdnNdc1PNbJlwJxqwtOjgpstvUE3
FU29q/sXXe71RV+2JMVKjRT4dzp3d8hze9loKW4r6BJJWW2QHBUD7JMaJ6BFraYU
JLt/nFI0f1NSH7IPmuR74CaTsXZqmTi2jcFetRzX9hzibU6T6qZqtSw6oVlYfRr3
FMEjQxTHvJexUpGUy0xviD+YlkaLydMi5XhOEhpN3ry1lN64DTcGkEZUG2Rc3HIs
Jq1EzPLxP1ZwQki5pHrXcFNt8c2LeeTYKvvP2Nf21fTTcv2YfhYLxuof0Y2KUboS
ffcOgQJ32ChX9Te2Lu8aB2TVWcctziGSml5KmdxfNZb+qATe/Y1ZXGnQogzEkY5H
WU4+WVVUbOuR4JBbsCN4bY9Kmk0h0kf7eg9dVD2M/i2s/elNRpROnHS9oUt9u7+O
Zx7GPyVLNhB4ZGu/jiubn+Ki2gOmVCWzQKGiMh/hv6RO0B7ttD1fg3nVot239bHo
sWLADE9NrMZ+UU37xdttcH4vcR7oqFcyRNGqMyrWBUlVzn/9MexNa42PwugQMzt1
Ups35zSzr0AL6PEPz7/LMbZatIH0RWm+nnV2ea1Si3ZF6HS0VVRFIWmloW1QZ77I
ojG4rZgnlEPIJ3KcLBT43RoLKoa3WYapVgJKubXGy7qcBoonWRWFFiv9UVVAx562
lX4pCTLJlnrjmDajVyZ+JcnBhGKk3ilPxvnhQpY0sHExu9k8Rnx0njW9mlLibjGY
LRsmzlViTCMdX7bMG2E/9nkfiG2lNIN6ACbDEfHSFYrtO2GCD4fEyIBdy0ZviN4F
eS8MNyZ7Zo55P0hg1DvtY0A1H9Ga4QiYs5iqUIz6Z8COY1kdTLv3b3Yz2ldmgzzU
06avwpZ+zL1MFXsxkaXJtfOmNhXMOnbC7bt8olsp+uOb6K8Y+yPdbgHfsnaSP3TO
BBWVm4ogEQn4X8BQE2AHN3aZHUTdOW5+gxYwqUHPwDZDdlOo2p8iUwUbH8tf63dx
IW+ahxA4Y8xf3ida8itykKNgHS/dOTwWcmnjyOjDNCA1M1jP1CQFPsdWAsmqSx+M
Lh4Pfjb6qdS/zMl76KuGbYnre2O7L4S/3mq28K3mogZgzDxExWHq2bzRyi+RvWql
ICqbog6cDnZAg/m41B3kN2KxtKHYroMOJp9sOD5nUc1Qz3hZsd/uJWjU1vaAYVOW
y/6sn6WmGL3mfjp564U3d8nybyuE2ynq31zchSDFza3uKYKHSXFrpY9I9DDVJZPq
3IDFvld+uXeydsxNu8Ng01a8JLE0QD4nF9yx0t7YsZHgKXtSoqMgBM7fKwV4M5No
OoSFfabmR6gUy5FbVfjb72qJzSbT18KQxAA5VceIyu+/F9CWFQF8gkdZ+X5YWGpo
87cuKtfFGHmBcmpk6hw+Rjx9vL2sWYRYpDvDEVqisGqruljx+IiFtMsa4Noq9grb
pFrcEuS8/CiAiDk/zQRd0K6vvRdLXCoLAmRZcjqk+sQ49nf91YdSJjCfGsyMa869
wOGEObp338XWtHx6s/mdBV7mkuVumrpKe7o6KBNO9ItuWiJObg3A1kCuK6WBw3X7
wRsYIEz5js/c3IBZsDGJ3RTHfMflEx33QIsOtQNX0jlSwd4l37HhmfM6h60NC+5p
kM5dDHsh8RRG+uIBqZA907C2/7s4LCnDreA2qLEMRcrRbZ1+Wchp7Mx1ET63LwfU
hkWEBdDw6LjEPjtgCaVocNWwqAqvNj1oYpWoTY61qE5wNOe/UTBRnz5MlIp2tkB/
NQDpgphvzCa7USAx3/6/uur1MjWxAPDbx2FefA3QQlHw8TTg+bL/xwvSVy06l8x7
4EbcOsW01S0xvuZONLFvosUfrE4RavcN111ZCC1iQRKLMQFT5ayXCZZdthnejQtH
xmjfu6TnNnJVYiwjnazQb3n5MX7BEKvz+L30WEiSvJQo2z1Tw1LxYhA2pfjEFJqY
NlbjS/1mcZQ61X7I6gUNBdbnQN/cY2tWic3fuGCealJDQ2BXEzidcPUtAnHZYJhL
c9I6c0BKKFeIG2eHX6/XaiyHfKsmbPL9rkHThpRW3uG3JnloF423TUuKeoHnyAlS
Fn0AEXH4a0rfq9i12KwhZgugyH24GjabBVMEunxype2UCwfNtsTUgaKSvHBjQITl
8I+zE8Y3ted5dr5VGebtxy3zf5k56qDQmUBGWcn6f4vPDv6UhLPv/NoAZMGgX4yU
PVHinaANU/TrpZ8CaCgTdZpNK82qop368FlgTK6I7MRrFlUDbyGJtI5G3ZMIxbCd
HCjKgSMSNca/DmI8ZdGkB1lodAs4Yot/FOTeJ1FUIRogFCaWj53OzxVN3Rb9vJhr
i9dxKzE6fI2WKKN6BwANy7019PjPRwqkZfJdZ5sLBx1bef3ygu9qrmYZGP8+7trg
ID1wI8vIxdgI0+45lvzlRIt9Nr8ZgIE9IuqRuG3IrvaDLUDRl7+bXBCnv4xsQaHr
JWsw0gJY2A4mZ4ZeJpkEcZ8vruLYIIGbOtOxjwicSZMBR2oIUvRHEFtvnA34Pduw
JdNIZ3fAOMbXqW2fPEyOZkuz6UlSL52l8V/x5QqxbEk/0X2ro7Lw2Nq4HzWydXY5
zsuYjO8hA27mKe065mN6/xlDZNIwwqJThmKQDcXfL+jS89S1RVPOEkpFlmisbYLq
xRdm69/TG0azEJLxmyJTpwhR4U7QldojlsTu5wNHrYdoUjyeUxYAxpWYq0OTDCBb
TtHONKrsnzHDGaK4wTSL/yAlThj3Azo0BUjPLxsGYm2ujcPmBXbYYf07ZGz2Rz1C
4HcoNMVCTffS+CK0fMpsSzFjJIThisdL+Sb8VTnq9Zqdeo7T37iFygmcd2id7WCr
ZZyyl99Iz/VMLMaj1AWxyjSyIg1EV28dfpyu9OcFsb5zqQBVdfvCu0kOrge1O222
8uMDr6VnlPtgxugJbYULDuLIyK5wMk/NNA+lK/8rRIE+POj2PAppEoSPTNxL6b9L
HThDejV3YM6pqb+Gff/oIScc5OUccSOWikEJbD7bBizSFCxPwsds4zTdP9ZyJbaL
u6kL2oFd9b/jiepZ4WgQvsO8kY/kprvLW2jxH7kMjB7P9xrL4KuM1Eq8P3mOctAz
p4KY5mptDKzmZPeyep17z4bNHWDaxqYLt+AsY+99kt+r1rUUzf6jwVsmR+9maq9P
NPp2P//MB6tOOGg5dWz7q3HbqsO9LlZcCz5Fw6P0An8fZYXX3fNktRmJgbfejuu1
wzqaxe9XD0OBSSpq31fL3+4a22OfpnCOgvnxGhyHVhL640/v0v7vchLLJGut0lJS
gLM+6XA6JJQWlhrJUkhMsdQI1iPUkH7D9QDoWq5UjZSGyfMWfRsEdWOvNGu2ABvi
VUHDX2rJysjOut0pvmK5779ErwzKkrqFr0THM+/RvUDmcN4Xfi7m0VXcWIsGzwlk
2q0jZYn0l2L2JTb4r4AiEWCPUkqkcJRmGbktCoWaRTmIuZ1zJOEoYAetbWPy2Tue
IpuOSaOpXJWRFra0j93CwzfZwY8VseK0bsf5iXt/2SUs2I9Ndmx5E+P5cciV/Oed
H/ltxi3WNe7Zel2KeIdM+fpumgSVHQ7ZHz29z6vguLceS9WwCbwL8rHKd4jvjpTa
zvYmCTbvscBEVW8coOrvDxUqR/2avj4MM5MFcVpQoAu7fHQOc6st7o9RnE8Xciyh
aGzmvaVa15k3fWukPBM9sYOY+uQd4lSxCNDkNMggpvPlW6sYNbdin9DpDKPK2v8J
o2YeCQeeAQI9ZddmkROF5TGiVFh1XTl82rXX11quNQPIXW5RB6oKM/VQQmTGMmVq
gZVwGMmvj98ZhuRYa3xhiKoo7LkfeNeCzKIT7b0CBKbfGXXBCvAHOb8FU+K/ASG3
jWSIhu6X+8w3TpQL34aI0w5VMCNRnWJ/lmgU2lWIWS5UPAy3yunFbtFIUhtX4VCV
6V+XVydZbcALOQq8bzIcOsrMwUBv6qCkcD5EnVonCtnn0pQAsR3wakT23Z7f8LJA
fw/LmE5EW3oTEr48WoxpBJSeesdGmWgqKiIHDIwupwbfu6WbEjIJTEpO4pYL2zjV
eLC2KDwVFMCfacAo4p1ANKc2/+gbrAZ0M1baqNSG40p5mIX7ThXrxZdkbhzs1ds4
MkXzf/rGtmZ0Vj/4QCf6IQ8rAOsH80KFJQgyeW+A7vMCdbX2gt/w0naDC+qfmV+2
R+PYU+/FWdIjUkH7dq8wElfSKf3mG0NBCy09g6JUsMh1DJRKk3LEwFLwNtIihabf
iWtsnkogDnOu9RINrQ31YR0lkffWAb348mTUo21jFO7aYEYyn7vZy5IuIIc86sA4
dxVmvaroxtxWmKYOOTh9JQ4F3IPitnFdTrZwXur4PIehcnajyRRsT34msBKqznLc
rKdce3Ar/5EFMZvlJ5nzTnTAa883vgmFFHHFmXsRzXXURyyiFJ9Kf5ZRC7MalInm
X92p2S407NszEBqwEQEL2Pr0/OapHsBbwAGHySMU4YQPiA1LQm4KUKc2+f2qBk/f
lnTWts/JfN8KTldDgqa4I3Jc6TkTW3xtcJhv4zJdNnK4XMFoqaJnHyGzN5VRcUdX
HJnkWp4OJkInRxZGnOlqw/c/h8iTc1O42nWkZ6oZzZz3wFJvakGgTbe70Qg8XtkL
IyUIm3Khh+bNZunVzlgZaffbgleJeq+8uC2zvYvXK8x3QqaYd4bm8Jjkc/QlJSVl
sick9PSz+XWDLgSF2QVe19jSu3Mow4LlvyXwvW52Y5LVpKwpJNXjIVMrD+fJHuMm
tc906u2qMRlk3NeZhA+HMX9Q9cik9fCuL8/MXTHPEuJLF53lWGPs1/sup1ZeUJTU
p6ojlf2vNh1Tq7PoMeL18xIJ7kq5rEVYhm3GGdQm5p1ab0vspSz4ShAD0Y+85O3g
LRE3375RqJyAx2GOAcVCJ7ULuPz56uHiETAZcGQpn7nqPC95It38eyQZ7IOCnc/h
HGdM5GVVfg2N06HSigIQKAcn5AwY3q16t0PbeVMiCEVmnXHIai/8pi04DVEwojoz
T4uqgifAJ3B7rYmxfziGwSnXxOYI6DWJ534R8SfIvBDzl2aHnup/IsRgw6FBMmTc
SD8wRzVlQ1AJsVH51LfN7IB/Xgbr4t5EFcGlGI5AZfL2JYKPx+FWqxMV6P+zLVWy
ZeYSQ6obWqiCEMhuTL60DwMM6OyKGfOPpnxsYMEEeO6DS/29jL8/TTFPygvlY7iL
XhYIUKLkZaH8m9HktWq/pmXpM7S0vpjcWBivX/nXmIMqxD9TSr+Dq2p7CyIq7yNB
XHoyb0ZyX8dKMCc5Ka1NRrxl7IoHKHald3guRV4JC/J/g70ocHOlv0g6TmybMM+R
ptPSQIKps1r5VPZFEx/2U2ngvTUNuRrwXeG6Dx0Pzg6REX3vsNaa1KyvsFtwf6Qj
6hDtyBG+Oth6fIDd4PsQcShD3I182C/ewIilUlBHVDhoyJnJc2SqyartmyUBzVcx
Lq4ltyaPq68b/e2BTjfi4p8ERo7iJ98StShIOKZd8VkdF+5mHbXcjqHyHYIhW90U
sQzYxV6kZbpuTYNUnYxW0UlU7+/N9E8LKfOdMxwd/wA6jSTZPo9eEoINcN3b+s1B
beAshWVVq+oZOFv3eZAGfOMQapoS1KqSb3tYgP4IW9M06XCzN16J4hGLMIXjJ/gE
m9VFSXSzbk6hqvtdviKsYxrQeIHem7pG6H8JdeAL9MAllUzbjLjMrBTWn+K24WzS
2XcgDG+egqLvHWXymFfbpEbUPNd/c+zw7YLJacBqSSuPnvx0tCMFTrpw9DnM5NCO
JfEPmwVGvoAxejY2q3KkUqJWbrVEHioGG1sTze+AGZ8G7UXm9bh7KLn4qMWKrP9V
NCJtMtU9eUTtuj2YhmkaTVm+y8soBgNfajyr/jESfgtqguhA9ugjUVeadibvx6Je
CGuW2xyvsj1veiRpRe8VKKEkrLajPDie8LkUdm6hpa8uXETsxem2T+FdldbyzN/W
q0QbR2X+0wDa07bOF6/KwnM386PoJFfzW+TF05XAnhhc0g9qWdPnhbRv+VJUIZJe
chyd0cQeFPbqUzm6NsgDR3LyfgZJbF0nkHqWA9RfebVJ+mbmpf6UQfVN9quwjAts
2GeLghXxlRq4DD0m1Njgn2NTMWGZK4SAybJwWVpPnxSfYcB3msWwaF9uTzLAvCMG
Z29VIaArgEd5q+TtwJ74hHEHD2sugTvr4jPeHjhZRmH0w5YwqICEw6DrJuNJ+gsl
tzYC4zw7b9eb/irpCXFCP/sNrAOU8EQQSBDvV1UgSv7Gdu5HHqsrxdxUur1KAb6d
Ehuw0biMPDxIAG7yQFUwNS/XdCAasSGcCXGPwiCzaeC40ljBwRu1MKfVBOW35jNN
IsxUISPQR8gdn3ZlW3J6CdlGroVUk7Kyta195qvs2lRZ0c5tKtxXI4UkEyMj5nyw
JJmx5HBiKj/OqP9yJHOE+8TTjZYWRxEv+O8cT1lOHFGz6gid/yMDL7sc7uDrRtiU
V/Iq7BBR6+FyS5dokklUMekrUYe1ntNbzFTXr3MHk5KgU+J+jvxqy19hM+J2w5du
fD+kKSvonmoF1uKyG2NT8ONKdamHD97IJoCWI49nB+xxDiw6x5ZwHFplZSpm2Fmc
xWrWHTiZLNVnw9plFdCxCk826gZeGylo3FhOHzcC+rh1eyzt1pIwvOmxzIXoEn0d
/oUo9aC6B9aXcDYAPma4AK2GUYZ3kWvApwvH0ozLHtU9Sl1lzBYiq/nv8G/PMRi5
oxcV3TYc3NAKt5rhuJ0gcARj7ZyM4fqGPZdogwNvSHZ4wrui9tI39200Pj7hrQlB
Ny5lqksfASyw2CXW5qwA0khS922AVmi7qNuYVgtm2YsQkV8iAazZ0qInSToYIwbV
8jHZc4FpRjAauE8hIUjpbWKMkjsAIHclZoC51Hs28dzxtGOuEcuSfslviVTfihW9
ywdEhxz3rVns1tnmgZkxx4RwGYDr3SjBgigYFiXAcy2CXJyX8z3JFpzrbv7J0IZp
+OVJlTwtj1KGY+WBdV7Cxf4kpFpQa1jqmHshZDtrUCS2bUbpXWXHe6Sh+bFJ/zqD
m+KmFpctmwVgH2Wc663dYmbd9iBMZgJlHB5zLfkXD9A1E2QD5kcqVx64ATpl2bWo
ExjfyvEFgeCqzjs1oIvEzPdmwZG3KZJsf40vpXKEGzuovb5NPPu/EAKwsKi0oQtX
rVRTF93srK0C4dWFJfXAc4oWEd7f87dJqczpxzCxSaqLaykPF3Wp3GQbJe9JGzS/
NwQZOM/mXQd98zRwA4/F4w2XfPbzcb6ye0yO0FSEtpbxDHP5Kj/y947K6krhjZsA
MOoDWVO6ClG2Tk16LunuaSARsDxc+jMOETQjla/NtbBGWU/tTLZ6LltI4DvkOe1A
r+FWF7YwAnXkH+/d+seStR5SvaTldSq1k1Vi2KrJo+T8hfL/mpWeQmGDbNr+nh2E
7pfYPa+IezN+DhtM2I+PQoytrWzehGKHd0M3hc1oVfk9sC95oNcw25qDLUTeWlCV
QTdC54M8PUrO41wj7GTlHSQIMliYz6Zlwl7pPz0ktGPaYg4z7LRaEvDiPQ0X+FV5
h2w24pu0qW+4+dTlttN4qGCGy7twZjjdMP3TeBov08W7qJu7A1W9UdZbMlUdfxNW
qfOENTvuyv7m3yf2u1tfSj0KupR+DwgFTjDMtkDFVgk4dP4nLxSbr+kapCUSJ4Sd
qKqUpj7Gg9qnkgWSwcCE3TWXzSrdTxgFYCK2QN+gUKzAWmwHaPAspygOynyhlxct
tT3VvR4TdKhhtZ0LYSuLSOvjPX0LUec3OQPqtl+tRW48ef/STn/IOwOLnzjmB3sS
aftviaINgOjmvcJ0sSFpd8ynK+bCYe/6Um76hDyUpV2omXn3jvtV1U0txcco9wYp
OoJDyYwiUFHRefTGkXbJGQjLDXtwzU6dZOmDIJm+/LMftHOu8cuHiwmibfwid2DP
WV1qrZ1XJWQ4Vumol3HUdMSFEqIdbVENPXC2/sm8HrQglpJWKHe1sUWnxCuiqWKd
ITJJl7O+M6v/e2oaIng/aeVg6YdcgNdb0lx6nXwqKKCbhEDxi83PhBzZwZns37Mh
E37j0heIVjcqd0bhG9nebauUQOnnoWULWNJZpu+lNXOOltjdkTpMvijjkdt0flEN
VbAIlhLdx/j268OXnwNbZE4EVLVVFDxWLjpAq4thg1kHws4aMV3ECUE7aV53E1G8
e1z85YN9luzDVOTEVucxp3/jc2QcSNY+YP/Qod2WoT0sUnU2m36M+FqVhSWApzN8
d1wDe+A7p9cjbWnTmkN+JMMUe6oM+N7m20Yunh/r/b0aDVYgmwee2Qq6hmqwKmCt
58ibI9uosY4i9vxmKmB39wkFKeUWMajvlTqVznBKFRyO8J7Vfco9iJneCAp2iTuh
YZKWcMTRchHy1bXhKY8Alnp0U77PViDUYcCZIG1xuu42dZX2ZnEHDspda7g3yulH
+AwCTiDQ/7XNMi5A8DN0jrk6NKxWjHtEV8VMufB00oE/yxN1MZvgkYRL4oZCSxUa
eHlWhplxCK+vdD8ojrHZhJdcX+VR4PZScrpp5qIaaUS7hsdRvnnE5tDzetTpqu1C
k579cHPVXQWlVBMbq+9sEzON4FxjQQfXjIB7WB17NnlE0QJ6m1J30AuNttk/AWw3
OKjvTiKeP8wclNnzV29FBTj+Ex4lt09mte5BWtt/3kLALGPrZi2b7okPAKHCamch
7TAxjc0pWNFSJL/YArGDPhBoICPxPx0cyosiDfwzNYadYZ7tFnXkYUL8ufrVPhzX
Q6rU9cT8HHMbQY2Y0ApG8CbE7bOKK4e+Vxup7yW7g6lYTNOrDWjSXdkGgYq2xNCt
vvWU6Po0zmbCWiKOTydmkiBm4ghZY6KaKJ6Mp4oNUZGlftyRUGf5nh0N4nuadhXV
SyYC8BUcwnAk5ZSXSEoyJalCcIvicaH7b10PMB5ccHnJe3nhw0I7o6eVPGByz0Gr
MdUKeUOfbmxpwF3xlzcnLKSIAAnmfWk/q9gkwzrR/nLugOf99BAmSHOW01C9NF7n
IGL7o8hikTbXJ174jHPov66EyILi464/W1xrDwMXPH/x2Gw1JlOeRcbullFNAy0n
r/p6j6zN7JfTahiXA7QVK419SvljcAhsAHPeD7Khu+0I4dcKAQFDzbxdbUt4xy0F
YBUwkUU2M0oMdj7wsRGJZfkEqfS6g8TQrfc+9tSJq4p/O+AzaKUz4dkdkQhTC1YJ
Cye6ITwiKsCGX3/IQvI2+w1eoNcx//rI4Ma4CVuS3GxiVP6OiH3fH1TCRtdLv0g1
Ji4m+BsIdtnk3em6zUj2rbC/7khqbfqguIJdUBU2MHGp2ltHRGeHgr74xI44jM0l
Sx1vqmU/pjJoibe44elgK097B79JeFTHKI4IejrqDdfU2GnN8IV8P8FMJ22FN7Os
jEmtUxydfLVBfLFhy/QJfd7z/Qe/ENBIQX1VeOnyDrAGWAm6mOmgFvydICIjVLDt
p9fXRF5LIG+/OGmoqNlNLevWkNCQjKIFCMV8LV8vW7sHLvOfbNM94hrC2K2xN6t+
3Ytsht0PdNPLv6ekxJuSUw11992GetgDervcZ/A7sbB/+Wp/IGU5Lo3eZBaX/aur
fGJQ7IesoMae4bj9TrpVgYv+UhiKNrM9laWuaIp6Fa8DfBPvABdJGcLEGfrWdi3r
7jOvZ/IEn93ygXDWpeiaJRxToJAppBfuEr6ocbpoi3fQrDqsw5OMXhB8Yy1pGsPN
5uP8oU1N6+/Ta32JFijAogQ0fQPo33pN03oE6cf6iyneZ6Fn3EqT/ubQ4vQwCjce
56v8hQcF5Vvi6D5qHcY/P4rbKH5fl9xdj0RFw2ygGbl3Qj1Nd3WFMjgibrfG3QL8
dyy+1wyyprkHYRoZZlddRsgP5Aix13S90wJQtzRctFVC/2qq52iyD06XrgLJQc/t
+YVWpBE13EALENlmj6SUsDGjq6EWZsvU8BLhAm3xz40W7bXaSJw/t0OQf/ril3Ad
EJHxcr7ZaU9G6obPgdTYBowVuYoM2y2Tmqqo8Pv+5Hj2TXlr3hL5zQXBgGPLEgRp
gu0lw+SV0VXhJjphxsJSH+66QMU+08ocKIw91Brm8VT16ymFAiwyvCempFdj8RBb
KjegkRvtwjG8qvNLgJlZf11yncWbvKuL/+sUUc4/y1rzXUm5kUyHYL0tb98wblGs
kSeos0e0v/YAuRTtJZks2UhnuzfW8Tw0VlNWfuqy0wHAt05oDgnHwvw541QIczzM
6UzCMjJSHv9IJ1650bZDdLxP7ZZfPkn/LX/Yb0es7qXvxkRWRemYWiPpQEnlbLe6
iJjtK4hEplLDNWBxvawoZs5+sgAlEkcUCoLOrWtc4EjNPj8X+yY9mjuqv3ARNjON
hbRTV6aAO56HtCgH18EaEhEKxBRq/wU8KSqHRxmeHGFYu99RuyjYKpoU1iX/Ar9P
32CpQznEtMCB60P6M2djCgLoQ2do7yCv+usjU4f+ODqx6wltKxAN/5qldWWnWMyw
0B2OHUzj/V8sSpN/Q0t0l41Jt4UxkXUCmp2T3AopaGSoeeU8nHohJZXNjGJrvgOu
d60gf4dOZ825oj52RGii7uN4T8QYoSG03JZVZjsm8kPiJQegw4H7LoVuwMwR9CrB
aqhX3oIlaQkFy7W9R3zMhS0YcAy4FwEbGHFBH5Y4ZBarKj/5sW4tEorlH4afXcFm
5mi0IsF5/5JN9eZVTS3qO+ovYD8Ret1IYH9FeO/2h5INX+ln+anTMoe4XMYB568r
KiLtrMZpTxdxoN1D61VNiix8RgCqN/BDRFfe9gxp9agJ3CHSgIj9An5xq20qd6cq
0V3CUizqR0dE+L/vbxUnE/coaIDhmPOaGxPvGMR9pjVPKy9OVKBV0tkhKWOpNfeB
IoVOfUdQly+KtnyM55UrAWaugIbiboDZ7WET0H6129BXZaslyHdmQaYeaFpDPq3L
AsCvjcgq9fuDQc3PmElh5aMfYFPzfwv7K4SGYEDowja3je8d5k1FZmPI37O+GFGu
q3F/5khCGtAcahd2TnYCaGthNKOtfdFJXv0+zcG0hRLPjCNRuC6KJpdndr9wohxo
7u8JqOEQ2HBLViihSWlrAdu1nigj/DdPR0GR6oXTSnl9/FDpN3PZBWtWstcR6VuV
Sn99EeTO5y+f0uBjArvQT/YvbmAUk1+P5riDWegv9g1cuZaXKLDybFIMTq/MFecn
ZatQ+X5gUYMBbDUHc7cKlHv+xialtGC5z8oJ03R6P4epKRWM4pxzS29c2Mgar54e
Yl6ByWCo9waexL98f41i0A3t8JpIqwE3Ghu4KPryvMdUu1RK4tjr6+WGXQ2G4BgC
lNpViaRSfDXFiDNkcH2tYmnDf/Nqn0Jn5BKkirHr1qLxkWDI0UnMDxdlGqZ/KuFV
5Lpx6zSDEZH/rHu2GpFM7CWjZiwuZUgnxr+DxkGkMLzYApmCCxwAnIo9jVU2eHY4
3cNwWzW8zpoIUBbiCbx6KqsZCOa+F675RDg+QX8d9x6OKEtnUuM8cDFWM8+AIUqs
rS/dAWsdIEvcHYXPowy7hQ0t/9+Mb/1jDy/QgpIIuYZth+AbRto+Oj5rtwROy+lb
krM6Q8XYcHRAb8wpr3paiyBiJwPH195LlGpaQFp9hW07KM6H5B1T8gl2Pw4tKXLw
dCyqU4rngN9TsLXP/rtYZI7xCNde0Wt9pWvRI71yzYBujodLtuM++q9ANwMS6HC/
yipzZp6pzz9CQVa2DUOKeXhvMXTDcz2hUOUotRmxV+pyCPHPLmKUvGpExAPpc7/P
Y+Epdont4ovcZf4m/1FFih0VX+UNpzS7aJGLBBEBgAsbrzxyWp+q3qB2Rtv4aFVd
ve9AaFwN4mGEjLXZJOMs8Y9evWngxPaTbb1HNvuSbOIpQGZIx7eAILcxHWoPtIR2
hNezyasfc+JhDEJhpcqnM51/PUA9xFlFQUNnLuuo7hc5d2tEWovKKp9ygkgav14t
Sl2+p9CroTnrEVHHcHXjQc9JhMP6ZByJ7Qo7OxQeNgtMFY3ZxShMClJaeVyrALM9
WiMAEULmw8ZvQ2I+/fBoForZmda/Q4KXXGATWzh2O9XnbQFjHSLuRGsmNQaSlOb2
j96HR5Bw/bAVvAqBWWs3tVfQK9waV9rVe8fAxHdNftQu7EMHwwtG1nAsaiG7bnbM
L40FoF/SERINuxxNwYG/OQ25azQz7WdQEWYv/PGXQ+wLCfKS3J3ZXVKtROr6TsqN
rjWRiIaUev/NbYGRimH+O2bECaMfQE+qpz+OouWsxQf7pdprT1djQVn98OBSy0q8
vEFJS63M0BsQboHE6xkPKbj+T/frFas+DiwkIIYae9MPZuQ8OhH0m+TZo2OKc6wi
+X62LvgpvyRwJx5KkJbEf/p76ZVSPoz8p7swPwN3VUfnM04UjuGrDldC+fzMF1WI
ESycGImeyvxJ9I02cr6oSedTOmzLml3AN0ILKSIjgq1RvR1PTeLTLWOAG4xDS9bX
TLT8HXsBADaHjpS5H9fb432hbUPmf5c28EMDTn28wWaTQ1Uxa8cF30dKXw+Lj1/M
gfSbWTpmy6eTpBvfObjhUTqWYjLbyvAHoOpQQgcvXZuxnmVvlcZX1vos4cy9FuOp
TIxJfliyomJimZE+FIMZW+D24BTAeTtirjzp885yThIO1ybHVJy71nCjyBfYLzDr
Qv8LkxlHKJn9Wd2bO8XjwEizRFEfb8w4VNoRS9a9Gr5WhSuDZZHvlxnrWskiIsUh
IpBqQ3iR254CpqEjGIcVvIUjXYKFO+O5ZggQv25Hft01pu7PLnt4d87D4tSHQ9nB
APlQ6FRs8IdgO8wzw+0LvoCmQ+E9COQm6tYIpV63G6t+VGvwSXKioJJxniCcBrHR
RvEWg2+2r0EcmkR1fGup5YFQtL3PlGWqturGh+/wSUxr2H8Rrd2eoiAaeXAl45XP
1OwuRCW5AD4bXl5c1V86Q8+5uLNTN/8XvSn0dK+OS6OH/Goq1fAIeQphwtPri18Z
wKxFz2V9iUpEMj9Yl7bsFazvf5o2r7/6wQbzA9iEj9dqIdgx68TYrtt5BHu+1nny
mSCFLl0LYsU6soXuFfJP+lmGVNyqJzbYBpaR3BXWJTTFKEigl194HYthJDb9u3QD
UoDJcSsI7lNanx0DO+M9je1rJf61kSPqu8BiQmolqyzO4VbRjVjKthMBDFNzqRBt
wBDZm3SctiHUljAjwM/tEsbswH3NLTCeZNxgj8wy/Iut/b62N5IAyOZeo85SY9/y
iiaJHROXT2Hs2Vo+Gh3zGlTaXapUQYWYb1gGBPS0B3UdOf3WBOUbgwgbxLr5lWEi
C7gyNF03ew9Fq+MykXE2IEfbUxuNZYIykBlHPyBJjV9YdtXgnRuoF/lc7Fc1ltjk
dH/f8fU8enZJFx9N53K+X342eyniIPan6M63qR1UQQwIELDFpOfExpgnVEFnJSQd
rttU0v8eKzK/FC5L7N81WJ6DX3bfPbiE3uucvgbnaIVIWa8xFugFG2vPsqDh3w42
huFXCzVC3bg3xnlDkRaunU/CJXAFTJKT4A92Nj/1FLrj1gGZuBgWEh4AVeXkJrhL
uzM2hygcLXMLYTaN01ahQbaGz2utj3Zu4TlzoY+i8xyp0f0t9oTnSW7pH/sBH+SZ
o55G6lOO7DlJHLSNs2y1BchzFwkh4FJ/9wcC6BvDO114UH2R4dv9TsErLUhbsiXw
Xssaw15R35ppuilWB9/gHQzFxPDyqUSQY0e+8mUkd1GQuZUfA8dSpRp8QagbRAuV
grJzvvqckd+XDrNwDrSKbry/cvSloigvjjggOA9N21dP1vK2FUKbML2idPmCak7V
y9SjkBCGVpJIiJqJRKFnvmawL8V2zcZJ4ipBLNewwZAgn82PFI1SxPUaqEp3eol/
xpOo1gWGiLm5n5UDDXbxudVeYZMSqjSBo8HIdLjhX1UYIq2CnQTIeTaowUIJed+A
weq2IzFJDdH95Nz9wmqW8thZ56uGDVcDywlF9xPVEIqfsjif+mXVZpBIJs9LpGvM
d2HEIl+AJx2gU0XmzywLCmSxogwd7wR8dR0Xhwx1GNm1ukhLpUCAHcvMlw49YdK2
8Vy1Gxd9ghgBbND+d6+G4pzTjrAiikhJ0GY9iXM2swwe8yaVzvKp1oUd316Xe/Ku
g4fPnNlfMD0NymKp4adXK4ksR9PevPPeqNV3pqAr/EeabfwzDb82YsYRhmNg96oK
amD4VQsztIRwWdzmaww0w1cIqL10b9opbgU/5ujf7roOYUyq1x9LYIQGrCdNiE7O
2hP6bc+B+v4wZ0/GHVnllLAEpofXulOwY51iX0JPuIuZ2xFKHPTXf8N3FpbEyaas
++9boRn2RQziX2o4j4lQwrBuQOF2P26cD/qQr68qiu8I6CWoAqh5kI3gLK9wPMEg
8xpKNKKb4WiBYHc2icAqj0cLxdrBbSEMDQKvegJkyL2g+mwzxpn2uoiDh9QkSIbL
llJCO1+/xkNwQ4Q9tUWbUAm4MZ4lzMHlThu72um859fHmNKHuh6rXVwmWiTeSfD3
yXGfJfbIxrwQX8s1wTZun5cAkfIGg4cBioKq7tdk1r+GRLaZLqwY6RnBsmOv+YAJ
6tOYjNq01+S4cF+FptDi6Zj1pM9Q+PN3SMzgWdjK0m3/gUXfQGths6gnJaOHFlM3
fgmpvyGy2FsUvmcSl9iu5t99G2COD5EnuVBXfnaStpT0l8vhg32y/U/i8LjPW7xv
wzpJDW/0pGkPQAFcQZnrfKHfF5VdFqMUAsW7rtY1IEsiHlsxuJzeGeC3JOHcPTab
uOYqiV7CkLQYmmsL9kKkom2MStGrUo9hZW+m/DeQL25D3048q3xPmk+a3ASubV/J
Bw1LxH0z5pVUyUieWSLR9XBHTzZYemxmz0eCWxrfU+06dKfKEYs+Y4qe6puH3NMZ
pIlAv45jdg5fpxdTv2RNXeltoC3sK2DtLIz85mYBezD/OfVBDx5HZ2QVE7GuE5I0
4jY+F58GuBCRkeIT9lGg3XefqfaHlRXPSrA2DaFvd8DA+0/n5qQtnSnX73h8Ux1K
235GEEmsqAOQaKnD3QwjXLPsTVImVIUAeTAWZd9Zg3gNClF13K/V/2r9z8dnj5wG
1Dv/mq6NLLrloftJi9gU23K6DFNXBDQj0Vhm6c0I9/kaFvV3K4lFB+Jw2aUDFRrP
8n4T/TWWXjxNQ5MUD8WJ1/RBax96zIJrRqbHpHvF1/MDz5jWhz7I07GwLShc29a/
X6I/j7ZIvuUJOOCIrEvanrflsMweY6gCufEblcqGB78s9YZu5tcb9fAhstWfSz1P
5GTdtNREzt1RRmvE93TIByYM2Xsp2GKnTEKQzfwPzFboZGCqAZi+9VJPXUB8jU/b
BsDM8/RIgMlzPsxI1XHirbBJhv2uNmdoOvur+6Cdc0S4j7g32z9tQRGIBZie3QXr
VEOndlG/Xmqn8hqwI9HN8MbsTGYrfPkXVdQjUYMto2ict25Bj26xb2aErBtCvafg
DKxtLTBlxatYGZhpJ4+HCNTeysbtmtU7QTe4tvxR0OnrcaEKNl/EAgzc28OmaV8T
wotauDdpxSgawLhmfLrAVfKnmkUv5VOJx923U2LRp01/kD3RysMJC7BmeW3cW1Te
MrmMn8YsRfGV4wSvIlZIDPTKzGi3TnsZQ1LHHSuRt06fz1iHfbtZ5x+I4xlhNOpU
OA3ixI34YBmXEhw9jMLZ8voTg6HzFLU7JiJ0d6G1cu5pJbCU7k7KR1x1EKJ78mH+
5zhOnVxLTD98+WlfY/1dZAXHWLc0DmNNwWzlYvDHzSY8a6qYUj4cdDYyn+YiKTRq
y7q6DIHw1yRnGzNc0c7EIfHORdkDN6D5kuJ0VDIgiq9ScOGGthhCrLfWf+C4D1Xd
YSUsacWLifs1XFytF65DfKiZHW1Y2FQsGgPX+gEjmGUX4vr/T0peqRlopiVtAUZu
yFs1yW7nhvToM2ibvvlO7IkykNnDWL5VVNBpb1a4kLmW+LuHHWzM1aR9dNEVM0E+
P5beOMUP/dT90pzWPaNyDzTD6lC6P7QdPR1dtKANbPXDZF4lbDWBN5ceaOloOwwH
QYnOCvRoFcccdgOeqBdPid7c908Oeqgd85sUKMI0vglvIqVpR/9iuICjNkXpAM9J
kbAcJ0pWBgglSdxAcJ1EXtSS13ot6Zr2KWpCpuNohZ0JJLpJ34yeOBcf3Mo9aCzM
blmgxYBgcmYhu0NB1nHKoRvXadRDiGvHAAHdA3HPxzeYAkQVrxyI1tmp4LZp3b8P
kKGqI3byv4C0xj4ZtqatZHh3lLtiE2SlfWofIxIMkqMjDUu8GvAy1diUQlCmzcUV
NwTWtpQbRY5gUbX13UniKPVNlpz2ugtMMK7o10X7MOIG/LGVR6PMSLYw2QMxG1oL
q1CDSLuMLQdztfcsZrxSC2EWrTo8wXygZSU7RKAfVD28XKxbBJTidGZptgr2uDAP
GsZSEv2KIoqrnVQokNeb9n0xHsN5feE/DZE8fTOs8YozaoBEPEYrDJKJo8M7V8I7
ugxW0xkF893gsoYYdhIQ0OixjgEiIMBTJqECun1hd8bRRPvpEBcqbq+Qwkfida7o
9v6z5v982FJfLAaDxYj0+E8xX3EeRB7z8fFAj1wP7emaGU6X82PiYXtYcxmgpBcG
6OOatIDc7tJkuMtGE/Osja76YQoZd7iXCgGaVK4TG6TAS0H0i25T8OQdLxaKo6q1
K1SbAkDi01HbiDFKh1ZPZHB3yXtQxB6IYe77fr8xGBZeMmIjmarbmVJhRyJgptYm
1hlyPQ1Evciv8wMa+gFcwxNv8L3JH7wRYFslwuvlYf+9BpfI8ILX28jC3X37tKO2
8uIrEXGhX9qOgfBNQJV1yEaXGD1yuyHy97lXTvQGDWu/tPfNLgrf6sPI8ExaN5Ow
OENI9A50yakppHsP+kr/Qlu+5P2lxxfwxaIDqR1sDaiGnqLEj96x5VSMv/kiBqWI
DskmpKz9jxhj0z+V0smE9aHcv549jsUiTIq30fmY1irQV5KfMnRyh2Je/ZqMiZGf
uUtg6VdTFL4yE9z7ns5imiBiEy64UNtx2tbiUxljwAOijISlOEdej52izmroarhJ
dhKy5Q+PCe5KryK137zAYv7vJE/Ce6pKlQYIYnNCFflfKUxT9b5UTJC9GEYJ7V0H
ZB76Ri2haWOuMOrNJKmgKVKD0rtSnAwGMAorz+nu7TEbwt+sEO11CRpf6w4sS1jK
hpAOcv7FXEnTPJcdA6xjMUmAv2qA5PN/CdxHoculqNAtpKeFHg4Hbk2WhwBo1196
KMkPilYixAe8KzehNhwIrGP89xc8xu9FZYpdlP9aulp1d7dYIlPzQ/aFIgumwSHi
qSUL9axS33V9Ld2ZTQ9pBQITMJSeXW1CTr1CKGi+JA3ucQvlTj0DKvCO+rs8Ead8
tsVcq1/UidEVndOCscJAGHRdcwHq5MR2oOCrA7cH1x0A/lTLoUcbj5LDXLCTp+Br
dHcBI2pBQKl9Z6/dWj6BtLtQdet+4iS24CcbHuxTHZbuQVQqCCKPc+0qZ5dM9IkX
KVR2kSmkjrZTbQR5sE82Du7Ok2klKENuV0T1+IRixU+7ri2wkBvT+i+uG/csaikU
R2/KE66OW9pvKhSIZ9eU84JVHqEyUYBThTISd+EKPSq1+ZAhVWWEb17fX/mod9vq
nAjGZ353HqU90KIA4UA8zFPouCmBzJJO5SvLN2bzDibHec0t4sdNW7Tr4Qn4DUCI
p9YsYeEydQxGZfZg2NbIk5zr+5F0+jHyT8/LgpIXK3eSdf/Xvki/smiwt7Klw6Vb
fYye8oh6GAvvUyCdUOgRKpXqtdT22Pm9xZTH9apnUhxt3CQN1rSQ7Cb23O9wnrxo
8c0w0FhEcm578biayCuSctm7Nx/xFRH7ZhN48can6GuMs4NZxz9/ewvmj6phOIBG
vmp1yhwRin/scSLopjrnoYUvlArm2Fv1xz1KY8v8KUMPYMzVVOp+2Mio25uzF4yL
D4/XAAP3ifYXRfn5fA4CPHTAhM9sKPWnSa7/dDSwLCtaaPA3QFGgKDBtqWCARD4v
Sq3y06TRPLcZx+owr5yPrg3a95SFxurv/+LHwLLvHmStUFdiR70QTwnMS1t6urjR
gimYP0SJrS3Y0HQHNKGe+k+DY+viiaDf6AlKerNpJa3SxIPobm4XINPY2bdMp99N
4dRESd+6rOk9spLe32115e46gEN7tv3H2K/7nL83G51jZJdSNEc1nk9v2cRgHyXr
9Si5rHMqobdM6tV7BUl04W/85klLrUdc0PSkDEybJAFIOz3ZeUuBWPnNhf29BDIK
NvwTugshZV/Z6wsy2734tL/yCkNUMeKyHlhOtaedZ96i+OV6u7BF5MmMDnutctow
H0W9LNswH3vnqfCqU9tjLx/JMjuxpVGJ3HBg0e1XzWrcaZN2xFZubhwLoWI07Nes
YSAaXhuui8JwHIwBrYIaztksnGQrCcRBxBrgXHQ+S6fN4DH2ikkjzsqwwHmWLKvY
bpcd/VVPcJHDLblPumfBBOKOGt0cPpeVh9XY9nROXgkmtOo9M8hTmfu/tSClHf6E
xRT4mO6GPMuG8wGz9ItdmcfPnR4QvtmLKSvMP3nWRLOGuNfp0C+D346wsKuJBYNF
qNdXnxsodJoBEWaz1sN6F1wgaELuS9Sdb4u+uVsRWN8ObunVUneFhCK1xaPNAZn3
bqm+qrVrjxZLrOzDVzWHNwezjgfQCuUeMUcc8nBV1EKAjrJChOrKiVLBfaVI/BXT
M2Jfuww7aeewXgpUuMqRpFI5uL8DuSwVbIugJ5zZDakALLz9LdxpSpy3AGBuJ28k
L9/L52jQ+4ise8n9FzTk4QmR+trl5RPJDkIbfgoIB8jYKSVxwGYSsZSgqxslFPhL
Ido6apDOx7R95OSmMVpG25RSZqGR4nC3eFvcykjP+890+AUo8wdKWm+YczNpcQKY
yWshcVuBrMDhLQksRHPKrX7UVvaD78ugm+PNW3RnPHTAdw2NmBwL4EZcsPhi4vO9
Ond/0wb1q1d/d/qFse6e+R9S2envAkWOKPsGiNovNLphgwt4nBZBdAquSqKl60aa
c4Fe1Ew7HnxIcJPLc+LytwOKgH7OnGhnRX+iPiJCtkAzYGAiymkWTJHMvdZisRpP
naggYrqNwaSr4rJu9ybXHD7it8OdXU9RG541MOEwDNCZHRtxljgSZc44/SwF9m9/
BVK+UJhYuEIWbupo7m6RoRpOALEBatg7op8noyZkENfVDWVfsnzheuHcz1Sg3g/A
AQei3BKCnnKodIZgTzHxBfYI6salv1Np3ZNoGJgA0iZjUZfjqsPVFZt4bXX6BrqC
+z9z15uoVJJPGpkees22SKKdBlUV8lKcxWedE7KrDh5qYexl33lNXIIxPCP0O0zf
WROOfJdpjwgR6er+RSUQXGZFb5qylX4Iwv8vp9XhwOx+wQdxDgpRFM4nunlPfqbm
S8MVpfEUa1kzDa7h0QtO6+/C70S564AJIIUQs29IlVkpWwpbbZQDaHZbX9qnz3ts
uMNvB8GqPBPxphsIcmjaO1kcf2OVIME29nwh4QJlEZk+U5RoJ3XFcikmOwuqSvLl
yW5uf48SrbpdVXEs6xKpXeFelC3tLEc4IrlaB3xj4+ym0PB/JsvDCIO48W+0w6u0
G09poTPCTUfycTfLvjawvYwk+ubZ/oKqtm2peo7I2vsfP7QhRQ40Y991OzDCvGi7
MSlyjFSS2fqw31IjedFB0j5mePmF7cRoCfjQxVZQp2sZGiH3oWdGfKOy2F0mg2nM
laPWV+z2MclNWfcstn8uN/5aXyS0wJ6eJRKpYY7odVF3VJ2tc6VQTh4v9OfmDHZz
+4YCc4vGt42+QZZ34zbukjNMPNox11xM11NYfkk6S7BuiBC2OzWwgG7vfWfJx+jj
XPmwIgsqqDrbyz/fNlqyxgMxEinzamu1twziEtZRzCr+gYnxMOc15iLq9UAAEf28
+l6ISyos3sgTRdkBnjbV1nqK2Cu1xHFZDC6eYHp+tqArQjtShKyjcZhIgoAwH2/s
T3/gOINv1q4hr3r6RWNHnzzjH7rfC28RZiDDqJP/NSUxoigc5/9SyJPxJsO1CyZJ
fv4s1q96wX//7tCsFPPtQ510Hl3dRqfrmo2DhII9BYz1R1+DiMVBGANuF2/mf30Z
DaxrLvppZ0mbtL3iPLKaxi28YaSK9wv0W3S0cCHU8zf4BdKVOjLNNz/Cr/nUcLfM
7drzIU2ETk10SVWmdn3UZzI33DubCwOqmy+Wdckpec8xyjaGYhWriEZBBfqflM9x
Cc0/xlq60b90eokN5aeRYlCS3Q+hmMED+BMJQVpjBC/cJhXHXAvAU3TaxaKb+ivX
M1DYybTWXpZqJ6VRJ0AnSxiiASsylBOYxBea9TMmhd+naYpIpIgDo89wF0ED6AtG
LDbo0SDIexxL32g7GDvEbfHVtDoJpk0zvkiLzUgiHyWH4klPhgxGGO1Buul8mxwa
BL9uNSTvHfuWjW/hE9CFvhqruhr3IVUaiVqbZZGXX4gufjfjMjo0d0w0l43O5tbg
IUED8P1GJ4MEWMxuSw0dic+HFDqjgVFRpxgJaXfALl/oYMx3q5m/kVeWVOCvQEV8
81FCd2xJM1NVRnu8YWTSdl/PIgScl4qkD+VPhKN+SCtc5zohunoSoXJqfPFUv1qa
wN8A+yWnigfFOGwpqZ2S5dgAaSV7JjY4VoJvPZMN1szlSaJYR0GQvva7hl3F3VTV
QoxuIea5Fw8HpJE3jnA2qQpa01daN8AlCO+nqxkxaFsrd3LahhTSUQ8CA8ND8TOA
ARdcb0mYVcXzJAuUACKTOd4SfWV3/TLioLEC+f0QPYwANKdjpYGcLZgwq6MqzDoY
+S46n5tGzYrhRhqSw1MQgoskYx84LNoUxBg0ID44z/9LwZHIRDoEaR9V+EBeP4iS
+dX8pTSXPCOTAGoXYDK8vF0s0vTnNyeu756uh2hnHL7vQgusXYOLEccfMErsKmLo
NExIGKxYMWyj1buMyyKk5Vw6tWxGeevaVYjmbx1FZmb6AUvL1EtyrnRJbBlyK+Fq
qFSgLFlO2k8YIL2aPAsyCCFKReIp7O7yrgtGhZXLYNlsaTC9r1ubZWwzt0LBFjRd
FXR15C+1dxP7N1+ycGBj4WEoHXxd7F2FRlOYH74BOb+n89MUnlngBmEtPXtxTt7T
0PtBq1toN8mRLP/+Ho0TsDQkBE4LSswkL5dX40g5rbJp6Z9kc4Vw6yQt/uVNpReZ
7K/L1WRf/JUDDa9Lc61t8NlpQd5SF9zMov0LjLQl03SBL0fTJVNM4A3GMqQVRW7E
ESSu8xsCh/bbKj/wK28eBiygQy9XkmU57P8xdT9A7Gkoc2SQD/SrIYyc42yqVYP8
Ld4ypuJ0DhOi4reJM0ApeIjFHMT4SUclAEe6+SJ7fa2eJnZ8c3Mqn2uxG86lEVsX
WwTubPv2KTn9IMozVSVcGsZ0EY67S3i0qtjZWrU9fhPczJquWFrvdEyWmL9VsCRA
1/9kJMRAJBG0zl8sgyMwyeHple1QJM58D1jFanRTVhBg4uyQm/ciqZ1Tmn7ILyOi
homH7wtju/De2Livsgyj0eRaiED+YcdopALkcpQhiZCdcENP2HDvsxbw5Z7aR61/
sGdP89hxVkRx88OuqrTHWOa10/D0doMkDGV7H1Eu62qnmkIwlqKwWjTefEWRpMbe
h/Z3YEWAPtGtfkJmCstF9Ri9gCuxMa76YLdFABPsKBXGG3oMBfgi0eSUeU2tBNiQ
idd0yc0FDIVoWiRXdjm7k6F88yxD2S5sbZYG2aLH/YmGZSfHU1K3TbElx7Gkt/gf
nOEy8iSfiazN3hRa7jC4oPmXHa0Se0N1GsCMSoxlCnqdngSG/3N91c/Wc670EXcq
k7Nd3fZlKtXAoUfOLbSky8zqfj+BlDNG10Cahx5CUEp0u/9+xdb62ZDXM80lh5Cv
GV095Udy9obAG/KwsqJzyl94J0YA0Cs7roFNL9RrTfENv70cp1CYVunI2GTyyPAP
EF20MdzQcHwIia9dE3r4EqGRbFnE/debSBd6g3kiEgaMBPnsYkNqqerSukmfaQho
aV0z/Jux83uon0JJeq2V9IQL9HDTb6+k11ObjPo4jNlc+rYr77jJ497y7Q7JRjA7
W1DSE6+YUWRxttRB7WzcBoaqbb5TRbmlVY2Xdtds2HEPiUVxJNFH48hiBIhCKBql
+2DPanlAqx796qqMs0BWmyNS1aRfWhKGDH/QrymcWG3kGRg3L5gU80HcKdtnpwMN
JoOveEDxFu7FPw2ONeJpeTxv0901TqioKAQtmpMt9RfVbbe+vyYC6y6zyrTOaqxo
eAlyvFZfeYzKrZcPXkcuk4WoFN+aUkk1cWRRK7qb/ODjT5S9FFvf4m7CQq2CulNA
3Lvrt5OQZQOpuf4WzH+0bLpappa8oy0Cw59ZtTUBq1OrEAAHqgMSajo+f/5JdEL0
IS1RlXFkpP4Df8Rj4QeQp69gTD4dcP+3ceVJcQjS2LdL0gzRjwIkDz20zksb+kjw
UWt9CtZB5m+aBrZ1QXR/DwVmSZKekiWMdQ1MV8P3mEeCWYjcZkRHocj27ntiFj4e
hTPXxoDErp2/Vz5yfQGbmJ3R67y0i3dEXgf0PvR8MzancdJGukXnZNBlZ4Oo9H72
G2PSe4STEWLljsULgJentApXv2tdeAkK0wE8Ljt82VTJXJ3H4GdBuBn0Sxn2foaF
doyC0DNzAUNpioPBkfFS5F3djFtHM7SIc3pPokYlasm5/m6FQUOHdoUKqKItkiCR
4TPTmnXI9lLf4B+iI00ZqjUeL16E/ydAzHjRLTgoxMQI+s6rpDDA1XkpZQt2SAyw
B3bhuaC1Z3WwIy31FOwrpQHHqF81f1d6QmnlNL/EqYvRVIy/3v+52a38rnkIdAih
SWylU2kLdtNp41K/J34EzFNBvSIBDy/A1PBOXcI5EV8bA+u2J9ksE0C76lLiFoyV
PDB//DCCkmAlYKrim7hathTCk2SOcjEthZEPaH7jJyduT54fxvU1Q0wLiyEbM8Qw
DYPtOfpdICdW279HRTBFF1OjIF/p7i7T30tZzUH9z4cgD9U+JKiC/Iia4OoxPhN3
ytoYLOMVTD2q+fh7wsAqHNOgIECYeqiDq2N6NRkIxGC4dTyUQTQJqxmA7R0urHzi
4uZcb+NsYVPWCYVeqejrPVh/meNYy4YNK8az/KiTRo3FWo6yPgWEIjssWiG+Qlnw
yHOBO7XFENGu9BQqevQU6gtAZXyN1W24/u7h6JVBegfH4X3Ft93FjsRBJ7ouK8cW
XqDKajNUpleUgZJhG6eCIwLU4vMzN54G2nNAX6pwqWURvzroG+QymhhXjxEQ2z4j
IgJLPj8llq81OO0IQZ5QHNgY0HmGH2ppCE4RfuWOlqfT6icQpwMSwn78A966PO3X
qh6rKU/0GVgsoWSZBx3DX1ph2IHx5oVLKWFSU9QhtSOS+yFs6VU/4p1BH9qINBrX
07wysc/vUy8izW1ePUtXZ2PSAMwmCCZZ++zQk1t113S5xvaRTTXKnKADDq06gmsb
GtGz81P5O67dt8XfBBw9bUsgN/PND/DtyCne0ha2CbSANUlXCyFpHvxAE7U/NONu
g8M99lYjNC3+EXWX9y13jF1LZqQU+YOpfjIOQWdaAATzKr1qVQ2tu1cPJywzSnxw
+524YCJF62jgiwb6JWKtCi3YCeQbEXJVptibdAk4WyTrKqg+IpJgyqaFRKGqqQAW
WJJ4YPNfcO8RqSKgy82A5evWJcyzQssjIz61zeuDDAHPtPOmds5FcHd586KNo1wR
dER3Iaz6Ul3p2Ih/ep8/K/LoeUCBIM0jeynU+va8UAZtiwcsG83hagq34/v7dGj4
OCYXLtKY7lxRIuTLPkBb4uhWmBCe1W1pWgesb4CQRq8gWHurNUVFeNdyIcyFmb0g
j6LcF2GfvgEGFQyD92nmiqxKmZkHaK2x3Zdyr49DB1l+5txLG1qeMN1kTwm5gad/
HfDZuzhtLZ1IA+/m4dmkuGDmog0KAXM3DbIwK+vq2/SswT4GJ8SoyhYWej7YCqPg
ZX0YOi9IkLUwOnVOMf5nVDg+z/N9hcwOTh2auJ7aach/F3I0wJtC9iN29SvzfFtJ
nmTOsVZUIf+MOs/w3XwRpiGOoZegLS3j90VkqvNOxfE2fz75hXorCMfeYpj6i9Io
BuOPWDhT+4qfAjGzWbqkYBXFQqYd9MbAWhYPl+/1BNtaIx/6hec9sYby5Mne5t51
pJp+N0sP7UzZshDjUq8hA+WXJT3TjRI28UPAHzgq6S4q9hBKqYA23oZw8mQBXIdj
6ZT20Tg0ZcvlyRtKmdGHC9ZP1nNtgL+U/CvHn+ht+bqPtZE+QaQtcuZesmiy2XTx
blrvsi8hZTMpPG7np69zdsmLHtnNEhclZEF0hx+B4LFzPO4EAOdvF15vcdPLYXbm
s7yRVX4rxoCNSdUTwEO0tREEitNpFecttZDdsDvXxpFlhpnJ8nOsaPVM8N4pjr0w
S/QUlkdY+yhUJiudI0Kwf9Lc8tKZ8kdxL6oT57+uhuLix9fGesfga4Hmn0xml2Lv
DXTF1jdYDU4i4NtDpzlamGA40Na4Hzhtvvu3kvQEgi+hDgDzccu9WSDwltum6Y/p
TDpKRXxsvR6uhKHsu5kGnIuY5mSEqEh8oN9z9rVYTN4A9h+MucKr1bU1QRoyAgc3
3v14JujYyFTa/LpdFuvbkwQOzsjq73PTsOk6nQGz+8ajFkaZTy4AprZjgxuQYUQg
f3PbHQT4kEQ06bSDgm0t80bEj+Duykk+GvZtMZRdR1PjgxL8x57TDk2ewkGtj5cP
z+1wQ0hqKWxjby6gzOhwCyp7t2CS0WXw24KMlnpJpD3wNiTaP7rpvqzCSXXf7nOS
6fnrAqCW/QNf8RMPYLhCey/xCInQ6//BuCXGruPGy8U4k6o97pittDlzX/DaQjV0
Q2zIF8+3JeN8m0YJnm2y5KdL0rRqefYKF2sI71VjQ1ZZ5yWI90/aZtFGA9lsn7RF
JhsRbr0zeC7qdspPNfzwMReiH8MoPsiXc+pDCFVIx6UEaKsA9dcXVCxTx9s/iQLG
Jf9L2IWmuOp0xdpTKSXhguwRNzP3WtleSRbkQiIEsfl4k0oTQqj3wSSjvY9WK4a3
ofUtmyhGP0wLcNPe89lM35zjZFTs67ud2/KpOf3LnbE7t1FsOR6aEnievl+GurcW
iDhVBXnDK3rAydDks5XmfDVbOZS9i8QMR5U1zh/aoiH7GTVxVZex5i4B+qEe+cvE
ulu1MxiSuK1sCkhAo4Fx7CnOMtthJ+q9rcV8BpTYhzVr94v2HC8xVO3Hpi8hvdF/
2rYBuVnUYN7m8Uf/5k9dAFSzNDDiTs2Zz8YiuUmht9pZE79VLsPldqCnIy0azy8U
F2ngAeqLFTlpc9+Y5IExhX89XuYPtVtAAAWWdFGeGy8J5iw4xzyvXEozgRkkeghF
jiQMUQgqcXcsmBbjQACIrm2/br9YfjIphJr/Ql5hYLnN4HM2r+eBM4ecwRitmWid
yyMHwGefm/xLbGzfRq+6J5WDoD+xl+tz+6ba8qzA+f78Ty2m9bvb1HIPYExnOCKQ
di7ycqv2zovAfZP5zx8lOCP7mBeBH5Qxs/IJOn5hjkNiQLwiJOxjlvW/9JwEQ2DJ
TOJWCyUcxoxvYpSc2f95hVIOuF1AxyNRviLVSPgfuDL7IMcRBwSeKwplO10WqrIg
SgbxiAIiD5p+Sx0zNFEB86x7rk+j4JyMyxxDhJlALTiuUfnZWbyiQqb272YNfDJB
yINOOQ9/80lAcAmQ+Nz+f+tqKp+Sv5sVFP9Ixgsvnyg2ScxDjW4eFti9MnJlnWpN
p4/59+jN19fmOZGfUqzBijsjfQoR9n92avAc5BHR/SeZ6JNMkcYCnESemq/f0npQ
g8/+izkAtxL9pcfVHlvlUnuTJWkE/VlkXxLjgGRAbis=
`protect END_PROTECTED
