`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8E9uGRazzizFG9Zmy5ic37q5/R67MWdi4IuqoCYouBIUa3dwru/UdmQcSt12iNqU
OHHbnggdSiJX9Bjw+Eg38eEy6Bx9jEzjUapu6tQegdCyMm0KDLv950sqIvrXdrcy
K06XQkHqZiQuWwYReE2iXzEo76Cn3LjWRjdKPwQnt2mrJ8oRYQYFFvQ4YukhMJnn
7cOoGQJsNwxQlXc9eJdM9my0BrbxnuK4HYImsWMeb9+mYLIgv3s4DnVc8lGc5XIu
0SMnob9yCcACkTfcC5TNNyRVMfmVmEsI5ZSaPBudP/CSKGhUITW4xKAj5I/k6Htd
gHwe5mKCw3ZEFR6RTe7nvq2pP4ow6oH6NyO7zmhSJZo=
`protect END_PROTECTED
