`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZXn+2C38GRrLLmpwLnLTyf2gmFs9bioXkMsaPjqWzc0eekhQhbXt239YtGwLPDV
g27UMkgplwlIAIvde66Oj6t1t9IjufrSJy7ShjRzKgCQh8K7N+MZPKKCPrunDdhi
kcda6LH4/4FA0HOy0wC0eHFNb4v5GXtO9tcqDHFUQoYg6xsHaQK2i/ssKx/K30Xi
rs2rO8ZPION5Y3yk6kEe6dc9VdcELX1xUKzNx75+DkySY7WiHZcf1YyYkE2qIpdU
wDy3vPqJRCDvPQHSoAxsqoSeg4s5vyamthOiekOX2jWh+AA2REym4uxPS13P2aLM
XVtDpsBUQO/qcMl0mPBenvT96fwpGGNkGq3yk18aWwm/45r6juIUr821X0IWbdW8
E3toXnkC0QUjYbTKckcycshcLuSWx9e5sANAyXSWjZyYLBST70aGCeqY1NTpSQIp
DIBw4ca7jxD1P5XkMIG25KUf5Si2hc1PrlFkLJA72IVO08yPDGzdCVe/ZsujYUUV
2IHUz9Mr9wvzW2kFJh2YRdTxbl2MjHJVVRMufUnwuDox6ORAPmtacPSIn3kGUyI4
vWfFLzxsXWW7mUvipuM6MbaPzmLgiFMjWkulpWJQhK9zeIBRy/ee4X1QENXRH6nP
EuPlc8algkDn86cKHgkdRg/6ImRnTxDRvZ7MhDHRlFc+nZt18YVI5gPM14Z6rrGb
5mMmPE5jdGIlcUFrjU95+TYVHflUQg0rj/Sf0isay/s=
`protect END_PROTECTED
