`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rlakb6r5ktEZq9eYPub1DdI8CSNHOIcxWjcA9HI1PkANWYHy6nwemHSztzx+my0p
c/MJrgbq+a/60sKuChH3duI4CwEsHFNS2R93EKq2uaBchF6g72yzM69swyu40Txb
rrb2mekVqfMWlwTMwQC1HUDAB1KkdMWVNP27Sfj/RalhrR+mpb3XQAlcVO6McF1g
zdo0PJ1RkPpDw3P1SZMzeup8n07DafHYNk9X//5XeFqdwmgQRADdCVZgGs+JMTEz
thWGK3Bx2oFamI8s9/5B01I5MwR+nm7lpjeNS460hHPGxFWbfBHQJniP2i6u44Lb
hOYN92tF37l8kveVnx/E/TdZMrSD8y6B0TYPAyFJ1J2l1JypYlBM05wYt+cwf5gm
uB2zxc+sbMM4ICLZsPi5zY3hu+7V+/n+Op5a1AMEHmAFMlPkoUYCNKbDZhQlRU8o
sL7YEZUFKg1biYR2RXQpL7UU4ZsHs+Vxq8kwBEK5rWMwEq2TzZIMtIADzim/E0Q/
jNOo0XgYFHesvS9sPH5ry3KBKRSYG6mf+yejFiaI3ok3K3uQxkDBd22il3TeRVpa
+qaPEcQpCuYx12JuHNSsX1HiFCtAqn806zn3wPxEfbbnM/0MeQZiGou2P/RSYnYW
isyCFRh4ZVwCqgk0Muew3l0KNC4TlZsVtb5JUoJmK5ZdoKNUeOrqsskuoTwqX7vp
f9QS9FPE12GiL2Km/xv5IzAJUswUNn75sajq0l2seU80VrD4B6mzCx86V4jwQWBS
cZU4L/gYzzsx6fyF0HsUCWhSlTy8TXPSw5MT1g5E9r9PO3uGSOUxzDipw1PdtnNw
d1kv9a+a9vBAte2jBOwqW4cPQXRiqvFmPi+loV8U/pDsX5BglWnpkTfhkpMsd2TY
aufotWVC1r2KV2h2NJFLS7wJrRQy+xjRNwfCVtT4QGfRSmbAgQ1r6UT+TB7O09vk
GIywyfntOqZRjmr/KrSfed04XSFbC9uDhUa6VUXGNtcTTMl6mfZv9cdmEnMC/Tar
jKnrgK63l7l3eVglll5mp7ycdXB/paO+aekJ+Zcu8+dr0ZyTcCk0pyEFHFU7Htod
v0x2hZXgPnRgfBxIcEaa7PfwmNoiiAM4ZkNeyGwjBbFQY5+JCPAGlgU7Rd7xvGeH
hwjxdQr4+Oixn3lcBnZKmIVfEtlnjhV1k6PZC2maxaeTvWSAH7GC0y7lsPbv82U2
O3Qizyq/ESNJ1kcLFbZ7e/Bvz7X+7kaTRqo9+KC5VAuH8E2+F7ki3i/I4d88dSk5
BusNjDJWrM13dydtVqe2+68+v8EXdn43be4o31Qo/d+Swjn5DX/tpcxSnoBGg5hz
xqs5vERMQkMvLTThp0Kuv07J7mG4E9GBKgAt6oPit0c9/t99nSZGFs4xxOwfpw6S
/3CxSrq+YOgMKqHYgBrZ5U2YfK+cDHm3kYTclZGH9PiFc7yyTpgo7R7QESggMX6P
W0AzgFKGap/+4MksASj0UC0jyEaagC9Rd4r1wk5Mg9Ns2NHE9Pt6lXsduB6Sz9b4
OcZ4Lw6HQrAQNRPrzts4HKUPi8mJp6RYrNMnOS6Byu7z1JVZ/Wr3lLe8P/FzT6IO
Rg3TMUJM/Oi02C2PXSvvn+swKGyD8Db1dcBpaCYWbaw4qdSalgqruEizx6l+PldB
c/wc5iin6zR/EgDDOtZVZyI9PqTj85apB8viC/xS9ZTNU/EY16SxfanBXqF8vnwa
btPU9LU3JHKMQrVAuB+nwSup+U0ievabS6xuQbJPE57SN8nt81WqW0/c6+hl3t6N
GqXCn1b7ZxOWbkHP9jryph3jdGYPYypmNbIZJERgq0StEYTvYbQ9Ewoj9X9xrhzL
sJiuhaFr8nDFJdIL8Ce+WhZi62qgjNniUasyODXPRuWQV7C5avYBJcmyvS4iPycx
x3aSYJ8prl+RfWKUMFoe3cf27TPrM3fj3bSAyziqZBHm4cwwZwyVOPawN2jyJNOB
bPvd6Cpkx/pX2ApthIWC1GE4iKGDbvZSVXG4j3sbVzpTi1pRPxp5UKr+o2H7Qbxf
OPoF5NqM8Pb8c/7nubmFDc7gk+PoNTokWLXehXalE545XvwzycDWG9gmW1rOPJJr
oTq+zFDlk1/yz+Qau83v9gCoR0H/DzW0hhP8gApo96o=
`protect END_PROTECTED
