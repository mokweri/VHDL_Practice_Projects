`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IjeaEj4fwEGlJlZ+tDlItPLmjeOWNfuYAOKaJGmp6nRO2jrcnXc7E4RUBUWUylF9
6/Dk/qCX2gVktKySS5zmBf7xtspNi3eK5li9E8qJ9vSg627XLsYcC4N03qkKgKuV
xaiKfKy49eN3KRGD9hY5UtMCexZgZbOwutuz6Z6WD7smNPanvKWA/qTHCPW2Cn9+
2qrQTZuOyj1Nf9EBOcQ+nIO6Y80+2msOqdrKF4V+3GSzA18D8KHWLJ5jfpeusX0O
eRBh+OLg//+Ei50+9IS7toVRfwwQDnjebe200orSeJHOQtHnDogyUr86KWM+fuCg
2RcIT9Agps9zY3q+qYpVvdKSVho3JxPSOph4Qtd7AYRD1h6gNa6j7A0LBZ4se1W3
te9r6cxKCJRerqGR+Vfdb+VVxE3eNI7p8pMpr6RG8QHSYe79qTB1VohCu99lBFcv
2RvPwm+Ce3CwWRpBFJf+KFdx2EG5HqMu+jgufigKoO3qNjlzOXA+IHJQafQGkPtV
keIN6FuQISC8CekQLwWY2klf8cf6BCwzKhKxwlc8xMM0cLXlquecddEv5P+VptP7
jTqoYs3Sw9AcucGClnSWJIlJb3pTJ3p99aCX+l+08Bjn6bquvH9efKxU6QXMmjZM
0SnlyD2lWyvNk/MRXRWD/fCzeucuqfqCZgncsxOQSADfdZUT+SAmiaiOiIxKAfAp
IH35tyn9X7PZxaQRHPboyXFjcQY7v+Lv4kCiEyfA1VpuprriM1J0HzsQ4gw45lEJ
yJ7W/qUWaKFRYNB4Bgdej9XfmBs6DNvsUT5YV9tTtf5m0brTsLtoy6JuVzHmUZFL
celEVBfTYZipIJ2nblbt6w==
`protect END_PROTECTED
