`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+5H0tsaKLekqyeqR88q6YZ+WRfY04V6UDNS8eAB0ZhiVoITEsYs3dzzcJsNYuAEq
qJ+BYWWDG/cVXhB17ETOPDH5+wSQgdEgY6tM2mEv7ci62B/SPyHgY3mAlouWwG7c
tV6GC/RSx7KB9BBvlWDOkVs02+pRDzqFCCXASDpmCuDEzhTXPY3ajzYD7pHsDjiw
cQwl1EiNbs3/pw3o5Ww4uTGv5zei4oeps/hrfLXFiQAOqG/aVmYXeW+I6blCP6UM
4riMX1z5ywwb/hxthmD/5EitZiRMwLOzrFjx289hetgsWKNkOsmC/Eja/l1VjMci
qeAynw9BUqJxEYpIUt/NecLBSanUiDuhV1bOvFIRbkxAxxTTQiZVCokky9tPkPeZ
q60cq9Wu5iOq2XzgE8QCAS5dee359rb8F/uQlH4X5w4/2M2Ra9LwvvpLVISsFGbD
`protect END_PROTECTED
