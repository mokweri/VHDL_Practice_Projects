`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+aL468Vohz3UQHcey2bsmdQZpnNJtBz5na9I9f4MxslDMaRP7lZo7joKdFY0WB+
E14jiGEgYsjrCcFHaleAt/2OLKMXHUQPJ/Xds12YQ22jDeTsE/0xrY7yg1nS/fo4
UF9ExfG18KElXO1rYY/2OczTvb+gnFwD5dW9C+mUnOFynHpN7hm5vdrBmTrQG28E
LMbsWSNTr6mbWnDKUw8THXpQuX5gGTPjZS/COxuPfPtWC7sLYNbFS+THDeHZ7Lnd
00RlSnUyUAzW2cx5FFa0IAc2JdnisncI4BbOj5oA0Apnmh8pHqbdfzK5krG2Cccm
mHgrWZZsDdQaEsUz9r7cDlLlNaQJ79iEU4R0StWywrLjAHty/hIvoEDMSZJEBa+5
kuNU1+73+lsSZ8PP3d8IPs5eg295cGHc7ZCAZ2Fv0rwqIEF2YThfbsBBp1EF5TNP
U3t9NsxKYkxd6Z6s/+5NjCcuYUEc0C3m/rgtj5tUCS5jBYdIk9d0n2aRPUX/R4w3
H9jqIFfb4nHURIt4UNjKSkQ0zmbluAuntfzaZCn+LncS8djTI33OPqpaoPoLSsrK
cR7B3iVCUlW5s4aWhkr6/abmgZZLxpXNSi/rL6UNmZZW6lkLJR2+Ub5HCPofZWbJ
kYCkOFVCUIAcDYNvYAXCu/K3y4G+IippKEaki2rgEe188S3saZDC0mscnhndiBAD
bUUJhF0XDcJGjgJ0v6/vPp7ctiNjQJV4WSRy8mQTW/3MYRiggnEMkE3iMGL8j0Kd
NGi45S4WtcLpJye7EGxyIDpGKwKdLCgoz25KF2KozUp7NOxTy3S8boFIig3A7dB/
uzudJDufrq0E4BWwiLRtTFwX0rE9GqVeK9WljOEdDb3tjhIq4BE30VI6x0l+fg+d
Wdoo0T05duR6S8HaoQ7xCrpXFiqpapQODyk+q0i8LB1AVmB/VOFoHKZtVRIrNUxT
StNFvd2Fu6ZXOJmY+e7Q/gjzkSFLA8dEKvsRL8b3H7ECTlEZibts6rckCNK0KAh8
LKNFHXlm3pap6GFl/HC5LtcfE2+m+SxTHcVuXWVKt5DCzLpT8yKL93seI1pJrrRZ
plsvPQrmf34YYSq42ugsywh/Wjn6qGUXhSqM7TIAR15dMXHsTlbTCFMEgHxiZUhT
3VcsiL66ToocQnpce7ErlNl2dS1PQEPAt/x8z2f69fyJF+TcBMD0SNEWCQKcPewn
hll8B1MLMC/7KnV927F2vCq9j31Rk0y/55lkUwBG/SeZ3RjJDxGlnNzfNrWqa1jY
SmpwSE4w1ftTGyIU2qAdc94t7+NjjWMmggPeP5n4V6nCtd+Me26+xP/d2xFayZJL
WSHokiru/+LUR49w/ngQ/NmWl2GeTigaIFwwbqPTk/J7PDHAhnJ485orx5KJq4tL
HOnYUZkYk0W79Go8wVuEJh0pVOb90kpnF3sxIfS3dX47InstrrlDcdxeAPQsL2dl
tIimGZp9pt97sNHR++JFyqiQRg2uxx9tEAeoI5cmHtYXCiZa6ioQw7S2P6b3ZKjI
UMVm5q26uRQU3MhD8CM6RFC5dkAN5F2itbu+elmw07eP0txzXC0FRypXQl90uDuu
mN3+oZLb+kYs4b1dPru9HCJdznRaQhVUj7e7mqPLxvAcOfD/gR5Fk7sH3LJAT1ZL
KK0SmJU8KW0zWZYA/28HmUBiLbWy1tda2AL+xsNC4gfRkfOTJGf6j3DUCppN+XWa
Eo/mP/TuaASxfd8RTHzXdIvM+TdYrbNJgqET9pjEEAAis9JAC9BkDqa8Nj3vB4qu
1ro8ZcQPVM2qV4NCKUO4kxHfmx4EH2/mDlUV2ltuVK0w9jSnPWBhexuEOs+VzGnr
VDa99Hl6hVTnMHYECK9ijb63WC6r184CRYn585nX6ANaGc2lethwiDEfsOMqDOiL
oqUDhzC12ucjG06X5d483JYOaTHErGi79KIQrhuaiRriLjbUaH1rnz3Ie86lB51Z
bffL3z7Q9wMKog1C8jZfpXOSrG2kGTxsjMA25/DXFgoHkUUlYJm08tgQQ+hK0FuK
YfgQSpMbUoo4C8zsQwCU6PloW1+EyAoXJ3D+KnNPsLDWNr34weF6j+RbZ3GcTQNA
DD/Ji8A5BB4hv8WKX3XWMoDUcrb/S8z8QcC7FSL1kZcoAiZzH+zRRaxY1BHA++0F
W/rgKd7aXFvMWa7Ymshkm1i961q4iB1oZWGSuZj2yIfIJtyQgiTSseXmN4WLkR6n
K68PN01HK32xgPnynfwuRJwGrK4/inAGnE88WnvX514eCF3hG3A+zlec/4ZFT8uS
BSGsXvI+zIG6SIVf+axTDTuBmsta7dvxsC5m7Nzei/ZRgp9C0q+3Lu6rJPfqfFjE
T2N8TzUTQHhzLexnZowTQ7ojexkRxr5w/30PKCVMBksHUSxPM0pbd+ccWmg/QSwR
KBcgpDrVdgaN2UMT2zJKOhSim6hvLbKGQvnSI3nv6rkJR+WDf4jOX9dBPs2t26k2
erfNThzJKVT/hig39egtKF+3wlta5F/s1cVG5oSrNO/kAFrDt0AuPE1Bu0TNWsRr
ECG6RPlOTT34UoBbCBt+gdlcT5553Dsmff5Av9nksuCYLh0TZ9ryekmMtatWmPET
NEsURtVLVib6y+5MuIAA0N0ojL/lncDlQ/LYlRo0Civk2KTeXSnOzgQUKhDstonI
nvWDd/jbGU5NOGwpSgkcwixGabdq/sz2KxTYGYKAKKerIL/dYWg1xOjov663Pn/n
ff13QLMvB2SQwPha23ogpdTVUei5HoowSbeMNVRRWOTm7lCHPXRVBCou6HGih8BQ
aZH2urkVhQbxoEq69NZ+lgPJvjL5cOUsQ17IWmVNyKQAnH1vVokbVAVVhPctbMJo
BXulYNtCIae0iGK5kRjchg7sU1vMzF7k2XjFhmmKMOytFCZGgtESv3BT0ju5pApR
we2Tvtyc2Drathtks8ovCv6CNsyfa2PWN4vPkY4ollxd5OtK1PopxEnJKVdib9o3
s9kfPH2GHpKXkox4oN1S5c+1yb2NqMNX82ZQEspwOBP+MiIUf+1Gm8yrnppjFCSo
FLnvrjdpquLKeYgtFfDXYwvZY+y9lcyLBGqe7AJj03arqBWV1fwzsQg0PkaODJhh
Uin1Sb48NRSdSNq/NvoeEC4hNc+dymfbIuLjWmjLcOFHZprAK63cohVzH6kRVKvz
NglO8uZIMCtj34TIwmyTocoUwaOYjpKCKmxYQeTRE1fe4F7sHAxtcgqTabUMf5I/
ZvrDveVb0GEUfUCylnMI9wuyoWRQ1PS9EgL5pIzGAZ9QN2bJKCLSHcUjGY6F46ak
C20zktZapEtpGmtPw6K6Us1Xyr2N+h9wFRbgxtnlzqzqHPMt8XtYgEGfHGjQk93j
Y564M2gE88/u+PYkOpGuWCjNRm3rFG+Z36DlOFLCMq1tymEVau6wj3Ayi+ZAKzXE
HWzN1BVBcNDNX6WeWtSJY1l8zBilgZkTbRI8m6sfgNfdfc1sNGvk4Juviz+nm1oT
hrpcN4M2V1hZAjLcNloJPlJhsYtBPdlLWQGy+/JnWrWihogeoo7+oco1wfOn7wPP
8cTudNEkfLIm9EZkz7nGJvjqIP+2nx8Z8BAReMKC7P88EDljxLXGaY3U4+JzniKS
gweP05+X2pfzUHXweEYmHUeJoOpd5XlDbqsNt7L7gagTYeu1QGt/pDrPCfU5muq2
wHwMvROQ5+rhoZeJk82qK1hH717erPnbZHGxn28D+icjym6imq94MGUr6FE/Yl5f
9Z3qBm1cB9xNhsKUGoTBRTXIyIaHT82HxLz1FpzURScHgrRUtRb/jxndl/5P/IbK
mgD0o7qg0R+JLI0Ve5fZJyQ6vNhKi/EPQeZlqn8yp4t1QrOWUIQ0BPFDVHkNVObZ
p0XZI3TuYJn5+4M02O7LGBjHDpFSLQtmCdD8X9kgbi9qcMpQvWt3Nr1OEWFmrxLx
tPQZfMk3DkXhOaiadBlr+YQrLp+4lbou1ZDmstCX5g9GipOKXFe82vy6PTlh0Pib
vaZ/tZ8dNQtqpxAnEfq/I4Qdl3wtsZV5YE67X/w7pIOYnPi+zm0vlqNdec8Y3R6e
582EXjAhmGsx3pYdPShFeRj/x1mDuPU0fCqZJpYSDswayhqpyUJNDcbh6gQPqxJa
1geX92JGDjr5Nr8k/4Eeu3JOOMYaV079FhVBNZVvvSNmQR4F58OzcTtnK5OlrdBy
eCZQGbpmi45AD7LWeuEzdggtJQLFS23SEtpRjwn6IiWJi1QPIsFCTaPrt18sUJSU
MBt4LEe5Vn3ZmLpKx98M/mtDS5i+OShS0w1WB99bQZwoeqfAW4qFFeGiFzmwtFkm
nm1bBYrPA4EnHjRL3iqE8IAlWxIC1RBxVYDsXEvlvm9ni8HQGiYGg77ERL61+JkI
iaX5NoI1f7cyITgXDJXiZxDg6Hkgz3esbZNf1N4rbr0YfXC8+iNv8d/VSCwn/Bq7
afp2o9OFLEuZP4VFUFQ+UMwgD/y8Pj/fodN0r4H3ultAUxEJPdS2p1pmNY8HgFWF
I9pyPk1g7UC3e+6FJOOZUbA6+w7VLzaQgbaQaBFG4hZWLZFymPDGGJd373QDzToV
tCxKfngOC3zjACHKJs8rpftqPipQd9gT6nc7+/KyRshErpYaixT4kL42kQGpy0+A
NMBJ8kboYZh6oFYGjnK7DPwLAAE+Eldb4eAxmnJihEU/bBM7ElKXvaaph1bq7Yb9
tq9+BfzerDZ6Ul8X9kxPbkO/0b7Nmg5lbqxRfoPZdCN6VZL+RehQaYbEm9chXRHV
8JlTd+XFClGmjCt7OeAiebj+FvTEFJke8wPSxtVshe6rDeEsGSk7KtYDJdfelOUA
j4rv+HCtUiYzVf8gfCEwHR8x89aue7Vz6eJriP7A6WumpGezV4rxdRvvcWUMaUxI
4tphYTX/YaYurVO6PqDVrpKvk41JMrwpi0uohCc8DiFZdMae7QV9x4qHUOcgm6sF
B72mOnn4lW8t9ZQLSHouorqeJSPEqu2gBhCKZn9WUEY7p1yuNLB5/kFt1Z4cFw6U
KuoEG7uypgQiixuQuR2YGNVKuVtl8kYU8EtCbA+Ki84ipl3GWqnwE6ft22zC8mKZ
27c1rKuBDjCdsV+Ax7ixSb0dShpXMjEX30n3vgUSqRfLYJ44jQN4LN2VW9aU5lQt
Q07D/m7OWy9M6KH/ZYJw0mkNUufC5e92+KdqnR4WK4IzCFlrENS5Gs/dAZNuxD13
QlKKmtBLNQqSqwieU6/G/JnbXF6zrJbDFcI/K0/lY5GHvvOMb3bp0xKA31ojonaK
fNQzFktngGaUPa3VmbJV/insKh1TnW2H7rf18CI2d1mCjpu3Q1Tu3kBjZUPggZwZ
sKXsfoJoBSIMWXjoHyDLfBxyvBX2IFVxCWcd3k/hCJRHCJAr6XrYl41xox9BgM3L
TRP5Y58oYbs/GLgUE5tjt+U6fGG/Y3PV6R9EsQ81b9FuJjwhcFAbrBCKwUVb/mBT
3b1Fik0yohTro5oIQwbXS8hyg9r1F58zU5/xcJcA76dj4Ey1P8ZO6H0sBVM78+GD
3BLnDq+R667xs3mCbjlqEsaTBrcGvTFFW4VOUkhosOgtfbWvpGIEEKUYzY+LIDGa
Iko63IWdpmeRaUVxJ2SlTYYXZkND6c145jAQd5AyRdvKERZpimez3mbGDIx7BNGs
P6Dbw5eaJ1DO8nhAVcQGZ4iJaSgHeyTDOdgztoW/HMQeU/bQJ0o1DRcodJSZ27jp
rzmVD3FHF1Bcz5daUDADCEN97xqZFG1HwSjalftZCn+Yw+lbyYLzAfiT/YfwhejY
Ja/x1nHzfX7QaBPHzqVmuK1iqiW5Z8bq/irQgDCCy4qDzjv//RAjORh0mKO5YLPX
2DISyHBaFgOobgSjDsfegFSruWfjenrv5LQBggcM9iOGe6PSszsjaVemtFSx+AxJ
32XexAGsslUNPdKJWeAXDUbEVRIitIZihRK/r9rnBtlkouv5v0U16+GADvIeex4f
4uK5elI70rPXtojI6ufkvg8KComrxv3SQOozTXt8J9OvA+wQUti/PD1oVgQt+6j6
WCsPlncZVTQCb37OZKpUpHifit15cThMfcymWeZAjPIHLWbuXDrsj/n8iZJWQAXH
jK5awuf0k96TTYAecUW3ooN6aMxPgJ0YB6QSRMnoqYltF/LKb7vrIYz4xHfk0e1B
SMZ1izF/A0BLO2skGLwrwqax1RLE8uXHFjjSJaQTGrg/a6OEoRm9DXTIgHhbWOYd
3ceoKtQfNkxQlwkP9Rz1V6s8JeMuNZiRZRWUvzH1sZaWkZfQVakoY9hKTUyBJPMP
fKV4xprQunm9WMyllL0+iJts9LwI0bXy33qFI+m7hYYQeLy9NVEzYnCAuJeXl/7x
+oaVpfYXtB432u+QezkSED2eRzWxx7dLwlwy5ndu9lxLqsvpo+15ATYZdU7tJaZc
PY+VM6TgmpWwkPCLKbHrXSmTgFi9OZfP9j2NziChKy1C5k+KauJgklcNYAABnkh4
NDiNM6MlX+F7vem4SbWyln7qZstYgWkZipDNz+Sw7l+xC2l7SLZt9f/AHKYECMcv
MV0oDg9czSH6vJynH0pW0VSY38XaaiCcTtftOrkSpLpk//uRUu4YzQKu1M32nqFg
MjbtjNWxI+naplAQKPL5rT/I6JJ8kOnsusIQdRaEQZniyyeeRKsGpRTJ3P0i38ez
NA1m+28kNCPbwh0PeMi330UNwsHC6B2S3yYLeBO+F4A/lFIT2N30x2ZKCw+8SvsW
jRADWgc51fLtknX3sqnZRt6FomqXqBnDTfRyhmbVvDhIo6xit0WKeEUtJocBDAC/
40UhY/tSJCpu5cN+c7zwC5TsoqygsoogYU2Du50Eu02H8rddWh1A4/Si+klPhYT4
EKNgPX61i77eOXyoas+wyqWYV8NZNEnkim8g5y9O1aHMZFluwwc84EB8dZ1C0HmK
SznMI03SXMtwzOcCu5QnjCyN7UiTG7YaR8v43OqsWwrlGWNis4LfyWvNrCsNa+1D
FQ/Y5TXm3Dqye+IdPEA+m+uV1KaRfhrxQ2IlXXuQALcokUdg+fmj289OhpBEG5s1
KNW6VriX6UCDtrKy4k+K/OtKFeYBxbI3XB8ty3KPBBJeJ/RP8l488dF7hoqf/hUA
rT76DpfBF2b8jGb+c/4dleD3dCVrOcNawNOLebFX49EgqNWSdnzUl7mnQ0kqrEET
vE/PM2B1lqxUpMQ0MAePyNs0HMRQ55N10Wq5/QvpXYJwgxj+3/OZ36cU97i4qfbw
UMKUJwLHdzn5DE7805COZ7NKdXTdUYf2mARd5RBejwAivPY5gnDDuYyukRgWJwXn
Cngm0Q2gyU51OjRcjbO2cJCw/0Uf39V+k7ZaSYAEyF+nc9LOdmVGDzMcoQafzA/f
PgZhN2utQc8TS+9ek3zt1tOpHKPuEMg0nB+OEAOn5U8dkYM5dC2gsdRvJlOQkMXM
kBl92Micdp1lXH3D56w+WDbxUR8/snAyJQ78bj/IxEXmNEGo1gYRtx0re+d/s37q
dUnYXCsDeqXEp1MjMo6/u2waAPpRF63ZsgZfviLgFN+wuw9jcEk6Mp3aRwj/otXD
DiPv4qQZmOCp7quAyG/13N6HMXpvDXLbQ/XBzuY3SGc+FGw3DwIGIOfPK/+TJyQY
qRTkQtXz3JIl19AQeMpBSiuDloTqCvNQrbz/Rj5AbYgiL5L8WSB9xQ6+E1EpcRRJ
4rfXDp/JQgujCmRo/66/DIW0gSmPeBCM8CHTIiMo8oYcy5koU+74l5kX1Z8Cj3rf
JcyjNudNRot0m+Aas6pGlQz08AGT7IrqWJ29kuN4i+AgP5vdnXSGdF9xsNZ8hxSo
fov4K53hh0cg3/3phQuW3C3HOHCcmn+qqeXjZDxOo5YcWAWHoypAGt2D4otwBRUA
64Vdu3FuMsXRDgVc5TFtg7z+B16pPafY2OFimgQ1sQyHMPGdvuS7Xg4nI/AQlUNS
1DmxvkSY8zDaEWDI/LmLTeufTzYTUPE+vRfjZDfIwC597GzDxy3uJmATD44GTuMB
exdZz7uqfM95qzj5XABbFktpJPlTeYt/pyMkL2jmtclg0m6szhKaQ9IhjSuMXmzI
PKFPNwes6m1eK3Yw1N18UVTvaQL3PghFYuZ5L0PacuNsMWoQPutaljJ2IePcVyLB
fd1TeiVD+jiWvUktOg2sBrbWqv+jZxO1TkWeH4ts7vEHIXg/7KzcnerujqrskHBL
jqWVZX1xon+UC+QGa0i7gXIFSSwkrXx3iyflalsCoYAhvBi1vF580WkunLwxk1QJ
ho8+88XmhCNJtbR4H4vRIiqMt50cOhTwyPO5Xx1CSwhFLGJFGbsf394SnjTW3CGU
z24/Pn4xvOb2oV1EgOZv9orsJC4MvAdVqB7gYkiLRJ4X1gFkhek2G616FJBZC3mw
O1D/KxGfPHKQ/ed/Xn9h/XINnMjk/1yCyGOYBbyH1woza6AQXz5ItD4lYo83AXKE
MjlqENZ7Dk1AGMxplU58B5x8ddZabtHO8zPmvFbMMFBqhe9JG1DLQfDmYRfmCTH2
W3vRWjzv9k70ZaRJg755QxcQuapHhMDpOJLTFiCldGxNrF/pb21U2KyqAidqbo3t
T4D8+79UxcoOPyPCkPfJSDlh5SWsgf/QGvrQ/vwti8RnX4zeJy7UkaYQn5WnNkmH
MtMeZANTLYdCWV9t9P4zMHS2IkJzE1S/JDUgDF2EYY+78AqHMPKvTBqtRnFSxe2f
y2TZKbUCYmdIY+OMDNWpqqqt0IOo/luMLo+ByAVASyfJ9uxHTee2DUfauESQr7gN
ufKa3h595q8peFGBZ/s5iAD//K7afJr4EWQIxu7apMmoNA4NtX2FTTbzyX2RsOq8
nUguEBZ9MqWBRpZx62OulbgJV1/kD9p/Hg7XKlnm5riwUJhhUOTE15moIjgbNDON
LGS3HUpMo0S4h2gL8uOmF2DtHhdPvuuKQt5zvDzFZSv4O3CL68IaAnWINIc9+GXR
1Mt1gZjRwlXY4lXKRwNnZXSBfsPiUmuX6XAq+Jr1sxT4TOFy1yq/xOrwvsS36Vv0
RFSFgNrAELi31ZzgxJgMg2cEOSWKe8t6pUUwgZ5GmdnMYU+ikmAvWw2KfCsstSIK
J9zNvqFF4k0mCyl3zVMhXmQ9q+P87fpx3yD9b2Q/xbWU2NWQ4SiqE03S628fHYJx
7JB2NiV683d/7DFATxPdKyLs/vNL76PgB+b+wgI77ReL7sC9jmbdU0Ond4tcni8h
T9Bi1gDQS5EI9TC/VDBGLur/mYp/YL/klvjgJfY49fZhflqeMbw1obNR5VJmCBML
LITUnir1OUAlmiuvcCJsN25h7ClvVMML7Icc1A/+fIZYvWfM7nZFhUo+UgDCpA06
Y240SR0Ql+Inc2rk7sEEEZh80YgOqBN2sztyOjWTLXJVZI7GetXzrziMVWYhYlUs
IeYtezXurlWa5inHjyMgOdWx1A2UnGg/EngkkgM/LDSnZQ34F8uRvc9cvv1Gk4kn
hdYMEMd3l0PvNYiJPHw+NLl/Fclq/YkMsjcabSnvxVb4bYld1Ir3TZPVA3ltG8+M
8fqwZvMFIh5FoMKH3DrtayUcOqAzTVlKM43X/3AvORZ3wL8MmTb3gGHn4ZqZ43Ct
QEINgdUWQ0Hwgm4Sv7JaeFNmJb52KBIu3IOIVSlky/8o2G3j9hjmz/ET/gR+bgOo
E7UjDwgTmPp7eycblq9Vlse8F7F5UbZ3DXahs4UrVTfBSnrszu+sFnjkaFYs3DYH
uvR+ApW3998qirPxvnYXtA/1dhpM17dBtZq59QhOhFgwO5I1kYTERCOx8lYf8xiF
LpZeWyGlPZPBWUw2XqE45RkC9mtq1hpn4jtx43pG/Xzr34Uj9ClMsSFePhttYXDG
94VblFcxsXwAiBWzxk+boGrb7QspJCQiyMxkGvaV9zfxG7nlWGCxZnmzl7FYpcin
r0nu4t5H1iWt+DG8/1R/4g2obI9ARLHEL0YR5OXTKLGN2OuK0wNikYUUmQVyt3kX
eQHnopKXZgkCqiDVT1olf07dZO3JbM8WlvH2rsur34PwARx3YSKTBBJQBy+jG2mJ
366qY1mm6wZxOQ9ltRXaBT0F+tisfEe1A/NTb5fFfERLOgsuNCbzNGif6lUY0WUK
4aaCAmtIcnFcby7JoHDrNuR3HwpyyBZF9VwXD1f+lKUidGDif6Eyj0y2AHfOzlNm
JZlHFia/x7O2ZRUYf43QixRwdWCDP16bFqVuSa41tx5S2zIQoBlRXsFsXBATer0S
bpqbMSSK5ctTYGyC+KatGzvRvm1fGBfYqo+PkcmNNIrPMaZHgfEbuiqIQH6gJxSw
LIk2FU+3MkX+rF9x2j0DOLkp3rqQc6r/UphTykCw+oyHVnBvDmVHG7YZKJZKuUoV
ikg9+0KvYkJCTm0UOxJo+yzJdpHAWP3VqFcGHDB4CdzSlORhmdgV87qEU9VVOMIn
QYoHIqm3isyKG22x6eIGDkw7x3WIfRSEDbu3rLJKgPuHn26tq0Lezk3HGjKq+/CP
gcRZce39PWB5+sW0TKJoJWFBgVillCARySCPCbCzEvbRLA6WYgukY8ZK2q0eJjlJ
JyUGrZ+MX/7Kc17WjmfpuUD2XXC8mRrebqIag28I9xFzNH0VC6DA99rNMd+/8Y85
o4DURQTlxwh2SSHMQ0DLszdN0lp0FoJsQml7p4OzofRBLkSewIyf0IGr49IcU2eE
tJMw/ZqPttOon4ZSeUiRYiL3lE90pSDBUgmatFi2UCBt5jXW6OswcqadwScdHgJR
q7S6I1j4uKagCq7FytdnTRJV/CEnUfKhYBIk9mdNMBO+I84cCw25ZTV7NTOJH35F
vNlyDszYC2rbuYJTZipouw0hmWwtb1r33n5XoqEKMNNFLhMAWX5y1qCvJoGd6D+7
mI+VrzNnjCwddvhbRq9ZtGJI0iyi9Dtliuk10ztOs+rC3VQIW7wgsbGTYnWRRW2W
9VD8Qog2bTdsiJz/ya1NfABjyH95FdmpF1fmGGeB1cbPSyndBHhVVIRL85PyDNb+
0f2qDfLut6Veg98wHeec/ZINgt1C5P4YlNECsUcrKx8Xr7/zygIoI0sJ0INRoZom
QraJ/BJR5BcAwlBchiarMBITej+XKPMfefLXwRrb0zAfHHd+umWMvoYTjM+4/MTL
tTCLn4RpbRbivthJHwlisZOOhzqplfMVNIRhkk0HTwW5tzEgnOPbkYV1K/5SAFVM
2/nmFeVSw0wAwPXmlfmps8yfvCeUni8ENMaBitSVjgRE1qWMq7bxXSQPWOaHQVj1
j1Th4iPmb+lYhyGRLTeSeE0wbx/OWvjXs+MdQvRhOwBDcn0RoX98apmL8kMUs6V4
OhtZnkPoU4O1fRYOH//flAXOG4Ok4pT/NOkIqX3GnSGGXRnx6v3EBWqlhAkEdKyx
U9e+9PFUb6tG+nQiNxYhQzG6a7e3/PsdhOZ3D7nNdfSfxEwreUknT7hXR96hjojI
xqPUrBmEknrpvUQcFdYxT07YqKh8tUVgvLJr2FfcxeExIs+18ntp7zzqgDWWL0aZ
Qye9rX5OxyaAceO4VLpjlsk0PctBZwhki6lh2T3l2QgORZmyDauVpAGsembesPlI
gOwrXWH9hcjGG/duck43KhcC4NG/Gbt+zqXHQkv/S/sBFm14HpzUqQSvWvC5cPzJ
90oBjol773t4TuDHRh6z2PEu7LBU9d488x5jVQd9jkh2j2dh1ELF+UC2qEpoPYUN
kIVg+i/5+Wno6kkB0OLT4zme5QAocveFzHHu61yGcrTAekDKWtFwQLySVM6O5dAj
riJglhb4KruV/VtTggAlM/Wtg9LRFq6GZgD2mfOMSuxrEI0A9IIlcu7UwVInhpCM
xUpXVmo+kNPzvCYCk1MprnfdDmXplgPJH3VXWq2qBl8vRyyhpYleIRg3CNxidwzS
fsJfyshn87sIDejtGU1gm+5TFBuLGN33kXyKx/RQwQyMARyXqnLFHRfc/kDV+LVs
vnX8UJB1RAyZ3m4KAaxxfTwj9dhAJV18jFc+SzkU273u/zUgzaawQuQin3IyVqt0
JIwvDkVyqM+M8XmqNYDOjcEj5TqVfmKEIrxRZrWa/bgYQvrGnJyFBywdkpogAcdg
2636E0lAfkHq466og4ehRM7NyU7qWOxMD3ea8fohGjUQUWc9V+yM5gGnVx5TwLQx
fSqrjoHV3mBgA3h43KiN2YdB8iQpIXjWPY393a7TCqTnJJibaB2lCDjp3v39kcIS
teOVAQMgO3y2D4cnszQ7Z3NdxUCMsmzNI0zsBIxTf+VdlZ4WUA+tcoLHIsN1XE/S
bMi9dgUXhmi5UqC0BOVq0On0FIDyG/VAlkJX+53oBe7YEPTAfLum++osZDIBHH49
8noCS/4KxjO35+P5udqkvNZ8eROMpFNRodm7g8T5HOyjR8XAekHyj6RztsOzG2va
7A4CxsdSuA1fgFNy86Am50g8ZwFprAVftXDGin+hKrrGg/qB3Vz7CbeUGN6omPHc
eQXU9n1yPb3sF4PQ/vkAKA+c26Fab+GlqN0hZvPMez3yDiGMI/AYVyLzQaXegGFq
mT1tB7QCGmyQXoE71fV6vcHhIXD6icPgit0iiMhgp8k4xlJkwDazciPWWyfnwHR1
FQFCS0low0BeapPDZycxRMjh1w9sTNnZJLCkj7jLXO/0E2rYZkDDBBnf2njBDLUU
otKc+ZfaYpOp/C1TJXpbb3rEHEHILUlwGjK47bntEo7ULueSjFjJvXrzrccnNK9F
x9HmhwJ3WA3xqjrc4hKNCRo6yKMUS7Yg3d6MFUQOfTfa8aBMkdxu1K/5A6RagLzU
Sl4gKTg7uFTztdp6g4l7XCWAwHJDpdempW8RV6LL+S793mnF4uytIZnCy5N4RsbO
iG69uXf0ojXNY6u+RjZNGFjGfKsRiiFr+ji0TB9LXuvPOzA9ufF0mB14oGkRXumL
WlMq7sViiZgkC1ZdDSC9o7U80DgplEffojX9ZgE/QGCtOf/mdqMp7Wqt7hvalLh5
Z7ZG7RkbS2mmB/QB9BK6FFxYjjgFAdXq/YzNWsuc+iZTO8jMxBSYk1yU2qSC3C7v
zOnhUfxPv6Upkn5X7p75aTQHjdsEmS+jXbI5BOK4dP6zirOWl6lCY8/2XPYblVHi
YHDrj0tuB5k/9Of2MmO+N+n6J6SiIz+N6nBCbzd01d5qvAobhxPKe8my4eQLwZwU
VhIFYYrKB4phM1xc2xMUGe1elBFykKyeB/M+rvuCEdg=
`protect END_PROTECTED
