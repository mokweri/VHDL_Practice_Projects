`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xCPy8WkMQY9NFq6xKADMAsxTHN+bGQeBBLNNPgnZdJw7JEEGcsXfgJk0/SGsMKc
K0X5uvTCe7LGl1j6F/rWI0cSviL0ka/4EsbO2vwvrp79yUJMMLJv0r6uRr3PhJH1
JGP7cgOqT2njP3P10VuJ07vW2B1pVxCDF4rDVIS+r669lUUW/drcvJxAtt1hJmD5
Ebg9cD8sAqfojnjAXYB89wh+QCjGjftnSdmgAy8TWOyO8qPKw4F9gdmhyo1w5RUt
rxemaQEcHIDSFZvdlLb4jSiQOD06tEHqFlCpC9nANl7ObYWfUNqq5/mUlYx4QYl1
cyQeOrraVLPXukbl4EMUH9QTaG5kdVHKl1qcKsouHk69ix2x1FJ9TrY0ZwawhKOb
Nwlj5wj4uQZLtH7fhKh1ZsSo/TS6LBvcjVu5kuK9P59v4kSTxY01kb9WLYbooS7r
Q+9Lzm7NFPViSQoTMgaAVXT6g0RXTpUhVMZ1hNy92vToIO6WOqMIemeSQHQdl0I3
NUUOhoLNQ1RSp6cFq6iNweXiRsMveRtKZ9jggXGhO04yEKLQpS/5Rjkyxz5weF/6
rkTZ8ktY9z5WcaTw4FApPoYxUIXOSVl5Cr8lZL5kyZgDfouj2HjxLZ0TM68nb01s
qU9MIK0gpw7aiq8BBv0w4al345yy195tql0bOCZA3K8qOwRpQ/9BHXMb/dFXCkX6
Pv72r75UJ/v6kdY2RUFBIlSRA1VOG/SDbrxT+hydlzUDUGKDcYJlhpZ+pUV/2PXb
CHsybTHtYdFp850dWpCl/rXSppeb0+a7V1O7dp0VX1ce+Dg+BJ/ysD/JFJ7oLGZw
E743utxiWmAOpi262HZweMifRLhsgEahSzgHe9+FVo1EsSs6uzXuSEQDJyOAt1s1
qw64IVGPi30Rs3Nk3zhah05nDU/cJD0FhJp6sB5UW8XaJYC/X6buA8a2vZXNcEju
c/CsWL8MQWjvbTB6vo6rAoHiePKPo+rPAphBQZNm8fehVJ7IxarYT8Msr522rtmP
JuSdPM7Y8t0fX9Fi8cpiN6WBB7VlclDu0y/llgjZvhL1qv5eW9y0Rvd0Y+i2mr6e
rk4zA7rOTwS7jYaxjWsKf8CBqnLwSc84bltU+e7/ESiBI5ErlP6v4SvanFs4awFN
Qu5exk1E7wQP5Uya9uB4x+N5dF894M4bavZTtgLIiMXOjoR+3RuIHkE0FmxwXoUf
BMPmildnOmsOHsP//vNZsXgdb/dC5UXZnIPu6QTuWN55bNQkEaflk4BDkPjZJiy2
D6C78HooO0SYpTKS4T4rA52cBcm64OD0cNz85OberyahebZ6cFwXQk6aPD7h/nPi
ukWcRV2umzoPhHYbyXD2RK7fZhxecLEAUxb/II8zmxLo5FKmJmjDnX5LGYRcLzd+
IBwmnXE4UKNWWaK5MYyL+ir4znRQL73QG3YPkcHTzXAocdTDL7GC5V1p2hYFI2xb
bpReLqXV4HTvpZsOFfgwjeCoPWy4LTw7NfZMPKZxwAIsHWYD7ZlCJnilssN5alBg
Y5kAbntQ4mBj0152DWy8+8gGYZl7szBdDeo4T1jBL93jc4aNGJUYfXFI+p7oKX66
eULYVkySfad2E2Kh/R1gM2nVuCvG3mrUBDLJjtxUsNxC48Syfnl6txrW+FDCNsfN
`protect END_PROTECTED
