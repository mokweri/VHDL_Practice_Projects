`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2NO1L77JVee36b5vMTI5nyEp/NChKVLJgYnzrWRw5SnZHpJ3W4PeU5Y6O06Pibix
0YNZh/7hrNm21Luj9/vnxGdThMGKMQe0agg48eUuYzWrxNJWrJI4Zfs1qFU64LuR
Us2AJDFXVhL0i3LKbBQq2vGdRvk2cueEcRgdxZNAcmFB8AgzNlkJ+gfz6Glmc12I
rhkSSokqHc0CwsEhkFn0L2Jem1UYmgSZYIHCACvBCss20tPdCbbcm0o2ASSe5buQ
N0FjZuAAQSFpT7q2IZetBsTV7WhxUgtXW8aySaU988+zk858mBght8wBDV5hh6AJ
9Q4RcclgaJh3K1Quzy/hXmY0Ykc2/e9vDvT/FVLdGASe4crcAGnvQx7XmfVWMq4l
GjHLTd+Y8N/fwcLs69ylOsSRli9X1lIuzOmkFYLovQDQNkMFDtuDe95VsESb/l5T
tyXAVj6YgjHtegcKoWaEhW6FV+7Ap4t1t5vdtQAxVJxC4j8Rd7pTlQjd3yjNT/ie
O7A0WTdAuN0q9YVhNpKfvVXXbK8JK9Tag+PhgCpg8gzGSdpSrWrfYOSji9vBJ3R9
/rupBa8R9Sw3i7OFjgXmNslyr9l3N/lSPWql+YpHeT4snYpXWU027UEbn2mPn4JS
ig28OUMwoy+bb27O8RaIHoXa5FOpeB60r63a7GGalcsvZDmr5EFp67Uw9WVTKUZK
ibkQyCYcg/Lfw6HDimiG51QzntKbyYpSvEIx/mR/0xiYDBaJG0mif7M5xo0Jk5cm
bJ2WGys09sTkOdB2REwTtayZtp1AzLpZQ/gK7hEDAtCUD4E5h7x2gxWESnsse7U+
w4YrcPIcJEdXe2IlnDIyOuYvoYNchQhJ3fbvII9BCSDDF+qsjAq0nus47mgxomTW
Yhi52Op1m9jqrXFfwkabMwn4KaycF1stHavm7D+5NsaiMiTZfno8AAnmezKHoVCn
zS6/7SsmeF7azUXwi0gSfDAcqN1k3eXqZM4ppwnshuYlJZvtlHCMq9olKV++ryR0
jHOjyB1dNWoawsIWKG+jLaCNpGwiECVIQNMjDfaKH+XCP388/sbHMFw3TiRdTIRX
VXQ6RrbsXW5QrEB70CNc7unsuY090X9I4spsjGlnc0U6hlxVKfuL8SyubleWsCG9
5aTOxC49NgHYoYvlIk2nAq2mg+iQJ2RK4X7Sjwr6Ag14Qj9ApATC6xLAHcZp7mGT
FF12lESvMSzNqwLkdt33fHnjRKkRz/uju+lBbmVB6Y6tfOc/zDB9ZjkEiRiOLDQg
XQu7gn//2PVnih3KFyg7CpO+nBnX06cSR8L8STikzeUc3gVXVbRnT3ePxZ9lOkCX
WTX/Lf4vVgjZMptvgPCpxxbN/t5V/bVYkiPu+OvWH7dyD6mXf4ploJxXezWtW1Af
nXt8mR2IVSdUsOfX7RZPXCrHqdylF3DoOumEKQvzNaUhP9XZedyFjaDj6VY2vCsC
5Q6I0cdayx6GlG4xeIdSETjB9mjEkui2CRXNs4PAX5IR1Vm4l7gYOS3EfniGXzVv
VfWfDA1jXVoyvCsoNHVw1I+lEYp6HfKo9zVNWcnA1jMVCYT8gUjk5BVD0Xg82934
tXdJNVLQR3QtW3mgLZ9Z6nq1OoC6tBP1aP1ethCash1rLBoCcaEmGNKrYkuEpz1a
GuxlCQYclhbzCZsAnvaABMarbs2UJgvZRFsPQyu2freg5fvgqGzzVmStHwEGpU3j
BlYu4/60+YFfzyFlNBIZ4KmU9TIYcIRPRas9iD0HSRW33SvAUCjSd5Tuzzc2GN2T
hhU1cbMImm1XoW8YqZKPx3ROmBz6fXBccUcQeHemqB17gZfjK8luuVAzHamAQ5dl
+jFDKEqIdSD7mR/h7RT9xr+Kci9ADnUYESEeZNbKn9dHYoe/XvnAA8ypquayKxLr
G196QTQIEwfwrbcc0gVz4d48vYkRTymT6nXQgdhS78Z1Py6sWN8nDr1Ool4kSeVR
OHFjxykANJfMvgeTgM/T078vmitRdiqGSAcbQQDYcCzINYJn2n0eVAc6x5YZdbjS
KRis82DZe4cUn22ixaDjT4Or2JsJdoauWAT6ZbQxN4Q2gHjYRJc6gB4BFqXPGPU6
A3zIVF11tRdP+kRub2z9I6V2CWK3ZK8ogYxNZndll9OKWC13lqFoYsxyG9kMy302
+mKWvouF/icKp7SUi3od3KHtY4IvniPTg6rQWZmOYo1rZsuisdVjDzCz6axAdWzP
tFhv/eVm5862sF0UDUSDRqddLnci+ButP8Wl/8k65zDLhhZa07/B7M0ZmbPITysA
dh0y8r+RnisYrkJhnxTG1+Xk1dY0I6ADmGL7rDnoaHZP0tNyuyta5LviMPnhpLJv
VjUAP2i02FFYKbKDtkJbYfs8N/LqyW79wpvjKNY0DIK6WnKdvvdwXTCvt1uQBRD6
czUFebnUjyJQJOp48T9IsGuJyiM0HyA8HQ8AwYUj4kuGFhfJqvZJaNYLiaNJ0Uky
s5U87pVgl8jM4xkymEFiDl2vDpzmqB9PGoi1+vXNJvbn/SUvpJeJ47AgUtMXN6eK
GkpGP/A73kFKFQ+y3dUAbzH9uMgb6kUDXWlRioqmNxSx5APnICeCN54zwiLsNl+s
SFYUmW/bT8XnXWLsHEsIhlYPtLYKQxilqVpEmOsUTT0B2b1Af0BnhbzHvNZ9wTF2
p6wqjWfqf14a5fnJ9DPB2C0lxunC/2QFALI8vn82QQW8mTR+yCGy+obTAOC53x15
v9N5m3lJrn4AAkcDraaiEi1SwXKJ/RwzvC+a+Nbf9p0mS0kT0r0czQlnDNCXzWnm
WOBdGDEO2XEaTmTrZ9b5PjB2gY1oBkfVCwTMPTpAJ66kYr8NQ7msF4JKs5RlmI+i
7XGOWBNjcY1b+Ak9Fy/15dOx+yCGDPwhKAHvuMdnPqQB20Zfdtir3bbwfHFC/nkN
L3v130gf+8s0LNAsP8LCqSJK0MmccB99owkdQymsUV8VIQDXyAMwMG5D6pRDtd3T
pOYRpf5KMZBVgdRWPVRyUL1z5Ve9LNdU2DGncDthYCL66UifqGgnP4pxL6OXsbpA
Ftu63hP2yHxBcHAz8ifB/0esvXYZ+GewfS0x3+BaMruQMLBpxRzqprbBpj4FQhpI
Pi/FUzNd8EAJEMktlLrWI9xnrf+k6wkhsdq1Tc2czNYowxGLSozXdA4C5LSrqavi
nekg6tzRnS1Ge0+Fp6hbSqY72a4RdAi85HMkwapOdHHWeZ/iFrlnRIPum2j8l30s
I8ajtMFBmvd9LBCSH3dc3fxlMaUKNorcck+UXjAiR7EiiJHGJu7ylEZGXQi/Qnv6
S2F4NRFzICaDdrIQx1Q4U9PEfh1gwTGcsDZrDEB5FOQhLZiFkqy8d4NEE6j2plVx
TDd7Mhr6X+tRlOp+yMwxal9JdK+vVzeVMI5R4DaDoMc5/gYtyGHLYFJXvi4OHII0
Qbu6RAMxs6wFNv0ks0OMyb2/B17iclUxEZDmy+2EXmU/yj9Ng+a16L7lsYltuxyx
LKSQDc0CVg+E/BWUZd+xcrgJ8Bsh5dIfunclddv1quStnpwb2HWW0YsfwqAEZrW5
szMrPRD4KeD4eAZ2aRp7hkbgD3QHvZGugVt6rR4U+6JJBwyGY0shvjo72Z1gK0us
azkxbJbvTQIeZev0B0jnuQlxBTWStLuAJCptCfRYQyyMUwPMyHeJ9NVo3ao88xjC
vglBgovuB1gv+tM3Iqa8OBObJHfOKudskYifIraxOpavthv2SWJFF6TGurH9ApcM
0SBB+jNSpUh9yO/7QV/tffBT44xKLGbPk8QxxqP/RRXbXIlpaMHzmfP9hAZLGr4I
MTsKDoCINamT61E7+Iz8khHjWR5ENbBFHpBN9CRdxjDNZ08rsgEAE99BESJ+v0CC
85wE1h8ZnaCZBOoKrkVAZ1ZTM1FuiMKpAn61VwVoLWTRlgKiE50yzuDc8Yxsoh+a
gl7xMT/+TVND0/ieHDB5AMS3Xt7YzWQuGMjq9H2KDnFOL05Z9UEBMyVe1vgrwdX+
kvEhgjU/RGjOnkm+DK71kTkZng4ta7tWA5/NwskRnWQ=
`protect END_PROTECTED
