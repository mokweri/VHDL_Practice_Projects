`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CZXQffgDhApu1tqdjVLgPLEhmyPE66wQcVlhzgQNZaCTiD6E7sN6AcXjAAjuXCmQ
8/AwffK7r+lsHPyiegJIU3A8abGyqje60fzGeqRNnfbz/Uyl2I8Od/Tn+CYbUUFf
3WnzLBkiUMNo6ZQUenj/kMOR4Z1uoO0iKyDTVtWsRvUpoI8CqfLYVD8FtnbuAR+x
iiQZAy6uI4srlBCnG7EKkKijq3APcrGXD57gQStUG1OHOVsm9svAFCfJ6WmhPq2d
sjMCcEJzqUzisUZJ9VwfOlyvGyqMOVziGx+qbszwDjQU/ed2AyzclQ2LeGKY3H7N
GsnAXpTqS0kDikMmXnZ/Mg0yL1SS9ucpXBIGvfzQhN0IpxT4PPVJw6n8KUnHtL9x
DkOJxu0Q+vizm0C5f9b+xIMiGtqzZ8ZjMLMrWyB2lq+Q+PiBwk6fT1y/eWbPhLXs
i4RsKocydAVvcbGNc4xy4PaZ3iWrZdnHftobew00WGwAsN/O0SlEtbXrpFdxG0GP
DHFinAH7V/SwLoW0mPIbOYB9AHAX7nRXcnS1hNn0AG/ifd4G14U4AT18kYYPSu7H
nWOqlwE8KW/zDVugMb6//Lq+08r19LuIZsX11cCFou99TF+YAvG7rZzv35dDdYHc
FuID3JVN9bqUvd2wKjXdpyGIlwS/Xl5Q9lvg4pn2JACxK8LLVKTV/6XRdQ6wAseK
qsGuMCyzn4VI+gNsRLR4uMapFMJP4vqlCNHmbQ0Q2c+UAK03qBuoZ2Oh2KY54rsK
cV5/Ycr3lnMUkdl6nu/2LcQmPxqAN5L/BaN+pMp1PAGKyPED09f0sqexrvdl7sHS
8rch9fUCr561AIBSWV2/ve31dePowWvsls9COVFE7/vDTIQqdNaSE2/4/iktV9TE
5NQYqO2H/kWNptSLekius2Gj9QnnHYcc7/qUZJrMBz/bELW/Yl/13h+tViisz+++
CvoWc+lWM09FVeyhFCI/5NIOPCIXGoFkIxEd4MPKwx1qe7n5+4SQ0BxX2jG5SWgg
7TPlhQaofPbACLB638E7DHfjSSu78gLgoat3DhxgDxVfiEFV7crNmGAAQZ6L78dP
fkGx2lkTyn3ngjBx+UtFyobJnsn5jpx3iPJtE2HPnXEwNGTg5T7P8pdPn6Qp/t3T
Tchi83pAI774g5ffWCPYrrC7lGzLN+CwpmLYTRO+IR3p5U1jMLoPsjMns7JT0jWi
SnKRI2w6u1T0SP/db6WrFHZSaBk6aHHdFllCklBv+U2QN9UAyu3oS6xpx2heuBnr
dxjYRWjPXPKlBMH4cnwWZUGmxXXFXf77/lao8oHI1GFuUYTjwL9CpZST8NHMoKbh
dEhyXuCFNLuq1t/O4tuU+kOARiAJEzk8D6ACzsC11L84c9/UvbKz2KqTeHDkl4Ie
xUm8s3LWVBThFlno0LOzd55pMjH1TllKxSCxeGTHyXfR3Kn8E/5okUTpgX6aPwIH
/SSL6jOM9bc9JMUFm22lhB9AIL9EBgRAgbp4w88bfjpUqIcVWWafb19Rtkz7akz6
t3DA9WM7lD+KOs/WkjcO3mHWzZaXi0xqe2fiprsAZIxjED7yelyqEKJrC+KpJCuh
Yn19PHYH7uqOeih/g+cd0ZwHJ4Pt+M8jWtm07SfQ7uO1X6P9pWDH/XOkJ3Fuhc+F
H34DDqCrvdAtjKyCj+NgB7yzicq0TpbWigWOS38SzAZ8er9a717Z6OpJgPirzPoL
iDXyvyvRKeLJXhrvaVKiuygZiOr3depGF63a5MSN2NfKL4aCU8a+bnNEd6CELtXI
qsAkUFeqEOFFaaWCf4yH+Wffom76JkOmdVJq+R9sgjEo5C/vXJ43inuWKFmdgujS
D3pNIpFg2uuFe8FGDBC5rFu6zROGfuUCIbgHom3nkG20LXb3xTJ49tdXud1ZmtH7
Mn6vv2r2Xe5UfJBNGG+5Vl5VdAaxsnDmGmepoljptQNezTrUi7TBeoxJaBN345wP
fUBLgaBAZlVq1DhZ/AbInTmymOnWxkvmfsKHLx61wn/ZxDQQlvreR2PewyIRuSde
YUMLTDFAzz94PkZfEy/2zg5rMgVBxOORXdlkIxbmufJF1VL/DIk4Q/gAa9AtHSIm
YGExUBxHJnAnZCYfJgKEIViVftBiyXUkY6eW5PaTlmuloFFaiRFtruYfOtONqy2C
daoU2gPdG43P5AX6105uP90LVB8fmrA+NzJudxViGYAsMuJm5cjdFuYzy0qkpMny
8c+4UN0C5AFlK0bbFF+PZ7LHQUpSWVNxW2oKxjvYO/yloFtAZwYwLJ/pzSOexAtV
WGUlUsvNyQjYSpoYgCV5xfFe8xALeGE5qpxsbo8Nx81BWka3XILY5S+9khtJz8zD
DTVrfizjY/8qfEPw2ZVdPuykVO8E72HOEQA3PcFZctl83Rg2HGizS2f6m7R5axfZ
AtJZQfmqS4/RCZ1CX7+0SToGx8WbmSW3Lp8HvpClqsZ7/bwzl9+8fp7fhk/zAUne
62NZJB4UNQrcHyf+hqMUByJZwPaOxKNRfsoiW5ctBy3e6HU5354lSSkR2lIXe/KF
SHTk97yFYOGH4qfrebjppgPmXm2ISImogYf8F33ZIhdym4vc0QbZ7/LfalOhrAsY
uamC2AETQLnf5M7p6sEevlWaEwkKw0W8u1W5kGsPOJZub4rL1NVG48n73Turio/X
qp0h8LH4O8DUw14dWSTgpdsdPDuMSU97vQz0/eWXUE6CRUgOyC7XaaP/OsJN3bwG
EECk5cfV1MGvJrlmWa26e0XUNb+x2d+uC46nKHHSpnbQ87SHLvpg334An5KF5HL3
4Cw7VnBnJGBS7aI4dSLHSEvsw4ylT4TFHhJKKq5aDSXymUNjNSHoGItvikm/xIln
7wKKhNqFcSOIXDdD3D3JiA==
`protect END_PROTECTED
