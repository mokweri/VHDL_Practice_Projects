`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G9gCsUMb2oBy2mmXvm1Yg5aEEuTnG/WXX1gLpoHWMcjBDRRjv1GQxdpquYvXUmuL
z/y9ijXycJ11lq8NvvEqxAVu+Byis67YYy4rctLiUuK+dYNOBKhuYuwlZgPJAwEu
EN+i88WQ5Y6R8H9og65bf7YgGI+aLilRHucAPgph/LNpF62Tuy0HzB6OMeWSgc1A
kEyZaqbvXRnLuRqNrF343brjT7E4ZvJb3PUTdb/DS+ekzbZ6Q9RnZnCqR7TNvKJ8
MTts2CGKgkqRb4/FxOKHp9mg2couMJdLwkRVOtMMBFGGrA0uYOHtGnE04H/SoZPo
KIkyQiXD+E2/yRyIuDOfqBRsvViBDe4EBSS10THO3M96JV0iFnxevGeObv12wAuW
lUpDuLRMFNemN8WMqS1cIFJZR/mJOb4i2sFubOjc+gutMbI50fUOHbhyhA3Y8YmP
89abYoPnN6fTAjXIxlyEok7nHJmKMqy6ktP5Ydel2YbHdPUEnmEWL2orVCMH7aFx
fJuEBR9EkCt5iguyO4l7tS/vSJDeo6KPa+uLKQljRwxGkelIA2GCYgaA6Tzrm/ye
BMNii2oCRBb4NMOfPruQqADmUqNBaIIZZ/J0+G6nK2KB8xJ961X5h9Gg9XeAU075
b9AL3kFLVM9uV5SF6m3LXdDehGc0kdhftCq8t7QS4qRD81kVnNL99kXMqQAQlyug
1JOLzXHuKF9d80myegG4sr067C2e5TfURgUSvk21IyN/SLrPpcWSsvcVEG4VidLV
ZYHnYQmN1NksRYb5MmsXl6SY+MekHYe/nu/OisILTz0g3EIj89rsQYSYkUmAXuXH
erkkvrobuwY/ApFsUPuXbrNSczUT44W+11RS4UufNzCgJQOiVZJtVN+pu1UozQWK
4qiaAJfK/nLS2w+tW1Y9XtaCMEbSoDCA6AiZsjXZRc0qasRnhn4gAq3YB2NQKYkw
F73aq+BfG2AAYvZNh5MTEW3OJAh6l06/d/flLxXtk8ZJRFJOzgqbtrJ4RVNYzpLf
o42J/XGvZlmwDjIh73/R7KFuI3RS4+wIiC7n1nZHS4b41nX3GCZaZtKF0o0F/LZ7
to31gQ6OvDyf/2USBAZrFBI796LDyQ63WKNGeGfqviUYGnR17zzteoybdHI81BMA
1egzJevNGUBoH1eeGBR4MTzzKY9/TFXjCpvrHr1nHp8LZA9q/NVhSYJA85W39CP9
8T7a2o3OYsgX6o4hK79l/UCe74nNoSYcLhjpPsnfhfWLDShL1n/9ixCjARtFtOZC
JiJ6gU/bkF2c0qbCtFgCAgrLXxMzZAl2aHu5zG8OU1313w/7ChBZeY9PnMObhhim
GJqJGJ7Czn1B2eFU+DJL/JNIzvPPWvDo7jv1QkmdrReZrjT4FG2wK4+f8UlQGKp2
+NX1I/P2AVH0WN2PT4vlHHB+pXrBfjoB7ysPB5bBGHMlR7N5uwvb0gYgm0znCE0X
3B1ALrltSegeUPYaUC2jpnuSdtXXCDJL+DSod0FKTQYeWWhYyulRuGaV5kOiUB/g
Va41Xh8GFkB6OjcsKD5qLxa9F6ztvfLJ6XjcmfLMcQg=
`protect END_PROTECTED
