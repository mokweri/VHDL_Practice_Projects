`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRsrbYChBgmCw64MuJJAVtU6bWZlAJt8nlWVXZA6lgKMjIfUB9eDRRF7uW+ohNn8
gLJmqMZy2YrzlCB9cR8yoE6Ng1abnfpD86janx5KvkSar4AHtuD42PI2Wf6nZrmZ
oahCvcpS6AGGZWsyW+km9mGFfBpxvTBuIruZ4V7H5BJKK2imq+LDsUG1yHjs/fn3
yKULHj3wdG1Mr+cS1KOUQtVEtKXshgKsoH1JA9znOaG+fy4R8RU4b3o00OWrrgh5
CfyRECzVAbaSdqjMyPgJ8aklp0d7eh0d0HPDQx1vWDENzszmU8DWAbxqHnqplo9W
WYWUhDbru3HMEEe79SdVFxzbpTCRq0cad0yOmgDVAa9SBpKJ3nDp+qjjTQfLPnM0
6bZXRjqob9QThxi910D48bigMByvDJnmK5Q5YSU8KCiEglJFPshJ6iAvOV/Miiqa
nxRhcjLaYwIl/opCmgWy8cUgr3RePu1//losp2ZzNEs7oI9xTtkCmQIQQKwmr2h2
mPkbVDNL1sm/trbX8mRveNQ5pOx6kt40SZV/qGrHm5EDzjATnE2nC3FcV7yg5/7x
JfFasRGznGQCsKPtW/4PySJUooEifHpWqME2qhUVG8E=
`protect END_PROTECTED
