`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvCuKm0QmtgZe+Lqg6p37tloHMLJu/b7EJtsOFrjtL/Pn7PMs1Y9/zzLUkuPhuJF
jzPEAgKqXrFckj+AOBY4cDPWEyMYuKRpBKtBUPCJBmAAmQ5FfBOWRNHueFMKL4ab
ZWdxWmwXjxLxwo4Wtn+e0/u7pMd+hUs6ieHfIrWj1HUifxLf7hK9fKa3G7ubBGXF
UkjoRgkJQ7Ck336yWMnN3+3tqYVx7ijpy8T9uoUNiMniXJYRi9hEyvp9Hp2hOwjR
o41ZKjs+bz9GqyhZB6igjaBOyYBPWrCCdcaS2d5tQsyTICl2eQWwmybyXQ9GSCdL
MW5czxK2+zqlhyIVrR7MXM9fRRFlB9MN6Yym4ZF04kJOYMBUoDqcsxzi4o8VT1BT
xhNzI+eYjt87k8uW/hO5KVhqJ8CBHWxl3W/cDCvGXQtAHBmEO2Fv1zo+Y4NyH6dt
NjlkPsKNhbKm/0+11yA3w/9k0uwURSNA1Jz1wbZNeQ7XdJONbtCJhgRkYWiz0zTa
ut2KbJ/4d0mxo2igDGrn4IWjM76Gv7ZD3vS5/sHAAgyaaqURnjiinYKJoGButLTZ
WK63YzA0cbdBUf0Oz3VuFty6TA7s5J2vyWxXtOHXed01Aao/zxPbA9ATpjtieYl8
13ZCDv5XDj+dAMp2gNWEW883ZMFNhd5LKdbjMwJrRvSuJ3C2cwe7E8WFGWgji/rP
GzfsLOnchms6NgeHGRxvneZd7NmZ5+hXq4OXhQH1ZDdGBb0KPf8oEN57PRSaKOWn
5hQmiWjIk1I6emiR+hV8gFReyEy+GXL0yH/weAWzgjMNCvAGa0ghTqJizCdF7NUX
Lg7veCE2MlAbMv0dTgjnd9uOvbU9Y2zMV2xB7iDohPH38MttOXfenCgo7C0YvIll
9CVBIbc3LoeV1vVGn7Ewt/CyDEDf3MUz2CPGQClmbqqD74HfXc3MdFPpygBwXHA7
cE6PD9vuci4o0SL2S9RR7jWty6FMlFGq5WPDI8HSB7ZineOuA183jldZ8xRPHLQE
+31GD0xwXh0dmxVOMMnG/sMo33CeCLxAMThajHixk7bOdSY120z+ni+Qg6ij4Xc8
DQOotmMP3w7JIGnbsiKDWSQKJVTR1tsbxEiFSP6yfhFlzhGrb2t2bBRDKJTbSXrE
bmGXrWexmb79tSc863Hl0dGdsPqkWSezS7Oqxvp7MKRX0Av7TFDxLBmRJlsQ/1SF
3+1NerQwyHEKmpIsuD9TrdcO3NwY5uS6n/HT5wuidW73iE8q0tpZM9jM4mGaYw1J
B2oTzVeljqT6dcAv5u4Ctz4uFj02AZt9d4N3hov859g2rmxTFWAsm/e+Y1bJoQFV
YQ6OkL6GGIlit4BDl2KwFKcJRNEaCc2J/0vt16KyNng3VrI7qoIxGf81wU82zaEF
3fNUwbk7sW/wWP38SaE94IdQ2TgbJcpHs6UsOhMpISN1Ke3zVO0O74aj2Fa2LPmB
2I12/wsc8RmDr8yqEc5v/hyT8zHT5UR58yBKERLIaGmsjOaPk2ISq3qeYr4WQIFq
NuhGVqDhTkgCVZDMTKp01n+tjzBczRctTjuaO1VbgOIos/C3jdZ/5WAMZ7Np4n51
6IDKq9qZVW72Z/q2cTm6Yb7tgR/a9u+rgj/GoYBRQYiuIykRUZ0YAsg87UAesVzl
AVxGwv3d5RXfnFXCGAGz+4+cPsEdCb9e/FSfceWPHY0rW026I4RrExLC5dEWHcjP
qu435D+4euY+vT6dgYAWxQ0mYIAHMlt1+0g2eeAuZDZQeanWkyQ72YW+14vcdyR7
HxqxF2nhBZ0322/AHbOrjEyFfKjDPHoSU6KHk8GyZ+MpxflwX/3G5DEtIG7GpKTf
IGDzXbGJPmuoSlpPniKvQuMIHwy0cxqoZmlXLtcQMCxR3DKxmbkffp4LFaYMTi5c
G7CNTfXqwx6H1m3JUmIWi5d189D3YZI20wdGoOlxTXCR2Reuz5PlZvW9kn0PRZEt
A8QiXeorzDLms2aD4zbYjmfEIKssAm9ORLWfQJZrY4cE4LryxmSj3MnE2rgvWoJS
Gx1HNCM77RF5Y0uUsto428QLGwsfwhwNNkrJ5chD0bPvv+bSAQ/np7cm4bkLHL8F
pT7c1ia+UfrYvNN4XlwcN4u+9pKrbei/F0Y99t+TXpcau1G7yHDzfUwdnnaY9JlI
lR8RkK7NTBGHIJ9eFPxR6FgxxQQq0x9zRRgS2VVbI/oXOHsT7dxowBSljIOAQIDN
3hQx6jghjpTYksPrzoHzww==
`protect END_PROTECTED
