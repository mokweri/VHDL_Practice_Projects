`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65wUwGs2zTX5qJQdspsVTEANpmRGEh3S1s2xFcUl5Xskcbryl8d2n8H7H86BkV/8
wBRhheDtfG36FvVMz1R+t8NLocZvOJGX6Vol6VrwDDsE88YuqrY1g5MCrsnp+5NH
vmQqlgrVSqYYY5o0egc3xeMZbGoZqhfBl/dEd/yF7l+DKCfPD2Sy6SUKZ0JZzKE/
3PLHMm/MqOOVuwCcUkf2FFTWlRB/6tKe1OeJSm9kfVCZAzH6fMkJnXUNAr2lN57p
g8t9JQOrkDnIAPy59JzbOJSicJe4PVGalscIpoMT5ZnpY9r2kL8XkPTTbOBrjqQ9
oOyPZgKt9Uu59WHnXiRB8/NAMD+3FXNrvSAF8UMxetwbio3zJjddHjqynqA8r3VW
2nklEkE62C6AZoAdLZrbCctMFTCbNWTiZXAqAbML//eIPmhbMqx5j+Ykn2hziljb
TCrYinhCDWBWiWa0deRtASvoeX+dK7/3cMrbSJ6OI7FmITObfSvgOZJYu73HXv+H
fGNXIEprWobnn3+MMzkWmrdZiruOvcM8tgI1MF+du9CLJojqAzewDHh/6EjTk2Mk
TQse3jGqTaNjn+z7JCY40bhY3+fnze32X+DzcOBnqR04dkJ+3rIz1Ef+OMuQ9SfS
pN6pw+dP8Qiy1Rde2i/lhKOsqiA4GD/XnrQaKgi4s0GEfK+7e9EeFW50ZLVJqgiz
hAEegVoLGZycw08BzfDyRR/PfqxWKKaRL28Gi6oEMbt2OBOtjtMv8cGYGVXW+p70
xAbm6op2cteWMuv/htGbgVo4+WEcRVlZQhTbI2HuvWOMxu9RSAt/M+74SdptA8xe
CbR2nvDoYgTd18WQ1lBLY1/HZot0gpJ/Oph3QB/RFNxSPJa4I7P0aI5apMoQygyj
quTG6KlJ+eJDXwus8HeFpw3Tg9/Ajw9W28b8uQywzETov1V43VQ9/W6FACIeuKMK
rA0y9DMKdeaDNeRi1D6KgVjBQ1easog+9rqU9/JXajtyTSMMqaeD/8UzXxf7C/kD
1+wK99K0ISBlLgitAg+qWZ0i358EcYXv7FJ+8BwySz1xKZoFJHKCGeG8v4Iqieyc
+P+K6pG2GpyLMQX5WvVPP/2ebx83q57EmsA2TD1FYSdMqQXKmZolHff7jTDh2wBA
/CmxJ9uKm32ZlchU2p/9PWKfxHSs0E+kzV9k3giCkpP662ayS1MnRiJehsZsmZiP
f8UtpASwmNMyosEjKYalqsObv1ph28D7is3DJK+q/hsFVrzsv/NnVpE/9W7vjip/
NfH63gr/zBY/+SU8u/o+/fH7cNnJ9pXBQmaXGY9aUSiBFVpNOKHBoFewCHPGciiz
HRUkK9jThuUl0AlDiFqtbf++/UBfBYdtViiy9GeSof9q7XpmXLkq4mmXuycNeA/2
0d4Qb9gTbglqK+55DmiffNOcFjjm7Aogb3GXw6u8uAfYIu9wf7bU6nzvWjscKpmn
8ehPIb+i+G7AFTzc2XUuG8ve5pbiSBc75uY1hBtoUgnmWpiEgEFnpq49/CeSe2wZ
gadyL6nuGh+5/ipf3qW0cc/uCbX/v+Jboh7YXn6BS3CQQ0fGsfuTTc53HZXbJpYJ
lCwwej0cZaQ96qHcHTYFWfgNix8aOYnfVxrCypn1VDznjYlT8CxacEXcvBkuA1hN
MViKxXMwBQVH/ocmE82hgbM9A5SvIwNDO2owRzZKTSqe8WzY9SjEdWGOkImJ1TVD
3KEa2YaizXNz6eG42r3Ho1xVhVgZFUjFzJF+uprNUF5AxZQDp4p30EzWhoCA7QMm
6PmhBdv6acIH7j4rBY9qnol6BuEGg5z2HXDkfJVbB50JM2l8xGTPuCwa32TMo+Sb
sSvBEPF69ZO/dYeiaRK3XhC82eUPTAZTDtAqPUt+pGtaYdGyXT/kJVWSEw4dnZ+H
oI3AY5mZS2+NmbMhtqdVYg3lhSp3ovBGMx5ddv4GCTuzTUnnXKJovYf9uo6TrHCd
4ZSbmuaJsEfzgZUrmDEHfMbxpvDfixBug4C3sbjoRlsp+UnO1f3I9lbqa7zpuVL2
GY8DD42bG8SRhaln1IARCnW2SGom5nWMIIwjKr6lsedrm5ziOT7V//ev9gMOoSlL
8AECaduj+RYeCnaen9WKRu6KHKkSkujJk0giG1OZBmAfjA8ALHD9w7p7s9quR2yp
UURIM/WQGlunKnw0Llr3nzrxBlr5+VHO4i/Sva01XNams/htS90Iq1fgSm8A4idK
9JY2FZxIU6cl0T/DHX4V3xB5DMQuLvDFYJquXEiKCnDQ02GvUI+s8dTgtj32GLJx
VmrpGwNmjJ5wMCeR0VBwaptB/JbyMhirrnREbDdm8BqMq2Eb3PcymXsQooTW9lYg
uc1e7bww3N7RE4TR5DeMEq8Onu+Uq5vGOf6m5uQE6lglvVfv3xGT4bOc39JyCNx7
szN5H/A6AcS+h/nEDs756rsCQ98PFO2qVvYVSMbJ1LhRfAgAfzX6juQNz/oZbgLM
E981wAUi+TCVq6QFNRkroQnb4CfTNpMsZavPfXCe2i4hB3FMMXumlSOsj0jvGr6l
Gdprjeo8aXdAp7soEcZBWEDUnnInno+z36qIkLZxgvk+WvDSR7ZJuxlMngXOpsTY
Tz4iUM8oVeqekRbhkRqOBIZETOsAbY5jB+uF3D9/kCNyQcgt3RorJDtZiVm7whtm
ec4G+Lu1o7r0Mux0vrhJIOlzaatrpIqGkgnF7muAneQ1LqvMaQ0bfh5Cq+03MgO6
4gS7aFlc3PwRhttSc1Yz9bxyodyXDjNRc8VABkfeIttC6ZMC31JiL92n8kBSE/LQ
zrgeMGdO8RUqFy5sWA4YH8Z98+dgVIXGNN6KYYxxFvcwe9aOiHA3wbt3l2t3N4D0
ZIJ95U+0I4WAPs9mT4J1gWCn9RKCPMTDKG4ry1j9+iXntW389aF8Q6xfw5SqWeA0
S/5+N7yyDjH8n/i90yjbgHFpX4TrP7+KuaI/PiVIw0MliEHgVl9EC2BXoXc/hyOJ
mldaMBWUfvgma6cXQe2/H/vMihMkD+4tEa0GZfjFQaZiqwgvkCHpGUTjzvdFVtny
WCP/SeojbtrQWBBrD+PfhpHwJvF0+BC4Hwskasd8xkKNuMZ2i4qh1W5K3e/MpPwK
I0odJ2UHUz3BpTpI+blqgsHn5WVjwio+KzfBdNNKrJwPPsOV5JWHf/pHteNx8ZAf
SVHc4JbtbBCD5JL/a/QLD7Df+kQT6LApsTyKJN/m+1kmpI4aqj90Kj2OhYoK9EF/
0dINfPrm9iPUdaidJszH2rP13v7TG/a+hsH+X4GXxusJc6fEC9YAX3szmYywRkEl
evWh17Pbqf5H0MwgiGsBk1+QivFNI30tVmcTcl8CN6jpGiAbp267ihA6Tu33jyD+
0dQJ0ysdhxpdWcSTXncNaUIRKHRB+XmLTjGH78MURym9UerpPIWfOxVLNGNrVQP+
KfDGGnnuyWCFXeNaWneBMqTmRxmZ9eRrk5zbm33UBdJWVFduau9qtrckqfdEihDp
DGLa3IGo1bkuqXt6GHXU/+PCMQAD4e5rlaRPn82rrDFCk+U6eYBWtjNvKeQn/1nO
6iBJ0jPBu6Nzyj+ptU3aDMzMelYQFaclzlkjglSh75NRSjIHwf+ql6mfzxUoDtJm
7LT6HBbsolfFhMWwmeGvxmOtn/ry2D1bYWUTXmQ9lSw9yCZ4rsQSa6VPf6H+QAuF
mt3GwL2C6FEavP/CKA1pLRGgOas2Bq2Vdm1leCuCso3iPfD1LgQxpZz5vmL/UIVr
jPqVy6Hz2YP1xrlOVPMWAWbmXWderDFqvLS2bLn3I0nsoFE4Nkhk72L1wyyI36Um
CpUQXTEVFZm5ynQyUpUZ5dwkjsnteluHs8LkTpof/o8LtHxOoqKTZSrw2EuM+J1G
4hQUc6rV10KTN/30aYkzAEXROabO9wtjjlXXGzveeZ+DQ+N1yr0Vccln6URk0FaZ
rFYTp+nwPZRRqPS7vaVS46otSEI1WDcJ9j0Uf5+0ZpPFVER0XNUqKolvN6i/3H+s
1+7jhvjEatM1mefwlmh32ElEIAksr26JgFY9OM/FR6n5Z0SaOaPJ5QSvEVPlp7Fg
w4fGeo23/cTfCXHJLSb9xsp0lEz7hFTU3znKhpR9az3NjnZVFuGq6RL1cR8QDVLK
o2fGbC9JuIBQ6eNq29TXlmHP1qgDpXOuC+k5wrKkeX1ehy3JI4fNzxbbU56jPftk
`protect END_PROTECTED
