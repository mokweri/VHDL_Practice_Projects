`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bW+bW9L0W+6bDC6aJXormYIxHtgDS1YdqHz+09OkW2R2Xneu1GWLZE0jjkKVWq1K
xsnh3Lk9UBH/k7jgh5mETT5fLRTjlw7tpxOqbOOsNwpazM2Gjs+WqwoFbu6VzDAU
mCxkYnQPAwReMd5oVYAB3b2WCPTVEYosaJJLRxtTMiBXXHYq2QrpGnBXGWf+2cyG
3TzE/8j0Ex//eo7SYZrb2oEglyJUgZ1UoeIMQG6GTUWIyBSPgcrlRztgrMVGCy/4
ue/91zj//7IE9HdBubsIqYF+qmCQIVavQCyGflM6HSShcbVpn8SnaizjtCULau2r
wtgyGIhH+lFZba/YGJbDHuOnShA9Jg7NGfColF0rnBFXXDkoYIg7qqpFkrlG2sFZ
QFS6dzSpw+S9Pbv98O4mfADEsEl5uaQMFBsgrKI4JXTOZMB3AgL7fwjHtJguuvfl
6g+XGQV2ZuDEcAHeW7xES6ZEIOgeAuc+1y7/65mLqdLNjMREh+rfLk0GxqeO7xpJ
zpNFUfePz80K49MxlCwdmFClGMi6PrL9l1sVjZTF84O5t57Y1e2VldhJlDbRQPW1
JeMx+63MfQSE/3Q8Xdpi9QxAU98uZ8Evb1o42JqSQdIU8CA2j2CWRnQXZNxRKcYU
m7VgHQyTRCwLeAd5izzQjmpm3huattZMl9cvBnWy2Yc7Xq0GgrGEL9K2QT4e9UGv
gI67qG/JKs2kCSKxKLq37iSEzFPqCuKxlCx36ggBzLk=
`protect END_PROTECTED
