`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
No1jU8YKOflaDy+qsKSQAGR3ED/mMa0x0YeT7dQnRaMQFjDfYu47jCkBGNZWZRAu
bSASLOKvDAj9IhMW/XPwEribh5vsWKf5T98R/OBiLhSJ/Y3KIkuXz1GODDmnRR5w
DVN+wglHahCxUlXerxZkVxMka/xMvxrHUROAYDggQZrozF2e7M1bb/DKa4ICtUOM
fl7MySuYadnKT4ZygQEQiCxJPLY4BDr23TNbWmQsSzm7p7ns8kQoJpXw1tOVdQva
j3+xEIbkC1JSqoDS5ndaEygZ6kEdvqMX0Yn7HJqs+opXF6J10B5EmRqyHUvCDa5P
j4+m6oGnQe5rl5Arm26TOvVyMfbaHCww1H2pg0tf34Q35KYVJr4c1RFZwTu4H7s2
ufCx3aYIpcY6zDezR8S6B16U7WgJZgz9fIip95gC3c4FUzgJzz/CmXhOJsJLk7mX
qpFL1Ky48vdOAUni478s16/Y75Hs+eKdC+CO2p8juKBKr2CwBFZf2RlkhPs94HZ5
VpH/4Qq6A8StaAEOVT8oHvdPAWwBdQ2m6SMG6LCENt3NxVCcDGoxxINNxQk+L9gG
iAfSD3f8yq1Z6b/yj9yVbn7ZThbj6iGY+SYkAUqZO5NBXfWl1jP378R/FzHWto5J
dtezmKN+I+9kbzg53rb6lMDKljusn/WGaHF+mUslJNh7A/+ZF73A06RRc2PhYVfw
kSCTrkd+UVcWVdg/bDuUhnuV8y3fXKRtDQUM2ZeoHWVqzPctzw4kzNsjgKJ/WKrJ
54m6l3TL/RbvYSMK5fhhW7fbV4GWme2/mdgayhqcwgzvsajVoNQk/b/w76cj0rR+
a2Sf6qv+V0LFzGw9O1IVDGmnhfw/ezTVOXEXVsqNp2MyYoJz4ZbTJ788z1Ig+4PH
uXoh+tOMXU5I92gDSSNcFzi6rfPK7K2vUYDrd7A1M4bp+GELUdplaIbEpjP8EavC
bIMrUN8tZFbUgvshTqwPxv5aIzPURXoOWA6kd+fDl4lWpEGNpBBCghbOyWnN+ahl
35tgIECGIxacWnHZ7h1ruuQoslMo+hjnyjqwdLXDfTCExkkUirsSNmZpvbeOMQg9
peYNbePrHGWK1kreKkGDijUB6+4wJTxkh73qcMxGnNDxmHDhmcttgZmbWKOOCvAc
WH6ZnQEbr5LZIimwkB6ew3pGFxWMizw1jWw9j9LnrhwFv+GmHZfxFltd945rPekA
scPdJ+5zG3aGk7jzJ/Yq24FKYk12UiSVyo9U71rcE+ZwHOzk8fRixwY196hChAab
LPfpX/SQvTG5tVcKy2GhqcCJSVRgf1CMui3k8cxQZPFccadkyrtxmwy2WSdv8nzs
aygxxbheek5gaxVVhxABvyiI/EmDSYqSwPV44D0M60G6whupGcU7nzkzPOWUX4AO
tPm75IBcfX+d6v9eNEePVpYBzpO/pUH7KB05002Y45XlXTwiPrQNS6lTRFdBZVbm
unlxgKxyQCXDs+rMkm/X6nKh5ieltAtQfkF30VRiDNj0V04TdPSG6c5gEquDRlzx
Af5HGJZBJzHo/h9KM94bjIOs+m2loqhj4rBgd86UPzFidIf2sY6G+b3JyLilYre1
wctk2AHQe51oiTxE8pdmGroxdS1lT9wGH/Lqd142zNAF7G1bX8MkiWPoKaHIpe54
Z2u/5rriVHkJI+tcGMk/+/uZwFe7nmkYtT+3iH6QJr3eq8Se37DffkRZ+5Z9RBvB
RrmIHztNR/DmZiqPRLZl0khK81z9EtwjwDafEyDndKTYqy5SSsypY+16LYutqMu/
xiy39LKSVhckN5qfi2sde8c0NLmQFCJYSFlpbbwye5sJCqyHKGxcOvqjm3M4T+LD
gYkrdj3BEZKjovJ/GAuJNrFic6KlzGEDmWkn4U5+BIFf/BW2TLhlNwvcsF6tNur0
APhUmCARXjOSkRxW2eI5cSUqcjQ7bk1Be57k6OHweqSONPrGzpj2lNePhSYLXDcQ
gLQ+XlA4Py3mzYxrctsalr7ZmF4PVouWfUZwSam2Wkir79/+mv/Hoa9VQxnwQN0a
RxznfWtDYjzzqIHRBQ5sfUN/43xt4QnPR3d4I45CZMvBW6rrybqilsNBJ24bqPB1
rJRa20xHDVSPioa1yfkEowWRcwRmciQwT+zQJjxMADGq4+T1ICAMnByIDkjRIw1R
4ogMtrk4MgHcMN7GD2e2F8K9EHgr5HhU3bjOWBrp604jELuo57+UrL3g3H4DC0xd
rbuchXTDjOWjmocOuunBa4fJwSOhQSEEuCAN7IL0ua4t1MX7CFGxArRX2zcRwsh1
ynBx0Wo9gBASK+oDAB6bUNIz4AEztHrobdG+o0nlIt74yLmROMwbbqvu1WZ3NpDI
diHtZW3FZgSC5NSQJrXhb1sY21VqD4ZXo6hdwGWqdP5lYDoCp6ScSXm9inz8J244
g14UzVe9dM6JtQaPbLgxF7Go4ozwsg2ATxyICJm/mr0mrYsCqHykm6pWtLvPUOLQ
P2cMz1JfOr2ngyPmsQGREjOJwn8EzqKgyJ0NN/J6Wf11XT19iL6Fm77zGNBZe9+I
ugCwp2g7H5oiNAWlF1mS8e0S+zFjaOq2SMnsSk4eruD+rQJ144MiwRmmba3elG9F
2Qa0zCzV7p/uM4qQpwtWRjQ3jscRmN71MsyHoDyUZJY4dLAOqlRVTC5+JjALXe8U
HhUQ3tYfS11XE9TiTOxSXr1fpkWDqNOz8FIWHoToxRjPq4RZwZng41FIfVrnY/QF
y1qwOI1Q9+Jzpv7C4XmrSJ8rYShme7tXbpwGptD/i8Q4kHOqjFt9vLmHn0Al25Hs
JJVHzDkJ5w8fEtyyNdwXCm2GWZyal7nXBY7tgbmpjB1KP2EB1Gw0IpOqM5s3iY9M
3CnEiDzQ/mPP4/kXmZVaKsx78ZdiGjYlY7yOZJ5Peyv92PzX//MAwt0o2Zn2vWEm
/hjUMr7HjyYt0oY1r6b2oR+A/txrwNwmIE72OaZUCGP/DKgjszsUxD1rggWQrjg2
n8Hrukv5908AIdyVWLlmCR4grK/UicoPIMghpfS4gzBirZdDZNyx6OXohT7Foq8N
A85UBcpjpkW7RUIJaBzMUrxiHoTGBZl7z4XsaqgVh1PPHbw17Z6fxe7d1gCoNpli
vfnYYs5qDgfTdp3PqTkYoaW/OrAi8NK3PwydnIvxxC3AnazaMaApZp++A3TXkAWY
SZp0o6b29+kDNQcV+NOLUewsYEtqYtzJztVloRJW/VeRv8ShCWqbnQuJ9jVh2YLb
/1+x8Zvp238mXAeZORwY4M0LrgH8CLxTuwstuTI3Ga2wU4Cvme4419hHSJnh9xZW
Kbo/dzMYgAlsTDQ8xpXE3FDM4OMLwjXUB5BI+HJD4UeX8k3B0hhjSm1uDoPyKWWg
YJgICuCuKjbBORjBQ6x6aOepVCn9yfJXcBr+XdfzpV6hb53UhqUBpxQG8H//KVJW
Uza5oxwB4CUPbb0uWkZDF18YXYcPI2D4I86tBkXOxlfOJ0woP7oJj6czaQ7UfrLZ
76BkKUK9wNZOW+IMAcmpLbyATJ3xBVzByiLNMkFvYxR4iK7ydMH1+VxlI5JP3fCe
HPE1vi4TM4gO+UglwlVs1SyTj/YHBfJeIkcHUnOawZtu2l7ree4ZK1vjrpt3YA9l
HXW5O0ThrcorKkCzoBgtsstk/yYDxo/DlQIFNlhHhbtJ6tTFHgq4h4UDd/U7rJXA
e8u6vN8K+LqFNxfoyz4KYreBcz6joSt3vwmggT6OqbvrJcxV5YLnaxLS87rni1Ts
c7rWzgBWvkrmHkpk548P7BFojIRttywWDPGiFwNpPX3+/AqM/YS7AgMg21gMEe2f
X/kvKwf0/dot+p0zBME56lT46J7kUXeR3QamDbu/nzxipkg978STl3BVzJf5T+A+
yBp2Xyk4tk1s7aik1l3LYXl+UTO4UBwvSZ24cov12zggqJKcj/+nRLGatIBCQVkz
ijo31eWaFSFeNfY8vjdldk1HdMNw8ZEY+/5V+mPBcoZgjzpGhpKmXRt/E1ZUd4lD
CMDgqQgzVhtmFmhwXxwSAYEBaB48lV2d0B3Eo689zBg8+UkqPRADHqwQClsD/1Tf
Ct/w9nX7WsUol0xaWVk/1gJCIBGBdx6rwxkw/W95eJOcLLonINVYtyfeL8G3Dgv1
CinvsecdTzqtjK715u20ZiLZAEYgi4IzrmfkXGy8qc4HhkVW3/rLXdbObvyfb0rA
G9RHXwAbQog+j49BeopS3g+3gfbFX80pnyvCaLbZ4OCt4Rid73BW4Rl8iKH5tnfs
TA7OWYs8ZoNLwzaMEWmWm8nMS9C0VXTFCwH8ThUnhJC51KbdCR0WQqlHXi3Qp22d
Q5GKPerwawtrol3KP3rbH+lDijLDOSkKMQokelqovH0Ul4cmVWckq/IDVSC47ckX
uz5qZp/LP9XNC2Ba+RMEbNnJTb2GFB1HdWU3YbH3QhE3eHEwzSa1wwpD7BmD09o0
Fe/FSvXtxakGE+fhdJrZB0uMz1F7kGP3MX2AAAstwVTQ2gnHB08cBSWXh7f8+ay4
Ng3KQNu9LXSOqFfVVYB7z+VFriHqb6AMJzvjJzfDg81FC7TCxm/G/whgZ11RX2Rx
Va5qwQ1JK81743VKl1lA1/QKbhUbTtC98xsKT+7Z5B1aWeC+2SWlGjDF64r68WhN
evEqF/WJNccAI/2I/j+xyUNBcvsTJGEBsOH8KUSIVf4BRZiW8reYiImkaYEt9sz3
/v2Qtupc0ZTuy/mX8ZFJ1nHJBMZzhqEnifVob4ONCyvt0MVazhJZof+4DQn3ib0/
zvRzrwSAv2gTkCZhpDDMsrsRMNvWa7LXUTTbpqCXLXWqINJhpbcm8uIbn7CosQpB
NhpxzoByJg2c0c5Ic8tj0F6naPu1vf3gPrmm1HzNOY4X3dndL7UyBDS2l4qzwJVc
ZZyJhh2nNBazgFwXgBI8kIayAHO8IXSyZaFgM6BVj3MgwrcwKEpa5maAMTBWngcJ
eemlD7mV3OUGN6nBU0rWJaOalmuTXJJgDMjjZCTwVWYFakTPNiwHmRuCUIHq6TuV
4GsS1LzQWjiwvG45uDWtMcaHDPGu3HLtN2MlojdJy94Ttjv+ow340eNFOmKxnLtk
Tsg9LfOq+M7H0sQM+DqVQSecteRXqR6odCkUZNlCuvw6STvgVv3oBlHXWbuWeqnR
FO4zNXKzUlCO1TX9wmYjsJ0mCBtR52W47HbICbuaOA/jkuNDSMkS+Kb33QHjvyZM
+8f9BnvlxK2oDZdKsCuSfrS1R6ae99IFHnJrhaPeRkamdoYkj4MEOtM6jrrYYNqY
yYzy7pqvjccfydqR8TYujXt23767XGGDBv7oR/3BWZJY7pjIVFdyDb6Y81rOnZfV
dX5QUrP4vDG6c4ZS6uZrgL8YhB4ln0mGMnGzMxM3WRGJx7106ofqPxsd3bcLpFbt
E+pwMcOItXk41Phz9HSJ4S3p9qQkFLVpj1mu0tNO1WhiKle+99u6A6tWhizSAPEZ
malgQ9vBUnY31H4RNLyNdrjFaUm/3Vij+dDNCh0RscYyurcHNkbtRTPiDyfkWF72
LZcnbilH+MIRto3gkTQLi0vTkKHtJb2Wh1xTjkVdJDMGIydldmgj8ApXv4FbFDAe
QANyCIk54W1+JWGzNOmD0prJuPC/U5/vaR2K9CkcD2aqPClVRqWN1LBCdAzhmOkQ
wsXG5hoGbh2Q4a3k7OQubD9JfB6jyb4Taroq6G2vGgqoZ/eZ87kHC4WbSH8meF+b
YWBDSXDfGy2aRrE19GuNOFJ6+YHtKmdOIbxaRvM1W4m6CXKNDeR4P2SQGoIJXjJu
3DtW4qb8VTpSJm3SmkSWRl+M/zIKSV+AMO3Wz1B8gbNKq1RcR43YefD1QJm8+lvR
35DdfKDnoArsYj4RQ/2mkl36DBHpdw2X8AbojOPW+nY3aY+gBcRzf9DfW7q2nRcH
uU6JR7UDmuZ/iGutrXRHlqSCBEHLREkmBtCIjYcWlX4=
`protect END_PROTECTED
