`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bt8YUc8SlLHNs80b49vXOCN7YVTLe0K/5yUOzQzu1KeqHl6+oy/zK7wvk+wuSLCn
NqsZqxGRVPY0oSIA6Fh9oshKl7x7tIOyoiLh1rCf5cq65l7V6F9Xsi21PiUwW6/x
popofXWn12HkUhrHS5rcy+2tDiWrfjXvzfgE4VgYvIbVnPPgY6I3tvJrF7x6BrT1
ZHiF3DboY1MDo0WWxFJbq9nPv3weWs/EF2xiqOFVQ2NLOjgnGcuBMl5zTzPWnsJd
STAdSM1s95XLyY24KxnRTIgHrO1YfLXU/5W3kfFWrrqtiRdw9GDYdH7enYiBMHR5
/kz56refSPmqBCFDnmaZEeWDvKr4FWw6eXMXGPmqEUn/DhkoNooPD4+pEXAGt5Jo
fqd0p1hPhSnX2zf0irgXpOAiNburY+iMoiZ6wwtoZ/rONcmWp92/1/5igBdl8o7M
eY9MHyYWyu0g7pvXHH28DLR7uRLHWmRPyRU8cwmFIEart9BPNj/Hm4bLkiXt0Pjr
`protect END_PROTECTED
