`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y7489p4I7D66KU5Shv9c78rDCM5UAl1j7iaIOvU9giobxNO9/8kK/RTx77zosEOw
jqaZCCkKNZFhUhO+BPWTSvzxryKz5JIoTLhuPeUw8gyJHtiRhcWgrkHcwS6bC0f5
rXN5UXjCm7MLPHyfUgVUTZH9vHaTgmYYAqm1dFfioCQT4bZMrNIoiypDpG4SwqXL
Qx9bk1UVe9QvdErOLGOUL9jliQeWPBKS2ioBTCYkcqXIe52kCGLUnGk2iWaj8wBp
bWRhQ9JUPyuqdsrrIrdcusJAJ0caaDn8gDcnKCX5ND40kQdMLTTUcPX5zDDX1SOr
G3YJNHRyfKE4XPmqcsipOzqCOQ68HAzAzfGbjdcQUtOxJ4/IjSfG/qBTX2Yfl4UH
duTkMxc8QGKnEm4JaCkT8VmGEIhUpOkGEla6AQOoNFPGeaWruWMX9MUQonT4WO8s
c3swqyJCVU29FARcX1fxLXSYmoCz4EyxTZP8YSiNdk+fWQ8Zytro81RI64/dycnh
3Ds9Sjxiz5xk7n7Eyav/4NyWSq+IYbRSV8MfRCE9jlger8owUHhRmpyQ1XlpGTNZ
DTUkxlsod0JVqRfqbqJvKJl2/iDyAupKiYy1EhqFOsuXPoVZbfCtHAwRo2kAVnUg
aveWnwBHfBp8W88NgL5FWUYsVa4mhBe/tvtZr9HKQMY7et+S8D45Fg7ttrhHlXSy
MrMO0raTLdNPI1bmg2Sxwp4ivm/GSSnK/DfKBtHGpJx7GYjbEM1+7iUxDWdXXekO
nlh8DkkCzTriIt3JmpnCbajzHHGlLSAEZNeaOjuBJaAI1C6jln8vU8nMkoih0ZH+
Mo4f55MsGy1q2TlMe9qKMwtoH4l4qeeycmp8LHYy8kQpQfoDHqA9USz5w12tpLyJ
AnyoPhWKfKDa9ZknyKBq1tMFTg0OX/C9mzhrlkDHdoAtQnkUTu0VnKlOPV/phXnN
bwnZbKI7ckG0zDzuRJ/AqabBsz9ILqyMUAsHAiewBCEaF5QpJc7ZszECUR8/2VJE
nmpOIX4/TESaby9LgG8x0t5rSwAORYLV9L+jpD+3ohtVaW/ojfFFlBsgdsGAki66
LdF4JkzPk+usMq2tp017BVOd8aeAbNjQcX3VKZiUefDpPDqLSi1g9lQ59elVP/nY
KFoNYOjPMyja+cOge5ENvg==
`protect END_PROTECTED
