`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDOXxfPcrpARymT5wyjEtUZwfS+bEgB0q3ho9s6DuknpjLwXAP5/9CrFALDs/A+f
MwCz5YvJE3jjY4ZNwHB4pqunkyfK5veGryyhaQRNmFCTbG6kQahnNNu/VXF2T6T8
zdLRLb4e9HvZvc/VLFSXX8gTYn58UcihiTDg5s6WTs1zNG5ChFt4obwcQwwQBK7z
xcAj8ZHE4nb7bXcTgmLHByfGM49AWqUsytDRbIoM+9Fn9ba2HaKV1g1C/nMB9/YO
+bKg40JnbZG/NlMJlmnnZWZ0zd7QXrfbWrsUYviSEPAvIBwVV4KHHQvHVuJK+xmx
9DWGa3/qAwO2Tf+/QL3OjsSBcVre+IrwybrCLYL/+SWB0dDhm190AitK5qP+TJhT
AWYwguGeE/ptbeSPEczkUJMkovOj5dy0LFiG41EWqNZ2nsfYRxfbLq78y1aUCdnv
oy0LTYIEGMsQ1t1D2OukWrQCU/lsGodkQiw25ukfrh8rS4apwPQ1Gfxsy4VEN4fT
yKkb3GF0lgJrrIrNe/6lJw==
`protect END_PROTECTED
