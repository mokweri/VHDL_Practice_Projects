`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJ8era/IwvO2CxhLD20TvoSPWiq1KOpVxu0n1BIvbaIy1W3h3ZutQ7wwvd7wpvk9
JGjpglJZ7d080ahoRg+9qRow05+jJ5lGuVHV/j1mPWlbGkI5TgaPLkhKn2TcPR8Z
ms1LdyDi4ytLjyDs5ibGbmnLDkN3CWwZaJyFNyZvgTOW0nlL8FTsRmnyhMCxCGfE
LHWgx85nhfBHpanxCnv/2xkrTMbIPlsIBOLq4CWWF/6DtAf0ReGVcB491zSIOz4m
O1bx/wrC0hxEoS5VrKHcuwr34DCTdIp06CWo92zm+LBpS6GUX1raCZviRZ0zrRkI
J9tun3BmlIqrnJjZwJELVfMrhq8TJXnDNXTYCBqVeTusempG9YHZKZs8s1NsLbYR
3RVT99ltHhIDtPl5uCtubcMqLAU09z8uvCV5/rV1pOFPfwOgN5Zf+PzLtlHuHnX3
Q5Sm58qTJ6YEJ3LqdlC2zsAX7P+/Vp1cc0EXtdJEoKrzY0Gq5TUFqoleDqbwkytY
E1mNHeI0tcOIzBuIZKnRUzRd/sYrpTOvEvDfZTL9l1IxYjwdwE/VsTn8rEc5C6PV
VC46aftrh86UltBp/xwE3J+AHIhT5WvO7HWgC+Cxjm/R15DDsvQEq89X4GDYOwTo
4feEGMvY9rhzmqXIaQy+0omSGKcbAmSuOVkinm2l7zqpZDAMan+wNF4PiH4bgXxG
uKrgQecfa3ESJ/PrRwUetoq0vcPxhLdBrM5gwiAVOyWNdgjIEzzCI5eiKouJr7mo
8ZYjoqaMBblY4ZAPElgRlhvSlu7RInYWx6vLjp2cCO7NpNKo5ug3u4J2/UQSRQ3d
X522C6LqIHVboWHhk7/jvRnP5ekyHcvS7lYtA/N2RJcnGZAZnmRo3amQn0WaY5zA
pQOWJ/0TGIezxuF0jeEgGWTjKb7fOhM0m10kh06/WbH3o7q4nzsZKGMPYdeWZpuy
ZfxRzSRebAZVVZxoF+NHRU4SBRstWxRQ1ojq1Nln2nEvjuqc+0SMQ6szheiiu/x1
SGjbvPiR3yZsNL1T03hWLmBsai/l7zczMnoYlPzJhUKLCBU6++ajnnHhaZlQY1s1
PLZYYyYgnzHn+albFLHC2Do0xbmdAVajP57i5P4jFCT7tldEYSpfi4iLPM20gi+V
Y+VFb0agO6LVMWDpqo5+Y0jcntEpbt5c8dhlOTpAJt8DbbvvLoIwiWbGXckLuH6C
usQrun0PnONhFcp3OfAhC7JuDkeEaITXB8S7FMzDgdH4XfMYN0iDHqLYavqk24qG
vWk2ftXL/JhUQN+/N1ljK9Q737o0jgVBsboROC4Z4gd5afwm6OsKhYDdxKIe+EMP
WETW+/IaH4RdhnqsEStVC0gMTqBDXXt7+uDahA8JA4nGEIJnpvQzmjhZYUkCnoba
msdT3SLkdo/8HCyl9+Owh5BjWmL8L8CXAGRSJ/njlIyTz1/kK9N/YcmUldYeJ9vK
w9eTMqsFiz6XwO3QOaNFoVYqlUHg7CpzX5nCy07FkBWPhtFMtCcyaUDBMZCU7bzL
8Lt1Gvue8IG8BaYYH2I7H71Y1IUa9WyRVV9HCvgTw/mEzgSzqvohwQNwIiw40eHm
+Ys/Z6DX+6ezf7LkJza7H6KSoBEfw3bDdGwSjugj5WtmJuyUylmYdSKQcOiU0hO+
TCuQC0jO4F6xp1ccYOFvL3xvz7exIz2MM7m1i3vcCj9oGSv/I89Zy47cbNHUWFov
IIl7D/PSCCEcEVNH91alUgT+RrBVQRHErP7Q3Otr4ki/0SsEuluCp++rpUWO7rlc
XKgw2u/9+64dmbEvoZ7r+jeWurQcqAudELQS1eOudCFeMLifGxjsm74z5KD5KqAe
KgH3o3OBayJ8ACGix2Z9KeEU865WTXxGBX/qPc9IiIDMuk8u+hMA69f03PMr92i9
JBm0runH7bPG8y+aGbEvHh9mCAbBNQdX4E2iHfVWVm2B48ZpFu4/sURyVs/NcSfq
nDnGU/wJK+4i4v60AXkCCFoXK1x2ryYPWXOUqwXLq3ekrdvIa2D0hQRifH3PHtC+
BvrhJOuxt2L1cO2hh3z/qugsR+nMmLfp2/kZe/jfP3qZ5srqy74HkAc1b71/QTF7
VzjSoXjkIPf6chBF1ij1EASgIp4gNVAUm2o0rxb3uPYEaHRNZ7IBQjAP8o2eaU7V
OPtwoodBsKoMYWFmV6KecV9sBnLbd8Mwia41+JBOjHlK7kY0FQqp+FFDkIrmfi21
qMJCDU/RC6tbi4I5yYgKcmzJLBo52w+18tdcGw229UKSK0Nm/7K1t7o5Rzl1b+Pu
Bk9H7DJ3nlpkZHvtddtZ91rPcJ6QeRen2fKUYphqv9pkyxhNrbN/aDPguU+5XyPG
nh3OBaijqIfbVPHeZM5JyojWFxOgvs3QqMFD8NKqtYXza/gurdwQysNMBdhqvASk
EeQ0vVnrFUb94sm5607xkyy2FIhjmUI97wEo2FSnixYG+XtBVwCyeRB96jkDmHJD
TB6U/vucHf8GMfAhLC6duX/P86fdGMbz1uv6+UPZs9sV0t+xpfLbebYc+uhhf165
JPdwxqS8OHJNmjGlZYHdwG+eQC3NAGPT2nc+kLFWk0QhSTLtwCIKxwfKFbMem/Tk
Ni11DWPm6DSpmZFwZnwV2HJBSW7+06uzLp1DrnsaQTZsuEvibBvItRqfk5PTuBm0
3/tP0SUiwrzhyVUtlg5uiG8UfajQfexhTd+jOutgKftFRM1zNzPmF28KC1sKl1eg
Y9uBiQNJv5iIzSNLl8J9T/RW5EzgXK9NeFmUV68Mz1RDjGh4j3kHeRGtDEUmzn89
3stPdMDBvvloB2iyqsz6twhfqNOnKMWAqWGR9xmNxmR+Qv6Kw5eqoPtI/eqsXso3
Df2E3dNmfLl/aYNUFD3fW2ztPiplT/KEQ+AK2ioEkY9tHty+YIz9OGypBjTqvH0b
Or9IShxVGNKGSFSr/qVwfQISJgj7aI4cCpnAQWt2nV9Fh4TgWpvAPj0G840R55V3
bqawXspcUuk1Pn+rKM9YGVkIHI+z0ZTbL2quBYapz1xM5sSxSGtTouJYhRFrBZ7d
t4rAGxb8UCZ/RRQN854XzpjSXQ0Ekg11hS97ivb32ypIBAUEvJp3TKFB6STEXMrb
kZHw3ZT9SdW+llLESRcXqBEPsxRMlROX/CWvEqFXOmw6rO28YNNoEnPg2AWjYTn4
7Cmcr8TWBVm+xMHn7YBrOsWm6m5wGuIyCavXt38aq3i6uVNqnPfe7GbzZbOnXKiT
zBDx/k5n8TQxryZsxAVyB955+V4tQl7dg6MLf6glFPqs7nko8dATVTB8njFeFgpm
HPinEbd/2zkfQA35aOhc0GpSqOzGPV85xXgVYaTXnjHqNBYnsD6w42MLyz3omRgA
SKtX/8GXef1WroQzWG+oPStV54Rv5fxMc2F5b0uc6u3uH6pqWjN3qmqAoD0Mojdq
OJAinHCUlVq+E+TM3ed4GBAw8lZWx/JiArmJyCZcMslyMUkbio+0t0rZPKHm5XzR
BDInNpW+XVW/QZKHh9hhuO/wxDmp+apb1zbgWnlISMlq+WO/Ar7kRkP7ObZLnztP
YCK1MAdvAVGozywlxeQQKuRXgy8BBRT0XWD4yQGmXkaWJ9X8SVVNTZUNYcq+mnxG
XTL0l+o75uuOzxgO6D0Q2aLRT8Hrk2xy6zEzjgR/W1elkywDVxPeLBDTg6WsqJHd
QZzh0TByJmL5H4N5MS3pCTK9V6KGofZcUAUsUBvXe0q8/TLaxkQSiS+dBx7aoEi4
OGgiflXss8mQ/UPmI2NnkzqeMF9e+rBohKd5VO5UjTWrcuS1zCncVswzNnbpyIq+
JK4BBtxuHmfZysuhJOgo0/X9Suj+jg3cAiPlH8BDegDRkya25El/A/UEEtidc5Ug
6RqrKI0szk8OfPvd8iFxaNCzcv99OBZAWsf5AUlsiBRcq05kcYDKLZwc0+mEPm90
ayjHdO1YIB/fQBIkhlZ4jE/GERju4D85QaBZi8RRTIdbfpeyBp6nd+bpOeChwinZ
RPU6klwcvU9o8jcLScHkU2MqrSLDkYfWSBRvDwWlfr1DqjmrURtiyh9mzONqu1aU
Gqm1N3+KGwAgFCCYCDnBjzdpvJz6FNvpK+4KBuQ6qfd2yBDzm9Kff+oA90yi/dTO
9X+EjG619h3REHUqoVlzXWppuXK81SlO6Rh/B2SWdfUbHUV0plnzhFNRKVF+YFyn
Zhi/qBTAgKAIPh0YoceRybgYkLO8QxANgI0dGmOuEYlMuXSPLeEi8+t/34EJJcP0
h+pZ/F7j0qZY7qXjTVInxOq+t3Pi/FG4sPcsRoMTFZmqCuG6l8cY6SmJugMw5sjv
uP9zvgzLQ6Rm/y6LUNyPrdhP1QU1hZ7K40VDkuhxMEfqHBVlvqMhTaYOTMOOXDx+
RHqJbmD0ohyXrYv5w68+3w/lA2owha4jBL2F8W+NP7OfEl6S37r2R13u69dqqsx9
fCptFB0UO+d9q5whLAMeLMcxU7/ePsqsQAszihIr+Z9J5HwzhtthKUbUAcd8Ni6c
U/r32xL4DGrTaOAVD+Y5GiG8HUc8Jx8se8mqm/jtWebCyh0NE+E0ev6Jh584A4bU
UmHfLyXFi4ey/1+MO04sGnwaOu+qaIvVUOPkb4fCq6wj6QXGau1cqQyc0+7dRFUZ
BAB1SmT3OVamUKad9a2Q2M6VqIC8+U6dD1Dx90BkDgdfNCFN6W0qAixEoT1KmSCO
AUXeKgoAIL2iNcbcO52C6aYGNDN1IlIJMpw6XkrOc84fNNto4KxovDFz4VP37WqH
NQ6OKblcpJ0m7AMpiYi0W9I+T/qy7hQ6lh2wdlImtDdmJiPNb6bvwteUTWkJldrW
QQqpOSq9iPWK7uhxkTmqXyjWz0/Mje7aIHpvP7wGK9oHasT+2tIla7ydv72ELqE/
eTDziCcQdhypsz+2F3FLm/qIdUf5o2Aplhjulk4VVIidQS+6OhDLJBAXqdYDpJyn
9UO/5P0G8GorLNx8VNlRF4OFgN3q/1xHo/8JcCYOyAf6gxBZ1qCk/SNa+qIgxBkT
c4/wk5YP52ziMsSlmb7EPXOROiZAMG6beeiRgmsJItI+SzJWX7dB0qG/cziCKtfm
UAq7Cs/9ynSH+yQMhBYU1/HKzBFy1n4GPea4Kfy6Ixtkyv7QvHHWLWZX41/mhrfN
jxc+O1JQk0Bqrprla+C2PmZTaJPQTxC9QNTsaZz83oCtYsuYJVZa3hcQzixwtV3V
mnVvSW1N3gHqEHwx3CJZJn9Ua6R4y0KIzvBTn4ycJT02Cn/CuONQttUsmgpgQaVN
ijXUwiC+rlx25g+ojSTTa4t7oexHxqvtceMEbP/T3GVAZlkZ5Y5cF7JvhwuoihXM
33LnRdTO24SJdQFr3SfekzokmNoIfLL2KSv+dTB2juEW7VUXCZk38fc/oCbTQpwf
mlMhK0EfePngFxAba82v3ZOWGsNUWv7uaAEYlq9iMGuXgktqJzdbA37SuBlzi6Kb
RYczgMoqWlVcqG8jJzGPcLVBL5r24aoS9YmxMQgP5lxmPqQl7VkIuLbXM8gEhPFj
oB0hswC0d7M+8SfTCdkoS+T+IQ53ImlXwJK4a5KNqVXvPHRhjbdZkRKrCigsOXSP
SQTtexDKb04iCZNlAFyOKzdUy0tirRQS8ueYCD47P1GNfFK9MaSC3Mf8JKzTGpfG
Reppv0H5bQjPAPY3WxE5csTlsz87k1rUVP6Zw13TbycxannXXj6xI7vowa0BrFDw
iq45Vm/ScsCsQ6jrincFNKZDnaawe/J/yY8lrGtqioyAod3mn/Q5FTp2C1ebDyha
u2/f8TDjb0tSOEYrksGp3fruW95n0Ij4CCeBLkRweCQNg/x4AG9hzNgqVq8rZdX8
DxpvtUuYg2HJkzqjCuNzcAqjk2/90VxPPQt2poDin52mWM+tI/9eY6bXTteJSTlW
cZVFbCwnNl9I/Hk06izIepHiVQe3DAvXEFGu3av//ZGKLZi8g1GG8uGwmXPjn7MN
+Z11iJgjUjpodKzOP63RJwUaHnLQQpKc0ltDJ+Gd10rOI/OjiwsM0tFs9LopXK3k
pPj617/nxMu1HYP1hKjZ5akUwFf+Y8fpFcp9lh5pulgg43qaZGuqIwnjPZi7Z6dY
guYvCUCaNxSFng0M5aqFmmEvN7jKitfyAtuGmCwSnoWfjFQqabN84sdNhuzEn2Pe
aqCQdQ7P/m+xGyZNg0A5Qvh3J4uhyD/UNucTmeJWLDCACzzQSMylZBAI6praVUhK
B/tE2jhOPqI52cskMM05pJnoh2lLJ+17/SY5fm4OYsNqqwmOtoDuM6+cWN2VBNWU
7H3SEAsVjBFF7z4xsi7XcPvD3GuXUH5x7kFzMZS3+h3J2lrNBeKulymAeLo2Jsap
Ewu1CA6VTvFJckFznAbTOgh6dVOhcNX1o196NbSBKdiWghOrAweOlBvVRfUI2s6H
O9Bytkbn2kTt9UYop4srCMx6XUz4AHtwKmWBD+w4jm2GfbMShrHurUTkWDIIkBMT
IS+5hYUysVpD+nsQgxOVyuqABVTGD4yfTioiREl0FZ90jRi5ePUtR567OFCaoLJT
IYmCoWeRLj+ZdukbJyV05Szi6RY+6h29tX0GYR9uh98fLeyzqwvsMuG5QlWV3Tn8
0yH9NcrmvPPbzMhuFywdFPsZFtLurub4zWGHRcmzJRTkjk9YpcJ5tNF8xAoIF9z7
CD/jHuflMyp+p+U9j9wOvquKDNTBXbJM775X5/3CEtdbu4R8PnkvHbbR1At8askz
7Oab7VnFZunetDoT+B3Sagbh+YLx14Vm80Y2/P3cxSa4wcW4ezN6hsShtFpY+iPc
f3ehMdPaq1cL3UG3G99cWfUn93jWqfJlXxOrLArFoeJnpp8OrjU1/BfhSiPWJLvL
+0RTNpiKoAbxYhgutwr/kdrBuz54N3YZSd4E2IzIS/CSv8mY75uA50LOAKzDoatX
BeAAUjRPwEK/1OauaT/KUQosAoZCQ6+hVfSKmlxEcudWHMxeIt1EnE7pOI7DF+5f
Y2sYbURopqnOYLQ5eCbyASfKQcPS2hWLvlD/fhU+Ttn6sW1/qa0csaJqL1Acb53y
FP7VJBSJ9D2QFE/kfuo3lgfvrBVY7BdXVrgUORf0/Z+EpwCiHlyYY+lj+4J98Kjj
uQdDyWLWkaLc6VYybzGVzJr1rh/gDLydlVElTSpBhAjJPZ2l4axtNovCNSejqq6j
1txfuGX7vMvt4Z6ofwnDzBRRqjOinkR74SQv22nLrE/vG6my7LBV5v/pT107pzdG
fqtsCvpATlIqecLQhApcWFCCzoVPbyiAx0YSoSiM3DZxt7XXrXW0qDQf5QLnhv7P
vPsQpto1HnF4i8nfl0RbQqxY9/12ZdudC7Ju3N52IhPY8D1mfOvl/byZj4czl+du
vNb2NUbxJdDCUosRg8X6Ows5UFzOBPXpJYJXJEHxcOWSS/ixBTLVEwOVj0D5dKRw
yTj9qpwB4B4aZV6Bj8cjRqNNX8rWe7Vdsf4R/ceosrBmFDmUtHE+x46X8GYBD9FB
fpgQCxjIXqIyURIv38m0P3U7qzI6h9jR+zb3OCa4hvEja0Wt2+0rijb3SlwS8IpI
II62Zr+JIZizmf/dLMUbGD0ZSZ4IgRL5lCrG2BnK/nYpbOq5V3FF6IYTMGf5Gp17
B6oJvTTCx1pTSev+yI80R3lVLmodcrt19TxduXs+0PPTpWdeO/+39tBDi57yv3Yv
WmfH9mAY/OPuscqqP8ygqFiUFFMqgYSJYocSOZ9NybawvDpW1xeoEN6wIg4UUUQq
bLXgHi/kAzA10WRIIUUbYrmPBmCCCCeH2RsJHnx7LvsEcNB7IOeksCgzc2U3mlAh
Ti6izRox0x3/7Tc5bvvVAJ8qi2x/f2r6Rtvp6AnhgZjF3fsNZx+Mxjtl1RWhe6+T
OkHHdtl4pkEmF75fy9wnKwOtcfcJCzunmCbwljuGgE6jmVCxyX8INecjAmgsAXTY
PM83Wg8M9yilMhE0NG6yoPK06nBAr8B2v46K1l0wUGE2TFzfTu3oqTFwx1ROEZvl
R00v3sQaabTiZBXJ/yhE36/WM7lsZ2q3oIT2lWUbDvp8MjI1vfIEw7jmJ3suyYsv
jTOkAci4MDjug2GmbKMG3CWXsjj/hQ8GeNjD4WmxDciKZus9TaxxBeLQ4jHhnEbL
yvZJFqlXRQgUQBLFU7P750cs7WXFBsGKWpAmI05mF8Q/J4/WWInm1BiOIiTFAU5x
8+O09Ymza6I/BoEa9BGZgbk6z07gabBmkX7SagSTuQKiYuj4reIVRAh2bz4pZF33
z0FPpiH6ouo8ImoC737fhlClt+/rMnBCOmY/aA+oEE9UQakL0E56TPX+xkVGpUcV
z58htyLJF20YpHDYY1XgrBBy7rJkkM1yMbS7ISz0B3/OsQ1+Lgspg96Fpm9AZWEA
VBGszKN7DTuht8Jg7hociPft5APLTY7PjCy7Xts/jb3BaF4EjvzIp2e1WDiWdt6N
YHkDvU02K7AK2eTtm6jcgxNa9ODxX73PM9mU89mScIpjmEANkeZwF81SHX7yFstg
VRqldqM7V0Mp5zOXWhAb9iItL5jWzTfmFLoRhxbzqakfExknXrFmtF8LNgWb+M4f
tk1/cm8MfeY6sRQ4HVd8CG1Hop3PtM5XWaHmjoArTp/fyha9TY49H9nT+QaiY4So
CqfCVyQ8PeKQZFJFOcTV/MnLaeysRBZkt2gvuQv7tcewzw0u7UFMorRUX0U8nQqq
wURHXApZuw0SYolQBZH4mGsFRShlbtWaJMclehM9X2yaAcFsy/oo0IaRJegde5F0
KE37UgfFoqf4oOf4s13ZpPQlhIKwAEkLeTe4g21nn57WuY/QSspMfWmb/KdKfqLA
gcEm6DbPhL2dFOdtPMGwGNRbFQ+JxuOkZ9UMeneVnCCsWveMVma+FNc+glJMVJRm
cgwC60MUU1rRpu968nmFazoq9Hlw1sofPncuFRH4z7a4PIOeFmLGbd6QDwGQUb1N
4EKqf+EHvfmUsF4PTjjSpus6Ewnx3SASB3hvjxvyKnb/9h754gC9g5/K1QPzPmNs
iTzKR+848e3cB2lDR3SiqGFND1ZkDVikWq0RG0gqmNl/UgHC8aurM78ssvWYR7dr
Ykq1MnEmLOUYcs0/wYEoZ4Du8VYtjLCrxAhkTd4ZVLorZzdnnsS8VZ+vZqBLs8Jv
GYCHfEx1x2MsZlHyAGrsvXPNXA2WWqY2zHXVgnIbeCTOtsp08xGSv1z6AD3TUJcv
j1i7xJNzmtHViFL6/KwIfdgxywO3ju1zpLebQZivEPHhh/sUyz4IySLfVRGl+8jB
f3vphnWhkjjpyJMRCHwOEwTjFU3PatOg0HcYX6BVgK1RhnKgeXOSpdOv50tAECcv
0ZMAFVIC8QLmlKJ+uvXyFVnH2B9dBBlOKI3Wni0hLtU3EPTTdDY9Z/ioHm1ikIx0
zPPOiB3iagwUOulX4VXGtY2Ow0Vzz0PzmY+nNdTqd3xr+x4vNRWonhHjEaGthd6x
T9C7Y5ew+i9MqR02Hg/J5HW2GuB1JEIlisJ5nDd7UPv8vEBiiCTibky8mhgTe4pV
rL2gdDfTBk5x7kLB4JiTY7ktmZv8tawJl/6SUBgAQ79ce/YHLkbizlUfuMp0UDpv
CJghiWTe3n7SHQe5LwARDJRu9FB8eGMM3FbIuy2e/CxJtKOaDixF0nQRdKiLNQBM
+cGSxdzJ+g/1xlvF7b+zU2QmnFiHlv68TQCL591mxpy1pQQMuzQGYE4XHleu4OTe
9wshl2gKtQ2uc9FOAAl2u3aEr3q3GFl972N1f6AEKHxBABPuPOsCBByTQoTGjMfS
P4L3/OmdpzkSy152v8sUaN2LmvjMJyZuOns6JNBMb4qTz/mGr0eZVqWFTycyE65t
wvIs1UfkB2Cd2/uUgnc2IlbDOYMvJpm3zhAPMPLtohO1Bf4LOpAYBwnP5DR1UJo7
nzivLxxJUF/CypOr+PGQfUUAPiQt4Ajg5KaWD7WenupeZFhxg690B9xnx/sRDhBe
HuEnPO++XAVdIo7qfXBFaaHTLBoKWiDGOKlYv9H79ALSxe8i9H+en/k8/cO2zEam
qrDZxJ7O0EYJk0rEOC6YNYBU/04tGSAUIjTV4gnBOIOzYhOckMwvGGoBQQNO9pyI
kXkGM2S2uH/ijbR0v+uxv2U5dwCaPXVYAvu5dtPsmv17U9KNPNz8u+pWaXA4hS36
tTp57p5jqOCzJHioCmqkGeT7VK5x163Er6Ng5rtccp8ZDWI5HnWPKa7HUiaz2dvv
vdbkiYwbcSxHyn0/uLD2lbte5vkCYQHSArmewnAc4GzQKI5++6UzLBdH1XQI8gnj
F3jJ8Vc9M3YPxXfJ4URzY/aG0F5QKF10wSuZDQpY6fQHNs9ir4L5p+IUwNT9p8V8
Fy8dfhDOqLNDFXrYs+rQAajP8n357v+iidmWRQHKjqceb9MF1g3taAKH57lFFwG+
Dv7iz2/goPxxyHmwPEd9YQ8iI3LaYt9cy0RMatP0JBIv7QwxPnx601Xpxq7fenPR
Imv784xHuERRqv5Zef7fCfgpqPXmD1DfhNZN0uo+CDiWYFEf55TfgilYSF1Fx9Cm
F3HS85wLeBNT31zuqbXRoKngd4o4Uq0R7d1G1mMBvVbCzhP3XJ8KMrsjVVF5NShz
Wh9H0CqW9C19lkJ+2oRRkWhjbZw5zzpUtku33ESUJ0wzR6SAgSwV67VNOEwtGTOs
VDwgz74OtcLjuaxgv/UJ+X6q63ZTiFNzUOJMdYMTYCn7Wwu/C//6U3CVSI5GjsG0
uUkVf9qAPKaz+pY/tTLBhjOJ+bTbfD2Ek0qXq0y9NhdVOEJTJKC91+r+elD4yS1T
mW4fA/Cy6M9eDIQbBPGdErdKpLF725/k3cYimHIr1gz7xiR2RnjUK+GPgjx++Y8L
xwFD+konBlAueNsTtSxPJiFMuYjXmxQIV6kizCMjvpTrWBwn9NTYiYEZ+BYgDqFI
vFQYZHzW0R7SdTTB24rCd5dTAKPUcITmBP+a+Izn3sIvdbZqfxjCdNLX8iEwC679
sj58DHZHMXl3cXSHe1NspU40IFBPH8JbnefJx0FK+VNjeT4u2WfFza90nueyyi16
6afMmhatjJOEf/qsC3z6diIE0712H3q4OsDs/DTpbWH1nL12YWj4X8pR995cG2aT
T1on+K+M/HIwfCAEF51+PHdlbFceA8OvHwb16VLWvvJPfmYpIxkm5DNoHlopP2yt
yRjHQj6ULa/wGLNYhrUT5WvRa+MP/lP2wgNZQgiFQyo1ZWZtXRk61S0BiD5VnN+l
pc8LX+ApE+zsuIEHICO9uTZyMElACpGutC7ytUkUOnf/ZAww38rVJ56yqu0YA3AP
bFH26dv/yAbdZTg1iFL4KFYujbzi+4RvKvVM98hPp2WcDFKDUvGzQuz2XAchR4MP
F/Jdoxp+5/Z6orCjM/0/gHg0ovqa+CfzCwqsY8NkKmhlLzf9M61pOG9SMr6Mb7GX
0Kt15rzWzpyoatxPotmPqNzEYOUB25PZw2dDZ5CFi5zzZOYsdzFAS6EZn8rMnFDC
FuoHvQZWvA5ok+3/R4fbVu138m7IYmSK70O2CnpyZ7lMUa2ZOl9FADpetwm6ahSq
cXruiSNEzwIETlIl469QB0qgqv7G0rZgE9wzIhmddzMW///3EdLmIewoagLjaFLw
5hXFJAb9N/HyKP4GUKYOMv8S0sBW0RjSh9OaaTpoCMqEJlKXin4iIbIarsPNXfk0
XTKrtYaj14G+UefIE7Rf8rRk9wIetFBG2qYSriK5siD8dvo33sEt2Jaqzsut3T6u
vcdqZps3KnGnEqS+wuOEZn/jARyOroJ79Oo9RhK3w5k+ILgrHlQOog8jCnNk/L8o
kIFPOOJgTo63SVxRvW5RxtxXYmLMGHhOmW45HY3f5OSlXCg1AH7jQcJkPWj/gBi8
283BhBKXFRN5Tm0txcHFS4QCkjxI+WPESzJyG+rCxd2zUiIOys30ucI4nYpx207A
BzjRLN7Beij2fmfqLe2ft2AtsNxFSSMJ+R4Ag8ge8M3wnrvYcURL8t0RD6QByNiS
aT8get5+PZrwWURbCCr+YFvSGuYQ8sGhArA9/Q9sur5bbIdgAALdh8VsBYMUOx8i
kD4DI91hUU+HHIdhj5qjojbQaj3cND7jKyni9fuQkcWrIZDEtnNK/sj7YF7ZU+OY
LmrGqbxOHA4FxZA/jWRLUtJV7+rto4RFEVR9VnxxEDoS9URQruPJ3hrEaJR6oPQu
4jHJLUIKxscUPy1Gs4hLgiI2jDSE1zHkAHvD9Etd3poQfICJUVPeTszUT5lo2k8w
nHMNmhfmmDDBrvmAITMozU7hz0TwVHIN3PxNc0JWRcWCik6TDt6WnDq0o4HmjWCQ
gqWdidlByQRPbbjm/kxqzH0mwTYtXgVOIUwrCoPQPx3XGIkYCi7Vk7AHZD4JRRrO
4+x3CSECo86KkesntIRaAx8pnsj+KeiBCsR3UCPyV3nXDaBPVKWgW/+5DKsVqN8e
1gXbyrLXwT/v4EeCfaSFqRmUHeFoiI1ExfQ2OOm81oefBTCKTFnpbIcN9sl0DH+n
32OjJ4mF+THM7FEqVvwEuvaVGRPzHLHDZNZgTrAPn+HFWRDgjbE7iVc8V/FhdGgp
lI9StAD7JAMt8rsj+IG66kNpPDs4i5ViBlJtidijwamCTN22P7WDE/2mja3aeaBh
YDOmAL/UO4Xvhnwsv6wMGzF6WgfNd9jF51hIJn0QqKr7z7oB5M4KQcB/ksSLa/y7
IDbmVg5R1m8xx+XWY/hIC+JUR3eQ1MY+Pie2fR7NRdPteAr9uzCocv2+Pn+1WO7+
ZJdpmTrVhn7vryIwaqIBmWiW6D3499enterLDx0vMb29BJRRoFxkwoKKjjCJwWXK
uqJiSROINP7XZdtkaOY67f3KHJclLPdP1jrxh1TR6JvZG86tXbd1XqUGwy3LugFO
mstdnPXNKqXUwjGdiKVA6IhBLoXIoV64cOio46NIlMxaprNG78Rux3x5MqBIEMeQ
rOBJBKzH1viaQvIc71rRQeDg4G9pEzRm8khbokHvA+hHuwhbwZtAxpRMmlD903JX
snSG6dhyrwIz7W+ECcZFZf3CXA5tHzezMDUewVRa/nAjR5SsAHt9NvXGxsT6ICj1
nNUIhJu9D0SQNFgKRfTu+omjDZRjWLi4uOSEOpL9LIQJz4dqE84btk4b0N0eBU5I
S54MhSn9Q+8FRf8wrwF8HxvJ5avLRMY5+hiuuiI6JV9TK4/7+gXtWLmikfPO9Mwa
Uoq6KgpKweQvJVNRXUNjfSlUoR/oVbFKyBTrKiWk1yLmhFsbLkDJNloQ9lYUgOrx
wZ4OfayUfOjByWyEjsJg267b41UKaIrx6+Z+l01rdPUogpw/I/L7nbwBFNUCQJ0D
j9lEPRpBz6sRBqXJTZ6QOqJ3Isp/FWgZPqWsTwdjiQ4aNI5stHoaa25xvRt/T2jo
reVALj7eBlbMybJ/GMCd99mu4GEhP6Kgs8S4ZGF2fDGCpVbAmlL+SKECzGPQeXEx
VvDTV6P3PQAoJRU3RfvWUo1uWxdlLYQxMxjiXxS4XMaBo3S+7y0Wxf+OqNklxLKi
Zx5BaFlahBXTmCBFMQC0hsO4ncqt9lNZN2aw/p2izZozq1NOeXOcXrnnGSiSq0zs
RtMjj1E361fH+FExGhUTXTuFeHbTz2kLRlaQHn7u0b1lo86ICBuxH5akWV41Qx/O
akh3X1P3I0RiL0BtxNofippk+icdNyHItu441aX641p4bDZ+Qixf0EkuV0pMblj8
cdcd1i78KT56pqI721qB3PapyV/f/KcocQuKX2ll52GcoIx5qlhwlDQY0IxJK8tl
mHK0Ao6Pu2wSk5OiRBL2aZuOCkHIa/DLXnBxr2mghepsoEEMhcAikZ5QS9b7GjSF
IxXekG7s3LkDbvjPtjrou0Bfqp4qIITUn+J9w7Sq2Ef9kP8AFarjF9LKGSDM28FB
o4zfMFEiyOnT8GictRWm3HSPqBaxqyzA+Oa0OIDpQ/KOX8Uadh6bfu3tLkw2ompa
QeyTw6HNKEThiVgxG4zY8L+RklMMWBLv/Rh9h1dV9F0k+iH/HT6f9a+dSpSyn9S6
+i5TJz28qRzIuhZPiS867dqbarl2WcRITXeHBDwGlfohWbUI9XunWkaxXDf5Ato+
SmC2nnyybv7bs0ZS7PquHHWgOO01Qj+ogb/5Tmw/BMPpggw/gpTubbMcEPN73YIb
UT4U8wumHB1uZxPH93gka2yMDF4xLa0zWXXe4W0vbBJo5xJTkZ24WjmCZqO8higj
UgfD8WYOBaCcHYH7Lu+fvbh4Q5/bnZ5PcMrjSkSdQnSiGIYo12rQCsgyKkl58u8E
fPXpP18ogkhEQ0SSR7a/fgfdhnW1leNTTD6KJdGfio7hhtoqvCqeaR3IhJISqO45
6x9Aa8j1x6mpMhpS1jRM28tZrY554+s2q3pVgfilD86M6ozaH8imRIe8OhW84I2w
kC7dlOjKtOAwBP2gPIizdNP+FuVjn/dE59P02SnLx1285wTho9Efm/hm/ZNfVgYT
XXfbEGbLQx0Gfw6bSVeDfinKJrOhPvmNvZAV9GAGyNHqq+IT+iHXYxhi5s6ViWDO
NntywXA9QvVIsMthmU74VEXwEaegVqJTjFqh/JDulZUh4A4gStX4vDdjxCKzQB5R
zEcz/SdKMnm99+db3hU7pdpCRaDalHEOCK+LEwLOa+XSJLSndmdgFBTs/Zys78cr
vXPnwZpsAZZUPvlP8P/NEOQMvljuSSunnd6wE9kKil//bbRTQVepaA8l45jsZ+yf
cOB4Qlzo/k0fD16CWwh4f1nmpR0+fjwuG7jXTEMTU5oY7cgrjDU9uFjEl19CLzky
1rjOP+zZjCfmtTakkQC/a+zHUn06uZ1B0h9bbO8DuJMZPzmt0KkpZS2BddNewKCK
xsnnzfXz/Qqzn6jf4ms5LyJHGAygDPFn0qjE0Rpck56pp9Oj4SL0uPsIO3Zl7drq
j5HTVlFYutMZV78aHWjCwkH8dtp+G8wKP6agImdFHokzDDwToFmx/rp6Z4sA2VfX
0b1VkekMsI/qswTl1aJnLB9b5EN9d+TLI1Dz/wlWxTtD+LM/C+HjSunonrKTJxMD
O0VP9bfq+hkUG8UXSFb7/GDTGgGfUOhtTwZ7gv+6PgWPiHXH8LrYWWFVQH+5Tv+v
XMOv9yUwIoGjHYr3e0max38axp0023yZ2t0vyK+vcg6BN13CP/HKvik4QZIbk04O
B4JorkCg9NIsplnP3m17PPVQ1JM/IMNgBVJWbp269F5iSBUtSUZaSegpE4hTqjvy
u4RXsm5lhvAoz+9fPrDDnbuUJQ//CBMQBSdEd+4VQEG0p+AhcOwilsErGVaswcaS
7aEUQ4I/Rz430wylappSUKw2gYhFKOuZdUTp3OmPDenSn4ubjbNO+KvbY0HMSzxo
vHyhoId6R/QMLy3lgTuHAb7AkCjTs/e4dnh2fpFsTgvltqRBL1wvtrLteI3a3Pve
BVul9fqbd6i8AGYD0qJe7wJ3ycDepeQYnN+ECkB8X2WBT73t+fNSRDq9h1munR1P
NVXIz+uUEqSzXLJI+wWNyACmwvefZptc7Ju4cvTJLkD9Q+trfZQL/j5FqliLNjQR
pscPuB4dsaYTr025VWKT9DJDUmiJDpR9OCK30zf9DbhjjhKi8KnlYiOn04SmwC+9
iNH+INv0oZWhp2+j9EPR/xhof1jW6dn98NYop/QusD8+oRiT92COIvDprwfQQoGp
DYfAMJp996upBFh29JvRWzxlIdvUVU7/xCTmXWUva9+B9UGgFEQDc1TBlsSDXvCP
cxbARcnrEpOmbTUnVQ1lPciXCnj+/JrRzQAyUGjp2JSVDWjgEfqxjSaU5/DhopW7
ce3yTDL3Xqhq4VTeGaoByyGS/ne4U5Tv3KyaKcJmGpVBbRCz8riTb1xlF3tminYG
QM5mjFFt2kJP5eYsvavHZJDmGcWoO2w2od1+kzmme46owHeDMrxI0xLippjVC5WB
ukrve9kvzX33mtM4Xhf/IkCS4T/Bevt08rQj3txgtWb3OvmKwaz4/yCjTRFzGrrJ
yb8DlFa3W8IobsPbn9GgLulXG52hCuef/aj4hm9dkhABw7sQGHTnDPItFJYeguPL
dFVBxgrrqmsDH3K57vfyt4uxbIb5KKNhxTvQB+lRIMSc69X1F0BgHOkMuV7CAQOD
21+V2il4JzzV1sxepNw3b2qI/EKPKHCMhuP2pilxhnxvzNSktzEhkvBxSLcV0jAT
dpkuiYcR6m/GSSAgFq+C11w4UIDD9Ikioxuzzq0xNFMW5qp0dZp0sSLMsYDhefRF
888Bfh+NYieJkqvcFPFWBy4WwHRhoDZonnwvPdo3xSmAZipyPFZ//2MHZkKtR8Ti
a9jWJrVM5nUCOKs9WI8F5RdFsGpnXnMjjibi2BT8CbF96d1ytc3jH5spkza5Kfo+
WSnj8dv9NEFbwaLLomE30OrRirojmYDnxaow8jDyOYXUbb/cm7/Ol+wb8En9TGht
pmvgodAqU8+vyzWZyqC6Q6lbi7FlDL3bNjBpaBZFGNuvyKK6Y2O7twj0rq6KwqQh
UJMRURvWfFq0koIV7tvs4syOOimbLqHM3rLc8q4kYhkHTWl/OPfdNK9lSMt5Tebt
TETfAEgu0xJVNc1izaYCB1J4JE2eRuNGLkfZY6apRvAFaAH2ltngUwoa9KcjBIBN
3eT7K2yvhzJqwIcqp41+NUT5sd1Cn9WvYgqaQWpG10PEm7WQaQPy5URNFabhTM13
ZsSdG3qQMn2PKnq2sl91fN3bZJyrIS/ubGIzKLFAOvdbfUnmKZ96wZpi8v2gdrRu
nyPdJ1PlAtwahLGbNWSVzv+v9y3zaLaB2v8Bzw6N4s5QIBP3Bm+xtgLVEcPpbbfj
RMfxA3gPPNsaHwhVWu6CZ1WXs2j5bJUzMiccZxvCkvPdirhpRk3zzjHx+dnBWx6+
QZrEptKnno19WcFjbfGsPA2jLMZd8hjv8q3pSVROeqgFjIBwJJRyC+PsAJz3n78e
Z9vijpYRKj/ik906jAXZIkJfYkz75vuWFoa6VwEzS9gvKwcAZXKLUdo1ATkxEas6
BYivKZnIs5o8rUciWVB2lYiEr+tfztsPvXmpHT8B7qFdUQv5kMxJJQgBoQaw5ZyZ
C1wlUObzte1VAps4eiwM1y0m9ZhBVupBolxq76rfeTjdBM/yyTEvk3Whr8sr7xPo
uUkXnTGy5u84c6tI4klRhkBnfZzp9lxPnG0CEsl3zQSbnWWefDXiJ0y39x+axYYH
usS+Tkp/YEhZ/SJQt9PVfGfE8a4c5gxAaUVYsNs8EXEyhwBtzV5h/2XcgBexM51c
EjOOOeYVc+BJra4mNBq+gDvWKmblFB4Ie8wpW9T/OabQjZf5PoTuS4Wh0q8CB7Uu
JL1F0H+ukAISRCAvxtR6oEFxf18y5T/zfMUtCXMTLqmrmF2F2O/fUO5gXsygf7Lk
kyK+YGK9sqV+cBGSt/aBjaYyZCk47PCWtbcmS4a3EIkGsImhDUTCgNbBoptfM0eD
emYjkdsOaJr233AHgwgmeq62YVy6pS9/K342mFVX6dW1l7mLfbVxKM0YGZ4T1HTg
udMvjL+DjfEI4mwF2f5IzQ7bXCHLI5BrhLTw8VXPHmI8nm2487t4tV+Mnpr2ZvGd
ZfsrUzaGaE//vSQ0yCuvtaPnPDEAU3zfFvX05CeheLeiXf6sthnU1oD8B8Iv5HVl
PfazcYLoafW3JLgW3UWzIASb8o+1CeuFc8wikCdww7yTmzzisTplDueKb3NGX248
p+fKMI+6QEjbKIQ0hTmJgntVVmTqIuD9qxUd0mWf2q9fhedWoiAxI0kHTux+WjZX
2xmhM2W02GXnhTePgM6h9+ksHiWQbDxvQ3GwP6kzSxzGxBcefqJ61XCYNUjDud2W
Lzk/XVq409aHh2g2DZIy+rgmoAmb2gW0EvG8oTuhhVCIxf93WOjVP/L7geEYlggh
nDrPZvNHH8rsJ7PHlgi/q36Zv9td0gmPEWxttZI6VmppKDg8vyMxamn+Nk7ZECgQ
ehuoP0yTXEyJ35LLBKNq+/eqD5Z5NlKS0Nn3TmTnWMY36GnSIVlxupRGShcmB4x9
KfeEwhStWbCGKqn6oGmWzS520Q9v59HwNoZxN9x/hPhaa78UnJ1gXdiPCzQ9ZlRv
jBx74DvnYXxSlvLDLzFLV1YDTcdB8MEqGUOdQX1zMDGW+Dzi+IXz9COjZqeCG7r2
/a85KDcOxmiu6MkOK4ZgPWc8j5PiqVH2E1IxL7Znd4cvJ8kCZHECVlgZ/Jr8Rm5d
tE9jHW0JgSajWf70CL/q+2zpcUraKm0p0m5Fo+WbJfHY9QkcsiQkECiAv9BnS7fQ
vQGg27dpn5fpBHsJ3CZTkOAZB+1mR0DzdHjhQaj6hZaei8x1QYR33+Z66nZnsUaA
Ewbgm+34x/FPLhwjH9HP8GVv7C6ek2aV5nB1Hx035HxwyWbrK1PLcnmkV5II1cQq
VmTUSPyj8uCsH0kK6+0AfKfjk2SY66paAYG+XPKSZNC7k7Ic0kMupRR62XU3bS76
yvzlFe1kuSphP9CQT1Ct+paye29P8RFNLdZkuObnv0TGioDdgoMOKYRqJ8FK661W
roAsVwVX7cu7rpYqHWTdEokGMD/s9ln4rRjggtbQqdSgFb2RpG/I9lTZtPJswB2f
s2IFlpHzP8mW7kq1tIQbT8h+DbGkSXwr2gXAEFNs3U4KvOuq1sj/qXrbRo7Q+3Vi
Pa7XygoXvCXIFE58Fbly4Zfp7pk0N7x3D6DGRZxx1zUbrVkDAGFlk7m/gBQ8qGkZ
kDKy5GLBjs+fKkUINcxZI8Hy0hp1ePZk/nOMqs7+SygLx9tf2uwvVtf+oUdvmGjz
U5l8jEpvPhMISa83T03UWemhLbdFIVV9iIPaKexBkfOCnpiU8RiXHwZvmB9sVmQz
5SBPE1uGW4UNWKce2TMQbd/A2H2CjTVL5ezGlEe05XddOt7yM/TrZ3rT+GJPjWlq
jnBiGZ8pEIaOVZp4NAn0/0MlFqpf8a3l9jQrl1LE6Gi8Vboi7THOzIRK8gYJfALn
5rogEMFMr1xbKL8uqgAhHsOOmYvvUdDHXDflGnlvb5zwZX+NZ02sv1H1xDREtLIM
ABgKKh8dSmn8IjS8FH8KJ3Rc8WjbBIkNxOanqBsP0QCN7fAa/TK2d85o4Bn8ySDj
Ny5I7p0givWjDh7AHy1ojYZ/aYKf4jopO9PaGIGwtt0tByqUTVwe0bqphcISIbuE
wfZ4RZ2WoD34Nw3MZfMbpziMN2bguOwUmrU2ZZzrCLFZ9rENOaVux0bb4GvA8Yj8
fujodN9p14J7MJ4tymUv7c+0okDSanZqtXxkel3PvAh83v88ZxNwo/lU/vVU7DPl
Mz4ZAxQcF4RFrzA01acR7m23P4VGpPMf5YSBAkaRnuhkdH7e6RvNiKMIlH1UPBqa
XfQQnvFqW5OFqdspuTYsQSqMtZguUjorhJPwi2w6YybimUpby3VaixrULSVnzni7
WLDorBfFZFJi9moMOfrmlGGY57HAKqP5m6s0Z0sVwzerHO+EQe4jxljl0x360X1V
+o87rxhuZ9s4q17erJeiCZJLqgXF6xBH2uNGOxhDyYVWXZgZ8J4TKvyvOOOBYgAj
2SZ5FtKibZy9hpcKOyCljHXIQGa4RuJYbhynL6CA6srURPGFGh84U/liA1cBw75V
G6S8jR8LHNN83Y41lHepmNuO+LE1VQBD9ieJbGq5JGhd7o2myF2WnUEFI/RrdMLN
Z7xNyd68vbcIB/mVhKkzXR77kvJcGGR/oZjdEoQ6j7x/U3UVLevAMCwdc0HR/Bge
p7aJaAcJoeYR/wS2tJnqlLTeO8f6wjnz0wykX6U0z46KyjaUx/kfBCFBAlD4AUqu
Dl/8OaxXrGI0nv19dPfhUDAZO6/KOTaeOd8nWUK7U+qb3qnn60osMY7/wIRB77Ng
rVVbAYSDrdZoinnUl3d0De2kDy196slCAoZCRp+fPWZyw5grMSZd4W6G2VyYcaH9
FKkrHmRh1kbIcFt/jKffNTGU4D9sZk8L7dJrX89u5O1paKNbRCeLt3Kv5mFRT/wP
hqCQFLdRwCqEeCvCxJSY47Ny0pnWAJRdXTdBIJLQaWy43mWPoyJH/yDqdBLR4AoP
bsKR3PAOCQ+OO4wxP5ZvlND/1Rzi+BOYENNufY0pWW5mQT1xaEbO+gKzYC3x7tEL
VjvImyIfNPfkaZUyeToONBkeuf7Zgf+d+J5EQMXLzmiCB1q4nMX6hrEx+e5MdlSs
hZJxyJWeGfgblCVHL593hCEMtycsJq2MPuy80sp5egbFhGwS19XXLvkBo6g4bBKu
EQVPBR3wA9FbyJipiHtUKGSnDmi1FKdBLcaJ71tHuzERmDxr5u4l9ewbIzMolb/m
Fpu3WmatvppXIiDm20OG907hUIVmkkYTvPMl3lttgyidjUpSkljuk4cO6D4Uq+1P
me8TGeLMO/qLomJhexXAaFmhPQ/ik/C50ae/WsQAzPTfrsIDIJoFkb6674GOMjWn
bMxvxClLxRdLeUUlkWIxCOm1Cf9X7S+p/+ThZ0wAGK12nKzkk7h4KQQP98J/Shpq
9iU/l8LNdG+Z5HSxIdRD8QQDg2Eq5iJrusr1vuig07FgIq3+OhCr2Rq6GBxKwEFk
GSxfXxWcZ1SlMrO+MivR0Dj5TKgDZgSMdGZ6pTJ/5LGg5bFUHJz4IfOhBDacZLZd
omvrRvMBHimUS+J4DlVQKWzjnKAFKNzn95Z6KF6rhP32b+4gBcQ8RvWB9TY+JrII
MYJZAWK6cpMcl7dkAArJGTzKNvMh4kbikeDIViEr69pST1vXHUCKpzYEt5yh6aw+
acldQ/k+5fAjIzYnoqW1GOSFMQ0G1PxiXsDVTaaVb1L3q9M/i5o5Eo5PjNWnwqLf
exVuo9H3EVLVYo2uRPWbPPBN2EnIHx6kzutJIjwbR3cIZ9+4sh9xxSzgpi1Tdlz0
IR1RDTEvSCVKtR0oe3b3VYskgYkP6Fzl+/gJcz8vaVoJwtL5mYg3V4Z1EsT+Xqbh
5E6E5rIVR2ISot9zj5ikxeNGFsbfQMe6UDBC5z8uRaoSxydDqmkivtNLll0sw2AQ
UPkorYq25q0MTFDK8GcEikzv6bFqoAROklRpHUzx9pPmbW+2xt3k2pigZvrOvSdm
bm2Kah/CXfNu6rt6uh8oEw9yd+NC27ZAjoWRfIS/KwAcix4ZWKU5w7Cp33KzMhbQ
y58ncl84IFEN1dQKOPfFpcuL8kXZPHtZkGza9VPJtWsj9BtkGXeI5R6+hh8cQze8
3cdey4+AEAZ1dB7EVX6RC7pW5a+YcMt46P6bDL6x8wwW7g9QSydGJt94xe/6o9+Z
2UZpDcMczPaeY455ZoCZkXYUkhlY/2iO9kkP1tkQtIUA5biGReVqpZkAUvLN2Tr2
4AUfXcL3AMTzPMra+H2V60nGojeS+VWNrqGKMxX04XAgl0Bj/i8dijiEHxv18LzE
6u4IFgVLPHIEBySDTRNMGCo3YWY4zWqgDa2E38MgWyGI3We/dYvP6uOXPIcKTcmw
J55eYKH8rs6Mwi6nSDbZOcXdUUbzxvMyD4bLLFBXfJcGrjXD0AzshLvQ1CW3xnoK
Oh7ZW2Hlk1XvaiulQSUr1DA0hiClA1AF2Oxb5U0cNzPHJgu5oRBSoY23cndBztJS
1wbYco2KTWYhX/usJ+id05ty5KgsfeLuqkTE6JswiT2ulnwuKTk42G/ovHKARkJw
nKv/2f/g7QIrS6dAfA6iUaPp+lV7PqzSjQpJ/zifW8o8SymPeKe6ow6lIGwIflvV
KRvuXzs/zJRuhBR7QkChhnhqc0XDp9ow/RGP+CYeKnsL7SScBm3P4RyO4PNTR1/v
ccRDasSozlHK5GQQd1rsq9wD3BZB28p364qpYdSlbCnCl3wzNkQR17EdbNW12EQy
yG2eCIuaGtCc3CXPEjjluj2BQ2e+VhTesSAI+9Ycp3k2LTNBaE628UU8j5iayx5/
E5YM+/F3yyqQzlJSM72Y91Ognwu5YwBo2qzTXM3bIoS22Z9oZ7PNtqSntZH5T61I
+Pt1uA0mo7agbADquWwlk6tn43nbcIzgbLpBK4QwREk7oljHINhnBgLcponOrgiY
jX86JfsPjcQIg/cvoE29FH0eGxqg7tck0G2jgT9QyjHkLAcVBHxXdRV6mejJ4jA0
YzhOIaXp8CyF/AmVxRYbyC3kbmwHZWOBHSMP/E6zWoPHhuLOoUVJH4hJbcYGDd5b
ojT/E0TujSawxN2AhoSFKB6YNqmBxvaRhOdm++yRZmYj23sgLrqidOWklsamu72n
psuz7VhpoO8bwfeFs3S28as6OexWpN6S6ozMLlSK2n2Ee1lKY0wqV0Zsl237R1UD
oqc/dArgFUvS/fQWZrTSfIHrcXaNzJC+QMS7e+hILGuLirMOdKDVTUYtYjqhjSat
aloDwQMx3pmRahCTAkklHp/7SxyisJoP1iXEfosIbKl9Eiu0P5ed4w35QEscyMmL
/6GiIc8/6MWhjVo74M1kIAQRkZjGRqKg++NegJySQwByv3MoyF1NDbDWcfkP9Krz
9kZ0ndXOVN8AI5KqSavicM/QDDAho3+X0DOB68s5zK4CCuZrd9RxyB/2PxPwwvAm
9zz/dhjqqv95ZkwCy3uN6O/hrWUMYfT+KnKqQC3kZJGxnNdJzlzrvdbSBU+yOHVR
WSefG6bAvMyRAbIndYpv9LS1XYivTVfdGMD+qFN2PR/7hz2d7uPT2AxxSfIwOqp3
RBRyVn9O6z3o1rEZCL6q3N9sYFVvBKIDBJf8S2HdLDT9gOV85XwetpC8isvKgCpn
kXSTqUHBHsY/Y5mPzv2klbd83TSnP1MhQq/oO0768lsfCGkts9lPspKbG0XOzbnX
/sfHMkBEuzRd5GX5zs/8R4/9PVsz99XcQ0Hzd4spwWEMTsqNSNW5XRpL7mAqaA+3
+oP80Q6Kh6RByrpBBg6BYjngoV0is0sa+6SRe2iYspB1W3F6Pmbwm8H8T6RqlNTx
smF7KRmcXtdK966mSKlq8yMtl2T/ekGhEoUsoQtknmLcLB3QEi+lE0g+K7P8RiHY
n9JnwI8d61UPbTN2uuexGb7AOhlKzo9H4rr8dTHn68q9nCQedPsluFzhpjIvuSV8
RW5TaMx8kCStTBVldKkgHVEzlzt0dpu2mcwbkvu3NYvDbT8CLLhGiuQkIlBkSTfQ
gAgEAfCOrHSEkhhZLnV8yqA/L8KdTawC8HNLFlsygxf1HdVPgyyocKx/teHUYvKl
cuQgKmGynEMt+9FCCseLjAqwFcuPlr0fONJImKB3mcM8RCkzqMTPKKBD9SiuIRld
5tEn7I78MH7pFkQvIywjoXpMDWDPvt7jos5s/taLoLKcrJ9phdKcgBvy/+0zcr4p
4xwb9VHc5b1qP/3CVcCgY2je/d6hUsrg0lFy89Xsysr+Os5rMtjrl1HY8poDdru+
2QbQnmFfIM+G/meSQFb9DizJll2JnmNPt+sXawgFj/yww7BI4Hha5zSfsHO4fT+p
cSXW8BfLDS3+KPnZZ6B9zA8fXuSoxaJEOrCSVQuzlKf+Dp0+fRWXZOz1al+CBa9D
1trTGFdIuKbfo6/cKTPigDN2zK2FK3Z5KgFJh5IMln2ccH9422eCcEhc5rGctZqH
mpKz8/4Aa6NwwwuLvTrKjgxF28qIxP+gPC31qsJjuj60je/zCSPcTaYHNEvjnK8w
LyIr+WicOTPov9QNctIxxyTSgCikA+IXyLQFnBiSK+K7eyZXR8cEuZKaq47V3t/D
7ySKE9Lldzk0zc5bpY2vhloc237Ea8qPmSo8Z0bLGINXsSjRO23XYnlkvFpOJh2P
wzIXv86imCyXogcwY38RBmAZnsE2jK79DCQteBnbx/dL4fYDSOv5oQ2smRbN3m9L
KOZC341nrzvDaOvTTr9QxSMhZO2MB7D3WQXXGus8QmWwY/PhE9oqwXOHQi9BVZA3
jjGZFVj0WDRg0OElfCdNWMyTpskbjrnAAqi5+pCcQd9X3iq1cnrnJySvzcLdaPUW
y8SJ7g6HbuGfGyEIcvbNRg8qEm9/+qupGjRNsN3LHRlJdxlVtcS2uW1bidF6hm7i
Ymcmjphl0Am12Q+srxUovKdT5cZVdH0fCMi3evs8QjkmyGvfHfMhnJReFkdOXyB6
uF1zqnmfbWH/Ntgcp7RWMTsVQIG65sq7jvkplOwc/rQZnfcnj1p/JYbN83K6dw6Y
VaWhCJAOVL/3S7TjnEv52qSWW6ei4n/yceSmZVqYiigo3odG5O6Acr4PZ+ekTfRI
aOh97geTyRJuu8IvP1Vgs0huTcIixuingDxz5uFffhqgdsF+qckJe+NKwx9JvQaD
rdH24FNKMzXnwX/l4KxgaJzN1kCrVyk+delnyY1IaugYPhjywOp8M8aSzY7qJz9m
MgqGmH7udDNDCSNZNcsn8vNr7jytAC2c6AsCq04ahZg1ZmsY0a1+TxQ1FFbnV+K2
fTo9TADmZu5lG98CB5PzHrzpvfV9Xt73x1EgYWlKoJd2H3ahP7FIQDI97tAeLahC
kTlVPkfxc8IWMb5HmD/s5DJJtZhmz9FviCy/OSN36XDlAhgBUZGi4Rr0fuIk3zb5
rQFUfJANLYCYcjJD3krwjGsB9eVeP66ltCdjED4rb5BgylTwOxUNYMozeuZjPXuG
1PW27XvISE/hC9WvneLVFXaSO0YqNOo9RLgDLJfsTocCv9R7TvCiufxHtiIdL+YZ
ysf0GdfJ/w/NAi62VWk7ani8/WgGcI9ZeR8Bd6nIvqMNTzU+evwtCXNWY6EBi9oK
CT0HsWYj0cNXG7WtRlncSeXg63qO9hH6Ltta81kF+RFC0LQNSlJyHsgSbcVmB5FN
FnQ8nZtyL5FlKZ8GOLTobxHTCyIxCdllM80+QQFJFW0zXISyJQFj0AFS3LzKXa0V
dEW2e0mLoJfaTBp0uzy337ImmHke0ESa4YPXq6EvTY8QUbqkTKZVScZVVdGy4McL
X4dDCKPG9VKeLhEm7VFqo5dVUsJ/5ISfH5nk7PBVKyD0bNMBoKO0Q0Rq/YQQgPbc
GZDCVR7JmUxOkn2CxTiqK+UKqpFGk2TREAWjg3S+tZqk9SyUXM7fgHpOPuZ1gmeA
IxnsM0y8HMg3d4KgZ8svn/EF9PFiqGb6ujhipIfDB6mHl5/N6fl9CB8jUjL9032Q
/XnvjmwOESedx+vyO9xe2y9Q79w/mWSNWUoAwOtWrFRCGA+B6lL5t6Ne12ZiTzsc
wyxg0gZTXB8gZfacE7WNwOEhazQtjDP+cl3ULEN2DZQOegE3Sx7R04h8130x/+y5
n2RvN7xfEk2NXpcnZ1CpbuitAMmCb7Hqw8gnp7Ooq14TuiT/sUe6tkVUpKDHjNly
5Dci4QF5NXjCCw/37zE5RqPp4bwP50yiq8RE1nFTjbH4w0rbiZhjavwr+6CReF9q
ymbDEzAWhvLudmi6FAtvgT0u/bAMNgWMkjjTCYRC7SUJ8DBDHOMLCsWn+8BA6s4P
5h8pDr8szxEGIsID6m7l8lUIJXtqAw8+WYDSPSj1hxl9A/VWwcU2HKqUJ8ybNdDr
TLjkjwXeVfCZ1nWMJ8WqVDJHpdjkwnOB+iUHtzrluqhKaVD+4vUh5D737NCFQrBF
S47nGjXLd6XV12NHCUE61LqF5cAtdylbdKuiGt5fSe/rDVYRecUNX75vVhRUifLJ
FnuYZDVj7pwxGWUCF3JJk0WLbFRyxgcy056cQ/eP7hEvMbSGAzc8Ap/k9EhildjZ
5GEDwhuxQr5elVdnZIZzSt+xaBXuCHUSE7up36KZmSxUGLFsdrv2ZT9Gbevu7Yeh
+xr8aZL4vPJd9GYVDMLyxlLy+R7cb6DaJW4Xy8egVBbxQ91rUAuN9psJf9Hj5HND
CMWHKyqSiBZirxG+IVdi0BeutKNkpPhec3iTT/EwOSLeK1UzkVwJS2L56QMVDhIC
kRytqfyP1rfsZFG8ojjgX8kiGvCFQoJEWXgV7K/6l2zPUNIL09GYGz1CB8lO918H
j641QCKcIoknkVVG6xBNRGO9vgFd+FCHxM/ctf4nA8CQxvOdTXKg+6QgZR4meUWp
Rq3AfLs8Ok+TpZNYaI1NH3jn9ISAIUT36V53ykeHIYb4KCJ1EkmIDgIqNL5PT3Un
Xp//sb76Ht/VOcyOKVC18V6Q026nZoqbnezl5F9/LvcUIIY9RIQGgDsBRk61ddw4
42W0XWlVyfSBV5BmB1pea76WFhhquQgh7TbgnpHASMp4RxwIvCheOuMeQJrd9u2/
2ZnlRQnKOPEWNzaMfG3goHtjQhvey2OcXVatgMrWbozZG7HbhogfmvxznN+jEvVz
hm17WM1hkHYoSP98gnwTQe6FBQLZP0zuDyEhPWolG2tZUvkxzC3gs0fWdLOMT9z2
1CWEVPIiurRH7hPOBil6Rws3Ph6aiix94HUfrXOdjFAYarxjtA/vYUm4JVFuGtc7
QBH1BvQJspMjDr/+1gWIt2ZpWhJrzWgUqyphFBJSUuqkIpRWco0mFJLqJNSYjQr3
tYrH5Ji9OO+Uaw/sjHEj3T/MSpMXFuOfujMXUCO8E5C7RbZyItqhBc5v7N1/qs0d
ejFYpYPACkq5lSyEfPowWii9Wj2issjpTFmDEN5R/vFCWmrJr6pdRdS7rx7VgPtE
/CfOphGXhyC8ACQpEpkVxiM6ic9YBxRTfNqpFz7o3FIiCSHBvvx/Z25eIv+vSjLe
P9E4PEtbWAHBiRIT75WsUFFbTZ8Q0dEeBMvLy3uRB5dF6DYiz1sxQregnDfXN5jQ
ne40iSpu/VY82TmIDYMD192Tt6FDRQzJs9eo/8rWdQSMnV1B12cpWqQnJjsC6qYu
ZPtxD1kbx+kWt3Eel3lL/NZPI3w9zY9cex/D0Vnt1ovna5DBGnpoouNzW8RLp9SB
fFxHL1AV9JG99OJLuS9NB4JhzqR2XA620u4HHV7A1mVmLzJp36yYZDdteOamYdzJ
G/h4F8233/uvQatQ5b7RlvgEgOufslcTOVJ/sFHIL7vJae7opUy/J6chTVyO58b+
DWULO191NAZU1hugvdegkzcpMRnv/7Kn6nve5A7YGVpKb0LwAI0ryvJJIqBthAZ+
nvGuCU5uqD6qzLBqdSjGvHayo9/O2/h544+Ooct0kQGPddSKXnd0zqIk5jfkna2K
s3nKjfTKYpHR/aeK8SdJZctcIxFZgGTVLBV+llQQB+zSaaQlrJQUI99vawzFDeQ8
ZzuGaiNquaeqcVjYSpEzDllJFvnAc6XILg9iC1eyYcEEoRfN3RY+IQW8lNakb697
An/Ll5KPIWMKZuAtm1DfipWtYU16RmNTM3Crh1sLVVdPi3roFta7DvWQ1I5Qe76J
g66FYT8v0jCnammoy69bgVblxcbMW9HX3c/MARrRWrKWgt5oPo0L+hr0k8iF9xs3
GAA1wl3ADH+mmiRfaOEcF2v488RbotuejCInoRpi1YWvqcb94O2JahbVKEU8oZU8
wlaIwhrqPPNnyOHZBRrFFLOzyebqzzivqflWa/zNoYpKEZXxsJxtnBhaf7n/BVUE
aJh56bWBJ6l1R3jinJmxfyeJ/u1Tm2sx9YDj/84rqWWedXZEc73uaf49CX0QqHjc
tNWUnMv2xr+KmckuIgpvyprpwP64S2uIxjuATzJL6Ru23NN1hZMoOO81+enmvxha
owHg8/tNLxjM2figSJElZDrVUw8dlbm/e7lgWcaAfemniNUsg5WKPc/WmL4dgqgU
lAXkBMSczjrKQuaccCv8J3xLX4USN/6qsJmiPC+4mJIlE0YHMpW0tp1iZZ8ThRcj
uBXLOyNGGP/rCLBgX7sQwnUrko1V95mmMRHlowDsX1yneGHmO8HoQJrVRICZR9hU
sq6yKUmzJUQVBV4MDrl71+8yCQsMGPQxmKuAkv88t2UAY9w/sKa7nNfd+Qkv6XUw
RAtLOR3N8QBc4qKdRibJq3MZoW7eZ8x6EEqwi293DFiNXl8S4zSkjVXoIhJjrwZJ
u6AGtVLDBBIZdRpnrmpsjNUfaEgE5fqTh+emYSacWqaCBdoE2+fZfr8Z1f5hL4RS
uHde9FqewFTh1SZeHEgi82jCsfJU57twbhG0YRey3hLi1OKE/VrZoprqkJpA8N3r
Bq1VimAqxZYM7bzFCVB34JsQFa89b+URgU5mSFQhYLtqQ9QOBhh+OmYFua2VjjqT
UrwuWwieBBQxuH1mlDMJUHhynDd2MCH4z0CcOuquMlTcJaPLOccI9PbXC71f6HF1
NmCJNaA2JinUFZZloTG/5D2qkKtJcsjpho6R4dvcWFVx8ryIZTkTk3CsTzzz5Q91
iqyLrHN4O8sKZDZL8lgzVN4+D1oHpwXQ42UGGRpcqBafLH9hlT3Gk5P1hYvzNg8k
WN7PRiKs9jj7bVvBmGT2pHQIEqEI6QP0RwWtBQMEESjlW6sQ8KljJXFGh+AzJCkq
X/dDzY9CRmzrlEoef73Ulb6HQ1VQDMMOAnt97XTePIaF6RDrdU5dr3PomCZFc5rf
xIK8m7y3cWCZv052Dw5ofXa4kEMyGTavMt5wmbg8Q2fOgaut4ojj6zxsQvmy/U9H
Lw/BCPevSV8Y4G9z2HmJLr5OpKuLVwgAoznIRgtFrQXqluEzbZ651vw680mFmcsr
5RSWbU1HKIPvpDBvXWjIPhFg8yyvjepirar9qSwz5YWT3QR/hKFBaeDH4vVBLnz/
duW00nE0RXFdtu+yy6suBks/c0SaV7D5cnqdDYyp5Of5uFpqNt6LeCPRi0T0ZujZ
tObZW4RX6mwpiX9Gl6hX+fOqngGUXE9h7m+FfChPx3U5Mzjma3QjmAuffbB+mzWm
fJ1BEV2MKmb/1cNE+0iokpgP1ta5vTofBnFlGaodupmb9sLImY6UR+WXf7CMZWJb
5HZ6bVJWn49R/FLbvSZ/9VzURXWZLVEM9WIZ3w1vEDYioQj8VxBveG/CBwHN5ElF
EXPuT1QXnHeIXJhnPC9oN9DIP4STycNTN/gE2E7ZljXHZBDkTb5onfs2/3rFbKO2
wQS1/UBw0FfCqgGck0PsEVIaDCFP9ckyg978/PTz0BI+s4D4JZABl/MFKeUqIVim
+iCboqQR8APNWJMaJv0GN4nk9coPhbSbluoK2HIAXRt7hMHOmlyTJxBHuAHRaChc
TWsRTieVRTO1QI7l6S99C0IMDKzfJbj+qkOxpQYXN4RqFfaVQG/few972OOk641e
wMRKe2Owzr12D5yC++wXMIQ68aRFfgkpv/QwYved4qssm81gX6kd2XO5D128Myg3
BNR64CjCdFqO8gsWNYQSQ0DFrviK07/B+xJCmuhWZCFx4uJViSvzRZF2eB/sP2N6
M1ESy52LZainc1K9lqKIPSfBdOoREjGGokSA8gGnVY8KH3NeigAxDHoYWzhqR7CZ
O/CimujM4LqiznAl64zaHc3N/LSszfHtLxp00HR/aNnc/c6zieuTwb9hmvFtxsIf
alQh+0KCqUyeHLlW3fipo6RKLrEkMaxVLSkxON0m1W0MTJ/hv5Y6k8WFPElA8cN8
QQoxMujTaInEjg9Nc45oo6yfPmY3lVOSV3TRC+H2Mvyt9GQ90VPz7KRCRm5MsF0X
yvKeeKfAdgMVhZ8wSwOQo1iL44c1BfZbzmcjo58xVILGXO+iHjaYcSQArvUQTTHG
lnnOnOQRd6sKvnszXikTS0WGM2rYQw1AerRg1DXywjgrBqfFWiN/9G8HGxUKbCD8
8f7Ge4zptnmlWqdjvW+6n5zIc4wsHgC41DsTVZSmsX1BFFyJ5sMtEJXXdQ83zOBD
Gqp3/Yz58afyEYyBmHcydbSj2xCJ+q4zluhL738gHI/y5zRUCHAGOKyRLjJ+sLiU
vfbbK11ha27nPkK/2qpQM6IbQt072/O+YKObwFWEytGPq7lm1Q3fq+35JnpD0g86
rLMpru+ItGC6AEzaJi5jK+WTn88rMaBulQbmjUuMdF1o0FbalKjchP+IxVWITy/C
O8fbB/vd4AAj9gScDuwowN/vkbf6vpSsAdbKAYc6pWWzBDkw9npfcQNycKk7TzFO
Yl17w1T50T4CIAtSxKRrp3pb5L6QOdL+9b7V6+lR2Pk0/ZblfUZ0vd6ZMrsgds8z
ONTuA4F0kxc/p4AOc+AFY/uy3BKrtEHQIM2QHM/vmOO6eiU8m/7MZ+dC0Aag10bP
E+T9AvQLGybsCIA91jA2alw1Khp0mEBQJS7wfJYd1GC/+WyBCq1i+QYI5Pz1TuoR
8+q5d2k0jzIl3xRtNFuk08hW2mg5tbkWRLdYt4gVy6bXyvUkj0Q9ai5siO/GU5zx
yqwP32Y51DysrQhJ+abuisJQzrqDd1SoaKU5AMlOXZDHYt8V3Vl2G64ByG4dJVxK
YF0HPt9AN23EXsupeOh27R3Pq6/VP2BZsslSesWulrDV53qiqQzN3x2On8yfcrGK
wbzSFfHXCfe+D6BiSSnctOT7HNl8NOYl3NT/5HPsbfS8DTQqOiwxcPsmlxNQXI9z
AG2bzhz7Me3EJf/flUp27IsUIXEC2DhcpTH2he4MR9ZR89I7Xnna6RxbrrYPxABv
t6/6QeCtUSEgZi76PXcLERQc4sUSSnEKLORIz5BxLcoX4y935JGquyofBVQxtP/P
1ypWya2ZMTcC4UEW+IN6OTbAYrHrB1HD3H+ouZSpkYnfwsUoIxUNEJHlcx2CQu4X
BPZ0e2sxW+vsOc5rGy4D54ICQnwXi0MfD7/gk/f1Glo/GChJN69aYAD6TGnj/r1a
bIWGFAJ9lEeoOhCpyy93zca9CU/vIEFAC0zW8eBqm7UqRzdDAqY8DLNu5gFkFDCz
GKRUk2Y4CKEvq1ADdqt+7BMmkQaEBNIeOyPbbvGM5OMlJaO0FTKI4ZBiAdILxfBt
bCR3CWcgVawfzod3wR/eOR2EVNDFDht4yRCaUHW+O4qnVe2QF5J7nw3X85j3Vfqf
h0FjD06wGyZ1uwAxn1rqJVlb6ec+gLvTQcvH8cbVu/+GXy5Go/aFWbNhE5rP21HY
ncogqqaNU9/l9EHTaWztL09RQbN6SnSJJrlkUrEHskjswIIS8F+uSG2OpaIv5GEj
AQHDUHYmugTLxUtWUOAAnzqF6F5rrik/hgjlMd0WEVieRKFg1UcJpUQP/svfFsQb
wlQH5zMeRtBF5bNrzQftjkW1Y8QQPOjRujXCjPcOlK4yhu9lbCBB+ZfpDdFNzi96
tlmusUUvog05C3fyqXDxcLF1Xxg4qVjKaAjm8/TuAEn9uEjYjQx8f86GyhpTquvs
bUxHZRcMOjLvbKctWPYvG7mRyU3nr1Y3LkJQ5WRCyOW5McdE7yWx1vDx6F4CumOq
nF6NwVx6zA3pFWlkncblGk10zTyPKGJC9xDqyeGq8VktLKsf1agaI0WUcA9p9yqA
BG2SmUDHYNelLr1B3E1o2VbkTaYKdJvO/WhAx61G52CST4YGZx5WZTJfHfC1zw6t
RSuZYPg9xniG/OJUQ4m7Z2qbnN4v66w8G/OnzVntSWm6MGxLbv3ifJ9Zv/gNJWsl
NOncumcWuDm8+ilgxjurJbKdBE2PhQNr/S6JEN2LwrgXDdsJ/KO7FeEmieiUkrmI
eZu7LoYNnWHE1Henx/LPGiCK881yljJr2QGtOzKSfIIcPaQQtXFE76GFcOKy0OyR
q5y7+hztwO1WnJD+BCG1UDioPqNBhqrUrfl24c7wWWz3J0Hs4Q5ZTq5sJ9ChYhUG
zp5PLEdgLciDG5xCC2HwUhtSzn1RaVPZkZZi+cZnxo3Bvo3NT1tjJCqc7jmqaANm
4iw5lY8LeFYr/jO7IcBpAbgPd1EKHTTYTm3AX+BzXcYzm9j+r32TQs428Jb+eNyZ
DRvYLkM3x+7+VvVsfoBGMWccfPN75tPUvb0gbRXvofBRLoQOT3F5LHSBciWkDESx
flEKjdkrRJv5uQd/r4yGRVbMamlZzalBI+BcTGkng3DP8Bx44uuFqEEJxRMJ+UtI
UEzRQmUlARm/wSKfPU9IoOXEDkcvE0OEIkRyOLdLqAzjNc104X6ngrBtYXpJoNML
z2YXNtjsImYHsGD4ArtBluCIDdLOZKscSKi0mU6iYei8JGZAfqQZr74hq5bAUS/o
/I3LQ/Vq/haXgbZSQux1O+FKmPy1ZhVOlYhbxtGkFRYdet+42R/1S66mv5fdnwSu
+yWFgjwiShzo3T3MISiqEFystSqHfHDh930Nv8prpE+9XoWecvY4baok5eLP5y9H
q2qj6oL5oBRc1Fsi8rvDzNH3++DtDcc5TCOxVmmPJzdT19olDizL5UySdXpRaDTA
xcl+HvoHviqH/dY5KQmrkfAn5ZnGMBz+sLMwqucB0kzgRYH2/6kYU7ed5BTuqrd9
qJglOpEOzHaKepOG+jrQZnKadU41o6o+eX5VtcOELdSrHOiyF4J0syXYG7hWjG/H
O9hlYgz1p/ovOHcZefinifeHSGxErwCuVLMbNIex6t7LmsuuB52O5Dk6Wa3oe0Yc
8/CiPgvUiK5R5MG0csthqMIrsKLroEbeugforRTEph4bjqdNL9pKUYq3zZrACjHl
0ijEaHqldq2uU4KpCh6Z5BdS46i95ENEBJnHepeceW2ELQkapbjUdNGD8PpclxuE
zRC9vQswS+iQ00f3uzcgApL4U7BGbcJaa7sI1QpOn2uRY4bZkbOczLhTrBMNtLXt
bQfbJb20KVkzR9T2VsIeuhU7tJFOd2ZDsb5gkx2XqFDi0WaegHPrPZjzyuDBycoZ
wUNzgbhXPfEJJyTspaofyFVp/XgtHoObShDnPwk/mI7o5vvHlF3YfSEp2LTWZEvZ
k9lme5dxze7lU2mOBp23U8Ri2Di1ljuqiInDM9D603oUMY6gqQoqQPd42dUwPWPY
Lh7qxR1GvtNSij4D1esvdua8MC4qe6GlN0ee3r9Ixjtuujvk3mtJtsiFkDwIYnuj
CKGMmwXE0hnEy/sWgd6jXGtlQtzv+wuRPSyDy4QyFggwIrmD+CQmMrRbfOiV/0mv
bM7y3aSi4SrRo/sM4yG3a0hP7YCvX1a4JVQIEvj7tfkJn9hMR2lITWtuS34P+8gC
1P0L0i1WfcvozzeEB/j5l/ry+bZVLZ1By7RIURjB7ZuRFDt9VNMWZf69QAU9lhhp
cP0oGtLvnuPnN7I1/MV2dQ6qZ409zR9H5/qF9sFYZb0f6cXXwjGegJXYipSAwhic
dK4RH4Ab9dp8Wq1ojtasasM8wqM4QXa7PpVV3jJ0hK9fBWr9k+0enzdoIW/6BylX
ICcLBsIv1VD6E+wb0DqoYSeYIipv7V314Z8KfTuLpUcBbLQMvr98PHVPWQZe+I+p
swFTsHbNozFiXF/0eqlrlE4MzT+zk2R5WoIJF+/6/+XIIhtnPnAd8+5Ii3RBkZgQ
TWijRxKQi8LmJICBUuYTm0CRC09kjqlCZ+2VjbAYOIBWCKSooGxGabbijog8NpCL
OL+qc3vXX9KJaNqny7SHXg3TvmqwjgRsa712e2dQg8R9yqAghUSEighEXRCdl1p9
3y4ENqxypc9QImrPHFIXhncazS+3OPzqraNpDBG1130NQtRY8Zx3OuMNx5/0rsf4
09jeAQtdFnSjFgqj7UHoUxHB2vvDjG7Z0abwEAdW7/+5I3SN116SsT7TmSTII9mN
v6NBVlLCJAW0YlMhn8zPIBB9IHcj8jc36caZ486Kz/ZhCT4TWMhpE1FaB4R4Km62
QLFeNNGey8HcTm2QFZhEBqZ9HYF1rLswT8Y84hAav5LUlKxUj2Df9C3j+vSOz+wy
CPbzICeFzAscPYtNrxcK/U661Pao2vHhGmPhwZCm83bmQZU6M6/TYl+AZM8bQjry
iki4bwq2gGtHndNpkPpAqXFhfAX+M5+bottHFyg1jxDzR7N/iZMI7GCJMJQosblM
Eig1wbSfbmhkI/26QlmWojUEVnXkQ1vRnhRH0DwxcWzU/O317PiOS+9l3DYbgq3g
BfFNqsqZtjTgRl61iDpYbfH86FbyU4DZUGlxs7pxHImmaorc+DFTCcLMWM1GurT9
QbCmAOoig7a81fo8W1t96Jt6+IAOvo3tNC/0yMWjpB6Sl/6qtRZBfcF1GpX54odl
23kt1hUYyKMfgydeLL6MPhrlqvHpZx6XoO8I6Ope1Ijn0DFRyprdaVUitxIG6tZv
UkrOc3G/STYQP69QIhbV0Rpt68RN0BLkB1UuXm+wDoxQQBc54n4maB9R8ECrUiEO
v/MzHYq72MUTFi7nNyETlG4DBczY6MNOsR06fnghaBgqnGMBEsiKc6C6PiG/Ibrl
xvyPQ/WwKZrR4kRr2NZKNHIdekAmp+cM/u0MHncww0embXgUtcDSNODkrmRfXZcL
U5HWCp5RwLXIRacO1sHR6Kw8Bnhl620CvOVEgDqVxjPjKcahNYt4uEi0FG8imtKs
urVh3Z/AJZRcKlrBHhGIPkt05ArqbjzqBK6bZO7oLd3E18s99D81FOOlSO8quHgz
0B71b2Xoip0mZB1mzbFOl+IS844qwz1hXF2jymTaksuNFHS8V1z2OYYXu9mtItFT
SsH7GaX1fja4iFwfbUPnPY9jzLHQp1+VbD12AmqZE6vlZSoNPhmEP6F1cFRVdVkD
r9fZW/Vqz9flA5H4SjJIgx3ByRtAhtpByxzYaw9vlqEUNGZN1VcF9RyJo7oVHJpz
3llfPq3l2xj5tOFMW0rNwo0jnD4kVjrUnggIuZPDrTxy73iLshGWTyf6gGJ8sL9l
IpuurKb6XswcqZoIGHoPUEAbgtvScdQBk1t+j4K+0Brr7wujDCFjBIvHGX9k2BL6
p8M0RieKRzLs2mhyOqxVQl9DYcQjxomPMyVI5PyDDT/CXRhXQIttyMdezog1pSlZ
tZaO7YnmMTF0kVjApUwPvV7EJMotuMY8i1bsKh0zkX2LrwFbwWG37gaCevHtdTMK
q1fWhIejNJvIZRZI8p9A1vWa0anVaFlkTNylNnUlKv8sC9EszdlDwapcj5tEuZ52
Zug7eiBLBhyLNoZFquFhC/sgZoDJC9GqhHfRTRdjt2QJS6gohcdg8lYfYWdwv8mO
PZpjefbc65aa5fTqfso+ztwPRc3TB38WFglBxatHkrbackrOzGo+nv3Mlsk1fzlk
AyGPeoICYIOpDtUvrlZZnGYXF61eeS9vtrLUjr+8GCF3En9WMHtvbqth8L0QldbG
55jfGq1Z8SicRmue91fue0/maGflbAp8REYgHtkP8Ur4dJ8dTNq+LlXvYuHDihsC
fUfR6dBfVp65YPNgP9t6xo0+Q6aD3BV6IiQ5qWnJSRB4fwP3zWNEf2x1AFNxvZQa
Ni3gpO54Vikoe/1+vf8MvpTh0Z8of/BpIWve/w068/XRwQRMWtPYf0QY0c/twOus
EXH/PA0dVy2ZUkHMNlPySQrtA052WxeN+NotwWBXOz+C53Btz4LbLeB/lWyT3cHv
bA1o+u6NK1qyVx+KnlHGPFNwde12a/aBYCreRWc0/BNWm+EMWHafvYEX3mqESJwj
eqs9F+mjkzy3jkE1p+coh2efMrV6Vdo6/AYYto+WaMcyT2l5MTeyx5yYKBCO60aw
lJHv5SL+o43GysowB3ulc/VuZEgKRhvqPcZn0d68ItjXEekA2tkZsQNkdMDR1Pjt
kYpE1BE2HHz+a7lUzth+wHfiA8m/kn1XgtRjpulvEvMsP/jn82Ct2R/n296oMpNb
ylcxbZTm2F4toiBz+POvfPLXQyMQe4VjgglR54zjmJJYNrCfnB581B7VXPMr/BxF
HgXIJf9Xf5oH71PGqqgbNEOYwbIvmw8UF5VKhA5A1lukcx4YF0pfwfhRnOdhHlE/
j1JgbHBec7bkD1YXaSyXJRTuTUhkJ0g7XGlUq2P/aHpQvcUXxy/miy/238Wkl7g/
SniuNWx6Hzsv9G+9Ud0zU8j3ktexZk+O7RvK4CQW4Hnr7gsfA11XAm6OpVyiCNJj
DZFhoQ33nLECmiLqPQaj9731QVN9sEt25LXPrGsg3ss0M4GFtEdWsYOY+5ZuBRrn
WsANfI9aTaMtbiPDuJtDpKyd6kiYECINq6tZru4KWcFv+x3825qHG01Sza7CJoAy
veeMA4IWKbEbCCKd6+NbBQicq5IM1Gz1n1xY9TVrJR3+kIHoekinNmqlI2y14QvC
plL66Xydy9zlCszb24VU1Rgm99QEE44ILfxQrmCAWirKc4m2LL9J4rXP9gyi52+d
v6poCmhI942I0CYW0niU81F7qoMMF6kV33bA5czvV++lDEk2uADURMs1ay8YVxa9
MQxjkvypg0tMkcVU5OqdmkBYj1L2Dlv+uX8r78ATn7cDHoulUQumZm+z8LGl4UJX
O6fo2BGIlfmTmDUZ6F7iE1Lug+69QMxbZvVkZiukuef/xKF+YMCzgL7dMcIPa4Nu
dbQjxii2fQwi7/NWGT4ZUJQaHwKcVnGRwaiTKdUgaV1HVEMjs0TUmmWDfzDhl85m
2mMU9/4rbZxkoy5dYWm/sh1bwzO7+MNhydD/jI4/UUVTdO21tPDdyAsfHe72CMJB
UIbyjynftwUt9TSMzPNu8psjsO6xTxRCO5yTELNhDM9caW7H1DPYD8WC2YYgpxUL
ovdG2oaMQtCJ7JDW0ofuJjRRTD6UCxPMeJF6XlgS/yG1codQRkWxwzQyZSGToNdB
evldB9gPDYOOKsbQMtUEE2gwqPyopFgNpk/zbJi9fThw32JZVULza8LzT5gWEgs7
bn5OtqSfTJ0RLVBgGjt4vU3SpCdzTjHdnWZN7Zk3a3gI3V9BIypqQ7yhBVlapev8
RogBipopBxKoGaLamiM/jcQur9DlzIQHTWiaflhL5qVDWURrpPgw6QKSSEuRc3iC
DcDSj1geG4VKnL2nyU0x17SJ0RPiQIgLr8f9vXpTfVvCKLN/Pyq5OB9YT20uTKB+
QwLjAyZn7yt8ee/dQUi2N7lK6isNgiFlWTDcnVpM4esUv2tV3oeD799sCAuBgzVD
vYoq4opul2WAX1PRayyOCDH/W/hRRm6E86FmjMY5hBVDirxmxOynaeD9hjhc/HWA
CzDuWDQLdzAnlk/tpLsiraM+10S23Ufcz1ozJPgfPerEGyxqtI7ktJosn1jD1Nm+
w4ocfLM7+G6minzxd2to2qzbod/QuvOtIvyg936zJDpymCp4p+aTfrYO3vAkt2Cy
ORAOdR6yzS6uZ5w2/WD0bou/2EuoG0srYLyHvsiimLNo2555r70ElIIvZmeAIOCn
rAYbUP9jtufhe6HVR07ZFW1Mwvt4CppYVXwb0dUccMnC7oH6ssLX40YSWmJM5Cqd
Eg/uKdJsE894z4HrirHg0FjSPBHQWF3HLuGFiaHrzrlBsY95uPrFzzwjguBJfdkY
twuZs0i1KH/gig91EagGB+HR+mXlM6SKFaWMzsf7eYkAYLnMPz0FE2LWOH/bNAkD
Jm76ic7J2GMVp1UE80gJJMm/FUFbCDLIRqxgVoOXP0YotngVYoXKGwmQQv/slxgs
IvGZy47f2kdFJ6QY+pu5912MVu5DDyncQF3BMjBLHMxAh/tS1SD4QWgZd56oyIMZ
Mtg/7X5Hi1G4IoCK6kgBJ8ZHy783v19SSU8oNrv3TMM+tknTmFC5R0M8toYgOvNp
JkehSRyp7k5j8bBf9J+APeM27ddrTKc64jgJjIzNUM9ACilKjjeBXITZlvauDufW
adHIDHGbTFvAtRucEwRwZI0vcRD4gnFrcyikloARwoKGzxGKcLvn9278q3hZoYIm
AMzPJmSsyE4+5ogVlxxw0qYNrGKWxJG6YnNuC2CJ0jkIHpEkhGxa4p8mpAPb+FSB
hQMIwbVUqbnh5bYvjV03C4ernoFEBBw9WDxVOWPllhmSLko0SCoep7qrYflph8VI
ONf3tOXSpP7LjlpcWxaQduvhaqOKnckdCUsZAGNfFGVFJlSRLeCloZhya731N+5d
KvxJ8t29kwJKhzZW3iwIYUtEoyfGRoxwxM3fC6FprvJolyBpwKeVAVUbQzwrGZ+W
OBqUq2veHBOawSyDPHKlaG420BPCXW65IFC6BXBkdRaQgpH0EpKQWRWY2+MS5gn9
brJ433ujfZSqzXADf3oQYxvkIRnFCjX1vvZUNDsuWXjTiHSkwS+BqaXZ1muOu4vu
gWDmYdDxNjOfh/dXBFyry9Nus0nn7iDEdsyfzjpcWQLsByifavXV1J1eXteomiyf
b3wz9y1QAC2C+N69DpAlVIkWfI4P7wHCjZNsrvbm4ssVckzDCUwpb3KhBaaIgxXf
cUVZAT8wnDFosUviztvnxqwQHBSYidXwaDwNib8AeylrwPY+TCDWh91JSPXu3is5
vfG2EFxY4oWcrfi7XcYdeoZdShYIEZjgkOhjiQhpcF7CoAwdYYKJKmoyy3AW1/jX
khWo2VgQb5eUQ3DUYtVKXbex7csUbVM9WhNDEwH16sj1GxBMADL5P1tUninZmCs1
ZK4XOLylF8XxcwUh1ioV4Cb02vTXFRVyHVfjaMVZ37Ba3vm7Xcww+pPDyG+n/UjS
B5BceYha5/vzvhig7kpBwxMB3jeyuOFwLROe2G2WVjLpUBduKbS3qdjXyvTU2XXL
5kq1gudeJeelXF2wtIzRmPc7YgJRDvS6VKWICpkl/p04w3D2YAAwqScwewyl7kfP
nx/ZGLcV8YIgdD481mHnWyKdyzn14/DwR4yPEZ3LWAuUJ+0tSHMh1Nmd/oHnIh3k
WAzQOhSeOAHab4ViYpprsL8F69SEMko06MC3ZXmO4bYzRnzijk/rVzm2XmFtd1tr
gRJ2aV0XnLn059MkROVqbJqxuOM/mfuqzVbw6xd1M9II7HNXTmhDeFvK+osgwB+R
oGOkBH6E73goyfJ/K40qanWtblYrnzT4FB3lW8dlLGTmDj2Wz1gFpFaC2P3+z+eZ
RK93VoF1agFwqrJKP+oYaHL/EdhLgfzwESWv/qHi3rOO5bvNATo6cyVJo0K94lZr
VejazarkN6HUMNIBfhf5/PSkpNKThWiXR91zIR8dpYYDj2th4V6cSRfsgOUgPW5K
Zqj6evvQd390hGIIQb6M01A2V9R+Sy50xVf93Rn70JFEP0Hsr8ISE8Kzresxgfu/
wtInlDerkhoMzbhENtWpuC+F5Ld5IQBiLYZaYFUtPQ+gcfmy0rAHKcmveGJO44WL
gxvF8UEUq9IogiVxNZfUjFnsSgQ8iF4TiuDa8W9YS1jVMbpS+O9dI5H780LtYvBN
e08NnZqOTkwCpVTydY/0Q/3vVEjZIv8izshR8Se2PgqnlV5E4naIYPKLWSlMYgEo
50mEdSbTeLJIIwOc6c+WifJFh7Ds4lAOqzKMr8jCBwWeCk+b2pxynuOvfDArtKIa
P01K6qQLhesGZfG/iN59yLIDE8DMGuR0CfpVpXf6i6EP9Wkh4pTJfgmMIo700Nu2
`protect END_PROTECTED
