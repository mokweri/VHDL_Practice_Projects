`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DG642V/83qeMI1wols8Jijn27/lzku+ZZVcfZcAI2fsWVNga81DRxQRCwUWnTJyY
gZ/LVieOnasRVyQBMGF4fHse0LZ0UzPc8zHBuSa9OBwq9dO620k8IxLcvIF7+Yct
pk+S23p/muAFMfQ14z3eOQXrFhXjKTZfscbAgMGhziEgCJs0vVF9FnQwZSQY8Yyl
gCQR6RtsSgstdzOt3TsuglXYJ2tXfCB5iBNPjJuu7WnwTQYMKfliRiOyf+LPTR7o
vexE/DAgytnJgWu0aE4B1cMs5h/COIxUraLZMfmnLiodM0dqaiU4LbZVyEVQxlqb
dcDEYDAAlx5w5Ck//ZJD9q/OM97XCgoePptUbcbKA0L7bxcdJWszauPwcHUKByc5
31S07YWWoWIib+s3XXhkBthP3pHr1XYmUEl/p4j2fiE43tw8ICKrUxZ2uAXNEDa6
`protect END_PROTECTED
