`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lV7np9RyNoaau8i7KwlWUqWjcoQrtYVrE5GlXk+wq7cmmpq9jTNWoK+T16k6Vyvs
7UcoSH3vHMeb9PV6HQqAt6qGoFI1NaVYQK6wENUIjTPaPGiIuuzqyS9S4laToNJ9
HgF12zHL8v6Tr3/AvBRf7mTRH+5qcsQE5ZJVIH1SRz4/zY/jNY1LhhO74a9Bwhe9
HNdlgAFQcO3Q8nsm0aQpVqUksFvJ4QSX0Q7BrhpY6gDF87ccYduBbg0R2x3OKhbK
nrnR975IQSFPJFVC76a/Q8NEsijbC1qYXgSFsgjrXuGPadRzy2pqNGsBR6g5TqsD
r0Rkrpwtt/qzlkuIWQBMRVIjFowX6cFz8QKm1dIP93AvSh4xSqx6QSFu7TDvVn46
HUOmnwKd3j8v7q0YXy3PdNOx/BW2Z4lEsSkPRdw068CFHoxfighXf+R0JesvIUou
Dxuia6XXM+RnwJ3+yQwS6HopwropzFo5idsWXeGU5GM=
`protect END_PROTECTED
