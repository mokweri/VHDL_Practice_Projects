`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VL1ZXE89M55DC41ljhZwn43aP49IR68J+troUaeoQO3IPylnVQ26P3wLpOgktrO
Wo1VOuznZSIExopjw6+RRDWvDmm5ks+jb4WJniUJijmq1zYEKyQwuHX1cMPHyeW2
bN3JuwMX+PWeYFNcg7oGObE/Qwjfs6W2Xtqz9c192k19NHQYRoDQzuzOVGNv3Sil
WOB4YrD0jm/ewO1dOfmPmZO9OPoLV9H08WPtZXYv2t3nW7v69uGnyhF4qgSOJTv8
X7NpoPBrMXsddPXZyWfD2BtR25PUdUpmE+/DCYmpRv11w0AcXAo9aqphh3pMAzRg
ZV0iE85O5wWPPTP80qPIizhxR8FgnIegvmWp8a44W2UxmiX1l9IorrnHmhvCfMRV
I3r9oBVMAjxJY2JnIBbj2lYvMTI3z8q0zmH2MHJCZEh/dUI76m8e0qFpr6jUQHS1
QM5+unKtNhDQIoOqODVLlDM5/Vu1hQXal0Yf84qZtQnFA/bV87wdIWMSowgMfWIl
SajrMEvKmkknMQXnC/v5ufLqbJLOCKYA4l6FE7d/WVinwBgHyocTIIv+1ZnNqbsy
K66xkrfrPB+yhxepY7QfdH122by8fEAbDqmMBt3g45f7QgoF9LmdJZE8+TqUx31u
/1nJ1XhWFUjTz3aP8NqJTjRzybgmLW+LVnL4svEcAgxR7Pyp6R+EA41RrqZCpnoW
MsDblcMLDSLFm67g56zSaTFnrCa7FDdgOjAGR750uZHV09abwaBwJBt5JN1zBRbf
jK2QgyGxJ5NfwXlw6/iPbM0svCGGLN80aKRLYWhDwHePnXz/gYrv+5ElX6zjzvwl
TS3IX3Y1HC92mClwFsSx2q0MQOKy5UGapsmN+Ys28TBb1XUmStiPKBZuB9Gw32Ev
lVH9mmM5BrgTzklBtr3svwQU1et3MM0SauibP0rNkJBlv9sLC1d1AokwwIhzKFK6
/t6JHceC6glzIpmLWHwJr4WTa35t9KFWO4W4yiq/FK3uQj3fY09rBATK5ZP1zXdm
NCs0yvBNVlOwS2w0yEcmYqvRDwzaQshYTk1Hjoe8AUCQM1SSDugTft0ZtMyEwEs7
jxFSDhJtXOq6wIsaacAqF2pXG9mWvEQMj4BPhaMnJ8mLe7UEPB4LdWwp9frA9Zoa
yaQZ77nnkuLMnnmHLHrLtPAEvdiEzuU9hi4FmtXXVra4Vx99nnut62MRN5xF8Egy
BBiTHyXMiH78Kc6EWVjslUusw6DpbvW10DLJJqODLQoVeYcZS0Bt6ThnKtAAsxW5
BqDL9VffU8g4x5Z1JtP560R2ftLxiMXXLFlTROevaZpZLWcJqbBJ4/LNO9UFRmO/
hpQitp/ZDOR9XWXExNs+PPJlbKrWnEBkuRAyB6RvwvhfV/IwxrtzjqvtvHcOIwGk
5IMHlE/zp1JI44GMP7IOATlvs5tdFD50wEQAov6L8NLUQPqm5VrL8x2G60TH3d91
doscetGhHunVcX7iSQVLlKJDqq3NMy4fpI12v8TGYmQL69gcfyD3qagKavimye/u
hpoP/QaqZ3x17RHmjYKhAhLTluXWKwM+rSBovSEj+8xr1Nv1w4ERUCxVsn8pFJSm
Rhr2wr4nAHuV6yO4zssXXQSTPYR7lyuLCTNY3nbmscXF8Zr54APYzymsz4Z/pZhV
EfLNJ26rnisxFmhAHvofXHu/MRIhvyBrgQDwq9K5AW2p5ysGHSf8l552lXOPOKbe
1xaMrf2Zcxr5YIUbYP+YEaVX2Fh+ec5f31acCre7bqfV8X/h8KrFmPvqCaAsiaKg
ONXDFFc47+nbz11B3iL+DCHAhicSD9W1b8jLEUAESkEk7OcCcH07wahf6DKRbnY9
`protect END_PROTECTED
