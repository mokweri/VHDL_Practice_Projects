`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bkNZ36vGDgLhcTBpRfl/vCR7JV6VZcLX9GecX8P0+7OLG1IQ/aUAoZTscUqg5gK
yd1u8JRUh/c/jAamb4nL0DmFvtIKbllutXX6OWirloXgOgP9gn9Pd4wcw1/NBhTu
rsMvHf5g+j3k5EUbqECVk5Zr109roDUGIqfukK8kWbUGJTx4hSLBp3PedM/4k48N
bgUMKnvW6tBiY/0NPu5w0dAqmAVAh7TdU5aWrwxPdBlPUllranzvlqwTIHrfGpUQ
nhloLBpquzo6Zz4MinAMyOTvx8hAJAtLFW/610kIRD6P1OCJYRSQhrWz+SthBW0a
nTMxxMhstbs4N2PEEfeVUfPQfwf5GgjUmolUvOpUizq0hN73ySGdCCNxJi5RuWIY
7zl9rpg2+fhqT/Nv/Cq7zriXe1sm5gMSWgZLZ+nEv2nvsNvG/z6KA8GfEVWAGNV5
0Kz+5vpCvgnrgMH3LaIMsQk0OS/X6+1lb7TYiKCcV2p/jZ7F4LFbPiBy2dOjTT8m
H31ncXIELiuuut6jRd6ggITMqbur2fTZ9D59ejtkV+Ul7+YGiANhON5cjWtRFcI4
cyyMMyW9KVx7h6qm7x58h+XIWsVquaM3emfElkb43m4MAELxXHM3feXQgd+mtRTY
spL1ngS9xzbubsxuIAZZ4vcuzuKWnB9JW7u8KslK5+2WiIsHpBsUzt2hl6e76xO8
IwUG6VTuWe4CvJYJ6vCDI8Jk/i4QFa4NK7KJl5OT8ScU4zT2QyJX+5unaV/kFK12
y2k+w9V3quT84S6b/iepI6l8jxvfj7+bxg2pbMuFtoRHYxVogQm0DOkUIUSk/frM
4rnnmP9GZ5X5iKeHZPZtQ23vTnlZtnaOnpL3Rl+v2h3jaUXMShOV7SH5zE8cEUO4
riegC1bjlOlbOcN4kiMiDWDofDoYnsoqvegp4otPlbi387hr6TGopj4CQ1s5YZ3W
kN2EOUX8Cfc8iGYQyhcUQkwAtnHHZQqJKo8xkyO/rbeF+bZcQtEpwB/fconkAtz/
GhS5OL0FfkDS1dJCxxjZ+QF9vAU83nInl/mE+UuyU1/LVqsghk6+N/L7HOK+disL
DS4FbHMmdyrz1bqIH216eWPFEdtyRZegKEFSm+i7OC/nbNhRzA/Y8jnAmRen9nXK
su6wOwVjk5FtuH5OFiirug2mDR48ahVDM1/odmDEMAyilvQCwn6p84h+9yiRWzKg
ZmELl/bELaa8WX3MF4wJ+9/pXPkkJwGmh8Xcj4xcdvCGiLTyxNvj+aUIfiwCsbam
kdnIKRbTUdm0Y6BLMyoF6ts1x8Y3F+yRMSz786+krb8NYRPG8Qtf+tPtc0GmuLmE
foPufywThGMcnhRMTexpmS77bYVs1+3iqk1gwFQKeVofJVqDc2EHy3oFdxWPqYCA
/XyG9j2PKYZ4DrJchh93riD48NSrINYSAhzvHhcA2PRD+A3ks8gMHkZ4zRgM2c+v
`protect END_PROTECTED
