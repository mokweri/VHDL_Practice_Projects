`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sn1OLTT7L2XkVH33y6iqiBz/tRWCL5zbbToGIYEwCuYpZi1M1QOmKhZUym7yTazb
aP+hQPjLic0eC1LG3weJgfwe146K6iHaPRyH6OiWQME4RAlxFE73NeWRiAvfHZXO
54suFldws7WZ6kdMavOX/doorScNqfwWlXMfSBMcnYbqMHELsBOj4RcqUlPh+3az
+OeFZvkSIQrwZ7vnV7Yjo1/t7guGGL5F2VpHCxByqyc2fcdDXBGn6g0qXz6jPfOW
cAtOt8AZzO3TYgYWIliCFf7nMGlnv+8uJTSSBPFLnKwVpxBUFe4C/wnW8wxzqmuK
kthCcA0d3yKF23/OTc3pHC7idDWQnjtZLTRDU1BQa6jxO38hw/MMXi99HoQz/9S1
HiwzggLzc8BYHeuAnJOOXXM3tm8ivsxAldVj+KHXGELqHmji9zjA+wwImcc9L03u
efnuG+WQTrsYg50+Yaf+PhXhJ0ANMJgXjg7EY5WM4sa7C2g6OtLLjurLinU2gzvh
96WyCGfkRu6WmiEuYDjrJxbhlO9CbpTLKv5gBdO8W2KLF37dS7guye/ZmJa1jeoC
RV+c51oKQF4KZyCApofHPw==
`protect END_PROTECTED
