`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vs24/jcf5AoF5mpU7ZOAT2cr3vXdOE84esQgQRDxUNji2XREeJAQkJ/K7Dqtsdnj
dMW8EfLmKqPKRIsAVB2HEKKl7o/Agv694KYEQIOspdvPTCOr30xhJww7EbQ5f+AA
+e/gQz4H3+QWVbhvesNep6fHeCgSMDQm4eivqS8H2pA=
`protect END_PROTECTED
