`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9KN8SP7wkhGCO41YbtIpSY9nPikiNIC26WwNhnlukb6Wd17GjLHYzwcsa4/aYOU
Ree863J5rj5SdrpZwSrwDeNmgMQDP+PGPqqoeWZCE6BtlPk8973pN2AGOWQdzLQO
GxpSLC/jRscHFYFWfPe1J3jXUrbyBOya47MFWll4lc6KnY/PqJqr+tf4+o8G8UTo
dsyJ3tnNZ5AHhTf4q2DS1Ur2cRobaC2RPzW6ra4h7c2TC/VueEvMZxJEgDn/MpB+
lPWN03XRwbhF8O3tg4V6s1iraky+gaNONta2wwUIDZLAnyzakzMZdLYhdzbFE8dG
CIQl4+wTmnvZxuV1wgIcSJhFej7oledREAxb46poQCRCT3mKee0b68yF7f0jAAaP
oS7tGJ+aDKNu/zS6wzMYk+V+QIXMANc781WCVvJj3gXz0oyXYJFDMSFaTvWmAE2c
0cFn9JG34s1iMNMwQ/I/RV1Kk6gEKvp6XU5MOcy01ZOhFk1l69c/7nz+/LgG7o/k
CoX/5fnkX+KKKNomWKsaytXOYhz9MWafcjHM/WCw5Wv5VgzR0bud720ni/IhqTGa
in1dcl4FukvQtTj7EsiLPIPMf63t99ahT7G4oaKcsCIjZ1Iqh1cBevLEDyXpISxN
MrTTj4ojBNii1dkQ2UiWRA0bnPUeg9K9fYKicAbNcm6tuZbY23xsJD4ezfBUVu9Y
M4Irky2yMII6RbaF/gI3zhF5wyHWKxpeaEZzP0zxFS0=
`protect END_PROTECTED
