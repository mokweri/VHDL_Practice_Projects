`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3nqF/2wEGwjPrZIkYxt6y86siYB9ke8VzjQoJFptwvICKiRRs+u2nqd9j5PHgJp7
no8DXhblGTCYPtRSyYEqEHRjl84lTaNYqTQjLkG0lIReR0yYnoaU1tEJDTCN//1T
Pck/130G98G5cEa8oDWTotq9IALVuuqAPQ+RtcREwhQrqzheAnuEqdVq/vWTvVkL
VFzm5chcT3ayuhRhL0izxO285rRdV1u4lfu/7W0/r8v9aTU1bVuNxdaIdk5pbByH
K1bGd232yaEpi5Ruv1RwBu8x8IXQQThZcLfe6+XSkDE96ytgVOaKnuk1WK99PlgE
Dgr0GLVRN0ihoSRR1/rAcn4CBqefoy6Pm5gsSJKwmlXD8GXCOwxoagcIjcRHwIhX
ClV+cu99GBXKytVKiHM3scJB+J4SfVMHe/45Wm8U4GkXiT17oNwcBt/L6CTFxGhy
/1GVJGQoUAG6x3UagGh9WBv+jYxMZCgRwJJR93DRh7vxyPCE6jyxz/PWgy00NXJH
WseCr9f77283q8hANduLwlfkAXcoWMsWP5IeCnnTjxg3M7ij+UH8d/h4N3nPzlYf
v10Dl8YiSBDTUxm85kelnRiK0kInwaCHfZ6G1rMtvE24+FNbRgEiJTxocJMEpOag
+PhhgBqmlV28yOHMmZEyFvdAPtpgLr9w/zlNlDFxFbCqAFZym0zRVmCDW0rB/Nwy
o7poxC/wi6scMmukXSOczGTHlvgURfdCYLkeILFNXzdGDzbwH6kyUS6WrVsYT+eM
DDXdGa6id+kktS/sK5kdnJSWWdllCDlYZdMTqy0e4YC3wdBzlA+vS05ByQIJta03
ud7kGxgn+5JYBgXm3TyFQ3bPRJY6e/KjKXvLlvVjTym0rmrzF1d8kJEomjZZPbin
qdq4BiU/vCq7vSJEPyi2j7lL893a8nmspfPeLLKm2sgKmSuETrCwPXeuOdZsy/RD
HESU3TnW45nG3o+UsLFwnnI0NtwAwuVgIPSkMpGCCnGbD8j1bqmCtO8ez4GviN+s
bG53Y++xQRxVY7p9swhlc9dSXFMrJ+gwLtXNAnlEkVTHvIk/kekmaJIdfrlx/2cu
qp6+uh4nAHoXvwpuCJvRiQ==
`protect END_PROTECTED
