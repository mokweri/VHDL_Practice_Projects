`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xlceM/5NJny6WSWCYzOnvcV70o025WxEDktt4YYKV0bLtc07Q7rs31QR5akqDqo
Eu0O4k/DfeGHH/y1CyoaRaIJujgfy+kKtdBn7u9rMz1q11z4fzRIQ8yE93kiVHs8
r14lYoBGKRVKqsc1JzPjTEJXvB2qG29VsTVmu3X8aVoGYXxVH/OCtLTlCnjFfJgl
0r/y4QNA4kJfrubNvaBROGxFyxde0JwfDU3sS9uNjg4VdXO9Ws8r+6z7dr6ZRPfu
E+mSiIUg+f7UEQhajiWmZUD3t9Luz2hcraJC2zp8qxr3cOG9iMT+0iNk765aMANx
swJ8mhfupJ+HSCUXB6WNuMy8iniy1tOOEN6vDt6ZM17Z8jzZHW4xikwUcxGDzYf3
ynM56tSDe5pTitLMbiQh+QH0VGjE5Y16rGF0ucIzJ4N3ER+TmqtOiPwiN8J6PiA+
dmMAGjGNMhWUxqCP0K1Y3+hJAuibDsZKni0oCkVmshdSefEa65FMsLs7QKwVkkJI
qbD3D7KELZXuy9Y28OnwOzjiLyVsBI/Yi7kdscl1qaGT+SnUsM+Agi8zDFhAIXVs
h4n6FlTcjkUCdC64zWVP4/FtReMaoEagHMQCk8ci79fapDMBObscA2hiGKViJBRL
Gmek/4RhdASltA/OFtex1Rh5hXnPPvd2N7/JHyi9NVJRkFCu7U2KWCEs2nm9Jcsz
b9MmR70ZKvNSw1TS5LMlEqdID1iABmmjrXHcL8jhlLO1de5glt3GZPhXF293GCUJ
3TQa7oQiP1uK13M0ldZOBQAkKmuaimtOtyfHVQ79v3yS23qHjDZpEXpg5EWDjM9h
unE9+9E0/zkb7Mt0qPkLAEEXDZmKkqXpepohfRubD90WDN3q7JPjkEWZgwHBxSPd
`protect END_PROTECTED
