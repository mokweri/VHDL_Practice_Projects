`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+x9Bk+Vl9Ik5mfMXUSuObrd11QRHLE5jPs1Ryk9IGj8KRrifi4ObGTD0X/r56Fe
Fs7yyWp6YvG1FwVBGnX5tyIOIOrte408+NUuLoX/JeqzY7q2Fzje6Birwl20YgU0
t8d93BaDH01D7NedGgp6Pqd8vYiTGJa1i9GR6ORvLgAYRDVGRjpHR3lEj7/owAA+
AEZk/W6Ty4E5uA/hlr8D9NHVK/etOHLS59dhiPvsK5+yCuh0ObX8cDHFWWIiNDA5
jPOHxuWRGLQA5df07ZHBtuA4Nffxxn5lPTcfjDzhu/I9AOonkwvMIFPidaiWBfE6
+iRi713uolCB1Qu/taF6uPSR5o5IjtKNODncqu9TlhU/xmdJjRUVt+RCgVpt1GsW
NbnJxahCxqvoJhyFKDH0I6XYv9Sae605N7/RRHC+fwOTI4cPImpzCy1xJdHn6tiD
u0UfzFL46i5kw71RpgXQswPxLrIIqtPNUaxb7mQXpzoAoKfIxiu0Z4/BRvyCtk6u
EKU4p8Z30Y2yR5oNKbAgHsYJbCqzOep0lCN4z6x+PvJGdKQUF2+gdNbIS/n/q/sM
mh6kNNowL+Kq8NPhkXlQ/T8ejN466CrOQxmVcAdl2SmDb6Sn6FikvQsqzKgburiO
YDtnaqM8lSLuGijcgpmY3cr0BGX1uoRKySIxHy18EM+o+tUg0GUy2heQG9zkBoNs
Mzl+uh2JYqpntEa0ZrUzGi/jsgOzOfpNvQolkTT0LkazbdLQvQ7bUW/LXpZ6v+BA
zMjd5Fir+/k4+u/RGkRREbHkAHF7+XHCXkYhlsMjqMrLcSRiq99O9G/tl6Qx4Wfr
jSSQGlAYq8jyhT7IffCWop7OBeTR8OkKDPiiDpUa9Zs5q/LBaBBLziYxcn5/6h+8
QAIp162f4X7NbABpl95yWGJrZCu30mxsurT0222BW0TJFXrc8NK6tOBM35fA32XX
QCAD2k4zKw0uC3MXkNjxQR9gPSVYhC2OlqBi4i0p03cQD/WfPn51Ianeo1J3lcc5
6LMJTFpzQ53Hi8JcxdzRUVd72Bon+Igt0/2hbY6La2z6/9m5Fd0gFScvrf0qVi6c
Hz9PqH8jntU2HROrKC738PKkE2b1uGTELOtD/v6pb4X7OumyU1bB3FYB7icW1cea
UwqF/xMy/DtLcmcGKlIms7Bwwd2/hlXvrsXh13QJU7hwnwYcyDvWb6syDU9kNt2B
RSaLY7wcHpYO2IblbkI939sN3OKaxu5+mLc7OiJbixckWY49yNseNCydTxNRG7on
QaWa0GzXpFMUHOsxLFlQQ6RhvgOIMfIn7VXAJxS1EVTG5/+CG+zXVIrUnEW0vqwd
Qx73E03PdF3dVm3bDy0GvNX98eMN1Dq1v/GZ1ckqd3OcaLgVW3f2BEEV0v9YdE+B
ZxosLpuJ1OCnOI34b/gp1ZGHMz161dclO3TxbyHhTiS0jv3FhC6TLB+4Z/tB5ZEY
dMz8ZX2iqNXn3eHeGvGYaorRsQVPMcDoLTbcCA9mFPiDeJ6powP8JS7jhlw5+2AM
mUSWxR4gMfimkxJ2TBUSoZUI6ZbLiJpJsgM6DtnmoLrf0XPuf03WyEMBFlgpolgN
gfAVPROckAmsiHj0Bv099R9Gt/0DSjxPHfmb6bXbk45leuiNW7seeAqQ+YDBLwEe
v2qNU+bvCapRRRZQ27V1pi+Syz7guPkBGcr+gsCdrveMSK3bhmeeYkwXexZ986+p
dH9ByH7NizA26RF8mOLNkRYT+3f+ig2Hid+xTK5jVv0iuOrydx8ykRKMm6R5jH+v
WqoRXiJVrSkDWu5e/diL6MTB1J9L2BNCkRe4egznQdAcqP4EznNKCR1fIDVJXAF0
sWR+1TwQmKNrk/ZZKRMob+NFMEhx3cLEf07LUXLBfYWeKAT1ujmC5TXGaRqnEs2n
B1vk66M24getkwgk1xP9PvKbPw5VyK10DOLZ01ey6maWXX19T58Uinn05kf1o2w9
3agpXWSos5UoLmxclST4QLWlvZOWVTFQXnaRPay1EyuZ8JzwvCH7b6tPIyp9dM6E
7WiE7EhV5peZy444VOPJ7jLQRyBA2pjSPMEoQH8JnSzWcBalEDo80MSpbw+gEDaD
LEhQYJlaW/Zg0P7QdSdHlfaWNGul4a/Eou/k/WsjmKxegZuH1P1T3eue2BsgX/BU
xsXSyiHiXyX1ohetYwoX2lhE5rw9TJg9dhlh7+1/a4ZLB4mepUFLdFKkWvwBtHYu
+4+aC6zNXNu8J7X1HrdB8e/JWC2/lt4MZ1gwkrAahGS/I5j421HW+h01wGFEsQPT
dA+zaw0weiS0ABAreUlVEXGbMoC6NESQBJC3/0lpBKEP66EIEQbVwa0qLGHCiGjf
GzcjtTG7pgWkmqQqDtXbBkosSyF0y7YHJvqYJnxI97IwANApOz93xt1aYmX+vgrT
zDrZaneEuaZgQDI0pHmLKPg8eymyOrkAtSYrqhafKrD0Pfl7+/AyxPTdBRoVTTW3
aWyOHvDqL3ZGTzOYtdckXg==
`protect END_PROTECTED
