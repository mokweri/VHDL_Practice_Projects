`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zAnjaXaH7rG9P3OT4QnI11RmqXFK++7LblRQzSth0DNMPV+3Rlz3nj2i2ND2HD9I
a198QXBREMzDtQpF94YgnmQMJ1cHd6ppVcJOGdln1c473yxM69/9+TO1MrGIiSHd
x1UXVWZKReZCyYuGLhKVIfzasK2N/1MEDGl11ul+fvCN508qRMyzE/IBZyTqFP3a
fJjYoJqq7WJDVs+5zP0QVGq0gQwOBeXPTWN07cCj2GKren4XqCcE8EG3qLY5O/K3
wfOEuaod+0P4k1/xQyWSNhxPqfOWgZuqHbMcpoYoE49/5BUsdm8hH/AbCvy9YC7X
EfWrm3exEfJZoy+QmmC0SPDw/Q4D5usSUVUM9Z72WqrlKdiSCEcw3YFUQLg9r/b4
xzNC//V8UBVSl8HYzhP+IEa/+lLeiAML3G9G2Cat67A9RCHeZBJuADIYPgviJt/7
2EZzMZNSk47/J4uG3W9+DBU8lI2caIM+xQz3aGMWZkCvPHBumqc1nnvz8Zve1phI
OtmuqA0RVGAaq8BGVe8jZLETXmhgQV56/fSphiBoutorZreiiuoB9ouQKzXz/GDy
Av9Pfv35Oq5Fc/slQmLUuXTQSb7fMipWpsPFYblociSpCazcyv9Uk8BkTyiLKjtD
+042S/n/lKEozoc++NfMLperfVtVIHnXLBj2gSzpc9ZOpaW60mqqMaTXCFJ713xB
GHMHrR7AtZIz+ScX9sF43xp0ZisFNq7JnubOZR5BDEVKbwPVokWlKYOmMLyzIMrI
Dk/qFfSTJ+VtpIXfAPgIdlgj+jivspY66ilIru4arEXp/yRIfKKFIKWXkcYOi/kG
QG03qC2wmPp/rlWzGcurU7pG0Hvk0eD5v/6HrZsdlW3hIyWI79WgC3b0dBujdVOr
kRSeh3135Tov21agDXYIF6PAoyViaQgYy1/eByRAq00ZlKjwA4sOyGJg4aZnrzYH
W+pwds02/1MQZwhnVeJjux/IAn1mRff0P64LOadH/vstltOUhmrQuWDWfCMJzWyT
N2cT2S0mhFmVsI4NIUoAjASEW2dKJagnY/HxYiaSNMV7U1Lp9f1iDRrC/c+B1Xmy
cBME4MXw61oF3CP1K10cWphe77KAftjdhQPzVr+9WwaN5sRXlYmiAa1fzd6FC77w
QNP7s25WQCB4PN9fXtN2klV2e6w+bov54Ky6tqJY6LNA+5O/8OnL/bwlGmROZVqJ
t+N7QH2Unk3v3lqS9GGjQMcpeHlS4GM4gd86bSgY/N1Uo/dDcZbifVhLanrwRX3l
FkFGmgrcynP/7dBPqqnN4WMUDHYQUgtGFFxFGL5jtMM1e3Y/wm1HK8FSdcqF3jVu
vxief590DekediJlq5UjaOOjQ/4Vq7ObhAvt7ZVV5GdYNgtnE7mSMLIv/QTN3e54
tfmhuj03IY4BY63marOezcXUprZ+axEz/tnjd+IyjyS3dd7cW6fOYMeI1HKLQG2+
eNeLvt68wRQqI7XEukPknv1lnKxW+V7EmrQrVXMBsaOnOcpHiK73CA+EMFi0EWy2
aBwL9xHzeIu9DIEIsdei1QBg8ot/aEmKr/DQRqt3HgTRhRCI3dfRTJKfjGxKnAz8
COHLCFqaNTVcZ8HHDzbWwPqDUaIERc94K4oD1jb3vTI9leEAuPl2s9AmBX3FqMWI
PwFaeDyAJ8YkXbtNPUDQspZh9uuiJfHlLLxktMjfWT+Duk9Jyum5demoG8bVtcxe
lBuLIBPwNkkI8e4izeQFap31wDQ6icazW0/2WWp6tfTwMq4dt+xeo6ojvYF4wGmV
Y1Xf8FksX5TXUmvkPT0Ex3MZHxPY9VvGJ8GNTfoizO8ncHS0D9FvvkESkxXLh1Ho
nfLc+XrUW0RtQ2yRfzQz5V5LP0un9ib8UumfzEapRJPPULg7+JGPi5aWMqI9rggv
69OSaX67QTuIxf0gyRi/I9EdGoh7VlszUg/1RaEpwnIjx+ZpsCqdJ5/wtAb6Wued
v0zmRMejxpnIMlitfeKqaR+uQqEXIF9qc+v3Nn/lJbFBA8LgceZONrX718Dhchis
Rwybp6bCQLe6wiwOVNjkxYstn63GuHKKPVNVaD/L1wEfDmus2qypSvNi2SECN2gD
piYVMFEW+Xzs7Pmy5kz75yzkbi3xzpXHyfWFMw0oiZMCAqjG7/jyuu33ZFeQPvfm
ZG2Ce8fH9zPhvgoF02LCdpNVVt42bvEkHZvdnr9wbI3i/6suBP2xXpcpkZXc8+EB
zcu8DYUKQmstqaD9FooslsBERaXJULzULZOxeMO65akFRmJYuMb/aOMBuEXMj8B5
6fuWdpFzGCC/eaooJRnAzTTFaSVYdl5Hl+QGWlIcBr5EnanpU+s4M4BqxAhLl0MA
qtVLeAL0EwNnJlWts2ZuT7mu910Bu/+gvKC1Cle40009xVUJtLim40EibQpISOZm
+lvwOeq8YILGRhkofjpPXFqvbS88H6pWy5XJC2S39EQbPbf+UMj/byU2zQPBJwOM
BzgY/tEKaPwJgZjsWXop5TE1mlVPKnoQ4XPrF+IMULU=
`protect END_PROTECTED
