`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMimCj70JysC4ZnErLyQ8XxsDTaKx1UtaoZd3MKtqqwgHjDxjo0Eiemg/wphjoYl
L/+2cZf6NUid0J/tYffix6mCqP9t5WZHmJudV+d+3nUKEiV5MJnw5NbvwbedircY
+VNFkKU6aZhe9gS6IYMyzCphbaYv9FKgbR4hYwhzSouKea4xDzUcEAi4E4FuEMvJ
1tKjw9mOFnj7VSllMJMPL0EO19VPA4Jx35Anx0J/Q75UCDM5549Kj6syPSmPMKq2
ZLJlIegQBZ9u44LJVK96tM0zxGijWI8x7S/+rU3EViCxJ9pVP9SEZ52HQNAc2J3+
gfl8Sp2sej85QDHXXwTyuqcjMl4ATzES6JhzZRYvVYMA+7ZBuE4C+aJvMG30tF6K
a4slrGEEtHDOUXznlip8y1LorUh15+BzPf7DAZWVdRzrelKoeSZ3/vNO0Bft0BKp
JvkhLPNS9NwdLVaHsbj/8N0eMkeMGmw7Ur/osPj5uqNj1aHcLpH/UIzMzkUw03QJ
YX+2rpNt4EDr4qQYdwdzsXrw++Uqev31JZfdRN6piQwRrbm+277uQsV9gVUJTw0m
72zJ1F7cJ02sbVJBwql9I37rzFnL9RUfVC4sKKNxD3AU0l0iak/Iv9X+gd5iLhAC
x1nxS+PF3Jlh1myAb762869mg45oz2nalQ3c+/pEqCnIq6TX+vi86LgymH/Ec2WW
L5qczCoXFb3bw6R0TLuD5fDI1CEqJkitJHzJmYgiub+eofedOJxa40IXg+oIQs2z
74SpSVqnpRRePfvLzC7H0g==
`protect END_PROTECTED
