`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TE0hCEbw13jeXIb/niSfAVyLyMg5rfoNX2vxvZSYLJHMRNGjpj0ZYVTC9gkP2JUJ
DXHf7YRiKRY4uI0FUyFk9rj2RwZBxvLyODsWeTD6fW1f5EfLKZ4DjTLWCNyylgKA
pVP6DL4+MDoaZo2sScS5uTZTypV3bBPKi87g4Y76zMQbfgnHNIssaQ04wZbSxvtR
7Hb9Fu7h85m8hGLW8afgrFvewu0LtbaCfNFmYrgyUrjoPkLwjEO9c8nY+XaGN4sw
xIinDjYQBObK8SIoAF57ED/eo9UoCRIrI2beAGRaHpc5Tgp2bNTWbk67fJBnYWeM
fnAlFBit+3xZqFz8+hdR+Zgua8y+7ore8ZtYx4LWGane10eDzg3RJ2ZRkh7VDGsK
CjAwpc9WFXjSucUoQDHc2Vpr46klh3zqVADvhEfL+zY2pFrZphkLkGtlKqFiv1I5
/g3myenPZKEbhKmFr3dcFnzOzsoW/t0wOpz62/unV3GrBSmhjw9giwXw+5fY89ij
eWj+CxqEw4/bIXhLB2L6jw==
`protect END_PROTECTED
