`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ToQ08B8Kxm66MDkAoerewIUN+aPG9ymxRFr3kXTC0Rv1jMNqFQuHDZ+CST3+VX9P
fH85chsDxlN6t/r5ofJTIOLJKAbV9a+jfwjOnGHNolvirgW3kOSTeTuXp0kMdSZa
H4jZqfBP3MdT+O2xDb1hKv1ErHn1Rp88AR6mD10RahJd7NBaCTEfd2CfrNqxENnD
IIEZI8rVUKAkAcRvuxk9mJXFRtuPnz90CMiCAZtxeee5YsYesjfZ5XFsy8j6q2Zu
u4MWYa4addv7zvNOSREjjHteJTUzkE3tC3bAhQEUKqjQlleAcjX9FgYbwlczAqBM
ulYvFcfrzUhdJ51UA16XSUVZZx3Vpr+/ZOdQ/G90ALUYwkOmZlLGz8qWUShaUTQH
/AfRi+HP5Tn7BrihQocusxV49cCpWgee0Qk3vL+P0mkNFYdJaHN9ZaGz6xIO4dkp
Vkl5bnQB9p+GS5zN9ntjjtDbbD5TAXkVpmYtZIahmLojehTmaCyj/an7dD54/dsR
/xtIotbMzAiE7ZctFljVMQ+LU6r1XaPmWDz00HpEU6EfoEYkEsJD90fBLzc9wcYJ
bSI98bvWQto+0znGEwD/uAOAhpFLK0QXNJRzati8jBGtrrvYTe7bLybSyLwGpYct
i2XHjdcHPAB8q86V+IMGwTBgoReCajxgtnBIhM9CWGhzG/dIBxcQ2B4LxfTv7iDZ
aEb0IHiE4VeMRcji26kshSXfjTh+/uC4VnXwaYJ9g1MbOuIECg5jk2zpaa+B9ULq
NInMtbPaHwPnrzraxFvD/RITqffgWo14ME6L4wNsp+AAMH72Tr52L8GV/zGkP+c1
lVq4zDbd3GYqEdAREW4P+WciNKKHnjaYtGo7Wke5knlonwmPy0+JfVkkiOB8DeZf
9StlcMJ1LCGJO7p1tCN7Gdl+srVLkRrT6kegjm5l8tPj1eh48F1Ue3PhgvAJ8+yS
Lr8ur5yv+4FH4R1wVlwcrdV2BfL/jtF5vs1mHqrPQXIFR3YrtdpWbwgRliqR0pgO
8siaz0BE0pYkO9aW2UZ9yRoHGDLfmSWnea1kGQgdpSFhIhW7XZNTSWVpZjWkzFBL
+6OHhJG+8F0vEaZqrHCbmaJJoJjJ6INYRdTdsBCkDSg+Lr5s9mpryn/Ps3xpxkww
Bm6goTUrjnl+BxxmRTcTrFuyKgdr3AItkY6jrwftYbulCPMfyGSRZPnPdg0UgmIU
uJ7PrKj61K1cmksk8mBGaK72fJdd3LLc6JK7iEDtUFyqrq41ct3J1/oYUmeuge/k
XBSak31frSwjOSQt5dCLbQ==
`protect END_PROTECTED
