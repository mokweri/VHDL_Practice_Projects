`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1g0WflVjKUXOch6RkeUwEJSsQ/GZF8NXveoqx5zxmQ4RKFNlseei8nCmbqxD40dp
YNCmjMT8sC2VEP5O8JakaYrrIVkLbRU6BMOPizzFcEFs9re1TNa8wc6nbEV/3Okk
WTYc81DUEggUPKB4zQtDOxohytbj0Ocu6w/+2aeYQAJs8y73cZVroV3+cob1VldR
lBKwwQQ+x14jWC4skfLKMzOA8+6NHmH7HX0/X7spDPQqYqS0jPWSsrWiRpspWdPI
L2gCinzvXYrzr6934qkT4We0W20WaIPBXl7efQTe94vQxsFa6T0sUIWjuUED/W70
vEu9gAUEY/Wzv2XmC81t6Bfm6EResnM3LqFqz7sMwKg/FhGmbkDdUAkWlWYeYllv
WReFcepdEu6ggZ45x8UYF/jtAT55cLhwkAGqfkBAJetODmU16YvUJ6iXMvM8rZl3
fqe2TisfXJsltnzO6Vsyp2ZpPyO6kWsI86jDkGETtQV78p9ZJdlX7XenH4RWt06z
TyEbMUL3KWvvKamw/+uNgVllqZSg12tVQCIpVq5oeblQ8mvD1+ILoIU6JeASc7NP
+AiUjMmgOAVHlaWVs+672cqMOp/DoJpqCS59jXh7S/pd6oyTVUZvl1Ymv5ghUM1S
zH3dRBOJXFEVal+xHY6rG0CAxTPMOPxIyFO/I4qmjP4NuhE5f6IiW7ysqkT+9Oel
P5PjW0rsNMCGlH3s8Os2fbbx9xizMffbCKCX4BtB+KkL1hdnKLJ6zaxH6IDA89xR
Ar2QOsyxn+Cx55z+bwgEmIMeghpWKJ7DDHqBWyoAsVVVRARVawK8ErUd5wLtOj2g
cqAmLU/ARnu4KWddPUndZ5JS9jRE/Li4jtApE/LJuuors+BbrFk0VLbAN67iDSoR
0K337GaRU/fLlHnR2uv+GWJijBF4/srOW7maAYIEgzo=
`protect END_PROTECTED
