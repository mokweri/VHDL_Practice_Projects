`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T6wCSbay2KoNpp3bd7RTgU63w+eRUIDaRMduv2toclmikkYiKaijxXwOagHPlWfY
cQcUr4XZ/3GsPXaQmeuKy8yt9lvupdTSJyMIfZme3ytNhKsZnMdaCtzQwbFSvMov
PwndhBkJMNBNzL7ulQdSdc6SOGTQn/ZkPSgDta8mCO1eBawtu1dBdNpl+3Oq13O8
LXC/nE2UXuNB2ZmFqVVtAyg+8KSft6bjR4Ha1DUC4vukf6pipFv4ruEAwFRcxs+D
/ILpsc9VJYFhpL3ivqshQ0UJZu/lsw5IIZ1p1DdWyRl4joFRu+jIVLVZxNIb+QJN
AsN079q/ynjIlK9iRLZnkqKffmwAPh2iiwWWkxRKqLBNPE2RROhSvcqvJ4xkWD1i
I+6xx4Ua6RzZPSXFjGl3czvPIYAK0giW+o3+I3Td4yK6rQ2zOG+MTkuC9OFzcYtr
clE9L0cSGzbKNFnSuCeeQHdHOlbqrPyW24Zj4b0wtQ2BATpm2LCD/IYpbo0gEO7Y
`protect END_PROTECTED
