`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jZcUGeAhauOUk6Lqyba4CsYPxuKwMTDtS+x17KN+/LApTPpOu+TlxX7mC+G9F66q
/fZI++MIvDf1jtudzVbZqvwEPd9LRetJf5e5/MPawvg5GM7T0GiSvboZCc3/0O3n
kycHNLU7gozRg+j8MBnYceLdOuSvZPLL35E2beP0yDit7MpinOIJUAXzVGPOiJyp
cjq3wnNwkr8g6Wj/rCzyfz++4/IudyLbRVkrSUjAnLNzKrC2ARxjtmfkHwlv7JcH
J4HVMSXYbopqfAlPDAKuoZyVmb1wjhIM+AeYnqNsyE3KcpAHzHgqaG7Wavq+p7bg
8so0QBjDBOZ8s0xoqofDEKeqiZj86i5gbh/l141BTH8cuWHhoOo94Uska0ra8RJ+
TioWGL81+m4i+cKrTQDb+y1+ejZ8W4SB+6Gzvcb/hJ9z+JTOAgQRy6RuPtr3qFhF
hLxdkdC6w/imx4rKJ1RkTFQSQg7rh7k23jleIa1bvTuZtyw9X4zNuGQVRAswB60m
dfEAYtG7BwYkdBD1mVknJ8KkJSyo9hltEF7NeArjHjFWvwrztusA1T4YouFfVpEU
sVK98PAaLf35WlQnQivf0XQXu1lgovfJg8osqeyx8QEkEfoFZlT16G6wQ7AC74GY
AUUYZXXhpq9P32hIet/yT/cCCHtWEt3cLIMNFGkuPqYHRqMkH2Olfh63KB2o1M2I
y9LvdfrTibBUvJhPUAT5kOJmgt3LGuD6kFr1GsB/NYBS4Jz6k6LfdXQYf5s2qYuw
S2J7wlXHUbHp3/l1++69jzA8XP1aDhLoQzWelQ8RYAcQQp+t2np6jTNkzjhvWuKi
`protect END_PROTECTED
