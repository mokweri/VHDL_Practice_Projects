`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3kVIp/gP48aJySIJEDpYzgzGwM3EoYinq85PrdaJy343QdjVA6wyu2bNfzIPrtr
L13V5/UtX8wB1ZWFVWePydNZVGDtCgas9PfDsMh2y4QjOh2SxBK0BhF/HaDwZ9GY
sO7rVQdGUKvnl56Nc51p83KTDl+ZszFj3TDrmMBMhUqhrkk69zvisH9Wqmr3gk4d
QpVl6g9idqVrkGLLJVKwHAfR+VdqMZJOZ05ejCNFS/K1WtCxJ5AaaiQd9SRm3v46
q/5+qAhz6VO8TEI4vGXfg06Q0e8pf62OLmcrWlO4g3c/UfCb686Zs0WncciBAhvb
T0J81sm3bWPdLqIGr1My2mukDZdjcSidLBW7yxlEMHfY0dI69E71mjoLuUjQqKwU
Q1y4CKnz/MPKR5mvEnv5FKIa9rmS4Mnp7NOaM+Jj50QlymWFbvGBNGkucs49RQkF
t1uLg5qFHw7AtsMEMXDiAcNy1pBH2R+legqggiUy3gYxbbsxTsVSjO6KqbQCrMtA
qH0ujp+aLQqHzYDlyjOULU45A/nO9nAGEUL1mB0me2+FJOeYJQfZ9AUXnZKVg5Is
NSZPIcj+8sA4xbipQCrxq7YzGYLshy5ZK14oxaAfZ2TJMliRdDvzwbDkTT50Q4rT
n8JKnNMQ3zePYp+gfSNpngOEfm5y9cIInNk8G5LvzhzAGIJIHA5vjYjQ5Y7J4zUK
T+4sDfNAe79tZZEWhbIcYrVllN84KtT2DCDWsmKC+bs4CEkhUPGJNL1l409BBdA0
eyb0CCOlIeWbOFD7NBNKG52gLonoTZwSRaiq49VlmZenRZXEAX9/ZDyylqPS/nky
x5+odTNsK0lxNgUHqh/Mr+1tYGmVc5ynjAHmIhwpohbWw5tDGRqYEkE2Xqxuiv6g
9NeX075ATAW+wtNUT3ny3nJVTXmxhMz90irecsGmtahrpSPQ6FsZAu9plOOB0FEg
KZCKGhgvWAzX1cqS0QzFetH1/ff/EkNiRKFYFKv3Ur5eAX8qULBW+79XTO4EKP6y
zciwHtg6KgEwxeIuaoCNYEu7xyK+aKuhES/2/HN3hPRvL1LSZS6ur5QmmqKxVsG6
sGnxYbSaAVAc0maZV5KCJ/5j5fbDPPERiSqAhVuJiIHoWqO3VNTfvmLs5oN91Sig
HyeTfmofh2SVWjr+1AxORwbLkkwQnbBt/PsQtNqZN1xHKH0VZKcQagAlSUh6pRJ9
OSED+G/15bJI+N1Q9yaJ9qijhNmQN9nFimO2oD9OC5vIG+cUY22GoXv5JOeb+9WA
bptDs/1m43r2ICSEnzfzeIdXIp4dLqKng4PSSkRYeEq4REA5IhHxT6NjS90TDvYK
klsdYhdDMKBl/ksGMksDBo0EbE40yuSMdmgzHoSsMk4sgtiuhA9X6NvPQ6GZiH2a
PXFQQXFrOYIL8iuoYG/xm8Yya/61mVniy6SAoPMw0SQyYqCyaDlLVm26z7yysirR
xOLFCWLPM4xy4UCCGsXb9AoLzsh4zyJ9XdQM/HmHU70l9hFl2m1fBzgCm64swD/s
PC2zBNYlSL2q572snEvhXn/vEb7htgcjsCCdTurzEfzKtccGg43eBQFvTZJpksn7
8f3kBYQjNCYqEbNy3HKbuZFWTkhHMv16dPJSUye7/Nqo7E5tRHD2fDxyCt3sG1by
rS4i8/40xK+Q9zxz16Xue8n5sbSEovVVlhZ/tsDnhm8NSSP0aSJaCtMsQpe1oTUK
atxPQvH0RivjMVqXxbRvhAOcZcAId0CoXywwHygtc0yPMvSv8RCxv0BfbSkG+p7u
O5GK+tMC+ur88RAEBFVgKGPJLdLHZQRYkoxnFXtEIHHe5JJiw5CMSSw7Et6BlNWB
ijHXzkvKWB2lHwGa9VZ8l42oQZ1Vh9CfFNXAdlfBe6tZGOcMEwJOqdNFrg80JFJt
gfg1KpyfRYEOGMZzV5FZsuqidWr06JN2T1yV400m/VUZY3QxhgRmlbMkaqyMVj3b
wAin4MAZpigzNCAT2NYD93x+r3P8n1halHybxo1C5UXwLxmsDO3qWbRqAuP7F7KD
rp7sN+UleMXQOhGqsNqVnE4LI85bifbVhVMXNLuU+kjAYHqtknDWtz8CO8mf6SAg
Qfve3/VnJ/Yx/u8D035DSVbrLnSOnTKAFzSSSHVJHoeSVixdzxeLxqJvJXplucw2
okDUlOvnTIQ6Ikn3YV5hRHPqS9yASDwfkr/R5yK88Jo=
`protect END_PROTECTED
