`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CqUxxfl9vQJgP3SSXHsThQD57B5rqvn/15rzoEexbNbcTla7TSNItetfEr/nPJC
g/kS4rZTfbpw01mRdspoGCm3ADyjp/NhMyHP52AG4O7gSjHXg0ILCmUj15lBO2eq
9ppSATjn/bLukX/wCiwiTS30eFTMl1Y+/UuzJPHcjLiBs1bbFIKQY+ZFTGIafcPG
wj5S/6BPQnNOo3/drXeNTd0KgsPlLonQkA7Hcb4RPWV8WrXw/opfiGpIY6FBfvcZ
YkmISryOsfW5K+A4QjZ1YFANjkUaIOQ2ur42HJS5uoSZFodTUaisXfG436otd9bA
tcia1IVaeXB9On98JB1auNxl5FfJmg9bmdrWqQ5kgl1nkGcXyfih+988y5a5Gh51
Zd6lGyYbq8ehH9xjT8IzZHe69wg9nTEGGI8CQ/UyBDpZheFW3rKLk9IalZBQJvct
OG8FMF4l5XYXD1ZuE3/G0HLM7GHrVsxaX9WHbah3rZw4rtBGtKx7l+j+doMbhRWK
vNPZLJ2rWx66EvEYiyx31kr7YvoMXHAOx67qWXJ9JlPP763P4eT+jwZuR5RG070x
ahK+kcSDWV2LnnUKObXwdlOC7OFB7CWtdRJ242ODKbnHqdLma7zlHV4hQ5kftL/M
l4eQqLbC4osb80nfPMvkRJcDI/jx41xJmzS2boQBOlwrYzhQTScgJqoywMDPsXsT
Hn2boldfs+ozO9k3fIrmA8dJD9VjPwIw/uWzqvRtIk/whJm4OxqTdQR2CWhnNUvr
yqeVeKJDXsNbdNZHoyZPF32lunhAV0g6z3cP65CSpyHOTES8/9WH2TT8i1oKDZqa
jNiAZgPDVEHNDFNlokb2vBRXo9JzrhIM7Qoh5bEdJn8kHzpf2hixb4KToML+uNaE
qz9E+GLyH4jhgF/3A0z50ZBcUcMM8aDeXGHSufuYsIgifWxl3pKBf1Vkn4D5XqQj
ViV5eZERC4dLxFRk1O9vUweQYjBSMvWdVXrJsgagiq3/+EPu1h13iIpGkRMRBRcu
5db263TPtF3wC75IMB/SpyuCqsNycYiBjyf3UsH+i88S8cSjPGXW+EMUMPr4yW8I
y2XDq+wJW7OfjyuMmZ8PGIOHIbZdRmXediCVmvBmA5CZDI8ldbqvW8PvsV7yDN5g
dG4q0wZv0TPKxzg64hMOMMRQNXpvXwrmf9Zq2Qjy7bpPWmq4J7Vw7L6pZsEf+t86
3Po5uUPlb4gEDNgSTeStP8mBpksGV7EAN5aDILKig9nVVHAuy1Fs/bqdCbZ9PYDe
lv4a0MQHXm8uNjkukOd5MeM30I5gPmwtX5WmeXufTHi5t9Cg1ERF/nBxbVqlsWUe
JE22nSWZEmwn3xAdCh5V/gVA0yPhUcXngXhlkydmolXDJzQOFYcLQb7vxcqk84A9
8K8svX5iyZCZcL7K2sxscV8wdSbH0j370niXP0FfxL1sj4xbvJdy50I2ZUx1saLr
zD+HnWmdxdnHTUHl8SFQ/h3DZ0Al7qWkJbKz62atp9nePLLCJMnJ9sqh8BPlqOMt
VB4Uji3KOUe1PV5tWLDknGvQ39QE2E5p/Ksnoj3bisXxh3LY7vH+a0lbEoqRYRiA
zQMNNK6c/ygdpgmvMP+aOrgYVheKSwPdSKbIcjsoK3c9XI4G7wPmVGXZJipSvIt9
WLV0beUrp8iwmu/xkNTc9Vi9UeQUljqEgH0Kx9O6tCo0zPFMEPJV6yRkWclI4KQq
dV9FWJnX8315R0S48YRKaLNvIuyvj5itPEWcFKaGLqaGgwuhGuDK4Q4Uacmfw00C
EflE2IbgLkcw9POev39ujUVZArd+zaCWoqFhTtFEyUsHo4PSjjLYGq0YzYC9QLMD
aaPWlcnIZbnjsaXBA0BVBlT5Pdu85ceeXNUQa3+fL3VCdRvKhWCHojqhAnLTX/Nz
g7T+oOG+rb1c8odyuB/yxj9/fVdKoUlhp+VLLu+Ej4jx/mkCM2Gmw4xELTzQbYvi
5OqMiIijm0y/CW8kLEn636G3Oc37IkQbHXOJbdTgw/9a8CwCy6RUZtzP+qRELx6Q
MsbLrG45BfyOUx4p/LlxQoPoM5g0qeaceCTK3Sk4OEItBQ6SD0INegq2tMS3/vGU
ff2TqLBHkn3oIR3dCk7txTjW0qLk1MCOx29ja6K6R+BANL8orSBzIf18YUupShQk
jQ8mUOkSgRzpmETu3eJzdy45/kmUAgYhHTdU+lsQvBkGvwAaAWNiOgvmW3QmPGSE
rztc94x+2hUncU94GEbMHZBdrWVnaglMxui/Tu6LtahfJmsiz/puwRSSPndYrup3
uoZbtxwODVCk6DR4XzVqh7S3jfGopB/9PQuY7SQUCl3e0+qkPWcpuD6eB33l4S2H
JCGcOjPgg9Ob2XSE1NdCSfpddBt/Krxfl9u280CoID2xQZmALQZn7Fs2vEk0q4Cw
BY2n5zA24EaMKRTTizrRROYB7eV3j3+0xOMHvuPyocGYSdKQ+3nJqC9WqqkyODv3
nSoy022vsKH6aJdeL3zqLUP2szY8MfK6/hbQNJqivcAxW3uJ4poUG7nOnIW5wr5M
`protect END_PROTECTED
