`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30jGkUEskR5xH5duO2j52FKvoC9NGDcvrgvbCZVVN0DriFr6ZaqCSCsHGELZZeHl
5PrKknaaJb3l3HXP7qWb61iTt72mc10Z6e6XzvLmZ0bXSX/PhY2fQ35kYCW69hkd
7JCc5vc46ZmJeiCL4nInbrQX6RE8/brARBmBwpMUQrLOp+C+gFeComiGHjrz7hb2
nXYcqhWTR9oi2nVQPIg8fK6h4GuOoAjXKs1NTd1UtTmIp56EMhE2oMl5t9l++8Tu
VC9Fr3CcyAmQ6sWcYkW/fv2+/enEMZC3atH3U5LZr0Ew9KnUb7IAY9VYpYdGV0VC
kAFl3CTwTvVynDiHAKsJUH2QJYqCfocT+ceC+Q0CoqM76aY8yKn8TfuFf86Yw8rP
88ltmX87oIM1cWyXJph38RbZjb0Pc7xPL2uA3dPbUW2LES7yMih1Z24zXugH8qEr
XDYJdoICuOTWAXYmlV4FzRAcx82JUc40GIE/omp/k2dB56kGnFFd/8YiDMixUSF8
Op/35Mm3AcBllItwB2wNonr63koTzoyBYv97ZWhr694uw+2EOzMVqMUwXlEWMaSF
J04GCYfhQ7af5fUI2HsIRJ78CmNrNqH1LRCXBxK8NFbRIsiMWGUeXi0p7b05BFwG
p85I+81ofhRIAIU8Vl7xnBgds2mfDxNI3o05mwhJwsyGALiXbVuydMjwiBpw3Ze0
/mnecSTUBhwDWEGS4fLVKbH7FyktBEjaSxo/PoFuJ3nIto4wlTRSo5Jzn1g5ahPV
pdG1JKnd0oa5X2ouUQOKmjcluMTiPH6JkEputZnbl0Brdv7gn4IW0ECl0jxWQSDy
6aSZWHYZorp7AYkMrLweCtjzas9ANygYy0EbvCRI8wRIXJetCeSwtW6vi4igzy8Y
cImA/LvXgPgww5wvIxgltlYvHrviahh0udIxHHeRdkTQtSNy67x3qAGDW0P6zlDG
zVi0TyNopqEK2Ls3OM6ObG2vxYmgBh76NrIqSkUFlspv35sVqdTEEQdvejQ8IrTM
DPsYftH2as/RVjgX7//zV6I3p4HaJalva9OK/1oiscKr9Y7Y4nSVEY3m1PUOgBct
pMj9UcVj0SbbUt//1iIEmfON90vwJGFje5PnHT+CEQR2sor3tbgPpgVzGvuYMt13
uxTjc55zfTI+dJss35ibXn7CRMA6U6T0M0Om4Z1Np5t5/lx/I33qqTNs3j4ci811
es3cKZcQY1L/q3FLvXH4H2wMjKE+R1EDjd+MGgXMbkqraoDgP2lPBeZY+qU/ZIW/
mId5i5qojENmnKT6Z4P7LrAUrzioe5WcknrCJAe79/pMghicpoua1me5AkFz2ogK
i22q5wGlxKB54APcnFBwTClHfpuMlpROt/CqOzBhpXJ8PZVx385RqezQMEGEG/qW
2T0SeCxRaZMumdfLHGxlyxuHLWJjv5RJhXDvmdTvouJGFqAIPqJKLkkm71XWjZ0W
kpFZY9Zh84HMf6SUGR7rhQATBeQACcrjxcSz7OqxA6sM2XTDt4vMuKGJgTviLaXG
b5w4sPOWf5VSsFZMirjEhXZzGq4BLkzMXC514PNVvhu0VZ5OO7OYpVk8oyssR+Kl
LDu/Cf8XUmHrplX9PrK3qb9jDVwG1fYaqsJf4qOF14VKU0eJqwsr6Qyo9h2udkqG
vhqtIJmD/hP6D+FHsSDCUAbVfzlcPPXCCGuHjpNSKiAT6HSZYE4JGSLv92MUGGAL
5wo/At+Kg00CTIDAZ9O9gEaFqD8yvBG4tlafXWddWe9pS2xsufPPfNqcKZy7dZWm
plnaxpB5EEvN1+il4lySurX8pz1CHOjbYHMF52MRy2DIf/MygIQ+a2xRowVJ1RkX
eA39KVgoYHizLVv9OsO4Snx4zFDMX2De3IKGcCL7jVHoSiIFxQTzn9Qv+oTZUDBt
6b2pV9UqA3alCur348DZ8nY+XpDoCQNeF6w7c20H/w49mHVUl/c+6bqD0WXQtvgx
nIGjYGIPh89QDzxAoUq3VQaNZPA+64v3vQJMsK4JPyi/JFRhXGi44xiA8OmuFaeS
tCZz5G+9gmitkgPgKuBXdwKrTBIDa+ck9qlX0BBttWLwvJsQsePp0HS7HrVVDLPm
E4xqktvNLuQzKgiFdctsW3Ii0USgSIrlMM5KwsIod8UN30Hk8betUTcna9In5TBV
Hr63LGeBakSVZhj7cuiWFCJGhKZRrvsng2qF4cR6s6rDlUFbnG2jeinRsb9Up60c
0X5nb4Y+7YaYbc+7nRnvgA5hWeT3rwATFhTzRQR+LbOEApPNbDTqpA6ARG1RnzUO
ID5smMGuUHP7KzmjVQA1I/ONiuWgWFuxYUgMuMrmJfJrNcywO8mqjN4V6dcsx318
0gfbZRRAy8YtGjwPZAalcRaVScZwCfeVpJfRtbJKIRioXccMJKTqxy2QARtuO/zT
iI76SZN4TXysXKHQ93xiZwCW7jAiPElShWwsUwt4Qg33Bzf1QEw+GSc7f2Qft95G
pwbDwECJI5cBItpakjcCC+Q1MoGqihkit0/tVPq/sUWgdUuSSCwfWhx231qVAb3t
uNdPyRPPuip5HNkfrw3iUk8sQgXh1PooXGSkJlerhccpJsTR83//yUW3VBR7NU6g
ov16DW6zUFDGpfLmQCKyHoSl76WgmR2NoIaZcP4EQL1riqMJKxbPbL2bgCBtKb8L
vFwQf3/rhjgk2WZtw0wX39cJaKp7jjmJneCCvbY8cyBcRAmvaSGmjRD3cuKywM1d
3wS2xtOqVDuzE7hp7z+bvIbqCSHBKCaFXmfD/2o/YxrNVcKBQIlNEWbkmoivVdUq
HeJVrUCm8YT5zWvVkiqv2ZcxGRZOYf5LVsef/bY9IoXg1C1tr8cxu4q3Z2y7Nb2e
/uOu8iSWLWufve5eGhLTcnPvtfaTUzkz/Ssz8H+6Zco=
`protect END_PROTECTED
