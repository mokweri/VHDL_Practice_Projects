`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhwtFrrOkRZpdVTp+Si62hFugcyO+JiUEBKIecajMzACZV2PMGt/5luiFn/Nc8xn
Uh+UdfCu/Zd2EqZAbB5VSyINearqxytb9fYpoT8ro2+OHbXsrGUwtjhL8ZnAUn4+
LxPVYrXLlsN+XPV7hQuRIp0YCIsnVSFnVZB+CV0Lari224vPcpvepuucAUM84H3U
QNRoh/ltcXivfzweY+akq8oQyKoYRI9WQYre3meIbUCS1sX8upFCqjx0fqUWEko6
thndUXjdBKBhGzgFFxBYJyEqmfWvTCDtZwJi2tvpqo2XNRDf/O74HPQV4PRmp79H
Lzcl08TWZmdnM9CrC0zsrLd9YYWthDzeIaOPOWeoH2yl783wb6d4o3NF8J/J0Mkd
MPK74kguLTJw472lAJvFqgu1e9x9yf0g5rRpWd9GP/Y+eTdIdrbCP7mxSQ+sU6E4
uV6YBJU5EEqrMYiefJESCjMqV9CttOW3E2r4UBZPnTyrXjynQuS9b8wsP68/HlSA
c+e0zXDqeguFNM0nIGX0wgLhoZRTbzui9kjzxZTYmfGvygPNfNvjSALSWJyQi32u
twKYhaaqX8SPkIz0OJEPgkiW2x2zZwrG7y6RhImPJXk2QLJMq4Fk8+5oH8QevnvI
Fmk88qIxPnhUILKCDz3a0VuUQkEo1f1LCWEsSN8Q+1ZK7dW0KWXnUXdskReLAS4X
0LhnhCrQ1dlpM2i3fiuj5uT7ijZXoQBNBlyoXbwoQ+TVYAygUU9E5u1RY3mQZLr6
0AmHOpbDISaJsv1g4hUdqtKhXnPdu2F647sld0fYKs1bqtBNDAENDY93A25OPnuT
oHRB+TKen6Ey1BaXkqLa3AG+vuqllVyIXJXesJc26FgC/DG7DtoF0na6xyiONFeD
B4vXtHbBjE6hHmsoYvZOSM56B1JUWUuOaVY1GUr4DueHLFvyRnS4mJUfRXUsNsIL
IfhGF9Hkv/q8epoW4o7eiljpGlU18y1aw40/Tt5vyV/ti2ZxW/MdKrM+mig1sC8T
av1+CoZl9xgDbVV+MX6IlB7rhzVQPRHkK9DRj6BJhuw6VvwJmgxFYov14datgUWR
hWpglkyh6ybEt13RcsF31ET2Jc9u3RSw9o8Hlr61eDyS+u4c8TygOhtVc7fhz+BB
2TLeBdkzQairEaccipAbXKhectPcJDkmwsx9w5Y7AvV3DjsyKGPet10McV+eteBO
BpudAQeJJtbn6mQ+u8xAQWyINVMQAWV9KU73rT//btcOAoBaLa5uNXN55jLvbBj3
23DJZrQTVSsUeZxatEXnRYOgIf37Jw0yCzfOfmNM+8Fzi8euMFqaS0MhshvMwUVC
RBCqd563+8pMshZKbKufNBwjzxZndGulDBdDj4eSYXgzF8kYC7FAzQekoqw8DuPS
mWiYR5ox00uYwnbkcvnagA==
`protect END_PROTECTED
