`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qB2faye6eGA0b7sQOQVKfGc4nhqugKpG0rWsIDJ+YpADRcokoiIiFjMfJjMhO6CP
6b03D35X0jRNc3JnuHlaJxUrS9vZROv6mMDBkHPB+McNbF2xBj2Xc4P8oTZuUJaO
BUD4x68zHxgKSaoNuMt3K9xomqKhkcUIrKAtfVISa3Wo5brrBLKUpG974pWXgmzG
fx+Km3nSL1ZY2b4DROPNwZ50KHpAmWQRcR/ws4yyLkFvm7v6VV9r14757TGmdciL
DBX8hup9ltvCh4o2ZZ8AMuSe0+y2DovIvPHhkl6l7MvsyqbXc7IXqjhI60j6c1qc
orTiM5f/+yGql4MicPzPlrLyxh8sDNU3lf5MP4iQdfWdG/ktWp2Ycw2z46bi+wn5
vnfGsSeDMoRmpNjZE/8+fOVhMAp7zk6VcE619kcJnM3RATfNNOFlrqGRgJcO2RNt
5j2/SO/63XCmWhB4k4hcx/s5Kv+vNgZdgEecms3iUn1f6S86sa0f54k4yBfLkXet
kGPB7K1pqkcRXw7/l92OoWkL1OR/uvVgSfAlaWgnD88I0ZUdliivi3FBwhfm78F5
5xo4AquwTWyWtHJtAVghjSZWpu+LdBhM8Mq2kod4jZapY0z0ACR7rJY9lQP9a2VA
agaJqz8qJLU7swPqvCYr1f1f2g6Kyz5r4GY9GqFDk/qL1/M48yVVJxTO7hC2eV4Z
LThX+gjblLT2A1rJr/gniZUrJBcT+r+r50uQwT4KtjhRFCHhlAUr4wvIsmLSqwPV
RNUjy8ohv5TcItAq/nbcqEabVMylrKzxF0F4X6w2bTVLA6s3gdQxxPVbEcHxrC8J
9CyYZZemLRtIPzKYRVyQ96/Jbo7sU0r1mrlLcVi4Js1O3wsmbyX5w758J49ed8zT
8RtM6iwYLs5ZADH6sswzfht6hsxu4SmUZm3+XTsa71XjBTUcW49BxGSBZcrAUE75
1haJBs9axd7wPhtkyewi/VvRASVd13qXjPzuqhIDTkQ4Cxor7FoAr3VOYm/vHGVf
PGv3IY6JfXHLm7LQgsQZBQR8hdQ3tyReHZLrqMQs5R88ISNKXuKxzVtRelMV9WGy
3boNfSVowO4yipbYF+EXD11gRAzn6rEMWiUEVU3KU749He5Qfy6HOJJg24rjSZvH
pzsx+9iBzRNrmLqMq2EkxmBIWL7Txwi84eDwpw11Fl38+MMk0cj6jT/KufO/7/BS
pQtV8BXyYweMv7RkLCZuxRmywgnoKTDcbU815m20L6Y75fphLgYBqrx/QbhZmzve
Clq0pRbcCKOhNEj6mmaiejG6+RknoXUnMFyC+3LksuJmE9PKG/ViQNhYdIxWOV2O
nVGC+n1fFEeZujLw6xBR9VZXHAqPJJED6Erra7xIx/Gs6GID2RaXRZp5d0sobr3w
uGMXMDjod0UTm8/o0i2EoDwQdN5sTvDsrHBtTYdq0ECIVOYyoc+rlBtwrM837Yhl
qCe5hljjdozvPOc3JfuPRYc7iJ/k8XZfACcM/CFOQrIVRf7DEhXQHbljKHjibnNL
Uz/pGPC+VV0S7zAqYm6Wuffcv8+OKU8phmlAzu8axT+57Uh9pE13sMdygSwgv8dN
8q7bITW54Xgbvz0SaKdZG93KjJrZE31ni82pAblmKALpZV5T7fr/vhCYAPfd2uyk
YAqtotEbeWqH5PDlGIf0EX2f8Cd+j7KLxvQj61shZGxNfsNXA2p6zC0e5KoVE3Jn
YjpHpDeQUrAXI4eP/8ghbuE304typ3pPNi5h+Jt1wixycn9wBhJaUDEjg4+3KAAX
7CAc9upMwmgqvofypVJWdbY/IoXDeUID9gavD/GY1YjlV99uQDWTXZlM6JGakGx7
SwUesNUH6qkwVaY8TWshMpDtCgFgGg3A1IMwtbdnqufTEIogH3/6UT08TI/XMw/L
vEsBdLjSFGzHDcFX3l0i8nHQEl39s5bYzDjWBE0aABqk/GFxs620v/H9BeGTT+eI
aGubSAoCQ7lKhHiDAsHxWkJKKvg/hekWqUk3ejpHplYZMG9wcGjRKyuKLW+Mj7rD
yeUyF9iDvjGMOzl83Ic44w5UjD1GK1lYnxReRhvqnROhU0RvLeQPLii4lAGDBr3a
HADRMvVtXJ9+GwA32fY/guJ3QzaI1BexQohix1P3VvUsyjEkztd3kHj34Prr8Alf
TJSl4rNcON1Zjq8qpPbqRbR9IkIxoc+LObZ5yn1mPwW5in4DlzyuTLHfbFFNMIgM
0BdPXc2DMBTermtme4GZ97FhzkEDIOaH2UtMlrzpd7YEvYNwLQcbH9dlY3cJCI0t
lLJ2B6DPLMtjpB+yD25k/fE3BKrBdZ65+dtjDVIcRtBJQX3Ky0JSsx/nvAUtOrw8
T9SJ/worK+RQphCbbgIbKNeoUsqtlDODzePVkmamADNSb9BJvra9KEZddj0aE+qt
8Ithey7NsJW/iOfXt4WSlnavDd5ZBCu7theTWg4iV041oyDeTKm4z/7+vuFON/sR
0kXOtZ3/SQpQ8QJjyt2BrJKYCjFMpW3bNTWxp05Mk/oyprDiSEs9MtkzBlbiO3AL
vpV9K60oWcCOwp3f5ZxH3BxBJexiecaVKUmGpItEFdlmxJfW2d3MhtZ97RSSZ5ff
LGm1CKluxryIFTasZhmFcdG5PV9dgLOH2DJRJktGEHL+IA1hd8DWS9wW03vrhk5P
BFpVnxywuW5KEhYREThOYMOjkdgUZnWuZxpOxnqeSJKeFvICdQsBVuYSJ09AhPYP
WCyUCAkYaEa6o3jnxRvzvN13JZOBQr5WYWO0Xz6oY2shgUeCoIxRvoJJGiIXzRQ4
/E3efjpejSeK0a4pmMBv40Q+9no94eE7WqKFPynxYdwSwJ5ZiJQFlDK6lH+bRlL9
FFo/vG6ma9WD23RIBAcN16G6XcHyQpx0fVCaCdXWZguVgfg3F+3nSdBG8ULz+oCH
tOHkDgqoJMKfWKr6lR/lqrjoGhQxHQy6ADlDCItNmm1IVBdBbILjdFS28wUOT2fj
ptf4o9S1TYn9OFzLeUkpJYM3xchy9+8NIx+2/RT+IyLurj2fG7ftiVSDfqAbAL9B
mGIZ1zHI76x7ZhzUhoiz9/3UUKtBmgKIdfAuNG+DpBmViaSkJxhi2NNdNHUHiQ3G
ZpleWrrIgsPp2Bxlj3NHLPkMClTVUVN/UKwShV7BT/Za9mXwR346ClRm6DnsR30S
OcQiTW6saQI5e3xnBKesyX0tMiP2Umb51ziRdNCcV97yDtf2A7yMFb1YtGIc98wy
DYJf5SrKR8wO/FglJFm+o8AGsXTA9k9D93B8I+G7l61wJqr/AODIqjGSxrFJAQ+A
NgmWJ9BD0Gd4l5XiODjIAg==
`protect END_PROTECTED
