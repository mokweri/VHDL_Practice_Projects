`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qr4u6dSixWx2vZvFDskUbIRbthKPn1Og6HPvDVEDY4QaraY4a4z5mmWVN6plUPDQ
ZocmI+8yp8a2ak5/+b/3gcwHQe7g3n2vu+aekgdlS0TaRNmE8k+s6SwILSBL3CaU
scxyz3C1przgacCksAsYXrGNJipV/ED6XT2wtduaYU+9SMPDw9tS9Ic2iP3YEYyR
v6u5lNqaZgyGZV31K0TQQQUvjD4U3DJSsu+qF7XcbDxtOG3EV/2TEkk4t5FrTa0C
S9fcvjxu2yCiYgO5wgKTmWNwIQalP39NtBTg7LtGUymICDSo7eKemrwnbvTKtoot
L2WYZvWhtSldl6rBwfKd9BaHUG+n2SXXFb9/qrC+Kke+cJQ4rjYG6wQJgMzp6BxZ
LqqKStqCwrQsSRynsinIrgiOn6ylG/URuF4Gfjgix427zkwIeGA9Uj5L61zcRis2
OgDNJ0Py8VvOGWbDRC+ROqn85mp450F0HaaPe1x4NhslrTHZVylGOdUDf/PsJpJF
5dCsYXYvKG03nkwtIuYsA/+Utx4QkN5WjR9UPHHSvcGREjyd7oQlGC8NAaYWltiL
q/HAjO1Li6IL3VWWEudbvViYXvsukD4UEVIp04RNve6zT7oniuS228Imnr9LaWjV
FLN+teZ6x7xPv2DeTG4SWsGQ7uWtPvmbHptlEsZfA/KmiI0qSc7Uat4leEUgE8eS
C+6zudZSbbXk2KntWeHTE3s29pb72Z2C7X520xUK3zxUzlqZmYZIy9zLn4Vj7CkY
Qm8r+Ghj+x3LDFHYa1yHGfZ7OuLMeix0o2jn3Q9hvcV2JZD/bg4f3x03wO3Jgv/g
KcIwNFx1FrnPfU7JIOWsVh5bL+XyY+b9gbSwAs2+3E1fDEGGovjPGJvGqtVNHYdO
+NYzh7nUkB1ojq5j/z+QaVnHSg0vUGHSF80A4DVKEP0CKos0P7MqmN1c2AhKuYLz
cOx8hsNpBFXiqP4ARK4cHb3Oo0maKa7RHEqRRMfduhnZhWcAyXGZo6l2e56uTon/
Tx+AmwnFZy/2dx8BmsQyRboY9sWdXMB2wjZMwnHfXkKqwrXu6n+ZKToXU0A0f5Dv
UZpKW1v/q74Yy7ic8jDpP93oPtEgEVLdomUUPg0e4d/+pCqgDJ7QXXEcnN8YDqj8
zFg4EvmZTNfclJDtBwRcuEMk1+vz7E+/U4dFEIasNFsjXCJi6XM0fZB5fRr90dJO
MEgkJo+sr3ul77saE571rboJtZi80X0060GfGBWpc2BO6kF6zJlCfqf9Nplod6ty
H6EW2IEg+YvbO47P4YmSJ7o1K5OAixecqjGa/+qrux6byxDGLe656AZVOpAIStbi
G72WT7FUv0Jwe716qUxp2IWmKf1NWMpqTzDGqhsb1PeoBiZP/n1Lc0VNS4FAs2Au
`protect END_PROTECTED
