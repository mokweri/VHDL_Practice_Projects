`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPhxOzeDDmIOgx/mwTmQ46x4H40VEVZL9RwmjNzzkx0Y3zk8HRDGcfj4vqHpnBkv
VH/xBVcJkusVWYTsXLI6mmVbtmafB0KCmOOMmvfIECeASayMFbUAFBZlPkvNdTkv
/JDOdAoryKjmhhWF9aTlyYYz7lLR7yTqkqGiP5Qrr18BGnyc7Hi+skpcXy4a55XR
YYmSwG4UXXxDojSqZYLQ31AoRsSGkKurTOBYeTQ2RaXoiq2cjkJTwoVFNKfzLHn3
5qdP+8yHpPJRw512lfd8Y1xWl+UwKI7Cwipq1qXzTsNXd3aVbYSN3261C9ScX/jT
gXaH3sze7el8KMqSr5eQ/JOsTqiDtLZc7LVm/kxM9x+WG+m28GlgmsJyS4XfMd6I
E+fP2PMOAOv1h02M7zMHvJkT2qYqmdh+uY0r8PhBjCNoj5+fbpt7Kctf6CCbesv/
HQJpSJXNzZrJQwvKH3s7BikkxHSUgKfZ8yFDX9gFL4FPiXC4H5yn07SYE13xwuN+
gD+txD6ej2e0gZd4MBOS0OiYHRWenujNtoa/mFcVq/pWDmwgQverV+NAR5/Zzp2g
2sazvO+zEtJVtoqQQ5JRT5vQDqy7s45+PsfGvisT6+m5m9Edndc4cIJwdihmoM4e
EjDJIIGzAJ49LPTdJJ4QgmntcJ0wF7Nx7/SRgRc8ORgyo3c/0ljx8C9J3kGAdWiX
0zdVV42a+jDS72sN8EUOmCzQ9eTewel1o8oucnEcTPUqcSO/+p3oel8O9MwTHQtW
kYF1VDl4zbFyV3TQMpC5DnUB5bsIvuU3cOYXE0Vc2ZHTd2A14MKSRZ+ZmeiYrxfX
BIJvdXb07q9cjBzVjfSOvA+2oM2lHG6ctY/aIi7n5FE=
`protect END_PROTECTED
