`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2GKhdGGvRzCX9v8INLiWPSJK27Pecgjyued4FhUI6cuMXcwP3VxuUwZ0QseBCG0
ZJjfpgibs6gdsBDBV5ndwGumx9NZdujEJ0dK6mIZ3je0n5x/gKGbXbtc94//ENYC
+9Hqnd4qi5V6g0ooFXKB06nCGWjkbuqT5ZDr91xGazmFLVrPLm41ODpQhB1HLDbo
erOCBJ91VF70ZwJ2nfvfpEhL85Pk8gRuIxFk95uq1AALkMBFZzXSvL5uUIxyLPDb
Mkb+XZcVk2pPzzilxIE2rmWJOIn0qtIGN8/LSALrp5geyJZ6fus7GKsGNfenQ23l
n23Q12tC8ir71GSV4jTE54dtx45l2GGQtd8dJd2AoHeeRmN/5oKrPcbF/iLbWWHx
T3f1ve6jZTZ9vH3brImIFT165EG/Mb4xY2oZx6SV7SYlAIFKQ7JcbBvP3G6xPyYX
8vroVhrd4MIDTUxdusUU8/A4Xqk65rLArzrcl9eKKKul3X9Mh8IUCY2E7zBJQzAB
Gb6Z30jDoSU4yo9i4z2rRaAHG+35cn/GnGHS0egkIcva9Q4uQn8p8k1BKJlGrHD+
Ng723OYXr4muzcF2xDny7+f1eLUMKUEHBmZsCEXX4cCSHsaTOyx/Z8ZnYXTSUIQM
ORP2AKVOUvDGEKvrHaMVIJv+1D7uv3K6EtQHjYx4CBZ24FGwElb8F1nh93t15EVO
rDFFS7xH+qvr/pcqsaX9wlmaGZQdkb/o+RerBEfwFtdnyp9rxSkokM8zRWMZzeH0
/mx6nC4dssm7WdsI12ucYR6tenVNZk9ykVT0hr6/MCtpELeiAL5HANvx22HRriGi
gMFcPQSQ+hm4ONa5LxlCV7+Pa9U0iDzH+/+XjASC3zCLBAst5Q9XNuATUAoYv/xx
aGSCzUjiuXL3TA5Ibxo59uVUzbPxoMU/mZdwjeq14dENlQq846IwpxjYuay6+p+A
`protect END_PROTECTED
