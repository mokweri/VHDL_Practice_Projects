`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yn50TaagPQ4Wt7BaMKVVt3RETMtyPf4A+iirRJEwl8cicVWDJtHNtkDzNHPr7zVn
qpISkzf1bSc2e21jVvJz5SnjS2mPlzzw6x4ip/yWqshn54ZhwQLJGM7Gmunespn0
pxhu0XBXb1hvaakzNmg6dY7cnUXm86cpMFCaeCMD/2NJ3jk6c0fTiyC4hjCMy5hS
JEsBNAMCc62YVpR9vi8VzYBCJpQ5/iiNT7wDwQrPpe+2viH3nH37xNvoQwt0cbHv
1xzADK4F0Jfl4kblCKA+qmxaLo4Mli9LyBJYLKItXf5nEeWTf5pHoBmnAzFe/FHD
x6XI9cH3PO4NDXpvMM3JzxMm3wVjjViyHJO/PeNqX/zhamh/mRYw0PTULXVfnD6W
gdp2cJRdpqQvhoHdbae9+uEEpeLmlM8O1bYBw8Qww2FFEU034U1hH7DBWKApHzkC
5hYIZndBVhKHfuf3e6xWS6SH2Zr7Z1g9er+UwL9swYscnbqYAFPVr+mxiUCSXQPZ
mk9CXgWeKrZPNhP6fvl9YQ+8ZOUyLMym2xkupXVnPcGp7sbRxMsm9YD6FvyeW8NE
WoQ0AMOP7GrnhT8aJQmrHL0Dl9nX0AVgfbr3uLw7eskQjLpdPKtzBnsthocGy3IH
+th7gCILkOwKQs0738/UmECPWFcOMTmlI41yzyjoL2Vrwg5n3FXBx0nacWEp8eXt
h3TfKxTu4VtNhKMvfNvTR935uXl/Im2vpV8eYuiJmT0lp3QfCDKtIpJTUppg2M6C
hCJowAZkRdwfn4t7r1oHX7ou6z46rmOg0g+l3LCJEMqu98bI+hGepDv06U1r675e
Hz8LmoyBd7gukV63tQuWVmb/+6OLwv2Ry9DFxH39DAK9wzpEoVFsV/SG3hCf5LND
iTMJCTYdQh1W0nm4IhgmrueI1BGtLS1uIRzJXaHOs1YKzQfMQEOVcIW9NcBTy5n4
a/LWHF6R36BzERJSL1AR1UxZ3wfAMsIisYViNUgPfH6z0oAX63/w0a/wyH7KFbhd
6EEg31iUVpzb2PvRue4hUu2CKgBJ+B2KbeSS65W5/iPmwytYuBK2g8JZoUTZpBVc
+2jhRHSmfJiP7c7z6n/qKUCbz+5oM/kF8mfpyXbkYPJKoIzI0VmI73UAlS1iC73q
obrqn+Hs25aQzQtiETDgPTO2iUjgkIfXcEc+kDbPXTRiEi0LQdTIwRvfD0DbyZFr
oWaSAvOgDle1BIJ/emjw/mE602IDZ93NZfSz9Po4zkGQcchE+HKK2JZ+2S6JQNyq
Dw6nXOP0gpKpuPsAzZRZmDKRbeSeKL1CX8DoPYKyioCEwIjDSZEGAB+GanRAghC7
M8MW6rMXz6T1Q3o/GIdy0YnURhO44o5sK/+V4oMWNou+6kUcLxWQ5wllYiG+rb4g
x7gzFoxraMOlnhLAPdYPd8jHWoBcTgXlJ4gRGfKSDt+Om0D+L5Sfz2WZVOaWkFH8
9HPhlHAlJEG8DNgWSGhrs1zb6aFapivPReZGhSw4p38ikZnNLZBQyMo+m7q6GMGJ
q6ESzChLplP4NCZBFfxQyg==
`protect END_PROTECTED
