`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cgZ5GBvs51A5oztlpamHt+Z4tLF9k2OPBi4cqhNC65zkjbS/fN8DuMS1SC5tq452
/ZQKF3R5GUCN+CCWkUqX/hy/PsPvfCIPU3nN4qeDQFSAQL8CBVKo9V7kBO0XBN+d
7Ma0oqnuayzbLi9J9b3Jtd5UaJEzUM0sSb+EPtSujZ6WbX9LCgWI1+1ggnda9EEp
cjiXJVVvUqhd3iTEqUTZm3Mo8K/BzEGKoZc53voJ2JiYYLigH3NSkW9aFT/BJs5b
2LN1XR4KxINVavwRRucnrugVjX21ZdAXsfg/wJaZUGZ8TQR2H61/mvXT7S5R+8gW
tNkjye/ey29SSarFk37gZLPJh3J7zsJ6zn6jMRrchtv8+oBZqkxBP27Mt8HfteQw
FNxLWMMZcbkFKH3Gp3XYIruo/PzMPEhBuMxlb+XVPmICgio9qDZlzdDfdbr+XKDg
MKPIzJ7idtxPSlYsSbd9yourKQJAvDGOJDfwoDxrQRa+hdUfWYSYOiQmhGWmUAMs
giV8Nu2sJj5HbX5T55HohjEZRD4Hp1CCBhL5dBaJwAkK5L7edPTVytoy7sEdZuhA
uktm8igARlL8qmCiEtwmJ7AQMNe+UXq+7rn1cTAKgayyOzY2ym64HzRNB3TRQ0/R
+OLl3NgyIhhy4Qw9c/RO6ceTqhiOyHZ9RzYwMSNN2UDUBG7jsBF/byuJQ9abg6dK
o8FXpopV5wLgyAcvWkejAo8ud+z9eBzSi6pg3hKLL/fBHLXX8gR2zkDsPbGBNCRJ
kfVwlJDkDnA6THQm8lqVVjaXIEU1Mykk3FdYA6d4MIuqwgqr+bEtsBVtjz1a9wFF
l3aETNzB89H4LP+RU3o3CKhL0+hdUmV86d9FUDf0hzyyA9QovWe/97NsmFdJftad
OhvC/d1yb56F44BXsfNX8bSdAgHO1t2468Yhg25ISXVDNtx3vG3o26nwn7KsguPc
sdQim1xxrmB6IAZe5EDR44EOpVyj5ykDdF8Mipv8KiFx7pHlmfejng+MIYka7bil
9Y8Ob9aIYJMxyEUeQkZGIjXVuEaGk1WAc1kqs1Z5efp0oRhKgRG/YN5rLlYs8pI0
Avxh48sEh2j9vzqImYCJdxCmNtlfOc1OGwqq9bLEZVvsuqwRHUEh4Fp6jAg4WCM4
gqgj+vLy6fZn635slyZV+lOLSkvz96woSe8IOJzfzn8wfXwLGuKt6D9MxZktAFmA
giTWkzC+VJQ3Wbqc2mW/4wJYQ6wHqWbbnCyMBXt0DI1sSWSP9/cpXM+hb49IA6oJ
i+LU2i40ytIpyhuRGDTAiDKOQj+p2Nh0kTEdZzqkqn72aM3aVrW5/ghk6Taiz4hH
v4w0KBtqrfZJehAttnS8K5tvYSA9ibg+ond6IISYt3yZlEn6DXL7b+tFwG+hykvA
hZp9edGwFNSRvCbxZIGlj8P73xXeJDLYMR8B1TAehXcSM5uBRdY8fTxqz0K9PPGe
O/uJUayztQj1wAydojnJybe+rkPbnUMDwEe7h/tUfkBECK6GVK0Br7fwR0cUlMgz
PL6s9DCbJfUyw3N5bmKgTnls9IMb3aDh0iTGOR0DSWIzmCNJfxfcKhjHUd5zsjd9
KOBgAsksiMfOq0bcyvybVdb8sYN0f5HfHnsiq1Ay3v4X7M7GWzC/sM6E0iXzPHca
s2jMtnWoLM/N2vlWTiAm+RhJH2nzILkWsBgCRjzi3YryyNVPcTH4fuaKHtMryMaS
C8ja8kEE3o8sQwZcc/JrOZP7n7R/DwFY43k6C++rlbD1Vskgf5TnZ0enMoZs7ZwU
xF1Cuu13jFdnzs5iJ8BhjD0L0kH8Ht8xJxl/WSH4uErZPHdAdDgcFMYVm0+vgUcq
OEav0mZs1pytyOPj9hahq51dTF4ZGIiLrnTnVLNYckyAim7qEbVj4c4rMd0pII8A
dd7LzPjHZtyZqMVSCIGNrFh4nZmpw0fBuH4RlCpdBIE19bmK8P3PWkUsnDOeEjNr
FVqzuuVOYOT5bF1vUDJvPeuEw7+U6M2UFJU/qpwOM0ESf9bT0TuIz4HDkY4SxDRZ
kddm/Bu9rV2mYxL7kuaFp/gWvGxSiybYKNSEF9enYJ3yJYMGJc/k0ETDs9KxIxOL
Q4UMJDq68K2APJglcWyZInoio8qNi28DCmSlS8cf6+EyPIsthAbBmWaZuunyyEjw
32d7brzRND7/zSWQ2qRxPHNv+tOx5s3lE0Of6BbhVp5DP4nFTNaEJqroji1mC3Qb
N29TThtDcrOLFaskVho3ov73eFiSOCtVhuRGeHiScj2CKGK8njAfsA/cOd9MY4Aa
nurzUlw/zcBGneJQqC6+A4Xr6APLywSk1TQiJQ/sdlTMhglp4HvesFLuUxoDp+y8
jSpwZNX6KdeJ6BTrPM2M/dN00d7J+4IsGjYJJpDhTrdxcQWBXO1PLoGc1FrlcDNW
hqaLq3BwHXhj0Ndlb59uE/FiTJnMbUw/AyDvLzbELDpGZ22unUOpbQMUyjCD3RwI
xelG/jTXdUmQzn1Ji65OYOsATYiM31+pomcecz9aGkwJB7ox91OtQDwnvn1EcuiR
911vOA6fh5iCbz4/9M3V0fNS9kTnVXFalRd66JKVx55VIFl8XWJbW7IF5HofDKTC
lZoDuQgU0cJHMteIWy0yPTplNTeZ2aaB9I8rzdXKU5E/ri/fFY5helV2kU3i6JIB
Zb6PyIGZgUMnrr9gvK0b3HUnFTgIv15Fkfxj0tMP2vtODb9mGFRtowyoYCIEjFeP
I+A4tnolrT/dnO/16y+lBd21HOVN1JpEqzyunjs6wgTH/9PqJoNpMkbEoYlwjudI
hcfbP3jsqnoisD5Ap3+ICNmsNod61NOeBZh7Iif0cBvoZA+B7cQ3iHiR6VBH6tHu
COlhE8QRPB1/xc6xHc7i7cIiwPdDMxn1VxZHLDepyhQPtjsBA6yMy7MRPFQzt9bd
+JzZ6xBmnbIJccPjw1ei5GBdShdrwVbJCWr7rVIRKSlTI0RhzxGoiccdXYkO/Dgf
S6m08K+mrmsLMZn2mbDf9EM4M0nDDAruutGmPoboCw8rRYMKxGseBy5showyG7wp
rVmuMKiQSBPa3zvcMoYvpbp6R0PnyW1FL37UUHSX0vvKmHvVI+W5IvnuF19yLvRb
Ra9X/dy8pfxmbohJMFeQJipj3AlyVKzUijNAb3Z4dwYQUw07/4DcA1GWo5eE0JMG
97ETEejdNvc2k3lgk4ZuhfWI0hX0PdKricMGIjXdiyz3INSoIzUH8gnz7NAK/DoU
wd8i6UcHtVknrCaAxSk2Gda+8+noGCAYMh8D2ZmRk+66FOfaKZL5btOSf359sO9e
i1HbyaerQWqV7jXk9JveoyqshTjqXDVQvcOnXj+sxG0ejf1NeZicZ2b1q3E/DJVB
5RM52SbHs/QwxYAJXlj+ZF3rvTPEXWc09FHHWrT0pYRIHA3va/+5trYi1l7VXKOq
7QrraKkAFybdgigxSkJGytV1GDLbHHmLRt+CQJk4ZS24rew7bt1lkSXBrwgDK5h1
s5v4CqVM4e+B1BTrgCv4VKaPU91Bt9RnxPXkBMhtInxB66p7pg9LwZ1/MqIrVu0y
FBNUl8nDCRqUak+1jbzBltytAOB2xckwD6MBhlxaG7CFIvmwVJ9Y3xTnFDVN/7mA
3yr2einv6PV4XvBTclwPvlHwxOj/flX4WfX2AX56RKBzaTFb0arbgDUDCS+NxclB
MGK+oCkfASEhuZp1F0g5SJ9omamC3beTAHRkZBy4swT82Lv8pVaEVFHBl6w0pfJG
ucQi5UpT1QAgIwZo8s8oKkA7bwoeqrZtRLYE5rstFeccerp0LjIW488Ont7Lp4v+
RvR5JIR/ssS5+G62L8F/+kxdQuXBUzjwnvxa/ZIddZmJoKJ9eld85VBinJaZSJRO
Mfj5KNK9h7IAMCOObyPNdvfPSzOkt62wFFennAzboFR9DExrR4p2TKxiTqIXTNnu
wCHf7YefdeGoWmDY5XMsPKAIzfNjcWvCeeSQX5coEqdOtAGF7Ob6rj6osQIJLb3f
+NhNNDk7ECqohiWTog2eYzNiwFCJqHj9v76VAqI3M7+MnqKkPQDg/gofLBrCT4At
k72gbi9S81rn7X4ZPTEcLBxiZh9x130AQSMi+bkoZLi9e9UM96fbxKznJkZuKZgy
vc7CFF9+/2/lidtsoytEH0K5aXWsAGd5iEihO1+NYvREY01Fg0O84wUCd0E29dbC
fFPqfC6//9w2o+fVdzj03CuJilOfq/m8owILS/yGaKG5FktfsRVXAAmK2umyiL13
AZv8smEAPHJLluw7DUPgv4iUMubrnJQuP3IVR+y4WWuvfGq8chGsZj6W3bLg4cLw
IgfgtDaWec1eRJu5Tu/IUfFmR4UcC/aTnkqQmhEp0goPs3m6MinES1dbfvQhu1FN
ndNDgYYsg3Fwhktchg8RhtVIepPS014O/F2XS+Kw0GlyrqUZQgW9EF31CRofAdq5
DmPNW9WG9FzxwC2TcSukm9G5Rq+mK+S8pEfLOi8wU3XmXNKf0bGUR4fh5T/Y7aiN
pUPX0gzuqiMbxPApPHpKnKZytTs5TLlovbE9o/YfTeUy2iwpw/t+I1Ym5oc+OZ6I
afNOMfRaucGMLlXehzPHC62+RrC8Fvx1wQYuhGTYI+wPstZTVl/mXbhYqFrq9Fj1
KcHPQJ2BwxszFBCF/KDztSOlck6jDv6EdwMCOa6OjmxXkvgYiwjUVZ2FxgGexJZl
RLh8siKEML0+9jCrl/2lOJNoi2Ov6POA5PMoowU9jqHqRxqZ7ofg2OjhYpJRFMIW
zsHpll/UTBL4FIY4YzJCcGZAbc7MNVmfuBSk8lVaCXIjFrjxdD6tpp5KyOI6LEh0
9Cr1fCfBwZKTCKPL9s9ZJbpOKMBfigWfQiZQyO5FM0yrCMGmxY71BzNZFh8jNfJH
CgMt3tFy8xOVj4kpYpsNmPGj1Y4WVP5ZrH6W3owvajb8rsIyKLLgqEYTZQOP6O4/
MUUyeN1ZfSapmDtJjNYXAZqsMENFbhx5VFxEFcIFPafFqdVt5IEnhrsskvNAOvl9
X/2TDiT9QUpLWSHuqksRpBrgT+XqJ707+fNtiRIY9KbtMbmbvRY+cwDpWN0ZQoxY
rea0ehmZz0cIzTYNfEk7BBdjZ0Ga1+DXmVP5ILMT1nQ9nSu3dj3LynbSykB+T3fr
DPKPHhEbUSGVPd2KPqFmxITxMDsUPBNSqzIDJgVEs9cRgCO3TS17r9bf87M9EhA4
ZnuwDQ3nkgJ9AK2cpsLv47PG44shACBwHKLtD+w/C0Xm05UQqGKAv5Sl3dqfNDS/
iDRkOcUqsNJgVGiazn3+9zH7qZyvsdHA1S8T4AshaLLGNOHNORXloxdHSiOZUfix
FmmloGD/qOS3gVkLJVMR2WwTVp+WFhOSLh/KcZ/LMxP9spDzFJUTBYcdXPLvd6Vz
7h5DmdBybqxv8xiljTLlNsNitN1NSfyiwBZkBSjdaPXx1cIqymihb5scw8cbjXV7
tzW5KeQ2niC6RXu7PqHw6TQ3/0ED7DENuLe1mKXYZIyS05rJbSi4iG8JfFuSiUoQ
sxm2WsFaAelz1wO+mojL1XNFfCUMRPTijaD3jOm1PrtvFMbN5oHilaHLvuZejQvi
9NS372BSoULd7sgDg8KuCHqnBeg2FqlqwaLY82hiNdjCm6/C0xkB1yeZ2jYNTtf5
njGAR2EgeUWuKixPbEe8F66QMAMguG5xZvJTE7SjVBe1eKQ52pD8gellV/XERVmw
MPXsOZBIxgmxNz/fI0s2/KekD6J0so2DJzy5pDqzGMrFM6dyTgX/eik31WpkdgWj
J5LbR6KWbSFlTY6PbjsiwMXLkqwBXptbUpZ/6IKl6w6JFn89y220xGz80WwT3kEC
lsxGHPYTV/bjcr2Vy2iwElybMVUO0/Y9XjE/VdT2hBafnMtMwO4DLxIV0rBPQIly
GJtGWlNFajz8s8LSw1jg1WfAa6QIcXlDZk+I17lHGeVHn7uRSDH/ggLDK/pYj3Ax
wdbg/b8M4eLvPq68I8HpVXLwB52bCZiZEInBfPKu7S6xY9RHswUtNq6wfwTvxciI
GzFtc+syG2VEkoUmjKyWWpCG7LbvuiNEewl3a+Cw+KkLCq2Gji5KNHtxCOsa05o0
QGqRynRbPySIo7jCV8jjcRgn5TpobtVnwWStRjuTmiqDHa15MiTHvD7X67/8hXbv
BoyCFTW+8CMenQK60YwechoWHqyL7cvCEuwnlHvydwXW0niiIyk0B/P9Z/xgHs82
1rPRkuI7xzLd2fFSQqJj7ZZGz3yfwAHkWUlpTvpfcn5vo3DvcKY6EikTbwWfQBHP
xjIn4T0vbC7P8MJjRnRN5yM9Bfvl7oENt7W1NF2JdXFqiYbUFoo1VjwzAc8UKzv5
BgiV+mZpaglZqxEKP2BBz291/u02JHm4q3BPfo0fvGULIXH0C9rNYcR9Ve1uYCdJ
0CI9qDsZO0s6yQjrtYB53z36uGQvfK5CVz9sT9QJqf/6NZxbfsONvswAeZy1NA+9
3jeVC5k60F/kp+DkU+ejFAmv7YYQoVE8nlc7VdlB17nmET5IwKS+D/7XQvATKjjG
g1wxCLG7NKzlvSGDzyuNTnxk9sQPWLTUsm+t8l44B6FZhBHA/X9wPmGb7XooHl+B
8AxYYEK/Uf8QIJIUdFQDTj6YQGzABRTu0Y1L0wYkZm0Nq3/C3JhcLdJ3IB5lcXwU
kmcZPpl8j3v1OurQbliSDxpR3TqVhfnahdIuHVNwIdgZdJ/lGfrYtx/iMhUSDwnX
dnblEgS0J2Kvrjn9fpJdH7RLO7lRLUfn3Oqe+wuHcivUQ8NlPdsvwkz4vUwQFj6p
3FZMqwBZb5pzxq9h+udolH4HzOzHsit564BK7wWxq1W2tB4Ph0/s8rq5b3BgbBIo
7Mc5agoy/McaqyOgonM1Vi7B/0Bn02IXMf5O2mCkcl3kKSesR66ltfwts/imcb24
qBQEemFKlAWxeHHpbm+O9OHg1o4PzdWefp3kYZMwLwJf+BqLJ9LvwJKtlwiXXSp6
PQqsmuqFkhbwwUJzrSR1+67Z2BXfQsdYtZpKrh7X2/Qw9cib9BcQcnkm+j85+QMy
DtlYXmKenGoa94o5+Dur4RWbVdtxRqntXfJtopN9ZXPEsw6gbbdd4SlTZdHD/Y2c
3ckbFm5NIAfMNfBrjbL54UEA+aYVSSGXW8hTTrFxmN+z9uNWXDFl6W7jhnup35qR
j9TW6HmMCFbMi+16bQKq2ZY6ekuI5Vr5oc5IGK0bqFIwp2wUQBE3+jANm/soO1zD
I2OfCsEiFn/8CJl71EUzlH/dU7RweCvLmFPO5qFmm6DYm0ALtwXuxsq6ZuByse6h
qsYIuR8rE3W33WWazuG+P6D9U4lZz1eYYNw2NM+Wu7zAGr7K9PqWAiEbBpKkIkxT
YUgG/x8zasbAT0K7PNSIQyhxfDXJx66/eU9GqJT+2wwk2wUDdt92MpPTrK7mTLU2
+6Cs06uVzCv6v66tHNSAfDXqQA+3r6yuHi1+CbHlYJYkpf6tbmtfaEP46XTPx72O
x6rxCOCQAcYL5iQ9jO1Glji7zkGn+32cYkEGvIP+KTK5F7Nov5Il+hRpg52egAu7
znpCUnNN36LisKJUe/BaWI/iVZ8mn/7aCX8FOHzyQ76CWRQ88Ec/hxbL1Ogc0/9X
37SRXhnukpXROYjjP0eebbvSyyNQYjOUpUcgaGp4C386FZcHlZ9rWP+OmttqJLHg
uMJ8C0hMvi1A2a59wyYp/Mwi44FrgAnK3tCvX6T++/LPC1KLjWcfhyj8ocD5WBAv
XKMaLMu59g/G/ilJVqKkfztEtDV6YZyX7WXcR0zfsZu33RW4ujM6wb3MSmwhlWUf
GK+zVcIgLZ2VWDC7qYRRdNTdTH4Amf9FbSGGHGgrPg0Hc4f7ZDc8dM04qQUGDPfm
uWEZU/qZFf5VNkpk1E27BwqRcsdEPlDRbJ5aul0S6MATyQA+nwG9x2qxhtq2Q1+d
DFaP/7HdQ5+gyH9tyWBkQiYLgv/kMODePyGw9h1maZYPzT8KpuBa/v4J7va/IIAL
X4x0obW/eLxPVyaF+2VUFdHYzz7+Nak3ebhtiaVJonet7ZSlbdnOKjT9hf/2SW4x
e1X7iuhN05uay/y2BkpY/WLmxIkmycCKROqslHnRqE4vUNduRqa4kkUE7t9aekpz
V/B/npT0myt3zZpM/7qAQeO0lI04c0jUD307FQeeuFK1JLXv9NWSrOxtVAN2bwAe
d6I4Ks53XPjYh86LQOymldoqQjykf9/diCK8LXJrAhnbmkb1x18fz46xR7NtJx+H
/SP/cdBSXGJefJIpbAa2up2q9R6Il3yAOOD+inm/4HlUt9WuVURyVBNCvwCJ8XeX
sQjSylfy3rJ7PKDf1z+aIuIgst7+vkHgiTA9j4NJaTTkH4Ma2HxIwEznpw7+Oo4A
LhQmFFXTMVx1R2GIjXB5IE3XwOYNZNTVXLmTul7uWv4Mu2RiFiYO8i2LsHLirGuw
T0+fJwWkPQTqe+zyCEg1dcsmk6c6HAOzfl5OMxVJsed6AI9hN6rxNpURGsu9b8m7
JHX6Ko2/NcH97gPoSn6NmAzOepJXmSWotQY/iAU1EG/AB3MYmZzoSKOqSX7bhNna
p/UCc6Nege0yQOL0wv9LTnNqi5s7no0FlEdHQ4fzWGRQreN0FDsuEF4h2rccVGzQ
EGOYJ/x3FmJKhJI/umW+US1auuT+AbExsIttZtNvSyw6EX8X/ULkrB/z3D12PsPT
QmYC3z0o2+Asjs4/SWCjrCZOTtAeWK/8xqxwijivM/G0KxqhMUu4zNFe8lrVGdWs
Wqo/Yxb5QiBh9oLEqJKBVewY/K3NIKXTJvM2+DGc/nYk8tv7TG/M3y6jFsqaOgP1
/xxWcu8hI8cyTMV1SoZE9qKLTzQ/jicQ5d6sh4OwtHTO669Hb8/Ya6ELkjuM6DMX
bmiAswX07yk2nTkYIKeCZ+rvawYlMj6DSV1x78GeYASu0K/ITVlRQLaO/cZg+3uf
oiOvrGj7oUksrsHm774/+ERqRBxKNoyJVr4xhmMOerd3FvlcWQ7QJB2ZhRBtsIB4
oLmgeDi8rRj75+clr/SkHSRzkiTL+6PnZ0CDRgyo2m+T6dqa+EtoSoRYKeA+Qbj8
obInu2cTjYFb0Sv+zTfq26jknnTaM/2xPgpIM/W/D/kSCXzPv/ZPb9GoYtX+Hx23
9tJPI5TkkGAKvAbfkrla7ORVqy0tKIorwgb23Vzsd9gRquoiyR+3hdRqSwQ5imZU
sklF5jOVWB/SJJMuOlN2YlEy/7Syn/5XuRSLQ9BR8NisNK86MrZATMU2Ogm/PR8M
2BmAT9KA0av6nr7ZY1rd8YzqwqROk8QD94XoSL7e/cK3sbaefp3TwGSWMqBWNxJ5
+CMONNqiy6RiJWYrEljtDavH1sn63LzOqobg8VKp2gDDBhVB9eY1sbNY/sE9JNhq
Dkcgpp5u1LfD1KFX9/nVpxCZ1VPOWLX2z8yGxSc/HtAPUWGwKUnWrjGdlTCeVeLq
kJ6WGJW3Je4oiK4lSqUVPGACTEtGZ75pHdZDhShBgJIgknexvkmh8HpedFL+qzkQ
xnTnK7H1skzkaOt1IeyMA8Lka0/udg2Gdqai23MdxaeqLxMW/1qkp43LznKL5bKX
3GgArhj8/pZQZ6TY/Q3IvDbRarCBj2mM0mqPgJukcXn8QApL72Wcv8yjuVN7L5Jg
mHzIHiqJZzi26gf6kvqyANKhXGd81asMe6DbkTp75gDBW8DYpPvG1yjmUpq+Lxc6
z6g5RyR5QVol6PRYlMPpyGP8/Q6/YKcf3XLeteWfCHgUz3F0N5BVr6Qga9nJsh9I
R/AsvOctklw207nEiKo4Jk5AHqMAt/ZXTgl9byIJ6nUn0Ia9oZoa4vao7HvD7xhJ
y/ES6/nWQL9NdKfpmP8HsFqfsda3xAqurh+naeGIOPaf3kN3Rg5z2IUdfOANnxW5
k8WNp3gpAiB1zfDdBpiKlDB2iAMmUBk9SGhxYV43oA6nNJf/jLp7YEXRKj/We1mu
ay+qI6RBeKDbJkqQDL5YT/edL1lS/uib+zBFb2JIpPqZr2yQgeNSQuB54gIX8303
mmk8fds1xy9GG4P8G5Sk3sjpORXepKFgfFER6IeOIfRxJubaW7yHPdyQsXWrzzwq
+tS+59xDp5Ou2fj/J1y4jR6JxU0Cw3xbcRa09jX3rup4DzVrW7ERr9LJuJTMKqEG
h6a1W67zBTEj5ENQxXpmzRlxBaK/omKRkDGMND9Ky95VZpckRoqvPskGs1ANUXdV
osWvshLmW5O93aY8HFeCBbWZ58OTsAGqTYGvT+/CW3MR91OhQgT03s1OWmv8GI1F
T4Q4GQN426/MRbOiqSlDzAYQ3wGiux47DHawJUmcL49L8PO6I7wq7SQRTDNTzVP6
gTinF+G0W24/KpRpWZfdZptb0bizuz7L/kdyfDVAPtT19hku5oQaQjRtqKk45Kl3
xDG19okdTZyOpvM35Byd9ucmUIu2gzQNQTgp2rti4zTrpzQCflf7xhoMeRX01JFO
1EUtDoInZPHrfm5amo9b9PWiv30oQ+1xvtCXJvAWzBdpQPS4I4MH+5oolvcbSmJY
j8tg0gz86ch0OPEZ3Q7FNiMUWXmHNDbG1uweYXg/zphF7wnSAz8mf8JyW+Ctm45T
9LuKmHlI/MEvvTuPCS1MB05uV9PqKI0AZlPlvZowXKfNdO7d9FrCYpv01ZFU0pD1
unF1OHP76Y1qZbjy9z+OrmB4XTFIwGn2frcIRvrMiEOYt1TZJ6dixr4ZlLMSu1LV
2UOnyYzu6bQR4LedSYEyA0Hm9m5nfyMckn2I1mJsqyehL0LxK1zrB2WQoiPeQ4fg
rsFLD49e49nAl/OxcKhHw46WAh4Dc8g8njRie7uuYbY5z89gqxUwh+5GbR3M3wx9
pIagyAUvHG8qXMiT8R1WCmsS/oa4nGEE5cv2gxTblbDIQjVJ7gvk+SEykr1IVG/3
KJjIK8b4NzmoizaKrlii+yO1tvFozrPdNYleUHHgT8euh3Ke9M0IKHY15xg/+WJ5
/IWb3mfOGRrgXasxjSwQnu6+UHxiagb+VF1rN4yg6xOvS/anJPjTtu/P2XAgPoP3
BHVQldtm6HxOB1WnaKXr+DUtLDwhkprspsTbOQddEFrg+ZpcqsGswLkWkzZf10je
SNEsnqwBourFcz4czTdO5aJOSYq6QqBwmg/k+DVgAVe1S1+zgpXv+6KAVHgp8Mq6
ZmEHQX+ZBmdgmnw354avMHplVz2QBWn/q9N5Rvr6Be84pGCxBaIEA8nu6wFV3bZA
l0WQBFrCt55DYrkyVhyw0+zBQ0s/Tmo9WNPnxkOZwyYCVWmmP3+vLIQnwnWrBLAu
B6l1ragjMH9heO88vHrokMSLNu/sa/oNzNNpQX0QdvEEZU3btxTSx17FRD8UVIIw
egg5s+FmddmIG+dtRqWv1yWG2biPr/CSojOR87Rl5OImcgw1+hhwn1AS4ZpY6DZF
BsiLdBkjliS8Uth7U3dE/dtIq62M/uzIqp+jBPFEmpuqmlNDw9URf344mlkdca+n
1IZ5tyhvzstpFu1l7cePjSeUKsbxkg5Xt/fYXBb/7UoexNB4hOogDv1NRfXlC8wb
XwiIlljKd21Xfhc5OYwl824m0SXlyRP9bRXBy+7cOsaViRIxZMis9gOkWJI0//fI
BcoPN0I+ABWlpFokwjrSbPIzRBSaqoh5KZ6iWZpcgjGH4Mi5JKanw24o/DL51vSP
EESTa29Ivqa9StybYBq/OY5mYQfPqRKS1cYduT2YrbR7rApzAy6fC6KFuwrAOgZd
Gsa+zocNwy5GD2YT33/YTnyfKFPRaBn4yQa0k6Z40eS0Fd9r5T/NlAFD+apLFxl5
uXVcZ1BZ0phB3c/rNjxYuRCs/c4LHJUx6lu8bjnB4Ig+IiPfoJy13yo95XmQBRpS
pBaGvMxN0oUSTs3p3mKD3nR/XmFr20aLuZYvCE+vF1z9LIayAmtf/GMlOiroYPnJ
FPgju/QTPA29QmTiS049ug2YgZMZZePhYOTWB2WKC5jLVPX0tg8wu8jBUa1EW9wN
ab6q3JNLaueJ6Gka0r4yvLuYchSP3B22YuNiAhsYpNVf+gDZLpaRo+OtCwYZDzSe
4oO5TXZ7HNzc6o5cb7LtWtvWAuBWJga0LuucLbn89ln/Tl8/r/0RM2cDLgrzwLxM
fbUA8LKxyL2htE5MZJ9Ibau2LTovTzoKidVSgtZvmiPqo4CSMyuvmclvsQ78VQAi
3FvWaLCS8+3dhM8tvem9vUq6NoCHB8UOdYkQkJxyN91TwJsYfwqpiHnx+dPiN0Xe
EpDQTSlbIwjR0sgio2+ko7WJ/2uwugXxgbc8k8Z0pNg4+YNlA1mWVzSPxpG/zcx9
Cl48aTyWD0dLO8HKhs2RAA4i+hsklZ9WgrpZfFuxZsR47g//qGNuUWk+vwCCtYIa
TpXLkqACZ30H/PeOJqzTgxqMoQVagAEfAoDnyY0vbZllxUx41mYbvZsrB0VqAoAl
hmDhtDh6y5dj7Y0wsjFl6pyl2s2MimPBFeDOdR+rcU1PeVS4erAh1qEy+IwznoXI
CuRE71MPZ1m/vAmHmcDxpM43AksVBopJy3dEYFBWsFI1oslMnPGBYchGJX+cFGeV
45sTvoTqq+HzIJbcDJo50JDP95QcMxiP3RUJovarx5xILjDwJIDu7bqUT6fbj6aM
TSB5giJsq6nKfit95vfKqGKIL2/mjnq8KOP50/iUDRMIxvxgSzjLTFa3DTV2NpjQ
ULwFyldQMaQvk5pujuh1uz/boxVKaOcPvxI6V0dc3RpaSuvi6yJ5RhaeV8W8FC/m
OePLioc6QA0K2P/m+BIxLfyIyISjStxJuXolAB2Ly/S6sclZFIpeymUYtm7J5F0I
rb/fCwaZ6vf8jVczJm07SbomXg0ySlKQltY7/tSEG9P7qNlyUFBeeN2rIgmCmUNW
ye+zFq3HF+1+IWIcwtvasaZGc9JTAiuWKpiFjgqbpO7pLgChQA5vn4+nCG8NThMG
M/EYExLegZXOyEWUyaW8g4HAKtERw1ScUnltFGhWNB4iaL986Jc+dolp2TOO3OIT
fIW4H2YC5d9lqap+KVpM5oPA5i5k7h089jZrGv1b2tKIs/Tg3XauV41myw0crVXu
WgiSVGDGHTmvnBumrnXzSwOy1U8mmvZSneX4J+MaZLJZk/VxnBLcx438jjlBu5AJ
TgFhjHwpIm+m8Kc1JCM8O60OWve6Xk6SGCRXAmSjtaXLUMrn0OkmcTMcAqk1To5r
i6UxzrBXL9+EHlh1IShEt5+DLh3f2zroopPpL/EN3lxvXdCsQM1JtiWsx93vqE7M
nwd9XzE1ZvojZnRPV4cC/Memxw8oPEWUyd9bgdhcDS1d0AMpTaYTm3QXn/2bH2Sf
h6MgZae7gq/DXgbik0DhEPEoL0VMzvL14C4mi3Ab4XG431ktLVtsN+oGPLmitEh0
dWs+g/LeW78C4ERZo2h4ZWiKq7NXRuN8DnzmbCKLwpIWqPh7J8L37QNkAwMh8Zuh
FJ2krslESIBpO0y6tp3uJRaSftRLugeucW/rGiHMUzFhoWJkJxZ0fXt2Q/4Qmm1O
Q0op9/9qX+JQ1/8/a7zx8S7SurYgHK1NfQLvP6lqGqghnd+OwtfjY3bFnszRZ5hk
8B91vNr8g9cR8B8FsuXb/ZCcl9EJ1VHjhiXTDRtVaW5vAy/w9Z3W8No5oGzpFO7I
Fmss4b12GH7iSLoiAfQD2QUDu+ZFXkh2C7CjDnblpo7Jj9SbxSYAFkpqYCIl6rUy
gNejXvIv6VKCAQ1N3EBY5+FWM6pZftPO5dbGEgdY1plN84NvF0qIwQFkkh1EIJ3i
pWDz0HKqniX+cKMnL60UgF70Ikr5IGmQ9Vzr4f7z5VdoWuEZpEwx/mIB3tRqd96s
LJwJX8gGekPyUSLZ8LfZR3pT4bINyqmMc2OwuomIxfxR7DyQEsD8J9co/3DgkFCB
vsVn+zxZBGPDgfpEzzC/oz06i+hple1TnYR2tIEIZx/r2aJMKLg7pNvuHGdMi/Z3
7m3LMQxDYigcR3DbRzHIwOky774cg1AHEPQoeOvKmGLEs67qnwoKcHS8cHUuWCY2
38IxtO3GzfJ/xVK4D6fxq/ddr6KLbefgibHWauTVvvHFSZkx3fbQcANqe29+lu1g
rRw41mmJApFdPYje7wHghOYOrZHZixHyN08MCD76BDl8pNUIbXx1hhxLhM+JYflC
twXjZVNL7dtw44IgYiUVB37yrIOt1NlG85F5aL0c/yssl0octQf1wPTK+81qPFbn
1T1bQrp5Ko3Mvy8EBggJGc3TaQyrDaQyGSBIrnqiJY6iy4IifHLeRlVOIJCqpxD/
+69VKSqE3GCCvsb5PnKInFVDe+0MIfY6mBaidBTUzSzmnYGuqB/u8KTfAy++H51a
jCfDGtZyQ9EWq1YJtoDRIttMrBJ/rZVaX9hlVzC7UooH2mQGNLpYRlzkFYeYTsrm
2ov5dXxwqah6ftxeALOs36g5LB+6Q78CED7cwDkFJZ1gb1cZHQ6J5GFM+MUWCAqf
4FSVagQCUEXo21nP9CYiP4cImkCQB/7SBq8ycaMLBcNsPYqx0aBe8GNCCF9bB9HK
FqOc2648dvxFsHlC5UbpJxYyAf1bZrJ7OnuOS8Q/4Pdpz7JcFCs7b1mDMkCleW1T
QlIck1i80cpxSASI896CgWbJpjaV2hdxdwERZs6tyGUEQU2M/Ry7bUwPSrdy4Byz
BRhNEaMOrI/Zf1MyIQHC+9DXzWbJKmV3AgrzNPwp6bnos+rJ8B22aYlU2gVivvn0
t7P52wAlNH7JN41cmxTVOIghDRvVXKcF8leGKXuMC2nSdPOsSj6dfHb+Nw7hcBRv
0SBooNWzNJPFDVEDg2qbRFYnY79lJDaTFvk9mvht6Pa+81PfFvErac7cOZQzug8G
ZU85oxCqtTDnISgvxSkF0qV4uyUXdQXwg6ZfWQG0GPTMgRGNae+HgHk7sON1EPhU
ftItSp2K40xULpjq6BNG1/PG2sD1HvtwqAwyiV3q5CzSqRiapWxMysAu56ow7k+r
nA3v1tN0zr1PHqiGft53S/ktcureKqqbtQ2wyhLr4mTG8xe9+pmUapDi9pTslSYc
qw5XE9iI97d4yNZGBnIRKBZwrBTyiOf/Am6fa5De7Wtc4qwI3s7ZnZ7+9NtlKXBF
wc6CYgOw3kwC3/MHlr+lFD0/61CJUyKRsoSU1h9TfwFFo4XT/gY38MPIWmY0ryWC
veBCVLvLZ3E4GfLOSTH7DhWi3DqXY+N/djnKXUrnQpAk0y4bug4Wh6Gzm+J6fydk
khC3JUtWk1ZtKyg84WXR4N045VuSGbfYNpwRQGSe80Zw3L5moH3K4s3ShoKujOFR
j7L9vwQ26tLhPKH2Mjv/ivYem05d7GMAGyy+sRT/GeVqY+qpeWNwSEqRUHejuceq
RqMDBITjzcQmTG6MKTp8SyI/aFFPdcl1UDqdEXNZw0eeU3CQLEZeLbX7bqtW5Jia
QeEKHGqaO7s0Pj+X9HhPYC5jdhHgcyGmY9yYdKFd5smg5GjnTlOX7pNOWRcLgTbp
PtlIQG20rIraUDQHSstV+/seQqv1INPUNEj+DTp4GH8Sa8c6n6+0MFZpp05bnQIH
uJjP2/u2U8Bv2jr6rWM5hPKkRStibKARbLk9zc0FMU2BrKrYizV8nWyLDkCcvK9t
WyMbLQim+qD77vZCT531Kws08b3GEn1fNkAqfbohUvL3382OQVQtqnXHbHWlbVQY
+AjO0XVjVZSfbCq8/1budhCJndksJyx3/M4CG+lrCOqSFDlTKRBp1HoafqP253xh
7cxng30gsB4B3QbbkMvQUnbIcY2lhuxJ+kI15+Dj3BLoa2LslMAUFXqIkbUMPF2h
+OitN9Lcl3FFp35M4ZipwuWe5cegAllOxJrkZRhPdnDiZs4FQzsHKfRS7y0jZG2W
sDkT9aL6zweUQejKAk3gCsAOUTitRRQj982W7NLy2mISI/6i90xzuITFcXsBuNdm
B76CPSHroecmjj7D7/ykbwiLRhiCAd/AAgszEpkPHG6/eLsSYQ+6jEHu2sxFd0D7
q1fMQNgaWOzTFumQJEs0l15m9ULRCf7K1MZc6Qbe9DbDPuR1uM9wQydrRYGOsC+/
6s7BSf+aCEX1aW1P6Jrivi0A1kLhhAOqQFtYb49uoUPGCFpI73foFNsYdYjyb0Fc
FMW+8JzHezz8FsVsUrFmiI/UFtWK2oYugc1dmqa0EMMZwi94tBTwF5ASCTyYXXSa
B3A8HUFmjCPuiBiEHjAdoe+PQanboXlO+5a+89SENHBuNsNhKvR96fBOtLwJHZtj
itF38pur+6lJL+YNyCDSipEtI0DyXNGh6iaKO53BthPvo3TGQ2cJ8E0kKJiGVy1D
xJGdQPDee85FVJwdrqJzDJDMM73tfww87Q/2x6Bj/XTV3hRtwKLhEM+Ua5b30OAe
bkmGMSPTFZouc4mITqD1C2E+ISfQ0dO0/a/x1QMV39hV42476hpU65Wtfc21nE60
TE0e4iKeV11fYa+co6c5QlV/ORozay1yWoIGIZigHlwtEvSnxmcM40PT3rOBuOGH
33WH6H+UqdHEMhUZWewpymLa0FscJg1LPN0+PTw18ci4FAig4+4xfOsSgzgS650h
vkVyWEtsRYwD5UaxmTDnejCNHAlBleBKwqdG1PkzjK7vqI4TBO4y2H2OmcYKmR5b
mJNjpQyXqpCBy8IkHCMRz/okZg4wdM6zkX65HMf5OEATZ6ihMCaMXoP9Gfyz3dIr
ZvLxPClvwW9aeHMDMWp/nnejBqgDlNdRRkXZ5uMkwhaXWzyC3QbrBTlnsjTsLPBL
C1drnFP41uBahZq8nxd9dugNzM3cqWyG8UfSOeWJsvdd3t0w9fhHT3vOpN7iCbZv
WoWpSXNDIVP7X1+vtftM4jvjMnxoRoCZU+d7pFDl/AlsBdU6+L0qw9lsev2+/EII
DESZbmC2N03vbCYSn94NnddnmLuZXNeMSipYTkTa9nUF3kGs4b1UmI72yb+OZ0k5
6E9xFt4vdrk18icnDTsPslMIiAN4k9IkX77a3LnA39v3n6B9lfn1JlkdWT+8cBek
u/zkXn2F8Eaa4GpNRCTb2aM4rYFBa8pcVwvc6fP/NHGvDBYGdqFlkWZ9eje0iy4h
aVOKz463YvhnxuFLOt+FGv0NvKmsx40xZbMWW6EDRMuMLdr7dBuJAycG5VU//slT
OyzsyS4Ig6wpbD8MerUGd/3dijpj/0evuVeMB2nLZD1SbUdaM55Xve3qAFCmNuYB
FGzYl/FsTi6f7e6njHeh4mIV/sNkZPQHEPeE/wa1lFjXrajLt9Ue/C1w+QwWb+xD
eqIqQ8uTpHeyxrOY3BsVWJJiQv9rwIZo0leChULcMxcveuB7BUskOwO5BsaOsLQh
I3QuD8BrAXBFR7dRiB6x53WGADcFGYtY4BLS5b948pyXZ+qHu2UVuLitP4LHawvB
Y1cxWvZ1rTo5xD+Bht3V4BIjvHVsbgFeU2oLBT6AOn0MgCppIDyoO88NtPRb0ZeO
pii/8rtwLyIYgHv8NJwAOulwYGhEBXeHS/hRpQJxPkSGVpqt6MZaNWctdrVmjmN/
VMs9ItJd+PY8Ylayx+Y59rQI4DSfVbLbhE7m5oF2I1uSxo7B7va0zZu7//hKYNyb
QLvS9oHQ0PQXzmXrwQeDz7j92xaXN14ZY85McNr6pCzC6c12OKoVXnrbTe/eQQSL
rCnJqB8+FLGxlBIc+eG7igbTNnkI2YuwThkgyhbkA1aQmBXstNH5FkVAMAYimfxm
P91AMUDkanrKHO4Dk4K7jz+/AWfgQMvtmZvQh49Bj9r40uOSCForI1AUuTqWpmcY
oOaI89LLLK90cV5DQQ7T2axRF/S4KQTPY49P4Bu1b4HqmUysFd1WOg2ZxlTowilj
Ooufn9lxuu+hwpF1QJKwlQseX6Ea3gPwdTuEdcLTQ5gH0Y62RsGVGg18dxEGIoYf
y7Zgwde4W8jwXnPmwNoQwGhoaWfzbWnocPAkEROsnqfKKmizr8ao+QpmYOQf4zPe
psmRWzXroQs1opjFsHQhYtEWuqdH8ZdtzuCqgAaCO8vOAcGYLLbnkVbQ7en4ihWM
CB4jw6ZTqlWpcszdldPCWUtGJFq5VgRSbcwAEJAHySATWQMwL6v7jD9F5aEXfcQI
08CVPH3bksALEYuw+yBX+KFmI9XnwWbK2eOYCZXNsjdi2T32/FIadxPKgx08xdgu
U33RQlJRDaXChDaijJyf1AS7w5in//F6hfyMW4COFcOHkg94+ho2DS6qRV/XBIMX
fObr41xnSQXOk7c8uBVn2NScn9cEFtswGP8DAqGnAJn9NTkW9tSatiMhMjJWKE+B
QQAA1oP1nbyWxLCnwxsEhBq7ypFDy8/V/i1v4rboop8MTU8kb/wxvg9ZNJhaPZbo
V3Q9K0S27QJ6g1DPjf2wjbvsfVwsI+PlofvWqAfBhxp2KGNUnDMmcjhxPvsP0Krc
l+Q81pi1cvexKo0MNu2BO3M2F/8afR9cJ7EEAE2XsQJs8J401FcE+O3sQAI/unml
gWcKT3Ko4BnmRUOb+8MYvthhHVxq+QxRnIMHf8GbuWsFvOfvG8Q3OHXFN6bZk76l
arxc+p4xgdgE4AFp628jK7evZ8JVKjiFk2MTJRJ7R7+Ou6d+Ydst3E97ghEXmI0F
PuVV4K4k4VCttBsJMYtG0o9RyGdL0O/Sz17RyL0U9n0fSIsHljnPD4xQQI3VXujC
lZx3eLdAIdmZM7bdzXIpkDE9v25Hc0oBlSgSGpvbMw3AdcYhWfK7V5E/Sk9jwKmL
IMIJwHeXw2/iIaKgl8xCSVOww8WDc+zqFXCU5EcwTrL4cPjWwdyAcL+HVZf3N0Bc
uVi36ql4qBIbP6/apNT+ILD2vTScy2JmRFDnfQZhhZx1DZW6SDZdrRDW1Zxklk9B
gIoprlV2ZUpgqTtUYX7qRxGvcdF4owT7LivV7lMDRRoJ6eJif+8DkTuvU76RB2I9
3utOMV+NqD1trfbglUv3XChlqptxsxJLV9BfSTKrDG/XJ+ug/c0VbRWT5NrU9qRh
UZeSNZZJ6l13ofvJYjfpQhnvvyFKgQEl/RnIu+y2VOZUQ2nqz5cLYD194COg4kjk
vZ81VA9V8BRpbFVRpZ4xQITmxNq2QWra99/IBkkex4bx8KRJq7PPULRQrvoaOFca
NiiTyJPZTDTERHwwDdR2Di5qQm2gC3RSNNPWubtrnEBsF19iGNZgKTmAJxV8ZYgP
1AC8I0z+zbgwhASt0uUL5kIwqLID2sljaM3rc6kZ7pluqV7adcbGxB8kPKGRNPFL
FZ+1NYrZbzD4vz+374/l4ZhxSgyY43Eop5zmnOHlcI60mOXpDggzDtX8Xa+tiDrg
vFaz/zlhIE4T+5I5H2jc8A9X3fR2RQqeHWDZV/AoTwrbQ7S2j6UAs+RDIBui6eA0
v3ZEz+Ub169qWX1pjdiCXAZYBIJjd+Cq5MBvQHZTijEnL7IyG40LuHA+tgS7enfI
rmZ6QjNGT9dNIP4sq7cK1mQZdg4/SdyQ9BMgh0iWTc0ruaEPtn0p3JCYSLpR+w43
a7sYtTSsrQdn5XfqlYfebpt3bhAD5dCkzBwxpEDLDfTeDSPHnys5CxBh/2MVHaJe
5e6hMOptPVHIkiuuveWZhhuI2X2sg58CYH5f7smKBeJEow/cwT3tOWFqQliE0Urq
QHYRkecwIu50niTpRKvjj/UULOvD8Y9cM4QuNk3f2HOcR9p+c67j1gcqTK5Ar8cj
mNP4gVDz3DNfNtvjA/0mb/0x+szT+vUP+8c1jOxNYLJSR70w41Ash5GvajkaiTzB
Q51BAUjQZ4Doy9ISmfIyzT5sJsnlXWa67+551uh9aaKdmD3Cg7n80rynw2AnFT2T
+59mSOB85hiDLnoMxMfwlNymGqOQZ8h76KsqnnV9XDBR14b5IIwXHfPne9xNZEVc
XQCqzT/cUGX2cjCH4E+fb8v8Xq2MmZR7FNLisE9A7U3Hhqi2OaZP7tl7SEKzRHD7
K+/zHJTLmw1YmaVnOui4z43NkguslxYNcBxJjx857rlWsuIXbH0cLKUrq7xSOcS7
QQ6dI+Im1FhRtx8fweARDMrV451uzpzsZrCB52B+YqU0aJl3nyzHjLh1uwI8i4tF
Ff2+KsETeELYua3o0G5Wd2KJLc6jAm5W241nsqe3V52A8J0SvYEbYq5ckQCQLCh2
IECea8x9X6D+jkcVlneqEu91GxHPHuoe4Y6qJH2SvkTxdAqdSKOXw/35Yy+1lqYb
sY14H9GEq/BuAXlzFttOb/yNP6TQ/w1ztgNnKiEqboLFW2KOmLOjI3VbxFbh1R6h
QjwrQz3hgZifnPtwiqZCfem3XWqIOYaOo8azCz07lqHuCwxUWV2Y/vyBavVvxIJF
xU84CqnxQsdqNmZ4MbCUhx8d9rR/P/AnCz7kd/Cq6bWdDEBc40xzD0uZMVQYvaDe
5dwF8B6OuRMtv9dJ71+/+QuqZcxU67KuHYGmR+7E5JuFczRxeG0LLSYxv722RunB
wIk5tc2oqTnzkAEhrMUl8d17iXnh5+ksZtSBJfLZEc4bdOz+qFs5MZk7fNFgl6hk
kdz9D5yZMZA2eDkEAtdKjg1R3R042wC215CjrcNFLSAwmRlO/KtTLZMj47QzI20D
rOA5GMNue9eMFfdoanzBB21C/2jIabzRrmHQ5FlTcYqXWr5OWeuTxmsLclBA0ONk
2ZWqPRadoftMIsk2lqAid9XBs1wabnO5qcwuzI2Uqe4DfYOBVd0WerFud1zTIn3o
qzvQQ+hH6/9f92JbC+JqGdMvkvYtFwPm01R2NGz2V4Ry7+yAfMmCFDMdxXk1NF6P
HecIyUktvy6rcgr3ExElWe2D1fWlr2PvpxAqJh/kELDVNQDOSE9R+5UNgYDi9O6i
PC4Rk0fAHLSvvVEQx2DtXEzWe0rrjhLB+j0ZlBfCraS86a/ZRpgVURB3x3SQtdh2
3NzcaF9rTNJk+dFh73Drqgg5731aSYmLDP55KB8Bmx46NFSQ963Tn+Oc+klwGWPK
PJ8QHcx4pA8ZBEFlMHLkN4/8yS/s6SE95MK9S1Bjb2g=
`protect END_PROTECTED
