`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dUd0ryHDUcdfNqw2bgU/cSzhSb1bmSE6540rpwQPcMMxV/32kJ69o1fuSio5OvYd
btKGlkJVwf2dK4wsOS+oWFQtL38datB0dD0bqT8YPpP4o4vQKBDZskdBfmK1THWE
zR27qSVSziVJVZELZ2g6xtDH3OHJRiRZ+MBi0ijZzqITrV5WrpZ5tIzBPGFGwmi3
Xga9Stw7V5jocjMtBk1NiCj58sVVXKecLtuLX9G5eYmQfcThDA7QBr0MeKYHhvKL
Bv1qdR3Gkevvy4Qr6YuKdZ7QbnqQKSq25+ErQlcjjiY+1eBHIf0QH9WKQNp2KPrj
QPQDQ0A4/839mTNlFJFYHyZxngfUjev7EAmGRKv13cCVwfRgs5A14NC4rRedkPOg
Stb9CFckMpQcy78lGIWKb351WzCSwP7xxL2MbrH/ZWReVOgbRjEPxaVN6CPz/SLT
CK1Q0GRAfYaZ3D0dfLEwCrEA0x4QKMSocrFY6itUq/OWqoY2JRAb9GY/lvKPhe2F
fbUfJKPTFxLMuH2y1Yk5K2ybgK5E2Tu00bb42zwKsK0WdzwhCn/8ZbjTrFjG6/t2
4MmeyGcZIo7JrLz/0BChnBfP2G1f3ZnvvIobFILMaR3mo9VucyKRSgDok21r43me
uhZXGSdO3kaZ8JMQIwttP9zrxEY/5mDvGeDQ+K55E4dwrTxysbyumUwHDGZSp8TD
x1raudABXMSrPMdvUjJcXjiJSV7XuoY3l8AXZ6KwX/l9koqnzm+jc6HLGch4aENp
12E96UrWzYeqtF3A33/Wh1smZ4X9KixpGZ7G7bx5GyOp9co/LR6pks9Ike3iH8tQ
2YVGqLdtGWTvPlb8K7AOVgpHE786KUlTR7GjMsm3d6YsnVRDWeKhh1MrTRP6eVYL
YdaabNtp+Fkto/uFB+cDkd+DD+72cJAerFSaZgIt4N5QW+G9truclcohQAbnAWZY
V9KdVxcYBlZQJQzOCF2fO9pL71sgMCoh1fj9kmbvUhBx+wI4IIW0F+ULvLdP0mb6
T437+fVLQWGX8pvwas0mQuLqKjYXLA4/Hp8QjuXDkbDTEelRW5aH2Ikg0j7JGLMw
6D4EyVnVqaZ60NjMW6iQ0rLjRKFXoVrNu2DrNCCKJPwNGxhEMdZHZXM4ZJeyNpPu
sLzglNp0oTB9ozfJAlDmFsX8I9p9lIi2denTHKFzeD/jmFqSzG7TYY3ClgSG8cPv
F5xS4JPl8l4U1ngbZGvudqUinXop7BcijBiUuNfafW4gSJG7uqQjrIX93IpI8Od6
0b6hHqxuo/ucah+VRWDu0W+hwAsxd8SnMdJR1kJ9KvMpnIjtg/tnIGyL0rRX8LlH
iyYiDTdXIRzdCRtDiP0owGz8ft93FApZv00U8d/Sx4UC6SlJgB+CZZqbqu1XUz5x
SQRfDl17MYppOEigGdTXsC7f9jyg5/qGWCGMhU4Ix3EWIRdwUlEYX1d7S1Ysxe7z
9DE3aV0PKnmj1WYs5kBepcMHkMlolSVjpKlOUubfqKa30SaSllUecvsg1pb6x7Rj
9iPSgrXDG5BhZAmB/UuyXfw2n2yDmBs6is77kGYAVegoCbEwWSP0oB7i6Jg5MrwO
xMSSl4vd/7Fx1qWZLyPnYWtryc5S+5ZERzHSTpH8FktSybanUnI4AjWWeorMlDf5
1jaiAtc4stR39db1Qw4t7aE9nIcrshtNyMU1j8d7NQukhJ+DXL5rRzujTGnqehJd
ldWE6ts7CTXuKQtaRD+LOzlQu+VXanJv8bZI7Qt1a3KF1rapfIbceiKkvIy/Q8Wt
P+W4qFv2RS5gX6OUgBRdn6FOq0STsLD3uYiw/5dZofwzei1yDdl2BS4X4oCqEe7V
ECBVOFSrk8KrLN0oPpsa58U1XQfFhuxp/0nt9Aez68WbpqaCbY1vCTqVQU6GE52n
NHubn7Qsd69vHqGeoaNP4uPaqQb2V/l4lAduzWMMw3s8a0n3Y6BhybmgnULGrN0Q
o0qL2kaS+myNpd2EFY5R0UN+/sVxrpsE8ntp1RJjLB0w+s3Q7CnGplTJygxbPmkl
gWSYfdbmaIFXBudB2vABOshdb+ZYMUK7e0lizZB849Q+eivb7lCkvlvZr9lyn39l
jfg0lOL+s2koBzpwafwggQPoMjyz55BZH3wtiRsb02XbWsE+jB6/bo7Fv/ShwwPe
obrzT/yRvz8eTVvJyFjWRB3Oh4/BBtsrx/GdwgTyK4Z9afd5WJpGLNT5NSuSB9uG
QGyAva4x+79C9GZ5xEb9NeSNriTJJIMRTDqEjaAsrBxUSHToM8CdgVTp8fy6YWFu
EpPuTzE4qmWSyItrWuB8X1KnbeSUZeeV4VLgfQZyJeTAvBW0cSX6rQbNE1WScKz8
0ByuscAFNiAzocTiBdkbKNFdJ7mhIax51TTUO9sP3DJnfPIMBzEio9M7PSuGcCFo
Xb5HVmSNR01PDiZNwI6JOT4cT3xJjEgRk7VpwpX7dFT3mx1A5ab/Vn8Y16NlolC9
kGid659Hhp0s3+E10jBrVY3rQtOT7TRmLusSWFthBoDqLcdNNN6RcyzlTZ5kiV54
8yKnkmOqnZqB+nDpU9YV1ZgQEqWp0ZWJps+yc0TiN9SEFFtxox3IUNYbCd5ZBw3B
z+XAHz6N64evd5N6Qk95IBV+4WvaYVx640gG+hmwdqKSId8sv+K+REkBcE789C1c
O6U1UVR9zhaLrvm3a1UHHSfwCkJmomKw43eTQwQyyQSJZXYwOvFvpjKH+/qiJ1Ej
DbT59YJV7SYzGuYePjwqqmqLYLt+iEqXDBUinv5vyrEwZqKKwAZCH2ZKXudTfKy6
MZgzUs5XSVIRtuVcrgQMz84X1kBhtQN4mGIWnusHtP+RBpR/2c5MW70BU4Zc96uV
35cimrpxLLY4AOWHMgn5nQuP6tG9EO/IWTLh+4+R24HDqrYtbQxGRV1o7rpP2WdZ
uctgALhleGeJYNqMOYHlr9i5GT6QT31ziy2rXAGuQiXxyUUUncnGxpsj/48HKthU
/Dz5DC2ru6zF7ny/CYjonwVAY1JAZChUtB5dkwc0tesPerwgT+fJ6k8Htzbv1scJ
bqPFwyZ4LPVsOvXY4u6gcXCDeWiHDhEEaHNEopyMWKfs+qgI8GiMwsAEzHFEVim+
mvJkiimPkj8KtocRUIOHa5EXqY0UvpH7lTOaADocyYQbbN3LlVYiOy4swzCzvnJ8
SUlKbILD4oCpk6RIrKe3Jwn4VZ13H6+fQj+g+TTakSotgBTU7+84VMS4/lg3K0Nu
t94hdtFHp/FPHz9F52w97os0faKAKlXLtbGgfoXlR8OhfG+xg0ESv3yyJtn7kVHX
mp3jWJ5lBGN1nb0rQqoTqm5lkykwO3r0Ig0OHRBYMgE4fFiwCkSNQE1LoU19KHkt
Y1hE6s8fTDQ/oLgIR20FqyOmFv1pZW3TOd4t4Eik3b9ap7HYIxNoYtx0vl2gafcK
59ocE7FrQ1x72ntPeVMXty1fAiJiYF8uAbozL35gdIVhO5caofPPxBFftQRst+vp
u9RV+hBsqKGepD4x/OTMUiFkUew2wJn8agr0/fmR+E4IfqxSogKv5XD8Y9LiLaEZ
7kDI+zQDt4EzwjG/knlu128rSc+CUyFj6tv4L+oXFs6ujlcYBM036fmHiE6bGbTI
V1zlG4tIcISm3CJ33jO+ouympYO1hGraQ2GRbg2SsvgrL9BkWBdHJv5xUZppYdWd
3sJWi+R2R+UPn+GPvc/L8f3t6a+NY5uiZGQqZajNZ705+WvvsnJeYGBcinFePtJv
/e5oMcNrAx/MV2Xz6jiLbekrgTkJRSefLH6g03fccEHETkWarfbpYiAWX7+CgcbS
QtDQi48F2KPH1xXB965yFfDZs9OH/jAqaVHPjEHZxGaYWXJUQm2GNIgLgLVwYUSQ
OVqSTbBBUzaZUiTqEbFB+wA2oV7H+tweonSuOb1XKbCRinCieXFTgBzmgxeB26Rk
rCBCsnrj06wj3MMQeN7oflbVfxyZmTPVrRTKE1z7PBCYOt+F1zjw/MQoQxNr3Juc
9SJWjvxUE+MHU9zxJ4h3Mf4CMPJIZzPRPgFyKI5pl9yVjKvzL+GKjhd/VaXC5TpL
YVQICZLAnEpNfmUxRqGsBVqYKugHyIcUrvIy660zD0kYHk4k93Wzo1SAjKwAJJ7H
W23iNh+S+49rS4cJt8TczJB/6p7EwkyrIpSKXPzqU3SEc7SL/2tQX/du0jUYalWA
qppLsPXx0RjN/LiC9wiT+2hQvXsFQD2OTZSlq2wyIQq7cTVakhwiQuQ6i0W3S8rI
J3nf/dN5a1L5/ZJ4gVAyOchl4e4POrAQjl3o67yKmKj3yzNyxhAbOrQawuaAYR8T
KPrfZR7TsAa78dXmW7vdnhGqyTYBQ+N+TdplJlC1fFkH65dye6EgTF1E+z5MQVqs
5Dpr8jt5LB105+9jZ+6p6eXa8BxfYuWlWbWdueVfUFT3P3EFJRM0FzoC6qUOs49v
3IFI4EixSEvprGarHxNqdvdTkwz25Y0XAvE5CgEUcptYkdnTH7P8hpbDQQ1W4YIy
2NE0YdubQSai2BcWgWAaHGDak6uQ2t9o1MYGtzhIZkxaGOnJuhV+52MirGf95PwK
sH9SJCcYQbJrcY9exeV1wEORQLNPh5wkqnpM9qiwbgZsAswxn4ekVJ9qbk1V01Ij
XUMI5YUP8ItmqYRR3TFvLGDGoiW+TBopt70huU2c8uDqb2zm94YNib6x38IOhWpM
9OIiZsZJXq+5UzwhbUapKPvYMHcoVMUCRUERdt4qOqtMNDRBtOhw+/jTU3nPQj5c
3tJ+jEBKq6SQwplANjfMsKykEAEtT89t9aVV+7ZNIFP5NpxhIC3tBnWGwnratrW8
GxSm1MUbeeVvDcqTWBhRJi65cHQ7QYnc2KcFoQ1+0I8CUKNxqepjHIhQDLYeW4j6
LSOgw0T31fgJZAjGjMaIouWioi9qwKZcWudxReiydffWNndnDO0k2S5bREhYI7A9
+ZJwzr891ciAGc+8B14W2jPsS5sA/npxVaiN3UsQlQzm/niyzTuP3S7VebKYMMX3
BgUyDlEZyt6db1wwVjm3LTJIFsI+Zq6AOdgqbU5p8mstR2xGFroQuES5yOKqlkHc
gfxuUg5Hg2lMM5LGFZ5NbRnY+M+91Lgs9jA6CKzAXHH+oaqcVv6L73YE8S0ffV5l
vHMIKm1ZeosJ+NSAB6T9mClgx2pa+cXIaLw+GIiVghN4oEdOmGafnQJc9gmosDia
U8PF+b6MaUHsWA2JXDN5nK0HhpLA1j3aPi5ZW3T5z7qLiiOJcYksFB73spXNexuE
9iSfWCmyUF955aJ+pa5CGhJkZkbOK5K+rBI4qQcFdfal43IK1lTwNgJjX++TjxTC
Y3qY+cxPzYypL5z8LxuVvVUxjMsGbFuxMx8kVyWq2ZnzYvr3bdh3S0g2ijnGSupi
Q+NtxwTbNEPgJ7G+XvSDjlLs9jpgJMRIMUETX8F12yWk8P4PSnUrczsp74GQZ3fu
Vy/bGTm75ycrqHZXByTOZqevkdSkup2EaCGf6LWMeqGwYWpoUfOEcMl54B42QeRQ
axrNZlOAYTs7WLrktRbs6pdlG1C8igGLi1zU8bLwuzep+PFtvjiUndJEHxPtkVZk
Njz6t+hVEU4RDGJrggYeoIfWDJoJH4M5Hk3oB4nVw1TCuibjga3aDJGo5hyuLMDq
93IkWbz3fMYs3at5towttqvChnm+1DXyDgS0UKnxm/W7TYh/mU1HjLaDUfIR9puJ
fZG3GJJay4Z0IwKs9dXgswnvbjgGVsfG+LqpNxJclzVfKKtO7bRB9qwZGJprbwZx
dnrWB5kvRrtUPEUTXJezzJoHogQfUOlil5rEVXxK2orS9v5R10Qhs+Ruo65Xrx+T
X5jI4Rg9FMIZCG4WAaxCyD/eW5+lLwWqeb6qt63lgC9PVdhs0+6B3rB2FTqx0YjB
q3zf7StZn525U2nOotfylqWJv+fkzGzVD0AziloLWorXqq4WhDkxq9ftyR8g2ehw
U/70xJxvpWv4FMrqtoLU1WjNgABNMWXfRYEX03SU+2lTv4JvYWyQqvNz0dz7+ex+
4BkAhv9CkCpj45nRmHHPp+W4hQPzE7JiprOnuQZ4UpFGRZa785nZi5qfP8+qSCAR
5g93KzumJDo0BDBI88EJrla56Vg1sQXZxmX0ebiCEkGYwJVpMp9XCMLGXYrGR9p6
qZTlH3ssxMN/jUHxr8Dk0s9iiyEgshCSjzjvoQLINy8/+XlTUvjS9XARtqdAV1UQ
h7+b7RSRj7FSHSjExKwT1PJpTco86fD/Wcm6jffosEKUo5Yh9OlySbflWdPOpvhT
1gZ6/jkhkXfL5dd2QE7wZavL19VwoS94/zGwPmCUiHZcKL1MZ5lxdhysM7FhB7bk
s23cce6Gc315WppOEMt42lUL1U8ZcqS50rv4jtwgnIH/JAZwQjp7FQh8dJjdJndp
nAjx/B86fKcxCKdy8eDEHEK581HaqwK//EIhMwbimspZrQ2bnq0ZZMPU0wPvVG5p
5EXbzJzdYZafCwEyGcZLr3CAi3++sTCIRVh5nF9pW591IYdiLgquSm6ge4KmHZZX
gXifg6oFT9NbGuVd68kY/RngHySLjBdzFEWmZ0VZkLYxAl3NK0YuJg3eeS8xHdCY
FYbjmm/Xhaf4K/8kRzxmndb2lwAi8tfbAgwm8ByMcaRGI3Mgse1ZkEbwGNDjzC54
j28MlNuTFKTu+5FQecCQNGZUlXlFMS8WHkvNwBBKucF65inglHchNjEXs9ogayEK
/S5D9CoaV18g2ngLCGRe2MM+bayINWAdxQjqLZ26mogDwQl0EmTS9OcXu+bypkWq
fqy31X6qtb60o9cLhBj6RsrxDodpmXPNiHC3JE5u0ct+Ni9SUgLAmRuqwUNwQJa7
k7/ZQ6Tr4CBRPP3oNdh6M1ohyuiuZkZx6uUKLLpXIMAc83mZzEyIXZJhzMnrjrGb
U5tm8i9HoPMgV7G2O4tVtPC5nm4pHvx2CE5kHfc87NtkIYFQJXjTe7IcmRhVLCtX
i/kMyjoFtHrsuuJsd8MIaErnRUcZyVGsj21fhrVlMwh8vArmDuEQESe75YavzVIF
hV9tf/qHCgl0SwH2q6yib7uzWQgIz0vvMWfntRun+vk6bt6GIg9bvM4tai+u2Rw0
AmhOV/3W6c3WwfJZ68YWSlFvXKrpb2UwmqD8sIMezbVZ9qLcpRI1CnEMCIM8ogiM
YycGRAa+1DmOpDrxw0mwlPRe6XWIERVbNjRpFormaJxxIQzNOhVL9k7JLZS/4Goj
qetaBsIL6mZ+nf4+CRzdMlv6SS1w5PrYJEAnNeg0IqCOC4nOoFexyGu2u2XiwU64
hTJgVqwExcQT/lTVct7nsw1dc6AesbActJQGUmLzRJvTubYp8PLjki2gJnESCa+Y
UIBbEHJ8TS39kr1UULSWkC92fzKdQI74BVMJ3zWoLLoMsEHiFYBg04smzrfXhU8Q
qXNod2pNDiyfxhqjjS4hw/198dgNzMYRBbGK09PhqFBTmDsODhg2QGDQulWQgJwn
hVpWd7zkSujWkMXIv6IScWuR0nVAXzJNAk0q+LkD9p2bgW/IplwTM1vN8xDY+40O
781oP8HlGbwSPWbc3xs0e+Grl0a0XVk+WzbrpNOg3TYSu7RBy6O3XHol/Q9wZ1w7
JyqCSbgoCUT8h0bWH60kOh0oiT2Ud6xN7//Sn+GBrp5DJo8vEx3lBjIghBsv035x
82khm9sFfWKoQye56lo3h7VsssupWpOkXPoKBPBdSEMjDVfiQLnAMzYLttlV+bil
jkpmg9mdcjZvI5wnrOEGwUdBQ3ROod6/tmd8zZC+cmYZQ0IY8FP9gHB/lwqZl3di
FiqIQf7nFGSPvjiajCTQygKOhyaE7+lWWOZZ/wxX2j+WXKtjwlNRRy5tHItTAuOq
GSKlco1rHrx+CkBSgBO11Je2N1ms3bi82xjHcZzAs2o6hvJO5+xmexnGoAWQ7xke
PjNhMBHXQEu4R14o4Skp480gx6gJb/Z6uIf9Y6wG68n5F8iYAJIamvmlfBNBTq/k
aavkijTI2Obz3+2BYZ330Ru4LS8iG3C5x5AC4a81ALbemL9QhiD+FlfGfiknDzhh
yL4fiPxf1IMktjk5VPoR6AualT4iLAIEuiSEV/c+mp0JbqSQjZCTjSEzQGBKavIn
HhhC48xlxgTtzQCbJjcsTUPrOqE7zLxCGqWWbXwfYjj1cX13bL6/taJrDxeX7aZ1
FgxYPqSDzvONm9EEplY79t6MwqZrHEJ75jwrms2bDiGxaUL0k3Aa1uz5wJXRDgcr
+raMphj4EDTIfyLJcRyL2tvf6hC1fihXrzBdZ7YwFpPhwDPQ27OJU+AGN03BdVdY
HiBCD0XSoEEuFr29MiVzv+byLpTB+2J4nzU+0pUBpOhgKbeCHJF0aMSs7+wt7JNv
1J7mFcmrirLTzzBUTYQJvQbqd7n+5DPayx6QkSl9RPWWyb9hkK9l7tajnJSPwNBp
reEQ3WeCSRtibXnKfcfl53apjrw4owrd2+o6OkPYQfYzkaqczmqi08PaNFpIK40K
QotAgni5yawcRBt04rItFzCNlVEBBuECkZyJvQQjCndb7r3byEHepr0tHbJn2jZM
4Giy9qfSjfDXkRIzQe0UxQwfpK5fEeRVwAHolkzKlNnFjndl/oy1dwgd56tXbwSr
vQzGhtpUNAdVIj6fO0WR865DZNHXuF1dKYsVXr9tKlgMYcBxuo0s+ZBJJudgIy+Q
ZOZX19IXFxdKGGkE84AJH/krxnPxBHxmMmENoem2rCglRZ0lmaKFev0wVhweCIQ3
n8D8G6KKgZypwUoPZau01h0hOtZl6N8ZKoY/0R2bTvuRNRHKMKHvbfLXimQ9/tIo
JU5Jt2OqEZrCrPA4aVXgSqskCL/of7ymGbanVW3WsR9UEQbwYN/NXfdNe+sSjPDx
TYVBTep0m1j/ZPiAtzt91e/e23HpgbCmc3g2FqInXfzQ6kUrRODWguAJWAZMFZ8l
/hQdkNJbDVUHW+r4FLwxhEaA9g1wGNzanGB6ai5r9G9C9r2A9DQOfxMlsh/s/vyA
d3pVzpiGH3PBTCOdloMNfLn+rLRq8C4ZqS+AJuvdCUOaMJ9+hto8FcGLZSZs03rD
ypST7CT9H/VK6D0A5PDwPaTNSYbCOalylsuPAKA6MgdEy2pKyaCM7w9qoQMu3/oq
rMXsDADKpVWyvdDKLfxOaTV01BapAYY053StEhrhRAvvAYpjGg9hwYjTYKNx9azT
7KZvkspXw151HSsbBXXjWcNKqisaJ+ubxCP/tFLU75SyHnrcRsqzOrGtsZKNnLcp
nUvuOI0XSwppxlMMR3OmxQloNvLEYf4hedjL5EeLJ3Gysw3JHv257EuWUajQ0YH2
DFAdPhYvVfAhxsMUpHaGDc5if7oGeD1JHiRGcnQR8n52SkEEiIxmS21bJ/zy6Aok
PBfCS5Fo9TyBQyWUaZoVHaK1nE23pnewXo+nEseATvF1B5GmcXKCucpKgOosOn2h
hEL/tVryEd79EufMWKex32Aivfk70YNTWbBuz6t/ojqcA34uAIYStLy02AZq2rR7
Gi/SEDwkCII28oL1F//GWtpPcjou1AzPqtTmAU3bKGn9a7ChxKYstU1qMCCTbHjf
JBZiFnSrjNEPxVLzFrx0JamsrQ3c9zIA+VomrKHVNlausFWYQXXf9Fg+cwoh31vm
NniDnOz8UNcspIAs3w5FI21tTl3a4gHMFsJBnEhOMGtiY/2MYcV14jZ4ZYUFVDds
Yx86nrSi9c4XnMEj85qLq4qVO65Uj7syEFJOh41eFdkplGahcxgksjqDS9wBvQlL
h3hHxJ041TGaGKHzk47ifAwlIAjXTL4cwmmxWKe6HmCTG+k3bL+TruM/YazT/yXB
QGo96xs74zPYPAt5OhjdS4s8YGM+C5Pv8OTmpWF4PJROTr859sZIsVR7+9Aii+HT
QsWp68j8/1KATEHAL7wgBW6Rd/m690EtvVZSKXlxLzZTGNYACrSReDC8pSvVvYbh
PKrq4RLvw0ShJYSGQU6sxWkL7WeDSDEGEyyjXtQJ1M/LaZxh9z519MZXu2wSNgp6
erUdCi7QluXrt0OYex/z1OHuBSIvk6qc8Bxb/IvrSBN8D0w4dbd94o5BueeZMJNI
Kc7cEJ9k+u61ThnwhaoF2OAvmYL2jj9DDukXOn/fs39sHuYgDzVdjPvXdPqmym9l
YOS193P56LJsxaQ9al/k3ePqI7eToVNiQ8UnFPfJeI74cipLoKcYjuVUiRXD9/Dm
4YbLeEOJIj3JK22vD8q7h+ffpLqxzBnJIt6wnrWfe4f9sP6+bEHRHUcke6NpOROK
b+9BALshPwByO5Oo5DPyMK4G39PI6uTDX4bAxBy32IxyP+iro0RtGT/H+sM0nqp6
AIFyI///lJ8QPgxPudUJWwLnpK5+IOMFuaYRS77aZP9eTQZNlcyydJePXJ4A3CuO
91HQme7ZRcQ6xgj+oRhfdh5rCPaMK5XdkKhVD50woMyQt9WYn5ePfBD+kM+/wQ4T
iZ57J3/Cfmd4Cu9CKstmCX5t4Z0Z7xqBBcbgUdUwE/WOiV4dkYnsXH1bnXmL9g6C
E79ERcyzCA5v/867un/AD4CczonPyvGJw1hIzBWvokFRQY4v0vWqacLHO33mriRC
X2nGfIJ/EXZvJOiVRCn2MsAroxQeBW/QycJUgav3VCYJ2CJm4FWXbXcAPzWo4XSr
M+3x+GQYC+qGRzzIxhbUMOG9zgAD0QAa5Mts5VdcRpWDZi3EZKM/UGtL72ynTj8r
5q5BWJ80SlIj5eQCeTACxYoK5gzN9o+4JttszI03lvK9TgQPFN67KE/Ngs1uolcR
fW6DG0i07qQu6qAXf+8dluqye1Da7ibjgRugQMn8M94fDO70oBSZn/OErmgVjzwv
v09uuJq0TX+M10E6XZoQJ3fc8amZco3IhPEsHkVdX4ggIdi2V2Qi4DCRxAlDBfsf
vRewAoK3CD4eXM32M0kMP6yUGJkR0Ms2QGALyC395kwKRgEp/kqeRXYp0IkA5Sd4
AvzyDRnLcv34w6F6CtEh2HsEP0HtbmnktOnWVeJTtH+oxwp4qSljlQ+zslQAUR98
Ik6NqgKeCfyFG1ZgBLEOmWn4KNAchmNNmpXpCecgo3UYW336qaTBuleI17Kp1dY8
hze7hwd1hgv2/HCxTBugzhv8fFJB93O69cNZ977fXq4Fhbkj3i2p+KgRZclq47eQ
+chLzqlyEdzudRRLl8CsuqjEk0nEmq1ArhZvHyCWmooXcpMOHK7lxKrzTwfGZjZq
VPNgQlTCYuTUv4ZX0sknbMImgWOeEBqsGYZVEKUJOIXkpCsEPU00YEXgKJkIwtaE
UPKQFCGwfkSmzlTm41qtw6BgrYuVWxSZxv/0DYDHBVhH+t6Gr3ObDsiN2Y/RbJdM
6jFatxkdp9Ym5INN5mSoAzrxbR4bWfS5fpXUz1tM4Ag64N4AJgsiGgq/Sq9NJz4c
6WENMBcefEl4VItC1e+OsFZ9fvMnvB/KUyr+qjbbIfcIspeyC6l40p/4e7eJEIpc
RsGYCiCFXyTTeabvbl92I2gUSkGhqqrxb3TwRo8N4Zy9Evrrp8S6t6dZVWr9PDxJ
+fslCQdWVKuB4RaHXwCUTrzQ1XjxrYNgjUWAi3qvNyjzANQuD+5MY8uqekirfN0W
UsoRDQe5PcAbO4laikXWnWsHdXWedYv9rEKM1g6qf3gVkBPXj1f+Z2Rsin6BRWEk
WLJO2DG1eYVBgjpNnqmwJVMYtuclVZV4ttJMbQgR+JZ7AXGXTxMesMzG6v3eBU92
n6yZh9Tyr4VwDtpJxcYccHzx06b3m94YQOgfsKSjYr2XfEK3wZMehmPjCAd/HEHv
ZF9GNuQXRdzdm/PwxJBBV84ITF5p+SKTO9aaKQSGeDCNzleH5onYWsc/qtLB4qId
z/VZBLChgAjgSiJtfN5gdUr9V3dDfVf8jYrRSGUCP2/FP3u4Wu0Plki3afxhRv4D
pI+ToRbec91ZtLs18v9tO41n/jHcEKAdjFMoy5MgITgkf/g6wR3pqovMAZZE0Pu6
ukQKKlGZqBdWC6gAP92RZk5WBnysG/y+UsllNmW902dxGI+MPN9UIutjPtd1ls+j
lVDg3pLvKcIjKvhuWFSoYrWK1y0BU9DZPMv18zhzfEnKdNgqXAX2pX8qS7emSeXx
iPCgJYR9Ye+rpAh+akpBFpQFvWMlNDAJoWGK8oddVeQ4s27Y8m6HUczGAypGgydd
mSQ/mEGuJjQXx6j3W7lgS9Dw3Ql4Ge7rN3uEsTaZNDwhSG/GCB8BWgYJJkzFk5NK
T2f9+XfQGnRnC+erT2FCNOYaHtYVwHYKyjwONiy5ny4nD9mwBfzlKIiuk9h7D3d4
dcREKCS5pkd/MQcP2TcJjBpuMtUV00jSAHloJ1uoZRf903xeM97mW+3sYDQyTzCE
ZEg7YvWOXBfcx8FDp1NSyEFFDBQKMEvviClN2RiFrkipAH2K3zjspDI2c5lBaOkS
x64tjWWTuWru5WEIsqf/xIFvZm8EMeT0ASTTfObMlIceA/HIiny8FSJ5zV8EnJfq
E5iZZtvo2erSomT+AWRuiTaY1KDc/gZ4rRGuB6HNaQDE3WesdCzKcx/yctUZupFR
vmoTjAVnh/odEc3KyUU2ssJ+0hsMHihYwjD+J3kYeFyaUPOuBnwu5CjRc8iazulO
O4tvytXoBQUVMqI6fpa4olvn3mSYANmdXwdqpc8/Ce2oY1OSGoBklyjofbS3F8M/
ZdW5gaIlA5D7jTifThuIEGvC4IcPktENTtnqIhSBF8aHCLsYTtiStTjb3UZ9aiGx
3JRcbcQHvPAESmFzBbgnv/oD9VcLWGci+TihtCvYBhczxGNt3En6wpT5lSH+cbY0
kEBlX3mSa90pXMZpD3XXnHRxIdCaMxBM2pFX5xglY8kUGJHTIhYDUqZsYMlGoKji
K7LbJudToy+WkZ6Bh4eBOh12Z89WRrK/t7HWunCqDIz7a3qtY0KJCACS94K2jRIG
xS7rg+cYDsyYuww1l9+R1n9wHBrE7CB1pbIZ9I0GtYmNbLnMIaS4TP+mSPq/db65
4Ni+X5roqbFa3DsBT2FbGBUy3A2I87XZqg6cDN8NK2KF74FiwMmFpV2ATxeOE9gX
bxyOZwWoAEDm1sALg2atQYGKAPA0kqSyB0peFJ/e/sc3eJaXxMI/lTeojZ9MesxK
Nj6Xnds6j+onkvp1Q+ymAFEdAPcFDsn2C9mku8aU0cyhiXklVzwRY85OJxJFkrfZ
CIMOIM/aC6EKppOY7BJXU7tG+Dih60SgYkJhGLyt+9JVVw+6JhpM8yvwpDcgp7/W
1FWfkSdeBvL9b6jQ3IzoKeqrHY1wXReXcH/yCOn/J5IZwhRNAl2ajpIA6kHfEypc
v28LjS8vfmgbQpqji1YzYC9dszApdTQerS5oWwi/VW2b9fWAUWnN4b1jpbQ+70T3
HKQRbOksyB75CFDEaJndOyZz2R7nLNqHHgqveJZ4tkXm1XYgwPlNRVuJVZS/6hLS
LpxR85NVB2L5OABSSg06qOR3gw1EVjV5bHGB7hHkw/6T0qDlrlKByDpvPOU3c9Nr
SeUy1exLZFa4DsjRBfZ4QxTvM4wqXU9dKu3SagVa42GsUzhu2E+VtIKfg2R4iQjT
UDc/nAz1UcgkKMlBPg422w2qQFKmXdPaWDsL9hKRfgsjH1cAfAA0dAgPuO5MOsNk
R+vy+M3H49B+pcdkXgWXM/vTBPdwzsso2Zq2o7g6WL9GkrPgoUlZ9caREEESroja
LuJTKDC7Y0Q3yeJDgvzfKoJ0UcwZPXhs46UJ42YtWDKsRbLCitrYxZxVhtuJXyJE
KE7QSsoefpwnEn96CxxkIE8YreFvoYAoMLZ3+dbd3JyZYnEHSmxm7paoDiVQdvn1
6f+nUjQLTvEYTpV2Yy+KbOqji+Ijjr2ClUJLLZq2BZMZZiKi7TgrQyxLjirDaCre
WGHJksLxggnjHS9TGnkOXqS0KXIf2kuJQRdJi26/LkxaPw0Vc8lb5Spi91nCX+ll
e+t9rspGgneZoV8JZi1uVVUetHiK7r0H2VHo4cxm7gVOE4P1vAGS4Ckt3koHaf4g
0vfvtUO1mAC1XGTsSi4rZLeCsxn91D714iOyCLq4/tDCIDwnF8VZVzJ1RkW8Aoas
qZH5VomBbQZh732vBkTukbBV5bo25zEwiS3Tv/5Q2l0XAzaOYdVkKMKERfHXMSDW
4gsK2+zEfOfBFHtQNqnQeA6VcYYUoXog8J6/LsonZiD95jxEXir04yaJPQoNduf/
bcQP17tFjo+XpR9MYvskeUJAQR7ZKnhmj0YUEOiR3L7xgAVKHAYzQ5qI2pjrLQj+
G9mzk96s7sPwtgZy5jJ5W7A/Oy/mfHZpqeIUSAYbtqnx6czhJaeMLa644r7bJ4fb
uC8v4WBG4wcAmg4esObu64yaJYpyRtHx9irsmGNmv4H7bFBrvpudW+ARs11m6UXX
E0x3aDCiXgNXA9RnBwVwHr5rP3W5I2iHZmCPOzgEPCRTHspbu3LJgE3VSDZEmD07
FiW3NSYjpz45zxnKHaGuuOpv5wrgvqz5szGyWgQRrAMPYsOESSg7CK4TVlofMVkT
jUQgk1rf0SXOIC8Xk8QptPl5M8xE8b4UfB31xJY5tBm8W7wHQL+MoPO0pG9H5cR6
B227BG1R//LGmuP1YcuyDEZZZN0urQqkEKvUDDrhhEQscEzMQUnM6UsOTHAabVKJ
ftwwBzf7OdUX16DKBq6BNNuW8pQ0EzkDIc+w+frjJ8p+SCPT8vXdfGtpUkfdDMYj
Bxp9vtrQxEFzWcGjEtoGWqoVPxFIN4HcPMD6OcN7tASMvHmY/Petv9iETKmVumTN
3XPJEFVT1+U1bFXkPLReDWpJMqkiWZnC2ZAdC9j9Eejafp8FB5qNJs4Nc2flpX4b
BSCJfpfOBDeiPiQMuOVGSyCWTl3kZpuZswPAQxBOKqcCjOb2lIe3ftwaEPiCV78j
X+EoENkzuyDlsF0rcEjfHyIWgBnYDICPyxzLSJl5+y0aGONxsU00ZlUyEbM9DKVD
9E4bkHda03LjU1AoExxEv6WuzQwNnwVRCHIsPuWbVCMp8OIy0v1s+uWiIYJCid7C
EwOJghC2+rvl0i11TFJp91mPidJCufnRM7636u5MfbX56u1abj887IigWzNeTlAC
pX+g4VxOV+dmcLbZUf+3qOc29HRphgrRGCriKgoWe7Ys6qqOR/QlNga9sQJO9I+v
erAmlk2M4ByLvEyjBQml9dclmgP7pL6HHQyGmNR8AtHOTGaWUxc31hLnrpQeXnXO
QjPNvU8X70fuQ9fEDhVCXpFNkLAIHZbxNF6nfDqQS1QCsGEY6H5pW5UbtJsMWLLO
AyKWpNet8e6s+9McaKztV+JBPy/WsOUQR6o+Bi85C1y/Ek7As0/py+L7ZrqIqARb
Grz514mEZqJW5bmUWnjdz39D6hFoGRVXyztU+WDWgyYukLLOIVEQS/7lSdEW+eqB
nEjXYJ19naW6q2mRNtBV3Ab09GIEEFq4iyFA2xOQUyGTeabTktlaw8iICkF/D46g
8V+fRE6EfiKeIl054XhqYSDZ1gwQ/2Sh/TV4BS5coX5eS3S5pG5NdjXJdU36uv1l
TC7NkVD53PWrfPRWzRtBx3yFRapBOSTUl16BGMn/4PUClaE4w4yLtMx9wWX728s0
i6I4m0vBVDksLBFvxIA3D2kjKvRnX0RazZ/ZvVFkO9tWRoDCon7k3Wh7kTImW5qo
VR89kuwhkkqscaP/5LQWXHFRoFG+W2CNuCXUK959vA/Jv5S5Cq1CbYkynhUQxI5i
X2kMGzydSR+h0fqaat1gFAuZKp+Y3RJx/p5NBFmHs9wLFt0dd53xWvv1oa6gsdFa
tWzG8nrBBKDKwevctDvJLSu0PHhmNFiqFKW7spD2MlqH31y1MfEkHwy9KO/bazoq
cQzX/GuWCgQHhs2dxKEk7KidwJb+d16EfIdzYyAMekHGLDHvCGGZVOCGN1Pxu0FM
Crq+pYaRZJHPaok14okGdFsB53TE+dWHFuKPsmJNOfDVHo1PQxUlBAANUsRtNj9q
XAhS1BEGtmjbIqBZeBNjH3GNH4BA+4eYD5Sqb7e3+uEfbE3pdshf+hs8Hhjv37mW
072bFsbJZZM2yAnAmgP4QP0NUoULxsGmJYsKh2KxQEtRaAM+dS7PDWA+2hCS1edp
IpTaDlc3iS3jUD9YDVFcfm8Y0TI9SNFRJfByXyk/sZTWrQXp38+S73Vhl8KSM2wS
KDYFxxn3XJYXale5e4wUx26BxpLKdUmas2QCkKCMxwEzP4ndp/w1uzRtDzk4P00/
EuqymDszvefYHj5RZzZXSFB6FjtBV1KK+K9gynEGoaeNzzXYqyFhauvkP+KUH1/d
l2GAvt6aqwY7+4X5LWE8jxEjQ1zwyl2okoD0V9PVrncFjE9gv4ayQmPbIZSec0iZ
SmrRIQIZq/EKYDh976Jxp7bKz9OXREyiSVVMqJ2Z00mcOdn/wM0Y8jii7dVP32Tx
kDCpSv4PZrcx6nYx5ZJuVjTnN0NOzvPq654JS5ApXJXL1VA9aX7miGMGiFhlhRKB
vmLgeNMQj++TDXWDkHKdOxpmLaZvy/LJGH3WWq0gZ6gb1uKoijvh9D3l/5ZJejuH
o++BeeZZ7mE4RXtw/jqjM00WdAqY1Ubx0ZUpyu9fn9McSQ0x+SEXja242YjqcKmn
+ygLWnlX0/sc+ncXd5Wb2LQEL7eTs8gVRO3pO+V8s9KI13tvbLJMpr8/EeJK2xOC
WUQ272snlIf3BGzO1wWnmeATVDGi2Mx4Z5Vf5VPEfBJYYX6mNh9CiO8VZ6uPNP1p
ox07bBB3DlGYTv6lU5yaLGrFkSP7aLpRiV0ve3FFFKtT0/lD7QeWCbqgdGd9nJLV
Gyyid6snqaFbjLOFZozg3KYZykkdTPW5oehCKmCPCFQ2I1me+xPI8yOD6api11p/
N3i2BS0CjCdHy5fPwCBesrJgQNGjXFKLrsP70tyVPLMzLCAoq0Wu5z0pXjZFA58x
UVudgic809ZGEAhDUViD/63RudhmQGO6ZaFd0VxtGFH9Ti9qOPXcV4314McmIa+J
Bh1G6Jx7HwQX7BHDHwsLELPMm+kJg9svfHc3X2+OIami3Lc5qM9RAPcSqT8MFEj+
A/ZP1KyENN+Bvaxr8pBKcPG/fVpM/YIK7Lbbc0f1hYgFjkr/WHvAvetcsKAwHfbJ
XPFywdoy0iAFiPjSrb/LVttcfzhi1jsXkTihmiBMJDDVFe6IIekGmc2m+85tbUB/
kfyvreLlCQdTbfDRCc2aeIknk1RAJz8Cc1uGnvXxZ9MgKEHTDTXvBUOszUFW6F8U
LyGCBwnxDu1jP/Lojr4R/yozPoyi00kwrzpuSClxDt53StvUi8s4o9Gy9CzUQaXT
3et2dbpGVjkJ3VwiElYicoBIV3qoVNOB8tHRy6WQBpqNSWEk6NVJ3XcbQoooi+IH
PyTD3XO8RQ3YyWgomP898aZfeYrgQgc2MqpOd8WHXEDCPatD35nsFcEA6LXW8wrt
pNz2mTBl6uzKFBSr1owG6z+CQ+GRvWkP8Nq2u5w13K3kKhJT4WD0VPcMKDnw6iCl
w8morfgJyBL8rWCoHWqwBNtuayy8SobNbdgsZ3OaxdJi3+7DVr56ZhG1QnqvM+hD
XJi8k25BucU/WYlrCHN/K0I4Z+PtPOCdbf2hr7dnyOWMQAfyuRC3o53gtUDJF0V0
0W3ZKmf7rqUm4/89ezBEOZn8Rkk3WoDJ8pG3mVzfssYWI2WJSzUCQ7zqYYtVoOyQ
xmSkaekhgDJsRZ7mqZzHyuzIEhNLdzoZNQYAzZLDjtera3HS2XdFagtQ1zOnYcPi
I3wD0jQXXfaXfLL6HZK/KwV7kbL6U9iyRpewLHYpzO2YdK0+uQHdGafvgRtAYYZ2
cPHK/3nG8qru2byB+WM7tvM8PGVfNv+rAHPLgAZJSLc7dl1r0YSgjlTdvlTDoMGJ
wn6gIGZRo9r7V2BlBiEKvtjItTVnCKmSEWZU0JiEESzlqqhc/gvdc9fwKIK2t1Qu
pJA88IsJzmvKfal8EuwuFdul5tGj7TsYlsYfS8b917X3jk6K0+nFXI1AgQPF2+iG
04w2whyAlWbAVur6dWaPFQhW6bhdjDx+TJJD/wyANghYSrwBcr6Jb5Dp01r0CG7v
sb94lREYVP8anjT2ZgU+t75g8GRc7rO1r0A5HYK303M488E8MrVaam4J0XzqbHLR
hmnFZ5isJqoMjMir2995qK862WL/mFJpEtshoppDSnH2nbBTwrjL0G820PTPBrQZ
iOgka5LKjONm+SrUyUOvGuP9Ja+KlbaJyrUX6KYaZmsPAsx903KTScRmyWvyQPRU
ELgcQihq7065X1tZ0J2GeOxt27cWjwt1iAUFXynXcpqx264CFtFyfpZb29qhcs8r
FSgic4XT31DAlvwiN+AvAeEaQ4aPid4Vu1EOyD9JGWVwdnAJlBDaYGPBAq3FDLIA
fB3RhWOVtQsH13uteQV854S+3pv2w0inuhX+6omf0ose2oUqUyXcFJKSpzT+cL2l
4OqBeo5agKKbtsVjthRH8MJ9qwwPm3mg/5ToCQf5HHFzigWsesqDE50My0hpN1kP
wYoFq7dTC+CZus9uk3biWzItDzPi9OnGKurrUAw1U+LrcbIBM+nE8kS3jlddn8Hc
yY/2+IFDWdscqZXi/YsJ6S6jkyO/fIZ9L0QZ/iChLU2qhmgnFi0fuU3LWmjVTd1L
QJUc2ljO30TxQ1tgoOHRaOOv26oJs1G1WyOmNArPlkW2idCR8fTH5rj/HBp7NEPA
3/qHK6BDdK8swBQWb6oPukFOOxdBBM6IMU1LQ9faTKS/lKbHM9hpHT5NOAsvCpRp
0aeTKT+a7ftcI+qKAzCLbLCdHd8Jvc7YTcn39YzeF4pJSrOH3fa14raHHqQNJQhQ
CQVUvim3tLQlQ8eD+Gy+AJuRs5mXJM2PVKwg+zEto4/BD9qn8YvQS5Rg/OhH1VaU
ucBotI2s1F9IexqDFaJxEGrxXr9TAtPZceSK2m5+UukhUVDRoEWaMIGgyhN+qEjH
m50XSnCzNdbpVmyRjYLN+2KHcdQKZetgeRCPCKM8je8KJwYhti1WrWm+ikNHVAmy
DRQQXPiEYcFSAViFFOnxcthsU4hnODN36vjW3LyoDGsO7sJktIcZ8/y+hsDoPvcH
C7uW2ZIOZCYK1NHEQzURnoQm9ATmv86SlBugWSj9LUqahmZoQhuMeRx6pGT4+9oM
hfG8yeP0neZGiKbPmZjr5BDi2NjmbSURznyHlcCy4I9X9KXp0wisTvIOrt7xcsWU
gKkImryksG+QPHfNFYLnGzE3m8h2/CjeOeMWuxNVD8ldcp6SVsEH5WuOcqgOywWY
ES9qvbeadMNnMHVtBQEmfUrcT0Hk4rlF6pA6yBp8D541vyxVDeKpe2qfunOZD4F5
McgFKLwAdvs5jw1fsqfAwWN75M90mPreRUKc+SvrgkNkJwI1WCVtW2m8ZTWBIn82
B0+M+rGhbAGsfMzl3zUqs3QpIi4saRnk/2D0Pza6Hlh4Qkoi0tDabARdbEFZZt4t
OSHe010w2cqL2E3Nla0Kg57zI1EYtHllG+xUDT7q91ZbIVcF7jn5WCTWWXuvbMoF
tzZqTv2hqNE55AJWVst6rOvoY2MlLyE3W5r/xT/kPpxIbWc6ni5V8UuZFvFxXsFe
pWxiUaVPQziUk8mq315+Rh4V/2KS8EpE6Bj0gxNBKVr8eMPhuh3EJPe5TOHq0Q17
wAdBCXnY2xMXDsvCa6dbbA==
`protect END_PROTECTED
