`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IVhs2Egbi8MbWWnQ9j1xZDnuVFI6XpYkPI8FiFmSa422Yb7Tb9f1uYWwjcZmqhQV
epJ3S+/yJ1ABqLcSv85goQGaKDyKJvP16OhkUrKqBIwUWz3mVDC+ozvfcUTQci3v
OtXhALog2jWJ/+RoWyPEL9SF+nnzjG/qUaMcdZzHcSInK4LqCv23DIT7idqlV7ry
StdEcCw6ZRN4FR/ezUO0PnKHv5jkv1VpAequePLUaY880i5wvhne49rMCm91Jn+m
O8a+keyasPVwLZkvTTzpzOAoVDvjjTeEKFrjhqnOkcwqnLANkjiAwxi6dCvubWhZ
MbCqFOS57oVAYpy3l7Irtt0ERTcUCE6551Vub1of2JfggBEq8xP96vCR+aaXYrzY
dyWlgK4fN06ypgmNK6K9u0nlDuFCN3i05zoBTC8FJiALbWsPJZ+HUv+q2WluDj1s
GFsuuPSq52efiuoZI0DRhCBS8ZD8L3fv/P7qQzozZNYdgtSxCz632SE3cwsWzyJe
fjUHBCqt4nv+Xl1NXURv0tO7IJES6fVG/3h/k/QQHdvSuek/vxkJifAr32V8dFmA
ijJAmA6NQtTB5qHBR6KaWa2KsZzGJhEFoUNgbC/U2AWWps2cQnUit9sTDEDspLE6
Jy5nm9xOZUjEsWYPyAuXLQJDXmCbKk9UJqzvrCRPjESdO2nw86IfnZYKttCa/cHC
1TUbe7g9chHZ3M+Xju9TWyrRJnES2PoylKP7hcFy43nCVEHPIWVNYtzlMqKFw4Xp
aoV6OL+z45GULuOs71Eg+HykEgYRFGOySRoXWR8YPkcyxMta9KgfisBtqPeUqegu
sehCoq5L6IyPWP2ZROwsnOD0Tb9kxmpae8DY1y2bRn4TeZHXISmauS8N8Ubt4pM2
m3UIRQyCV8uaqhMRbs6f2dzaNtuPqYirX8bBdNi5hRzQ73SEfNerpuMyYvXRM5Sm
3BnAbWHdQCPKXKbeLE5jsG2KBBMwmaeY1s+n8iPzSWJeYv3E8NUK7TN+1KcSEMeD
zVGv8De9RdAfn9gdlv//8mOORTOyvb7eOEtyIxqp8aEd6NleAbUwQewfqeiHksAH
lEmPzHiAZe82p7Nbd+95caVhjLeEbLPxuIFieQghVcTYWDz6Yr6+j+Dmfqzslyd+
N+iEoct1SWPhkJMnd4ALH5GewUHI176kWx/f09guF5TPCyf4zjAySFwNcIvvnvf+
Uh5BYM/VUO9S2gn89CCqeQabgkC7ucXEe8flaCV4kI9oFvGKQh6d7RJJ6wXvk5ju
Oh5tDVcLarlJX6uGBvPBclgbGYU8DCkougQLve+Jv90MEGVnG8aGC2JJsjcJ6aAP
cEQg06QjYtLx80u2hCLqfGQuwQhsSTBOXBp7kjU0nQrQ7MIPzMbT7zmLnB+vdcZn
Ape7LiXhEsIMtjDJH1DbCrMfjdir+phf2X3n9fZ92jNC6jJU5Oca4Ft6AYPl8fBe
z51MWIIs0kEmZ9Vo6YsMKzHfc4oV0PVm9A0SRVDxLBShbKJhNPONSNN8uKBiENwu
d+9H+Cm21quESN3Ob3YVXUXqB27B1P3Iy1+5uR2xTSINyuanLwBlfMRD8lr1G3jy
ZktPH5QyjJkk+a5nhGIZ9YgzgyUyXNiCNoLQCv6tHCNYwStvk8jNAdSwq3YoPFXj
PNHI4q4bKnw00Nl7evgFMN3qEzRt5olgRbLb56Cj8MmsnukjKXJoKwkl+tBiqqIz
xOGCm0RSC8kKMp6XS4X0OFkVEEezvyFosmixR8H+23ZjbYxNOfS3zTkFZOJ1z4Ws
E3ZqVb6vmxXNnSKrIOp332EylnWkHTPENdUIQod0HJr2P4IHTqE5n5aWhTKYCcfv
I7vNY4g97+OWLiF84H/0uB1WnEHUBYG863jQXu3mIr1OYck1T9V2xw7+iICRkyT7
R0i7YC9yzF0ZHI2mNxt8b49dy36ZtRKmkfz1JCRrupgQv64FZXCtfeDxkmwYK18I
76IgiBbFwvbPE3MX1/0Q3YoQYc0vzk+iM5UCstJJUXpZShQ7rMyQc0EowM6eKffM
K62rP8Gn9C81Kntgthqfaepwpge0CxW5xwOo8HeDokolo/lTIcsfSAbKMvYozoJ2
CVBGJEDDzg85lh/INZVoYz9Vip6aplgwAhokyrb6jKVBdsZh4Hjgodh9qM2VYRt4
3uttA4S+neL3Hnh28t5J1R7somdpH0FtlWLH3tMCb/F2TWFOx9LKub6TGqhsEmks
zHdNBNhH+g8n76EEZ/hVPmMXtFMlsqZdO3jnjrUtOeJZS5CYmG/xPAsYBul8abco
7kJymEhiLSVLLIN2s94YYd1baCdXF+nsCBjzcjfBaYuztbHhBYgVTNH4EULx2kje
DlmaJzxQ65+Sp4q8tu1hF6xr+l7SSdy6brK1waX6OR6P0crsGja7IeYvlNHaGNRO
f1VZNkxx39r960odSxJwdVgoe9G2zsEQG2p/bIwdYgq3taHKpzgoqmPYzt+s1D37
50TJcJHuYbxVh7BtnEFEfdqlhCSHfWlr9XSXdta5vJWuyfqDrlee66yTkAL1km9K
nE9HW5cdHO1VrkGqjsRwWRU5tW5HHowb0e3tNbOT+73zwdyeAYSc3O9Qiv5N3B4J
Ekrf0P135Fh6glaai4/qZXPN9IToxykTyn3ohQbsvUJ/JbBUIT4y0GnHtMGYdWK3
y3osSCQkn/a49mdjlg7oZ8wYG/VvC+jjdhvkJp7dlkggl2p357Pheo+wrBQ3tXVF
LoeaICjAcm7YKO8n8F07F2N7xfVVQcVmMghImLWZFmsa5dEemQxVDGxNnF25TM5P
RTufGtkpQkH2GubIV52J874nP1O64wQOeb0sPlDnufGh4APDVH/Nv3EpugByXnIC
t3xt9LSvH8xb4f/awYv7AaDvMR/sPAmv7lpO1Yp2LGA43x+YrsYEb2C/fKQqlIcL
qsM53b40jUZdWIIiI5qDe7tLp+h9EU80v+Gmu2MyVBb5s2a/jVQs7lI7s6J5vCq3
LYwTTTcxzVI70PyWdKWQ/MfTVUVXEmAPrSXIJIxJ8TYcWqzy8azJ40MJBrgYyUcu
KT9mRIHdiC7jgnjimPBNEavSdp34KTZ6rTeucl12wBv5g9hYo+u0temGJKWH6MRx
Kx4clQyrX8kU0/malCS/xd5OQbXaRaNg+33DnYHy+LMQva2UTKUVoee/fWyvyZV/
G2Okf+qoHtux4ABrXq9xeeR80ZIQSAVDGBbLANO1mKuLCK2ji1HyWUYoPIOfk0RC
7BsXhnDDwXGasuqf+1h9IpHFQe9bygSda9fZOID3D9rzgJE2YDgioREmSq6lHGGF
y2HXXAoiAMfpBaGApSapAM6o8RrnoVNHWB3AW5jzsmNjtdMnzP288RRZq0OB4c99
pyqhbiz8Bkp6Hn5ysPgpCWYzbeOBVQILWlxl3HmWrtDQpUARhWm4fPLRPySzseNe
5MlEZbLYZ/cSeGbhjEcRbAWPLjzTyjphjbP9MVntzwIioEda0/qi5JClBr7ZOmE1
lfaFgby0eebyTWT5oAG/yOb6XuS6k4W5V5kUTepSQ3DmvJHUO0ZuwTpBUTfUBpkE
DUxzYI4IhCRsgOYJ69y5wVDuYPDfPoNfFBHf01QL85P0Ygg3r4QJzUJHP6l0NrnP
b9jebgXsyl1Dv9AIzYovFoxDhUWww9w7m6edYUAxirMT6tnqo3qXu2V/cXhQSYJ6
ajh3rrNii+osjIAfh2zZbiSjunYXwyKak1K7PHj6an6FPTVRQrDX1DIfaDTK0WYo
O8YA9XYDSbE7BKa/30tUyc+I1UhuT+DVZA+wgDuxVAm9Exh9fNZHJhQz3XBwJGZr
QcRu3XOGou5GwE923WHiveUnW+tBWZOrd5on8guTlShJ58XILBZ17hpkOzr73sFE
/+Ik2OcjlnQLOXtMjiLDdy1l+/pQjuzvbrGCv1dkaNcOVkKwiEaOF8Qe0pZADyqV
ZNtyRIC2dwDR7jMRJYrAYIRBtQ0jdFnCyoZH6Sc+NQFCzokPhYsjUcwjwNHmge2i
nobJ5/rQpCdExns6KJ6R0JkKUFeGSw4gkW67VCkuATQbV/OZtURTv/onVgW4zvKi
1z3BWZ3lRLPOPPct/sCSYkkGyYpVjMLhgZrvSzoVxIH5cjwrU8kFyUWmHc75Q0/6
VkNLTEmb7nw/LbEbPJdvIC5m5PZyYNO8E6LarsZrC3FkERxhCTgFeQ4F/2Gj46EC
ykk+ZbNTgyTUhcurD4OYm8LbyTBH8GUL1SzQ8V882o1rBHVBnKffXxsR1fdXamBp
KErbXca5cei0eEPeuCCJDJgdvck+Ula6jhtP5F5Aeow923+xb+uh2ODCpjU97QgU
77YoblfoVWPdgWJX9O6aIzYilwUSoC3sMdulhFzt6L14HxzMY3bKxciRX+XNc3OJ
WZieUo62u+CKVgnHBaK4B9+IlDjZvIsEc7K3m3o4HSe0xedZX6ZAw/w+xnxNcml+
ZsQmFhE8A36t7uRTIDeorwxKm4iK0KN/7KNcm07h37AYY1xAzjjvHcp9JPLmA+B9
N2+Vsal8/BY5HdJACHSN62iv48OJxo5ODEt8Wr7z1xfj0rGF44zR3lNZeITLuh8F
zoMFwHT4ZRslFReJafw7bA5tMLvA69OSp3DbnrA4Wpxe092w25gpaa2mgukg6zyb
TcHQfdEEfz8y9HDKi5L8WBak+qwxQSaO4yGe5ut3F7GA/KjCpcpxByilygUAyQKq
eCpv/PuRF3Fm0KCwdyqwpGrTyiE3+u8jyBHMHO42YmMLYoHp+htD31Nc0QlBG+k/
ohZ0Cne59g9oN9RtcWNiMQj7eHLsOsLSqE7hDXn+GLjToQe3t+cv2/VVNTztTXdU
llpB6KA37B9jiWa1OPU4G3VPdSmfknCsoHbDF3C8rOaGKDvBZ0Tg+7V4kyxM9m2/
sBjjKBTMzxnDXQsJOhSt3UUrkETIFgDGtd/hsjCnXwXO6IqRNcxo/nSiKWuCwgD4
jB0dS8fuLVfqH6nqqj06KFCZWQ+PJ0HqJk9lsqJximlpg7htolQ6K1J9KbzIsLhN
FfOCSiYGwxi8L4SKOkGYDiAoREsIbziT9gsS9lL6fNKVhE8HpcEK2q1Tn51QUHs+
HKogrPb0NZ1KWqyGC42O6sidbDTxVjj8o+c2kFF3f2a1Y0P3bqa8NZYPovKKLesN
JZZVSBVgHsikN4fGDEz2r+7wbptC+qqht0pvT8J8oCnPJGXoAQ8ChKaL4OubdQ+d
Cck7Uv07gt//VGrlA8rFN/yI9rRGVIncKWsVnf0nNS5l5NDAzVCeGJ1nJT+E6X75
2ON1lQexIrLyvynm1qhl7Lkw+vqfDyE2Utd/Sb5qI8zx7KuJ6B8wuIgvvjYzknLq
OMytsP0h8XJJKcz8aX8Yu7YmgXvRan/NVkDQHEgIMMpuZA1Q2LhKc+p2P9LbS8t/
8d8TODZeYqofTiiiBYiTCAkITJK3GzsQEfZYjn5KWFznhXxPlgr0V4yNPdcNLG4v
6Zmf8ECUShZvAaiyJFh5AwX2By2LRCWON2G6j6jaxbEE2evfLg7TBWP0hJRK9P10
jABcgtJqygnSbE/j1XDa0vvwNbotjyYmIG8X/JKKXlu8hlQwrlhbqQzDK8Bw9geN
NIrPkJXLizeF8t3AWcFZkFcB/0s+HE/2yCOXiqBAhQ9k2k9jnN531L/vIeJlJfne
a+1C243cSuanA3FLzocPa1DWujCZs+QUSSZf+r37q2+dkdD49fZHiCSCs/AjHdzq
EebNeHSh9o8Rox5HGTnTyNmmyQU0BuO330g1sWOQLz8wa0cwgPVbB56X7Nsq3f0a
1psuAw5wv9ZssC0S8NPBUU7lRbPDMWVmPvWpeIfJdpCSUMAUXuK8usSFE0FAKHO/
WAZS6EXThoq9+OsED/dZmxyHbrmgD2GZ3BM+QX7MhN4hINqO9mSMVJlr1TOUuAWu
Ggd8HHFCEIX3PnGY97nv9xKgC+gJ+bRng7xNYpxV0nBRauVn8GpApVi5d+XzQvvU
8x2CNP5lQyneWo9fRlP6xv6qxsCHYes0cy2C8rnn3xyG+sMeWN9XtgsKNl+HhWOg
6z42LjmvS12swg0dMrvyPSZ51EoG0i06rGSsTmDVJ3DXojKQN5+oO0siimzK9wWo
oMt0pJFfEZd8dlOV+QtybKl0eoCzVY3B2RMjpLs2l6rhqx//kvsTtpZd6TMuYIZD
BlVovWd69Z+Y1cfsWauI3zdpZO/jlo8yjccTI9lwI8fxcUK39m2k8xA+U1cE+Jga
aSnsQt2UEucumETOlA3HpAo3YBi1/79OGCOsJ/m2VCcPhQKe5VrmusAX1QW7djT2
2QYVKXwpNSO1lMB3nBfryI1NuceOvzmaDDbHr/Frj4R35PcfzQK6X4bMAbq7kPpi
gzjRG0jHKmjxhknEGCeIlWJQ2gR8bqCIkBJazFgX0RhkHE/1if+2gZc61C+L8CK/
brd6A4/OVPEvzbWpPpcxuBalUc7bdQJ4MJthYA/0S9GftE3e533HkFmRYslngoAl
pxsSRZG7ep4vmuNLHXJf+j6Sp5zpTgW8IW8LIWS48W1/UZV8piy+7HoYQnmS6TAD
2kFNWww6FTv4fJNtzM0N56+Nj9GkDITOPlgRBQkAN2rJIEYS0FRA2YRNaynNdd5Z
/pMX+csPs07l5yNHWrefslpsr/wlePSQUYmDLvw62cPIeGqZevOAy7Fr1rYQvOEX
SsjIrnK0b4wNzDXJ9YzLYACzuWBAQ7409eCovQtD0LMJsuukbxsJ79hNwGgiyQg8
6oWXdDMPhkgfqkJByYUlN69YWyy9XVo5iqbm5yyOJKAaUyYxKyZGuVu3VFny2Y7u
BsJVgEqyQh0PTg3CX9e2RNsDPC3umZcJh5v8U+nuAE/HB+pM/dEKJ4fhr+5gRXOa
BYmVcw8Nrp4SwFE0XpGVDC1fe4tIufIDUkElnnHKor2YkmT5Bs9BGvLKdZQKUJ+k
1CuutJimgQ1ybx8LubMkyg4LUWYCWQo5A6US7lYMuuvlDxKCkJo49Tcuvk7lY1OK
Mtm/0xVqPt8xrwxVazMcCd4M1dZUfqaqgvjp68T44yQgX091c6/pM8kjCvQdkmGD
p5Ai7xusaUDjvHaRWgAP/TrvW0LVzfPUoxnlT9Boa8qK5nV7RNMoOApy7Yiv/U4t
+IISS+/7IEk0lu7p90BQRsEwX1D1jH6xJpwLmDxB4kMcw7dKxiIuHr02PrckpuNr
n9P5dKNOovAczyb8HcYvNMdR1pNjQWb0K9079mIEQWegD3FDsURT54mFS8uGkrXH
3TJmb44xnfKPKc2dz4XJ0XSBf8P2SiODxTegZKQ5bj9F3fR7fZaT1ERARMZ7TGaL
o122eZVexZhy1dpg3R2osVhdwqCblUnSX1xzEkVbnuxdU13ca9/mu160o/z5Ys+y
KgqLiuvZCDhDxkmFOyi5obYUpI52q+c5zIACV/joCruUdhCUFnMHEGl61jLIjErT
35DrFyyaYtSrZDfHytCHakMSlAfhP9YjDcHGfC9oLQQcaSwTIhgcileCal6UUFY2
b2Qu1m63qSLkMRKIzifw5PUSfqtyrhaVQb8sQCAfsiR5AFnQD2OBAokCUkYOGoPg
m6iP3aH1MrnSfDcPh9SUwkBnMoLqK6rlfjCWvO3NuwmM4vqh1xylfAIcvf66AQml
F1F+A3tjHi3CYl3rcMU+Ozt230IOREoQwyT46tYkw8vTxcq14DZrlD4rNv9nvyqG
lu2l5gvo1KVO+7JscO4AvqwH+s6X7ekkDbyK/XSpUQqCy5F5w5AgxKFTccwOeDvX
Os21ErQAUM2wFsRkkXP2S0hxcHhcbFplUPrBbiwKENf/04m842q7Ntll6mNxxo/y
34sIufimUyTAMOX+D6aaK63Whn+3Dw2cMwKbCzpLelg69T/Vvauq4J7enPsaKQRc
wz+8z8Cpo6c2IEfMKAy8LqsmJd2j49v+I1Zh9xBZ945BxC8Iozjkiq4b2hZZ411r
ZavB1dLaclkvcBojJiGUc5tJ8tApiQo2vLD8mzj74v7PpnTE20NfPuwQL73TkHc4
4+IRml1w51/DLO4vDNleJBMcyB+bQr+5QoC12C/ClEp3EdK1Xy3jcS/ip4E338CO
Qe8gAyxTi/4BHybIoolzZoIJ3e0QW5FLaeXLApJb+k9aNTDoiIXeBbuEruLRnV8Z
1mkm1a/FXMYCWlKMSDWwKKdwV+crJNKjqLn3SJnXWCWTM8FjfMRqsFhTq476j1yo
4oAJtC/LTklLKHgWiEV+50k0IqlNlwQeyD8OKRbjtA6YZLQkw7+1jklDa3briMAw
j+CIhrhpmeDwCL5i2PGiPBl6NS6Z6g1kXm7OiD9qmE5bcQl7zi8jkbgxV7yC6Mvg
ny7WOiK+AtNqZUIcIf8pKKHfGWy5Tqkm6lhVwYwGn/rz7bFcGwrZaN4AHKEysLO/
ugKX1hjRgXmDc3kJ5WPhVm1rMDGyV/vbsyW8QSu/XCoBgjtd4o4Fhln1amYwzXDa
/uNjlY6EvgjByo1/lGNPYIuOsZInOmyAbJgzf6MKPDAYgNolzke2grcH4ahjNdbg
iUZRVABT4N8/DTajtpDjt7d3tYxR441gIrSs3EznyyBNaGPV9wvD5pr8XCiMVgDX
LRcoyAO11GwaDwkAxVF4c2cwvL1U+Sj0wQM0++peIipxtix/+41+g1qqXl/6GEWg
As0oDrLdO8YP3qylYASygysu6fCxRgPlyV+hhj8sBksQwjhZlkwsmSDBLvkyk+be
RPr3p6Ri+E3MHGvATF4+EGQMV4nFcHEMBa+inMlgYfsS5ieHOijkN2+nt1RqWLQO
z/MAsR7o+IwMGJouOiNsalllbPa/VpDQG87F2ngS7g9DXkAcr0Gxz5Tk/hTkfTiM
K/Dpn0dKrv0PoMTbDMcJK9GHULL35Qu4paZuoGz2VP3wxrvHRAf9L8r7WFNDyo+8
wNgsyPB9Hj8DMlJddIGl8pk9xOPhISKf1I5kQq1I0DfjTiDqaiDv0cmVThfcJvgI
TsFS2+h6dhotArcptGVVnI5UFKxs8uiIulEOesCeQO4kqrhIAkIs37gSS1ZiUbHv
CJORLayhSH62w1/niTWbOGFb+FjpouKR0N5zIzmPjcZMtE6Q+nkTWeNXs5hgKYOh
Kds9rgv5Ex1J8WIeoYKiS5IqGbTnD+agVLEPijpdg1T0qEXEokPrpH0P+pBu8/Xv
Q9olgMvgUhm7ITZlHRBcCw6c7hOKw6blZ5su6HkxtOn6D6dhncIF9bveogjhA7Ox
MZvWfUwNst4v2Kotq4VkbT8JmjOwCqJ/hD2JbmbQ6qAf3IrLqzeZBmpVV8yJYAX5
HTN4Czl44cDG/9hP70XRvVm5LEk+ovW8ROOB5FK35tu9+KPBUB6CzYsWjLdbGlZe
eRKCx5Mt+YcaJb+R8qR0DDc5YmB3WCj4/u4dQYWRWS/ibkxua4I0NGbFh57uwOxG
`protect END_PROTECTED
