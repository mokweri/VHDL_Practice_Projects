`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/jX62/P/Zq/E2RPTbJViGICI9lgPE1GVEJ4m2Stmv28UZchzUVdoJuaVEqzs5O1
Yq16jdEwTcdpYjsODgUHehQ8zwoUvgNP5AGl67nWmHUgiBIbdfBdpUWOeWKWQ0hB
CnyHelWPcqUfHa6NPMl2xgbwNFCPNHjUToCLYNvOAd9em6dX1mDvJfnGl3mKHEx0
A45yKtnbgr/EYsaPCLpbRwc92eER0SieBTXIgujbm/wodYzZ6ZbaoWcqJ9e7aIGw
0L6s9lTr1Hpp/JaxgMAITqLu9tPKaovHtfx6b51RIYixMteLD0sv1ZtDgZrnWWQ3
ZIjIauCgxWIF8XrZk7VDQgMvxJZ1CfJwkrNNUrkZmu1g4brR5okOpm+Xc6bd7hLp
CWMVMEvXlS3mYLVfnlkP6ea1XYZJASJjyGRp0ELckm8C0ZKOw6Yv2uoi+kWcIT1e
iVAkI2Pv3KC4Fk/EMykZ+qpQVT/rBBXr5C6CbhkN/bLMYt7LhRHzddGl5Ti/QXrb
oEUiRUnDxXwRw/KyqslsQY1J2BFhHFVVXmQblCXa/1fxJi8/mZpnQjMgJ1bEsG+U
IyA100OFOS+3C/5J91yC9WFvy80Xx1ZjkEUZHzwTQJynIFYFhfa+z/OEGSKvFVxr
jNkgPKRaCpMjmtHYMEzRHv9wkwFN2RpD1zGh9r42g6x/NV3N0T08ODTVnnYN+x/+
XrpIaXP2q3fwfrWut99VV6G7d6UhHOjPqVyLZF1XM8hYQ19Kw1syJGL8eCuPJErT
axekfKAyngUnToEsaa72gzpmg86xsb9XwWalHxGEgPXwEnmtZNuD92oKJaIRXxUC
opokX3i85ROREx7smLMbQqsoRKio30TJ/b3a+XXqJ9N4YSoYrqVHhT9SqbY3cOLN
Lkckf/mEsTw8pWbR0BpcUh6AIv5XJhr+IhZ/enQFeBO+I/Qxi1jPV882CiFiVEaq
4xjxsW5rik+C7mbqf41JK65z7dAnNmZJrks0Y9QRwsX9gcyMiKjRRCsMsUQyc6pB
ZzalxoxD2JvNaHTG/NvH/5qSyGHdxJ0lioAoFtRgXZ4g4zwuu7FUgFd062svobu1
4ZW350mVYNhi4KUvblxnjfTf/zVKxiVDiUkjqGofmibE7CoXU39k/14RLvt004/5
miEjJOYGlMC3uyNWog4zwOU7Q8U52jF5JYsOBHaBAGWK/RrDqQ5kgGmnShx76bRt
iXwk4Ra+sd93YYjks+Eg79MabMYtWWJhF3NX4vBgNoA/yT2Rt7lbSttTru4OA7XX
WJEPwBcDTMX3Q7ePUsooWfr2l7fxN+/Ba8FWuutNXLv/YnxaxX9zNEGEQweE4pLT
8TMfiI46rnjM70JKjOrIMnX1h4sZtvmhbwBbYIfobEcFdm/1BRfUs7YLitm0JXp0
oNUSTquXlva8Nrri7wZOFsghXYxNoTaQucDcf11kxVRPeUerizv3OA9MPdZgZywL
MHdQlnUWorWdX+vCDJcJDjkRGboShTYXixshoIS6pAq2rIuGjW4IZ7z/KiJno6+n
rxat25Liwm8JcAmWMjsAyKy6AISaibJaY/r1F8aRWt0gIRhIlgD6Lsdhwq+t9C+Z
Nzk38v3XZehVBkDVSd9Pme9mp0SVe7uuGz0vGrlVUrM490qxmYddrIZOKjLYNnAa
+mNXt8aZ8AiVDsKqA/0uzuvWqIzJrEiCswIJtTiMSTy9AGsdKA/bUuaJiwGLI+kQ
kbKTlQJsrEAtV/8ZzLPWRePxJYArJIFnBxKldJ+CXWdZSHd6C0hdYXbnEAGqeXXs
HgH1OCGE3SN3ztbG+f9chGhO1ae1vAxB1tay9Hwi6mq/GPbogGXF8SWc3LiIDN4x
l1WErqQRu6I0vDSEy3QeLTTkvDpp7q9O6sveIepMJcxLoJ8w58iuiullybEkq4ti
BMatvPFyulKVJF8B3cNVQNnaiIAWwySIWlGBh6+piRyXgqNavlZBTuWs75utwJLP
okzzl+lG7yf7W5lAPu0ia7u4Lj4PgTglXcBlJkxJJEHzjbFROFAQFyTIT+fZnTJd
lxcNStApA5ngEgeoNTRpvDg5QTvYONOqbV7CRkPe0HRoZ+KIHRA/LWIC37A3TrLs
Rjaov+gYlKb9UJGGmIVS6ix58TsozTYoX56WsjneaZU3hvIPHdv9RglZ37vNMfWM
qfPjZKGdasbl4FDHP2EmvPp9pKAkQAYVOU2MxVa1ihdscgbRzYQFV6ZD2qme7wpB
k50m/0NI+NyNdiW5GNdeuioJPIpEVI5V6A0VT9tbTbrgv2ADA/ijuWF7kJdaK/s7
eMmkUEptQM0LETIkaPoM+cEGXiy+7O+ZgWVD1WUzamEjXfyNzX5Blfg3V9oVZJ6m
3UPSlc0lhZBBL/D0nSvaKotV34KtyDpVHfpfEagtIHm9GmTvvkObeNecoBpqKlEu
BZWXbuzrJX/uF2SMMpQUZ5RiCTXih1mA+J2mTzbw9lXd3TNz/IZfmWkOR6XkwBlH
9OYISp1jRZtgH8MljamJtrk/qBzoHtAek3PvksFpznvEhAMeH9sK9V5FkOIJLbOy
noRpiDh+inSpy3MU0WN0WiJVXWCB4HuxUcFuoQO2AzVbHuKSnwTcJ+o/dZGwlOpC
D7akCrxwsmii3FYt8A5v63mdC1bW3sJrQajNajyIW4XaNZxNyZwoyWjfcSqhkvp8
I3WW7bxz48Aw0KAdat8x8c/HGE2xIT0R5hywkRkQ4AMoIyyZRZ44x4/IoKlkatQb
KdkrJ0XQ/29itVXjk/LrnwiitJRT2HdQI8Kbr2CJ8azZZpCIHk3uNdtPbnXUb61P
a6nri4OPjCEFf5/X37782aaf5R8jIMrzaJkv28wYyX5bm4MaMqcrz7XVF1SzDwu1
2yvJz4q2R7bfWdNY/nS1dtJ+vokaDKOxUJfCNSPSbYRm2a3ta63v0sBj/uOaeUQQ
yYE5Kqu4kVxzNRDiUtctlfpOf792g9BBXnyGd8uJOgrDC0VkfDbB7dDoQH2lOez8
2mOf0c+Zpfa9bW8m5LiX0fZOR1UYCvCDbwdVmA4RZFQO7oh4AcGyeYQsyv5FBTkq
OHz6SO6qB6zlM5f8PyxDtdy2kvbntFyBCDb6id931cSvjCcQx+b8XjcDFys50fsN
mh9wZIwBmkn65sUwpQeN77xjd8r24ZPHuwv8/SRxxU8LBPHgCeG7t1K3fUfiWlu/
e3bexD7sLzqoKiGqCFL1ivGBNs+Vqnd08pQ/E9JLAiLgJxm5FEAUxg9i06opkUSW
+yrmUGpxSl9W4t4eWKJxv4u/8B6LwWYm9wl7qcBsXcG6Dc6j5B/cDirseB48Qtp+
lta/bqWs7lGGobEhzbmx31vYNJYDNeTQ+h40eZKMXqYf/OctsmDQj5CbPVM9+rAC
4Y5wI69NKl6jMkREFS3QGSM0Rt+9lP0M0VLbxf6oAe/N/L5eQUT9SN5c7qVNUf4q
Tw5qIWzrGbKi3kaOd20gIlaZ7/+OqlRxhsK6wTFPYZEKmQBdcAsStT8lA3m9yBbd
jU+OVQWK3mntYBlJHFX+hF0AkrmwF+FSPdlEEVbz0X4W8uR/nllXy/FzRhj7lItP
HMzq0ZmdOyxExU4Y0X7aw1nrX1zMnZHRjBiS2q6hNu8f00+Rmz6IH8d//FtVaHna
9eUyK7t1yUzFq2zNCIJuzFZxZ4OoUX5gTQiJ+PZp6kwRRQ6E9mpMX5Oft70ccjAH
p0oNW5Ge8sRIB+LHiOgQL9WeOx8VBlXLBdID/4kovx7kaDvArk5xMuQWGeuutsxO
KERrRw1J/r++ui4UFAr81KbTxjGFGXbQbW4V+EpeDNKnxHoRgyg1uyh31tcpWis4
duPvPxAO20M2UjB/yRBcXA4kfagmzLdFyNpoHHnVQzSAdzHPC9Xj7gCszumpx+4l
xYts0PeujGs8yzWHm4r1EQaN7hbNA9jUfiimv2oprzXiA7CDr5jiANKgfcqQjmNa
VwSRMwR6hnZJoeePDGyMS8qK1dM0HGT1XeH2K3T8f4QGe2S5LWql8oEuL4wYryAA
st22bONSLcn12rdEtV3l+twCi9vc3BPtHGSrP3zkBMaXEDaYweEPwD7m7zvc8G4c
VVgwTl/VKOla+GVaSOnjhwVZr4rUw6CcylTbYUzSK8Po8n3VTBAQG5Kd+PYdhZfy
/8lUBkThkWGy6kdFoC3aXjMujLFAg4YppupzZjsD1SXwfqBCuRyinxWAViTsbK0Z
OuXLOF+xXHlr8sPKeHYqbmxnj5GFNLTyamW5NxdYa3ELKxdGfngLzrPbfCWTO5/M
tOJYDtm0VhfXON7KyliYpXu5b50zXSPtMCWCA6OycW5vG9Bnro+/qHapK4jDwg16
KHWadfiuwzLyLS/HsHC3XXolfGeJ1clT7fVWxbIqs2H+sFdx/XlLfgVtSlSXGzhz
LNoB4knNTx+w05ttveLytcD7UBBdZj0X27YG/6sRZrPnfGxVde8WHHiQCE/X0yOJ
++ykmQaNfHk934O4B6BtYEnqU2OqCgoYyv8cSI+heKXDQccP5TV5T4qzZIuUuiiz
b5pnXApv1oD/6CkBy5RqICKhB1X9pizY4nfgsVxGe8Xv0VTM22RXJFRlXYmrZGxE
7gZDz5LkyZviMgeq6JyBqHw9oDyhQHadbfgBZ3LVhv0OzRAWnK9vABJ5U7HUtd+A
rY+QjVQOjXL4wEn1fBGEZM8wC2T99v9l54kBFf0+hjhpSmC7tXV7ohHfJwoGd3yb
HDiluGS91eCji7vlmX3UMcpxJ2vuqjxgJuRpiAO6CyieE47yGu8XzKLpZNKHIAsJ
2fYgOOFgmuCnYsSr1G53+ZK11X668XHeeVyD3hPsb92VnBxCj8pXYqO7MUC1wHBN
y/Rjwt7ZrUQuNBly+8YMhZBck4/YQEPCUxzkxu2o8480K9z7dfvHilp140fBv1uc
bcNIFHiR1L0lOoJAuB8dox6ieJVqKu2uGhU9em+83QGvBDl0sGQCJoT+kpqRsR4Y
6RQaXqBQoXysggP+VNR3KymZq13iaYcVjA4OLCe7OsT3f+A+GTcflh4JgEyQkkdm
GQ2XD8IJmwRUZQGe8XvVigiqk8ZxWdBWU23VKyo2si6uKTYiroCv5Dyg159uym7J
uowHZ2oZq5rb7i+McXbK20cV0Sl0NM39D25ohr0rrr++d3nSZ4o4Jsbm1cn1ayWG
6uB0lA8sL0+Vk7W1OYNWB45VGEU6qMoSbz2kYPSqFGudfgqprXg1ZxCpme8EFqpa
bxkj3FIsdxeXw08qwJeXZIBMJBuYnbzA/jO7E8C7RrbzIADZKLDH8rtif582ZBAN
uax4y0itonn4EG+1HI+DdnVEBaax47WJ1Ywh4ZVHnSo76gT0jkH+s/C71KS8+JPU
IIvt1DK3xY6au2GXHGXqS1V9D2GEI5NDWtsCcvgVUGTwLX+oFPBQznk7MHCS8E3T
V4NT50mVKzA/oTC9GOikHA==
`protect END_PROTECTED
