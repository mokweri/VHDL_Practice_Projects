`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MgmQSgHd9nadQ9k0dFdFVTjJn7vNjKI+cXLVaiozcD27zQz6ngF1mRbin092JtH+
ilIAoa8ddQ/HaJI33g5pgtQjHR5UVHZ/7H3dn9qQ5MCt88facDXBYqIb35oOOrSB
DOuR82iNx4gom9Rg5yy9Cvwz3H9lg1k5NNglhvF+rx5LEcaOIpdq1raLPxLlGJZK
UviK7uFpMjoeNJMB+h6Xo8A909OQ2Ti1O0LxIenL4DD35+HpHnaxRUV/q4VYRKKK
uyVUFtKIdedfR86y1who1ZDQu77ctS1N6G1FAEUH3YcTOmm7EbDhElDMwsiIUxOi
G4Np0JJIwsDVuUpT8YMkHYvJHOLT8+ArNtyxOYp7fJjutRo6bYHaX/KT60Jslhxx
46V3CckdnTojhIDA81V+VwD1ZIkucbeNYYbarR6acmBNk0kJnq6hjf+gP912cnQW
ytsKjgwFaWd+TmO5JLJb7b5DFtkKOQtxEJt3ZXWtV3cL2qKneXQbL9R4uUtRhkuv
xsfjv0cx/eRHzdgKVshbVjMnRlbMLLRAgRYuyO5ZRr2WKlTdk+AOwjY4FZtmp1/T
rxEt5AkK3vLvXi9n7B8fkuIJy0trKTmsSv9HrykIm0VrFaeu05Mk1oVkza/PpPNC
xqvPF/F1TyVqv/1p/v/NN8eNw1pXK1Thdd6yS3ypkzG8MWJ5i8jlAb2d1Oc9z1jm
UfR5bnpFN5vGKKt9ULS6El2e5ItrxiUFDWR5QtpyUarATcIrwrFKnMQFvv5Rot3y
KLtb5zAJO+MXKw+P7KwGvPeP6QU13YQwL5tw9KscCjep50YUkN24WdA5Imfs9AEs
UaWvNaI5Cxjw8deXbQO/PdIZmcmgZvcJSZSrCwVyD4s6U9d+4WxoQbAwCuWytCox
EDYxh/DVBaWY8TIwyQvCZ38lLRzxppw/n1fGH0HCjmwWzl9atp6SQXa70PzOhLEc
SxoMSb0t8i0Pi4sEdWiLyQlpaQC26mBYR5qMfiebfm0NtzZYiVaMDJFOl5piHo0v
/feYxAJFpeInxR3ZZuoqpPkJAmJsSLT3eHrkkk3IQqXA9cyRKvxkNHEuwdHl32Ip
gIfpxpssWZvaoHxYG4EhH8FXi82fMbyOHtipbhzvWDonsjipIuiz6XJNCDl5hCba
0heEhOITKUB+CumzLL3/cnY5sBmBx9UPZb5kXUGFl1Y7GC1QWiPSzV/LQxiI7vVh
73mjcChpqEZjfwqXDiknhI4r7HsV5EB/s7PN7cP1qkXXozyTPd/HOCkvhh3dHCCI
KAwKk9dqjLThJtSjuCdGUPKO2ktb6otSMC0mj6FKzCvgDUz/4OVmEwRMWmGz6l2u
bw1qPVzhkJM+FQgJE9g6w4TwHeWC3Na/YgOY+jQ4nM9ThQTSizLFK93aWWGVB2If
2TruTRVa9vnsLes4Wv/lzoKmmro8uON4zx0ot5KIhwnHnYpLEPgLlkTspx7IiFui
5emgNf6sEDJhx8vsQ1dskPR8CeVUAByeWbXFeWuc9PvB9JFQkGc5gpFiH+GQHhlD
H9P8q10LMYyKs5Hj1TTBiztVoHXe8DB5LOCyK8IqiBIKHkjjGFEMp41uW5A7FUhN
/+vUQeq9DaPBR2LZfzF476IgvkE1nQ57BVCdIK5efICSEHlClxWyYQeixbBmt++7
aJtenzALDgHPFcoegD9Rq7KctBvV2Whxg9zAC/1rh3rFAe7srBNUv/ynUhuRbMQM
WdXBWqX8IDa1UlXZa1A58Ma9Z42j9+WHv4k/xtAeZv9dlzNdjSDcJG9WuM1k9Y9J
NiWHUJjQGgL+z1xPz3stlQFjcHsZVcvDplyh3elTh+p7YkdiiSd/mHOvYX0nudiq
v/KwBAlsHPz3r4NqfiY/f1cOFys/vlxZaDd+gLzMKy4p1rEJ/HxD4vnlgR3BS2fj
fY2uXjW71avQwZBSnLxHcey/ELc6iL/pQVXn0yKcwAB0dsOFUxl3RlLkzSK7CINs
ZZJdq+et/Mw+BJgz4GpX9E/ECNmsyTLLQTltMU/BbLUFhKFC6oEr8Hh6aMIz7EHq
L+Mx2VqdCqxU6VkT45Wx6gc+DQ+GPGyDlZJ0ZIcPDrVKDjdQridTKtojqTAOg0QG
r1cGwJThngpdM/CAXO3BWINEHkpgdTRNMRwZHb9TPQJEIuKOshGlqvp2FL70wcIt
JYQrJNBxBF3Sd/rDsgIgrswcjHvZGAYdf9/ZGrpuPCSgxAEUzaWOO6nkEy+AIszQ
hTGLIr3RJTiWVcmuEffgJjPkMKB2+yAENLevMMWYVJvW1NcQpGBoLlXczsoqhVc4
MGnsMg53GzNBi8M9wRwywT7W8RaxVPoWOKDrfgL4tSP7dy692Zj8rpYEHlAIfqb0
TZltro59Mel0+kb14mz/Eo2/xSToAtVR30g02jemkqnkq2HAe/XnrDjy2M5+5LMG
JKINB8GFizpzwG77W5Qai7fMUkz3Dm8KHGCRjcldAE8w4GPYYvupcgmFTTjzA6wP
BkG6YlyUpzwVCXFYM+AYe4ydWQXt/VWXEcHVa+j73qikOOmybZ5KINW909abxTd+
vPmntvnRQ+Q62gXyzMGq+bkexCJjeGK7PuRDO7BaKsNaA19Oj3nZ0AiROh72oxCF
cd7mhLs1aPKptcKAL7x8ygtjhnBBQyb9XoNqx/RZ3MtZYftM0PWuTugadCZAb9yb
kSaUJP9sjUisEg/NglL4duDAcig+pATBEo2gfXqrZAJGIpN8FH7ywQxG1xc7Aj3L
aZxzPzBYLEOsA7yHOmNuBsr7X2ccFb3kjtWFqd5VtvCW1bfpIU2ooGznf9HkqL68
TPAgL0iJ4n8+6WsfzziNGyu5ZE2TeNn3bZr9JO9Q3Ss/L4glUnpsdMCxgyxBLurc
tvwoRCdXMqtqPhB9Ih3CzoqTwkYiJkaePK4WoB5C+ZJEFE1AT3qvYOak56N6GcLK
b5jmpy+zjhyxyxt7q/4ZzG8rHe/YtApgTAdyaL/q1QHhRk3d0QyAjGP0z3KgadLK
vh7w4akcim5SlIHp5ofm2nXd5XoFYTfkAHT7pSl6eGth62MvkXSQjTVycKsgzZnA
f9MqhNqPtVt4QeA5pvfZ7jl7jjYTgPUnhsfyucmhjs9jkp4BjpHvwqADCAwkRNU7
jXTvJLEnvW7voV5FE8PIuSdTUneLppRD6wgV5ag5K+wYA9Si8Y7oglk9NzUfSfYn
XjMsWXpoCjVwWfse1UQ4S1gRLLZCUHBQIo8VhfDsIckWWvrmvIsL/wVofoymI2Yc
tX3TDkivDNpRWna3e0abuc2Gt13Csk2wtvkkrlbkyF9HKIg3b4N/Qljdm6mUku/I
Eq7YPzfMZ/Ep/8y8Ec9oA4HUdTGkdzFj0xNQPUhYz3iWqyupEvU9rd3hsdVzeOGH
TIwjSGxp5H6KsjdJka6FrLxx+R2xPz9f/C7wm7iVnl4d7QREL9bSB5vxVqBzuxK6
9AY0VzMIixTVD+tSsK6dYXCK6AdjM9dZUE/d0Kjw26YYM2KmcDUlHol2THWetYt3
jz99iHKFIZI1HIN+Ggvdc2Np8TTR3nw/0yl05gjDJOnh73Oh7gyCo7MIDGsQymcm
1LVk677UcpSLX6vzTXO86EAobxIIFKSQjz1LdW6QtYjYoY1K3/2HitmDR3553Y91
+SGDdiKcBpTM1BHGtNe3OEPZh6BS2F/z2CmUVC9rJs4ctvbzVSz5nOHOZ2af7ZMl
1gchv0csQ0QijIIa7zUcD/wvg1kNzEsaN2oCUNnlnvLIJ3VKQtFDvXKnUYnxBB8o
9mP9V7gkkFBOndAlYtPLmOrNl0j4JTCxwdO7BeJ8FTT5yquM1B83jGBEmBZLENaC
cV9qGF+n1jGycMFceELrZw+/8rr0gZ0XuchpU1/uHEW1gGrV85RqOBzgqk3zuEJ1
Ojqu8/YaLyaElhPCFdDn6/LXChvQbHLEx3kyOHt5RoP6PCpdIrjhJuxYfimi4Ljg
lY3cbcnt3WaRTkRfeR76zQ8DCSzW50xKLa88te7IwQIqFG/1LBLhIJX/hA2bEE+k
d2DHWOfCMkX7i5YLCsISI9bxGfZpRHUyCLhaS253sHNTcDLT2BQRIWxOm7UMRFEq
p6jvAhqFOssb+LOUM6NleTWR4o5zWXvr6G5MMWg6h9yEb/K14+JoURsOQKYHzwM9
9qCE8CUMI7Bq5hTo230BoMXadnvdOD97MDJ5+xusQwYmd6o1aGZuXeRdMcdDFhza
/kk3VwCB930hu+4l41QDqpkz5lMQ/5BLVsQlB9yPdOAebIzFKZWV2r681mldkbXj
Wk6ZrSvHxVaxzaY4VpBDPYh32i4haNKKT39EPL/4bj39LF/96DBUNl5Y4RQCoGVg
EOF9ZC1sX6gr50iUuKY3DfyoIiRhWUWO+aQe+Dlxxvr5+eNWBeS6wtKFBOMwgYOm
3tSLWGoPsfXSVUN8o6NLTB4ser+HDiC7n94ri5hTKQUFA1o7vYQrucplSp9Nr36S
ZfFtVzMsL6oWSWizbrefWmw7f0Mj6BubHRY6TKKgILrH0ZoVtXjWES6abOVJsxOh
8t9qT60C8bSBvkFBAX6SixYsxa0Mv1va8eBp4TSeSD+mAbWmlq+BJBEMKcCShMY3
W6qLAeaa3mj1rTtgwJHOJz5CFnORL/q8kJCU3uWhDxp15n6HM0/kHpFm7h64uff0
4VJb86lcADAH//JLNEm77aqDGUjn6g4w/u98rJ6SiPrWtUnie8cqptg+Ib3LNUjS
Jmft8rq4o9wIvD5nNP9nNHVn3GED8Og5YdNxiqRU9BSRcEoguvowXWHZVA10XLbF
Li8qvPRvfcEO4XFBWjWGcgGm6UE0txwvR8AABwUnQqii8rfHBqcO1vdxQpye1G47
iGx7RwieBNZZQXcWygjRFk22SnrBXc0bSRgOu5i2UIAwQ3jwoxMC7bnQyt6rIDr3
JQuCZVLcuUK/gHPUE0Gbdy9apgJUd6KZNV/tWLBoH2r18qsSAnkqm1dbfI+WY/dJ
hc8OYemqW+GiSHf/e5YbPrursjbu0ZH1GODrNHAuORSi/MGtBMcgW4SKtQ1lxUTP
EcCWiRnFAxPJDH4HlO00p7BiVUllSnqAFhWpfhx8A/scz8wD0t6HzVRYFpuSphzv
J1O1QQ3k+A1oQ4PJGGJDtaNmPwwxfdyDXHCIQM2rDIjfnKt/yRGn/Q/g3vngeK2Q
5HaX2mSzgnRMaySjBqFHMbt+QZSfhl06rO/7+EF/ciAtb8WPCwHqgIzCzDFyK2On
OX1/wnbTZKT3TEBYGCnOT0M3MfrqkUIcLWuFRroJ/nvvz4Zz/RKn+oS5rsM+X2N5
ADIoE6Gn3BJTNU/xJcGVfo3nP3Za8CCnVTXd5dWRAnjz53LDIO3bm56xOycigUjg
Hw6LyVVuvPhlpiwNd0eWpUtL+aN16jP4VPjEZwe/7qJbHThJPHvgq0VJa5jEufEE
obiNTjuqMn7EKD5rUEYDh6l7apZxumRAsI0UFRKuy8QEuRKYXAh+kKRDZAlMLXO0
dn/V9D1UnFoLlmxU/u3qeVf1T0abVgLet/K/nYJ5z6QHWTb8Rcd24jcDmFnjn0v5
By0Wea/bF33xYiOKrbBTeO3vXAESunTEhtPRN1OrUHQ6PxlJ2f+Thh5OwjwLxG9F
ALktYZL1h7wSHfnEnFXCdNkN4/ifrTo+EdpXvTMZBMrp3t9HWjxt5oe2vjHXf7QR
uBCwrfUL81ao0yG0Zevx3BassgchC46Py8TEQrlsw5O0g9YqxdG2zr7/+NdnqUCF
P54Nlj6qVcoVJURtZ986Rpn5szJBzODfdEE7CtkSoyJpqtixNmvkDAbNfi4yZhvT
Ke8C8pQhd/O6xtufSgdHFvoOr+/9LcKhBM1sZI5ZsODh80E+BCS04y95uk24ABWT
OQpwRQEjZzGPEcDgkN0f/7UX8z8lRvC27sFqjR4hC09ZItYWAipzV9NnZOhnUFr2
QUiPREg/NS6swl3MFxBkkJE6J0/Y/nHxB89CPZtGvzOzf1e9dr/hm0EPIbvL8H66
3xfmbMciqr44u/1I+irj9kncAUCvXHCfvxNxsOOEObEzwgHNSakXpPx8H7iq7qht
mWnfJd99KObFP5Th/xpIG2SDNoOsymfk6o4PLmqN01q4vOmdSaVcFLrzaDM077WY
hAJao2My+SETMuhhKrpS9Gd0qBi4TH9DDHgxvDeYNBVLppwnWg5SiZpRlDah8STf
6w+XTZ+6mjJQHZqWKUsR2E12JuoatmLnx4DZCN1kuo06ZIJmgbj4eZSzblKzmg9n
KqyNKeJ3LZW5zplMoacJxCtfMgEtIe92Ne0IEux75oZ5+B2kC9PLXa3X9PWWQtwg
YhLJi6zJDE61BJkelXwpXaGsbqLDL1EjvYt8XjEglc6crybnLbAa5yib4Dnj4aAk
GCEWww26FG3ACuD8jgC3SdTiuTdNQBRZ1esVKOXgDBpRf/3EPDWGv/O6gAwe1fvX
DvqlosLeIreAT8AYjsvVeE21z/+nIqt6KcxHRSi4/Ux/q1HOjD/cVqGfD2z6ftyj
40Pi+UeZ3mhyhKZ9kQzzLH4+xHBfQ6Bm6WmkyjwEiFydwF4bkLI+x/ExvRwo2Ffd
Huwwsmki+gNialC5xOhIAwAS2GyGJOb0mLUsSxMvuoWICQs4svRUgMBRaLUg+vVK
4HZOGYoCC7keYAnjDoe5WvFSa6kj8sIONROWXvSTYiWVcF1RcoYBBdp7xmyk1Nn7
r7/ZGCPudErcpoIeMkbsoxALYpTpxHoamjg8gA1eHPOhdyT45ANBt2BM+dkAoBug
unTqbtMX2iKiABmTDBbyotKk0Aua1jNdZMY8rcyoosv8p9WyVDJ5+VpDdrKi4SVX
C3L3j92CUXf83UUU1Ukj48n9xdEnwsFjTWIcM59tcGtt45cGVFCfm8DFe3tqKhOg
qKDTGKAizmgYNdcppfDJfQeRrT645T2kH2iHXPSM6T9U0Q/OR+0dhPjm7DzZBW+H
F5wURHWh1AheIS0+YMyLIwAggfdG3BvRsvchE4kUuBc1FFgL+W5SaIKfbkRSLG6Z
3WDx53yHwnLPuslY1DNJpm8N/gD+e6wcEFVl5DragpV3K3dT2QyP1XC1psy6xGra
EUO6KntWoUhF1SRN3jHG4HYBoFb2drm3G+wDzIgv8vQVhdcVzrQGRtuThxZSpZZt
UDkpGEYI9qbnz0lODCto1ZzH4w5/Dqe9zymbtA/usGwJwfOgCfkMwLWyrpgOWLoI
tjan/fGbR6HAhupC1Nzm0JA2MnYqpMGGA37x6Nds8JNw6dwjbr5EN18FI7HHl8MJ
Tm0cGDNcUUJ4tpggSmMnig==
`protect END_PROTECTED
