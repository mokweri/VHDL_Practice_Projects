`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpJNpFL7N0aTyuxS1dV0A4XpWJpJTC/PG59YbpFKbJEkEEHrVXQn0klTXcuJNGLm
34tTeOjNv82aJAwn5s2DAneGrnKmmxk60zao70yYOpsU7Avxhhf41f5ZBYpagvyQ
3V+A5zft6LkoOWqZLwFMO2Dpw6lOk1rFiiS+u19OnQaKgYexMp9/knHs0YcVO+8d
M+5QafI1h6fs96k3MBSRdufEIOpjLc5wrb0BR3/tSqBOonWpyOS+9GZdJAorKsls
l4qrfR8dLQdG4OiWLSXHxTuWI6R0ZZ3sP+fcuzBaQzRZuhrVZmMe986q/U8iBoXM
8jWDpCkTZe09kyQyGTRC38W1z+O281sCdO1zaWrVcgNtXNXa2lJX70NImv9rC/bE
AvAylE0yH6g30c9tsM4c0PkJiRXx4DvFa/5tZ3CiIs9yz2Axhs9P8Q2k3VMrdjod
06wNfmgvANfpV3EYO2g40Hd413bsBHqQLSu3/c7R55olJa943OfEVTkbNfgjNJ9S
ol8z6dd2jrwEyCgowte4nW9PBAOxwm0nIp2NI39NWVw5NeTo437awcbrxjnL/SuC
RSQYnpkzPAEaUmqzzWnjGVLB2BNt8gBCeL8caF1M1j+5a8qvh8XQywRgS3O3zcND
G3CPr7m7d0UxWQLChblM/Q9e9gXGHuFQCLZpFB0lIsAEU4gjpJO7moF5ou9v/QG3
ZQTBSRfh9KoMg6NdEcsmXZLLGmODvuiIhHjL562uaFeRFiFCdXgx0aSwuJP0VA8l
RY1OmgeolXMKrWUHbheBg1TXdjEWrX22QWu68IHkZbC5NWWe87kKefrTo+iDWv49
ktaJzJglaOWEvR9gEHlE8qgrh+9NkYbJ8xZAsOnK8k7+0O7kD0CthZjNDkGc1diD
H9IuWsg9EWyeI4LiiTJlFdrVropMpEJNI8veAJQu60X8eQyCsJ7+91aWnDWkCluJ
z73Z2mCBRQatXnnSlkwHGd9jk8fRcKYg2yNGxg9GHk197CSnJUqHaTtFT3ScQVKt
p3aYtRunOku2Wumhf/nCSEkLs+hhDzF6uBeWjO5Zr7SmhKbc+UsAL+kEee+6NUtY
Jus2suPahi8tn2W69FbHdnHrs6PkBip4NwVjAzrZ1IOyij1tyT3VJCK3149ezsWR
nt9CdQqrrofCOkE6+dHda6V7arbXyJMeVDmdHb+tHMbC6XWwySUFaYdsOJq0/Amz
DCwsGdGfAWbTIqg7EAGRbkycEpns5y2gkl3eq/2KJ1uudhmBsNPzG3zRB7lx2S4r
dRUZE1XdGO7rb7hofGkqJXWFnq33zm4SgbhhYiGBXLnymSGPO5tPs00GreH//k63
nd2y+4Aep60Ha6t3h74P7X9iWqku69jgsxjEec9Bi7YRHTNPppGm4DL4fR+qOrN2
xoj9HCA0vYXk32D6H64PtwqFBGJ2X0VnF+IQ+/fL1egiQP5+5VyxImjsZCA/z8vE
mMn7DUaj86tTmqgWSS/2e8vm1p4djAkhUcZ6B5IJu5u/TdHHzeovl0v0dkMupjfB
945pSSxckuAfGR7BAgaxM0TfZ0fYAP5HpmynlRCgapIEZqTRnL+edINDNip8PXo3
XiPpNpH2acS3lWv0Spnr8qw+6t0TBHCuK9cRfBSz0QH4MU/K54ukrSSFARaAJyOu
4yh+SF1cjT6m3viUb1RdK9lQf6lP6ZT9QV3xk3hQDuF/ZoKRAeMHnFp8hjq4Z4kk
tAs3VQXGLbrXvFnQl+IEY6rQUulOP1WCTBTCnUZb1zAfVoTXebp0vEx4womHDqUx
B8I0CFxt2Z3bPOM4NALrFrwAvu/lAGTgp2IKaG60dO5S6ZyXWPbn3LZHVJBXR1Rl
6rCcu3/6gMlftYHaThMle+6Rp4j8WKdUe6Ek5TbZGUbvpH8KPLPe6syWRTMJhden
PHX4ZkaAkpIaYmpou97ogvYQxhNuiFRSNgyFf6eZu00AbvDIu8tp6Rve9v6cL+r/
GU6ZULicTEqRdFbn+OtSrb9SEdRkFxccIi1KQ3kEv2Q2JpTVa3sZgT0RRn9VtD0w
yKoZOyKPigcvEmFKWojaopURBKwzd4ito/Ttd3yXXmyr4v7NfvXHRMRcmjVnsoc4
t++pdk0bjz/KeoNt360fgcBzYiKzVgMoABFSq2c2crPdLqNuErn7ddSOQ8OsRCI2
lZmAjdAZgDkYPusT4fSFEqgAf5Cpwi9ljIKFbF23z6hvUh4EFAa4eRmDBPZtU3Kz
u3oeu0uRToxmEXxx7lKiiYLC+M4EtNOL52684wmTC2GdrFl9GACoHvsiIJ7h1Vsl
nHrRd5T3q/1Ervn5Nb/bZ7LF7Vwe8m6wEvpeo52TxV6rfbh3d1EGlOD4gRugU7x4
VwpM2w1scGEcBcGHiTkCXUkKBLiLBvMJ7GEoROWebGoUU/sMKwtpVtqi7Oo4dnUT
gHryu9K2n2uJVGdcuhQAZkBcY96MN19xrNdgQqL09m0lGl55qYRooeCCS+U9SucN
AvYtFghYqRxDIxoV+cRhgm9j0Yq2ZI7uaNxEJOQDYa6/PR/3R2Hsm2ebEQN/JthF
C8YUzFBfxiCZc1Bmuo2OwzDYqZ8/rYLJLHeTTiKLUvsdTHWV6Oks21hLPEJC9QGs
I0Vr/N60Jr8SmaY6AsojB4lJK8vkwlx7DIE5H7ayHlltEExDCD7/1IrAWSvRAnal
5Z6oy0ErbGD8KE4owhwdCfc2jQC++FzsXc2KSMGPM1nSJzRpLvgk23jdg+sdwyZX
kQ6wG8YPfhWv0F0xmHQQPsH3kZkwLPtLB3/uujF/QZx2XmMffZyWijOe2uQ+SnQW
ebZVrXaw028GktOy8qaWk0L0A9diF4VHevO6EdBHX3+Gw2VNHdlonopD5eXN0eNO
ueZC35evR7oj/4XQJaQtIlscwpRYwQVYwK0HZm9MlVheltnh68IrS3PILSiOPwHr
9Bk2wHPaTEJKpHADun4+fIXKC/Uj0pUXr8nihxzedgG1uYTnGvwbrnpf88XW5YyR
Pc0j3vk3tTDdYeaTvQSCbBkWMTDgwwQa+RrffnQd2XWJa93mrPP30A6SLyICvg8C
pHn9uwPVy/paOhozb3dfVhmQHiqFGBePvqCjUuGQ98beLtGIGyFLSF2xa6f6mabR
aM0O+vaCanlY/y9pzVq1MoRwmqQ+sMvlca7M6qkV6Z+RcQ5FO0epKLUR0tF3cYzE
GC8yF2ut0Zd1GNVg2EAgDZ0DLcydTNFt7EZZ4WEF5WF7qPHm206rixJ8pFzU4wzR
OScURYSuc/W4HStBm+u7fNeRkgBoFq77JWYPJ0cU8AN5LPd1kbxVDaIBtXn3t15u
lBvkM7daBx0CO9yIfSD9E71JQOowoVmrGxvIuJu7pmZJZVA8HpOrBCa8cZiePw65
7fHr+DYxBzh4iahPOTunT/z2rcmxziIXyG+h3RX+mB2aq+vP7YRaCiBRGpZ+TPwS
PzLnI5YtUn/1tOeHytD8vbqXXFDwPjAkDkEd8bRJ/zQAbNCNls0rAq1UcP0mDuVO
lWhpxF+HNdNhV4fPg+O6dNS4GB2HS9FV7uTbbCcWBQtbtYT26u1a4mkdBTiHkPzP
F6nB1EjshOCSqk/svwwxKyaAqILkFEbs33/yJUNvu9SrCBjhVCyDGiDClqlvFsNm
ZO0zDJnZGX8Dt1xKaLFq0/SRz5uPxB4uLzhg+HUpEzC+ROIyJm10x5hjTHsHQ9kJ
gQheA1qQd8cA7rSiP4yuXdoPBxIc1NB6RE5P1HWTEkQ9FERqNTBk/IH3nKCY9Agj
BuhqkMe0ooqyKNahEHzqXYOJdnEB4ZXwBUU7SH4jSq/I4TOJQw+vnEEa3LqBiyeE
scCNoG50FofVKa9KjmxU0AYh843MkXXqiDlY+7PmlakehcyDbNf1NY4uooN9Pbsa
ZovFWcY7wEIrArXp1VA/31TWrnEt4AGuThttQ6cTv2pzRdRwoKBUbjZtaZISiEcZ
dmLY9vEJ6rqIKqNLbGBA7+Htu72wbBxNwzjITXXpMv2d/htCDwRuySxxOXXxGLGN
u73vV6+Ts+i+CnfpEqO+k9q7b9/UBMepOjV0DeMo4/LY8sNEXYA+TyOu40KiL9iz
/itNjNYgmTzXKC+mLjwX7JHSn6fOIEbhlSVfaafNvXlBy1exjOty1S25LHKaz4Ug
8xKWzk/QGurN7k+TiEl/MLY7mtHUiyQarPQzErhIzhs7XAdYh/AzBqQtSEiWRPYb
tj0tAAu1WPttRblAjdIK2uoa+DwDijR9e63le0N7Q3hhrlFucwEF1xdCOZ2l6Ta1
Lmj0eB5YqLpOiO+MwhBDDJCuNdSv6ANxbYL6C/GQdWzvuqLuiDIsr3KQlMo1gakk
srxFdV2ty0CMpa60KBFabUwvHDn8OxvePmhRRcs3rCBvGWUGSCMUdooQWKyFEKPz
CCmq6MqOLadrlY9lgXq5bNxVkom5BdTgsRzY2YN1Lg51CaUcKjm6eNXUeiRZ76/k
JSu8OJ+cJibGDNUKv/rPkekZ2O/RrJbpaLH0ABHlnjuJemDTtXysq3VaM/ZnIPci
yDFNvZuWpzw1FDJgVkp8bmOE4QdNLo4zTkb0HtV4AYh9P1XdGZPL99O6F4QVupsM
rS6XG6ubksgAvP+ZtSbr2CRxw5xK5rlUssdyfKweS8Qi3IuZiTUnjj3X9QzpllCw
ujIZjBCbSnv3srTjWOtVLpjoeXxbZuOLs9qgvTFJnnZj3uib/zN2EpSjMuBvC2JX
uzHp714+JQfJZANjH8R9Qb/KTPljf12Vbhbiag+Qaqobaa5jmTIZNykyQ1gjAZ4Y
7a9Mg5VTFi+4Da/8tsXQL1GuLzankPq0a5f1Se6PTZmPPpna1onkp+LJRM81J/pi
zpEZJfKoiiqdK7aje3oF1EKUnjNnAqZ8DRQBE1211uUJqiPzdhI/7C4u3bNPpNkM
DSBxwoUCQSFMxpKghoyucKMSIO/Ez7YANsmEzzrAPyLY750LrQ18w6mlt2ocV9WF
+es4bLd1czeoisKBO/OkV9N0oI2+ZtmzK5QMYa6jjBVQWMdwwxpyo1lzwOz6+6gH
kSjY7l8dP0Mwu0KDqOnCC46cGVMfUwSDsbUCHC1Es3T3JvmwRLgloEqevTNPf9Zt
v1wCrfouP8cYl8wFZ7UyScj1hrDB0yCzzVRYMw+O+Y3zg3b4ZF7N3r+Bck0d42Pl
mOlzsBR7w6McfMjftsTf4ccSe8mpc9JYZ5A0p4MFcH0r88B8uXVkKcCHdElKRvUB
a4L9zkguniA1ZpIwKOqZRps5HqK9ur59T6deZCghQq54L6WL/h5pKGTAMdllWyAm
QMX0YLqDY6HNJbHgJLNwJL/9Bu3PacQtew6xu8wG1FnkBCKx5W0+pxlBca5/BJd/
VCDTIgjxF7TmL8cMKdjQiVhm6tc+LwuwirK+UnzG1bBK9IbD8+p1VcMLK33/xVR8
TU4bHXe2L2Y5tDiFFn0MFXUzNejiMQ6xZPYntBzSpZnkfgl8xMhQd08dKeYxTHwu
+d0ojs/b1vqnX7g5TYt1wL3bkf2Rkq+2xBSWuE2ZACPv57LMkikEs3+D/9ovqQaw
akkmvKARHD2osHN5WevOPOGiEsi4d/K60ki7IXCZhDBKc5d9muuhQU0SZ44AMe4K
I1SfP6+71X7lJSaOfsk7Kn92gWKtbahA4Gv9aHEpwBf5+C5TAL+ueRCKpeEz5MHn
smz/ZPzcZkGLZEeslb+BLjMwgg2i2VkxqG0E9zTv0POUwAIGG3A937wWZ8KGwtXj
r51jvvkG9wUurpIQ6ySuLJOX6bDwWZfdFCpd8H0uqr3vRsWpop9myClwXY/TJith
VDgEPTL/ApFB1R8qRWAXyuGF3qcEHwuyANACKHQmljyrfrujHya6tTZm1Ut2CFCZ
EN4iwsqZHrCXEwJjFgOeSi8zWVjXgUIOoemdY2yeFJV/ACZxYTNWpkTgdJDWjc9O
QNc+Ife4IYzIHLSOUh6dAfwibXKhCVpQ/Qe+zMzkI9pktqOcOzZvstztyshk0Rs8
XjBl2SCp4xJdOfivbWeoih7Jx4XTxSdop5OYzeWOPkqSqVKQirs+EY8c5g0xXNLd
jWiUdqDCMtg6jEoSylwGpDkH63oHd1Ql2hD4HLl4hgQJBmjvJav4oYI5lwp6cG/h
GaO5FzARiDqcuvYpdkRDCIWG6AsvPDq+nvuuIBGECLBcoE9Xh8AYxzgZENyeuYn/
OM54PKg9D9qZGTred8/9XvO/E8oY9+9xI+byp1Gl2q4Q8xmcS+VcPABId+qeNiXI
Fc8J6jHJjXkrX/abFqDdA0b2qKWfe9o9VFvSjTVcRk7A8caVk9WfFnh3I2VIoohG
TPYNr8ZZvbquBz41hY/XJ9etaUUKytzhkKclCjVypdcC4A/CnFE5mCttZpd0uPYh
JlQLWsfoY6OnNtQleeIGB/k78DySIT/jFd75M4/DXY/uv5vR2o4XZ5iDpnsARJiN
i9B6kUerJ6WbJOdj6llhijdRdJTziJEswnEE4ccrNAAaVf5sQDbPKRptOTYDt/Ly
Vv95tpCp11snfU2APWFIYFKN8KAEE60TMLDPm+MYyN7JttYdFHfDFAq7oXzYpo0d
KXC6HMKeOqeB4Sci6wrQiku7u7MY3ZA5hMjmeUy0utR8Xd6xJSNCSA0a9n0+GqJh
5MkWK2+Jvb6xG50ymNDUso1e3kHCADMX6KwyjR040pcSSCuVHbRAb/ythcNGxN2E
2jk+4a+v1W6R++a5S1xYmardfabPYEcjakS1Tm4rY02SfK+NQnVh8NIOBxWNenbM
2lcEEuXcWmXDj5Wax1sSrRCWHHWCMEXFEHJYiiBcmtN1Kw3tqGTblCUWNrxA5iZv
kdQouc6EyIdGdxfIRhBZFk73bqGDKev9wb5cmf677gFKCs1BiOr4ebzvddTI9xMb
9LkRLVPz4OI6zwEzz5dCk7YfpGN/M+8oXXCajxO0j4guvNS4hPQGArinF/v2yqwy
I8ouhWLphPgOLwPDBRhnJmVH+ePgsITouskHIulnAmSHsmPDPkNXFNPFAni+poFG
wYBKr41WdifDK1eRYph6gC/fEOr0Marb5JVVXMcm/yuKKkuLkxqDuxP6mbgua5jM
Bn6Wx58UkwF5bfcV38y4l7QhLMk/k1ZoUiPURSXpJk6p9LCcJKflR2N/vf6Rf3BO
r7/7XrJLVNWqnDYybj1TZm38ufHV0gCsyR/iCMJLaolP70yBCRzD5ratQyKYs+Sb
HZgeS32IFGZuOJEcWD9pq56i63UFV7gU1sNFzdzr/NgJVM4Qx5yrKfd199BYmJwh
GBMTidoy61dCIhZHdOwDwnmx9lkGrgjcRoP0BfHOyz1Hz9QnDaeoevEUZWKJ52VQ
xtbGvMUbmSE/sNvRhKubP+1m+eflTwaI0D0fLEj4PfzkFxOup6PyzvaPUCFX+MPa
EmbTQraEMjFWwb5v+sS4vxjnKDYeASoOVfS/D+/Q7gIEnk5RDz4G8ztKRQrQvHyh
Q3B07ZXl3r4zxu7CcCXLskxY2bj3fx5mN1sUdaS+K7hNwp4rsPPCGcFTUdmGDMnM
UPxFXCWgCnhydyvFUxIo3eZ6a+0XP7uAf2yijHSzgcBpRJdPQ0xs6y/cqjbdmlFS
heOwGIX1plOpEGplnjanhDAJ+yLoX98LBdx7FlCtUkEBkQkyBIgion17/LOQzaax
qNPJofW0oJ2ESg3zlU3QWKozVMRJNrqhWTQzd6N2aQQpBrncNchmifmx+kVxzRLH
9oxwzIrqsPQ17CDOkrLCJzpuio75ehWVZe3aXE8mUnjzaI/ul4rGBVIHg4jTqgMU
3dYaN3Y+Mn+1I/02Y4P8/zhpJiVmgjbA22S5NkEOCPavPTiHMb1+5ISKWSaqZJBE
fWrElBJJOQdJhCcsEJAlJzJfpZKyaJqfgD3i0WnPSabLA8/D2qjgRzzkuplJE5r5
sV4+btOy1Sx5FPrwcYE/nZuuJCVYCldgHTWiRGdzPie8L6yc5R6y78J1hOYHIcLw
tRq7MGbvJAmwndILjCFtC/BIxve/h+JqLijx7EAZT5oC+4oCD2Qt5Zmcdp3dJ3yW
bfjp5z6Ro8ihq/mmio3z15/BGSEE0QSBmO0S57/lhsQpwk/STzn6FJeRpyjG9wcP
RVEUJd0FANetlkdm8blbEqaqxZyuZLHEPVn1AA4Hty5l+bzLYgFWQhJO+mJYztDT
oEV86ohVgEWSVgKLFbilTsWrnBZMkKIk8NNeXUu/955MxJm4NsuMKf8tetJscK1+
EmIIqv2eF+XJdNNP/djuw16dqwdEgrkEq95E+OGUKLz+x1BOuufcO6YuPUJHYL1/
spaQ7zxPYSOsBSBts1BAXhWvo1MrZCVdcxSHs5JtI+jvld3bju21Q3ESydGmWQ+4
n8ZNld9SDXvsAhtF0SCavihJq998xtCiI8m38mTn9FdvUeiuaQFtS5b93tlk1thE
lgQyfEchIDfg14jaYnovEUtdTUR7BOrnGXMFOl/zE/HSOZY1EhclBLGiyNxnjQXd
MRqr0y1r/IVzCNC4S0oCzIu4qD2cQhCjQuAwxEwBqBheufzbWGcyrLDen9Msvqac
vp//D2BKh3Sm4yFVX5ANRVH0I73iCcIKNAI5yxBUXW7fOP1nVi/cUqWcWhpiz772
2mvog0FOc95uVayq1ZtBsIs3YR2m5k7a2G/JPzGrzj2l2Y8RHDB1nCqTuObx/Lm1
ccrUPorUQYsUFKAZpB2K11HfVfhysYNMg6hjOEDQWYNdYT/Bwbn5+1OqpkFekXIl
H8QG7QSTSQmw05Ktcv5HYTGOXoaDf4Wk0tMxm67aDwvWNdfoaQx0ELCZnUsGWlF7
oFcSHdRdcGHo8VFFx6RAACmgMMOKNGuCRAuM6UU87iHUK4LGu+WP7sqcSaKtgZzF
L0IngZcDXANNpSsrk942PEU1XFih5Opk9ZGZyNWjm/gd7i0/fIoM1uCu8P7ydoMX
zAFSn1fDyuFCE/Nl6is53xzVokmua+C8+MN1CnCjqyPMXMS8Fsw+dyhFiD2fTdFk
4+x/xRqGn28l6q84IvOv0F8VNCBnR4xLeGSOL90aQxHu1KEDsi/hASm0kbVD6O3u
8WIbL+e9/4cXuTlYHaD8QjT5HDToIZnDvQplEVlYF1niOg2dxjZiD4LCmKihCmgY
M2RZilddceVvmfaIBQeOTsywEriamDfL+oNpNcUhNZ59arJb9E65ay4urRq7iK7O
auikLRozOIdWPxLSzJKNhnEk9IxvCCNq5eWp7+utLdl/24lBrKwOQ/n/DXrGc6mn
5nbgmdUmXZUIoMsEqedvpP6+dHcvAepo5dHajjXgsxrg8S/hErfTvpw3TC46WeWG
itTsF4fzowFVwKDVtgB9BBS3B5610KVULXlSoRodbxrROy3PRXBv5a0B/xRnbcXs
/qRUIgf3tPU9klukKAyI/E26wgR68qyPzAsg+bOR40RBe8sJHxH1T9ccBg69iMHw
s0byM69ApUD6Jjy6lM4Nc7G93hw/Jz/qA0UzQgjbeDWgSOclfFYKDfF2jgEJNfL0
SjHxQHsK7L4flrhqDfQVi3nSrYulVoD+/wb2reXqvbBWAGu1AJduNtLLRIIPj2dJ
3bMcQtHqn7kddYS/Yh/cMzSaEpyxomUjWcwi/PcBMa7Bay3LQZfYc+Yuk0pvrc5Z
qNpmnLUkTkcAWwhoEITDdNcyfgnEfEiL5bLK2QXJh7AWsBYebhvqE2+CukyLGYh0
m/lr+LCESZm74dR2iVYeO60TE72A1a/+4st67sP1EX6T75OCWOtyz7A1PvLBqaBA
LJyZVENy80U2HnC/IYqAyDmpZ82B5PoPvfEfLOh+LZxWjt6FhW+Xow/GOW514WDm
sMHuSt7l+Wd9vJYkRGJ6imrQHVYBvftJ4QR6rU2Hod1GOqC8pPTUOUOisWtG8LDD
9f6Y80TSdYPaKhQteOVgMfWDr0C6aau0cg2RqulvrkoGi/78Vdk0JS0LreeB0AIv
gpVqSvZ++IBCFlq8US4nyhACKVeMKSniTfhu1R7mK2e1h3v9I87giXYZSMlbzZfy
9/3BnCWYNSIe8L6ljKc2aocpae+QYNQFwZ56OIOy3hrISfHqax/RGJOoRPu94El1
WHXy6Oe1zsuID8r92qZuo8Am5hYD7IkTOI+P56b1JmjkeF8S8R94D7nR+d8+wPFS
zBz1rVRyQV29MF5f+6zbHeh5dH2B2UvYN26iblNOjGDewgulTEPwuc9B+MpuW9+v
B8Bj8FKmHhdomBPBAtn7mVobpwtSRlVnKGBs17IBUefK+M/btj1KvbjSicyB0TYF
uBnPuQsnwpnMpF/7yH4Qz23NCw+4i3E3DguvW649ZnD/srl1BuslR4ukyNW0yOPS
EThr9mIw/vSPI1iKZPuZUH3tSjRJaweWfE+XfI0P8ttiFAlqLvwygabhqVViY2tF
txU10vuzBY5xiaIy+dAhPOb4YyO481lX3szVmq1pr9QlB3a6aaw52bH1+kgWKmKC
bOuG2v//wyEHcaO7O7339g9xjTOBkFCtnC1ALN+wRd8nhEXQ2HskEOpO0q+a+IWW
RljUCQbXMGw6jXYGqqeA73QNnRSJMLaacZNwjqyZEpFjV/NHZV7lxtOOXekitGFc
YtN6O7JjQMnZMY8TmSDSUCqBnZArkBRsK7lEYIXotYz3Kd2/IKA3t801gkt0UuGV
MvvIP4BRMy03Sr6GOFVxSzXtf1HhOOq2k98o+9dbdvnkbv60cigyv+eYBdYy5Cfo
JG4inVYf+QmG3BwkRvuCN4iP9bkcKzGOTvQmQGb9s/ISoYcPmSuKMcc4rXaRgRtH
gHvQ0YZvczYJlTMmV6KF3z4d+WQgFgc7GNQ7NLE8nvqgNx+WED8m9HLPW+8DHnGM
wbqIGw7dYqpXiRxcXrb3OmJosJO5sB923BpXiFe0/LBrJMD4Fi1oGlNjY7jO1Efx
l8z5JB0y+/FDeLbwVlVCHWjKODMtfesFdad4dkE5fjM+ry2HjW71ScXWi7yVlmga
fwMImIIremuI0n61JRpCgDtUGalSs7QjGH07kqER1O4bWdhFLDVUzf0h9yqB9GnL
kQILtTd3Kpa1/IVuHvwM1modUAaYN+jjiVsP2+NezqEiTKz5sTz4B7N28yt8YxZ1
tJ0XNn3PYMCtcPwojlYd0DxeaU/TV6ngsyrx8oMYL+vChxxAgwG9Nllsp51sRupo
4bf9uoqmTnyejKWXb6t8oUM0JWI5J2LPcyLU9qkXeSbVUvuXiOkg/LIEQH54X8d5
0dNv16Bq++K4eC2ovCXvAzob/jnKsLSvkK77fGXitPtSZbTDcsuj3VyKlVm+Uie2
yaXMoct5mDwWRA/nP4NuJ+Z2RUUGARgheNNsRLq5+r0THvptBF2dc3Xg1O5IO8tJ
2FPRU8E7b3f6kbbA4EtHxfZZG0W6lDI9pB912CrzLhHBOCgdn8/PxziWbhNnD3iH
AblCo3CY4Kn1Ud6HMQ7xie/OaC/p+wUuaaqAfyveBTGEU1JDROSYcx6dAXK60PWP
lZVG/Jul5Rp7HToQH/lhkNFKcbfo69Pkrqn7/VMs954RwBpJHs3cS8WPXNiPz/rz
bQbMOlZzijAM8mOAHD5ep2xfMvZCuuNcXaipy1OtXjzHdXvS/VXIIfBe59VnS4Zy
WW66bY8eCegvwMelRoWhu071WVmJiA+4YO0/ZW6y16sllwkvHoNNSnvV7vYEkLOp
fIFrGrdMQSW/9TFRyljy+4dm7NZuNGEKwk+C/fi9b0qa4hjW/7FppDx1vD9f436w
o9JgslhvIVKQPB8d4XOOmmwBCDfPHSUuTeTeTbykJHWR3q7ems6Dxia85qgf9m6u
3OwhsfTFS2EpYdNKtXBxS9P+kE3BpsErYHF89rAL40JvAtmzzdD/1823r7Weoh41
EUAQHgXHd6FbkhLk9JfLDADAa+as/PK+ya6mPMkikvlnC+VDRI1MJd35dItuVq2M
EMBsP/c0DvtzzwzMy9r3Yewgy5BmPPnl03Np7lOGobc1davIBBlxBuNBbXznaZEO
GiRmRWfPyDvwzzHIKhXcYA6vv+GwQ4cneH0pqlSAMxInLLG91OhhYqZh8jA+kvdL
jRMyf23AaLkRvDQ81JyBhuIwts5jV68OQXzMESNen4vnLfkyDoGf0zz5StmT7CO0
gRsAAwnCe2ghvYChHKM1CeDrXkJ58AQl41wX5lJZRuk3krxWGXCFYnBH9QK7CHr+
VWQ22TJ1CLkoehrm3OJXdsuJs/t3M2RuwNs0diR6J6QxaXxdcYyFzM2N1gVcSNrA
AgQKloCdy/1FdHnyhqoTATj1D0WBBJeeK05rSXGG+nSA7XBkdVMCe4+eIm2l1ReB
owmJhGt00uJCX7uP0VO7krL7kkVJGi5iToaNv4L1DJdafmxXJGv9AiYGCgbtTUIP
Uro/CLAkhwO2F3hgBekdpKJvr3DH5/1YBv/tbht3Y5oejFrxmJPYhelplz+nGQQI
QX0ctKSxNRswJQu6E3G6VM/9XCDPoNRq3RFYNCEwmCBdt1hMKxoe/bdgYX2QFRGa
BNbm0C1Emm0auzQZcRT4v1Xg+5DCy7IZnE/J2FatvaI0MvgF4MLvDuiAjsYguKx9
HyjTzPp/GkwxBibMrQH2iY/ruysPFdthSQhv9xN6FGgWENnXw/TWahDtDHC1QSOD
VepeLijAqPbq7EsUlFzzRsfq67c+8qbvR8jj/Zm0nlWufKlgm6YvnJwyNwSsvLMA
wHqEI5h9nhSUQ1AfKX6v1m1QLKrovGksIbNoeEl9bEkDSxK3aDwgwRIGAQKo95hy
LRCegC+tpRneDymW9zFlINn18CVZYrxItDKbd2+TWVjiDHX+ne156NR/QYgVXQuu
9KVGLLyC82+h6KDZwwOV33DTvwQsgAnEybCjCpkO5OzZo+Bkjh9ov1sOCs89IuHR
j4glk3+yRiAVgEM8BYAT1DEzWKT18AlQYj4V7E4EdQ87KJvnCapN4iXi2G9mAKoB
o3ra5H8ws2dzKajNkHSkJYAJ6B6F4ImXL/RUvvDpzUAXBCq3/AZ0UkdxFx89cWW1
UFKsj7+nYvM3KvHWh7qngSCy/C3tDF+up9f1OKvGUsJum7uZWr2FD/rZ3TDuBjhx
QNkQhiRtWoU0g3Y+Bczn1+ubDT/KcTwAxwHpw990XMRc22sHB5+QpCOc/bHN7mnq
qOvqZobAW6A6xJXszuI8h91gTebsGqM4dx7sc9x+vjLO+8DUiZfbQuD5TbAXSJkg
NtpjotHXnaAkcOrfGBVKthmFUb+5TTzGcUJQYyayLcRUkO8Jb+cu+WzJEaWvU1MO
BPhxxLaWqWw1P6BPlQXxAVb2vf2N2cUx2HpOmUWAuA0qfvsTE/LZwKSQYrLjwhq2
zwG95pPKpGEOK83KfTiHvdIlgHG/0qQdjYspKhOKSHitm1mSqX/kDByMb5glRB4u
5NJr/X9FOGPvGaI157+J3ekArQNzOqulVIJaxF8+WofB8vFpfyz1tykX5fxGUeff
86nL0h5KzOfgyBhXyqacIZz/OFCUhGS6ZxaLzj+1nKHI1lgbyTyqyoc5aJMTd1Cw
pV7wW18fE7TZBSHky5y4oMw072B9g0cTTeiKzlE0nojWRa0FoO4LWjbpR9oDCFGV
gx+Ngqq8iWp9BMtYGTWnOFVWJWwdKvK8yHVdfRvsBCuoHvdF6S7pDELDk+56TYMl
kwZb2qbDngd48x0rkGvjzwfTi9EKv8/68g6sJa3QSpoJocZ/wqkLbozAcep4ZffG
hSZSyvT6ywCkFv27ZgtSsKyBWXi6smMVAcDpsfgOJE4ppwTe/4Kzl/hzoey08Riw
Ju+X39bpIcN9fLMBplkyzjTWNSU5V1ySHKTQ6zvizyCmyy7WLN7BuMXY83i4dw7U
AmSE28o87NNREUJKmNQGV92SY9NojoP6JIc6FKfWQ8FV2DLzm89WYpnqfqeVnNrg
2BByznHT5AtlDfswdUUvh4rmr4dzrx1N4RGhKkP55L9YVP7zXHXqYaSdqk7Gx5oQ
Zj7LxeLOYREKkK+ASMJ40NjcxzhUros7J7pO/uvKEbBcvhIsQ1m0t5Ul2xedEZ8K
Hj3D4XjK15lf+KUqjvNv3cuft1LqS4M5zTVGxBXTX84IQrQV5B5QI6Rm1AsivTTw
XFKDxLyzGDWj/VenIbixkZsN1aoeVz71dTYAIxAhhERYQ7tq+hbTogfAFc8nrIH9
lluHzGp7Q1Dr6ZaV1uUagNPsCAQQ8Mh+i5nahRoZRkUaYFVwLlBULWfnytLbWJgR
lQqSAPxdpMkV9vEnrHbPMnU3Bm4Fb2/HTro3KG6Yo1NwfHs1D147q1TFJaHc3f8D
l2M+jXA4rA5I3Ag1xMnkUzL0DaWdkVR8sClBeirfOyAVElvf5GyFX/56LYSOQL5X
x5BYRviQTl8HTfSu4jhTXsKZsHf7y3IhjHUQyJ/1TrwrVIUXNgBU/NMW25/m/Edx
Zaah0fkGkI2tXgQ0eS5j6xHNatZ4yAC5vzJDROFZhiQt19SlQvmnsXsLtZzBV9ps
ZakhAIn0WNomolwNDQFmwuO+U1xW8QP3imRp4ADAHtVzZOPJ1PeAPcELgIbgw7UM
QrUFsjFCz7u8VC/bP+gOygQ1fELxg3774obuFk2f4tS91xVp+PeP9RTi1IsHkvm3
Z2q9S4UZKYX2VWpvuml6aRqlazkDygSOqZ17IAw6E1vLAbdf6RQPxjhpD4dJdNsY
5Jo9DarnCotTFf1cxgx7ZHWFo693+jyn840eGKHskwfpbTr/w7vJP3mqsJi37K+M
k7O9bw6UJf7MCViXLbW2YH22RrENzPUpMJZ9NX1HeMDzkipOCi5NQ68V4uaxlogA
lHBoCHO/pS7KxGfgWB8ZLvAvFQyhb04t5vDDDdsaWdchPLi/lyM2rSAm/U25J6/8
OUxkIbmYTpLthR9Wu71H0V2TQGHT13aMST/nT94gzeG/s/vRhO45MWwiv48e5b9v
NtHx5L8yOyg0l6eA+wPuch0kC6Rxgwi16t30sghQfG2ZdXlXxOTceHcnrhmCtUYw
MX10gvey+Mv0DeQF7YvCDP15asDKYjYz2NfdVn6AywIYKep6ukiLazyeP5VtAT/k
rtc8iHXqYNr3G6SiAXSnwWGD39GXJ5/gEVxKGMSQbBq+Pqf2DRf1Nymc22G0fhaa
jBXTnfXl5hJOhvbKAVHvTIx/0lisXE3urEw2wXimZc4JRgydtcxAujd2QZYArvW4
I89MJ1ZMZPhLcJeF4hLtywg8J9BMJjJzvP7AYlTVUwVh8xspSNODw3IdKD1LMEpu
ytjOrpUbiMTl1onV4ADFh6DeyOKfSV8MkscDEFNQwsExSUjAFEgqqvxSQvD2ELYR
pMyOS+kv6P2Bxwatv9fFHeVKh0ElQ0GlqDHLiXgZk6yaIbnrz50EG/mpgNE4xW2z
vNHE8T2BrMJchPMwx2BYvKRZeYGj7SwPjafIqtg2elyJTjoCuYIchQW2KaCl8WN9
n0VQJ5iPonG6QE7hLKB9AlyoBm+vNJfyawZtKexcK2LKbRyIsVUiOeVXxnB9qRFM
1QBpz5+y/evBI254poWaIbzNEqBUZBn9Q6FgYQkWOA6yPIJcZuNzvZLDJQFOfXeT
S3gpxTUjSX9tf0fscTAX8DZLXRue4GPjZvMMnRVATZStTxj8JuJ9wDSPpMIbfylj
zaCt7EoZgqh5EOIf0qdQf7Q4ZZR6zG2Tvz2bZHaMOJpzPDKVEt4xwN8kTe3nf1na
8FQcoFo7ofL1FArIze5d0nvPNmWU7wjf5WMsrFn96SPJRnc6B6pCWO7vLIw0ByeN
iGJLqKzxJOkxgpAg8burzYfdTdkquGPOpOmFd43qbCLGwS6JQt2gSIv1oW17ut7f
ZKtSc5ZUtP6Mx4NGBU42krEKg0nKMHYjC6f+vwOkHsPKz6/3+NEbN4iBVl7Ujrlj
8twRdcx1LcwfBBtXFmUueBTtIz35wJNSIKC8tmhLF+Y1bqorRSQOreihkW6CtZWh
R2GSl4atuvseWXWIcEnw0EJKqUI1fSd2REAynURXuRBCQRRMpWS2ErIVFlhJLsYr
lLCAIGfiX03srbb6BS/BBNEXu9+8yNc4NLQG85TCP99XDXoVVo2AvklfkQNgVHu/
SVYjlWL7YwqLnG3kpcma1Cg9EQ5YRZZy6ZZCxMeKq+3uC6Gs4NrggAczGuh119kC
2uSe4cfknlqRCaJTn86BasoB8W5uo40dhsNAnal+h5KJ7f0SfvkohqTJRBmMwhOj
gz2ngEjsQnJub9Q9/IQbVMV6SvEdbVOJ3eJ2apkuh3gkNcxDFpudJg1Fm+x2wDQ2
y6z9gqgdAyoWkVVlQsESW5POddlg4twRD9/DNLOamEsXjvJ8HM5R9jG9zusI2Np+
GOi6OYNc/HlQtBvylv7s4lvTZmGxUzOYNBNDuYKdWs9IN7j9vShuUJQ8c81eTfRp
KqDosoLkXjuJkMzkha0YGIYBpwKqZxWQzJPIlvu2emup/BIXjn9+iKYkDss4kZyf
kyfjb3QFVwU2CNP4LEAlw37jt+8jkdjQan9KaFLv3oi1/5RVy90B9NVEa44X6pRk
30awx6jV5qEvdJI3LsfIh44yU970NMcnCp+tZ74TFFHUEF1j9nreFNravdygRruV
tgc8k5kJxJ3EUjZh6Vspwi42ExHoRvyUDy/YGHqGE3s0yzVcbcmG9Oxt1sAN1uBG
1wvx/gA+nbPqigA+Updet+oWyvQVw3XTagjmPlOZjHusUCgfrqrjv5cT1btVQHav
sy2Dwlq11dYtA0R4U58zpzN9pwggu8CsCdsX5QPssxcR4cmAppg7ZEcLEbQ+CuEB
j2wXFiKiFQ/28xPGa+WGy9P22USsBBk+kSPtqxua4Cp7qX/LoXimvfpYpo9BRF1E
c0R1nkBGHSn6X9CMm7hShROg+s63PMkUXVVl9DRNrQhOKHIajbO40Th9a4oC2ODQ
o3uUAInI3bMgz1ipYxgIruO3mmD8KRofzBp7DTBbNpCj/fS86ubkay7d/v1dEamY
X3mledHwg0TXUOj3Zvv6XB689b/uXdJXB4cBD4YakF+k+n9ZvVsQVz7iz5REgLe1
SKQ/QkNWZ/0U1DcpGhjp/nCz22+yNV+/69PaLLUuFQBVuRp3tZkjb5i7L0s563DV
YDoh5EUw6El3e0XckhiYhYSDJ7Q5RDwaSYV8jDDDB4UtBO0Y5SiVPVmzxkgh5UjA
tLNKvYMjN4PSRUTetzM8BwdTAPVERP93U7jeQ+0o0a8gw5wQLOcx3Q9PkqMMHP66
dnH2q0nQ0rf4ZVs6/KKcdlhvovb0iXi7rd76ANOgGpc9aKQIZ/NKcAi55dXE/SB0
mxet+1a33d93Cmf9843/xq+n4Z3+hEKkInncS507KlWL0d1QFKzotOljXCJSyXji
hO9HKmCbinaZH7tGZ5RRGI3CDl1jvvbVJOziHIufK0D/lKPiVy2En11T7Irm86Ua
dViBrTi7g8EFOCGpGGooAdKhUR0J/t5WDQhImXcpdZ5PoiWT4W9jjGacmgqDMU9q
db2b0S3jLjju77WO5suJ+LsGVSSn9jlcjnyQ9aiiJd9S4Y3vnDKq6RE/31jfiwiI
wbE2aStH0bZeOEC3EHOH1isZJMnyq9AysDwBmdwvFcAKNL1x3du8LAEdjROyUzV/
QUExy3GAOnYZExKlnZFlkLe5kRMC2FTQEyAoOMf0FLyXw6Q98+GyujEXlgU958/0
LyxVCs7ezOhyzyaoczS4TNIzvLCCcv6fTawIP/tthQP1W2l77MtV7JppuwnblpXg
zwQavhJ6SEcC3GHKuN8URGn7oFQzoZm4IKMkrnY7xuPe3d976sBarF99dVMElpIr
8s/sqo43nre+KaMNLyswdlvnP50Rs5RZAGqriQa8Ty5fgAxV46TGzDd/sSoSU91x
aFPYbID0gvUHhlBBj2u+YZ/RxLFtDAFlfVHL3lHPWcqYfnm3wEca7JytlnRCt9WR
NLImkVZcO4RO8PCgpT11veUNIJMI2ZBIQdqAQuMKG+QjFGz6sZWCSXYTBpvjHBM0
rmYsjJgmedEmWlmmH4u5vsOGG80HeIi9RG8TjnpA//ukcrLH9Mm8aABfzfN4k8VT
JrZcq8VDYJDuRNGee82kdsDwphGneF8K7sPTBlu8eQJzU58/8lvWzGuzXI9C7Fbo
5UwJ0n9he9R+xODTHMZsRHhY2a+IG+WHvz5ExhpYWAMnYmG54NY0DkhjfyOaX7UZ
bSoTz8LXogq5CTdUo4U4IMIt83Ck9gx0H5PuQw49b5QX9lhewedq05C0FSJtR/ie
U5lq2aAWtO7u7hyA/88xw7GxOima9LLtqTcpdt8xt+6LCJW2qVitn1/f/5evRsAw
KPlAeiqndgW6y2xNFd4ZY86ZGFzO3FFMPPU3bTDZqO8mqWMPRq/AY0NJR33dmGgi
LlOLNhmhyjTcKj52/1fGpGmihNbnP1hkfDD1QSC5GSF3mXphFPbZ2Txz5YA9043m
3P/V0m8rMidpBm1/5AHRIS1a4WmtFQmQ6mMk+nLCFZtyA4JszdFiruueAxxXmQMJ
WwDHClaRI3HwE7zlMiZENidRZFU/nqP6r9cTLsAvv3Z2SaAcCjuTE05nkposx/N/
wZIcsoGCxKwE5F63m3bSGbBfClmFrafKrgFIqFVPGyGjn5fixLH4YD+deBmpj55R
f+ZomJwH9v+7D5IFMe7b8VxRyReHG63lL+2xmnbfvQ6A6nbPE+dpvzj26Y72z8uW
mSkhLCX8npWJPaPust4nffZAPvwJn9SEtzNIt+H7wl4hOLP41zH0a+ZAEXVjHUDn
5yhqVFKvk6Tr5k1EU7TR7UsPv648BCxKD6Vz51BuTNXo5or6qM+G7XrPzh1XkfXX
IIU/uldb4EBRsbQvKewgKf/zLWirEIrGHB0dyQJSizdax7Ts3eudm7u94RRY/bXf
CtZCAu78M06bE2CB8V8v5f6vYxvs8qskOnSg9QKDV+tSln5GX8dR52Efxii5pXMe
XlPq0VGxib2Y9iGxzhIUVWt8tF3z9/hXTxXI07DtgbdauMoWhS6webyAuetTs2Kb
0ijbrakHIeagTA2tR4F/SLFKztkql0Lit3kdK0ytc802OD3Fq1WI5cYyQMSIuHh3
pBmrsG8AIp8U0EMHkui1RSwDtG4HE3kVvcZODuaMUh1lA3Khiae6V82gJ0Yyjkqg
dWdRty7NUZN2J8FSy3ZY3GvJW2iRRN3mket2HYvL0JTcMGylHYl70K1KVRbCpeUM
GRN1wssGFrnPkOvmdrsOYUlN5Uz+V3yLyDHgAoJqI3Uw0jsiHSpcm9pmfwjsyDeY
8i1IJSpXOdrH5pD3NGWcNEHU3X0Q2qsMFHnbUvKesAORcK5kWG93ZVNvbYm/8mWg
ilTi3pUzkQGn6ybjoR4k+vi1l7X9xsB2nXm6WbmnLLVu+fFwPcdu2mhW7nHL/Zf/
KNOIVUkQLYzSdzuj4otjL32b1j/aTurrQK1d4QxYmCBCY5GkWc68MaMQO7za2kJy
AIYr5VQIgA+PZjY2P4vIlD3hMY032s/C7fqAh8kXqXwBgmJJVEMAWrf3Y6xat5UJ
aNbyJdrWU3pjxReNANPCfovxp+Nyrl6fECOPo7dXpDg/Lc6RVrw0kBHVb5Q5LnPO
ZcTpX0zUEe+/NRhOA/4FfQLefjV/WkTDX9gZHmsQoR464jERwBebGrr1noLfH8d5
iB//xdQ5eorJpbokzD2MsEgzHyDhj/fgk/k5eE/cfunTPJz1C7iY5YFEk+jiyhy7
41z1vGaYvgGa2CWFXgOhn/Nv5sGSBgGbJ8HL+etu+Zww3Tl/Exn8wFLqD7wEkFXs
PfBIbkV0b6mcDUBMawmXKeLcpB6hErLmXvU5ywufbTFDHlTI8E0P0/2WlexAE5VY
OFErr5tD6s1+71E3XdqjEvkSCQan8ykuCYN41+SFUoXAGTe/ktR/pDLp6B8FS8fQ
UbOegTvWsoPz/IT62jJVbYZOnoO6ml1etKpwPfDa1+r7CSf5G/sBWBqkb8ZeraoN
u2Yn8Broj8sba/cC91X9p4xc3llQzY2B3+y/eCy0LfGfrpM37LgPMIybIc9T1KZy
GBqpRdgzHFkIkh6DDKBvQ9CmoH4bfc+9M8xUnoh5eXzZ6ARrwfMaXNPGbjXcVa7o
ulXmnn6XuwTfW0RcF26BMaXu1gRPh7xx7vFzXSAQRgoF5jlZAzFGAIxYrwwkY2vK
0+FneBrP/gWA8VGV4w9UoGDC+DWEHGjuxyCV+lHcmoDepgHqRwTpcA0uQ69wEWOA
U/k1E1R+h62fdW3fAlI4wFQAJVHNtsKGMQhX7RF1kCzkMPC1GUWH4gGUt3OFj2Me
gbYCyaRq+TgYnhgNYZRW1usy5TXF+ZESuEZQk84gz8QZrR+AV3BhYanvo4tsmPPq
tNrdlXkqC5mUdY+dsdecs8f1fx0vLW0hhUAHKPOYp7pSBtFwuQqR4sBpZmTBzaOY
87bp4xn6cfus5QJEJtKAp9/P28Pjd5dmIoa28cVasO4mWJDdz0Q1WZTG3qUuL6ct
evWZMVHEWg9gSVYpqsl7SpajifqJODsnYgNoHehkzT/ER8OBPIety4mFJXjEqY4C
QxqlpscfBRm6Y/x60W9jB9mClAdVbzLhlTFPHVMjOBXVBUqH5vogBoK38fNcdzId
tUSaB7d4rdJC+DPMN1Yp5Hno45lkhLqO23wyF6oLECXdJO31ES7IZB/lwvv0jIhn
Czfi6rjdHUPwYxDYRMCe0fSezqVLhic4BEFLmfFdHDs13cDwJorWG1QgijDAVGUN
140YTNXkNzoOlFjtzhBNUiDs4HhGVK3ezKIGYU7wp/z1dHnfranKbpT8RgYmTK5S
3E89SA8JLItHTQL85Cavv0qq0nOxS0kmeGLUW4wgo2bYVrKgNrBygu8NyGT++AW8
gtYC9ABoqW4FpbWG+QfmPBcecrXym70deCn805JJOdB8nhnEecmmMEAM3QKX2bgI
H974EscmuhEvUME+8sZTmHZbERjfqOyJK98MBCYEjDT7TOcTeu+Uwbu3wNAyIgAc
uFBfhbw/jG7+vmnRzub7tPneD3sJ6wAryaYUi8z1pXfPvWnGflGzu4NCyrSn/U30
uzcJ82ZpzsjUmjYEdFO54ET0NgficEMJ9cr2idKCfgcJQZP9JXnACFeHzSxGER0C
yCY+huIK2xTIlUKgOgG1ED5Mx5SgP+cASQG0AKiXW3Dst+P532oAiM9nmuy3TA6x
BIxS54UYTOsByUhPP9uLoXK8SxzVRSHILdiicta7p6lwWxDUl8IFH+7rZwmWb90p
gSfzVX//x0KxSa92DHf3txCJx2fzYMEcdbAFXhDlQeab+Zbyav3zMzIjTumu6w4a
vE3JOU+saECWRRa9G9lU8MryZwlwhpPqxhSEz52YlNKcVPqkfhJT6RrU3ZDFhCQ+
BKChto9DiA4PrsRbrxqgERZ753gsfuQ5R2RaAe8Kzxno3xvLlNS1IPyDCBwE4nro
sTu0nMrD5vk2kQucPFVM5mnmbGiE7fIfFo2mfHmwuBCKex+BTUZuJAoq2Z+L1ki+
4L+/lsZ/gqrS8D4WDeAdBaI0fIsExJCYBEohtNJ+GMVGtaFglQnNcuSzg77CzzbJ
Yrbtcss4eOpLg7Udd1eQ0hRa5GU8bYEtscjyZfVwkdlrQA4J08f6DWfSMnE/NrTm
CRYjLo0oXKgP4NaHD5GcJebzCaNWwZy7oO2+0jkk15dmREDd6KloSv1YiB5p99D3
3wbCXG5EXSHMdFBZVb/6HRq3uQkDuqn52IGE3IhS11FN+r00rxh2/anoM/LXibGk
Lx8JyxYtRnNcmYCvP0RJuoz/HPMR/EinRkO29mGzeuIRIrjbL1KKsYoBgLEsnBkB
3+EyMwZWJnBkhqA4r5zB/JrKbvV8us4HG0sSs+fL/Ozqe4Kem8cpzy8f1CmfwviO
WHIU2NobA10A8jkZ0LmBWe5xxwn8fXI9M6SnRzw9TJlalEds1O3nVbA4GDqBB2LQ
vRTc6avSDvWgkqG/I8UPez/SFr6dU4NugGmcMm+YViy2Bnw1llB1RDLJV+5bK3PB
eCBBD1Ht/sRm+yQx0ILYMeqjGagzu4lDDqCLsv0lWS2Wsr/QtvIs4oxhinBeIQ4l
xvchTgf+L8K0N/3ADCu+EDLSZFa/j+Z4FYDio1YEuhxRaKF+dXTiOjEDUROFIVWb
vBkg5KYnH47s4e5ijj5d1RssJ9eWS366Y0vaEZW/wwJyVk1GtZnAvB+5bHe2qE/4
sIwtJMP1ukmyV63Jcp52Ea/6yGmLED8zZjSbZPPUcvPV9SsNV37Xcdejaaw2l8D3
qzPqrI3gaaNwtQgPOI3XXDGYb8fYAbSaqV7aqQ3PIc11eL614iX3n3zxT/oJ48X4
sJz3mCmb4zbJt0yAFSLWd/KweuwYDnd3f4QLFH/7VawsrSMTHqC7QBe1XwravVzy
5hm6O2qKBC/4aCunOrfS06sOq/brCx/wWB9s+kU2nlwU3yRE65eD9tOuINMfh9DQ
2rNUHVkaIeywMBpg2UTmQVCYFHWz4q4nkmBUbYMeG2SrQJKHDFSKmNTjI/3pfqr9
PbzNFqALMK/FGKJqcnZFC8/BmkI+798IQAN3hjvmSrrdmHnHQ7btJp2VpNLHToSR
qOC4xCQ+rJYQ1BybRn/QDB9+pWZm3GGLas/piqKyrtszvQjW/9lgLb7lfJPTeNRQ
IZ1aBM3R/3u4XzypiQ//lMjQutZJMud9F6stCtdMWPCO20vwC5Cb0vplULC+jjEQ
EoSfZfs5lV1GIcN4BurLWlt5C1Y6Zh6UaWX3VSYLSQY5y3O4437V28+PUgkw/6n4
xd8LjNpGdAO9M9DkNbYWz+Pbvx0lrkG4hkHdLzRoIldaFmLAZRnzuc3ivBYIazWd
jdSi/mAuQI8GLK1QmPOxXPquRA3ipvYW7KuAc01sg1CFDo3RaFOk0p1vwAnDR8st
UHqVDyLD5IGZOotPTuAa0upHhdrm+OW1zMcx5oYKC2mVxId5SFzUfQeW3Eg5M/xt
kWeGwU6isRKneTiMEDR+z/83ecT+M5GMQSl61Ay84kOEdTxeJCBFEqrAIENs981Z
CNgE0qCaU1hBEGfbwhgHPGJQc0WeUms3tuT/sLqgbS+T4PiaxXx2+4aQOP1mv412
Vmypr4GMMnVG6+vtAqQuPPFqjBF/Omrwhq2gxD6UUkQaoGqD/iRhkLTR4wsAO+7g
C2I9RIb51XlhmXH3UbwduutgSNvUKwz8BAh7aYEr+HjBzl3vtZkpmw9nFpfM+ixk
Aec1bCTWT5CZxSvdmiXXg2sHVOLwUXmp1CXy5qrphi5rkbbLMSTryuqqk3cStaRU
l/81hALImSIeWtKn56QePXzN3fEGZZE9mw2bu9RzUZki+bO5F4owIun6ovnBgqy4
+9H0tGNwyEr77a8H3y7swKaJhM4tL0nIHQ3dHJYBB/ruipPNaTlxA7pnFo9M1p4L
eKJ8oWC8TWUelyWah+Eij83DgQwgJX+PfBF9094CgfydqKqjnxMjl4+ajJoGZuwy
9GKgitfif9nF/zPnfTxTgsBO4dvpCyBBR3DWnrEuasbELcvsJIK8Zv6mb7IQLkbF
FdOLbd4w9uYIMjl6iG4RAw+9Ir8kUQM8zYCFM7/btBFqbVHxiF94rJ9p4W+3xVdl
VnrauIKt3BKBMQ1LxxuF1RxC8XvWwTj6VMpltxdzdLeiiYrt6H3OaybC0URGVnG1
sj2drC8cNkLrCdZYIqVvlK59TDyJRoLUohGEwNEpD/+zy2/Afuf42+DMXRmAo11n
JL/gPx4ONes4ixIo39s09f/2TguaEkWHS7iwtldmYX53KjZ17+BJiqRRNAeUWjLO
tuRs2c/RLOhoOsrwccvLwKFu8xFm5lwzlpTxp7RNHpzVvyy4w2USqTYE18kb7tpp
Gxz5xcFCvJaXChknqGw3eNc7X4D7XAKTmRgMqTzUSNRRwHv81uHF0YxSSGWZmlK3
UNBqoKUDURlMcU5vgjFlYRWQAj+bD8sBQU1ejWob2sisUe1mUF7p7fKFvTkkp4Kn
JnQvl4K+TvBkTir+ya4gIZGMmdLyuggfIzx2V8mTkzZz2RwA7RQLjDFejHkiwy4A
vtnD2M153U3+K2V7zFEbOSmnzLbuPp52Ehjz2uG+Va7AWl21a4/hPv0XxQP58PKe
RhW4fYcgfvnFsSXlJrzkL99YyIX084srzsgpWwqslCTRPuHbmyVeTCiGOS+UkDD3
1rI9pT7qtY+rHX3GMj03eeWyL6skCxZHkmX+dNhzKDfc2gJ/QL1Caqk+MUZJmWrl
FunWBSorlTmNLEc+VhA3KF6Jhex3KwKHAA1jceiL3b4nT5xiBv0xzcqjrJPOGQ+w
ybSTZNyQdzC3eEYnYpqs1S3Ar6vmtPz+PM6FSaOKbzLo8jypb0Mc6c/Q91cq7b1O
0tqbZK+D893r3seeMR2lGCu7zrEwOEpxhKiR+QMizHJMK/mvHzpRREGQGKix0B6A
nWQbl+f3Rzj7toxvF/F7tqQ/F9Vbpa/yBMBEZitrBpQQWQzzy2hQqDdc5xxN+jD6
lYrPzfrYy2bhGkjxz0uNcDghPVyECYIPGhR3EMqwzwc0cBvONBnLL4tDERhxZEV1
7onHvPNIRtpE2il2XIdXD4d1pZjX4QqXYSfa3AtNaXaKGnK0N09MywF5qWbHx+kY
uFH6uMXFW+q8fHfc0C5CTLm4BEyKEjgsOjXYHCL5MdC2QZKktgMgIqc5DtOnTHt2
ez8ZxXDhWTeua64n+8NEGWc5UJ2esKfvXG2orwd0stWUZgQyU9DT7wn8eOpUYYs1
F0KHWY3M57M4Il7Wl68nmvsCAlvQPzQiOyZADaOs3CHv2nwnbyGCLbBQ7za33TI9
LvoeqWlU1ZvviX2GVs9zZs4XjPYOsmA+ijyPY0PwR4sAWvLEdAeCfcVxLBF+eho2
7qa74YkEQnl3pvbzaLUJ/0YWOIBmBiWMyMcUP/Il80hcx0Z11CeYMpBjvLYVkCQ9
oqVNOnTHwLAhUMcrnjbtBq4L55G6m5bgwo+zI82M3nW61bzwx7EnJuKglhHK90bN
abhCwBeECcQ8ABRCsG7SU/MFJnmY4Dko3A7RDJvjWDUa5lStuP7kbjmBzWO4iLLo
9dOlW/f6VOoDV0E1rxreHh70w5UyCMvWoaTvJugFcE3etcVmVGBJt8q6DeFdZ2lx
Sh/9+aUqAAlv+wHgIZzOpRrSZltbMVameKYs9J+g4ySBQkPaNyEo8+usoxESoOwx
6d7N3XwOSU6r2/6tsFltI9jXhsnH45NijyNKRCoSCgVPndY+jFyStEn14FuU31xI
3G7B+C5mo1IbQ7B6yvZgcgFoxlCjSYWRKrAWJGOCKIE1MweQLliptgxLIkgoRcjl
Xwhzt2D6TmDCGW7X2d9vAq8rvZW+GPMBELnKRH7owF0XGPJrBpw9VAQ88UGRd+7x
qZp5I0FKslET5af27caoGLzmuKK7/6YPxa4OrQsbObpc99dNa71hZP41GDDBiM09
qLbFEx7kGNogNDyfHpxHN792631bWEnmy+MIPmPpoCUR//fM4XCUI5Jwa5U69LCi
5XjWeAZk/rIGLBgTBraOoXtNIx1MZq7c2Vk2FnDUTxA7+tUbJXdnDIEST/gVnX+5
vgjRDAbIiO9+zfGl53P7HIq8264DsKCbLXogXrrwl1Sudh0yr6Gj5bQlaooo2XZS
Mu96/KfneHjiuPpFb3Qu7/tWnd5Q5g231g0H1LOMr7cykifcZiTykq14Exfo88/2
XxR3gDmK0JYfD5TeZhKlFfxyJ7LvK2kZRI7wR4uLnNBuEUIXQmxIsz+y+ChElvWB
H0lHD+wTks7T8MYpKYEJ88qgYaAUcGohtQ8XHdV4FLqsMuOvi7H7Vi/+NydD0bWL
IPveFdP22x4toh4qB3CTn+4ZIRO/hupkwb8G+Eo36/wxERO2iyngf9XggSkeRTqF
VY83FcNOg90yEMNwy3+RZHTRSHRkyYjXs6k2SGmmtbik/8eGIqxL0Ro2Rq8+HupM
kfh1Wj3ezogoLIiiFR2a2GEBy978XSy4lx0nmsYs6sZQ4a3+a57pfG8xitwDlpW6
NuHikqwES/F9Q/OpdcfjRKG2eCY6zJpYz+awyBJYsDBW3hC6FkaO9v4FNhZlwlL4
h9T0nlzh202vxn8K8HJQyUxA5F5FYwEtkglwLTieeSezFKe0gzqHQxIOy289Q9FY
6jzvUuONkw6kzvLgpiQ++GIPSbBPZzM3EPKpxtuOt3OqwvYN9EJH0Ovaqg7k2u6L
ivhcxgh1dXHJosB5hRCTJWxoIld2sprtHVRTtxQVV0HKv1r9TrgLDjTvk+Ceb9cz
sRg+EhDl8f80iXzelimJUu4c/5e/k+huijD0W8eG2WvOqnw1X3HHB8KoaACNXSQq
lw3y/PvAEtg7f3hxr+BcvwaWMG4yDKPQ4Dbeos0phAdsejqaVS/2W59Af0oFaga+
pHZY+kxy6/O/UjSXdKLZxdlQLejMdkyhElDhMyKnJLDfkOnn9bxz9w+2Tb2Mq6Ub
EfX8uyrA4bJ+Cvc8cWeFF/D2DIcoDl/ICbVWN5WC4m4lyqZufcWfm2S9TCHPPpfb
vsKFMzBFZOLQpHw/hZc7JQ==
`protect END_PROTECTED
