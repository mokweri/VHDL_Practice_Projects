`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lX5l+YcaILGsAhsh50r9ZjCXsLfmWDbKeqh2YL8QiquXBrb4cZzV2QYqVdXCdE1r
9CZ6xG5xv4erx1haX3VxVjIRIyH+Uc3eLwv5ZzM7c0LrlRvX87OChW4AWz5k41X0
OYSh1NmycOPwCD6CtHAmx7hpe8ig1bvNLuDNGGElKwNkyxLfTcxSrKf/dt3XRXuq
P6aZmI8xR/J5+U8op1x+bLc/Y4oU1dkwxwl4BZYBAYi1GQoxgy9sPSf9tHid3xAp
PHuJVKm1YpTYnbOC6jG2l0oR5jXHUn7IeNxNg9exjvk8fmVNhkl1/9GC8L40qwq1
DhykiFyQ4DWzyhU6Q3ULTKA+nv1H6DcyMxAT+JO1JKtHHcpfSK3xWRwyq95it0iF
EkDyFn5n3mmAxSrZ2sCxxcjmGmG5rNm06buW1n1+l/RZ1AibZIg/+1m74mfxbqEs
PrlTaTI4nU0Taktg72sKrWPBihGg5v/lvIGt5A/2pQvsMWpB7Q/rCp+eOdgDt0oZ
Z2ggsSiM/Ra/VoPBG1cvO3WObWbO3N4B5MyjDR3K+Ea3B4LVM11fiQsQY/1cOzYl
0EADedhYMXHE4hMfUtPEWnOK23NRq+EDG6BaHd4rSvMqk+aCd7HPR7J82LIjKauP
FhlhaXkWBg5oEiIfDcZi/A7DEtpcqt8ieewyXYgwCE2iiixSjc6xSJoQWVzGVJ5R
fH81h7/aIPREbbVHj1FLiKgkOXOqBwWo8NnXBJsLyLbKNo9eyik2BA9FuQbi5Fvd
z9wP6xioi+3qpUzi1EuDwvzjxcd54C104HbN0oP8xTo26SDD6ot0sUkb3TH1MCnv
UgXLi2/50kFQJTOH+6rmORXPMkWG0X7+/fUkPRh9DlAZnGjw8OC4G8DSxfF6i+PF
8OcAxS7RxQ1t8dA9UDatluZB5xoO2pG1CInCoj+9UUI=
`protect END_PROTECTED
