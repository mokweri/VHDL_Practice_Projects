`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H0+81msntUMlQyhrOg2gXqgUOK0zXGHQmQqoCLmCi7FtNrdTQWA2X91YKC3C6FPc
lxk5fBnesWNeYqri5hQveSTdKodtdnYBN0mVTqkgbFkoSpV6UjPoKUz5lCJmSej/
d9W2C6mvxwTejpcHwLfxIM+dQJlh/khOXqV2wXLN441IGN44f0Dg8Il0AJAlWpeQ
6JYnp9YR9DYfsM7fqaxja+6eF42RUe0jFBrUuaQsIwXTCWwj1iI3kKi0D6FrsiDx
hrdxI0muUjaF2iyBbR7qElZGyl6Kh/3rlRltW8ucH7sSkXgQBLktrWqZ3rGQO/XU
SrC9/kvBwOed0iv6ZrS96a1loiPs3k0zjwxSl8WmG/iQSgrlboTXS9699hVXxt+F
NONG0pIrFf7J/k1BKW01uF2KOCYGxb1RSqPLhrQ2pnw3zxhifS1kPAfr4f1eQL38
B0XKf/BNURXZrbSNCe542fAgNQ6t6//R3YxybnQzsBupQVcFoTf3RTrcULfnxHb3
k2HqGKxKZj7J/d8R/5caJKsqG7OdbjbyulyxbVwTB3mrv8qhRtAXIou/DjSp0erf
RfGZE2KbZF+zpTQtdWGfOwYXNMF5xOBEKqOiTN6ePvOSbuLpGwyjk450Sc1BlRj9
o7dSwkNPTmL6G56bVSmVX+cY7A76gs0jYsB2EGX0n+dgdez+qSNUvsJkjhZ24Q9M
exzTL7fNjukg+9GYpRqOrPPR3NA1AzEkR8fVGMGRMgCqwHbIYZvlAOu82kIci+Fk
/XJDRgir8oakplTExLD7OAGwrSOUPtkMrUUqUJD48PTF5HyuNIfnppvnuN/s1yBF
cL5DeuZCecfgbTlsEM7vOZiNlPxgKBINtvLJjBonfve0SXYVaSL8U4FN/dnd9dc5
1sj+FayZW1VLuNkhyD380ZtbzF2YdIbdCzIJQm9gwIZG/KqTNkIA0AVsTPs+hzRL
lo2h8yGn7GkD7GrrX/JJ9h7GO6NH4wfm4COuzIr+Rxz+QG+mW8rYtrbmCulQsmi0
l7gqh6rjQ4hUcI9nPmNIDa1nHY+qJPysp4+DUtjb9jker0tgM0Q85gxEMnIstd80
K6AF/TR7grHYpIkt8Y6QAfcMGZ+u3oCQwDNB9l03GGdig05otQA5KlhmqCY86C0J
W6RpthHY0G9SUGreM+6NMqv0HUr67+vMEhUEM+9Xp3bchAhddNNy7SI2afjQlkCR
k/MBm8XKPxedV9m7RDl90Vw5oP0ONMXa0zzQgDRotwnvX/NEjQikHWSNUq5OYS4V
0jzQ2LLgz0ffcJ6NGfMTbPAjsOKKtM2zRQSHG7ZVGzrlp8iTIDGCzfuH/ErWWMHB
nz8xR3UkQawPU4NftS/6Soz/kOf5aQPtAUMoBE3YldSxIf6O25ldvT3cjQnhcQFD
ecjB3dF2oCv3Xi9OKtyuHSddEMiqlocJeQg/vhCBZgcQaTq2F1FWACONdjCDzCIH
Pvq+cRoycrJWpqCo+GMxlbTSHyToS/hR39Si/VPWgIiiXykVx++Ju6Nr9+NzHt/0
28OtMt+nXuqSdD76+M1GdeaaGH7xFduVd4uZf3jVV5ZCJCVLCsh+3RQugfLgSIbS
hKJ7Hvq14/8nGxYRdpmYwVrMub4UVuIwgzyohoSLKvreSl+EO2FMPxUaH0yDgbVU
xVmAE531jpFx0BMMehZg3uDB4bXt3IomeUT68eyW8c8OjqM5vAoquyZ77im3W9S+
XP5WZmeMZDaLyDP3xST0hQ==
`protect END_PROTECTED
