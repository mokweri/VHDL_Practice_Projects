`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oin0/MdBkTKQCXYzBnZuolP2/281/2U4y8EQh84HOd6UR1op3jPQAbhxUSKJNQQ7
JHLNHBOhLLMLI+4DkSIKtJ1t+qp+9BNWgRhuDDWTM5LCF376Rl+4q1mlY9KCiAaz
LnqZ2/Pj+TrVQWFmVvVGNCpBSeGKxOHXNxyv3h5UqhuH7Pae49HisesP/9K+/JXQ
GM6I9tnSs46UwxKhGc62F5C5SZv2ybf4gR0nX2L7HTfQMqMgx1B2hfHU69qMwuZG
pZdxRFdwLKaDVVRzMdQp2x5fg1kkad6ULL6EelxXaNforwC8uI6EU10iFxquqIfY
YxYsVfmN/zeiciWS9dY3lDqnDZNvtGOr0wX0LQmNHOXKgmnv273PMxZIDz06HBV/
v7ZHigpSDLOHoCFOJwdGFXGQC4KzkmCdcxb0+Vc+OT9p40YRyoipv4Qcdj9MedMx
9YJaTbtxIWdXsF+/R58YnzlcBpWyGxEwVh2gQ86EpV9oYJHxES7kMvibu43rsQsV
GUJMu0siggexgyqzVWKhlSDwwHAOyDTRvHgDPkyn4P1Me3b7wXlt3MrP6UT+yO8w
eh//Guhum9Idk+Wsrzc4kBY615d3nIAGkYYnIphOMPsCOM73q7PtDAo2kp7JfvH9
06CDkoYFzOTqHeV2nkdNsmu5G8ENzJ/i0Wxl+7SnVjZxtoyxZLaojho4+DlpK7IC
MlMKIt3ciLPuOgFYdPvKYmfLZGo4D1cPwOVy/gu4wQodABWydsyoeIp78Ik77xuI
vwWnxKhIJcg6MJrAq8028o7j7I/AwlFMbG/krxMyJWpEjmuedaP+Nivz7BUfQyha
go6h/g8FXpJww2vjv36rK7+AgDJ488QrORjTjcfUMbxCpvKAgkaFdYmHtLRUVcrj
Va4U/3DU6xBifnPt3Vz2Viy5nzIkSzZR07G7Phd8vNNSCirGl8MhfM1sxPwFk2/l
F7S6v683zMTahYMkOeRWHJeizoeAf0+3GfDOp6knaRpVu4ueuAmaLtOE/9DFG12G
Qi5Z6tjFm9wAbMqm4a3Dce6MhoOvWn43RWxpxYJjsuJNM4z+EuIqffIoyvYpVTYl
1MYs+LnIjryYh3yoPW2PxzWFqt49KNwftNZE1zUd0nP4xFpnxS7l/2CyLRsKXLr2
peA3xhVTYHSqiDARwm0A4nw5QVsQ99fH52AZkKaLWrOwL5JEtGVzP8yYbnmduxQ/
EUF6IyzSCFoUaKexOg2PqQqs4AW0JQmjQ2+eQBGIBSbbYNjdGv5T2uSyEYtcBMJa
KXBA/NOnzIbKioWjvJfnXV5LuIQxY/kM6r3oF2SrZ1Aybn1/LXyA0cCTGZV4UTfO
Wi7BXZC1fIFkYOtdUoV+rYTsOwO9DwBOC3QG8CcBUMCpvdOzGt5qQPR/j4R2+rn/
NudbwbIRIObPtIecSzGDd9MmiBHe3R1pGh9fB4NJU10oV+svMNQOCgG2HHTPBwDR
rvCzMNmUrn7PgVoOvSIKe/xG7moohgvKrIkXheMdmG7LquGI43EBNUJsYnixXNKa
3vYSbIP07uKK3sV5XN+31vfKw8SOq70yclpsYApODmpxbzbevHsEtTUvT/agQFuu
K9ZfCPQdCtwwZxB9eT9ElUW8ITZwWoQhKvXgCgJGdwM=
`protect END_PROTECTED
