`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PMeVeY4FgO6P9KS5Btmu7fKUsEV4mjhUt95ZF0Gz5cTgM4uohuyf7DZtpBfIAejG
zFVyRjHJCDiB7sHhwOw98s/vBdI11b6PBehOj/kkFArKDmh08GoAfJ+Lt5enkFQc
E5Z4cj+UJ5FGTKYopnJefoj7VW6nDMpfEFZpmG1HIsKAFfqeBpeIh/3RYvuhdrTv
s/HNkm2syavjkdT5dzKYClRD+GW2xWGvMD/sIGXcIffuP4RENqmumUbLIPS6NYTn
4vEK/+QC52J26BWDDdGc3rRSp55L4ttsTzJbVJddcpGEVFBMTFspQx6Z1qePXPV7
yMdvK8aS7YZKuTeY5PvMxfiBhM4tZRW3NpCCwM0S+qWbx70X47se65MnzGauM0JQ
jBU3NDM4B1Am/I9QQTJluEuFUtrohIqHy/ZtV+3JEmI2z/R1Gsr23f4LWIeAdI3q
xokGN9RjFUYkDjySGNAjvIHb0mHgHd1iX63SB/ArksgvS1G9ywBPOn0oEtAsGMRy
Kacx4N6osrS0jeKCizlpxJ1gKv2fkYT60bvJVJXqepJ6j0/qA/5N6kfa58z+Jm/o
BJqL6uhBR6gpotkxMsnxkcvGbq58GO9FoFc9aZiUA2aTExQ9ZlY8X3v0sYiOF8i6
AIl+B1GCnF3/7hRIrrTx339CHAeHaxM3iip72w/j11mhReDLmPfAO0fVomj6eUJ0
sPG63ujJWA6jWVTmi4NEys7b7ATKVh/is5jNwn1In+Mclv2vo1wyiBepzTkbffRh
uTXwa2kEfz3xsIcYEIDLSyJaHHn1eZ5vu5lAgWoeUpS4EU0lLPFsJmQSo2ykJoNh
DnymGwrJPaHwDXoP8sBDyd5BHNuKV02P8d0Z+tORuAw=
`protect END_PROTECTED
