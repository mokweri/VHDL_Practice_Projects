`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0neehC6JqGVXjY2n5KcJtiYj4XDKAbMVzVg9SuvLBwGatUO1JHQdmQHIJ0q4W3V9
RgkZLet2nX+sTsUKGwYaKl5AtGBjbejYopQsAH+zjuHehG0BazXDEGJyXJq3IV+i
wGdIOUfYmnnYgZtf+AluPrjcro4JehkXc91m0cL1nXqEW5zffMLGaaC8NBJjUhZV
6r6f3bRoIAINDs/09E1bFku5TM3a8YG4pIZHcJYYu6iLYGWQDOGan550pxU+hnqi
5VPvv2OyEoi1lgQUM0qevW9XQUcsjeJn5TIOm484KQGRF1jfykGcxTwtF9Q8E5AB
t/JfxTmBbP0b6PtRzxvNYiF/bheX9jTpJDmSkjxARLy07pC10+r0jmpnxMB/TUq5
`protect END_PROTECTED
