`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xu+CRWfyW+3G0ZAhhkU+e79oGEYa4x/yunuKDbOh1nPW1RV5K9widx44fnXJRdBG
ajTV+BnEvSQnXSn7isLd6HKKgmQtsCK0+f1KKPLSbODBFVD7cWjPec3g9S2Z/7BH
6TBdOwIMAvU3wn4OShcOj+dpZ50QWGsrbiD9fZs74AALVCpNGnacZ1B06Zj7bw8a
`protect END_PROTECTED
