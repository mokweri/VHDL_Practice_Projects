`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItHsi2JT+jZc3FfK/hsFcrpHLeisVb+GfivpAGyeuZmze4WprKgmpWnKKQOZzZH5
NGIPvnoSqg/uGaZ0TUyk9gi8YeT5A1RMYfTa4KttKVqEZF0Gd3rmOilm3ydpj4Jt
hZNm0ooD5ozvZVkH1D3ZVkoQCv6XliE6L2W0QVjIldF0Al4FAFf3iGHvNiQhdROC
TbJF7YQ62baJja4RkidfRxLiAwBnXtJdd75k+0H+yXoTZNPeVqtGQK/Exk9YRYK/
3a+ftTelvovhvwgmbfIG+mXM9MGMAido1hzXgLGgmznU1DZid8wkxeRv4O4k/934
jnkk/drQH8rF1hbpWbdBKmryAQvkPHER3GGd19m9009DLsCExF6sxArQRK8Zj1ut
U8XClTAfBs7OmG510qF7KNXOXocJZEqXdZGRcvZi4ZFtl7bEQnqswcKrd37KEKRI
+aBcvY5+xuq0cr3Bleu4MH+56okPmnf907UTXoiUy8RjiiEap/iW6TdaAaabRHa7
+BBPGYeGGtnCP/LrqLrU2l+nDadEKBdCSh+EbVSC9TjYPdBPGxPW7/9DpvcBuv+z
8+2qT4faPdkQA6M5ToQe8vIdIZVvYlkzWRYLNsnChuFCfpMEsfcpRoC9JYouaU1+
B9IEOwlJq8N6MlrLAfEEzvAMULPCS1Uu6e5ztwjiCq5bX50zIzqtAA74eAQIRxk9
v4FqNK/bu7YwJGcOGE73wb+UT/nPO85bFYnF4vgh14yUPBnZbCTTb43Fl2sNRaHN
kir5/UJ6bdD8isI7g3b8PTgAJBnemDXn3nbUnMMimtKuRTfetxxb3pFevmIZPDH2
UObAkzG/Lva9nNX/YdxZCRaw7JiBULdS4J5btDyIf9XL+fD4GziPCGDhN6UOO0od
V3lhvrAPB4S/n8Vs/OZwYQn7PnqbsECHV5dX/IkSV8YhUUrLmpemzJDjxiynytUT
4W7LND3cLL9BgNzEWiAkpc320OxddrO9vtNGuD9VQjPxrU7qSVM8Rty2Bvxe9com
SwI1j84B3UimKGk3hdo6PTUtBhBH8AmPnjGVdGsYkp9inojlgbFax4MNo6bqi+D/
br/sk3XwRTamdzXGb+/c3Af3eECuXFaxbfZI0n0FCORIBxbI7ociX07SidXottE8
8RV5U51sKge9NzV0jEPuCsHYdGbCEEhyhWZ0VghUYuBh0jfmiFM4gkT2o0/TTKBF
vbv0X1NlcEvtpqPl8TiboGKyfnYv/WpQvtq8B99zG8DC3DWphSmfmhwfHtz5S3bI
TSd48u2XvPacYF4M7/4wQRH2DtzcpT3roz3PRQH40U1rRBt782xLlPGbfMXl7Lil
yfNV0I8XZhZtLWlLzg7bi8Nb5xOqCuX6yD/2VbeyFsgdcIXJKaW2ukyd5U4Yq9o5
ZW8rtyaign9FokRdK/+uQMvPgXIE0ziIt6bkD0WYapj57DIhPBaTD/6HOxS39x/T
h2XnloElIXXgxDAft6AGK0vhFShcoRJydpf3cWDNalRtqRYdEeeexi3QxHy/21gf
pY1VayTE5ZJwKy347Ha2gA8pgkwDtgNHYV92FcnBbECY2Nf1/B7QqzedD+cbJYY4
ForVoms+cprjE9guNQCapeTkyefXd5DXpGLhtL+6ooCc7ei1mU41ApYtQwf/MyYd
THCkVtuRjWHCKurIOfPC2sxivq4mWdF97DTyLudaaJmAiscgjJGBfRpwRPJcoSU4
VfrHIrzVQJ9S/8gWIJQWL3JVjPIp4dfxCPApqAfHDk7xXpEGnY+jz5RPb8/XVQjU
hCAaNIKdulRuS3pdbKGmfeF5zhj9a2ize4bIPhdnBeaWdXJ3k5li211xaqw3APvd
mpsjVKDlLhzPVXgIa65VilV1F+DDYY5syIrGtfbW/B2JbM5iybetvTFZtzhYajlT
ooMDvLH+9XIaR/oXac6Q8ivFM02ysbefw5tjYtw1lt91WYD/GJmg4ERqIgSfMIQ+
4v+FscqNiRQcpqob7VErf9jOZD4EDDnAsYpoBInxPOA5dxcqEUzyoBCgh6j54vYn
TgrhoKh99K4oR5T3EMXJ8oB5I7BSNUaghibQLnUYts5V8VYeT33bFWrwmyxdRNLe
JlKcu51q9ojRm3eVFg9U6W6Y7WrWSsjWi+GmsL8j+t+OOj1Yv1XwVrBsMMcy2q/J
yhjd8QiT2hslvOqg55SWaQfNPE8n9cUkt5oLSGgS3uHTrn59OcVI7uFYg/K+h+nC
9wkehGlUBqrXViJ4hrYCeiHC4jTeAxEMsB6Dho58xdzHUO95HX/9WsdSZ5kPHZXw
6urnJX+aJ0e/Q96jRgJWOtMd/t8QOuAOpLCEpAYWq9eNp15hYFwmPVyORPClZMCR
iw1/Y1uAFGpM4npmmfx76EGlyBOgp+8aSd/G8BTWMlDJTtfR1F+ZDHiA08FK0rDT
nheZ4IrOWmVTsCkIyHpSwT4k8m7ZFUnygPO0aoZWmvEPzmW4SGSC/FBnGjOk9Ooz
N9CiOLch+O4W/V8rf52caealZxpgRNxjsB6jLRYBtbQ45G2YCJa//o6ASHcxuYlD
e3ir8uqKUvW3DFEZOpS3Cw+1pl+OQIl4seLXcrqaP/Oo5b0MA/bEXhnesxUXX1Qq
LUqdLZF2ZRpi+wmb7xqvMSvl35qoIdoUsXwF2uoekUI+84Z5+BhjJWp6xwU9Lqlk
07dwLIwU/iluOvVCWakxXH09i36hBwQa0qlj76AsAD2PPi0kZqo/Nm3bCFnSEJUs
MGWZ/HS4e5xmhwqyiLpTSe9PkC5ToX02P+jbGTT4HVyJwx9EdbZFGnrhHRPzk2ri
4LoP6SmOSqzpGNPDMncVZpvvFEVX4HxiuTXeVo142s1yYwtewDeNqgc7gD/gsajE
wunWM/K7i7oHKN6TMuxM4ig4dFb3HpXCbKLffHhLITIxJHJsOZp9zDm4C/0bdAJx
UtrOeameSPGl4lcpQU3mKqYmAwGbxGDvsbgaUYPjlIbmq2OHBBbPqXy23GhxQkLm
i2LPC69w69tVKmlKRW41GlfUEBOyT9+KJM4ZM8DyKX6nK03G709mzYaLNIVvwfXl
jea0IJfESEBS9QZ8KRmJ6JBCP4b1baZNw1tIFXtm4QPLPrtBoz5MLd/ZBAE67fSu
gbyK2z9mIZLROUFguo/IXsRtRJ5+hn/bT1PHmnGXhUxWzST2nV1sZEI5AKk58/aR
PR8YfwYY/T7WvRvhEwBVS5xNwScBWMivqtaO3eF5nrNwU91OsK9GtVqYJoIPctRa
FsfsWWBAslN3WdAUG/pkpHiWdfb1DSrvvza40L2J9gnu97kmZpvcqO/rXfB8c9b+
HZcCicjjbsrIRwBi6jL9+3N5p+E5IWjtszr6XMA9Ex2JsXFgRtYHy53IVRhCJckS
zoaEL4KQNWUBr3d5/4cLXfcJvuN1Hs4o63E++1FdYpM5StQttfG6uUC5u+ECoI2W
iwmc/wnFsXXHQEMXNRa4p/7UBKUzQdlPvadcVNQqnuBKZpTg+v7qxgwuk+0VVg1B
4k8qCLwkl1hG/gQZHix5wxUxU9mlBrp+3Y+ctGqlsbmDDRjTvcfsreKG/0Vo45/w
Olf1/blp4MU4AkgNCDcKbQqnZmDGPYYjU86tDW2yqrzPqU3Z9AoStMyRhbiIt+1e
+tDa1iNZ5DG1Ga2e/5zOwuXRJapOB9Yg3REoGQ1xiG9Hk2H6RNoHRrG5HkhwE7hz
yw9s/q4LU767gUZBqF6jNsTaJTTzvnebMroyTFfKxziH78fDmBwYoqk15WHI7CG5
/GlXInxw+Jc0g2ZOOfQQZ6UrZ3pIgcEmyFcbueJaRv3oVfTs9KgS393BMQvtkoYh
IFtGiZYbpfyxnby9+oO4KFnkBMKD2gFBZphEjt+o4bLn4oEetH+OQ+WoTUuhkjmV
ZQr9/Pvq+kxqGLV9XC11o5ITkmeqmBV/JqgwShvaaXWMMQQTvHzKquRH3mU0fJC5
oar/E/A0qZ3hl0OE28fBYaZvvZjdyKub4gQFKhhEkkgUPN79MkS2u+1raCqo+Urs
FCs8uR59BlhsBI8edCOKHlGDR/rF6f8RrjqAiJQtavNp+vZJq0LYaOAe1mFGGSTY
Aim1DkWENIaJVRd+vLx+9HyhMhLcKHKJpHKsoykfv+7zUaWdQ4dAQizZTRSzb99v
D9hxrYcY9rSDSXz7WN0WQfBMb6EFgou2+5Jlrla+j6067fC/F7sndY/aSyvZdUlH
JYiZrfnhvM0Hyd6l6zrUiBGSxr2gebjh0FyecrJJ90B4RWktAtsWAnlZmt7QbSZ1
tA720FPcWJwDSv5Ae25yjjpiNGr3Lunul3EggkxN7bwqobhLUmxkgsWe8TJsxmNv
R9P6HEzDS/7UCxMItqygidyTBVOI8IMYt9Vm59IWidjECzItEVlAhd1/q3CBW7jR
id1MTTXzH7z6PzG1zlZIJEKVfz+t+hzpbcdwXocae7tq/8sTHmSvY0FVi3bjGVb/
kRunlJs2VdyAWuJdZ5ycGPZJYBfLSEdVunCvu6RhrJyVpjzMJi+cRM8yiGAw231O
UBmq3dG2/uj5NxBni1rcL/7KNAiWBBq3/t0QLkFIng/4ayZPRe3PwwdBy54db/++
UFgFjNLQsdM/wUEvevoVGrrf/eiAKJcobt4VGutXq1GFak7dVKTZIFl1bcDqWTK8
qKrnItAgIL4yii0Bt2P5nvUhK4JbCvYk3tWwEXMPL037vv0JNtVWZ0NtHgWhWNoX
ov3rCUPJE4UBbiU3CemXcKO05GIAQZMob1BJw82njdKiA5j65a1iLNInAF5AJa98
65kjeDdjKRl2unP4XEbdqamuFHw1wZ64Q5akhaG2tU9vGuoUXW0BwHjvbpmZ8xxR
S5ivlTdPcymv8Do3gchg2NQP9eFcCA3aSg18GxXRUFXG9z7SCqrWJg9diIdo4IKe
XrzJjfN8BH3qecvoiiU52rAc98Gm//rL0NbNzzbPhpG8zx5VH9uTa64Ua5MMvgEg
18A+DhcayZPzPr3MgtqRtWdsJWo0ufw1oGfMa/UqhkulOyTdfiwFhcc+Dw6sF0qQ
q981LZhukueKdQRcvnk9+YvTmB/bX61Y5yBnPTcWGcu0zo+DbxQbe+WYkJbBjP8u
AY2NfJw10w01uFyS+xA90Z0AqVzLMIx2OFTV2wBwqF8T6tVg0NaPJm9f6PmU8exS
VonYXLJsMIs+ZWOV5VlFzQi1g+SpCtKarOrOvlasZvXlEJzS2fTRMatlgM8cpzoJ
7ZzodoJYBhGSZFfHqODf/sJPKm1UlhBYhKoUsxM1kGUQwzUHGv49Owpswy4QuS9J
KzuQwaybK+RpWK5F7Kcchp0uSxbbm6VitmtGhVb7ppNl2PVIcowpEWnJgFElWCHE
wvB4FufjkYkL4U9Cfnn8eoEbL+qIeOgWckP72CVZVV7w/q/40gL1V+i4i2b4rN4u
o+5v9XSfIJ48WQYSg7x/vTmlw6nfUDKuTUwdzaaW4w/ICwTIMzCaljLIwLe0cuCa
DwQzbK3lxCMywz2MwIIAFA+kkSU3f58RI946oeNOfNesNoB9e+TQKYFaHFEMugQH
4BRvmbdpCuQe9DQsHeFQwsINxjP2JCE3QNwtmrpfXTeo66/VjON9710Gf8p4RW/K
BXxV3J4ofLXIWtd6IuRxMkoBmXyvazriTAH2m/eer0FojfGjgpyALf1zwg7BBeVm
1mscJ0bzGSj7zNyR39EuslSzy1Ba7uwIGwf0YzB4jnCZzD9uIztFevpCwLtB6jM7
E1AZApFHYLnKAw3+ixdjLvKv1ayKJsd5Qsxi+9UeXRMzwnHp34V2Y01NHpeyIJK1
n655MbNG68pkSCtShdnsLyurFQk9sgODEVh9URidWbMXCYhAVkpqh8Xn2OqFqK2+
YB89IVhucaRPYTlgVkHEVZSzTotlT2qFusyq32jgpRkaHkXzZseFf3V/nPFWzAxM
MwzB2GxLKm1wJUe0cru0NWwZzc0zMGItayMMte6MsfeN5NZ5LUlMwheoThgxz6cZ
NTKkq1VSx/zU4ApcDC4ZAQKQOkKIg8IEC3jybxYV1PMBgK3RmATc7/+OVH6zCSsp
jzbFt/Bl4gujOoY3f0zb22MWF81feFYt8N7lfiWlYJb+e7rdUGBzRJFPvkGxrAb7
VUmawX1IfFDNp4hapwl0XsJzAF6rmZAJT774aXmvnaoHBp8xZ53flpMPmkQWIi37
DVJKmdWX9tlTSd15LpKb4/Lhkay7TtkMjfCEv2EroU2s/42kn4bZ60VmKVt2+jvu
aErGx1w9tJjc+ZR5lDKYn4ui/+iKLe1/nVpqyW9vSb+WrQ5k/KhSmdmoxlZfgB/z
ER1zXjoxRf3DOBkPcLaStQUw/+9ybFEoy55MBk+OV/9tKvad3OiA0XsBvehiyZDu
wKQRTZSBWZeQsdxYP7lTrivtbUCUSS/Sr5+tK5rEJGQwdWrPAaFA3anAqjzEmncp
NCgvgDV8JeEkXCM0MXHn8jAA/1PrDnkwYdh7ALH281OB5ot+AnIJ3lkKEGw+vLj5
h7fGNzxBwwxWPhb0RRtDy9Np8OmK2Oq2IzSul9X7iM/Obu+YDbs5aGAei6xPZUnK
QZ6Imj6leaTSIrw6Tu+bWweCuXmx7F9y99SLjtiGy9MOkskwB9b3VBOgMGtAB8sq
m87GzOXwzajQf9GUcgnmAgFBzbpsn6ZR+sQFfpBUW8Vnyapm/b2u6ONRr3KRaDEI
A33TvDWcM45aIXRywBjDxsqG3TE3QhbazPlq+hDrPBy11S0ryrh8qKcs64JzuZe+
0Nucy5Zdt3WdX6bLUShw2SIo6Wi9cNclhIa9EE7Y1xH8qBJ28ck0f53a2TJrJ8rP
EMU7ZSeB5r5RH2jTyGBY07mXiPFOwr1bhIvVwMzpF66Rds7uEZOyc0Ka9YpGgqSh
eJktTWlZV7H0+rbUgxOP2h5sGqV+H2Ju8lpvSPiurbutTd/S1yrx3hsgOT//xAim
iKt/fXoVno9cV8JMmScGfChe8b7+8Rt3i2ttfU4H8v41Ovl6wMHRyh4MHdBoKTCM
IucKLPjmC+eo3AAnJJcascrYbxEJJx5G8Axmnq1cmDY91eeVeegnGUZl2JYTzOgi
RiwtPPk90ukHf8ikhXVpv8azvgNHJAEvzBvZy6pU06mQrdiUUGs2eZIuz9dcvNVv
5ydHJqbSh/f/8rzklMLNte++EXdvUXtPAJhHCGZh9YnudwSG+F2F6DwGBBQyWBbX
YPv+lSoJqzbypskQZm+n/YGQWRednmBPL0nf+c+yMSQPmNsaG4AbtwBCDjFL3+xR
Skkr9eLheCxVPnWiBIiXSkiQYRmwGZhBTO4H1ErUjiyNQynksR0uJa7iIyTQ+269
i5qL4OZMdH3VV8KRrzcTZcKqoueSZ+CZdCErp6R3MaYfsgr9djuVqW3K/YMb7HLs
hP0GC7soVQc0U2ZnFGI2UVqUFrDY3Af4OcjaYxjtClggnLKnL6HoGrdAIZuv0AKZ
RMX8NkhwcmOH14PtDjyF/NnNxAuPkXL/tI+HXHuw5COy92/sd9MEDzKPcAXCcK0e
0zQW/KA5kVlNvIAd/ohnM86McT7gG0uzd7WBkeak+o+Kv8z6XS+27tgi649y4suu
ZCbspSNBeIjIy6TZkzgm5r8XO6lyXtdJiAx6H6YEgIIPzk5mliw1nojtL/Hx5Ono
uj4VlylZsMI7uvbX6fRkw9Xp66PEQM90GaJiN6olqiNaN2ljkiJGENZi8nEAidFl
OPtivk1Mh9aCmvPKppmO3sau0Zzp9pQ+UfQ7fB84kEQ7ZKOpbzrf1U7ilEXpGmRk
4bD6SR1jDeB8qnCFm0XV+f9GkXFfoNUG3RPkMt4g4FcoPO1CqBRzPCXYD8Y2v+Pd
wvHVqlMkQqGHSbEtErW3+C4W4kyPctBwt7QgpwbGHEP6rqW/zFCuzaPOPnbYK1B/
VVSdqx+VFYpNnsux1Trh6MG0eHxaA08yHNoPJPsjx3UQVWMRMFrNcY4FQyM5Otf/
zh1Wzsu71kiMhQbPyiJt+OEkdjYEm+OD4AchKV2n9+qvmGQsCYyiGvYR+zXMfb0K
bDZpwnHroQbxClAOZG23vTx/bwZea7hZtr8YLH7nQz13nGhvno/a/4EdP93Qw0l8
Vn0Md9u51tECo19vgnPOG4vj2hlI2M+U5HP0qM9x9fpvkpK2RDEgszc4PjyTS/QP
QPCSgZ2G9tnJryxiFXN4dSgUz6R0MYcrjFMvMv9rHJ537FvjVPLHVg2SHkxAqOa+
6nmWLsYwllOUIdUoclfFXnXQYVyF1LOLG2GtssPL+jwNcSOn1XfMgEV8dS9WvGb3
svZikiekslWexE8i7vvyfzND67ZOyL8ExRamVIbnztafgZyA9wKZIGowRSt3/tIZ
rZ78tfy5gnXWq7xByQenbMn4xUEvfiLGLg5REvVoNYVx5SO1wgOuEZ91LGKj2f6I
BApVzgVYLFNpZLUo4U9pLvqMr6SVi97TZbEQB4o1PrVfxAjZ1lBbuxUy+WYFscjL
MqxKtHzQs2tzB2q6EM+0pMFeJGFiHApGlAs0Qf3hWqgfwIgAtUyqGFMG7hJPcKPA
prQnEw91OKXMgfPMunPxAvZ9YtjhBbhH5Dxw1lp0f62IUq3wrJLhu6Zf4fei6RPK
1CHfAXv40e3uE9I9bs+VOwdpigH2p7RLT0A1QEvfslt+3/2unOwSKDGCGZDSbXdl
6rmD4SR97qOJknSyViI1t3sxoDfDWOnInmA0o8aopRzgkSzAZSU3FiyFHfi4bCqD
S50hgb1NZWIO6RkjBb3e6vTfhXqy/oaBlkY6bWYrjOneESrJhj63zjAur9Wzdh02
pzOpDBXDE037ZnLMXcieqpa/jm1pBLbdUHu5W1uSOb0i1YYMj4dHWbNep3uEIvlS
k1llZqYdxpArJy2D6BZ7MsMp4yzRBSpvrMR2YvPhYuEj9h8yJb3kRm9EDoAqaFsm
WUnm8f9sG8VOimXbuGsnmQurR0OLF14yS+mwjiieRmotfnyiMkbBN1JnsY+FsR8F
KEJ8KRhsNqkrjrcRw/IxFHkUue5py7bkg4fh9/gflhukKN5lSi+FptijfjLtho6K
Lb8Y2RA8lsLbE5l5Jissx/4XGJ/ekOakt1sB3j/Hl23BudMhq2OtdKBp6dje4aTL
L01F0KlF5CIVwRHGbvCYb81ma5bNpom0ueAZg8ayvgx0rBGzIAFYFOUyhY6E2Jqt
eVYMglvbSjiFmAPUJbWpV1AU0w1wuCAsu2hw18hm6rREMCtJmwcczqpd5ipoe+cI
gbn01uTXvdtLPYh6tA6nJu3+D/5OF12NsKMFGRt7mgxXnz9l7StiA80j3Z8o9kqW
EGJOcpX4iKW9f0e/eF1LY+JSePtk6dnwzRfF/mlRVRtsRL2dMcOyULYP2ZjjFa6Z
d6Uy9OaFG9FrmzRxxfZR8m8uLHv91i6pds9o+ZJLS0u3fUBj7YI5IYLSGvyo/eeK
NoQoG/14+QmzunbHZEuX04N2yGiPbZcm9Z1Kr9/R6eiv1L5JwxriH42td9G9AJQp
7Z7OIwKFlz4M+IhQiqrC6rBgRuTjxWwrF5lfOAVOS2pVSioR07okkcXXlyR0x9YS
0mu89j6bdOFnOphjRvIYI9I9J020RurBUFRGH8ccRATIR8m4ldy0cPDHhT0j1wIX
sZYNUGREMSLFtxesSUN/vhVE238Ow/eyDKXTvGW7sOgKVLDf4fKp4DzgA64xD6Vm
ZWhYNK4Ntgavu66AeVp64Or+lwFf5GnGpgLC2bNcNhBApFXRBPZwLBfVeCyGPSEp
CgIMtT3em/3+cnuTeBKBxKXFnZD46xfK0BdsmpFdwkiQfACXXdpKBfL5FnkTg0co
bpUVtdqqurQajz/JuIK/UTQX6uDgAmLoRZJ0HUbtkb640qiApZ9sB5KENq0lhlrY
UxpC4VrChCZpXr7BW3Equ+cjvRyHd/Dn5t6KJG5DuPKUzqGlMvD+F0QOFF0X9w+K
zsO+Lj/X2SBcrIMRh+S6AFnK+9x3s7azPfaFKLA5bj3077mlkgg3mXXPvucpvYQ/
WcjNX6D7juER/RS1O5XxjFMNK9aF6D43nJL9yGSxZlEQjuppDyp3HCzBLT1PezVM
eJFbBEmAu/E78c8qqNvzu2Pe3sjBNb+rJMuBhKUz8XK3IuPOTYr7thBHWWfguF0P
mIhUAlcfuhXJ9sZGaGyIbhFgs39wlASH3tMEuovCErKSHEkMk/dI/aEfCSx5RaZr
dktauFWVZd25EHA/eZUZfFfQxabLnpZ9s2ZY2K4wu2/Acvy7pYgzhgiBNIYjNLHy
4QV29cYzblGTApSoFOS6uvrjag8IwRlvkgj6uayZtJSTxQN7ZQn37QlMCHhMvH2U
5HVO80siud6fqtq+GSvDn1mLWOPGFqhChsES8AGXdP/I5uvjderOQYuSMp9ytqLD
7Q8te6Jrf8lNLtSGGQ7HP/jabs8YDq0JL0/9pJfdLeg1vT5MSPyDVTXte6b7c2Et
aMQJc0/Sx4MnBIujYo7fkjttKi/yz7UPhqcuTJe91Sjcptv8ev2YpI8+M93dL4Lj
GIpStT5xWXJu/q5NfMkxZ0szouXAnTzAimvZhTW2h+PObOr4oHC9/rehwa4NrMkk
6WaQwbtf0ddiVf2hHvpNkMBsqKKymgx3NF4v9TrBPZDdiB56Na7XNB+3RZxvzE4V
WWP5+JaR5cptKaU+oMOz0AHzdl6OCe1cCkRm/4+kaAXgX5BehSO+nndZJcCHOYRj
Zq2f+J4f5y1rIbeztsVLq85BhA28ImP2BYL9vm3Ok9Ck/PzRYYbnopEbjIgRKvvi
lRj5LtPqGu6d5NnIg1fKydYG8qPWporLtqlW+Lwys78=
`protect END_PROTECTED
