`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OHzOdEYlDWclP5gDYANdL01v2uqPiekiuPbKEddig+S/JQCUsuXOFi8+RImh0k7N
DzivZymQBwtZDEqeVmWRVF1o6Fan4RFla8+1PWoENXLcOAFPtoaXJjfAIZnInihN
wI5cl2LPv1LIOWQ6aDZFw6K1k/+tFp/IP3rvK8CItnHG0oy7IdFOHzhR+nAEqt0k
e88sa3US+SokHx+Mls9dECT5lLxnFExhdGOdJzHtKZeCbB7WLsJ/KEm6sZJqimTU
UJ83TUaabINxTUWP2sIqlAOQrD/vL9ACKWW9y7sm+NuMTG9/4TjW6+dQYOiTXho7
jn0SBZpkwobpNGqAIW7lIcfR/uQdJbkx+KC2nqEc1NGevPLrvc5+gAIK6L3ZjWYV
Lgk8VS73wWrRds9kKYTSiF7URu0uBLWSJvX9HbdcWs01VnFlVgIoamz2cwtLBH4L
b/hrpbxBDcNu5XcI6g64E+WufrwbWTrj2VsJ2BZyXfjPRGhLLCGixtzbGy5W8TZg
Dk8ERGHfwryD1PadYE8/v+EGdAwFBsjAfJuNPZKLyLVR5yiHLh9fG4dRyXnAJnjJ
YByDpDQwgDDRYy63xBJleAUEQdxC9OpNdpynd1ziAJeXQCspMjDhxyS1hqYwsojA
rU20ZUKdrMcTNj/6iDG3pb7dt+SV+gl5MA+ntdw3HpBRWvmMs7wPI+edstEBaz1B
axVXXrD9U1XgrReSqTARfVWrVGVMx9xJvtVG/VLqmDxrp2gyAsFhZs56Ss1n9rRZ
xERh1Z9vsPO4JDkwMjVwf9IivtoybQ8keh1h2P5d8SM4VtDhIVaeKy9Ulxy69CEA
p+aMKY3sa0+KsOtrvQVJoQ==
`protect END_PROTECTED
