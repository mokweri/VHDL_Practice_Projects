`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnfZBfHpShpHOVJNP463jGRMPK9rNZ9BbH0bL1CJWTCNX9zaWqV+C+zRtEldidV5
aYuqYsOKgyVGIyGdUiu//EI62DMFaWmECiPVT/zA4BlbeT6JWdks76ihyQCD7uVV
1Z1fghIN2DbMMiw7ldtZv8B+iLDutRpXDCauWEaGxvlNu1Dr290RYsSjhBi8zjMr
djBLuC2ZDRa/L53JyKkNhpEErg3mfpcD7LiUdBZtM+mVCGahcF9m5LpdzNNId69F
oLE519S9IIbtcSfKFDBbh708w7PSDKQfWgk4NMU70D0mwqL7m/hu77l2OQT1cnR/
aefvzNULJORcS08B664b8rHy4qw4VLeLEQNrx2jLvObnzvSBXfJNUx/MPHEu4SFm
ACj/1k+i9PNhSdk/ZKDIP8AxaKCBXyplis21AMOJalZhILsEzq4zr1Yyg8gSVXBd
5a5k32MHqQEgtE3gRiuwPsZv3WKFeYVMRvjupXTp7o0p/uk/q4g+/ocU3a8iivK6
5rvXfKNRwLTzZPsV2y3XQxKaPQiUOSEXaK8LKkFIM+S7lq/nD33EXRiiMfy3op8S
NKkVEe5BHVGhl7mekEDb+BDN1eRn2HYW/6OgPT/Hu1vrDthD+lqD7GZ3LsnTcVhh
jzw8tH4wmnoKtj5qaO0Fyd7YAJt+R/fvJlwbOT/ngicvWdr4uDh6josihbXyv6+K
ybkjz+ZI/IF/o+u1grc7iBstvDxoirdg7VjBlsvw4d/xhBB0Cr3KsIW5NXM2oQmj
FQVbBiljm3kSQJrpa94vC8YSByX/HqfsjHlzI/X+hqu5WvuCOufqYRZziUxJaGAV
SUWWFbHV/nSeHq2/JNUPk09NQ3v/I8Jank3HArrHBCjWllKHwkksrQlEchAeIoLB
VUPt7B4fBspwGUWM3MqpfaLau1H2/q6Lh4faBAYGANp3764yksqq0vJFZHEjwIP1
ZkohC61a+lxZn/DoWxFuFNnxkre4l0Ay0zTDcHZ3nQ1mQ3jq3UBOonQ30ookQ8Ou
taGpVbbjatnBrwF2cJUyoudFkiqtucAPUc6nKVfv9erZyk8ETH7rcUi3rQnCe9A2
oDkFXHidRj9xJ3KuUqvXYgl66TErmc+mzWGxjy9HwelAwMPM2VVOLBhqWU+oU0l2
L+A8CABAf2TOWBcHowVNTKlKDy4iXGgvuYZA5H0DfC0ALsh3Nt9yjQKRNm9w2b1O
BcDWxWYpjSsmHjPRObknM6yyXa7R3CcRVFTjRurA/5fhWDL8aC8sLj84V/3/IAu6
RwIn6Z0Gr2s99Jqkspxc1Da0VaQvcWz87oKB4zXJEzYHL95/Q4upPbnmEmmt9ufv
afQcFCfbDDdXp5th/NeNKwjFeBzDR/yWkaoHQ6EZk2C8iK3/1wSnHuUVaIf5bjgH
COI2z5BZo1MIyAyWIqocMyolu9Kz1uUeat8pM4h5ovg3d5GjKnYDJYJfrOt/FXrS
RQEtNKsE4ValkjAg/R6vkr4XDAXs6H8xt33+DB7/8efMP44yBKADMGDkv8KJpwC/
OXPmtSqEbKBwsN0RmhVOcJZg8t51OiIDIqhHcKucR4HZR8oQyGSFMsdvkymm01Vq
VFG5CyG5QMpnear0ChdEqGiXwkiY02RCKSsN+G3TB6+SZeipcfrnio8pToEL0Rgi
AxeK+Ob7lXXQEufgdJym7H0BBLlTYWA/+tJlvhCaPfmfwZLcdR0R1e0aOrh7hqvu
lVQ5xGNJc6+kVA6xdb8/SL3Bit/sA6xntNzAF1CYfnFv1geKqIwHX7G0Zu17b1Ak
Pf6TTvueAzuuWhqUrzdrYJmbq3wJEQTpmv0Qm9bXEBBflZPo15fRDnBGmDvWfsc6
CbF59N2yoaOyb3hkEDey+foSN/Vk306yZq5Aprr+knX7dB5m/0ihQNo2Ekte41g+
u1wWd46BeCwk7z6ePsYLh1OPR71vbYpTdXYsyNpQRrfYPPRcg//ZaxMCGE1PZYMq
rxdKHRJi01DnWsSomvLkiWK4NyaxrVf6+VblGt41YLmwltAy9+jSJPrtRxp7Qpm7
idrSwX6NJYzPy+v2Yp6jCMZTTmQWRDH//LZRfE5aQYVOT5D++rbHW+uDsEC6+eVm
Rb1+1R2zW8rfO7cV63xkMcXK0GwpKJQMSeYOUINJX1RKGK5MGFWDsqKy8+5WyTeZ
2vg548e6SmTaa+cGJUWFvrq20L62Abq9j31n3j2s9sDLNf3MQNSWMhMZpuL1lyPT
w/wvI1tboyuudyN7VwOnFj6Y+yOkEDaMs/qya9TzvA8FaVZeZMQic4gPQgB/bBki
V4Cb797hA7d45e2NmizpxZJEbl+YNVgOIRdX1BP3xzd5/xeAcu2HdbyToKpDmyW2
RENnfBQqa4h7Zm5NX1+sTFo3HGKgfQdKHd3H/SuVxYTAoPWfifuB2aUcFG5h/eHP
9xgT1WlTXzbjZNrc7P5quhxbE9VRI3KskLk2ef9EVhNnLaVFeMxYEhDyLI7t0N29
IFpbceqE9FpIdrE/VnjnpWFsfw4445WOGC45PprUI5AzVLKmhb2DxxHNBEe9b9cY
VE5d8mfcqW1rBtrhLvuOdA==
`protect END_PROTECTED
