`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRceL+brQPk/s2GYF6VPeIL297pG79KVKAL2B4j3uM7W/JLKaqiEUZUa2LeyUBoC
2hWRdEqnWHehLi1/25H9B6zp07ft9URZmgOE3YS38w0nrxqv7K53ih4ZdN9GdWOt
760wf1TqCal81qsh9gjx6SrHiHbJ7XRvKBj530d5II4dGYQ3J3j3Qcie+yby72iH
YjIo5is2rI88QDxT72zETYkFYrgy2GFuabpnQfE7DD4xX+mBMwwWehVdLilsPXP9
JJvSHgaZVmI4HMh0JkuThe7ROx9V7yvxuEWcVwDkrChxaY/3J25QC//7q//hC30Y
YF5Rs0U8JlduzA2TLGJeD3JyJg/4oQ5LOTc5hh2o+2/18/7oZG0XuBZBWbKPpmiK
ksRzjHCqPn6k+6kYhAIwcotx7INZjnqnGs2Hv4zFf5f4+xG2UKvdZ/fjGQUbSCWM
DnIqX5N9pRYwO0OOOwwUnwyIgZPL5zrzzT8p/FUWznF1BxMl8Uqj3rGivt5QxRjo
c8Wggkb7PWtDSmoOn8zhqEiNlseI2HvmU6QeYbnb1FWTiusK3hQMoVV1BX2HlDHr
HtQSMDhGewbkErRZ5n1Rk4NZzo2oDb0TxLb8lizUwNCj9JYmxXQB7eDexn81lHMM
RjnHiqcKRbylCvIpcLWQlPh19t4Jg8K2Uo2hcVxd1QyI/JLWIC0hl3p7dCEuGLto
L9Jsk4O9vDtZccQC4k7YxeVTsbn1akBDPHQsDlpS334SMbvAzNA2NXPnrycAS43b
qQuAdO7UqanC2Yz+S7dITeJ8oeXQ+Rfi5P4d8cmPR8AR7aFXeMh36poU7CPQFAF7
3og0fz8a//HVu/lVjdjt2QbXB/9KAQSBFBVCWZPhzY34ACkQO2CwxDjWxRM9nbal
7BTW7V/QfHpDzd1zyYyDjEMGIbHuOHy7simoxuDDOfNk0lz8o6tq0aBUGCrLyWTu
3MplyPFxrT/1ro0mes6iWYsxeyeAJo6QVemOxghd+L7YeZocBjCOIcye8vfCgbrE
DwZXp0z5w/BmtynxbMRMjmx57d3PdJsj59ut/5EL/dsFYGCpSDqbTyRMuxfi/B5h
XMzyqYRY3nJV2sXTHKJUWjFJrw6vKwIsLonmDAnDzvv6VDrdooXRvEekd1J5zRoV
fwOpBdqvntmNPNEGi89piiCVN9KGHHof9HfNAAve+CfHHqq7Ub8clntojOUEaRq8
go6x5Cdx2mlRJHSWmWTpZ991RqHPVmGNFQFidPC17cDfOd7nHTd0KwfKE53LztHP
jY6ene5h2o+WnmO+tpIdXtbjJaocogRPe1qDyaj0N33on2izm88Kto2MTvwgEQbG
6tqbcagWlw3BZDCFWghG+8I7NH97NzLcczAMS2chYGvBnK798yXc82d5kbkYudyC
acMUjXyHNYWBWXoctFGCBbqg/+bApgC8GY/bieawhTGp/9x5RzIJr8eKz+YNXxFR
dbn2xN1MDO/FUBTWyUsOpZCZUDbcWWZrbrYD/su5sDmMlM+K8pruLv/7Fu5gqwos
DFvcKFgLxhcLvPIZmRR4qqx6z4C/dvEh8cimopCnp7yLtD7br3E96GKpwThbQ3pV
VFRBufe9I7rR8z690umUPZWRFRlYIcuxiYn9hRBGsv5nyrLCFMcXx/3fdLihT1+P
nKVY+mP/1G1DWnLxOOD4hiBo4S+c+mJRi8Sx92XiRk/Rz4RQZsUVxv9p1Xw5jWGn
jxODtobpOHaSmapqQUt8uLVIjhVBlTXgqDLjC7kykLtETyZg0VmiH0o4XyBjGr5b
y2SNkt4tTEriXZ45wuuJa9ummM6Ppa3cPO/gM6x1dPIBBMJJGo9IChdVWb1jtjzA
aIgv0nOVguOiEGuY4cMg0/VKeK/e/l2dVBsjYFfUU12Ry9N5BvhFDFOv9jDUw4Qd
6ny77o/2FH7iuSR4WNE1+0fAi9D+uyAkWLpzP5TycSfs/4X9BOnHgFwsDXgNKUKD
8tpQhCYLVpUWhvakS66S7McDd3kr2ow+wkIchjkZLAH3/Ca25czZoaVGm1n90ros
7Lq6esOH1kLGi9TUS86vMfyDqB0cCFFA01WIYZchwh7qTGeR2zXtKXUlQCoPK7zO
tIyWQK6cL+KGbi8G29ibCyruzAbYZHvn3/h73FTU4rWKbI4UmIggbwBCZf2PN+Lg
/GGBi1DhS+lISrdeq1/pFGIXPfM726mIlRqoFBByd/muE7Ab6XkAmB0xIaSYimDX
9/lVIg6OVL3Jz3lfpEvc1jlxSIt9gE/gXvEVfm9b9QfkJR7/STzTTJBhfH/4AJ1U
ZMws/0igF4eDnJfgjhFUZ4I3ROCdm/bTL65A+k63X9qL8yPKczuwWtWNldeTsDQW
7FRoCgHE8DcbppNtnF/o2KiVqHmP6mp2LvHrUEIADDNiWt9OOaJLCeIryHk3f3i+
VOVxYx503FDa5gfUquOrkYXfbhTjgxPeC2nhuNJ+AyU+YpKPbF7RicGdioX6+C7k
yozwHqLcH5UJAldJTx1hquh/xitvl86SRcNDmELVv+ekPaZx+9M856uKx7j3Z9Oh
wIja0Whgw790OINDz66AojM28o0BanO6Kmt+boiDMHqJgfcuXd8pUZKU231hJLmJ
v0On0vnbPkCnCydG8P7lfH5qQQv2WCSIRkJpKXiM01LRGzCg8Q3g0tyUAcDR7WoL
VD1xkbCmoe+jGaQFO7ToukKDnGEhqC7zKXPpNGzXKQaiTW3ci1Olr3Z4dq1i8fP5
OD0kBfokcWNlqVeEZMhESZy2OQWHfdc8MUE/Mz35SxKIn0sJdBHMf35XRIEtDILo
iF2YagpvXVwCe2OYITHuQYAGCetIzza2+XZ6tOfmiWPy19PSXE/Xgebk/FltnnQd
9RIU/WHRuLNmAg4q95JFtyqf5CVXYNAXq5jFPGevdB4xjQhc1ZC5T/RvTHKEjNcU
DPivOTEVPwsko/oyJOTbSuqVbondndChczCQibKawMw8453NMAgLsVLfLBmtZLda
VUlNj71t+zrgXMmDxh0YydeIPxaetcArr3PVNDknnmUGpx5XmxtM7tpQvhihdndx
sb+4HgsSR+jVHy53RjpB7dYlOgRc0+rk8NtH2gS/Th22hccbXVwQcujfpP1S9feH
CdlcIMNPE68jsdfc34CxLGFjj18j/suETulzjmOOaj+/V/scATVVQQw8h+Tgsg6W
CJL7oCmVTKKPispqP7cKL7cRhj44vkZ0raAJYQ0suxSPnY8mQ97ux7rxoQtiaMBa
af9THYgP0yoCE1ou6S+59hh4PN90ey0qHuxmODaooQL/MOHcvjVOEuGWzXvSQ1vv
a4mszRNESB+lvOvX3CQi+jXe51GctVvldT77LJk2HR6FxARTsT6ok9o5wCJmLJBD
ClYzGM6R15HlwIj5FsNniQRqmSq8oFwSL61rzX2078GjilaLLX9NUKYWcH/NnDNq
T5qOA/BCTcJR+Z6tE8b1MOlorvkJCp2PckVvd+9O7JUypWCNZKH+j8z6+F4m7Vnj
VlpLsbB/ytP3IOj+h4Zb5CSMEbcWuFlEVsWsnFUUCVFgpxaP1Ru2ZtSKEzjskiTD
B/XhJDwcBW5kp2ISNJOHN4oP0ZkMauliv+GoUgpBrUaau67SWkl05stXMPbSmIwB
/9XpYXRS/QfyAVKztxKF0lP5WiuMMDyPHcVpMomwvNSjAVomtr/e07oPYmzcIhv4
rnhcjDVz2rayqjQHlJGNUm+TWopuBsK7lcQsLUdDq6awm8Vfu9tZWJe3PrWbFnqr
eaA4o9uTxgfEyIYIClrHcBCsfmTAUaaCp/A8/SCG7CeTqDtoAgiaNU3Xi5WMj3z4
lnJaPKITjsXE76FNdqWP2jVq3v6f+avWZADyFCgeebs7s4iQTzdFSclBXq/D9TGw
CV1z/amnnLkbu5JBLX0Kan76nrlzvFHS6jgGAqgdLZsSgrxLYmvRq6whbR4vkYtv
UTyQ07OHcTywt6yJ8ZR6Zrt5bmY9MXuzcqHZk8S6AIDfMY8J6eFSfOJu3l0JLpVi
5INqxHTGdKAv8tvM6YN4ts6+ufsDvC2NKekdCEXJE+flwT2l7Vkw8gPBi2jjRKb0
1eJx+oBpmPW97pAR+2kO719s7rAUFhgfszuwBZaHaOrATelqbfJ16kyCyBlLpxbZ
O/3ZHzCx39JAuR54WT84MHGv0vvTpwrbw9nyQ6b1jxdQaROa4lWbi+tfRO3uVVbC
lYMMDMpXW4wr1DbrADG4wYYUXoHJTzVsCVM1W+tmI3oRtetsiXdEWoIh643Qil3m
ZtCq9BGVA69xM/cO2yTe2bDUy456xhA76JcTeywxThZz1HiNzLq34nJQTrxhEe4W
nHnUKHQlECpOX/ZiLUzY/Uu5cfjunDm+wyK2wmMtQqmNsVKDZATy14EWDbzFDmgn
teGvkXbWpVp6giF1Bj/O/HgUXVZxP6KAPwMD0i0+ShLo/Y8DfZrTdUUm9PB/BzjT
`protect END_PROTECTED
