`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LTlbrP4kAtxJJUGXvaDMOXtBLlBRZCh1NrcPvrmuqz1cZ1/BKmiNMUQb+pWYsOkc
DJWrw60KWtRntA39zlI6YJmKEDtPqmvwUOrnG9YKC9p3KkIbqUhi14+IlyegHKVC
gdpZ6ucnKjqSussPqI30NIhwsnY57iZ2fbv+jSjcJV7K1mRQhug5J+dybNQEIQJZ
yflcexDWIdxsMvY1joDDIQfd2ZOU+Agb0u6+FgY6ElaPHI/BH7vf9iB3vnfJlwU/
2E4v+dRnxYsdpV9rGEuXS8Lk+L8KkZtZ6gD9HEEuj5F+Nr+p+SjUxd2j4isWyyDf
R4uBxfJIQjrh3/qcynLewOPvZRy7xK5yyMyKhO/4VqYA21eVSyxDcFtU6EJSFAym
LA2ZjKj5LIm6VGYMFbGrTaD53mj+CObhu7wRy9HQro/DIphYxax831QYL2RNpnyC
Q0A2lBzSd1tJC2XAUVzDg+IZUuZ/7wK5uup9zbwmriJPrHZqkJjn1sdtVXNBCews
b1HYTQUEaofgY8oj50VsRrGRKF3dZjyKxqODP6a2YsP1tcKn1B/3SVeh7AqFJXox
8uoxg2GBYxPhe/u+cOj2QR7txlQ6jsBAAKl2Z9c041r35GaOOHC7yYXM7cD6L0Hq
`protect END_PROTECTED
