`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZ3QU3Ee8Ykie8LHlOuT4TtCLgR77tf42C0G0D2FLFSuXpoY9vAjRoGmWJPK3ALS
mPxhJj2iNhIAdL11L6sfo98ej8ccJKohsYnSCMnHQfOf4T9v/19yExaBcgHVUYgQ
4Pf5ObFvUr+tikCiBLRAq7ibKExPQyBu93zD7OUPZaYZeieVsexc31+8LnBCrdOS
2V8y2Yv5YuJxDDOOiKvG2PBoMeMkNYuravfv5Qio8an1XoZgxANcfkv7W5USUiGh
ON9uS13iLzoLOs6zKPVcsLuMzI9QVeQBni7Tf2ddQj2J7oMH/ipgOZJlnhXuOLEG
Z0ZB3Tx69jxIn1VX+NB1cJLWKYTHMwr7vvnvTEjz2h+GozM3z9u2p/uRz0/KmXN9
f8XM1RekueWfiDsvb3owFCzC2N2Hp4DQvKTYDWdGpqGCqjN04a4ea9ac65vi43Uy
QCnzXqHnDi3Czc6IkvuSbUL6Qbr9lyLaL6smjQuo/9c1iQqwbTM1/0qobDPRDxn0
QJAbCEDUAz+4CeZMyqHVeHc4mIyCqpPsyYfVGSry9g2NFn2xfRpJ0+dm5GMeiZk6
Ski+KWJKT7fRHzT7Bs3TYB8b3z165iwsomAjZR54TBr33a5TfUxkIr7CsDkAl1RP
cZ4NVbmGKHuRThmsauNVhvCgh0EXHLMyCsLIqHG4ROGmrHqfR1HF+5uZVSihXrTu
j6Kej5J2IIOCPU14r1AitfgN5nG66fK+loFj9C4sKcYHzCb0KAlJwDI+VtGrcXnE
LRLRo7MhNyRvglSTJabEaZaXtytTxe5jMJAdHD4IzljGGWA/2NIf8VQcR8n2Fsok
wcZQJpijx5aZGLRycY+2hbykM1unRY4i8tXIk1a89vbXr+IV6Rz3E/3lbTEuhT56
XznnBl/AXh8gaw0wIVsSrakP9ZFZdTLVoeY+GRIWOXU7Gub5ZWhDJ+Zkvc9ynR/a
W+23tgsnHDSiK+OEOIiFF5ISO/GcU2viJ686pXkqJSTbhIXyWvMW4+G/hqzXJewB
2otd1ZNcEG1fFx3YVIkf+ahSBGG2a6DOYWNYJSOPGaRTboxK5FMlYZc23gD8dGvX
nH73vHO9PAPnVJqjR8Lx0BOZPcn5oIkx1D7nlFxN6anEl28vk26IFQL1CRLlJUk1
h09qWpF3LtTrQBCk1sT1dIzErzQu4Ln5fcXuQeMDyP6QNfSZsK+VCkBvzA8Kx2AR
16YZOFpAhtSAGpgNR4yj0JpW9hVSjUdAWAQ9fimbuqcciNW8HTFjz0uhCdBHuaMn
gRLptgaAAOOd9u9tm6yr2l7Wsiroy8+y2penyrXTMdrt+Vv4n0iIC5m3E6qnd688
hcSD8hrJ1FxhBHP9mhtbU6Tibnf6MjJva1pS/4WLBKLwIJtYMZbpIL4uuzztcQZF
EFY2+bJc9d/rWp6ATN3KiQHP8roWWvUOWgYDca8P1Xdb12X3iFp0nmUeYkXT+QnH
wjz2wyHhXxRgDIWpo07SXeIOnJ0n0Oo/BDVMFe6WPUIED5dN0FvQhxoy+gncCNCk
xBgRteCEDG1K8PwsoIR7JhozlyU8l8k2X8GncbFsR5LOhzw7C2tuuQGp7ajhjP0o
+diszqIxEFDXo2Fe8GyysPJ/bJpyB9jCtHG9s0HurZdJ45Mez0V/Z9XhBVabsq/U
lo99KKVEMOhxWf8fXhha+R4yMMJKR6W+kWSoFwd3pjy864YMi9eMgAUTLd/DCXyk
Bjan6Ugn5DbQq/ZwA7C7QPfzbWlzUQw0OkNUUkscLf6g4m/3jVLCEwZbSkYC8HPp
XjSh3Lme1YAkjiRpdgFB/QabH3xdx7RA1wjkVaAdPTjO21m4AAV1g4VtHG7/TQX1
LIWNCnxI59rMONJKdu0g1NkfDl3Ot+/2euzMJXX2CxuRWW0fcCdbIunAZffKgdEn
FR7KrY31XVXIHJSD3qgX4j2v7bv8Eo6RsSHZfZteCxxVllmHJjzHFXIK9y/SVvNp
OG/m2OGi2GMM4brFBSYQOXJIqNsCFY+HKFnvZLcJmDJPEh1f1e9jhGJN7oYCXrDo
tZQhkFDJkWphRHB49nHq0RhLpbCXf5YsmRAp8m/P/CYFe7DJLAu38miqYaKE/k6d
HenYoQxhSHxr7Oa71ZXjAd8xX7ISCWdtj9e9COyRfSXr/c8bMx5GcrREDWSF1OQ0
cbRV8Upk1DWaCAR+otxuqRZVV73EkrCr2/d2WqCt5gKXqYCRFhfvMCZmcdQ8eOzA
jQKv5Fh0Jp7yHecpz/zSE4MSqZ3nt+GfsjAOIzNZlwl0g9aubmQY9Q5oHm3RQOiq
ZYBOkdnLdMEO8DMAA6uV1IvADdboTbu0tJelivFJk+726D7v3q/lBhlEZTyfsmyG
ZSVlrUg1qRHjXyEoxmYXPBqsldK4oMzyXIdfADnEtu++IW0Yn4MGwSTvnhcwHRx9
03zAVoe0+mmr61ofjtBUEcGoKh+fENoZJTj5uXZPQ5EF/J8D3xEQFReOzTDHJqO1
N2zWUAKlTBn04um3+1m6R5yEr00A/eEiWzAU9iJSbG2JxWXPE3k4s3tw1DnZMAme
0z0vXeLfuu0c21ixZovoAKzp6LFd6lrzx3LmQQosw//mkuKDggbt2QVEkTTVC9qd
mo8526VDxH7W3oLFFEEAHFBCQzvaTXUDs3IcxPB5hYhf9/wGSas7bDDaPYaoNYQh
tggDqZOYm0XEjK9xGR32NlaMYwTpBEbm6wtQ3Hjg+kDWRexRTg/85EyWlqgMsPCo
7bNfYbO3jpYBjpsgLDxw4VsC79Il9lYLAygojqLXEZ4H0azRlq7mfY8JrGJCIg/+
IlysrPu2e/UESprvWEMzCKgoRds6BTJaZGrvWuqZsA+LEaX4hPX8aiZXvoufT01T
PShnml7Qbq8xCkB+o+lwsqbyCwbvqgz7ud5GJctIyDZ0BeLyvDNm+K0vmHnckVx9
SySjHvgTdGfXbvL5kCqelzdZ66br8H8ElPGPFGAKCUyVudAa/3AH/9GhXccnO4ek
BWN4zIhFHk9rHilkcdUKkab6nGLtmxkLief6PdwrzQmoGotMv5gP778CavnaAAw/
g9lFO9hrLS438aZ2uUtMT8NRn2/yiaVkEmYUgKIlK86gDHz1AbWjaBo5VmOCETI3
uyzwMGh/yt7ACIHwBVFORnQlqw54gO10RHKMZpUCKCBGbqBaeY43Zs+9HzYtRcjE
ThicACZYvuSxOvj7Rmtx2Sj+s43p5nAgvRgtmUGabKeC79E3Xdd8gSUkjqHI4U3K
j5W7Ke8wSD4HjGO0wHZX36I+LV83Hl6xpd5ZhZdOt79lTQCGn/We0lQ9kfB/Nbyu
FCpVOcPaGek5FS2w5aC9zNICUf2PsJBt9omx+La32G/NGGzfuRZ8AeeCTzHKVxp6
2m2PYOUDBfbzUjm1XazPxP50g7qOVZfjhF1dBiEf9YrxXTbzqZhUSF+Sz/o1IdGq
2cdDxk4EEuEb2bSKb4Qle8sI68i84g86Qj3GAUd+4sojE3ja/5oQ+rO+sATbmVn5
MpZVwXRSTkBkv4LNrwqKu6I2JIFEpMjeT1B7VLpwPcLIZa3K9ZJUpvNDV2eUljTC
pCjmTPQPlvhvBXWxkSPmAPm225P+WFkQOeGon2+Ma/GPphtUHb+w6l8kV0KPZhiG
ACRFzFxPzXRiTDg2w0pduSvVyk/ddqUhhpHk5wNdYZHQqKGmQRg3ZvaKiRKXMEQ3
MCaS4mUl27ox5pTx96VNqtGSiT9Q557r8tqESfFcl6KhGEkU4sV4UcAxBqMz2Jj5
5094P2Zr21fef7ihO+iC+Wfe2tv1GUmuIfPKnhEADc082/ljuVEzq7ZIdQVH2oUi
eROew/vmEKU8egzmwZQd+GE9Ss/kXj8gVlpMQ3jYBnel6Y08EVICQIu+k0/J1qG2
pd0qBeZt7LtJmRlujDEpiG9tQG8vX3yq/gV+RoqbGzMm955nivvXHoXo6SAtEkoA
1zG3w6WvR9PNsZVv8+dnhiLDstr5SGsLfLO7PmuXcaGVpj4c3lRSqc0fS3DxLGHC
a9cI0WQ0fYQnJRKZLHBBcdJTBUPcDamXCMNkrt2Pd9mGoGZ8wnIZ5fOfnofB95ay
Jm97U+agmCJ7os8MoC5bd9nplWLQCsduxK0Fk5wdEdiY6PdOXcn55gSitIwpz5dI
7Jag23jsT1xHWR7YUI+hzQKeRikRcGJ3+vAYDM9WqJSuc5DPhL5cm2YU4uyiaupG
Osq+PbuGXGTgOLD9+hTmQIBh5/pmOI8fJnJoI4bPYHJy0E9e2PKRGANeIddA9DFy
kgs1Al9uZa7ngFHH5dgn2kpK8r6FPyBAM8sq4QvkHwhiOiSJ0hivXfgvjQ2sN2DJ
36L1j4jHvdYJfbxcA+DsgqybKin7d6DgWIfi7SsOTAEQ0UR3LQgkvlxNeZCKMPFd
d83tDj4F0LjJxX7VaK4zUi9q+x4uX1jpHWSFaUT3vRoFPXp181wuO8hSfq5ZC3ob
2vdFlA4BHaUcnUseZ4bBSOAKUE3IPsJ528Vl76oFERhNo5ObPei7Aik1X2AmZxP/
OroY1LfxiPhFsaZKVrm9eUZCS/KzlZ/d7FFuU8PdWrWpl+2D+0MPku9/9WUbsRYX
M5xIthRjTC02VVrnf2mL3NF1RBvhBnP5oX6oLoU6WH4If9tf28PL3ECG/Alnk1oy
0FGLSt+HddATYKV6v49p5nID0tenjHP/RWYgqQQUl2AyrqwUGNMVzE3sZwWObdHi
1Za+R+hlmQmDTieYI1TyS7j0Ve+dW0NWOgnl5oNYZu4r+RLWqWUkULl2dHTn2Rv3
QAn4GyN8b9ckDabZADIscZKrFRXJBfZaF8SR4OShoCECYDlIUvRFhkTaT/jHQtVA
YNWTtpQmlnnbugJr+G+1xAxPwNTEuNus6d6yy0zJgPHOIAsfbVQW3nVQW27QyGLT
EjBJtqYUwnIBaJ8WeFh5T1jtkhKel8Svxnd0pJ8IHmNe/MySiU7t5pUlThMYrJMX
qqYsHVfliRYcU0vL6gdlFvfrCAKJ39sVc1f/d3Rhu/MGB6EofWt3evL2ZArrOdCc
MIIBDbn7cmppwfgpvB1x61jR8Dy2F0lmG9bWBVHQ8UAs31Bm79n4Sp9oqu1sg1f6
OESOH2Iu4Lr6qQeHV5Gy+yC6iioOh3AD26FYh3MlsNaNKX1+XDdXVVm4/JxExTP7
tQrZGQDgbquZuA+lYcN6V8rXxDHZ9hvEnxxav3K4+rCrbIo1kuZ/frCFno7JKEnk
5ZHO2fOPd+rh80ilyNDvnoNUZem+zyGUZmNzVQLdg8m5ev3OooZwjHPgIBlMna+n
j/iS/TBAcKSzbNFBvl50jP3oKa9PRyfyXwsh0JxThmX3xXjpKZMbDqbevFzYZqzD
/tC+5ECVtVxhPy1xvDmTAmLN5Ab/fCdMEiTeKkDll5DlyQBYF32VFR2eDkNcaSQM
aq8SY0ANGY6Tp1JDD2PmtZL6P7NnfSUJxvSmRguFafsAygAN+FfIMMZ+AMfTATSv
o7ZVLkcqaI1BEDUS6iZe3LdA0HvQyrAnf24Rzd0gECg7a4mecaoWsmNPI40+gm8V
v9jDDHvseC2IQgH852S/HD8ooxDrZZmg3E6vkww27NSUAPNquwE+dLpx9HXdB/gh
+HL+CeHLrQRnr8j8T2WGt8viERjeFV5fHoB2X34uPjt/gJGf4thx9sPgoJ8QbTkz
lbXzExKsXz72/zjXAUHZNROrr9oxOoEfMB57C+oo/wRTzoecrQ26lbOHJ7K+TR5j
1yoe7T3DAoKtrOIh1EVy6+ZwQImZHQRts8ZeZspo3srkiS2NKkmHPCLT7WdFgPNT
CpwaeOhXfsxA/9kV7msSQLOTmGYXWAVS6Ep9A/pMnF4fAMOLR8v/aSZpY8K5FlAz
4czRRzhEcUYwnsFpgnHJcTj3tJNq0tXhpNcm8RQkYMFKJMMeBRfw/a7F3mLYCVP7
0Hd8VtIvcvVr5d+zTuEGQKVpEG94cQFB3xczb0115OrnSE3cOVfxmOV6byvj+Qv4
flJJqcJer7pG6HDo9DT05Zlf1n0ccVs/WO0somwwqPFHUKalUgHEMVvpCXeAVucU
u5/CJS1K8UhDNMdRozqP/S6PhRyrgzarM7uBTOTcfD+WhlEbiMokuiyABUhCyPE9
7wgiTWi3HGeNoAFVvm/5SnMqeL5GWfrlNO1/L2xN2eIIGu4UeztEVkaW2GrRAhvf
8Ngr5vIpCFwffIyw41b9iIGZb4HtK3qwourYPhEBeQfhOuJnSmCB9SgU46Rof6BC
rPEeQkdD/w9JaZS10hZZUI8wRvEqMafZp35ifci8BQ1JNXr+xvp8sowe2DoEU6IS
p84ueLLLRM0QwOyB3ulm1HG0SWCQAIizvw85JHmUjm2qXItzJGNED/4G9A2LT/o5
puBkpE4tK77P27QYRM/8olrFVO3iLdeZ/tckHtUH81FmMceYK8Pc7aPyNKaehneM
BG7iaRRk4/wCyipVgj4Om4u8KLOPr9/m5H78JdiWeiK9Sl8XRutofXOPjZFwuXC2
lkElFCbQQdzASkPsnS/Uy98c7E8TLp5F9PClKQUaq58S/xB7i9QB/S7YD4/mcpTq
ZkNZ0Oo+j4YI90s/n9hqI4udUWZinMG6tnaChx//emJq9s4xHe7blf8rFmFlLLaT
JAMoCRC7wI9jQF5cWgcY5RDrFLo852tOSwBxJeti5WNdVTdhfWd/FAQq9VFm0fFl
ZiRPXeimvn6KhFx63nLUqWXzt42ettXIF4M6ZKapnkSRhERh9SGSeWSM58E6EshZ
kAZmJEXKM18elQV2H4RossSvdK6wCA22PsNAInbaRaEiSem5liEpnCCwvxQZ/Idt
Vde/kXGzbfyyscfRmZBn0pX+9VJiqkOQDARRt4Ki70gp+rP4NHqLTy1EW4fpjmGz
YMS+g9WoctS33xSy8fNMJWiKCfx1GdzjV98DYppmLbo06bf4rpCkhTrxGwcWnFcC
qU8IObOkHSE8ECeBQLUvE4IStUTdsuxAhC3VDYyfjIFDlYZEoL+qfHDp3zj0wb56
ADD3MbBQ18dlMTM9B85H55Lf0Uprj5QerqS6fPDSD4Xv09VKfqHVbHYsRuwHJ6Kr
0748SA607cCtir0piw1okfDmf/+rLYR5QAQK5pvVceKh+FFRkNWAXY3oy8ZsV49y
/QxkMpGLAx78gNmeHDqbgbMDtvmhzOZVFpnqeBoAJCMqL/zC2scHHHYKvKlY7jbw
Wl8CJpn1lDUQNwtLpKwVnmsBUen7RkCVEBbcqd5is1GhitzmBFmRzESapR14NUEg
RXy4ZF2LBE8alBMTKNGdeejq0GXPfcpNRaruexPSulJxaooOaiXtXq1MaAEI4HCS
upKB8m12UrKTvAPjpd3vr9JwiBJkBX8/4lUncYBSWgc/g3vIyp6Kpw/05Nd4+zXB
QrEjUHVTJfWLGdFK/ZXBjVBxaLdz59cZe0fxsFm5/cKESD6ONWs1hnwjZuLC960q
gJQMUm4vUC5YxxOAZ2Wv3f01/uHemQR5uEuc+aRyL8MdCL/pt1SQvfBw9xYUz3qZ
2FqTIlJUZnqeD2XU7SbS0lj0GIvIsdnGQuVmp9yCCJ7AZsxPlet1xkZXJUb4RJXQ
gxYasQXCbn0MOzA3ctLbnbfiMz2ONzUB7gFEiTw/BPrtw6zk7czW68OaLwfWe9sK
khn5LENoADFybeTrin9fImRDC4m93lDGHs4Jx2NJPwPX0voODSVngPQgoiszHDFX
N80+8NBBRhlHZvjmiet68WrAo/yst8XpKqur9ooXND+z9OC+UCcvrXjbpCU0M9xO
DR/IuXk/LBftGCVbtm0AN2oyYsSTsKFMOnQO8LJd+MF0jT/ax08kF+55QWV/ATPB
1vkOd9rQMDezwc1htvu3HXol6RGaa4647G7L2RJW6SVmVcxDX7MTMdN3P17CqOA7
L88yp3WsgY9l59tN2okj5rr46FAP8QmcGJWJGCjDttyLHrGC2gUn7HYG5foOCIFJ
ox2fra2Mlnt/vOab3i4ENSHqgcwnOxPtsdaTS4lnJyYYdXRszuL3hQu+ugvjd6Ru
XIahlpB9PHk7lkBHIqwuqgELA81BVFWHlMP6svJFPo6ST7Cl3rGvrUUV56ipuRfC
HERoWaWSsFA6L73yD+GzmLWPV2eaMtykf2YXLq42QnsaispgT+djhKruGZHjnivN
DRtI6R8uaG9BgyIKIHuvxtaUiUU5tDAGoe+FHo3bxEkEhVrShRMvuS4nypzaV4zJ
DU/mZIfNpVQZpFZo4iYhUozwuzK3H2jfiUIEv7Yoc5YlkQEyxiGqBGhYUeuXc8So
2vsqgCvXHe/QPR3XuwmLYRXrPkqgPRSVbqThbqSgEc6EZT8iCk0VPYUeii5mR6P+
CQNHPrVs/6qWpnSapi+4WcFPiKFmsEqmEVQ++YaE6fvtx71Pz6HMSgxTX6bJSaJf
/te9E4VD1b3gLK9sgsoqEBay0gCnq/R5/5NKOroZWSKNA7lq1DnDRYdrr2OYSu6C
8LeduOfEpKOmWlVo7/iwgJXpnfp6104t+xJz1SroaQA3gmH55H+l5zb50UIe/N1g
ShgOrM5rJYD4gu9aDqNLI8y6iqaG8Fto/hB1rcPov/gTtDMpfSwodKKO8+kRAx7h
517soTb5f+qUw9tl9Kfks2IRa1GEN0UIs2kdtpNW0KRCON1jzx45fupu9GDdIXnc
LFf0VVSBV/Epr1hKe9kR7Bn+JWFFuLlumQ7xynjKxmdD6wdqz691nLCTIP5jr6WL
2B3AguRZZpzf3wtE7AoaV6WmyctrHvVUvPw1rbGhqT4V1VKIMxlTeQpeHVZSqiyj
AzzFJmqLsyeo1OUc2UnA8buZUCmLbGHlkxhsD3DEbGs7guDpmBb1bvR8dzDJOXhS
t/XoDgLds3D23rjBVyaytZmdDtTorhV965VZbbwIqf/U3/Lvyeql3n5iTma/1nTc
3UE13qOgqBiSX4qUAKrxoDxAjdCDxLkJglu60R87i1MLHCBhRzRHfgwNMuWCmQ0G
+6YbvYsE9jhNeSNychU1vdu8IposV5Haf/2BdpDbb08e6+izuPF5RRIz/DxeMibA
Gt/25p/pmTEMejIxnzM75Y/l4EeueLoDsFqdM6g+AfK0c9oCfh4jmxVqmV9dFlNb
jYg3Jyz6YuLmjR/zQXQ5Uo5JXRRgsJXcv1iUDaKhI1fkuqxsnHB9leRN6rQ6VAIr
Xmj1lezO0xUM1IAKCl5tNqH9yw/Vh3daUzzDX8RUzKjkIsAGNeMzWz2vpX0Phego
P0QOEnK+0w393SIA5kNEUv2fOwXRG6L9ftKtaEZzPKsAYBsHLiLLAcAcV/DnG7T8
fQWRqR1CASwWmzdWPd/yJXvZXORGYVfEjSZRet5OFmlO/m8WIC4Tw68u1pF0m9+O
RNsbzt5bwrnb9WlLxMiiettbsrg0LSrjHHlWLdDmo37SHxmW5WfBHzgcXLai/7Uz
JOSpzA/FyfMQs1Y9/EGo8zYMQwiL5yKX0RsOiJR6kWRUZ+7gIhpUNIV3/tUF7+Di
bsKOD2oOFCx9ECCHP72HGc9wrjuIfwReXB15BGzN+Sa9mVM6ZKrS+22C+w0T/+z5
KikjpUAzChdVkC2PfAcHGCxreiPTFonlMd0X/vo2Soly9iPp2G7SlMySRysu/HS1
FK5lO+cnzPF0W4OeLWrZR+oPn1LT74/ngwVCp8EYHwS8MuHmBs+zA3oUeV/t2c0X
mwrbYXoMYfEcYYv28VAD51fCbL5aVDOxUO1o0kUafmhkV0fwsEuuTYlAiSLcyE0d
7x1UAjKzgKnyMQaxPjJIy+42yR6r380ISanK7R78Y+LzfzIByG1/Xv1rzxwYZEMS
4fJBcHxzWfMxG1dOQovV1WNvcidbqmk9XGJN9B+Y/C7kjKr7T9rwb7JoGnFcTQyY
OygtGtMXD4eeqLDwi/MGFnJiL+N5J2FUUcn2VGwh0aOyEhggUwxml+5L8o5KpDlI
yzm3sm+L7g89AToVK92gTi3RTqP2ygS8FOtrYl+N5CJ2D4T7H4s1i30lYimDvFJL
I6pG+7RnYdTFOJUj/Ah9SIpxXYB8GVt+ouLLZ49VVPn/a1tmUE254pNqTGkOOZNk
YFHlW+h4xhYFPCUOB73ZVvb3lFZwprkksYS5Inh02ILH0V97EnlpHTKTDp0XMKOI
SqfyZ29j59Fw+UGpnq39ekSFQ0qX2k9VFHw5PPOn0x34e5dvd3nkgxephOXiWBBp
Hmd1ztTiTmlgWdNYv9q/PVbY7a839KhRWDq52V9/jCk=
`protect END_PROTECTED
