`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX3B8WceTWyN21wjS8O5d0WsIbmuNhTH1mIvNqWg+wTk2vVctoNwGJrQ8gnH8AZI
VUZ3uDttH4VzeEj9YZsUTKlL0S67S7rk5KQjuILZ730ZqebFX4o41l4f/Ibl1IXk
9Que/Sl3c4wlY/wkTDUOmArU8hOmMyMIx2JN2NcEeb8PrNPIX7XNebmeCEzHQEC7
x+/7v5FOvy2Wag3lCkEZVkhXR5ortWhINTrmfXvP4gQf9+zJbBX2cKfZayP3FMHH
O+QHvtgWClavBua8TaTTsg6BD+XpIMmkqGNL7hNsf/PHmh6XlGTPYjk+JqIpTeYh
4RBuwBme2BK08KOKFurlqiCPMUAdQEzV5H8s3eh599toU1Wuq3ouvhZM5wlZkBuI
/hcCUpq83R2mzH4I5ofEz6ldxpVfwdo2vbyX6FVCNgbRuUKAfjeyGmoa1Lka6pmM
SeJFPfumlpH/GaM7/p5EMukhemphuFCYkJ7C58QphH3Q1xFRSyRbnaSu51WNHTdT
6mn1ruUbKq2nRKiJgRHguRwrvs2d7KPn2PBfae/r6+fInfvso7yWtuNEUxwvGVKa
WeOlTOwLUsABZVqxvGEhe/JfbfNYqfLXyYGa0NTvv8QhIbnAPz+eAGAilee7uYl8
e8oNktqRTubFAdFj1y2b0zbNjQd3kL5NbHJ5pi+raKxxnc97IZNhiixybZtgecwa
XYDn1c0wR0f/d+TNawUtpAvbv8Ng4CEfj4Piib8PW3LGsf9jNDTodMJIiwFR+dCK
vicHfDgiBvHSK+neAJR7O2PRu/g851EM6iQFLv1f6/mYazSSHuUKHE625ylYU9KP
FDsq3SGcqZPSBxI8ma/KA+SpSoKEdqOHiUtnwoBtFgee6kkVOa9le02Pmh3s45Dd
CHLThDAO5F+Mmpfyo38yZmFNHHmC+YT6QwfkAZGs5YnK8MbO47HBWo8yzMTQcyXj
sYEXuILXjizUZM0PtOlUpejHgwh/1A5tNh4KWLzSeFyPhAIqALOJKxqwzg6z0p3k
H3I+zXmpDexH+mAfeJLO+Q0UWUKA/uRgFfCZpYhhorhU3wlj2u0iGkod/jUmgWPg
o/LU2G/j7kEVBvsAUE2+JkM3ud/3417lQCcBy+6JqU6CQZSJhyEXyiSbA2udUvj7
GGjAzah3xF6M6Rcz1xHqDFfG4z2s/zJKkliwapCzKbLqdf5KUoSxZD9tS0arE/ak
UQramzwRlYD7He+fQdKGOwE4NLi4TdgV7vA1BrIrNf3A8P/591GqQGaPybjzwqpl
By1LT/TXFD+xLbD05Q0a6IFGqLoUL/iQK1wkEStYkJUCYYJSPQgNSJh0IB86JrYI
yRbTkFibobJ674m+Wqk2FJLqV0yhaxArysBfOhDUA0S+VxWWQ/SBPcmDp9mCYl0N
cf+MsxoP1wCZNTIPG+x/bEHsO+TM3NMbpNR0U5IY+MJWQKM3GOJcQ89vm4de7SAS
4fL5gKGihkGHPbSOv/axa2ERbylw7jcsikO+0OlSCuWbeBGxaVkBd01mAAU/FUKB
q1RIeekKA4yKcSJv0MAU03CHHdKQvcz2hJXyiv1jw/2RWqy36//ARICOHED2fJdE
4Wq7oMSm2RproJ7JsBOW4SePwZEE2Q8ivQdU9VfDXh7G6J9SPvZzUlDWr3xxaJJw
L7eWO8J6Vv/tx0V3SIqctYxHaDu8bKeBajGHp/OJDcQCGLO7rzDoHDJaHOEWc1JM
N/E4/cWomsmiKayG3Fn06GIBKZs4yFCJ8RgMdPdRWTnw6rSLOOrHKxvTvMnjuI8a
hj23hIupo+ponTGKFJJbDgr7uwU6r2ql61H1EAurX/YtHsfNcIb+olkOLetEPrXA
VCD6/kVhDEhgiR19nvPBsu4UmAQYtdBxGZ4GcWoecwGwNw4J42ymOzmJ5fof+5jk
7Kcu+Td376DQHDL8F8Bud4LoPIUR8dSDIho+fJs0EjIleADhkZdr3wCg5kSpnvOP
V0aQOLdBD3tR6LHs2TQSuuFybQSeLkZOlTsmYYo3EQBWDpTLEtvbhw3xOHz6QoVW
qFyNH4MQBETPJROT8t50aTLonpbZV+mKVaGAtwpsBRFgXk2iOLddgbFw62lz4wd3
nreyWyE6s/tk5z9J4HKIhyUZ3dOEcfTOZ1+XS+Fre9XUyMzThmkxTVM+03I0Uk+O
NTF+HTWyMTT26EhqEYAhCOTSJalgOuLI85ltJKtiHgP6oD7UB1ZUSXLdreAmXBrG
4lP71CIGzopy2r05gNsP8sAqgmzlY8saef+5dRdKgMv+MjcGNULxVd35DuWAlF2g
Wcsx2V74RjNdhMWF63E/Dw/LEaAfu3wekIF4jx+WBZsJc2InHT7i6DBA9PPzhowy
vKItIC2m3hala8BnZUlk1BnKN7tUpy5+6FnzbyhSNScBUaUPvcB4z8BqZLfhF2+E
6MNOGXHmfIgjCsuRRvNvRQ/8bemBTySddrLXwxdhEh2xfznG2r/mOMHlrwrUCxNw
YNQwMYKiPYVtr90nTH+XnQj3dEYq8HYIcSgug4a4EBtff3QbrQKjMgVM+beslGPy
dATni78EDHlmOergmkkkgW2mPRoBfg6a74onFOWsCB8lNQfk5PN56FX+vguFPd4P
DeIJdOKGAsNJLuTCpJ9b0lbTnkS7CCsr7aUl7HswnMAHKMsv9m5deoKBLcL9f8ed
x/c6evt/BYmWNpAkrELsyxsTsJyUem6PYPy5zLWYEDqBa3Ec8ULhcFYISSIJWWlU
vAGE+cuOZjThI5uZQ7l1JMBUooJWZt+affRTuNRti894EmcFSA8TlYvmacJr16fK
zzUdnrqd2Eq7xkhpu639U40IkHuQhqStYIgl0LdJ9BQxPytjedavWMhl2RS+kLYP
oHTue+ATlA6wx2sZcBkN1FAJF3Hu/bez9ynwKTyDJIHgifGCYdbid1nNLXfZQM6O
XySjfNdCBxHpDA4T2ODOdSdWavKm28Xo58DZ1SKlSqHSgiRpRbjuZZ6oTRaKcuTG
FwIIadlYM4TKXef8QIwJiZJjQm8YqRw6cAHmCEEXW6IqxzMqX5/VJt4Mjg4v7kUT
9uOtBUve+mSalBfX9ws3mUqyMW98B2S9CDYMqtJIGsu5cDht3j5NNi9j+e34unP/
NmFaodhOY7ao/rXadD27VCsr5ZRGLYhsdL3afRIL2IypYI9H6gju5saVGcFQEV/v
EnbFTKWqezlCIldl6ZamOv2IyweYL3VSDqm7Ng6FgochIGcMlNu79N5zlGMDgwhd
tSPWvtIz3egSSOle9S5guZ41xeEG9a2SwD7xtM2LicR9vD0wckG4ECGtAg+j6WH4
LSWsCv8rt5h7RCU2sGVQbnUyT6Bhw1CUvZcykfyq8lpl39dtkjqqbGQm5wFm5QAs
OhReyUOWF4OaORhThMUwtvBqY2f76cXJ1SJ7XdSGsHEeKHUu4t01qjoMeamlxXoA
vDwhSt77q0nfVzqm0gP/Fgmw9Mz4AObMXwqzwcO6XXOgCLZn5nHDl7obxpXuU2AC
sYBElwMKmv+T0HrFVJ4D0P6bLTDWJ2KDH9VF2Aefge2P1MFSI2ZzNwirfp67gsoD
QBwMZrRKUZspvFIPHxcFa+sgrKpjvXZzuTiCbFt4pv7N/DrNBBBYWaQqtmNYRpRt
TCOV6+3N1gQsmGio5fKKAkHsAKLKn8Ieall2+/qwkUywgVDu3zOWvKNg+D4TplZ1
qyy0sbNl/xQpDMJdq36C01bi522KIm/BmCxUGp5KIFMrz0rwvXLfWAym/bdQdZNq
s2pg9lmDQPhuJZlYOzB32uY609yHeeaUmgSTllmUoBrqM64S5eegT5dm+BMaTzXK
DFA7JMQYEs7v2dmT/7KluFyv0HyoJdD2X9vwJBA/Z0ZpV04OKp0orgui/lmpqCpb
1hLMYUgpgEd7mO+S4aBUZi4bRA0PeePLWGfDdbW/4beffpo+QXbMt9NSjJmbVDXW
2/fzVNlXrmRTZzp8Gs9GkQH2djSyqA4U4CIZR4uqaj8ncFd1UcXfeBjBu0H1XOwj
CJjSbRSueQ0RMhnFmlXospRVCQtacAnyV1lEhi/Yw7+xWuH+FEiJpFyRePoHuSt7
+6ekRwUWRIrZ/hCsQRCeZGuCXilAgYY5ZXGiXo5m8r0H1zxjN+m1UXfOajxRSaAx
y/iZT45bPjl9VVb7t+esjODTnGKJJKjoUaQ9KKaQgg0OY55TRH0HjUObm8OXYk1r
/pzR2Ji1ku6pOsQzsEgBTaHHmoZhVyNmaGVPUakHEickdPtl/pgEI/uVVIicQVBz
jEC51XqbjpmnbNV/m4Hb6Lf0rSk51UuYPZHcSPJqBExoCAz34WAZLWyDX6unptVk
ZOL2SM2dLGQY2WARzEck5xZPGh7EUhO9SdGdcaD+xz9L72kT3sSz+DCb8CU86p/X
B4XK+9UzUkyvdB3Y0ul6qexVh5w3A9wkSLkhfxtVZ+XozNmXkNELiMd5hMKF4wi9
dDSd6cAj+dHGcoNiE55/lcKePpddJ+xviIjRVTDmBUJ4h7rMTGsgZFWmAkD3TnWP
SOTYzcQ478w+HGfd9AL1L47RhTpw9qpM4dnLQBy+K2ygQtguohCnrCYlskdsonrj
zs2uDbCkAVYtnAKpWrwczvYmYRrMgq4SLWFHC4I5WIp8NM3MZEW0tXElOExkdiqd
qgLxXS+qPwX1J8j/4VWzpzROOtgBGaS/KfG/C+4FH//h0cExXKNdBge/hKPi2vs4
AqYnXRYNQtI9cQg9uqzR2yT+4VpfEcPmT8lMzUsHuAEckfBn5N8x4JqHSaNGiRxT
VGXX0blRElSw+9gadu/Y6/czk+VsCvjfRRmUtiAH63oIqSjuSMEg6TgHUf+AidEA
Vcg9N6adFTVGKKSIcpXGWjALqFKPN3SBK47S++zIxplLoe6mtLZndvzIGSwgKEhS
09sj+szOpekiDPhEpd88QPRS9arRhV3VkgHAPpT/n10WEC8S/FfjbCZMd0f627G7
0N7zHuata9KatCldERf3DgsVcfw2VAMVOYYwVuIq+luDoQZQlFiO43sjmbf2ZvCF
quIHG30ZKj/1rF4Eiwj0ubKhYBPNPRr/77bxx9wgvszCtEVz7gsF2ARobhmj5e3X
LLDSPmpv9qX1uaOyq3iKLxUvBnOimfu1bi2S8S0RPr9Y6YubSmH/QsddvmbA7Z1m
NYGsmRA+707AuWyAbs5tSff2mLXRkO9mNTUUvsYX3wSaiKoeiVqcG/c8OzRJycGq
g0cpHnu5qV6OyOHqmB3w2/0IciDglC621lAhIASWAVyQWAkJOgZPCRr5wOiQ89/m
AEOcgX69wBi3dOl1MxAVEtW1Z+q6n1+DKklZQn1BRpnWzSbBN7b1pAuJ4YxdTeEt
aBvxWq9BblnzZ7Oip4rqdOx2Rf3fmbJTSt2XLimnbqnpgEhyucgJxBJT+5N9lf5c
YG7BX69d/kELJJO6jDPknD2E1C4pBUyvDd9HLlEl8iSYDcAk3wXyNfse7+Uxi1Xf
Qrk3kzAty/CCXD7qLN5OcnO+1LQaPu8KzK+ZYx/n8ramSaap8GE7HUolpvi9/D5a
UPqPPWWhW9w6/gk0D5N7QMMIW19O30qgQQ17/qePu+GJE4SAqwJhrklZ6FR5t5pG
ecuwPcCn4PC2gRTrSu7oOxIZMqYBEDtP7QjuvRaOcYRWxXfy/4/+jBEkdEVAdjZJ
Ii5p1pcczcRcOeYBhaagqTY3UGrCcpA62TixzL+JmjWrgwXqgzKyS0O5UIarZW6U
Aaho/gSHNzuoJ+pJbincBVOauAIh2I6K3vJeEcy5J2IybGdLt5xwkYPeQYfPNZ+c
4oKYaoO/hTTnRiCdg7Pg7KAI9PZWCG31LfVDkzZiXD64rALLl5Rt6LwsrU0RI7/M
ObVXObuu47SbDFAvFsmdcj0VF5t5+X0wIEMVxYScZIzfdilWvSJoyYIDZkCBKQZ/
C9uAwKU9vwdsnAFuiYSyzo1ioKo58IzEyEwOAWaWKS73hIQS3GP/7CRVb1V3tno4
Ky/E/PcU7bg57K2J/djD8HZsFRH6kJjlHzMi/fjS/Y//ydyVLVTr5mksu6dPLgwi
bMJBP4avc613EVAXO0CqbrOeUcxEAHrfbjcq78BdJcRjbq0PdA/23fUroc9bZ3NA
9I+Em5d7OR0dFjMuzvDYVovpZzE6qUGmcvMRbWItXjWRpgKAyJg3USeenFiMWlvQ
MCVUHYg6kw1L7UbGDqK/Ig8TR0uxTr49rPh1/V0wjiwSXZdr/fKjnrFHXRxpn8MD
HsmVvhca+6OtE90y5V64YxM7QBIbQlMUaIQomToYmEpkK5exuKT25GSIq0dwspfB
cP0RRtWfAN5g9ljmN+DfGkwIA9Kv0w4+IXrPvICzdWFNAwdNAvC6EFYiURBV9JdE
kfLypve0AtrloRW2U3PaoFI/VCznxsKsDrn4u2i6HZcr3jlL146BZQ6w0IhL0Og6
TVpJitYJM5S60q22+o4jSWNzvzj9i5Uga6CdCf8JQEOPpARz1PYr0XTiyaYwADn6
YsuMLJYU2t1oK8+dGpEYRHDe7Sa5mbtH8xwruC3EKsOYfB00Sfw3MSH6SAyZjpjz
F1lPaZdCUwLcL4xz+kkZL/icv+UHDIWZyXeTXZ9OCiDljJ4F0B5t9JC75Vv6X+Mx
leh3oWzG1dN92brtUGY5VakGHfDwbxEjcv7kq/YXfGPhLFv15GuMB8Mcm8ElHVg1
DIQFGvWKsw3wPAoqS1Nd3UTtijAou7b7IzqpYwB0QIvGsSU8m1Q5yOaO/C0ZGVbm
FLi4UI+Z99+br7P/sOyOv/2kf4+mEIobs1qI1aM/9jfZSxJHuZwISmVPqKJsfEyi
+n1wjAzKs9NYdXfwY1aslCJS9loMfcA+nZfrIT8EIxZ3RfUJ8rgFJlplL0B3ez5F
CixUebu/XykCVqWHyZ9IM0ZnlgSqv8fR0fQ1gp386Vtl8yjT8FG2aRLsI+2mCBDl
XtD4KTO3nn5A1sXb4B/nBNvDXcLOxVrpJL1C+Cj8F0D3v+QzCySOlSTbRfhstsAO
axtvymuz9bIbDxMLoxGaP7cxbnIVs1enAs7SsMvAATyNQXv8QV4LNYzzr0BUb+P2
aaMi+qIFlQHjZi7mccgQ2SkRqjGTNkw/KWyMxy2RsmT+OwO6wV2RdlTyN77HbDGJ
ONtqEAnG/OqyX9QA5fC8ET62f9ZuhUG3UfrtHxEmNOaKi6+hms/DC+W4Y+VlVirf
RcrbSe9DyWoKy67PAsqIRBWSOTZ8bJvK4wPf72HXQQ+Wp9j76tMakOURvPbVp2DL
Vzh2HMr8i7USU+9A8ZOLpOvZ4FruAFK0Tzspjd5chkD4Jb6lH8+cx3HJ75iDkoMY
dGjKvUrGmKwxhKODCwCae67+UsXu1FozRm/f02Obtvqfv6T7x9H2+6U8AOCjccEd
+xPX2sjIi9MaIcIyTXLDVcQiAGgy4EaURgxJsLn1QFfKlu14CtT0Eta+fE6j0F99
dy+5NVLRj4aEuan0mxPNNaum/Qulm8QXODQSMtmp3febG20xyAY1yG9Ykkzc1M2K
iO6E8yd1XuS/NSL0loDq6MWJKquk04dh2JhdUNadHL5KXHmQVHghgZBNhj5gTlXx
QYBHspFRWBA9IoQlaieCdFeNDBENQ974O+1YIACoeLxNvEJvhwInw/LqQsTBi9wh
BUcov8CYyz3MkJdb3OkHoQbzIr7aPixbLS8A6LsAdY/FmLEiunm/AZNsmxas1YTq
wXM9fDhacYlfWORgPFanMrescykxHB4WnEjR/jQ/kqwB9jD0m7+jXpL2JYu925iv
cj9qLixuZ2flGV+eXHhT7t4P4Wupx1lUI5RnArOl/1KyBY1Oy7OH3lHYqkrqtgyi
q2hBGq8U6GCpspZ/qbujjZl1aNzlfxbWwbuaCPIOesoEAQeglH81s6oJRBHnpfHq
G7j0N1RfPdlm3h2F1SyPXK5bPc27yDBtv3AnCeHSJAHd/TItBXlAB0/HytLp3Lsm
x/EUfxwQZwDy8ZON1e4SV18gOUysnSUR4ft+GPOwj53yYfjpQROFTLqZGK6bBpkG
5R0jAc8TRvuJDuI2B6K6KxM6iBGMPO0E/BlSWDJBmRt2LerP6DKv4xw8VC3PQ9LS
+fdSUogQPdpLYZpCm5OmKpNZVWpJp+ksY35GlgBjT/jux8FLU1WVb6sF0IKGft6K
oMOazglFdmK2nvycPE0/iAwkha/p1xtD7MEKs4j0IYGrxq4xI1hZdj6V6Wyz7a7J
wg2pyfeJtnDxFM6UoEpnEXEDR82fO4Ili7CZM8kImQrp9uTvmR2WY+e/hQ86RpAz
DHY0smtAutqUW2FYPeMZ4rtPrSV/DwNo/cSIm6295d+dQlcjpNozDp0zdahHkLwp
6gxx3gV0Oip/EvJqV1aisGup5+VDgicoiAMrYOGqdx+5D5c7VFTK6lXnoXMSUI4u
irevOFZkdnrEg4gTzhmJg7NlWxRju4jL4GkKpG+LM16pgsxHnN5eUgE80OXC/sSY
LsK7jAeFLMOrRzgtNBJP11JQsINH1kNNydxM7RZwNPydkmegn9LDd1AlzX8DTCP5
18UgV0EU1mKjuIIbUSmLWjf30VCNFEljeaDA7gi/xroWnekzA6LDqe8lgceU4+H9
/F1mGRO5fk6mo7AE4uTElWVEPazkCr5tQ9X22ZZL3I6Fp++JUkilhFXan2ZRhn/N
BB1bpVDY8tzSBeVRPeoAF0l7UQCRp1moEDVAvveYAkQTLejJIiX7FV21ATqWLIv5
GnZE4W+IFkDmX/+n7xC5MKSCqW5p7u+daMLAajQTtsg96Wv7lCt/u9EiIyHVAUtS
muizsLKGmaym8QO4Bg/rjyAHwU6nJHxXPVRHlblEj/fF0Mw5wApO+7mQif27owZw
ng4QT+1k7hC9KA6nBUX8kUuFvtQSAbh5t79Jyc1DlbE/ZVRNGibI4RlnC5vGM7QI
BP0SSJhrEhfE+PMgBgoabIhm7GccEEfUXdZp6va3QoDkmKWZd3gu/+HCz2Q8A6ad
/BBaA0Wo0bHAAQKpzVF32SKRMiLqF/sjg/fKXNNniuGWaMy5+2LDsppAf4zl6mj9
OFuGX6aTu696gt8+2kXbumWFuUhP93QoHEI6nTajZ9YjBQOyUFNh5wnEoG8u7QoZ
wF5rVv5N7Cv2NiSY+l5VvHTFuBB1JLJb+Y1LyYR/qD7auR9Ja3TD/9uDQKf0w62/
BXIlMk+fjmVDWFu/1v7oOyQiYNGw9Xq8hSqTGAspfwAzCgaE07A8Hh11A5RIDmZs
9mZQAzPpw8Zq2A694BOklJWNLCUn1RYlE3cu6jerH2nS70dCT8pIJclOII9f1HMU
6GndrTz21EgnWlpowIbiaIbLjDTcQd6MZz39LG9i6lXDx+CSqHeMzjMvbvs4HjQy
zPoEGEEbFucZ2CAVInib93dzHsFxutppiEis4rvRiPvWqTMkasaGa+qO/GPa4bjp
m7rt1+CHnKwZi0R4+NiUfafjeBI08J+T9cSB1mpiShJSlzald1+oK58xd4/cuF1J
b+3IVRKd9/tEPVK47zBpQzJhsTWN7BQWZn/7sjhtgQI4NDwYZoXcD48Qut0PWCFu
zh06q2x/IrIBdZrEz6E6mnEXjQ4y48ra7htTnygAYQ5eT31alS4FA9rBn3BdQgQr
+OQX9kkLkvt8Q253trEA7V8lSWACwl/Mv9j1zGb77dfarGwi6UgUzEl1RaIx8rph
fv0VslrT5NViU1QfeJWZXRBLt6GU/BiPd4vbeqKueM54k1hRwBnDMXBOjJJ4UuJJ
7EpMtaNzeYVM4Qqs7kHBYUtjXjA6aVK1bfLpmtemMvGyh8ekW5jZI8goKJFLjGI4
I91c3w4SCu25STugERcD69WbM6ogTNfpqoEo+DiZgz7ObcsrFBLFiRcE5FlinN/+
tZUURbwHNYifj7lXZn5EF5sZa45zLC0bae8FzAblLr/ZXsJdi74Fh+A6ozIlAh4B
+5xIgLn2CHLU8gBUkSnhmzGO0GI0EjbZNtFNiqGau4JZaLlavJ/4wGmbk9Qbgo1u
UuL+QK/TDSlV1uGgxV08UKaKIwBrFjfQUS52Qr4QENP6yTo/h9RbmnXuaIwipo40
//Q0t/1sRh0R/fKzndxYWRE2uqsyN1sLY8Xw5WrmFgQjTWy46lqL2gAU/ae6o/k7
05BmeBPcM0qlSPkOxyMwQ9O1aKMfcmIyE1hdWiInaf+uQErQ1cj1Za9MTUgbyleV
n57BmxqKC3tCCiIITfSxHxW52HtkOs5KknbUVRoYGzlri5h9+yVDhzvaM2JChaUI
jdGIbR2BEbdd3bFOjRctz0b4niRj64FUoM5k/QQb2Td4oWrSAb56K7vkb6FjLdEw
5FG9VCDzjCub2wDjXQ6BH50+ra0x3kMCERf8fsJKtP3xGtO3Pm1lvslMTKSgC7Tn
j24EWMqjbPfs6Pd9up142eJUvEokBFDmYeAQAVMs5/zR2fz7zrFaPgf4wsWIeIfK
HcgkYMZhG6D8fj5FRPQ8V4BZdXPUf8DjAsT9zCYGKkp4dpReXfOozB3swAVtZABd
HG4bl2zDLpTtCunbt6/USc2sJte/K2DwhtrfEz08TemfrID1NvWveuSQ8YGj9q9n
yx+PV2/gFFHBJlVnqGJGQBeFPDFHriObq62ZqnOJ4S2l8io6dD2fxZ/3w2eLWGn3
9mIM/hD4AeK01ZHEnztjiDo4Fg3cIUJOyz9NFyW6jV4wf5Pdeyk4tECAIfCTNdN0
9WVPnfgGqsNv2/APf+SoZ5vukjkydlZ6CME6RVD6PY5iG3BLAYGr1o2dtFFWP0XF
XAY1KWEJKrQ8U3W6lo/PrucAh/UYYMWn/1XkM5LJ/a6s89U/UjZR6j8qz9KhsxnV
KNfgUnIB4sNlbv3EGTQa5AsqFkQBaVK7nsJSTphNjbb/TTT+kcx75nTwdh2bOTo0
r+qDdvyWfp3iQsXRPm7FVIZtjpCyusH9/qnNO8+JfZZRe2UCcN/riXJl50d1FuDs
qPFcx27d8ZTVtIkZ2nOrAW3Kq07d+Jm776TezjhrAO7Iwr9OXgVif+PPxubuDI3u
n9diUwQ7oTdhvuAycVvwxWP7N7MMlsz6KKsrYabhHR44XRXAt2Sy+jbEGKmIcXH/
JXbvLxgMlS/3PcqnCkwHjuSjmwuaArXNV3uaSeW6/bNc6xUocsOJj+vrNMxEoOd6
ejZea2k68Ahwb4WWL7S8gWS43rrOB9GGA3E5xZWrIwBid3VKBiwbVQsGMmr9j4ki
KzojG4MYjHTMHiXIGdKNA47B7AcOaY8oEc3OXqz4qU3Hk5EDCrt0aPFk7iQAhfwH
Yj9DlzlHwFSfQlVICwrUdZAwmPKJtUojslhkAAcSd5+DDyBlUBp/Y151KmIl12tl
T2WRYn3sZUe9PgLbmCh5nCV4NhVLtEPpWvoqFvNGGHly6x208RAtfzrupKxs/E4S
xUv2HUzU5rlvgXT3F4d1DC8Nyeh7HTmib/d7n0RNh3uZ6yOez25jnebJ2R+UhVWZ
V/2eVEHXXN9fTuJJJOCbnDCo88fP/oipfwAFZAS/gOZryAYfZ+rqz4BMDbFbRD/c
MM74/XFl1t39C08Cmlcg5VlWHY0lCMpxu4/X7wGefkz28kRVT+seQobjZGz95qf7
OzR1vVx20lYvvzi3ibSlv6+ZdswX3jL0GK1HOZDvFEwVbPQtVeOhfM+8ZIN6+Da5
rG7/sImcDQqFlk34xLxHAs3wy0bCOmKWWyEVE45ZObAPiHylb62anAPwMfqTt0/R
85uiRtI1IaI4fITLivMjog4mK9jrU0gC30wgTXyneSxmsvjumxfonESHpx0uKIbJ
reMFQX+dLxsQlJ0nMJolaacshV6W4LurT+5VyotXVI+h+kr5N4ld87VAb4Mlqth4
7GY+KkHNWGRjMXFEKA8Q2YKGwmdkH6IRnfgetWIwsLnPzLn5mmYb/6kLDOLA3N/c
0WOnv9WnGBV3xysAxcD9uOvCB9nwhnev72Ut76ShkB5p3qGCJiR5BzlXdBG0AyOb
cSu7nTKBnkqlP300SE0xSoWYhYmbzdZO1QoZvDDOtqo2x1UyvoQdjsyUXpJ/hK+C
HjStmezUxZriFEIXnJpGIbMCbfYrTuRsde5o+eTtDEg/DVzj/LHEBtuEf78TTAUl
KczEmOvKJ0t1NBClS0BuX67yRUrSAmuqbqKVSRUmJXuMQA0ctGh7/l6qFyqM3Zp+
Vd3+iXIZo3ccUP0VV6lXiaiBwrXvmsPiFKQ5CIoXBMOu68/YmR5RmiJlic9SciCH
Y+CsC9bHjm45EUUIVPywuU73lDULfK1dhwvt30bMP+QU6jEddfd0dXuP7nhma4bO
douwNEHX4Z70P8hW1chVI2TExfHpZSOVPIeHOQNXApF6gGkQLUCLl9B36UmgpR/R
k2rCjYxUJmUSj6M9CMVSW+NVPb3j/V+ZYXTM3lmVGLLK9cZyiYb+/WlNekOu0Sx1
DQdrbe4vrSbIs/rIwj46ya7FBqBzLKbgi4X9z2E2h99ODITOROvcg/3fWnq/E7Sk
lM62sm806h1ODY70BgvQjxwa5XBMX9x0q4UuGC7lRGEFLvqVqNKHOgtrMajP91a+
FKnaF9DY9X/gaQuJSNOgylufohy+JRTABaBW8eclpv9xbRwa+fVpCDRHqXpPOr+t
xslMoLsQSS3wMVQZwaWyQrnigpADRO4lNbHIm/Ec9QSQsLIrVvnvJvB0e8lxCO7b
xUkWk8GasI2v+GYlaUw3lX4H1Xstn4bQA/LIiLfA+uOZRqfyoaR/7Giq0E3bDp3I
yT1b27z7IjusfwgB7/r3re9AcZbvIRFEV+rfDRKWh+uPcYPp+5SYsYv5TvbsJSUO
lKVOPP+geBID/Olisb4iXZRRf1oNT4i6Wh3yViTAB8lHlIKZmOPv1t6JUzwQmERe
b0lJnOcIRNQzoAX4ZKgO65ut35NuHgRpQABqzCVjYygT+Egkps/y5hEpfxQU4xx0
BmUsOcEly69D0d3K9wr4qdaxQwZ8U9hKBEmF5FAzBVXkqCmtoeW/sEgFiDVm6yVz
s42cfgBX5ET4CpMkvVB4qTyaChy4Y3PRM2OMA/kHeH+68No7deDaYl/2rqch/lQh
4cvEwfC5iI2CRzSiojMijAaSAILlolXXuDWsgzpmvczEGKtNjTQCy+rpy74RUxNo
5PBg6JXkO5DKnExUIophXx9Ky0ptD0//YqwH7e5MckwPjHBneV4d791livylk7HW
Mnp+xbr73aorXW5WEoH9ydqLqMyPDwRHRe0y9aU9bxbx0+R28eiDTj6h1V053Nf/
DmsLFnPlYvbF/45koeqAzU2N9D0DBNrEOm2e5TxJ8kOFUk15DbILcF9zEuoDkSw0
F3yXLT4gOUwpMitOP3iR3YRIfD6Klici6UDrlnS+39HNdGeJssOEktXK6bcohmfz
HY8O7j7n6XJ0/VFxs/7OodTYSEA5ZWh809h1LytfT0f6sfdEvm2Dx/qt9Mqam6Tz
jajm5ou70vPRWveKMaWxb7CT+F/dqikLzXR5NC1GbACSF5YpzK6M8UzuUmaP/uqs
fsAHlgAE4mbEVZI1NF0LCW8GQqxJF2M1dOhPwOPAu+cjsADq2Db6zliVdfAwMCH7
EU3Z1937x+d580wTZ55Nb7z2HnELI7oU9vxH5EgWRGDID7GOiUsJY6kVBVNvhNlF
A5Nwa5KLE16yxTCLNtMtS5zZ0flHE+QLO5jzYmnFnQaRtCCQ6D4ub53bt5WC7HwT
wM/caGBH+WV5qFQVD7LmrLB+msoY+/nX308yhxUVWGozDN4ksvae6wqXWFIFi/vV
mUFg2IyraizskQC+uz2rD9cXfIK2pmzUUTNzQdPEXkKI+PvCXyukO7N4wfaiZJt2
tpm6lmdUbuX9Ff2J6wJv8AJD4P/NJJYXDoBOE2sgEuQBpb5akeukm/P4FP2DA/Mu
tDnye5r4WyZY5xhtmoKB1nBmljQRZ0BAXg8OV4B2jelq7SEfkAVUj8+f4lUIUoMR
qsPZKpn8l3+6dYDdorE2+mNW79NG0p4h5fRuuQpwCmGliCyy9djWuFEs4Pu3gsXD
2YkjJ+y1t7ZmtUyufOqCui/0+z3Qb5ySUQoct02mxXWP8BdIsq70qW1Keb7NHr1U
5hIA/bgTp+mfbsSPlulDNsqzd3Qy0mU7CNZ6tCRJHwKJClvJeQbjA+o8k3vzaTFb
Nke0b8IAqWVhk90jtRzNnjkUk+xCtGXamwymdPNtVynIfXuD0BL0r7wgWCEizs7a
47k4VPElmBDM8tDIsTMswnAuN4yNTM6lyGwl0ipzkBRWynKbO/cnamQqNcSLQj2J
EZj19yH0J3iNc9Vuq7TUnhJgjIpGvV0NTjF6hc6ymhoV+LTU7aa7FsjqTzERxXic
1Hqs1mDBmtR1uvB3kl8XLiuNPQQJ5TBRSBbkWl3+u0s9ikoZF7PfbKCXnIzKwBFp
ZDd5HGtPzRGrAwUQZbCERgFo3WyM9fFoy/jRYDztqggXU67zLnTRxjuiXDgVS7Sj
QS6YusHSoLaueP0BQ5krR2EgwF+1hcyiGM6BSen9k0l2CHEoxiVgz4Y0pGBA/gaq
Ug5GHXUp9b+iaPyC8zGzVxmrq+e+AZWqbS2hMTm9Eb3HQEgWBeW05P7MYOvrKxu1
VFmlQU5ek25lGq+WokI8deM3tgQP+5d63nj7geCKP9SbaANfIhlWyZFPpNyXzk/8
inJyAnfs3G1WARRjDG4G3tPdkCsKPa+agkAYKDss3VTQFbnPUibwKUPTBsjikW8h
PycqcJdkxQWfVfp3lPq0rg==
`protect END_PROTECTED
