`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7JlxKnRd+o97rfT1T8vj7T+Q+z5pm9AxqCEzbCtpwIxYjKxKL1SBBTDmaY7vlWh
FXVIDFxDI3VmWZbGY6J/aUiYoEJzR1DgUq48hAuJWXLRTt7AbGCKYQ71oYe5Q+VH
JEGIWVN4axUeHRFEwbIjeheiS6zkVzkoO/zFIPBZkBeIjvifS3+antLfQkNZOpC3
NxU5yHaP6qlWVcLoK8lGZPtfPPpmplaMpwNJe5xvNOV6lTgXwe6gDAbry0uA4ZTb
hOGRl4qRej1z12J+TVxqvq4zgdjyq3bIddvpSKbn2NMoFUjny0uUpjkfhS5ZNUs7
g7tdPL3hP2Tiafd/Lp2UqbS96o/rkya9K36Wr/kHaQ/rbZlARJWpOaStvJqc4ShA
SQZhgyhpsCKVrd4x2VBtrEBaPoD/UYsyjfY426xxZtHwAIRIIdEvIh0uN591x7TZ
9I8xi0g0uKtEzOm7yKt1VfiNSoAiF8dA0bYzfm0V3jxn0P9SZshavt9jUSCgd6zA
yTp+NAp2UwEbnBVzfLY3Xa6KUnri7kqBHu4dEeOyjUXPg47Sk1//mSXjrH7aX18z
F3XruZAzrpPDDzs20cXzDDPRzjaTpKEcFBoNOSgxdfq4/nPPZhhRUfdCx9sFKNS1
7D/O/DsrQZwprUOuVJCnexy21YAI9KrNlkq6VbtuP8raWIDunkA5hJGFsShmnST7
xSpSZSsNS5xn61CDYYvB6gyRRe9w3nFODVjAqXqk6KOsn05q04MZ0pSFX4SPvYsJ
V+gy1Vt+nXoaxPAQoMhfAyl14Iw7H2ePA2h1AY0aGOGAyHSQ9bcgfeDgfcTD2Qlr
lLkoGTGAwxdX1QK4wc+CW2lD5yeFq14VJEzeHLX8I40hlYBsoYShfx16FqqkcABD
XcTVN44xDrpxaoWBUAliRuFQYbnt1FSNnrum/m6AjWBlxKjdLWSwpaFo6D9HkKka
6LZQMooE4NqE4o+zTBJFlcfHfM+OTUK6bf/rzKohUmiWysce4RrwfLU1DY1yRchP
CmHR2xkHxiWz8X+TBWhrGp8b8jTzYr9OFLkVXTSMQFQwB6MKSNfv8zFpyg4rXaIk
xGoKhfzdkF0wpe3IGdfxS6ydneO6tW2vJs+1JCusrd0EzCgrs8fSVnBsFdwdsgwG
YunknXDhyrgw/nyaHL/D2jiX/JkG8zeFtSWwCfplS06j1a/aBXcT5iYTukkW4lPF
JYFtZAjBiZWeunJoJiUIDa4qBM9sFXm3zVPMklHrXD30mJeVy8NFz1HpmF/2uYQH
xWGaiAJ9dU7du5M69aQphGd3I9LdQsSFjg6MhAzRWycJ3ZU+wcCHImcKauXv1DWt
0C668pcI6Lc51ift/HWKsKWjqt1aOHqJbebalT+bgScWNr8KXg402nnZMZUi21FG
aH+cPv15ruY9pVPY6qMFOzSROYf8pbr7GvEpoUAMT8jy5iOGUItsNBcxCstoNl/S
Zb+ZvHH+J90Zi/JU2m3rpgtD1x3s2lmb3NR8Vmyhk9jRnsHwSTMVGdoQ919c4+5g
DSRI0WDtv7gpjKITgG8v4fqGXzp4pxnOvtjwIlIt2Wl5lehgfeMEu0yZVOEkc8ig
oluT9gMtZGxCdhxWpWWBdZE1smUyXBog6uCITl/W6ua9Gr7ToZRzxNXZpqItw42i
rytgOtPgYrKwzt8Ui5OyhJOZxm6ZtYOidtghoLgB6H6yhmYWBFvpK0aCOQLe7aCD
4VNrzL0//05jeEvAxT3D5PwB+YSVl0PNa6L5+5qZy21xp5e2k2z4f8IdUSyb+l0d
xDE7ikRKgiuesdPqGgNL7UsDi47EkqvltpBGRuNF6WW7j+kFCzrLcRXVE+G2SPBJ
EO5CbOsU9nOEPx3ccwbr8NWVTZxLj7I5cyW4i8k1y0TebwpXVJjIfnSBt9kx3W0M
Wi6UoRcF/1+3OTj2CFOqrlTdKdRvP3BwWwy0lH26OjSEA1qVLsykuuTU8285YBvf
8MsVsx6vCjTw2zbFg7xjHZiUThfH5pAlOkgMCP/wpABSfW4+JpUwQYCNhK/trhZo
zy13aStM7KgYj+enmXd17HZm3dzU3FSVqGLIlgRDunUFi04XEocDXfaMoYY1+oPC
/vZrqVSuZQF7pmmljtdAzEbhH1I1oX64Gyyvtm2K65LS1rEasReEjcV71fl6i+UR
N08Qelkv7Fh4Xnuf+NRcz/3c6+OImIe9fB+m3kBJbfwYUGOss6iBn2/qOMzzXfme
SRc60a9/qIxee34yGnTmtyIkjn4EZGTdeOFcToWPHcMekQgkJeXw0VIAoxaBPfFM
xmbvpeGYO6FwimVniCEgRBKH/0okoi+v764hCGoIchhtkGGtccDG3pZcnu5HUks3
P00v0l7so3MRZbrAxC4sUhxKHSdjvkQu2t4VSdBbiBVD7MNOzTMuYri6PflqXkno
ypHUcX7pSnjIHCfl5ZisoZ6OGM07UdDdgnaADvv6og1+6ayfTIxxOSQJSfbY24p+
n5uqRXEi4MLbxKsQ5/HSGmnPI7nw919n8Rn6XNRUXt8=
`protect END_PROTECTED
