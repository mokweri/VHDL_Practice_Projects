`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vEiEig/gKipupauTxmIAHzTb11EaB/TNkMjl46Q+1IiGonV8M0z2nfyZrtReqJrR
TL9kMwNOdNN29ntikUapossSINasX2hzZMaUn3a5gT6DtjxYyA1Dw2RdfsmgLQHH
r2RKHaOkyCFIoG2xXoDcLWDtGptCpBNZBhYrnpIcpAH84O6iuj20EaCwEwhPyRcY
OWkDvbuqFweVN9XB/ICcnmrpH0pn5yHkr3EXGIzWRM4fi5cqX2emMq1Otr1sNezW
z46gPREefBVG6juGqGEpqVdlSOZNtdeo0VoReN0oR9CxSyIOwAkl1eiDFhFw6ahj
W2v59HPObasbyIYA+pX6oAHscuDutDqQcN1ZQueb9LhdNYp5ie0jOJoGRb7Z3mBx
0ipup75xxiddbscccBpLC/63wFYo6G6M7BKFUnhodt2A46cEtV3K1zkWiVQtEg3w
z5YYGjy0X2UOec7GQU1q4OjN5BnNLJYaCMP9ORqzCDzKG15fQFubBXO2ZH6jo5bz
drB75q0GWzzj2YJ4h3vhNWphRr6s8WyuazYMJIpG6oaxHEJLHDomsWx8iws15HLN
nEveZ2iFAIh8EYWUrQCS+1VgqFlqOd4bbi9sK3h9oTWP8370UM5Hqj7NSn6siVDK
FkbuZoviRATFLkBUSPTTvbtBC67lqc0vp/T5pvmLGEjhRv0TNQK3zbvIrN6U9sZG
hQGyPkDJ94MfyAhED2BuIOtBSQh4c2C6I7C2Y604ULE4FASl/EU5RW69fjVBV9CC
lrxLxMHlLISzKNvT6l2DI28qTD02trrYpOQHjMzOppov9iy1YYr4VPRK0CR/EGr9
rnKRMRF99sRqzMKwiE3/IFRK0ghgwbL4FCED69ta/QnGJe3q335FEWyHw/R9wN1r
S8J2fPZwuKoPj2Rb11M54ibI/A5e8PmbrJfwzZQvp9YIBs0BiIAIzBPKTOv8+q1s
+BpaF+mZ27X0Woq3pq94mz92qZXIksNa+m8Ydga1rxhsLrALP5PgC2cEutlZNUeC
2zU3M0I7lqitzC97RiqJq+d5VjzMMY//2DTTiQjAvO/lHWtKa1TdfRvOX2F6xvv9
v5yiujnopoC2A1himoXLJvh+00PrwWsqiQJ6zFDtuConDqqh54itBoYPRW/c9eoA
XdLQSnL1D6CBt9lwqvrrSfD9XPb55Chv+9uEY5R/IHIkL4sSoVCSpc+a+3aPXtPr
DM65Tw1A2yMeLyR37NrMT1N2TNNEDe1nT9EyXIiCfJBhMGb/HCq94hXmAcUuPDQK
ZccgajThuwxbTPJfnKzuDCROAGs+RBJ+iu/Wi9a+48pWSkgIWgCB1Eo3hEb5yxSK
LtDQpH1Yf6D41cs8Vzu2XCJ+NTQ/I2QaaCtrr+sHtTeFFV10IkaSHC8IeEyc9Azd
B2/DrMkplT7nCWf26iJF5bbPyJ1icvbfYriIZVNehSA0NTWxcKVC2E//aWEngTPK
12e1Loy92+yrIFiTdpKukbY29ogWFomTzVy81bwBpQtZil2lv6PjTuxychwwwFAQ
t4UUk6oD1Ss91EmSIJLVxNAxRSZ02wUaIVxZfXdkkOqCHmfzQ/d1DxHRAN5ZdRU/
SvVA4WtMdtFxPMvuCSWuXkT0TWy9gLhXw18ThUVkLM7Yen1u1s0rBIHkIHBkK3B3
Q871MLCWmwAtcgsEvHS4HanJVafAL70xBl7xNKL/eV51YEVsQpxD+ABazG+A3zz0
GXiYyAyQU+/zhqYCENtWsOamW+3MHBmZndFuhvm1ybANAzCB8Wm/ViidERDUcFM1
HtEMjMzseLNCEZw3uIOEcTrbkYCdtvaLsImrSpmOqk8=
`protect END_PROTECTED
