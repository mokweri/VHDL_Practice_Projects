`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3qpcFTykeZcTFsoi3WexT3m5SsA5myrilALYIyTAKYmPnBM7vo4FEeQOql+JFZf
7rJAWMIsQT2dACop/e4B1s2T9w04LARXZkq9DfymsjBAYrTE9z272rZF77OGTjrM
bbbJqW1gcHOr1fpTa9VZ4Mb58zK1k366nYfAAqLV467JdRSFuVOQArVDqmY52sLU
m13jc0U9pY06ITVwgBnXNVXMKeMosAiXA22Fw1aVZnOHJycj1lEgvdg9NaQL+lSh
8QuBfQQwAyLM8ddjIVvWXAXc2E9EIogg2Mww0n0ydc0DCImc+4wivqXNTVxnp7rr
vqqvRsqnZEbRQBo+Ted63SInpVRLGJMZHGd7S8skL1D8ckmnrScVtmJG3AtoXytU
n3tA5tjjsMVB222zNkA0YNsWaEpbikio4CYJRa0CthNrKZGQEy+kqqxTS0I5oqEw
WFVwvcKi+F7B9sztT7kZJSO/FrSQe0j+MdtlGHTxqQhTdFipg1EXGThfMR4UACy4
mpgR8Ce7jynP0erLT38v9J9SRa2wiHR/0TKYg9tB9rjejJQyfcfxiH1w4dAUEPCM
OtLvkSkls7WODifY21hJjkxFaPQqQdW8olKxNqMlJvtSiuHAQBzgLvHjXvE+cN5H
PqrOBbAUxfAdLRfCXccJHwirdRGGCJ+kHTRnVjDGKgavzOhJEUcZkHUlAg0mZa0G
Y5fFU/3ewCTegCzcuhOdFxY1GbgTbfe07iJqwV4Skwu6n9iYHjtXDrowf0ZdXutv
Tawh1n+Ic2fp8Nuyj+aq2IHxZx4MtlUgaI1NrIMq9ChGR5oM4XG3PwoRDTCLXljc
YjNUugn0sBtk0hngrn4K/r0UyCWBcq/J9O/C38r0yiTD2YM0t+VHxlmKW5xrBHE6
8vUOgCSWRZ8Wdw7n4OiPcXGWL5019n2ZKn9mGRo8sAQ+oVBPudTtlhnd59nQXLFb
qtblSgD/z540HgR9k33JT7yMmasoF08SlSostQQget+6+nBYKblRyM92ATaOlAkm
vMczybGC9epPlrJESBM0skktQTfFAe4g5cBNbivJC3C8i//GDVed8SVl4p5unxOA
lNUhoehwa5OFTlZ5w9VdbhW9gaV7B0Eg5HPO3BfrW2+IFeU2O4sXg4XPI0V/XV/q
Szbx/yi+1DeZ44DiZlxdPOUzc1F+mS7sCXHXepqou5WCpaitfgfsqUDVPLidT7ok
FVKvXWXD/4Q01UTfl4379WDHWhuE3R1/Devfi/dSMWFu4QJkfKORhUat/ynscux3
qdqrBGii2kLlDMKpzeY+d+H1PhB9KFM97Y3mW3SuvAY7u69AcMDlSJGVm+F0ig47
bQiqQd++UDo+jb2FZqKRXQNo9ejmnYIC6llEe7bzxRuG6mZf20Wua0bdcUydLQjY
yjqtsWgEAygytDrvLEIE+YHe4LMLmTOh9Bglmh0T9iO+WCTjDcLnbAIrqcPJn6kE
IzQYeNclXlyaMJLB7Puf0Trs134A9GXqgTMLTaIxfLaxchIvXPThZu6w+X1qbDVK
MLtz7k3n3Koi/qPlQMMJwZVFhFdj1eHqx48zYyc8NX8Cr0HMu1kv70chSVf6TMEs
YAXy/Cs4oNXdl4XeXl7B7vcw2AycnfTNb0ter7I5bDUuYHzCKoFxz/tso7MbfhIt
Fu8QM+P9Tq3rv+9ZleyoNqxNr66sgBSEGBtAvQ6cD+TydwYdPU32tYVjIp225//K
DouNYH+EmrkhcgozD3bT6qzAMCBnj6fsXsNoIN62wZCCe8DwUMKBoblhUqIOMipp
/F7ujN3PUjzSrZYyqGm55rEuwktrmr1L/uwWfdaiiG/lTZNVCGoxl467eobxHB3b
43oLDnD+99mxcOCNX4gkvF14Y6ezzH/Qxo3M4osG9IUmTONM/1FHPSwaMhFo65ah
mPtpByG0UZp0NVcXw2nk67JWzudso5xq41l3b/q0ogmswE36aDVuskAOmWrtOh4X
HONJn8vxw/RY/UMS9qGhAOJrs10FRbN8g/96SkX5mNW9LRXYO8ATRYLLZGT7d+Vi
79TiDZkoYVlotmpIDh9ImZMVjPScMVED5TmWXSHRWub96dTTWhtgO3BgKYyscDAA
lKEdfCz9NKJNleofg3zfnKyws4IXBsfRl30gwvi7zB8ukTIUKeOXYEag6QytuwDS
Q6mgV1E/zWUEVy3FmVhh5Gu7HeL0OVMRmIRbymSNKRbfS/fcmiBAvapk8nr9Mj53
UoS7tZw3jSn600060oaHS2VaRlF7bW0L8VGqNNW7RoBNppiA0WXEvV5JZ0f2rXmr
kx37YPYOf6JmIwjBwK4MDbSdX2tAJTRQaQ1BwFoUzgHdCxUg9j2vWrs5fcvD1/E+
zodH5wp0D67MyNFLDVQHFXq+QTCvRI0Lk0FZbkfoEYOFZkqjoRSBYpEVVD/bXJ72
K96fHqfyo5SrflB1HmrL/NQovBFEdah2MVC9O6f2qVUMiaXL5TvE4fn+gRKq4hbT
CVX5T5shps32cjyaj+3DnWYx84/V91nFWOzHekOXxcv6FiVU24HjyrgVh/E3TM49
JIpHYgUD4mwzJaJPnG3TT5WQINIDzHc6xeI2UJRVlQBp4Cbzg+nOoradmgWBeVxK
xj+MZS6PYIOElm8eUe9faQ==
`protect END_PROTECTED
