`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ePq6ivd7aFJHmny17TeFliYG3FJfRNOlDmPCNUC2OCZwe+YH+C52GZ6JnXF4+oSQ
R6SNZ3cVxuyAMCq7SDJwrJCSRWtFbUoTkVzNPM6du6wg0SWo/mz1QCh9+HwHjAhS
nGMYtOVN0DPq410/MkOQiZ+HP3A8XJLnsHAmWHgf+0Eo6Q1JgEXnutsd5JbwTe4R
PMGFBof58eYdvQGpauP7dX79QtH9NqdcljbKBgEr8chiR8flONHm+Gh/inYYvYEY
nbOQ385ztx2bDZ3CT516+zYzjpx3+c0kIvAXek34IrqknUhG7sXSNvH7ZxUlT7F9
3oZSGkX3sTgGqXFAK8kHwo7hvO8cZHjmHKS28m8mx00iVdg44LgjqpTLVnUr233g
+R8k8HGmdGBEsTmzf7u4GPea64JWLSshJtRVxBP+6evgkc8KvFhc7GR7s8qA6NFp
eAHM/lBalAa0UzYEl5UlDcnAz1NUA7yPpLcn+EyZOhBuxoTA5YAbMXTMNXSrx5ZK
NKhotQhO3x8YuU1qGV2KWohJBGmnJVvVmGWzJrpq51zQjIO3abWDZ4uEQz1kg8Dj
wWlQ99/+MFCrd0h3sGSiC1w9UilHVqUtD3zq9xtMDnM+rKAIX4cASS+RJwzqQcwb
W+zjQ9259ChjB0TYGO+NK583l7KjbHCdCpjsqU9cPOHBwHJxsyRIuavK1zAOjMcc
GYF1+RSKT1pgnTVIz7z1EQurSDLVlvKGfZznNPyij1hDIO7owdbGGMsXjeVrQnLf
xqEdwmTOTgkWHEBXozeN2wETFdVD1D3i6DRyPuWcALzFIgHuDBR7yUF/g9O5uhvf
kijGbiCt1NzJpgAPBd7GRSJtfpCimLtGPkRtti0GPRv7xBvI5UJ+1jg3/40q9vrS
muI+ekhswKB9g61TICswxDYNqbha9K8fVBzSx71vjdsPAO+kS8zwtNW4vj8Y5NkK
0M9vcSHMYUHhcsqIeV6xo9NrL8U33Wh5uizQTcX1WGusynxGfl/yzGhukwELKWiz
FbF9vYeprLv4u9agWbegaUjf0VU/OS8B4ZM/rXvS7FL9TJNXCxx8dbg/b5VWNfs8
UMvG4iD/1R/CQagPuCDLELWIKo2peLGsGLH8gS+pAjBndlcJjddj6e7dSdMPIHHv
8JfkkL524TTXUcJeSagGFX7xDi9uaM5bshTmCHDeDW9JgmUVSZt9rJ7XHN1uX2dM
kl/DiC9g9D07UfQTawdcGf2HcVk4SvGE3fyj2sqEID81F+B0+urD0tIWUls3cvJS
g1MW0AvbXcO6IDzGZ9BdFYohgUyY4zCiD+3mjfpo1Iys8gS6rJVuQRXNLR7FhTGN
IKgEFsgKd2r3zXUXnd+dYBDWO40/Ufq2uoleKKI6AHOkx1b2AppDi2xRU7S6L/md
2HhQRtFg7owtEzp2nZ3sx9WoKJ53k2Cjo+nC1Cu6sS05mcrLgGjnbSL4tXpBb9hO
/Mucee1x2/1RKn+PTQpIwvc3rxpV2HrJrq0W9TklFbcrsb9WwvaeDL9pv9bgfGJM
H7h4TiIrj/pfg/uD6EueoNVWEdyFsxQ86SAY+zA8ZMcxN98jbrYK1RF01Rw7VbJa
jhFyn+/OvnWc5/fWElQGog9o8xmoE+b17JpISyMGg9qPW+hVCL6DCDX8jhFG0EeW
l+rf68yKdhrlUnKZLzMws5gQz5CUN2RQX+sXpPH7w32X1dD65M4fhE+tbMEc2fEu
UpJ2JaiIBuLKKfYp/s7EsiUO5oSnB3XYcawpFTB6F7hKCENlGgUyu66WUJjB8X5Z
WR6HXkpUv4FzE44HyjIATFZ0z8tY0Xj7pn/bATnNWywwjYYk1vyj8tP6woZVXLem
9xeps8ynXtJQmNC/tLVS8zgLy3eaFJnkA93DAuv4AVHluzHBcqVT161VRw7ogk9T
eAxPfEH9cUWkUn/ru5pjk8XwJk7t6rWRaS48nYL2uqsSsHmWosFMt6QN2KXjxSrO
g/VhdOW8o55TlytqZDeCIieIY5AhbxF7+6yggTJ5T4bHDE3nEol7Io/EU40WAcxu
gZUs05m2yAwpAIqat1l/f7nKKIb1J8d+7ZhrJyzpYLAdS/D13Rx/NbLRKiiC7ZX4
tp5oMFWtokvAiGXmP5D1cSDOdpY7xJieMswyzq0878f0lfTyxOsP+UxZaa+HbzEG
wFPa+JaJagTafhrq7U56e13RqY/B2+TxNaYnEt94t5K2Z7PHunNYaMPrZfsenX+7
B5lnnXR1MzAkzf8mNOkr29Eqdc6YZV2OOZLyNmrcxZwoJ3Kzo8PZKlhGFIanq5Vc
H8rvHoeZ0gbnOY3Ky+ChVaErBJr7hktoDNXnnRw0aOzLl9706tJQOzA8HxHOYsVr
2dXq3n9n8XLHGFygYXV4Qk3178Ny6IA1QKTuzjyQrfU1QtLL1v95H6seqXQ7RLGx
S6vSqOXuQVGa3a0wdTxuq48zMLEPOkwUCCyDapa6h3PwBh/2zyFA0V8wr7lcozT+
50o6YxmcS3rblC0l8DVMaSmj2BqOclKs69sWEnPB8OeeqBIpdnA/W3gDiRZLkWXf
vgotNZfXKYtvaPRTMrqaBT+qsoHYQsfMJk5F6eCGHjKGv92/b2ZXo9n83tcIcR53
n6ltEFjHzCmrUkQgxs5Ooq7jruIBgCEnZfgl9zcGmVMKIiExIDxqYg+tAWY1RC2p
Pr1USRO20F+mnJoEUA65Ui+Tw/NfGXeUQlnaW8Dk5nK7nITOtEsuR4G6C4Kd6h2e
4IIL2aVJUUHaiu8VfoiTWnj86/z2tAPBHzDYD4/ti5kR78bUO8A3lN048ibdX773
bcbu2OU2vBlwWz/EqqaO7wBES/Fn6qKesgbukAS9CD2pF28SOh54fTUuhLWrPdse
4TGGlG7bP5DgdCEStxdBn2c/TyERX0kA2xeBn5WRgq6HjLd1bfgMaVhsJeaX1Qk6
WzdkXpJYC8+xKMRe1TADyCtWsxvVhMHLWhYoJEbN8X8mM2qB6rutZ/mgcCibtlRn
XNE2vzO52bnNB+7J020TJw31+2iY658MdIJRs0MZrG4J80ykBsaydx5TB3ND19+K
ZXnNTuqZCO+5apfoinJp2sgORTpiimgFqhRx+BPRdWT4M6ff7DPd5dB4Xq373Bb4
j/9Yso0J8TqKu6QXs/bAitAhVziwV7QCNj2kqu5rr64/HhsNBHRv7bL+rnHe9QMl
6abWp5SRG0d+HcB+yK4uO1lSM+UmCfy6h81j1Sth4Cp0/8rxQM/wtKnYtm3nTHTp
IXBQ/2mFZWXOItBdc4StJLne+kb13v3Auc7Iq3OaniGu/HSM7EfeojhBahGju3PT
F8i3ZQYDOIO1/skUovKMCrW7nlKe5W6W1fwkT4C0+uC+P00ON9gNjJASkG7Vjg19
7iaQwE5JXzFEA9GnUMhzLVOQw3qIASLB2DjpNMcXbQSRU4/jd760lyM141P0gQbK
LHyEhfAMMgvllrSV+f2Cnz1id3g76JvqwjK/hmgeLbur2EtwHgW1NeMBQU0rsDyo
SLlDWTp2+MNs4AGYp3jO+EJ23fWguhNDmTt+2Wfyi3/FG4VpUbbz6NgSm+WkqXbW
ZJiCW3WZ1y2hE8Iicf5Oko2jrcsfzoJCprB9M6FhJT3nX9P6ldoG9ooCgNesM+8V
c7Kpycn08fR6f2nXibV6BElSs3ZlC3N3oyofdNyFykApgH7h15yP3HVa1eGkwX15
r2Rf7mMbXVMd6AZXhoCAMC3xjbPvqZWoyX2B346mYS19QyP7s0Y2LaY+YiykfZgA
cuwVYGU9x4l2Z0KfEbZ7CJWbi7ubZ840wN6UQM1VRvfoYdmD7vhCihsxdlvV8cdz
E89ateWrb9Rfk+FuqcoLhS98jNYadhKPiOmZnC/X/ZrWOS0xoYKX3jIxbBJj0Fvk
sPF3B3+rh1TH5HUOV6ShT5lXqMg6AIJsxdAWh4vslyZwt6BCtQF3lEkeYpXzz3n9
EaIAHCxOWNwUSwPb96USPd/7z6f/xzeJb4PvkbqTpIeyI7MsIDU1od7MEaJfq2A9
pOwKtyaa1YJX5q3V+FH/XT0WY3WdyVf/5w7Asvx0v28RuE5ABZ6ofR7lXkQIqWCl
rrEI2ANztQyYTL50uVBTBpNyaeWvEUTNRX7sc8mgGpgxIm8MBwsWYicbs0uxrvgv
vfsDMCGUsDLMpvd3ItuPjmrWL0qWA9xGBmxJlya0EuYiYQu1AqyR/I8IgP1JKbQO
tfXoZZbKcQja2Le6Y5mW0k9a99UTxRZSTUZbROiiXaGzV5+7Ob7hndQempG1Pm7f
zFs7r6qMDKc13YIZbjtge0kE1b3x7rpkKyd5OnUiUFQ7bKk9c6+7MMbqhZB3LArj
OFfS/09YZLlCKPMIcJnAtJaIS2v9euhzmXEDIR3BKohy6GSRJ7A/9tfNiB01DUYy
DszAagygCGTlF2O7rDDfM2DuSp+n0K7tCha2C/FAzJJInHEC0AkE9VEp7ytZ0giM
kuuVGBGFA/qSfVSgK+M02mr+L52FS+TRVptRZIHqbJ3nHk+e96aViQncmXAY3Uwy
RnOfsTM271mQNXUGylp8RBqfpeb6Z4OHZx4h3+QsbZKhgQHG3oHR1mykpG89ZD6T
tGiDbb4UlU5dB+0TDy4FZFO+clC5bSH6tGM7x7YIeqKZAGkAN8X1uhwoL+XhDWXg
lxvMkm1EHh3+r5+MiGNMPK82En5LBTMrIXN4WI2HbJpWZ6luGnifOUXB4TBOyTcQ
DfrRQg33NOlISMgIAq09vqawnjwtPIkHIAADAfuRCvYD3Bq7fSVGbybqLGOX0QhV
dCUrbSYe4OZZp26pEpqBHCNN502Pv2oThxyyAXAkT3ZKKeWA9hQuQ/CiUFFrhzUR
e8jii7BF7U2Y7n91Q2cv7qN9caJsH5ll16W1iNe2LYfaxb9PqAQVZ+gWiNwnIiJ6
VG/1PPLkFVw478BXMIlDrdECKpS2znTwwKeJBXnj3QXE1z6xjXb8X+QJ7nsyMSTC
kvQ+Q7dWA8tVsN/Mpg0aImCTK7XC79ICx1kICPGH4R4//NDyUFAfjIXgFKEa23St
mNUAkysA2U9RApCuZty4vQoMkmxnMVi8w6WxXE1mhaMhKO0cB7Ll0wZ0tsnha5mB
wfsRhqH76c64p4P52LIuVxkKVfFdYaYxsOhP6VFKa4MyS+y1wJv3PZvHBpaV0IwD
u3F956vnTvlkOdttTmQnIhaR+Q6s2h4ENINpaJOrlLAbW6eOH+v+smiQk8DY/s6E
HE51hiGueFV1PMNLCgxjB8MZScuX55P+Bd8kolx+AMPKUPrlXR3nEfpS11RlZS3K
yBdNxHMTsPQA7paqkUwokrtSegiWLdDeVZdo2QHWMGxybwU2WeEuHyu0/CYiyqVC
GPUA6C5p/9pZSR5QtaSjtLKxptcQOOenCct+5SZXBrGpkd4HfYufas/1kR5hH4iz
pv0E/lBv8XC8P7pFYxsVDcPMZg2L+ahpYjEqpDU3NKH3CEO+KoM7nMmNM755cjn2
AGPVfqjLMOvYVGh8gGC0veNRNq6om/b7Sr4vH9Rc1WwLItARztszwcGE43H8NuuG
GIa/ozmm0zun4d8eXpLHU7wvwgbElW/Xw6xaTBfIa4/wBBTXdIQ8ntVYN9rufPr8
KNxSYMSbhFAzG3skjPGF4fuBxoNxjgCIfw8GFwPz0RdGMpzB3r7wf5c0X3XKLU4s
e0iE20oltVGAPTQ1JhDLCzix9Wpyuh516GkABaq+42gxWjhVG7YtvtvSyGr19E9k
aSS4AyMachybtYzePTFvDPf1zCWHU7dBARC9gf+Z6XpOrf7gA4bkJik3sNlg/78W
bqo4Zbh+AH62Rl1HlJtZMRVOWIBMdwQqHtGAn3f2z9l3NCIsUzHLchGvv8BMpgY1
ZSR2fUA98Tv5VDDVp1ploSl7YE+dqFFPF82/Kzno6xkWV+z6E/b8VUymjaqj06aS
0bjtdh5duBIbPoIPBJhzy3gQ3pSYYtbk9FppLolfkbE6uUBa1TI9TSc3Ex2shXBT
wREr2mM35bMFH56tzlrwFs3klpcSaBr4kBXzDOm0d4nG+ZdcgK8KAkmQz+ie1bic
`protect END_PROTECTED
