`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJUT92Z9TdLeOF6F9lxRogqYU8WGUS9haLT2rQmFG6+3JEoYo8oLPbDORaKjYvDd
8KlxLMvYE8sjQxDUvZ1yRsut06kaSzQQjJVWmIP1h5ubQE9IC4dTtuzsr7QMv9Tr
+WMvEOixseL2zP8K3Cf6qDStpSIqeWPjUf/ZmtLrRz81Afuf3mxyazSqKhv6UsNF
RljSnVQKx4GHOr0uKRoLbBYj8TwFvE956taAaC6IsuYx5XhVUjp4JeauI9w7dmgl
dUsS6NYMniEuuZMCF29K+PFACCSy2NoRNxeMGnw66fj8Bgvma+CakG9Su54pe1bk
WIt1xfzsWq6AigMUJNbTV70kbWTORAhgUiPZEbeJZtpy7bHriU+U8Fj+w0Q/U65I
jBPShQiBxUrh5B1Dya/rPNOefdMRb1Jy6mD61cahSYgok1eyiBAWHUDycZCISDiD
cCj6G5iHdhM7nwZne8wYmkqCXX3bfzPE8PYgX/uircv1tNMX8+IYZ1QORJfy/olX
Rhx9ox8u6qpJWSbFQpiQSqbwrIWzyw03vUK7xTwmQecGbtcCtpxV3ZBBcM5gJRhy
9Binxfj/40bFPrkxZekIbxFJjVxvdOriy+cZy+7YLLYy7nEUujdRUqOyxd+KHJRp
O4atAdzUJhEJka4Te4S81LehpJKDDxBhv705z5DOyedc9oymCU80yrPTxcFWNrNt
O8bI4qyBFrKSILn0BovkatZmyGYHos/mX6Q4RBYZi548oKwBk6S5AoOPx7hFlp9H
WBHHKBjFwTC1QUSXm2myJl3eKzz+gF5Sq7OzB578kWeHhb2K4pjFqvko9ot8zL3m
+B2Ic1GH9BIFucY7oSnOWGcAN190B0PHhvdRWsBbrwjiAjRnYzhXOm9jsC6gGIQq
LKqzdhJdfyEWo5iCdoNkon4xqdNzUohrVNB+RYS5fSvkY8n0BpCMxZ7iyezYsIk4
RpfMIZOfGECrJUhk+JNyLDCak9d22UKpQtx+4oETHxcUOCUfeqd86LPpdKBamwl8
H9FUlpCEdCp8/Mb0FNKDq5J4KKqRANoDxvyHqOhkhO2jQs8DAPtmvleQKoDHELpn
38rdZrpLGnFxrJn1e5Uf/gb4mpX8bz2u176kxdJEUoLXLkfLnXDf8zAvpjKBWEzN
EAAmQaGamk0h7Dm/mc2xIH7ax50n1MNyehuIXdBcRId2MvKd2t2i8Xy2esVeMAqF
cZchzzVcZ/CFhosCFuvQ6xbLovuAg0nIye4KFeYqVbqhQrnGynGfsWX6kmZFkFwY
hmbfMWBwPaki5V8EMyJF36Z/weOL4B8H/QeH7v0yJJilxx6NLnobH0G+9xXrq+25
PADUICuDpP5nQvAA6dhnXwQGZpNf19V4DAX+t6ko9AvNpoB+51QFjBoWQ6Fmc+g/
I4GCyDRDUUgHxLjD0OHPwXQk+7wTsGS+I8BITbsA3/ayIgX0I60hBBbRoPCneRLg
hXey1zm1bBChE+EtHTmeRHP69gQs/UQGG+B2Jt3igw7PCi/UTWKcpfIkuAU1UxOs
4WGhZ4G1GQdOnv0u3GgxwLrvQEryFhn+HCUAGAwH4zLBvsyrYdGJa8nZaaLQPNar
kyvgiHIh72riPQf8vH/O29A8j62DZn7A3vmnbZxkrpQkfrV6HaEFIprhOcud9211
rgFCv2ncuZ5fjRfMLFSaxj0qD/hmbAzHz/Mde+kLnhwCP6wKEmUrKMXkaX2u3bY2
I/s1qq7wC4Zmda/8Rt6V1RLfR/sc6v38Xg0eCk6QjrrevdI0oTF6IxibdaXNhIDV
nfVdp+CxJ8oT7nASiAThCpbZiqoALU+LXgXLqkAI28FpV8/8sr1eaQpqIjI/YAro
IE3h42jrPfqrE5IVzRdaxnlTwiIK8KjJPYLAez8QH2zwWW3dnlW5UaZ6xQr+xEiU
mGhQePUkZ7dlHy5JnZIyCaZlUAOtNwkeiWd44zUc7wzXnGyjZaxhbqprKbQUj4fn
lbfHEVERmA63oLqbSbrPz8yjwejzYKRRQxRKNV/iNkGK4gdGPtrE72MI60srl5KM
/JFHUBjy08Iol0+1CIOZI3icmOGH2vf1pG/VHla04TNCivdY9a/7L1UKHkd6Xtub
oN6sZmeEmItRN4COaV9L3gDR5xc1lbVlf2Z/Yx2IQRUEoGyYGWujMz6PfFNQ/hh0
ZKhq48LL0H3EC3lA8IXW5de+D12r7IeNT5XJCx47KoOY0TBohS4vmpYpfcoHGe/1
H7yRRfKwlVY0H628YtcPSPlD5Sgo+mVXiEYRvdaXR+nUjF1Q/Pvw/sbMK8zGIJw3
Pt3xTo03WHk7r1ZwEYN5o7xerYmQWMZuG21Yv8mp6R4zxqLEEYq5lCIfEQwi8XON
f+/DNodGX/c1Q6gK25oHx3mzMWImO8oeyuN9mJUYuKpKrnX47NyQZu6G7ZuAvCHj
T4n3y7wuSVFn/ZIM6Vx68xFsBMIyBGVhx2Y9+t2Uhtu3uo8ks0JmoqcdnA7LI3G4
kAn+N1ZMrma2NMVUFGYKR5hG+LrG7yubYyHfqAtzozIu9m3HE/F7sFunF9NOnKZf
KUIIaNuETmCxcUpXD3G4Lk7qUBANCk3WOoILb8dVsrGosRrGx9CMgTUOiAiw4Thd
Iutm9uqINLStSNKM9yoLpWs5uVN1QrzI+XnXarFRcjVcrmiCMjWgYrfs5592NnCl
9PGdi6ETgISdjL0iFky+95jt213V9olYfouREPV3kqV7UVF5rOAJfzOsqE4sVo3k
lk9Y7ml9tTZ694Rxgtsj5L3EGddemAjMpQHsCKH7ty3500OCQ4ikdluYMEsrBEuE
gKopLEr4N04u6ILLpc+L5nKJ6tquUfK4SyhR+z5u8Vs5dzWhyS9C+xFv874iA+Bq
/oRTcv21eWyICy5a9TxF8IPp+qzwj2o+6q9Nm9kjoj0Un50N3I6e0QmV1SSz/dbQ
vFl0oxYzO+le4dp/+ToYg2B8QfIxP1erD4FMKwDf8WqQluqOdYbaXT5hMtq85Upu
ohGOyklbn/1x5qd/tXSZdNshcH3QTGhwi47ftljCxNaNhDiawU6n5hpuD5V7Ob2C
BpCOylxVSh0yoieNyrEmIBBq9BlXDXE6awe6ksQO+WCZ7YGeVn9+zmLgnbr3txMd
1mJN+iMtwvM8rpWQxLKjGq4F1qS9tNtg/bpgUqg/P5HIFEoVI0Ib8DPTXpiMaCbY
qfTZ0T251qPOiC2BeR8lnjC/RmYyYL8s7yUESDcHAgryRNtFGvriEOYV89XL8ToW
e8bJNGSdxdtElaz2T7MybH4POZZJ8Y8l1kc9WFM/9u3OMO7g/hjm16bL8yN0i4eW
rygvN+es+tAlZuptJbclcBUyIFJgmd621YOjhSuQVLYZ66Y1WR/WHsoFVCNwyH39
GhS3xx0bLlnL3G3N6Ad0a5LPimBQMh3/l9hZ6Z2U741qm9I9oai4Cc9jyGdZ/I9s
TJFBAyLjyAcWloyutYTErnVLuFrVXbEaeAaAlIpf7nFFfgb4b12Q9oYuOATr2xAr
`protect END_PROTECTED
