`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9Z2lAXNhXiICd68X7m0P/UIxnLss9hxEaMTDI7Ao5XRUhLrb8zreXlbLYefOh/L
AJN4vCW7A4zX/HQu6Bl58fA6WLVXHYqv0dWYwYWLYL/1LxxSSswqZiCBMtcFrvuO
DIPOzOwOHLFz6INi//q0qOqr/O6jaLB5TvnosAgVQhW7CcSVRtIoN28IDGqKCc1i
baaDMz9DpO5s/IttlX4HJGt18MCUJaAyoR/mNPI0/gqEBRS0EVjgwhBi1EUJQknR
1rDIsLtm11Ww6UrHS+IrrmhtnsSt8U3H7W8Q5XpC9i8BFkYjfx//aVRqLRg0z42b
Tu4CFpy2DFEPNAy31bZb/ga+yg+Ohlx/vD0qdF3uD+rCDZHj4T1zyBrwU62hSpfS
J0rVWTeEmaNzR2BF7ibNqAt/1ygV3JkEW+hHc7BLxA2NzPQd8EbTB+gQHw03Ak9K
v5KKWnIv6yyYhQvWRT2YXnM+jvm17cO5+Y61q30l1FF1jkBwyusn5SFjh0CgLYMl
1+BBy6vUwm3d6D6urSRhJjQbOrdIHPHLN2H4v4wwpHCk/bEad6HlHwwKLG4PuMFu
JBqvEkH+76TGaf4yoUBXq7ZA2c+0mYzCtx6Mt8S/NcCHHFTKHMyRi4J6xGoA2Xah
dC/hzO4lO5VS1hjWzvMu8EccK5xdp+5EGdcxjvfE1EBpBUM58NSXm+a6BInskJaQ
dAsO1kphABVUeXn/UWh9waOAye5XRx98GtI39X5KYHQiIZllzkudkblbnjCXCK71
eyzADENP/42BO+K4ddhNz4GUcb3n+PxCdYvaF9FgFECXJkiREvCdE/9Bl2m6ohF6
zpc6BQzGEICOSVEieQKhdDIkTjpdpI1aSONES9t07cLjgRgHTpthuus6QFrpEkKP
tazxBneLGhYnHkSHSHS9+o5GTY2IESw45IIZjB3o6bTZ6GEncLlVkQzb0X7hR2W4
JgXeB591QKE+Ji4Q7RrR/wLP00IYjPIPb8GC6eooRhAgrNOlZeUhh+7Ywm2rtFS0
XUqvLNbmL9ubEBmANMBfRzBl2/yWm0AUjlo2GtdBOMZx8FbRxNlLrSUlH359HHs9
WNKLbf6Yjonf9cF0NMEGLHP1u3UdH5J6yhzExSyYd/NmaAjGWvRtI6xr2mfLZbKa
mIyX3I1Yz+IJye0klsaGDY4YT0SJSQKWWo3TLonueOCGrKx9TpMM4Y80PO7fInHC
lEnPFczeNMZqLhsBZ/xb7suhZMnt48aBFYVzGIlm+l8pLfAH+XAggFGnWpBu86Mz
YS9qnLZncFZkAUCARwvaaFFzVHWcCRMMVCXYmlyEQwQb2IqTl7qtKctrGJFhLCwT
RW/MldYFVvEl51LPYM+512Ij6VEA2vkz1Jha8ZRDxDaz4ANA4KSPOvSRXfBLwRhH
XKp8vpkXx6GpEHPfsuYtxkPjIOEfeODNdEs818hMBPvl/jEAANqQ42C8DYNLVoLq
/V+w+GW/eak6o9Y4NI2AFiZmWCdl4gNwEXuOFkNDpYT1v1F7ES6tJBdSvuJA9TpG
BSNSdUMOYWTmzkCvJqy4ZFYMQZPYNAn18SXjVcOUOVIax92dsVDu2YewWUv6t+Qg
1Ovo3TMiUG8unJqCqbYEzGrBZcKyJV3IVzCEf2sq1Qe94GV1n2pRNQEnlt2+FD9D
fJgT+fym5cEeGC3vo209dvfwidc3ztW19rdKkxVL2fZNwspRakdIbVNIRug5DvOq
1pSqQO3kPYbiL7+7AHmZQM8ijH7bSYGpYu4FJ/UpLK68kY7VQcBgnWz5G4cZhzM0
Bghho/3R3Gx1jHGf2e3kEDXFr3XnrEZ2d8prj+ougcmHYHKZRoWsiSKO8cFpR2i3
j45pr8WRPzzVBMHOoKImKoC/XCwtzlZ+rp5yDhSkXFskYtWTjjEem2oUTBSZM6ky
nigLHXEDGMqTaUJcHb+eMZ48FWsD0BYXT/1hecmsD27WE/a2D9lxMbPWI9K95wkU
QOQfziCm7x462/KskFTyeSuSZ9qtvD+J8HOzJm/VRX55RtJ9Ym0cSkiVUJbPee2I
seJ8CitaM4m/AI40Bc1GfK2tAOVQchPqY/D6yvTjN4I70iBSdqsl/TxN2VxG3+t6
ALd83rLlARHS4tt4ctcQDle44Ur46X3eRnDVA/41K4f8ODFM/HCHLxnoeWqJIHWb
6rCPHlpaqOV+PzmJK3wfRYYaeHnSal2IWppnckeA3V/B2SrTdhHHDjWkot0Uhcp9
L3SYp190wwq6HvmJQ0HqEA==
`protect END_PROTECTED
