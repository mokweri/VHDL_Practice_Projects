`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cbp78AkRYmsKCpiBsaUYWKeLV5ySglsM+JsNxpRSIxLWQgLbLki7GzTBAPUcRAEO
NNoPlN7FKIcXDJ8RbllmN+iM0fXO3L6r8w5p/Sh4CbNxUvRgvuWn/Y5QES2BZZS8
Py/IYr7akDtmw8M53F7qKcadRBLnlOqLQP+sMEgCcrmJWfZZhr89wRfHUNJoXgZ8
c/tPSuPKim8AHMYYpIVoxdzmrSdDVJRVBS2yX7rOx4gFhX+HD1njdle/LJmC3+HL
US1Uk+i9U2IG099mc3FiugmsNU25N74Et2hoL+NjIaowuzvv1yWbhtlWJyS775KN
QCI7VoS4qxGEgt6SPcf/yOF5dWcqtuPs0qgJNco8+TLQho2W6008edXiU5ns0aFF
3gG+FjSvEhsoC995gSBUiS++yIvIa6U+jsImIAIR7lH+FLlO791IICzWKV1h14AX
EG/ZiI5z859so9ZC50X4QJFoNxl9cSTJfzCPqFtMeixAJvRVkrWHeK2F7JoA4ZFd
i+7C71GkX5kU1O+QZWtYD+Y+Jsv3l82wO+jEw+IYu5cbw5+X+Ktx0F6IknpqL7+R
T+jx94ngmQhwSiUWSXH5DvioMlY5cJItlwqtf60aJnUHxtHRUbCP68Gdky/x4ExI
iH6bnEZp4x/TG8kUet9QjnR7YN89sPAjO+saxgytAoiA7TxAun0Ul82XxrikRjBd
SZSc/XfkoKkb51QbBamQ4nnS0iWQ029gPbkMh9YblNuvW30z41exKwjqH0a6kJRk
nF3E1GGm5f+h9e2T49JFOzmbFyTB36fGzviZpraV4zTC1NW0hDbUqL9kkonJdtii
KVta4VDywyV+2e33Zrs3NbTWxIHEag/390IuT3c9+0TFrFmVGsU2mXNn+sSpuDd2
lyHZUqqj2h1Cq16/9tIQxsAhKH0CDdeflDSev2tRprktHVLfbrfouMtOXUrNCj5m
3ZRf1FtB1Hv0xlMS6DZl2bIQA51SNhs84LR49B3r4gSUmQrrNlGI8DPRT49hlpKn
q5qXb6Mzjl4BNNdM/tEc5Inj5yb9y6vraELpfvGiBiJSQqeBvwU7q75B/+pfJTC6
l+TbTPPr18a6zUWqZGeawg==
`protect END_PROTECTED
