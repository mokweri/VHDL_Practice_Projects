`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6MEZwdmks+Iv/9So82TWVljjbXKiAKpYGDkgotDuW/4rWpo2Spm29hGC1JHX9lp
oKEOOWqe12+SFTzNwiDtGnREkqTEJX0w7BGrKMv2OJ/8UCb5SJaidUQbXRe0+yEO
QgbjY8eJQfH/5KyWhvy+tZViJRy5930gUI11Mhn091gpq2H3SVjrgZzmfb5X7m0Z
lmv/mwXcuGEpblC1my6vn9zNHwWJxP2rIAtSsZFBL//L9mJTrKeZCa1umyI3XEbA
ERpCCM3iYyU4V8PVvuc7dVhGIJNCdfNbu+PVgNUioYfbBqjmJ/O61sUlKA0LHDyp
FZ8/7qCytB74REjj2nMJl2qLGHnaIPBo1IOfs5ZYyS7HvZDCrsQ7gNMa1xxKAp5l
BUXFdc8BLN6Fm8098ljc5UTBJ3MyQO1zgZ+bboFpztV8GOWGx+L3Wa+E4MA/aRKZ
xnk0z0xBy/3Nhn2rQPann8Q5DfUMmjoRItrWaIw01qhskiQfN4KTc+HFBM9ztCWP
mKW88XTAGi1oMqCtT4c6gStah4dM6yAau2rH5s/p3QOWPQKb9Ls/mgy2kmL/Z+Ef
pRlwQOJlUF7+EEYMlRhLDyDJCzHhORiLkZkLLCdYMfWGgkkWbTUA1uRmNz8unrdn
efGQQ5ujsX4SnZZw9dZ82X+vVDcX0DdG2xsoKXs1Su85eLWLvdvY6+pKJnuZewE8
ykBD4BwIEN6PXICMu+vvqj2U9+cXcW5FOHJ7IFVgY6Z8Gu89sdu23IefTJMUuMY4
O5yBnlmFQbmuo/2KwyppaOdfiHMNpatVK328T3cmyaZE5VVaO5GJ44o9W/0q0XVd
vQsFoTwSuZh2PGPI15T5xo1MRKXMvy4aRSiuRXIyhBKV4e8EFZnVcv2MNXnkerPl
/yKPUlpgkzSkZjO0p1Z9eX42kc5RhXKP6hpyp+nX25RQKHYLJxED8ml+kVyJf/zh
RfflnLTQvfAnA9Td2OUWlqc45EVFkdNJD8QfuOQ/FQXIOBGOSYd9CUTIkb59+o1a
EBK82CGW8Jc6ZKzLhqOjcGSvou9uhkwfV0R/iZrN7zQz5z/sddaagcv9kEVeUp/W
jcEJ2106nn6n29hyDdv/Up19+6PNrlAZClSRYqsagmiIiG5nIcW+fpAT7UxPcKrt
MvOhf3Y7tcP27VzcI3oCD3DTHn5bERfdP+Yn+9Tcq0CD9EZUfx/PYc9SNUgV6Ke2
DfYyMaNYsmpMo7nRFW4D51Bbe4aUgONROz7Xu97O0dHYtoVIBUl70kJqZRvKrD/S
A/QwknjrdW2OtxlNyHTQPOS7fyA/aD88MaNBbbnnqFGuDbMLO11GZwj2rHWf5J9O
Y9YN1ZpPHAgCYTA8tJ32/9n2AejuKAU80JSPc6flpTw7ZONxfTrFRR6BEu1aeCR/
fwPVEku48QPH23JBq5g/OjTH495bIAopA8EVP5j5d3h9EGoLTmDV0WdNL9ngduYB
K7EkpxJ0h2wGM7GeKEsLyLwQmYAp1M+AvG2hIe4PIN4N68hxFG6BVsT0AluMEu2p
6Loa9wbWBYLi4RarsCEtavSYKlOf1JryT8ybh93ROhOvY6FlSox1inC9jf0rblwW
fqQqPegTEQiWe7B7TjWS0sUexS12GRg//dRYJg11vMVVuQcgAqBjRypCfcc50QZx
xiq6XUgOKicqbonIn7fF17CZeuqMN7tDw33/ylM2dA4WY6caWJb0I1Pq01yFCy7C
yzcKeFiA8c/7ptsOutGsr6Ia/4AB1ohkdnH1myyoRdIYppRkpkASE+nVkQp1oaw/
btCoDF9mMHZeBzVCxAxCfj/RMSOILRnArxyuMTo4NiBqMp58T1LJ7T5YBNHiu96T
F674E7SZVG1CvGLMmP2W5llVdhy8qnzVXhHI+nZqUp+MXw6I4csjcIDCqZ9OSFTv
eGDGKVx802dE9n1BT47XVp6d6noRP4P8IjL/pOyHQYLjK2+dIGxxqM7x7na8ST/C
LkUIM5/g2B+PQaM1XgYiCA6cTA+6q1c2wzQ61bI+QJwgRAxTK8UhfoCGm8dGUdz2
c/sPhl96dqtPzBgMn2zmANnKGV++cxD7RE/mtjNa6XJ4COSrSeXIfYBdSRlfQuHa
7Zi2Z7ovN1d/S1Qvljjex209CCF+xZisuAedPs8oV/G1hk9VmB7qSOzpJkM9CKdA
XSG3Bb8q40sz6WoHWs/LHYXgmsQTUxCW7S/5WIRMlaWY/YzLqrBRqHDywDXpOVXP
yWYg/CFrrIm6nvXano2/NqurjrzbJ4bxqO30+Ex37RB4LZutCjRRDxlmqaTGBrIf
qNOBnZOYEncefxpgwT8bZHsPRExIB5olPExD1DS9V1e+NBS1fHWyG2IQ4dvuG6FA
iQTp3nrgm0lqtvDFP6pivOz0C/Djg5vOvqCvnekcF0K6RZYJhESyDIuxeDpUU8Hu
wYlprPDQh763ioBFCxKi3NocL4SiNDZ6ieLQhJt5Zq1xvFYWs0lQF9fq3Ec7TAvz
zEWW8vStK68bbKdK069liKxV0TXBpyjkb55TJboZBYpvlK5JcHA9oCL1uMl4exCH
+m0fjIXz3GTVi79HCkohkHizUgFlEhCCLYSaPfKVaPd7Lqe5arHQ3+IqBlC8tyAJ
VHhoAifC6QNbqRRTbq1MiqENsZDpBGrI/Xj5F/ueLkZxezzFAEEFzbv/VVm6awBi
IeEFx8rF2Xfsb5JvVRKeZjq/KYQ61UOTq82lm473jCbE94YaC1Vk5BmEXjIgw/tQ
9uNSIQGnN3lSFzemcXPnRQ/ZVzSI4phN0iLbxlZz/q8c8TMmouVDXBLZxn6NlfwL
2OQOIMEw6FDBdzSARKj2b6p1KEswaTtYK3jE6g2P2AEIuF9EnDd3I80oLyBt+7YW
7I7L2nzLa6ugbEeYereW4i7Wn8Ty5tVogd2z65iNGUsekFYgG9uhiBMCxENMu5xl
x85Yw4ZLurs1i6R6jTd8uqIbWc9OrPyws9yILDi2eMLqp8xEck8whsYIPIn1tQAx
Awma3rUXZHYxp3uoHJUViuTrJDNLJwNsfB74/Jtz2ZkyoDw5qkab2wgIKEre8qzb
/uHDdWniPO2opCPyn51CJY/75MBeYD9qfexs0PaBCa14La/o9qBFMoJtCrK5ndl3
xuAMErbOLxub/55wtd3/yOCDJYaIEnoF+bZBhsAmStENdxrhNY89yg+R+QGfW7hJ
glrugnjOUqrtx1m3fMUFSVCQ6PCl65KksiwE6M4p8+w5TiT+Jp5n9sou0aR5G8xY
3+GaFXmOhT5tlRdgcIHtphGpWjJ46A31vpQ1qiFiirojteRvKPZjbjXnnVA4VgT0
/YGWDVnZGdPDESxKgxFnMIYCE48Gsi4+XB02UIGmsyemhg8mK4Xe+ENINF9Si/Pt
CTUvnD2WL2Cw7XrzsYYmUUpL8qFRI+QuEUO9TYjn7xUZNOsmAn9jDRp2jrR/c0EG
sBUkJsEzNAeiTNGiufT0Xe6FgnBaWlSV7iG1Y+Kc0d0KcfiBYS3U0JjFLGFb+byG
OoNSNShY6+AE7P0iFHnZP32eHBvrLkUUN6xbOGmiKiUkoOKIAQ1iaAqecpifAE1s
wAQXs7stf8Y7/BSM1PkkmDcNL7ynmr58yI7yKxbVgTPU1h/zQtbKGYLRaFG5O8gO
SA6jVaopTnx4IJANthEfHxUU6GgjIrTqkdsk7ikveIj0J8jiEffe/e9/il0O2Aem
r1g1Kn+eMHowM8fScY/oYiOdcuO4Xqip91B7T0wgS3VEV6Is/WoPsEzPAXWN+Gvy
tI9HazAJM+KxoF9f5bYh4WwK5heU8ZV+hQIzyh2mIpol7t++ewAcMXRfBygf9NrJ
be8o3TNLNMx/eDxX84lIUIoL3eghe0/DA5NITyJwiHe9ROWj8Sl8bAqLcsSHentn
v4Dz8TKYZLLyInzYZQH+DkSIzpp01NQ4u/D48YyXEpmlmQ3AZXm5GppGsaH9CfUE
iRfLo5CIKVaImWXLWmCpx1/yLzSo41sLdZnba3L+rJUMZjZQbuv2I6IboKqfynA9
Wq+SEIzmgkMBNsns/73Pomy1NWpXZJrYbWfQJH8RKNmrG/xCC39KhYywJ1JPia3/
/z61kneyK+NULah19fAa5olfFUf4NecUlsTtOiEBLVnu51DDVi9oGCbSEpwoomoR
ZpkFUF1FfecHc9fkUHV7fx7B8cYQb18lNbJKSUhN8lv8bUfHaDc7ZsM/PBJtMOtR
ZODCNrEI4Hujh2Sw5Y8rl1mZ1vP65VCYUjILJ2TvLkvN8L+cP7Z99opOB2EHfV8A
1SNHq5Efx+ptd3WlpGZgPR8ty0ddX5Yi3Cn07IYHRWZOgMB/sWG83RlZ+11LqcLl
QwpK/ZnUVfVgN1By7cGCJb/7gMz/Ca+8j33hkiwRHnzYxEO4KccHl/6pI+6G+9Sk
YyahPvGy9fLspPJlqkH60zDU2nBi8moFExf+pWPSUbkvFp9x/hCZnEnLrnlAW/yH
KB/JCBUh8lWpBNS2seYK9aiJz0iGG07NDOzo4PoXWgbPGvs2qE8DDe51Xs6vTVKH
jNuVNc6xnScXQqko9DOUk+g4NFEq/iMTVHJ8kRLHhRwm/n2vowc/JcW+mkoo+M62
Mv8PbrxUzl0gYhGqjGbfScMJMY90gDSYzJFcLys3UDFtRPMrDcD4yvPD3JU++QG+
x4FuFDZVxwbUotxd/0zVYwcTp95K5R11b8pAa7X/h+o6MvozBR0oue6ESY7zaxhm
zu5Jud6VGNPVA2FOEMGMyvuMrP0TIzMvB/MELtxJU/+lAfhvGwyphzDhe+AwpG5N
0WBPF+1I/SONRtju7YtdWROPENK0D8gIJtKGk0UpI8BuwpiYU/Nv3TWxZOF1DnjJ
vctY+fcq+AhQuzt966jygkCQcq+CM8bH920A0B6Dih/acAO0yhgOgX4+VSBEbqTE
rHfJ4sGpnk+Jg40Kh8DTuPpSteQ70vubDDQfSmP9uQwUmJ8+UlKBekmcg1K7ZVZP
Gg0z9JxYq1Aw4jTKU8FSCfENmfoFI6D+UGl/hXKWPLNnIEllOizeyusSHL7Tv3m7
7vvRqkkp54cssqt9d/hgn6Sd8BqK2GQSix6yQ9VCaO2lWXnz06+JOsvtufdNp+Xk
jJXaYjkuc2Qk0Pd+6+55qwGY7Gny+W6tAHA1ZxqcKUQViCMpUbjS2kriccLtVg/b
h4O+pUZHVwu4W93kGpokkfCFSABWRoUaYsGS3/bvXBLPdn0TNcWJQskQfE6DaYNV
1Y18zKeijIxCqhcKdoQK6vDXjehfk2jW3PSuLwoVO3xI0Soi0rt7z/4ciVXH4kre
d352LG1Msjr9sumYn2LNiCl9Ia28mzAOBBbuLSU6xASYdt1y6Z8WUX7GhKluZNsS
MV74X3TN9GDcV1ReF0yfdR81O0fOzCeM8z0RmnLkN7z1E7d6A6wLlmSN/YVlUHtK
gOXW83/fmuVe7ARAJezGmtOhP1JPi8ziyseFJ6wZJsUzv5Vjt/M2PKnkV3/VWtFX
W5/kISE6dSCcgbPoN/fqRITq3FvjDPf41tDqkgoIVIhJdt4zuD7BbwSQyX2PRMno
/vpScuXXbBHehE3Opvf9XhfaeyUKU5uhiEV08XWVjbhSQuZ6sn//giiYCgIebBmY
onn166sOTWa8yjp1eoOwGjK8KRc/A1hf/on0NmGgZ6y1eXBsf1Q2KA5FxroTNtN+
GI2HBsMy2l74nrThwg4ua0l6OTzOhYCUikh85BLFjI1oiGLTOiUemNeqPG19nd/d
kVSGBhLUxtK/R0wLkakweshw/M1+pB2dfzwrU9pQqxOsYbf5mb5N4aGWNr2qPtyR
2nrWot2sLdn7SpFVCv1KCYyE4O4+cREvLp9QqTCqm57uoMsBNEX0hF72F82Gqe0A
PfTKCFFYUNGLhHH5+h+igSEPnfk0p45uOgWT4BNcoEx3eo5Ledw4d8g0lHwLKJAE
fJTspPhXgZJx61a3IqANdsW1m+QGoQVIQ55MwS90KhOskbE0TzKzOPIKqb2T9Ijc
npOqQJmLRygq4Uz+x/vPBla1aoXTkSnKEoyCVeTwu/J4h+CvT0DNE7BvlFJkAcRN
t371A3FL2o7Gh0GTN4phGsbwTacc6nTWqoNEnWICjAfMoOx74Mb0SCAkUvHev7J8
8Dzihgg9LIbZgDkKkGqHAfaPa+78eKCljc38uJTKhvJlT4aZWippwRzJhaRT2HGI
HM2N+eicTR0JGD7srkNRVRb3QOMSZPODYT+uG0OiU29OAVRapE/k80kjPPvG0v6G
Sda6jHnEf3kKZMK1MGFtl8IxG8wgXiXHh02Vz+p9pwbYsBSHMT+zrByFjou5SF/k
hYTQyaqdQfXzz6KbPUDVLD9U7eBbKMtZbR522FXkP8na2PeBAH8gfIwq0pl/acb7
+c1bthxYhi6s0B0Rc0XSERT/3cE7rzp0kyNGje1o3Fx1NMLd262UHAsrGi1mk7dJ
iZuxUbPVZTSg8AP5T0Py0xaHLPAkJrgypg7qiOEYXCLqqV2KHBbU95jwpBHdbk8b
N5aIjDRvlKOjCz2lQX2lq+RWVyEqVU5VFSrSuZFZIxTNCEBYJjVs+C85sBQPl+d0
0NpyOOrCMsfm3Kps7jYcopO/voZXGVgNReBQsD2gE51Gd8+Tt8iHkQJyTymF2cYY
Lh1djF7khNzhnq3798dqnXRIyvGKXNiXw9hkWCrKedO43gEKMIih8uQrgzp5LAOn
3zbLzp3ad1qLdK/nQQLXTeLyCP+t0YjIz7ezK6TNHZ5LNkQC0Euo0ns617+wM3Yd
I0/xJm0ZcAfjvtAOf34QoH0V3K1qSO9glfYLo8sGZK5/O0p/8oCv3CzZakBtliOd
hjCQH65mr2hgN5Nhj/BjcRGfkTGbV+IkXXEOQJzOEwqNUtnkqcaDhQ6RDyT9C/D9
YUeXfKw9OdaBvsjCk9/FZMc94X9MOIzDa01IS1Bax06KEPDeYmS6zuIadlX5wR/q
gTTLfvY9qQeY4aDqfcDCZ5EJSn7Qr20P77fTFCnAdAZgf2VHkMDkLVqAAN+7b6HR
kX1R8pc+56Y2otjmmhUgyywSwddjFzdKTw19utMrBGcdHISfZlhPsYS4DbyhEOqg
UJ6gtcgwj7epmPoFbPJX9uNjV1kVxs+sy9MkDHnWPr7FdirherSOtp660VmxUbDi
kkq/sk40MUZxzt/CpbskplPAycVbFXAidydWVZQ5l75OwlixLOlK9jHi3xNXy58z
zseBwesyIbHMIzBYsFtK7u15czbNGbEkJaOYjteuU4VCdBYJm/ArH1ZN8C0ZB6Jd
nxzfzBGpJD0eBDC8yztBEBtTMtPGqvHf0eLVVXtqSHvgvNopk0vgg/bqMT3tp5pE
/+/rWdbQkzmYVAKMpGY9DOJ4JmFQ8wrGD6xspoVVCGKhDjtBU/HcdkLr/E9x62bR
8ox4f0vd4GCLZG5Wt99YGt2z0qtZR8FA5X9roZsA+xFW7VUV62WE9ixQdbI4untz
RHQ/8e8u/dUxiki00Da1uZzS3yD8GqKJWayA7TLzJt39xBPfB4sHSl5daBydMJjW
BgldS8HCD1szcatVTAnWgf90i4Dz+D+WQdl44CUKGtk7EElm4SOeXJSkMCRCX12O
agvoJzk4izM4OEZIc5P0e39AZwXJ9Ji7HLfYLiGXzpNlvK2Oi5lk4aKtbxQ5mLnF
x9GxlJMyEowJeUp2eXeteoX0CZQ1arq2YUKra7GhTPl0ah1Uu5x1GBBrwMClH9SL
9lARHyx8iBzpf3IxaWcDTiolmWcfZNin+3yFr4tKqZV012bB/hntKZqaiV+K1xEB
yZDsbfW+FRcwoBT+AdBQXXP++9594oOZWM0H2Vtk+liMk3d6iHomVoex4j6Cxucf
ciJvIYgzGa/tknfL4XxF+vRoSskUQr3dLHZ0NNWK7luiwSHV4SGzYSvKqEUnsx7t
BCfW0kZpzyEAhk4KDjM0a0Id1LG22pTmyvg7VGFVtqyO0JXrctm6raGIOo3TrX+W
Qu1rQeYCciP3q7MJDPIGcRBdf5Jy4ZLGDmdxmScxTrN1MH18ZWknB1qLpacrCtUZ
TB1TwqGf+9yVA8nDQrh9VpORi1r2enW2VbIpms9lVnWu2ZaKakS+vuSjBxQEPcWp
sOXj3Z+DflxxA9yDnaQ4qEPRoT2vxmfHnDIlEUVHw8OoU6lce5VKq9aaWgD/6g8v
bfR2BNB8Y86gdcn0TscR1gQvDzgcVSb6x+v21lRomGltkye8PfGuQeLat4H9deaW
6gKSNK8oZ9bhoqUIBXVG987tykonH2gmHH7XeETFeQWSjFKuv6Snf2jE3A2Ue/3H
xJ8jmRgx7V8EvJZ3JOk3abKmg+Qp5IuXXkeH2Nmm0xRxuB2QnBz+bcHSPnG0qEYr
yjWiE4kb+/A4sG4apP0dd/zKy0jOUfUEtZuwLJN2zBYwb+xZjQg+H3fGDigQ5LFJ
H68EzjOoSBTAzf9IOglRNjD7IdzHA9sy9BmuMQTSxaGSPcIVI+8sYWe/XTpp1hBs
eZKCfH1ytF6BvEuH2PTOJ0pqZSnwTYIywCZ0uX43BIr9NteX5cIjUa59xahISqsJ
qUggd+fGhF/sxQIKbrXc+Qmy/8pVTV33jxFZ+2v/UeuFUE13xNngnxd+agt0YKOA
xR2aifzJxJ9BbTCG0Yhbpi57t8xxdqgwCX/h3SbszOjJ09cTXlgGkwiGblycM068
jWHbku9pTaZATk2pClpDL/2VTL9VJrke5/W2e2eG3dfA1eICBM2//J3xrrY0TiKl
qew7FCyXOeeTR0X3RvqWr1jzeNn6rdETYxf9sKGaYmJvKFnzfSQIz6jb5oxBjsSC
55/urpPUaBZOUtRJU9AK7uZc5S+k39kopM0p9Anuq467PHK9jQNNpL55ejLMshKW
7xTy2UBPgXrWJ8F+8hJ83Siuvxo3KLrbAZpUIaF40SvOIkvMMp6KH9792drQg647
iavptTdXHgNvlt5I9h9e3r5txLuTnyvN87xOuzz9sjR/B4zcuZu2q81slb+2Rm0E
U4pslZiYUdYgdZ98wYfp6ieiXlM35gBTI3Kcipx/V4AEdd3lAeZ3pIOgqsAz5Mv+
Im00Z8lSi/YszIMXEtH5hMlWnViEzP/0Fa34fFVAL2K32MI3BfWeRO4dgYbK6wwJ
EUkMGUnyYDGYJrdpRnVaEZ3u56s7PR9d8tMNPfTa+HWKnj3eJpcTUuGiXZkWx7bP
A6vAg9VbsW2H/jjTRw0EZ+XXrqe9gYJZ2c2l7IMCv8GBWW49pQrUd7LvIt7e0i+w
PbbECp8Eiz8ZkLMQDI2iKfkVRxW1OfjtFsy1kWRppUKHOIAnbjkfWKH0dnDBVQNe
OnPOyRX9WKz5/IfH9loZCmUVm/eYfEeenQ4drNwUFEt8I12pcmdCYwyeFS2Lfdni
RiW9nphhQ6xADXz7gg+W/USZFrPWavKdbaCJSCeiVwSBZwzyfa+/JER91Fojo3mt
`protect END_PROTECTED
