`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
681mJLWPxuwQN/Kze/8NqweEkZLOmz6UJ+dw1ERkiDg0GFWDFeVeuLRmxG3ULYDX
tnMpsOY6xKcEAdY99Mo/54qlDI97oRiLvL4E1W4Fxd6vtZhB5M7o/QfjjrfsRsKg
F2Lwbu526h9VQqPkleJoz2xZ5sZhJ2pnnqxVlt6iyPCQxZ/7S5cXvG810eSEti+Q
OkyfOnl4ivdpXfb2sEK0L61Uf8NRrPlgGHpoRDm2HxceG6e28VJrbow9wWLSgqe4
4kqk7BGY/b96JQOpzI0gQioLbwwqRi38LTD9/pn9Iku6uvXS+jRrepY/SfVx2UKB
p1VGLINp6QY6VuQXl7zUlR7+cnKjlHpTPxtKZ8xw42rDIdpxCeXZTn/q2ASX+vTJ
IjYpDlAEyGrQ5o7YSq0uxcfTGIp2vZuaeneAG539ro0pPPhpPRW2vKoCpauvCN3J
OhGuUBFXm/5Vrf1/eKSxOcZTBYz6Pxc+XEWGtmk8B9ZXIRsBANTaiiVQjubIWm+e
k0Bp79FVCPIjOFDsxCyZzJUVqGxyvkyxnOax+Qi0qcyyRFcE5fK2+3knUCsSop9I
ben3vTA7fFd2CtPR0xy/t2gOZd18cMtPgps5r4gxJjy5k76hxciEc1sB79q80D6s
XGTuRtj5Ayw3UOuIMggN/M22gUtprQlpNGiKxbOvfSgdDFJVPG+U8sqfKU4BI+kK
cOzyG6ieql0S5R0LCElQGksbKU1n+VwnQ2oWCbwpQAiiwyHopn3NlCMhJ23xS8nR
D2UER8YuiFkjLgHsqed1Z3Nlr1F4Ic/mS7+36Gy5+am08I9QSF4JlkxLN782z94i
0ASoBJDvsCkAl/UFBd/P62965km50iLs1dCWe3EOvJEnC9AzzXJ53UDuIpGRJ5yF
iCQDrFBy4ej818Tb3PzrrZdfO+LqqRCzxFxCTwyussA0vbxNZtlYdwbfhrK4VqOQ
qqLKMdhxof9xdr0RP/IUEZg/Z5NXmqqGIymz+J3TgcLQnIYIrB5LF8LJM5k8hBFt
TQ1hn55kAQX5ulhnSy1oAR+asg+bCl4p1mIPxkmy8JuWk3dcw9fz54bHIDa+J2eA
SiovLKn6pJ+41vkQzcxv81mH59hB75AHyZNC3hTCGFAcATaUVkBERzr0uemWoaIa
fGAarHv9vyxo89cddpX5TQ7Xyjho27ZdJfiemFxKGWCz6f+yP4Vj24W8bz+HUnDJ
+yKp/byYGSQ3S5bDX2nahJEeNFD8MiEPRKtF4hoSJWOj16tumZWJLY0V4ZCBrIeV
3RxvPGDTX+RmUS/w34cWUYB/cz5t3z49dXoxvB2t0VRcTUYSqMi+YlRJ5nTzSHxW
bnVvwW/zytyJhJvTe2CiaX+KHBeB+xof6nGzhrU9HED0fg7LT9b+PLU4hE7XCgJO
3rSmvzwl3V3fdy7xkAn0PGnXdyEFB310kB5G/2Ws8AXxYYR3v1n5MdaWhx3B7wK/
f9c0CljtXcYCWyFhTBJxLbcg92RO8iItKpifiOUsrSW5Z75gOpIPFr97+kki7wFB
0Z756VFxlEJDJ0QBqtVXCrFq9mLHgfLVTY+l+fw9z13rmqdmyZbSMQ1y35bSlBHq
+k7O8A8Og0Pq3b0+0E/89n8LlhebcE5R2PLJozIhNX6dc/NrNQF2jjOmbIcLAJUl
`protect END_PROTECTED
