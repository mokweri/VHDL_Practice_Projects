`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jwc3hWmX6KCFVUGeH/o5LXxAray+twKCkjvy+EDD175abkKhp9miyZAm9Cy42fh1
/ZZYAvkQ2/nF0eJLTYbAY2CAVE6Cck4UmKZzUh47vrpkfVwOgqRE1yg2Bc0SwyYu
ZH+VStVpWC2thWptPBrnzBPC9uwj4Kw56qzaJWi0S2pDJ1BOedTmnyWZd4V/KVlR
bGN7ZVzo5mKNPFXLPAUKLBWrjlNw6wq8SfsXqAgMGErC5WOHIS7HeMU1nsDLN4bU
gB3bUN29IaRep+DrH1f3DrMuomi/M87T6ir3J2L3haeI7l8/BpGpqXKHj5rR7LtO
dtTWMk/WqxfL4/IgnTK1L8smjVQAP7olGKyM5sdL7fqgfbo6GdeKBMErqQL8poZ4
qe0wIhH4Cd1OaebLgJkJiiW9o716Cll671lUfnir1xusLv9u+umOIPwxCHPEnDfc
WJpnO6z0HhZr2fUANod+YCkFG4vIJRczpta/Ok0iQl2V/Cl3GtrkS4Aq0k/woQ75
R1SILzI46eiKVEhPuF+QkIgP9ggz3Vm2K3FL91JHyKplUWGhZu/YRufY+0/WbUC2
L/o0WgQ9+QfnVj+mQnp0KLIsjnbkpn3Y34jN3fBMuBUaKPid47bhTDgz3qPwqASG
vibDM0MxhFYW3ySsItQ112gL0ZBGL40e6IaCmb4t8Kb6qc12izABuOCDwo0talBQ
n3pOm8ctBxI4GhJQd0/kWYVN8tiRFVGNy+/f8avbhWC6S8NurrdJ+09JtxNlU4bl
28YM/J/xZd48rFV/o1MzJ61hpnSp55MkJNMcqbFfV1hIoRTgNmGV6jUObYOisrOZ
EUKSUlHmMjG2qnwUlZHOK4ylm1gHihWgVQrX/Y/j2zmoufxY/OjKnuMkmtlWh8ii
WXXkoLVwG+uJ2UrlrFRrDf4VdzXDIc0z8Ewv//QIYMIZoVOyZXMzwYID7UA0vjpI
4/K9Nbkn5FxkLOtPtZxTx97p3UOypyGrOLZtmjVTEExAV289pWzDQzvjx72V86b7
60uWmTW44wvEyXFUmHiGITxfjPix+GvtkMUtHBAeQUIrV3rKx6elUBQBCfqc8Tbp
3ZYPM0Zn5q7bE2+OWjcoLKXrHANYr3gGSQZ0qSXx6xwP2nB7MG8iAJvfzSj/WhzJ
ki+rIgbgB2DaMeE8bPpoKiCvnhIGQvkbVDv/pytHtNyoEHlZZnAqgj2WakaZvL5u
BE5mMMYogZRcfzrquJdgcZjpU9mosmnb4qiSgrTg1jVkRqYLTPbvPsOvGS1oi/NI
BwKPcEN9OH0weg7oxYXb1ji3/bbooKuxnt5lOIVZf9kVYaBNG5tv7Vl7h8KfwPKY
FyGTtkH2/rtCXFYW9NPJ8g4lnP/5CFUVnkNG+XmIwraVVlxlUs4jYIk3Rx+SEIbe
Bqy3x5B3Bq75FHRAqorwyJsWKaEfD8HnT31SWM6PH7oVOYJzte4PP7nzvFa/8gXS
1FcRl0KFFvWCM1LK4+xuGftcFgsW1NZ1f8IKe/IVXNCeZghl0FdUKIErMYl96+/j
mcJlMf9jKAogQzblSV4vkicyfMxdeqzmRnv7XhL6LnGHtbXP79MVjRjW/2DBR7Yh
rq+Da3YD7Xpc3hWhfEf4lrYnWyINas8l4XCmBtXS01HYRjPwUuWnIotl9pElQ4JZ
dTUlxR1yGiM2QwL8+Mb8THDBKWjZhmgmv1M13h/FVnVZodZqORUtCq9j5Y4s3/S3
MTDQdINiPIcSCTnDkCCNtOdBaMyI7SQ7J6n4Eg6YhPxtrqCN57cT/fwI6Zt2SrQn
3lshcfCHRStGomhp7sC2569+VNktAh1i3UC/pftGyICBzavDzfhvDPdOnlWaAZLF
WHYA59yOrrUV43+5jNDauDxUxHsqsotKlhJIFOiSqURQxWwsqvKtYxDH4wYigtqa
f364jhr7mpfg4o+Axa7AuQ==
`protect END_PROTECTED
