`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3P2M7QkUpsCXmxN9EOyms3CE+pg7KAZ36rYKk1g2FK7HfKdrhwmt9suNvbxcFid
BoTEZj/H1TRN0/NUW0BOqNaLefB1rf1bSh6emnsnEOQ7Z4exqGFDOHEVKK263Fqn
c3xrZeobIQCUiOrjuq/D2MsLjHNHpB3r8qjCAwXH1/UDmncRNPcsaM0vD4BXmLhp
ciINd2ZmY7iWzD3KiZx0qhydH31d4wvrGlaxX6B0QjPgGGoVF9N4KcMS9e+wsWS+
hRPUIZpi+nNOYbyB0ryn+hvHqT7P2+0FEEuR1C+JHZ+TKuJkNJq7RdykeP8pfRNd
0ZIV6wpNceugamWSDMXbM7/1rOJjhTR1aRNtqdSIbsmGKYcZCkN+eiJVKgWIRGyL
9Ds4MUKk8O9UWq47IrDwVeVMQgGtsY4ozcpprYGT9O8aBA6f89eT5VBUPKZLRjL3
O03nBDCZpCxH7Nt0qBTTjBC3UpXK/C/DJ68omk9Wkk5t4P+U7ayTzP6Ojk+Ljl+m
GdU6o8sBv91sHUWe/HmwCtUF8m166I+I2TT2f36PUYue+DG7PMBQLv33BdW7KtKs
mKlK1mI6+gHcf21oZ7kQJmLiVcaFtKqIKclU1+DlSXlbfq5uAVHJN3HJ7h2m90BB
SKtByM+HjbpAnNYJR4xEHqH1Mt7u2qAg23Efq6wYicGLwm2+Pd1XRNhQxEzWTuU1
AeBPfwBPOhlfp9NGRxpUoHESpLEHqZxYt06cxM2ryaOj2dd9AGUn5Wp1WOliPnmy
9NcTT5q/UW3ZErFLjCCLTa6ccXpcCKlL+b+TCz3dxeXMG5GzPvWyOoOPlgzY3W/U
4MR0XzcwKyW5/pjKNUhFfYLDBQ/ZPvzHj1Omvwnds0u1rjCwEG4KVBpZ00DY3gnM
RCuozMpU6LSdh69Ijo0RauSLQId6VCum4FMiCcHc2gTU2KFXFo+NDPVaPT/j3j8t
9esJY+wBp6NaExueX6dbQPyO5QkwNB1pMZtJHczXwNwkGpFnEXE+Y2NlbDjjvuB7
ifRkmgHMrPSoV3v3smky0B79dieIb6wbv4yp2dx9Kt6HHER0F6vSHOHxBnu8jPrn
6at0qL/Ed9XssD4tMzw1cRB/YhxwJRTRya6NvuSDEW+el2ad83XFuAlJiFYLgTCv
cyLiIFpaZ4uG63slQCl9up4wynY5oloL7TfBpEoi7QGnS7ID3dPAaPrlgl2Hx5Du
RAwS/kOhBI+OI7FyZECjSMxoiQ9mweposI4FtMyMLHaQE04XTop5YA9La9GSlVjp
HDMNbC4YdWwA5gFfi9WYeyvTaZ7wQvJ2EUo042empy+mPFzisc4q4GeCbjD8VpoS
M+KdmSDpEJKtRCL6AGzPN0dPibUCEnKOOPtyVoGFgnFBHiXWGytgumQHCFHa9RuX
UsrVXcAQeGkKwaSW96jzwRxWYm+KCdES7xtrrE4T6PHEdhvXLvMHWYRSzVjO6tuT
XuOz9k1ZL1ZKQo3qxjHRB2rltGgvhV441LTlAaj9JKngcQlZhoOXIVb2pHIPNHLB
CCbbm1BJeo1yLmIHuZ+KSGYTu4WBbpa6MUReXU92WfLX+goj1YVxWnU77aq9c0Fg
A9aBv1fO03WFkp+BDQC09eljqZmpl0FFzqhbTgQiST6a3T7rWA/Ruyk6IKgYFXAQ
AzR+5kCubKnpeiw9JUiyXlQg4zUVi01a1ViHX6bXKUaE6A/tBdOTjdBy3VvuqBUw
W1SrpzCCkx3XpxuFI2ZtiMIc3AChH8okJiZb0kGbnuFlQF+sPNSoepmxeh9ZXaVi
F43e0wVgKS8ni3dRYvCIkZugI0e8LoqynQ4L0icuSCC4DfZGEhItyV2v7ElCIHY0
VUrA0wRl5Jp0HoB+hCqTlmbWR2Rlifm4JAMjDTpJPqP+V62D18QyC0hAd+jlMlHX
TuAis6KcN4a/Nxwljzb0Zp3RKOXkXXeW/aC5eZ3b+2nLDfdRfJrV5BvTqiYioK0w
awajJSvJzb/kb9oCsGuxAwSsCr5b1gxGN/IW0cf8zAyX7bwc+0C5S2V1ZoVZluBV
OK1cum7sgC/5RLnUIuTosk4M3n0ixXyF6NcwJCIUh0x+/bDFxJdBSJO+m5J6lU1G
7gcmyjk3Od6A+OVs9f89wYKUwSb0zhkNB95hGlFDBsxT0dSJhbaO35Uv7unwOjr/
tgs9XVQpjcFoXO8vjiuVeIM3451soTtFpfS1HF6yPSUxSbDfwb7sY2XBwS2kNB3Z
N9X/AC6HkUI0IjY/n7g56cIBqxfWZZSuInLnD2EDdI3MP+xY0jkqrVbJ8d3jFGfY
VmDwkLjTnnTMLc66UObUA2x7DTOBYgGZRl3pixqyUCxVgih7GQjbbE4hM89+Y64r
Tyg5DH+MbHPycBajQ4x+7j93E5V+DDr9iUBJHg06Kmbzm9NfQ6zLVqZqZA8XJBtT
Rg0Tj4iW4V5O3Xikk+rpSlBorZ51jgnR7+Icl2d+t6PZtHJmQiwMC1X5+EHXHSbG
qRO1W1w64SASvzJIBbPBQRgutOd+yZ9rfcujqmcyg6eYtcHty0ESNtZM3P6fBLMp
9/uyiUrSbmOsSI2lY3VhTT7UsC+IiYuQpNXM/hlCjfLOP9VmHgEZT9X4RVgaP0QF
s+clEfMYmRAoiCKHsXD6sO7uJA+mKTEI33kYu8XyQrmIAfiUCg6Ckii4Y+0dijti
LKjdslOrNwHW57fWW7xHv5StNH+d4tBcWooNbCU9NtqPSTwzdxnTZ+FmFiw9+ho8
5sK6EOzXmJG4x8L9zJUZj6x+6KMaz234DwXJEhXq839jJihLCuDk5Q2VMfgNwCC6
RPD2EAah6zcUDjTLz5aed+xUsZrUeNasCM9UqQ7tUiFg/Mg/JMIkFylEp2xWmvd8
VAfQY2RA78zbnTUhunjIEl+mE0CSI4+K/aAgcgrhZFK2mesu2/C0ic6UvhjbPtRy
ZO/rWTD4moMSo9khkLrPqnVC6GYOHcAK8xhDQINB3ToiQ/HSP50jVsWBuw+WIYFv
cpd0oyZCT+a8V7e/5e9C+qNSN59ZKdoSggMx9xsfv4W9TiAbxg4mlB4N13F6mZIO
mPbK1XUA6FAtwP+RgiT5qWcSVaP5C/lda+Olhs3+vniFq0cltza6alyWI3ZeQ1/p
2Xa56ZHUo4HiRaknUsIAUubf6XXGW6u2nd9siLxL5GV2KvhWA6Eaq0u7f1GqJmyN
4qNLeRbyAc1aJ1FFU+NWUe1didHsUOzXVLYxdI4axK7Ji3apBsp5pYFLhwtHninV
Z/7u7gLapTH/u5d8XVQ6XFYa7OVE2koM/un2rQTWqAxCfC8FjgVAE21Eu7I+L1kT
ZSJxXIIKXt3v1g82SACtmQUhlcx0xMya3BwyXYSR02kRIAntSlEI01ekzSP1wU9u
kTAg+SGc4oveCGeIIPg8661Hlzkk8tux2F+KbOIg5JxNwx06t8zGqXzzmdsft4KA
P7GoXCMup9iGGsBIpedHMQ==
`protect END_PROTECTED
