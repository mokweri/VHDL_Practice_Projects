`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GKezy8gcF1BJWRiG7xDoiUTTxNEfQi2/IfHNEqjCbM3t4Cru6rnpTUvsPs+Cs1F
+iLzq0K3i3FP1WB5V/p5k1rKr6hMUrg7NB9Qr7MOlbe53mmU98/XvKTcfM7Rqnxk
ijX598C/xMZzRo82DOGV69VJWEDQ4mxDCwB4MmpR1e2nJh59KlrhUgxpupOT8vkZ
xGYgZ1TuJcw9v9qaLa4PbgRYVKHwGagmXz5juaFFkPgmaEMjSTIQxbKfflWdtpsI
5S/lQQPgp+AKgJu+0lnVBNq6Z9Ngk3X8BqWuyPRH5yMWxH/bU59gY64dsMSyM8iO
GhNsex984kyu7jzCvTLN45H0XoWS+XAPuGnNnBQ7sovEINNWBqSxj6l0gXIp0qYA
5mjsMADpJNipYQQHlqKqiUkNj/cKRHofc349X3Ocp5XF4P0JGLjs72S1eYYcUbt6
QeC8EnSTK1ERbNaeBgOIeZYpq1VfXVFWUTg4mrxVqn46eKgR9KYHYVoEomrKX3G3
JxJQVjRVvyKBjnBOsEWFX+HEuqHVXUuAe2IAPIMEC1uTXMfU7vqTbqZzmFQAO56/
7h6uOBRaKdAgj8gF3C/EGT4aUw73MEc4VhrCGCiVQuqlRqONNQChnwtZkUyTGX3E
RLRJKq9Q+71fkGKgjJVkuFqjkvTvJ39weqAg4SSk0yISDyNh2mSC7NqReBBX/Ww5
WUs8WDmCM4rWoLI5fpi7bxBYDZNe0jNzQ6ryOWGJaWVo/DQXjms0fo8fYDSxgtvp
JhPqYJJpDi+pLNEPa0Nc5WyhTjdXxmbgz88D6GSFCMeTojucLALrvlEZg4KYQ3uO
e/v1OVpovckUmIRBpg6t/HesGiZlHVuY07K+3jrB6H28X3Ft7a9TzGV7vYJxfj2T
qgcii+mvZv4alKUoYYVbfpHnYYSLhS8ehpeHgnftZsTuJcNzFM6edW5UVqkyXjBM
stumh89wucfR68+wwgkBgr3v+D8GDjnDo/Heo3OfceMKCtlz6x3N9j6GdeJkADrs
Dh6pswkhvqikltsG3bBuci3FHw+JemwVV6rkxXdZ9OO6oG5AHN9NjwFkKKOgJ65l
ubnA5czHy7hwB6SGkApHXpAhtFbtWoLPt4uNswLDox0=
`protect END_PROTECTED
