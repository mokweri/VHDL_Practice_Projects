`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbB86hXF8Rm3M/THYeVjZuljEHwMkIMfGBBeKYtsqlKH7Cp6KVWDzbxKv2UMD85D
OJRgw8CxnYHsxFvelIoap+8kPpomC7CSizI8tpJp7ZsUn/85qYZamaOPv0fcu049
GVgci+XcWcvPrC5bbGSYNjcSk8KeFevN5ST1ipcdn9nbWj5GbJr5E9jQPFzSpyTX
u2Ts0tjgbuG4K97ve4LtZbobiwF7qUe1yIT1GJNPKkiDz9cy38o6QlFL9Zs+uhLW
WfOptnxtQTjmYLHSVHcaJmqti/xGWRaX1rHUXG1OFmCANRJh6Kyhr0wJaM1ZQ3My
2nzZPEezUWl4K3s9pzBOwf4cB1zHXJpzFhLZDmcamtB5oEHgXEb7O4EcNoPB9Rg3
FunOqvEEO7WOiXNcjcQhZV9fIQBmL1X+jVbnGZpLqK9p9uyc3FDIu13qvM7fxXw3
7uY4ZZULdYg9QJlS9UtJeJ2hUnJGyTDvaRwZIPFzHkE=
`protect END_PROTECTED
