`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvflPDhdRxH+gAvlKieBoTIWuRThwFlVlNQdRNAD9VxTJL85Cz/gHaRxxFSjzbTF
dAeojL2/BvuNAdNxeY/XRlhFj6Ha+U0TtbgtjEhej09aeeTTyP9g2nYlixY6AFHs
oJalgUd7d7v6G1DFUIS/a90YJz8yXoyoR9OGS728rG4oDocMbOZShLoN285Ci2ZH
1b7OjptG8mzovV5hYHNFqZHRtcr65aGuxlpcb1I4U6DUCPyH0C4o8Sv0SxAtx+Z3
yNXH+2zw2E8q4OorfMGaO78AUjN3bTzbqPRGdPqAj2q0c75+UEboDIPZC0VmyApj
12bkPRFDbMJfyFoxucdyRY0aM3IwHNaW1DyQXpW1wpkTI0S2xnY9zuOn6Sn4DZWH
TNZkxeLqxEKw+DE1nqhICibWLGgr86dXtiGek8PMXBqfsnLJVLp0+aBtQneX8fYJ
RbCs4NL3sx6qB3zWERZQi1d67LnTsjVIVB/Zp60TVhapMvPUseGJkb7j/ZxgCXBX
KRG2CdE4VCoGvXIZ7rPB+2E47/qpOPPen9OHMMKRudQPxkZbZG0lZ5IZfxIrds84
Qj9iEUPUOAS/yVhODrXLjryDt4U2yowk9W+dJ9o5/9z9fatbxeasg5sCbMFhf2jE
2e/GMtrL4+ttLnpqrFfU31qlwwemw/4qOcTq2o1fz1wdxBYKWFkA9fni8wbVME3j
IFvzUfmPO7tTTMrrYCZJRu36wJAexZELYUtDO/k/g5a84REp+5TLBotGee3WNVDV
E1K1yTUbtrqqsgtPwsKmWS+zhBScWr+U/Gzq/t+b8fePs24QxTMnq85b4iscF9mb
Yaeg8cMoESXkD37b0o0LmbX+FGx/ssEtLGbrwjjgsmr+U8uU1E4KmeEnV3hc3V+5
aS+dK/d50xyobOoCftMzwH1TE1iK8F8/cIUHp6/h/ikv0TVAe74D+OTUd2nmHEpo
M6zUPrcHYnuz2Hdfm3PRvescwURIA2lHVAzIA0UhfhunPfNqKqGHkGX5pxTa7/g2
a4zfn/InEnIFZw3I/QC+KVAco3cfAvSMF9gq0s9LgoKMhyOyBTC5qH//5v1olwXb
Qb4P/eyzC6D9V2vY0JO3nMM+adMQPIG/8kqShnf5FfiAJWezhnPCWIN2QN3dIH/J
MDpFvz45SskmDif/2WN3BXd7e0s1x879AWIRfcvkf3uVQhSlUfii4jwGWMjjTPGW
EsVaKlgF5sjcJWf+02ImOcnDblUBf3tJbVKM5aSFmlCbqTgQqRwqQqy5svQ9rFf0
dZXicy5LjC+tyLKjPsKCWi6bgFVWqiLAIKyewCeYB0Uql1LACCuu7uAkt7g3u5Q/
RZQh4HJFfHap1Rj9VgitpENhW3hxOkEeuoWYd4R4ahZQ36ZjDcMD9kwEk9GEgxGJ
4gw0E1oRccqR3ncbrR49O1dF+dxpNiaeTVHawrTK4Ga96tTOt+BZXeSvkB5dsdb9
4gC5Ut7ApASmsbEwFfGNr3RqX0R3HaPyQcm5Cf3iJ/zr91nxFDe9pqXrEGvCJ4A4
hSPptevWnAYCuTMOr7Ym12XjAHQ5qCLy3d8IADXsoflwmxEHgimF2XRJ2YNdegAe
GQQJGZnSlQXHeQGbS0hxWA76FVsf8xA30IHTUrqXCfMUo/Cw6+n2HQuOL5yWpaVD
xNC6x/IHyjnVgH3GyMwO1uw/yENayXhi96LC2zD5+WEKz1TuI6Cfer4pos3946I7
bLIsyf/UAQg86zZkD6z84gdBOqaHpYkafajdc3hBZEEFCwQhkWY7ZEd8rh7toqXC
gp5GlmGiaVDeLCg9FpMiaag4Dlt2WBRO7UwP8951T2Gm7RHzdZ6julzdU4Xea1Zy
PYVQvfxW7bmLi041VUrJsBIXU02SANSjwGiEw3/tkxctvs3bymHvumQ8WaDdvrHy
bTTpo8ySOUj8+L7zUFLVPicUnn+ozoliY3HpfOUtA/r7No+Qjt5yqNawupFECQX/
pryZNiEz5BfLI9+ALwZQ1RWcY9Ij18XoBkg1KM81Z/PvOQsEMXBBwFirwfen5cy7
URuA85YNqpScpCHF4fncxz94CjDnRTu+Xgq6wz06FwE+4rCHY0DvtYX/XQ1NW3cX
3mNIfrt+axjZ3fOtBvTYE+oyJ+5hPhSR1fVzN3khMDJZnJOzUtsPoO/01rEhl18k
8wj3inUHtu9A7EDl+FFOmeFvv9Q3HO3TJCkErI5Lw16Rl3KxIxxgoz17+sLvpL2S
637/z3UX/ktrUIkv3nO3B7/6rqCbThN0UPgju8Gf1+0POSq6+/q+4EVucW6RdsdE
x+yDiytG/aos1bfT1hEao9yVJ7KvF0zrERm1yOyZ/hR0U7q47P7PLhipVtM0xfPL
7XXESK5Mev6+ltGkKgxzyk1/MqZSRPDbvRhVzu2S/auNfYh/78HP+X4ip9vIWAG1
OC+gz5q8TWgpur6lSvm+RZahM68az5BgcxIdjsiKXKNt1hYyKTA7iUtmnNB14e7w
UD/ZEOWzC5TF/ob+6XZPirB6Vg0rSJn6XCIzjXoHqgVyC0XaNhPXuWQeGm4JDxke
igRAF26qGfgBEw/dcLXrODJyBIc9iEdALKp+EJhkAnZ6VmTnCopMAMaDiA3W+Ya8
oWWqpQ5ymI+aafElzx0hiA2M5f+NJBAJLlKH4rHRpY+hQagqOMf8SCpY6i4IwUqC
PN/AG+htUTbTouazJawc2ow0K+oL4CtLVNvmyPqyYOCIrO9IcQXa+C3E+xPoU4RK
g/aPeiAlR6de6Q6hRKhdyjtQBI2r5b/eJC8FrWN9xLDRBFZa1XFcAuScrIJv++5U
wOu90CPUYPsR9hlsYWdBbg/WK4scz4yggpSjAg+PGBM8n4T+R6qo7Pnqk2GcFw36
yWEC+rG7oH1fxz2e83y5WDdWf82rSB+4eB7d7EnfGLQ=
`protect END_PROTECTED
