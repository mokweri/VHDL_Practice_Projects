`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A9hOXAi7iH8iRcrJviMyGutkpsw01EAZbhfV5JLz2vOfI9OELdqpBbiY8F8E+NPH
M769EkANUuDipDvyQW1sN1dbPHlveYthilBeiwZrXSOsbFMRJDNlrHdcs0lrCgRu
WDgsqYV1k1pXueFfPOTPEJEuCH+1OKds84aV5smrZyqhlhFfETW1lnMK5yYRNwdB
HVlAA544Zki+zmlWszXWJKaa59QTz27o/XelEM4EX0R4WzaEcn2hcJZXtdW5D7f5
Rirvf7e+lz97bMESL+zCrKNJGEYIWuof5Usq32qwbOzqE8yo+eDDPsgI/F2Mqeyi
fPpmZ3K5ohADEg222MJsWN3Er96rOTqja6VtdXNJwNmqR99zufg9CpmfGEr7t3/T
enho0D5RncYQ+eCw5VKHwCuBlbEFknv2pCYCcFA6Pk3xF4i/GWDf29PzGSR7uxPi
bhZJobny7tFA3l49gs0RlMPLBhK4FUtFNOowL9nwm7Hi4NXFABeSbbtfrwcyx0Qq
WP/KmKP6AUYfPkpOq3VHBq9RiIuzUi1Qj3Hr6uIRL4apYlA0kyGQ5W09eJQ68Lxj
LyqdZ/nvDi1/BkhkiFuTQntiQ0BKNESpkOQTTDPv6IHT0oGqrJmca0sB0sjt71fF
mq/LorebSTTdKWC3Hp8xN552h8JS3Tnbyx8ZLtupvUdbLGqKeFLW7wXXTgiN9imh
WIKQ4i3YAUR/o0PmEVOuPwxuGsFYgl4PwEzH04O4qc39RoKAEX/aR3hBcWyUQoq4
jZlGBWYjuAzhLNR3DAyQQmWOVR1jNrVFJk3031HK3Fi2iSF2fl9qDqvO0wVdV1x3
FkddeUe4KrH3K0PM0yh6HLkZDlHjZApDzue5LQ4u68C33bZgnez62N0kLAB8XKSy
WX+MvkQvgKsq9yUvIGdIYda4ejvR0oYA1XDYsz8K5rkEWGfP98gcbkzUZaAGajOh
8YoV3/yiPYs8YO9TuZujNgmiM2ANpcP6cdU7F6okqPYX6IStfDBO24Qm7BegkpWG
7y265dVgL3jScRsDQ3ECH1gEzvJapHkvQhmzv3PcIH43ic1R9Au7P8tZJlIcHJ5e
6hn0dPasIGi6LvROgREVy36oKVB4UIIglzv0rbT88+ikL5O9Nuch2juEqqjetBRv
ynQH2/byGdTysvETXj+2+IxgKCpdMWceobJFzy0SDsz8q6vTK1ZEG+pzEnSslI/7
y95oz8A/D+Ob5gaZhuYqJjxv3ke5reXTefw/Eed5/98Q6nu4jddd7xWLxBpylY3B
Au+yUzqaZwZmZZpmg/XbndTE+tURdPTH2hPWOfXD/SfQFKdxglqAvBay5X2tThFw
wiOP6jPSywlmAhTOIgAjlTt7SbTPO1FvS5PyNEeZ5sl75hDvPG8V8GAN9MwTwBnj
CSSN3oQN01aJYSf42V/6UA8htn9TMI1f2C0KXDGX+gmTYpVkhH04yWrrB6LrUDI3
r+VmZg0F6JsGwa28dquQoxeNSfRycXWorv0q7V/VOtt/k/VE61v1HRRfUcau0AFB
EvltMZfJzyJEyS2QXyVKU/+VoM6CwPzgSwVGGSbLls9n5wwY2aGoiX9nfrjkSj5J
toRqNMuc66ORARzxiNt4hRkUGtMOry1N1yeVRvnVOaCz8h7oIvY2Bd5h+4rAUpwt
snc6f3Tp4b0FWZaAJTr3+75vWC3o0HIuRrVDp+wnHVMoe9pPJSgwuIHzRe3JzLbE
WKOEjlSaGEuAum0Lzlt02uS/6QeVD1KxP/kAYE4Jr5MH5DJnWi77LE7SzIs2+G5c
cuIL0BsjRg/vsNnESW//4n7rru9kMVcUIjUGlI8Fo0cdThheIEkj73kOh4xfGkrG
MN4ZPni1lHwLDOptyAazfM4l8u9qt2dAP48xbD9qoooK9lSdyhd6vzUE2uSnyllB
NqvWzYQZQFylcZQVSo6fE3SsNJIEl90lI6Qouh/MCXtDxZSYZSuu3bjo5DR/dFzn
SX4pozDMMrYkJNfj8Tz//eUasAy04mzgOSHAhNJo6QlAh3LtG6GPE1ClKhRbBohG
/lM7kWH3yDAhMtJAo+7Pf345gXfafA1qnbszjNrIUzoxfpquGaso09/lxIQWtDv3
/t3p5tAMoesukSdLskya4ZDzdZ+Zau/ELjeoORw9wdhvnVjXD9yku25lwWuqrDF0
HMMX7l8J+Et2as+YC46Lfjg4VH1q8aci9H31qijPl0k0XNGIlCggACCs3Pn8mT7c
XQYpbaZ9zPhn8u5GWpen0vTm/FGSbnpi0TLyu8vXCGIf5lAMrVMVZkOr923gypRC
sUavY04XHWMOwvQuJXJNaAGUB5RoGkSEyyH0OqNfKdS3WklEHdq67vfx94V2475F
mD5CfLdxFsk7hy3UYmIma9zanEpA0+2l7wxRq66LlumK+c38VlsH1sxDSzOS7cPs
4m4G+hXG1xYfkn58PXj838mLEQ7Qcgoph0hvKaCbql1OCXwoHQnj685VNPD74Ut/
CvgelHCZFdzzoCnplC7CUs6QbkLCp1iU+mSdvMX+pm4SUa7eUFSSn9BJpMc4NfzM
HZlx3uAbf05CbN3G08ZUnHJRrWuK64UVOpRuvPKKmthTWlBo0w5+CyBtgUYTTNBW
0l90lKrlb2J4HRbOECHC5zr7oO8FxE95GYPKKiXSpP6UclEcTYChDve/D0ZSxlTO
D12EW/MfbOrjtTwmQnF2atxiG85+2/eneKf6KSxgHgzY23l+aILQXQjW+qYP0UlO
tWXHuKVzdFIk2q9mlZq7IpcPifOGcIJCteRpHApHWI8hAuyVSYnYfIsPItX8/DZy
CklE/Bi7BZyQOUlNvvpx7AMvnejzn09XchRdIAbBpnoaEbuB3hfCcGuAbVBf1KZk
eicwaQ6iWVRKRAtKjoMQ4xFCyEZ1QhprHI/JfkVmieO9SG4NXNqmbwJs54zUbt6Q
kqWd7wnLGEYrFfXCLzcCh4b4G0vwntbA3jdFSby60bcCdwwjrjSNSpAPlxf1zgje
wtvLf5VmWmseK4JyXPbMkGZoSzehXD8pFtN9o/L0Ka5O1iwbQGj91WQekxZwxH8q
AUSqDyd7xKurxEvGPQ72a/MmEU6mIUSEADp0VLsmSL2rqBs3f4tzYNuoHBLnS/h7
JtbDcpg783xI3YWcRVhcPSyf2qzEJmQK/N++EOEBsXNgALgTtBuj1yLYz+qNGv8I
SbfJiQ8WHb4pvsguEZTeYcM8NNiQ5d+rvGaO9BZ7sPoxl2/jQ2NjU2I4oAALBOAY
85h/41EqSgUvaxp2HX2TKHOZ4tw5paF4qC/nnL0FK4v33wNK2qpIOm7YhS9YSCCs
5dLprYOynlFCaOKYGKr/8lbioFZBckTKyI3LlPrR4qb31FpSXjTow7eGOwW6m2Ij
5WuNJ97QHoGpJHCxDctYOZHZy32Ns9z18EBoffRLC1Vdz99Sp/TFkKLjdDXnOUwp
I0FgdGkoFsx6YHme4+Ls1VOS7N4/s+ywvhuaeKXn5Li9o+sZjMF1pSO42rsXLVgw
7/iKsXtdnxHD9OepE7gEIHI+q08nvU/9q7/2sFg0JzL/8al+U03A9+h1MqVFXEK0
JUa1yGPyHE+bGLQJ+LQhFOXXix+fFNi9gmS6d+u0x8IEmbD1YRcnh5sj6xhJVept
G1Amj52QHB1bWTnC0YqeAUqML0BcPQReSaI9WeDphS7DC7+mswsbkkRtspk7nSUM
Qfslc0mJQ0EtDOzfqhxc9ECl2lHANDnJGXn1guwrdxYT9hMfHEUFsACN6wXaFjX7
wQrY6+B8X0qZWHYjTRxMh0JR5RJq6wpkO1j5/zfiywEtIw50KtGAxHlugZH3alDm
UtlY5USQHhZ1oUHt+uBYIdd71hFUsJ//elwAQgQ8v84xx/dVS6kFhNXYELHulFV0
gpEk39s+uzsEVX56v5dmGkrgWNcIAv2qQqXEHiGLlE8nNOmZxe/FnWPvE/LhwCvm
N9MsAC90IDmV1q9SwM6nC5SnGOsNPIdlRDwBwYVvvKUAzrqeQOtn2sq/zBmKukde
Fg+Ppe1oIEVJ/cUkY3XIsezN3B5bHAe8CuFLjrhWEhk=
`protect END_PROTECTED
