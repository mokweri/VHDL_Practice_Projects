`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWZ2GUkeUiS8QrBGb95JoNirVJxbGxbmwXsUSaSDVpoOvKK+3iQ5Lw4hnhKVM5xn
rf+lnMPllnO9cIxyaQTEYpP/dTa0401Bexj+2xD+1a6qYpfGqFp4sCAvBlK63CsA
kWtbxS17tASTwqLtT44DHeFnuGyEqXxq2ZkR2WvtlGAwFnmN3TM57yAHH0oJyDN/
SB7e3dUscASGVAQRhhSC1q9gpmcAQvBi5e+CPAmBXBiKTv+sCMOGabIn0/sskA3n
YPUVghT1dBkeuvVWIRdyxuHPKiVLwADWi5EoLo7OzhvclLS7IXSGa5deT6byWPI5
B/RoTG8Z3uDQ6QxKwDb5aI9uBtBNVrkn/cIiCw48BBybrTXW36TonPEWNyIG4Y8h
JiwXO85RJB+xVZGSbKMpwChqlTQ9z6/8YsudSQNYZcwlvfGrd9OexTFL1xlQarG0
7qB3wMYbU22SBGlwv0lzC+3n0zz2k7ik8IDaEQTnDuEXFXIxFbxP8o/pa+3Twk5F
RGsc5kfn5t875EOowq9QfFUBS8a/36hTRqjvSzFuOBW/VcQhs9/mVmvdbk1aJq25
/990EKshjHgvTCnacarMCrmmsLlgSStWbnR8VOJnGtDH7/H0kXBsZCEY31gH8PfN
SvZvsd9HAhsjwupLWB4WrHX97UwWdI4PqYZxaepPXBQD/OxzQh4SIdjbUXXwdxea
4jrJy5rKvNGXicsbMFCa5h3nOaiclPbcsrRghEwZd7MWemvDAuzry9GRVpkzL8d8
9ny7Ncun6Np4WP/BwMZvSRLfCYgpxl25WHVG56JO8+jPzzRs5lpvbqc9ToftnFBh
pvQuw4MEpm7BlpTV/wuAZVFl0DS7GIB0muPHN3/1yAFPJx4/nlBtJ51OZSMVCDnu
+rLGM0D9vTmrWLqQXrjgE6569+h9PBeUnf5w+ey0ScdG1u5SiSwRLVGwefYjnDs1
iuaaZTz0ZyMoTh/Mrfu3AheL69w7/9T+XZkevovdQ1VFNS2V3rcxVfK57ZfS4luG
nkMQfZ/VZeyZcQErDmBq8O9EiVCiN6AQjYhFMuiLN9g6HAkKrkVRYx4WOkKJfjnX
eJDFzn4LNKXIvKbB+7p/pkV2MczNVmJNruBL7g7GeLJiy53UMnjVuBUIoACnrE4a
7IrtprXBFIKo8UcIOz5a6YMy9oMFI6UmXgDGPK2yc4XP9zs9Gx73Y66YVt+vMdlp
auoqhDZO+zSc0RzeN/AD7/z9eMRBWxUvuk+R2O5Z+32dcNJqaVNGC+AYG1Ey+1P8
It5smUko2B0gH2ZnSDS0XFUXcjp4ZVebrmvomk0eKf5tRm7TAz4UJOtGporeZKT4
i7esdLWyLR2Dm/i4ZAR5erCzwY9e+OMIHpctorZpqAM9ix363OOZpNY7VzS7Mtrx
dJKXOSvcMwH312ejHU0CXe9oiWGpAEpraxu6tS4kZ47h25UccZAxjzGi9URqaU+x
2SZnCLn+xtYTso27M3cGV3Nvphti3eAoaAG/lxn2xR7aQbVo1ypKYy3vyMlQw3Bc
5TSRkB7j8a3urZSxK6gTSQRHLVpW1tUUYTo2rV9pvripTAFWosjDNcGpK6mUPWn8
U7jqEmbXR86Ax6Bng573XZB0hVGavHZ3uWNtZGpL+L3h5SDZCNBYKz5mjrOKzabo
dqJzJj9DeLKlpNQP4/eR5ABkyk0MueC2MPND0q6TkE2PBLTVP2O3oRwJMGS0zIuq
woWdBCHtE8oOHJTf23hzyz7AycHYeGUnvKt7GFs37b+bK5tDiI3vf9E8W+LD60O/
NszDGwUC29WnQ7Wk3ACVKb4ToOBsyip+22u8FNyYnQR2dS5wemldfMob7oLvOUB4
hoc24G8hhlugXLZmaZ6nU/zDV1sd29G4fqjcuqnRU0wxqVh2HwFwUkDFVF9kBAo1
H6+RZbAKrX0EUI/Aj65q1ZbE7k2L2BgljHnWIF4DhAdCvi2mcj+F2U0bVaukzbCn
O7W0HC4VmjnRRrDah0BEI/KgqdQMYoM0iqfPiTC7igZwsr8eMUxdRfr4W2ybbwzi
iI5T9E6tEQbiWaBqzA6/j+OfJWa530cn1CIoo7AZvqEFrC/R/XSc3s5wAS4lAl5Z
rC2xa1GI6gzg5Lg9nSb5py6P9r2QF2RYUi06F90nOo5tGlP63Icsec0JOlZU0YOQ
WqQ/whDd8UWA24zZi5C0BNgaVG6pbJgBNH+U5J+1kRK4b6daY6/rrz61jNLJC0mN
gT8sSH/er7/NQC4OpFLY38mJBIZFOlyMzo1L18dOBukVOAxxSfn7ykajehNX1Nsw
Z2lssle5TKPZbKrYi9YUtj7u0CnFcFXdiYl6kdDq8x0xmICnslOYWEhSIOWENYbc
r1olTlQi3tiwgoknfmBVob/CawQCpn76Fea7jzgyKUCqJPWTHCQgb8jXMMEghtdq
sTJ2G/T2Y8OrSnku3pKctuuZ2iEVBllQF5PEAH5aawhDTsoBQeNUDLH8kHrS4eXS
SVrrUI8ArnV+iujkOOTXxjuwAwVyYtkG1qP4SjVvW84=
`protect END_PROTECTED
