`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Inq8H3FRLA3aGkFRga/Fy625VqbwY5WOrOY0DbMasqeB6B4/LmJuBUfVWb9VxA6
VZmM18A88nzYYmfjbG5gr2zLOkHLoH3homAob4Imw4Br68jgfbZIUDY0mbNRMbwO
2zDFbW/o1p0n5RgKRz7weWy89G9Hjk4FnIQLhq1p3yQ3zabFv39+uFYuSC91g4no
aDTDdFoi9AEofIYmk7/amIs4avLH+JDnaDb94B6lHtKnW+eQ86rLqQVaOwmiCcRt
8U+o4AUa2TUQkaoE97f/96RGlLaFzhUbnsZ5fjYM+x0bgG6InxkWgrmF014j+QLE
SbPIKDCJjAomYYqTjnFxq+oMFyFummrDyKkrSS2P1YcItSiz9/vb0aTAT59FWA7e
bqphj1I3MbZ1ej8eJgHNgSIwYezWP2E24qnMXbnlzTSff8cd50bUckbzCEy9/nvF
JOg7TECKX4Yrf/OmxFXf7eLnaxK9bDKeM51Zd7UWu+oNb43sjt0aQHc7kSZSHODJ
lvR2EqgbXqMfLgy8GwtKG3XwBBUOvjO3ACqljm/wz0rXZMCl7XqNLamprDAXMpAa
Ho+GhaY9d9DQbbY2YDXHcm4fK0yHuX6n3L3JRUN2cfB4JLVlocdchmb/dPOdePeu
eGfU/Pp47vcZBpvDRFYC1psV0PBLc3vJDlp9TSESIBt8GtHcVgARqWHnw9a5BY9T
ri32hvA/PZTdWSuuBcYrJ40ZtE1AUa9K1TCw0ypbT33mZ5HuentZRP/uSRxDgCFJ
Dmq3rR0Jms86J6YmNk3XqrvRPvNF6QtyMti08UbzwzmN+zp2ieD98ef3USWxW0mA
dex+xIGf0qQKLsyKH/q17biDtiDke9afvL51dWxE8XYBc2DCqDS07eZws9T3r9O8
7j/Pas9DiogyXCPkOMwG5fOwB1/xyN1o8FiEBdbp9y7tkpZpEW0T1blf1j8Smcr3
FGdoK5CTU+OyggcZV6m5K8VnLrMzrgps7gxlTOZ+U5unRfR2fBjK55aa03NAJ4FX
XiSj/n84EW7SnbGii1pzyzhMV3yrxj9k3CAaSDAyiRs5U9/kHIYAmdIzYXi5Mwut
5IkOm4rt3cH+ME+AWMLIAnLCC3/8GH37KcqSYYCKYy8bNPyX2Vh3tIzlbHddXvmJ
6fl8CpfblRCgtCpV2kALObmHE2UzR36XA1Cnv7sVKRBZnnucYf9roJmmHmeQ/zwk
YJmpgkk5EsrtAbGOD1nH4B9Gvc/sQD8UO2+BVCWanXqfmfZ2Etc+V7/jdKQBu2wn
oTFEa77nb9HE+thq+9PtTt67jLhC5m054dS6rGqLkCs03tcnrXiKhn+6B2ZOAYV2
HG7aJErRWRLjImQPBLLNQ4NPHaBczhOUmfc/E1i7NwGBGvQjUK/TEGh3QUfv57K2
LBG32A/Wl3kFHsfDfpiQwq38n2WxQeCvzwg7vWyxlvF3S2MrSxaQ+7GOBNQYHeAK
LDZx6/gK2W9DSX7TwFgNFKXcfZ6tdURK448BAGDkUKyj6tnLwfxMcex+iVOjuWuo
ZQiWyCOv6JMjcQorRChfoHkpWznO0mkS8H1GWkiRA2PBALLfGPduNM2MWCAAUveQ
1ZK6AxvUY+HiHCm2MqbKQ7npvP4UZGiylEZkf2lpXFpcwrxgKGug6sJgffI76VGB
5q9BHK2WCyga1odK/N7xcQ/tQRdRmdzcWdkzdjM8XZeLTBhEoOOw7ibKHoXAo+Ut
C9cGlcO6mtNM/2hIfduYSQ/PyspXmqhJdlHNPhcXg97yWMjkzXuQrPZiNujNZr7X
eL9ishM9DDZHIguOXzwFYl40n/Tm+k233e03Py7S239lYhbYgZnqqYEW4XfO41BY
Omu/+t9YYqtHyUkyVDUYbQve0tkr4Ss9XoKVIVboVM+PbsPEijCABZWCTYqOhwRt
ubQRKiCmjX0qMJ7fqgFi8nE5UrIIiZIW5ffIuo4XzKo3XmtyQmX5myHPT8qwZW0S
NSLd+lKrFDYcxhaUQ/t1MAwOkftGTHH1DOBXIysf0a9mrk5AONUbVRc4IRhWcuuo
OPuAHLYQk2qFPvbwx46/U5vjjyG5HOo4DIfxyfbuzs+V44k8O8edQi8f++mRtsUz
qZbAdxsAwFY4a/Vggq921evjBrpgJlHJXcCA62Iyb94I9eA5pcP9R0oJbzNyXtHI
KvPA0EYURxHPpOxNO5YOtprRbH7hhfIa34UConEbORdza4OjWSDlzfC90jwBVty7
O8qHF7iBjsbWN0Bsdp7gGB2EUeck4PFbfIE4edDnA7Z7eztMN+mn1C/jGcra1o6a
pjPJtt3QrctjPshcPfEQ7PxtE2VMxtxF1QJX57wdnqR3j5lJ3s4ICBrMff9t5kzi
6Ko4YRPJncygJ54UYhWZyMK+ld18Td4zAEqju7dI/759dJ7gC6FqYfss8ZBk2UnE
Em+e03tXOZEwg7uaHloICpDJ7173XvI2N/8Jf1Ss/Yo4cl1NDPOKZ5NdejFTmj1g
rJlwIckiJx4b2Ia7s3+Jq+ix+rqfzm+n9WuQC5bBPeUUEWk9+bKRDQKhQ33WmHlq
H30Z2Os3CHJp1F49SxiO5EpIP2NQVZ6Srbf2KjKKcmGrWB7+wbqHF4dFL+5zbqt8
SUGh2p9CGpM+rH0/kEL9Aw==
`protect END_PROTECTED
