`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+mImteBn9C5FcRFsILhkTZ+sanV+9TX0YO1PpBcKuMrFbtk8CEE5YEtrKqi80Bj
JH6vUnmFdm06l8ubW+m1RbP+0JYDzYskPjca/FSYr/jOUyUvdS4MjXgdlopPOZM8
GadfaYH586Kj6rlEGzrTuiPCHsbJnMh4Gyd3/u8tXzsfBfSQhwyqguFL1F1dNF9c
dUpeFD8BLhwzZO2oMyu7v6Vg5oVvWcXMsOWADIy2HhFsVCT3YHeRRd9SeR3asrrM
PjW6ASqSf65fUJFV/V9TeFMMIXUD9Cve0+Bh1zTCeCYJQOd03NLbcRekeBmfIaOP
qDQq7ILd2WUdfMDRyHz+DFLfAAoTXa0WxJc0R03wD0xGyd5h/g5aljdyv1q4GSmP
2iVHJpGLCCDVNDllGvg2pLrq6zo+s+ZHzCmWuQgqVLsr9QQnnatcyI8rCiuQa7dG
huDeSVsjFYRzo6yf8q3ubKbPan0YvBHGMjoSQqclzvZnO8Ssqb/NFL9EdGsXi1IY
zoyzFFfwsZH2FA0Ply8389JKZLdttMhvcM4VH8sHzZ5xIUoxxINDaoRWDSQgNn1S
GNzRVQQE0N5iiYCtkIPsmWVYv+VGPgmINJL9bkjq+vRNkUvv+FO/dtexNzUSD3Hz
lMIbZuHNXvgL/+yAxe5VGWceo1DhpV1vZjLjCW52dngUd8FMmeOPe98x9FhEb/fo
zy5pa77xgTGLswLqH+f9T9HRRyEH75ln/tjuQBcmc1YxbJXc3AGJ8EPv4KCyKGWi
O/sNdwzAoe1I4XB2kkTNovq8U1bz6ekfqau3PiOZ+QzbC/xCx0Pz+DVgfSiu+OnB
A1Nb8bysLiItBUWgW/nxMjfIa8e1vwQFR+1ajgAlbzM4fhUyIHojnWz6dV+77QwO
DwC1vo6oMLV4UN89HaIQMdBtdWZop4W76VgPnqy99pdYvO8cJgu6JXqmDHf6WaJg
4tFEpWgNviX0xcTA3R2PFyX85GTa8V23WQ67OkR6YNpnuBHFI6APamAwGIk/ePVq
0OzY5VdrlkBNdGm7laDBCgdAwBRO43zlvm8Hn0jLJnEM4cj/yvwRKnjOJgFNSzG4
AkWdU9FbQUkhLX1DzNVVZYN1T8mBpZb37G71EUmBvn0N5ctP2RZGCHewU8I7Tpfl
JfXDy805FtOh0d97NHqyfPtcwxI18bSElsWJo2QwzOQPLycuJvmJ6+GE2Pm4ZGzS
+xB7ZQpUpE1+6b0JNXEC9tQSb404yP+8UTAAYdxmUi0=
`protect END_PROTECTED
