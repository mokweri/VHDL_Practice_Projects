`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NY6S6OmCwuupTYEqSYUkB5WMwQ7qhoDcyEoH8I+pq5wvKgmhhacbQyDBl1TFXWc4
QgEs2/6skgdhWaf0dVTCZ8u1tF7ukwmQZxmFvb53ISA4amfXEjeCKHNNi0ZFbrW+
gPBeUlp+PBIF/sX85e4Z7PBynkPP9fN+pqKJ3fw0cHlB1A8cy+wMOrt1peDfmWuq
F28NSC2dxryTox/HUyXJqUZ2oKywObpr9GuvYn4zcBYUjBTbYNV9frbJV23376yP
VqJ0r1/B0Izm+1V0Wx7sOHpo0BJOFb3CM50ajXQnv+9YfiH1GqlOTcZsgrDmXGB2
qpVhHChTAnZ5ExQ/asOhPSHz2DdJ4UQ96yPCcjUnU+WO1zx3D170ObPa22514v5l
R8yXkOrdmm/YdNKEY3apcgohXlkEAw2EjFPDZbcCXZdAO/7kJeG4JM+gEKDD9ftv
HEVrDZh6DoNiF3ApAIbCWLwI6wkdujG4PNvlrp7ghaVqsDh9zpmIk/f90dsJnxMr
qMAwACJiLHywgO2QHm6BGTlphqxYULY5pjjMggkw6Nqf6Waad2KPPIlUDB6wz2q+
+xZIe5p+b8d/xMqUjsy5xxvRfnAqBItyXgE16jXHOHB/5peRBEcElbHbYjj4p5Xi
0kUTvGY8SYeXzivkhxQEWb1C5hCpNJrFfrNTx33QgACIxUFLe6z8NiPk3S4Dbk3x
e5dnMiTpjRwBQ2Xrt/Ou/vC0Vaqj7AXI2w0ON8E6d2M4UhDvE1pVRR6sjvFtRlT7
5WAwA3ml+YuIBZGMMLYnF+ku+Mok3Uor++l+uNDrR3kkxxAIITnzvMxYoY3Stee/
xay6RVkNjYa3icp9OWHsMyCCuycjSh3Tbjt5MVR6ZbfhY4me4zao2fqqeNUrnehR
lq8v1wKvQqhIZkPi/eFXpm6qYSvmU51d9kd8mE6TAfO/VFgqybf7iq2w3pl87WOV
RPaNdov0/sJDdw9cJ0gpPIwWEMd+TPTab94Fn/YXSmrNZd77ZxOK75yMha0AXseR
IX+ZiaKleG+keaWKx8wzFI5chJNGG4YBhylw+71NnTi+5xsoE75DyekV8kXDyh4q
j/Mm7tCX/ufWEtV0cTHYcrlgRSWpCpbhUG271Z7p7s683r+IeXfTDF2uyiru9L0W
UYsb8w15NE5kkyZ7ESUHzGMLRiIzfpK9eLg6ZfkHKpDKeDQ6KtnZg5ZDxednfyl1
y1YPt0pOwSmvwqSr9T+rtsjiS/1Q9mkG5mHFCecPkx7wJArm3PLcBkSp8rAuMl2h
dHH34eZsV7005vAFnuwItFzJWMk4JXD2igjuZz0hgGPXnEMzJFv6NeTTnFDIVWKe
r+vFyVPgZLzEfavavSTKrjTxO6/sjcuEwrMw+s1PGBc2IKtDnmbmehGPD85f16vb
NGP//WdhSS0a9WA5lvNgK/EGGJhEVDnPMNWA/xpO89/O8PfCBF2FYl0X1YVdDtDb
FifHTQb5FX2guZK/I4qVJmJTxYKpgNMa+iik57auJhR6uiKOOSKQngYCV3ekK7p7
lR2ANy/hJqdYj3yIiLFWFz+sqM7ibNfOyy0+1OOQOqzsH+B+c/3VixoGN2mBGXpK
SH3GedLQz0cmJZBEQucUzMnnb3NoRq+uzpSx6rThrsO1268o9RKv5nvNIv6LazCI
lIiUBQPx3C4ZAs0Mi/DL9G6PP6f19hB27eCJ22Mb2aKmhReC+T9MhZcH2sZd0Py1
OxQkby0rCPl9AMwuLagR6+sR9uvTmgX6ZXQvQq/NXtORQqiMD+rhrtnGh3UEHCB+
5Qha8zS3bsCIwMiBwADkSg5+liPA6UKWgM6DaEN5WqglIk2Tan8TiT1KVFjL6SoG
Ti8k76wNZKTKZZpUM9OJScFqe8gnPkeqE7fRJkLEWWb4j/pkSeXa9cR6QSVSM+9O
BW/XO+MjFJb5xrkTA1aFTFVSU4u7+MyIj1PZLVkfQLb5xR+ykAQOz6MWCHHveIgG
QdULDLABnc9ZjMMdv0+trXU6Np8vrLBLw5i56bgVXCoGz9tE5pwVUZUc5LAtlsbo
t/e3+kY7eyuHE1MqF+xN7i5/BFXpe6pM95dyiV9Qr+mF0PL7sIa19R501mTzGPla
KAhxREap/r/SMw48IERYvPwN+gbK9jbSs4NdTuxDl4d1SWeWo1q0Q5zEyocF7/4b
Rio1FKAfSXMA20NdabPqkrN4+C0HxTmcZlhcoErPhgHpOT3yYu9SseaYExkmHnSU
ZyLWUwc2GaBvkaMHnnD1tqDAaeSTDMWMHExojx9ZTCRa8q7/1bwVMk1SPpNIQ6br
cDmJQ1cDZL0FQrcfm593tss8Y2MOV3v6yM+g3Jh50x+L8lmN35oBhjJAW/NIG6xb
BxuG1TV6nI3WTeNs3oXu1hacLC2erHnDD6qyKNmPnT70f/uJ2IgsikBUm2cxEUAe
lBdzf9aVnH3oMjoyxDDOvUunaNie3rg+r9MUMuiHBNIPzap0zU0IJ2DYf2O0Pv2c
8ZaEjIM+uwJskm2v7EqVSMUGv//YaXtYAVS8y58e5LvZjGHvujCttxWl/OEVR0LQ
s7qULicjKvuGzgJXSnEvLVW8sjEB3OJOMaxDcCVv0byr8c0taB2LxBVamuSK6sQm
Epg7cyuldjEnJqZhTFhHYr/EmINGWZwl16iHayFettxJt3Sd8YOeMv8fhuIx1Qxm
vFJV7aKvVIsaqb+rePoAL9WSSG9tCoYoLMGdjbS5oGabMFvHbqtFiut133Tn0EvF
WuxJ0t2FSB8vG+XOuLMxzQ5gReo0THWdinbTJjKEaPLc04nEws1kZP0qhYqg+Lls
xlDJUMiHZWU7JNCoZqqtvt+iyI4GoSrJj1rO+3QUUewhik6/Q24wNSAYsOGqlHyE
F8YqezB2K/WKI+7wwG29TGjYCb0enT0ifoMOh5+HIUwk1JICeB/wgAXWkvh+/ysS
PcmoXxv2j8e4rNO7hRTdj+IklEGkkQENMrWtaRLU2ZVkotsOe6gZesQkYOA6LZqT
+0ggPI3jOiWTfAFd9hurAX8ZTqwiXb5GWjMsVQyLV8J4Rb9Daer/Ugi3QdUuY7TB
3zyrnSXMeEQ9zK3X88Ex0yuuN7pQKcy8sjZ7cw/g7VPO99NiBzFUnVaFjYhgNDUi
YmZlRQCB7FOHoEKrmAlcqXd23lmZOYUv68lpxLiYnWSymc5DFkn2O3+RlRGu3oKX
QYui1nPME6UtKiMRh1y/KV7lvHGHTSTxVzCnA6UpGIQ3A/JArVRnjfdEX6k64uOh
Hc89K+POBvkNGuOwXxG1CgySnPDgQKoqr2uwvUUlfOr7UWLFPvJC1tSspoRmmcwF
7uIXCgIZ1Z0bDbcBJYpVhqgU3Eu05diJSRRK48rvTxjLXUXOhpa68O49UR0rvPIF
zElWZa/qVGZ+Ft8up1gP6sVLgge/JsyDg/PKR1byEe6wLpdivnoqIiNDNciSq7IR
HQqdz/CPsbFJNkQAgRhKZ4mMeltkk5Vbcci+DuFELFXicDtfcOOu0BZeEbu2r4OJ
wEThTnbr53FfAVkJ9KqUexBKDb7vlBouc8gjaICWRcncPX/egw9YY1Ppb2fzWX72
kdbAOBp6bHeTBW8mWuJ9LEkGMCRNgBJJjy7GpXlLmLg5djn0nGE3aI0c1OH6fsRh
/ihn0XzNoyPlFu3SWaCorhqk4ytGePwOmbyADRsNtGhwfpqNY0rBruqR+4Q5T1Y5
6+R4pFYFzCzNoUe1PwZvrsk7tQRpLB/ywDYx7cEu2m0KRfAMKqJASKeeFsUCy43X
nbj4dQr8jX2uR3E15AgQM7yOQSNc/sFEfI2cBtgz/5MZgXk9xNgH2axUv4Rp/SYk
MaN+I3RaIm7603CjDZ3rRd6y1jlHpGYuSco5ss0b5hbpbdhm2aZ4jxCVz0lL9tqG
czlCykCLGuGRRqEHpnoYYHAzHUXc3dJAsx0abLgWpJIQqX1K1dgDJd7OG8OBTD6E
cXmb6Uqio9PZkPhYWXCtAr4i7ksoZgpVIpuVsJKuigO8I/nuu1OFhzzeWS9QjPwV
8OAdXtWlkAcGjvA3C6FGfqElU9swgokRV+FYRaHpFLWjO6vqy93aUhcDH/mOMg+S
wLeImpG/1jGHx0We+LzBw8tFYMRHCpLe74e0wwCxOhPztA09Z/Otyo8v3Rgp42Dn
UOHGh0snLKygd/k0HLeCV0TFLn7eZ1StWUB7ruH7s+HUpetvT6XT7T7RoegIx9Op
JVJ1OiqeXua5kkEtVa2l8pecpyDpbqF9ep9xLBihWutyDh96H3V7f3RcCDVo67pR
6RPGh495hFkvJphukj0k2TBwfp05KwmQLE7aKw9RnshO5qmIZ/n/gHzJbHcJIPo7
b34zS8Z5cf01PW9eybcljunkXxj32mBJjE7bZgq/n3kz+y6iKrUOI0r4/GcHpEos
ShYeamBeTTwMwgH+rvXsyJrUNSrJDAvhq50+Jt93sSUBK+Q+edllWxnwVW1eW6OR
RcjZu71HB05dFU/Boy5/7YWq7sDkSgZs5KroBb4bcfvMJcGqVzthVoEMCZhBocjX
y1PMgn9O7PSvYruZAR+8hQ==
`protect END_PROTECTED
