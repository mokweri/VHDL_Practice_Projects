`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQ+QqqIDacnw6UVYYf7zbX3XYloczNiX364HpE5oYtmnpCcYOAu1I2tlIGbzM7Xk
TX9wrEBqB6kaB5FiSGTsCTt8v9o/ytlbIXK4t8xw3TLYveo+QBpck+zGOvbJqtWe
c+1ePHLk8o2DdQVms+wOiTe/oT+Ku7t1s/8hMPY0yGP/s3ay4jNrW6eZ+Z/WgXb7
ik52X+k745jFVozwOvNj/aY5d0FeHwI0g5xrmITMYVX2/VZ6Degz4Zn5qZa+bJdI
MG332PYqGRHOMjCrFIbWEjb3mu12IV3nWTbCwuxI+jrJi4LeYJcGhOSKHVlPxT8g
fL+nsb/5e2+rQfCCmRfuD428J8SLHw6R4Ook3PBxwMxhINt0tZJ1qDbvMKN03DO3
lx6+u/rrhUc0ZSnb9FLcr5SGvz2deX5w4s84m8UNO6sis8vL9NSvDozIlrs0SXe2
DATunnx3brp4/CdfEELGcit9dFDQv5gggPn9QmJNv/k=
`protect END_PROTECTED
