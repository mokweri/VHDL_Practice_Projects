`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWEGa0eeIxROUK7X1Y3cMIGkD1eNBdHe0l61FcVBMO0Utu0Zs5RJN//8GVM4Slj+
KOJPEyZCYFjCkYwDPtzqO4nUKHbcq0c59F+Soh+Sq0yAFdV9qGB/I+J0gY71P1GA
cQ0FmDoFmTgBR2WwhjTak/x0pAdxdiy+g+eFOo+JXd/BSigTa/vs+6ZQUfwUqabE
y1YxrR39tVfaZ5la6xfE1hfBi0z3O7ir3kOPKvqstt7sgwQ1MM7X11ydmWxFxPMA
CNapYTcRAjOJWUQxYU4upw==
`protect END_PROTECTED
