`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9HlJ58Da1fBAaTcGC8O5Af8CQX0xUgLBHmaSDn5mP0f91C+PHQ65kSjTiHP34ZL
VcTJ0xeJPuStRjFXN9txZTJEh6LBCfNUcSrfcjDwY9KOp40mp1CfqFtzGqRhDsXD
WL2cTIxJxvfot/nxyHzqyYZoMxP4KXEyHU14mqFOLoiLJAOIGZRkJAKjR9XqItJ1
GneeLWc0RMQsi+Xn8vtsd61XemGb4P/zrr0ihdVXyyoRYowOs9IrYxrbBc2MTvjS
dQPhv/ECE5oLZwpsr1ABiIK7wKD5GyXLo3BABPlv9nwjDttzqX+XEMXn6rZcubQd
vCEpzYhpH1/eLl0PyiOig8EcD8TOziOLWYTTL7OK0Ix/aJB+thVJcwZW3X0qkWDU
9wQvwfB6QuuW7T0fRmNXgwdvmJfoHkgWNooDLiZKhO4XzW0/TVcVZt65TlsE6Sg/
XgXitgjiwGRP0hqqbkKD1d+dvmDGQwY9k28el6QBNtLm80CAcCK+0nEdLW5WwyX5
dbekKK8LMHjkiDL8jtdsk7aO8Z7Z0jP/M00IGvXivGfSv59hz8uGauxT1INYpyMk
NYP5/uiDEcjdP2KV5veNXqFcO2B2+n61/B6RAR9N7hyXTVz8+Mn4NMQiOuwQiJil
vdWXf66ZN1isIhb9Ctd4GjuJ7SQdIAekeo8MCyNFt5k0rLEtqvcPISCOygX324XS
rtmhKWTpr13/lkbNYifGqqy/UofflCgpyXct6cx7zdX3PEjMawFE8UdSUQOI6nn3
vM5gpONIYrAynAToEMjYMT63xRhRnVv/dtnab93TMRek4GMkU6ai18Qnqb060Eh3
ZAV5N8FXku7evQJFuOqXN7KVpssQk48RtIf3cI3glIQB+tgI/9bDyc7gPtA9g13d
egRM2jiVg1hicxrYxWRmqNQg+PlIWgBkHyokTxwvga40+MdkeFAiPI9vyksPaII7
eVpv6hDQHXV6SsvPfXs/2qQhO7p8GX+2zcH7k3dije/zfgCyOio1cRIB+HEOBIfw
3QMXmI5NAX/dQchZTlCtlgGTp2dt1wmC5K1LYuaVxht0ZKwO/2dnifvENGNcgoNl
4ZoIISxS5XEAuSHmeFhMBsqBgG2qCE3uRlvZz1MJQxAMhm8c33UITzAwDx8/8KHs
38VYU3vsdUxhX2wrhKijjKJ0kNooWNBj3qZXqlkvBrWwMbOP5bL7mRtMrhL1zZxT
d+PK1JV4khRtx9OL6o4A1TVD2xI81bu4ccH5tGl/ZRePCQ7N11qxLLFIFcH+/YOb
kppsA2W4VhWcD8XQhETOrf0VdnxWkbSuOEKs/yYztdEVfevAB/oCwIzSpRhjSGaU
Hv33Jb4B4W4PxHLvSc0YuzFmn4yRb1XxmKEdL3iEqv0k38f4Zvb+8MnQg/1gy9Bm
oVP/2Cs35fyr2rDpk5uqiFqMeLhE1NUZ+1z/rgpnR9IvFdXxoLna6YCP1P3Epi45
T4s8c03eoYLzKQUWrk0PJqkrHiBAg6+YeTga2tPkdCU6AwlUTguG4k7CvbLa1lVL
MiNLdNN5G/ZihsN8rnNZPj9dTnxTxJm0PR6If6A782EEZU02IylROmH8Ni4wj0qd
YnvHYPap9mkZRtwgE0XhM9xaEsgPSEgRzwQb0l2uaq0SRj1d98+np8saxuv5SAHp
F+yITjelX4JCQVVSIA5c7E2Pwpsem23t/zdensM5x2Ltg3g9O66rkG7/PrU4UGkJ
vOuJwWa1lVt0HxOD1vbIsu/WfYfw9YJuDck7AtHqbx7riZK0JO+PKoYhH2vjx63R
aGIkxdETz5aHfw4MZyXk6JQlHqU92DE2//qaiP2yhjTiQ/pDpht2/6taUyaiW/nm
rl5G418Omle2Ryjiy3H8gg==
`protect END_PROTECTED
