`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7rmoUc3Z+sMSf7VgfuZvrLz4HQLjQ5LLiRhS4NgAu3SirqfgZ5X+M8lFlWcCz/e
bRyjJVSkckSxPZok179sKSpjv5yBs9pqly4jYrGJS7J5HxUgKg8CvawfYuHwU9yR
+3vgdrX8uEelQT5/1G2owUQeV953F+Unrm1ejj11gfzT19yxOngn4yDNMKBlomZ7
l0cfXyXoEWzNqvQoZfQeO82Y7erbMQoKY0RLaNgGzBmTtRX0akZq4Lk8mxjZLarm
flqNQZRc4nVdQZptIme3ImEJ1rrRXfZlrRe64zHUCsxmxOrjqzsdjZXzFysX2sJ1
MaE3w/3QssSYt8ImZh3WAHxx8iPoQG3kj/FEhhNX/T9MZXw11ElaIcV2lgslyH8q
z+3oZyRxDFZQEyTkWAiNauGz9i2QD9QLLaY6+4DK1vSx7F4bJmm09NWWiY57rjQ6
rgEIx3F6YIf1hrJ0Ed+nvCFb1AEpwHPFyz+rfjZwc7Jga5WUDrNF+LtmQoI3WZlu
IN1GvSnKdVLijWVNSsJ0lXrV+i8bpYAqSnEoMTEicLNX4JMH2AVvPBw/BYaHlJNM
tDMFvMLPLCqTdmZQ7LZ6/6cnHpUm5sd+1Pmimg1TBkS4YyjktMXX2Z4qoCFhqQrN
BRd8qWjPlKaj4iv1jqMMtRr0tShp2BaUYkxd81eQJDgwcjxDo1Md2rOg+p2foTCQ
yoIR6znIKBGrzcwiTpd8PigCxKsSEonnFRF7FmsIZS6WatNHLM+y1ADkie8eqBD7
sa2xlcNafzXQf5S+rLF8eFA3k6TJiPgrh8D39JscoJ4WCIOd7x/5VasvhYbk+KnY
L2fIRc9/6Iok9KQVhdUe9J786jOWmK9t+zK88pSNGyOk6rPEaRKrzIYQHqORp5XJ
VxDPt1smLmaCyqZDK7LheWocv3TiRWqgT1EIBv2fyg6dc1caDVit/6hfKCfyqTMf
bICTJr2/crTbo8o7lX7/8EfLL7lcnnaF66JZmZfH/K6HyplEFPDZ2wegAYw/QY/T
PUl8VSxT/KYi0lIgnytReZxM8/okcNVCfsxLu2xgjwnfJNl7VaMhIvpB2aYHDobG
AsiOHNLM386zokvj87tm2fzg+RK7oUHgYhi3B8a0Rfh674RSSyqHsMLtjML8BpME
XU+XpwDGDOaw8rzqfOKtUJdZ+VI9C1DiqsMmIOpKYSaMXrgn8got61rm1S57ybo0
fFwnUKsvUwZUJTSPiZb8EstO3qI9xZs0AWbDPNzzUv3QIc8uS6FnShvpLnRdmtYN
q8goOtefJAyFhQedipyOlRp/N18uuX4zNtTVSIZni+yZGUdtuPVrLG544Cyg4z2a
5uhAdJ5L8Ahm9d1rr/t8ORUrjuHNOT8hGqy74ZSdh7YJTtzIHEOwcDiSCLO+oA9g
q+w0GDO3WqeI1otMsfG182ge8fMj4PYqhN0XTVXBilrkOZoMZ8VdlIzmeH2mBbKs
FGMesOIJJRMPNkZWc8nEGbXT6upzHDSmXSSy6ZBI25xmRKyC0F4JOkLKt1stdC6G
NGpYfweztL0+QT4tVVuxiicD50cKVRULqK6q3TTRbNYYBXzcd6QX+e6r7ZSNnYd/
cwT6PVFaF/0OJaBtMRKLPQ==
`protect END_PROTECTED
