`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pxktLlfhptqUu8ModTPMUJW9UK4keo67AlR1TlRG3LALYajd3k/gPgrBpEpBdEJ
XG91nil9UH2GVE3VdeTRz3RZFCM6r93V0bhstusuh8pxtIvJXcg5ie4BGBu/NucV
G+5qT+dCVxmtglq1bXGma3FtIk0n2vKgBU6+rJ3S4rsedWYfydxbdBSyWSNzqBVl
8VyGC7KFOb+hEm/XvSZR1440DeNNYJ+Qwiz4AYC2Yx6eBgIZhln4W/B7kOltqGTN
v/jqP98KOO/SyEpVXGxxcQHyt/o1FBxhFoBripOvQWFQvvvtazwrU/PZ7uVmwVHD
23hWskxFLTpzrIFTbS+d7pTvBgQEqT7ML+QaPbbqwimhJ5DmwUk30HgRp0OWO6eQ
Rzs9WIaU9IaQBLLJd+mqlIMrCZDV9hdL7u3Ui9oFJlUQFkZa3xlzB1xFafK6zDXg
4jL/SNSUzwY9ej3jrNnPU4qvkXOse6m3tfLsXZ1pNsO6DA+2tOrMQ49Mc5tLJzmF
l8c89iIo7IhC4pH/93e+DIrqzuhirG+L3A9F/nuoxnhldXp4dHcxsjtvE8OW6VK2
o8fHYUh9GpeNS6PckDd4GCanhB3m0a9dlt5p8vFZRP++Nb0UC8JQhFPTpHc9uQpi
qVETjIoRJ/V8HOcOQ8WKGtjb0NhwxUVDsqfMNGUbgFOmOH5oJkR8J8zxQ3XRQ0sM
Z6bZCVihIAClp3BADivDDBg68snFfHDG5VPfhBgRNZZg6W6LmifLEUlnSKKkeSwl
IbSQdFalK/MFr9h6l1mysmXlJrFY3a00ODFP93Eh6ePAVxx0lYt4l8dFcDMH4T83
cFwxLZEuvWrfH+Rwr2c3tCd00MJUMQ16vELJijqlPw6yvd59EKVdm9ttV6qAa98b
5C+vLpqSVzZ7D6UpwNnotgKPC4A4G5XUJPKXtqLNVkYgu1ZY/1PoFLsqv7Lcqnh2
dU84xPsoLjdS9JtCkV2UV3uFQGnqslPlZoxrfDdq/QCZoiXKFzj0MySq2HOiGtF/
fzSCtnehpu8y3w4yd3xV6JaaVY+uftZVGYFB6Z5HiurTE3jrvqmXz3hNGckS4Vja
u8g6v+rxP/0u5mLXWzcBBBuU9B7sbTZ/MYc2GC/xtwstpjy3geZmfMSr+MHzBuk0
TQz7Fa7B6+dX1hqTpzlOkDvrH2FSrLLoeDYkzQaHZPogaFMYWLEzLf+lJmHvoe1d
+IAUU/WOLN47Vn3Us4EaWX/Oqqn+S5SQW0R3tjMOymH6ArMi84K1/WMEThPh7/4w
3GsWlz8zwqGq9hT4RH7BxYAVBRqO4O1fe3IHyFS9DiecnruSBPmAu8uiIAS9MFuD
TMJcMVoXnaw4G9u7sKERocZA+i9XK/XPBMxuKI6BLOzrs5y3fiOAXmyJ5wrZv4VB
MA2JzORL8ylMmme5ee84l+rUT9CrCcmtfkMrKVqYgh3jNv9xU53JAzbQ8J/iaGdK
wmOchwRPU2NXLKVXQCdcjxG0bmyt6HjtPnvxu48NuJtRy6ei9n3f5bUxip8YBFSp
zwsmcoA1SKlH4xptZEr4zf1N2u3wcekAfx4f0/uS9b9OYRH3ICE8jcXmJJ99N2sf
`protect END_PROTECTED
