`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CyUMofE7oTGtN/A+6KBG96vrSbMIg+rCgYQMqWgassNMVqBbFlFj4sqbk0K3rcKs
t+opDNPezJ59zp6Y7HvvglN3oKnhI4Pek9Ku8rCkEZeMhtN2zyyAluGFNstX6Oix
+t68MSAIHrquhatFFNsPCEBX3XWgpsb538+Td+2XiBPkiFDdeGjt09Z3xE5+pTpb
PPmy7V262brgzNBNj4bSI67GXiGUleuaNeX2dCFnO90P59VksiJ+2fmWggAP9mwf
qabPDpHQL8NAC4HA2+WvYPso7HaU4wDTn2Or1QmsJvuNfjvxCxXksrUQJ0mnynAE
IPTEx5qMyYP3vDj3+zFQaSohA5oLU8IrgabCA94f1awx5cw/7OFwvZyYGPtqypTG
ETCWWTcFTClYHQ6XbV5OT4cozYH9KuAOnym3E1E0zy5btF86OTeUVgI6iU65pErM
LFj0PrAkAYLVdf6YL3r+1CSYoOxyyAQMHuccxzXK1elzabRY7x7YoKQCjmew+WXV
sJbNSQ/CfuYoV8lmaCOOIxrAid2Kc8nO0wh1XkZBshyel0ypIG3401FGj6TsJdVE
UWVmmDG4xUxj2HC1n3pt8C0Uvo18jBH/3pMUPyztyXiEUdvIQZg+lR4Icr9Jo0bU
Q5Zcut6YX9h45tPGLuY9Q3AJEpC5wBw1UI3wQvlup3p8GxrEK+zTK36m1tQRJEra
qF4Nnk5mWaEI60UXteoXvla8iVwBXRVROv+ujfkjEmI=
`protect END_PROTECTED
