`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiiB0Yb+u8mdFFLXiDFf3wWcZ7XhxpB46iPU14BTXGKJjNp8wuHFwR2h7uGvbce8
k08qQ8tuo+Ydeyvr/iIlQh8RQJa65B7l8kxbg1qKWxiTJZSoYq/rLZzMw16jADp2
B4UxjAjzsHzQ3qttLE/MW6Fh83HbeakLL4wu/PEFIeKgSaGe/U2W21hvfCUjrRP4
BlzO7pPByr90eGjzDuun/LiyV88VlEsV7wblPGsF83cR2Ys2Pw6SUxf2cuL51FAB
+NysuohT13E6U+hPXSJ6OOA8djYm4IIshOrdgVoR8x83g86TpLkRIzV91eQFFkpW
LYTjxP3EMcRn0jTBiMlfY1i+XeuMxJgkUDBr84rPQrziVV0byljV6SAj6eakEslB
krCZncaDuuFFK8eNQUqkmfPgwqwqfUvSCJ672hfaikNhOExX8wxoGMdgVnw+KCuN
x6ICUiigRWlQAU7HfsmFuraG/pNap5NaAUaUNNJeY3DLOfvqVvFmyJYVedlZUIbg
UqJeMO5nRsWxDlUdg73jGr3Ywb/J7ci/8cLSCrGIEukPYh60AdMHgx4W6vGVTXAO
vnb/m4QPof42r5+EH/DqoZ8qj1QHdcELW+G48qRGb6Wm9Dx7LonARNNM8WhbdzhZ
EcguFARXUKoH3cVSDmMoQJVf3ZDcrsueBoo2S2am2rFpXUbIvC6i5hYffzWaLG4m
EmWJWkd4mKlf6LuGWn3i6okonC12KMZjC/beLJtlRfRJpOeEKwoF4puIR4x3oREa
jN9rVWYeBj4trzmjblrEcNdanKyM8ti8ttwwmC6mOyez1F94gtJQhGlK391iQ6U3
ehckg061Pl02P2Bc6B5EY7blDXRZlRoy6LTRvqztXbyB18ceKD+K+vnnhjejQtiX
PIKd99tdceaQ0jaFY3O1wFNH4/pWf23a2GpcXMjrrZ/iSh7UAeIVcWdEE40nK0kY
0gCVhH3rxxuOuil+GG20UbWswkvLRxGtYzuZxjvO9G5S4cXa6ZwiC1UkWm0TG6sJ
Tkd08f1QB5gKsrgCGYlp5PKhGXGUWmguJ1mjv+ptU5SiRvBeNgc/Sc1s6gVt5OHs
+044epX8O8qsP/l+a8l8LdWf7O09dWSdQ5gxziUM/7yZtGa4HYbaQKFYuy7zDonI
Svo6iMxe6YD/QFatiQy3zzNQ2x+wMqPdveGos82nGeJFBpn2ixX/BiyWkfvJefsi
hrbXj0IiWgQRljxyYo7qprWIeDicwfWMMLkdY8dEW+DTVL/iElIyVO477mNocJJf
i5rT7WwlIhsyOPWLdsiohggV3g2mRe8gU3G3vI5Csyk0H1ripAuh+CNNU+hu+5tC
NHyST4fmOyxECW1PlwDJ4UJO23XKK//TILaOa1OGfRczBT8/NFVj1+Dn9bjgzi1i
4SDNHR8TWsCL0pVWcUSBA+FkN5qtuckGs29O595XFxxG8MJpV2zh90fDit1qebt6
eNtvprII8s3fsGzKbSf5BLv1m07wPeLujpBAbZQGa9BCYoVYqDSU3uzED8Unf8v4
V4n0ZExsEegDJn621yKL+T4kxWrByObBHvWUKBhflgeLGvsUIhfxClPvu1CXgM3W
4O2NqpIW8rcEfLtzR3B8LxOvBX7MzZQlFMKBoXDzeYE4Ouf4hBOL3fXgfUQlO+On
9B/pCGDbZMRRT3nzVl/FLcVS+7IobYZTA6jF0cZI00WdfTqfMQkesZtEhsBojw8j
b/xDmC9Ygk4rzgcsgg+WrcDbjE/+2DUNANanyt5z8ctvsM3uGEV53LyL5PeWM3/g
4nEkmXnH1s73opKxP4rhvSvsBE/K8iONz7t1rw5++G+ZMoZiuW4/FXtvSjWJ9YrA
x688LoW1NdxZRv2ygqxMyoVK6YLOj50GU5fyHXVj7pXNfqIQLojrN1XvAvIV37bY
pHdE5QTOP2c1zFznvzAxAbzP1D1NFW63Thz850kCLlUYhoK6kngXI/lCGrSUTXbM
86HH2e3xDNnr5Hal7OzReU734y+QXIshalXM8YVfy5SAXCesIWqX5huY/5ahBGI+
LPGM1KMeHEe7IUC3KpTIj2CF7gOOZe++M08TlmtDOAwEf69055omTfCUcukMgOGL
24dXFmCwXYO/z8bS/k9WPBMRzV7GmhFbVck/S+PFdkXT4WTPlSr6+Qf3o6negkTo
+JfqPJkvAw333IRUgjpamruC1pqA++9fRjqrWGIXcCzAmp1ciV+3PFjbv8LyonS5
/kOdxezA4GqPdiK6OPknZgoqBAHsdzN0WwMyu7dx2q8C2S8NgCYGagSBlVVowNw0
+h8Ps0FKKTtP7+2rvudvRcIgXIM4HEG4/TYTAwX4dvEh0HJH7NMYLW9h7ueMG/HE
mEny+OuHHAS45IhHlMRODBP48YvTa+g90veXKZjbximcM80k4c/MD628dT/lCVRC
YacTWahwUUsbH0vVi0zOigBTEY4crpPXAX4+ftwRJahBnosmJXPRYEeQYNoDt2vZ
6CMcrciEHleFaoyUit8F6382/nqk7plzy9SkyO++1c56YhLYBB7HdHSKwO1Mbw6r
u2wAOfAi5H+9YEE11+YeWRIkkAfyf8zadPgDYK0Uwh3AOfED4oa+G724SVfqTsyH
GBvjm2Ss/IQ0JmMQaourpEmGUDI+qKqNxt3VYruruOzvzK2XLUSEkGXzJ0M95aEU
c3n/15TifqXonkorjy20wUXmCcPLinXuyka0b7BFV9caXPgwt0rJGWKnSQ07Q9Vk
xeJzV2LBq9DblGcJ5XLfYpcPuEYgS3xxtbK5heGywnPP0obR+6+VMzBQ9WcaFKBr
zKEKTC/F36lKpwfgx8r1qBtDx03hQgXVm+pzQqoxC4BE9GkeCtySihx905YlTNF1
ur+OI3fhACJh3Past1KX6OO3OMWLTWoRDVTZjhwyoU3vWLBn2rWnDZHnJBDgPPuf
E6o6X9xW+WQwcAffKnG06OeakW8IEe/TfG5VkC7AglRhCvdNkSDSteERC/VnYyFR
a1jVWLDpLOwPDSMuWGo1Ga0lKDpm8jq6MtRRaQKdOkQ53q267AnmlBL/t0wCybp+
VfA/00Z4XrWglCElpaMKVIv2iCy2LnpHvXjZQ+MrXvVXuuS2k0W8MGK/Ogf5wLra
bvWSN4YIK/bqefwxzgYAuxI9QsM7aJjehO8CGFnbNdG0ETN2C9GlsAA1DNIeV2PL
F5b3xsBdOlIFcAHXbwscdE4csW6HznqQ8BtADRrs/CKo+bJvaYXmverTEwerfh2u
koe0jfq+pgLqcjb31cQkPZp8PUCu+IOCKr5+lIYhi9e6gu+ZovedeZpg40YreSiK
78ukopSv5CUsBH3L7J6nOXTEDSUkMrr7FxFZyZQMgekIYVhjIhGR4mJmvdsAgYET
rly/d+wPeOTAwJg0hYdj7D610hARkF7gHxwfZ9jsyN6PYszkbF/D+RIb2uzqzlyH
OYar7AXM0X1Q4KYRbtJjRW/EYTt35qd5QuBj67fbe87d5MRqC9t6YFaA53zBwChR
Zxn6Iz20cOhHOxZd3elsl9QjxA3zt5x/b8uGpcciXDlabmc5AwEzURQn7ze+IBT4
G5hMJJtapf4+LokSXfcgThxSggbHIlwxBo9uZ0OMTx0EwFWD9x447rk6ep23tnpl
`protect END_PROTECTED
