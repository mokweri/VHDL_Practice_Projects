`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GlMtZ2/24itLhFviNTOgKvUmFE1xnHRePPf1TqPZi8idUiKamBQD+hSJOqbv9d5w
N4mXxUqeK9/fWQvt331hD2qoHzx+3+2aoL1oa+EPMnGm/kGnC8e1kLf+XROrz4Mn
xKN9ttQw0pk6qtMsQbTtYmm3ruCkOLsnrCF0NHVALBWGjd0Vd0eifpSqjfeufqOT
MYtQ4OsicdvpUnzLE+hrqUYjuuMUUpbYspVc4RWtgC2N107x49A/sM/M0vPBau5d
8hlkr9SE5jgIRAOgKLWoBhgm+QIm9aabePh+fO9HdXCWNtKuU8KVIuE6KTA5K7ri
ctpdjHL7RdAfa4rs5IVZqKQDycKuA8Y9o+uiKla9HRGKz9HW6YbtcshY5+QDcige
o5MJl7KMTXB5UvYz+V9cT3ITH0kF9NT9kiACl69OpLVbOlP51Oxowry3R+MWCc5C
uhpgJEoQNex8OfAG0vUuv/CCkx9EBdVhujdixEhMIJOr9iiWMQI7rMKrSHr8G/Ia
ZCGNgPzvLwzK82DtU2gw1TzVBht2Wdl7iESDGD/SUWDa3noR1ADr3XIWQuINYhGl
hbPNRlNMwSxPxjKb8O5Y7ChGE8iPWYwXhyZ5/xxqGaziDQTkvh+qZtk87bf28gv5
9fqtGrtHasUK++ql1sP8VCLvDdO8vqRme95ZU+fT2JSeSv+njPwkLvbcxez99h2Q
hO0zQV6n2nv/tYKmZEnDJ3eyvQ7pYWYKDSTUFaZqTYrCyuASxQdL6Ks5qPHxoE9j
RhgmEMJjp5SZFeiqxF+tnn4OxI5LkPRETq4rPttuKsBfwe9LBXqZqGP5AEu1ZKgR
uzlCMoVQdk1f3peW6lVBPRmnQgHoLUUJIziGGf6lA5h0KP2PaFiqi5MQZssuiU8B
OSM460hC3IIFqsT3MJZjJ1svPD62KCfaoPcYZWpaqTrGLPuF4z7A05ZGyg464S9i
ENAts0Ixf2ZDhDF/4koVEvm1BLoXiFZmZ46/7ftfwrTkxju4TZu4m6VRaM6+w7Og
qnIrUb4r//lKw11l68jf6du/y6xvVOmPT78SJSslTCSWy9eDq1hCEvflk+nEWtzI
DdTegTwzLntyn8RtrXVvFi7enmrIX2sYhLNTdTNXvGZChkLxe9b/+yC1tfctkopn
pwvv/M8fF496Qu6EdGeQ47kCt6xxOt8jp4HqDz0/WB1TAl3O35nhWrJJEXKH87lR
tg54GYPPIlFchQnf46GhvD3Waky+ngMS1GfKrQjAzhRd8LZUu1WrV3jW5PNK++O4
EWUekN3TI/RHlrzxqHm9DQJojVkm2Ztuec4exuZSYxeo7myV7UJCL4TVL3Su5Cp/
nYMHuTj9nV5cUOcz0wAIjMZaj8vIsxpuYtRrUEgoJoq2hY28w+brVaLsizbh6Tiv
ojRunwAahmuwPJBZ7T/L4vRK9eXVhuPBpe+/JFdS/sXMRStJChCDYXKa6r53DKLH
yAuLIQnB5I38RbMDUD8Pib0AA5rkyr9RZFZrpemBcFe8rFxFKGSPXFQC/yBjyV0H
4TpBJ7ym8kzNHAX3zlunzjW4PrREfHYenhsac8/QJWXfTSivqhwGw4/ctDrJGztS
NySOdiBkjui1XaNPkCdnHIE4+vqi6U9kRjAXQ2kCPa2x5HdOcqtiYPf2ZhrDreJ2
M5TtXWAYibqndeJx77lNHKdDlnMXlGmy/81w0AmvZeI8FLBICN2cFY3iQGUeG5na
2ycqoaC7tv7PCmLqv8mGL/fYcSdcmTzvJt2xpj72AgQGKS458fD0bxQgyut613EZ
qSZ1n6iFPlZz4Gn0aa87LmznYqm7PFYTfGhcOWc2udE1f6xYOIVn4u4pyS2Azoyx
G6YCaJgAcx63BeWxcsQHC8x51XDcCxK1cjoHQQ6fKgGiY0Pt5OC6GfSs17jRv+uF
uojmRZvzcTk90crWI1qFXTzLk9B8GpfG/Ivbh73z5+c=
`protect END_PROTECTED
