`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/Dsuikmlu09V3uS6ea72zRpNVBo+LK6wFG0MvSmTxsZM74NEXUjGF+eBCE6ioAt
aKMaTW3oUissdSEJfJeeXZeYRMmbn0cXSaxKhCPG0lyeCj533gGpjaWewfW819fV
lvyTV++HBJ3ncGB/tEQiH3ISCsnUzdKlw15Z1XLY/IzR7oNftkwAc758UbBSpMb8
oce6OrYvUwXzHM9Qo7PrL+wtT8CO/U1Y6jqn1azBfR6oL7dba2koYhCcNHxsqAyB
hWZWJJgSDAZLiidM6fXYDYGI8oVQAd9ljPeJDYQr7kiVSc2N8mzeF9RrJwhycah9
oK4m0XBGPN9NxXPqHK/RCKzepZuGmUmntkY3TSTQ+Tgy5Zpp3s/nBCK6ARBaquOY
kWuI6tTosvUgv+ljGihgiiU2I+J48tEtjwVasqMz3hgKtBZQffaOEYezhwYLEZsG
/HDIG6Yg3I99L84DEbmum71tSEA+yo/topvDFWrr5XDdFFwgC4/nW0jVr3hSjVE0
frixCiFu+i9YoodtkC7ytZoIf7EfYhHJHwLENBBhEYM1RrEzCdecHIqk0DuWtt2I
AYk475hgyyEZGiik+AxECPn1jzethJ62F3o6R/viRUw7HFoVt/bNjy7e1FjixNkY
ux/XW0/ySoBvPCR1ecu8yTztXJTbMTu6oQIUyBO74PnlvPMMioh6WAQD6v42erD8
fhNYYjYVhsFIS7GpoeNTxDUaczBScbZKabwY9XcL0U2+rmIrkOli+7/Qyen7Dj7m
uiai4o1gpb/tGrUfYGn+znhyxquUMbg/Oh80lJ/si3o5MgS0Y9u3CbmDfD//aooK
ajHZqxY4l/KNGfuvPAE56gIX+XZvfXUWfoWcLsQlhY6omOxYnMBRmbpaVOhT0Oa5
2rwFyGi+GfEsUOJ8ids+RV8ZjiMofWaXloJuCV0iOzptL9G6XgTwlWG2J82Ffrax
i0FftGCU6QLm3dTttupkAalHOWmq87QZtgdTUoMVoprRVFEtb57JE//ni3LjnYAz
Xd4Qne0Tc7cEAqRYtnfwhY1Li/L6KU2IuN1gzEKltemXidUrbN+9P5VlgF8YvsG2
l7X1cB5ZHzRSjVbvpEgm3OM1wnE/0V8IAxpCBLu5ZFy/fdufTtJraLBii7D4+Xnq
+FiX4wz8Fl2wK8F8AUVn1chSla/Vfeu2rbFIN5X/DjFk1Q48XeKWZf333NZtENX6
jWd0EoevMzex1WXoXC4MMJBY+DLsjV1vSRPRrhcez0yJIYzh2duj7ND/NH5Ch8D+
NyL6a+U52M88UaRHmoJrfh12m7pR48Y3u1SeXhXZe23fpTDk+ng2fMa7szidJAaF
3Uaiq3k0cJ0JXCFgvaa0LEGp+yJGEQdYdZJZDz2NM6jNduFvStxw0Egomc0YJCyq
BpT9nU9nOofhx+jtvkFCQCKHcPLyHOxgN8ivmrt78u/D91fBQoaAMRilD8bCgURu
6gyndbr4bmelpYo8oypABCS/BmHaPkF5U4VoUmDrWV/lPKst/9rEMmrIjKt5CDaG
N6YoPpvrrld5ZBugzpeG8J5JFnYfVLwst8ShNscgKdLd6g93n/ksiUJG0fImBIAV
RxOMt9iyLn9cbdOFGg4qthhLWtaumTcLXjuVI98rP/HD7VorktcbLTbQNRc148TC
n77PT1/ZKy1ouyd8mAOJxSJB0CfaFczdXHLEjuHoRRFIbIVLcCjyOu/5id3nEWOm
mZCN5Jf9an5rMOC2GahjrdTurzdqeCML8He/GSwAx5D8bf6DrhBDIVX3EDI0w/1x
REd765lImjSKrw+4uGnnULZsvoxo8EVCSAPDPVPSUbzhyY3mNdF1nwsucyC0uhtp
Xqy6LAfRZ0AmHgorvLMQUlcDCycG8BDOw0p5r9Z6yOmpXKy/cI5fbqbw2tcGPW8x
yd0VZGa0n93dYXqv7rfYvdEciDmKcDNyuZNDH2t6B+wR7fwBwIFvb+T0A+HgSmR4
sbQWs8bhFahnG9sTOAwrI2RJxKqpWlGoQq7j6WKWNeE7gClBJaf+ftGcXZR4Zhhs
30kHqu8Jmol85ld0znC5XW8gdPYlOfLVsTNXN4Mx6KFIzqvdgRbFAtL1qzvULcLR
rXhzYSFB9ZyvXSmXP/wLSQJIGQeZQuYgGvxI7/nlD9VrkAhmwhJ3ITOjF9Wq7wwn
JqRuRIUYiBCwiA8UShqCq3nGEwRZjmoGwFw/WVs+IK2UmQE0f5tZ7rsjW91lfL26
uR7YOiHv8C6RsL8lT21XAMzLvH2/ogvfuyDsw2BPwiUshKzcQb33LejM5KEiHX/x
o93NI7VZKBV+wbsZVkWQbu0VHVGg1UKmgSM1ORTdzRJRw5lNWA1ZlKAEqqnm8X32
v2vJIKHjZELT9dgyKB38hRbM2OfiX4SClZWb/8sDbeozOs9TI48WBzKnrXhGvHdN
oJEc5uD8duiDAFmGiKTIUdOK42ikweNzjKK/ZsjnTkw+9aw0b1K9BotLwJuAT/gM
olNuj1H/3kZ9kebybpH1MdI8BaXjsEpoG8vwQmpVYlelBXg8gO9adElCBYZx5J63
rf3T6C7Hl+K58Gof2JpbERJ3VHf8SbuCWn0UjO9biJR9RSQgP/DeKpxJcMzKIK77
3doXcSgh+rWruczOIsDVvQWr3334SXieiuo/t2UelpYtO6jwsfGJRkA3e+kJjzNV
Nl+kLVYvYK67V534O7Tl1jbH27yvHe9C2iTQ3YIRB56ABCXjHlJsQWesKiPSKO3q
echQQdxkK+MvXtIRs2oQs+LOj5GPPal66AVgX6C1iMld0vUnlgweN6pIVbVdqCAf
VZPpww0kDuIsXmbd1Bh+GwsjxANLvRWJl+2nQuCrxPyi20Lme3QBADRBqQP26H+/
uk+3IPWpGxpPcIs+pVh9srjQF14Lstn4tzrtotWIkGqwXZ+ojSYE+8giz4BIqb9V
ScIvGEx+1Z5IDsW3TbUYXRSlzBI8cv4jb4EuCmQSjyC4W8R8xeTKyoJWnfHA9pfP
ENk5P2QqosciidncedrPVQqKW5JDj8h57CMDYCdYTkNdY0JYmmklzYpAfzCVtHyu
SzbE/jhcLvTgWy1KftDPZX2u2sxLLg/17upgOp9l1KVx+QyBJGGIgVij9qIXtDn9
f4jVUbSy+oaSxh2EaNPWmQ9r1rS2BcNGcMu9ZIv3utLvr3QtBdHMXhtutRgsdS5H
hqaMzo87z521z8mIjf3wNSLJ82pQzxNpS/uk31NTqJ2d0fMt4oW1R4zJssCf4JIQ
HfA7F8XnXx38Yb6ar2O4bPpOdEWZNe8Az8yTH5LvN3VoD+6Vzp5Hha26DbHmWFD6
dNP46oYoRMuctmY4YvVd1M+lo66PBqyoccr8x95FSZX70yjmmjuSpysNIYf5tXCq
kifzDLRZTvgOueML+14qSj5EN2q2VnKqlYXrMs/kttDM67ZJxYcsLxjhzLgThkXl
2YjsTLxusQyNbAtyFoR6Gkxdo6N1vM4KscjURCe9b3ZZENRzpc0vG9n7h64tus/e
WbE2lHX6ysoll5MCUq3oX9YIwbPJMcIgp9/bPi64x2KieoZzWEDFQ2PhXcVaQZ+E
NyaM5YCJydTifA8UfQEv7wlLuCDYEXXt/PRVbsivRuersgVSWWjjfY7FcBM8Q16h
SaXZca0izCbCweCqhClUPBw3sifFMK/l0eXLniaO0isZbBjXKXDtY1HP3ncda0sj
a8BAJ/aYCBxVJKP2QO5mFRSWHCUF3XvUAtwY/E3Xo2YtYGYgjAL9/7hDxBfxGxDa
/3YPjDC3YrgT5QiSYOQ4qn16k09XrV3GLCWFBdk/sLYQjJSLYkYAQocY5m8jr2yv
gpDDofsNm7+AwA92JOXpPMw9vk2Y1aa/OQNG2Tjp9ivvw9hSXd40qX/npn7uQepY
zJFmGGXqPLffzhvLYMzALlpEZgzkVejUw40MTFhVPuS/xgmzzLdFybezo8Z+HWF+
sL8kddA18Ns9Ek9AP7vdAqOZGPhYvohrGmEV6ZIdDfxu1qI0EETsEuWsHzQoSsE0
C8RzE2N5Si+HN5RhoaTGHTXF/KM4BXnqpx6zbbAhWbOI0FOXo09SPBCzPAxMj1d8
0C8Nob+YXbhkjcFmlA6xu2alzddqJsQbXnNNjgV4sZhfw90YoVC8SakT3FDii0VD
4COnm9mcDSm9yCxWCcywpwcNhQUf7djhKTAMnsfveznHFuSsaKFfMGLIN5KAGvo7
fat5An58kNNQHLFoOZh7Iydu83Jn0QOPniTFOaZwI1EczaTBLz7x+uNxpA5bm3xG
yHb0jtlrKEObiICWlMsf7mJxcr7X+ns5gJW/wlWTGx9GH0Oe7zCtjnZKpy1zjcXk
OKKprU0/axl0GislJTwkOqakgy98Irt7i7E7/SF7KInnNGfiYASWPHNN6oPxShAX
agX90jre6HbR3u8W/N+LbCurnSLeadzOx+ug8z1Ju7FjkBEsoNHrsPpwpgV5WXuh
OngP76cisFQFCDpvimoS2pvolVlVYttjc6GN+fRnRyvYopigtDG8NQTIKlKK95yr
n9tCQyGz/nMHwSeYTtD+2rJM7xN6UvA3/P84FQm4NhmtrFue0v5sXgLXpPjtKbrn
+Sv1P0m4DkM4PJGSPM8cLEhbfVgvhKprcNYcsCGWZ3w/zgGIYZnUUbrAPcn+CDBD
On3X0zFEOBhd6Pz09g5tfWzsR86G4OnvSP6ONR4O8QZwYQ8ItF5Kxk9wv02Ph+vu
QgBAa/oz1eB6+9R/2D5qR5vZ8lNZAO8LuBUHbm7HVFY4QWptuDce4dk2jhP6gDTf
fgEGA8sJrCEB8UCf2AAyc/tEa6Uhw9PkNQmknp75CZmzCSsBI1zPfCDq+Y0uqZJr
A6Ailss6FF8fQy+yIfeJn+7XlCLCU5yyZM4SxF++gv8RBLjd9l2DkFTAYOoeJVnf
WUsVPzG/3MOrSleQTPbF+leWXUXoBAd3a3DzZTho2tzvA7Fzmn1YoV9jCHvNJbFX
B5/Vrqxs85lOY4MHo3nG0BTkEufYOccH7dn6IomlyKjMTtr5DIy1j1LdapuEP2/v
ulEHyU9ZpsQX+vmubvlCoG11oZNVJ2r+Z2fr3mvkA9bKDgD3bGOMAzxzrONVB6vl
tA65RquFZiozFGfwx4iDtQSe5YJUDKhy5XiAWzqWMcvaYMZggZD49jQgYrfR+ISE
oxsHCgBkXXWP65UM/FT5amvRUXxpHv0jCMqxxR4Ma+QzRNsJV5Jcvvt9GAmnA7wI
FNMBPC3GyJ0lDVspgVLZ+xf0Q9iKRkYqmFBHTCyfo9PE+h0kpA7aILmyYJhXXO5w
svbVpf1KHu+AR/Sls2RleTScl4Y6bqxqr2Mj3JNqLyEZvv5EMPBXQFoT9CQI7OFV
PPaPCwHttYlYim2W+3MhZB5BHld4geV5woOvB3w5B6pgsx2r2VhRRbYhLYc2CuZ4
pWILNUuKSLz3Odxm5iBic5N21NZIZMhJVm/ZJT56QK2I5ihb561k9vjSMtw2ksp5
oqxA7JQ1GFt9V5sg+im+V8MoJZOknsl/+aU28V00fy/LX7IWzSe0DnhTIXRpBJpv
71Enp5R1iT7HQ1pDN0DfBG7HwRzRW9V4EOclg5or3ZTlrUi/5VivoahBC+oRDH0F
gZ/HDlVO5r8XvDhAskLDOky25uI0WT89ceR0VuTLvuOzD0L/bFLv/gQqSNrxAQXG
Y3NZlwBsZR1C81PrtvSM2NhrQCRzZKkeeu2t6/a6ij+2Ra0FHIBTj5JPmaG613tg
ON4zhbz90blNyKfsflBaNhNct2RpMRBanNLVbqt+Nsfc5DWGoAp0cZHAiaA/Uzn+
FNC/A+XsGIHwSn7qo7gsN2OZEU/4USNSxTRWSGs1QTKP69y5z17Mzd5Z1MCSzj1p
jT1K0bPDbU1eVGRjebnu0eirIA6N3tf6MUSfDRIPxJj3g9CKj/dpHnOO394vywJ/
HeGl6l+RK4xloMsufa1v5IfgwWLQSIFd+1P2bRz7ZJ+d43T4udUYbotYCzmUBDmQ
LUYyt0uFAwIYy0sm7Ep8b24GXiiSpVN46/Pi3jmcAWlYJR0p28gyb3c87IakAD7/
sR1aekTINPp32qlxjQE8Mp/30a/2gBxm6IMcWRGVdA9zCSceogelrV5yaQ0ja4FA
OcI0MJMpEKgPcEmUU8LC2/QShD30ploHYL3JeKgjtZLlOqn0UWEJHR73U04jnuKT
ZhRpv3VhS7BNyoOVqx2gqtuH48mcATEeVps+m/TnBAbmnW0HapoeOJHS840REqwQ
7cEKVtUi/MqyeUWYkvINL87J9A2Bb9k3Nj9U+CIJ6Qy2twT0ed4Se8gKdbR0k1WG
34VF5hbAR18rqqu/pGAX6+TOhNcoE3B0IkkBf2PhgZ8B9Vf8qJCAs9EysKAyjmHN
xwCYhR0nahusE2hND9b3fbZDpviqrt792PC4jhtw9XsN3/A/yFZKWlXg1HYwedJM
wcdZzMTdeX/wNw0ah8XWnozRoplSLInJUIf5wX32CBxURtpM12+wAEkInM3gV0zB
GYHtsvFH7mpMYDOiiGlS0u7oVbP1YxFRx0vU582moHB28UzSTruHeErEcno+8CTW
YhS4AW0Wh0I8WcgZ1FlqStcHqV8v/+CZKgZBgx27HTiDA9zgo8HgVDWNhSRu27Tk
H9kxC1i1dlVAr71MPY83jQrt7w3Ma4xQGNsT/OR88SsehGh1maaDRJmQvGY9Xxus
DWm+zW6eKoK2aprJiUlmlI27Zf0UsII1hwIZGYRgg6b8Gu34yIfEQS/gtFQm1+u3
5KfphGaHdCjSgCw2SkguKo2IJQ5Q13LvwHsTE4hszUtg46zvPDJu0q160aaNxRTy
g9PL4VxcVwu5z8yfDJnbLknfdE6oW9zoRCXTL83dixZtRGu0AGcnX9s9/ZO30zFm
oXbtuFNjhTvHNDsztJyn3+OhBUkk8w8idJOjQVr1HPkuL90mQ4CaiOjPL4aV4sV5
CqvHHtAWgSdCbK6Auv/RUKO9ICZYl7ntUX/s5t/7x9M1ck253ckPe2MbCjraVlgi
52DRoNQGHTAWjH85F1mSc1a+U8llu086TNVEJGOfj4LgTVmCmv1LIB/Lh76Vep6Y
eadYBJ2x9Z2go8C1/P+yliiGF0mECNJvA4rg1L1ChRiZ6pvUABNjimkrBnmT29kB
LelPKSM3k4GQOhn0zvctwoxRVkm6oKY97NxxOkicLcIK7LP6e2lKFUyhH8/ujOVu
nTXkWFvZx2q6PaM1PbidDKk+dguZEW3lgt4vJcTWSG+4WRNK26MGqbc3uvlamY72
a2lliVBFTzS0cidKH+2sT/2yvmX3RyeT0BadYzj6hSNv1Uq10YHM0qwCnibutLvA
8KQNNYkh/lsAOwgFMvN/d0zlF8cboI+afQqMm0pC7E9j7HE0ajFg/dRhxI8coDEs
rg60zNZljnGonlRgiJ3ii4ofKcgFl5DIzDivrCiuhw1EFDyNFNdZEigjzqaF3wQ1
oaLMpuW5FA5hFEDvOqoQ69BBLROx91OI9M8b/Hi7n9OcSMyV08Ns5d6qiBP6V8bf
Z1GfkmOuGSjS+uiyr4J+AEDEFrgY3LHKx0nQ3rI7Qp6rHG88WwXWsb/15WtULR13
56ha3IxSVxgHM/U1p/BKN+uoyllGO+KzEQJXo8eE13MdNuMBgcv3DyP23IIUAzl5
MZBDUTr/J+I0eCX7pqYcYZtVQkR6A42LkpsTtW0eqbVgU35DqoVdTfHEoakfm43g
f2T0EpZMPYklYRUJMXZ+X51l7mPkJTJ08CszqhF/+wmmy5q0AdNeHgBJMwkWmGMg
ecuBzDMhcUKnzFrqfjnyseBWtiU6vCk8WbZVzvggSsVL6i30PKgzaGeWaga0Yui3
KDFJgq6PXj2Cbc6/5L3t5soFbDXcsX0rzR2C1iUjMJ6posgMFtNk0/aplcoQg4zE
OJ3dGPqODphADn2vxOhet/Ap9uQ+4ZvJ06P9rDCFcQnSqwZgijKPpKx5KS3COM81
M/TsWrgjsr3giRL89P9Im1n8ni1kMHfvGxGhICWWVVRKXvYFbgNfRu6ZiumWwxVO
iXedNGtdEXTMPR+855ErTkdkOcCnO2qtAw7q1FwvT0mvatwhhqhcerzNzQtqmxtV
fduRrb5gcYBsUUccN9RdbOGuAYlzLR0zrwG4U6odTQQnNbdQh0Ypt7XSBjVqMcVZ
W3QyIaIypSdFhEkHJXrxHPn5njahxPiLbv1FeZlTuZFr8sMgD3JbXZUcait4pa0m
OIehG0gDWT80CC8TN3boHwJIzxkeSkWR2RrrdjK3/ZZdc9VIqy0GNVphO/2hRhQh
uNg1RSDaHf8w9dSfKkktsZxxEUiqZ2SUMQum4YJkf7Cq9WaTkgOmcqyzuauG6dCR
dYf7YeovSO+TriPvNI/TyXftTtqhQDCuQBYhEOmjK32p3KSQ8v7VfD9GugqW3fNa
/QQNzr+BIbI3KC5EQbwdFVLzKrS6U/9WFednIwxX7qp4IMc7JGwc7byeEc+LhdSv
83K7ns0DbO6eMlYhOOi3ButOu/Us13MJn11bffJTa68cuuwp9jyH+ghpPkR/VDqC
ELxsqooj8rD58NDjJ8SCWUecmuJZd1KruKAV2zc+p0rGmi1B36gkJmXGVE/HnDS7
ksoSpYfY/3lxkK1R2dTK3csd44IrNx5vtUQArNYdMpblfVG00DgKejXicbVzQ0US
VasPWCe2pogvXkexElcjWCdcFZhMIbodeULlSPdF8fqow8HyytuH26UA266ikwhz
fOjWNxz6bNEDBsxxgN5HRiLW4r9m/kmcHmGSG5JESW3Wwin9N4YLY6mjCq4nc1Ff
sgOKKIARyujQwk4pRtXs09HoRHTcWcK8ZEOy9VROob23uJQUVwkyErnf7jLH1mnF
Y6UDFWWcFWwFtj9m+qTRrITqht/DxdauDD9AbH8aSd1lCrAin21rR685eHBF8R21
ASNSr6mJ1CX61CbJmuCJ9P//KOiBmAAzpu+Slwey6clm/w2S77RP5KdUkXrfqvmu
uBoMjdCCodscFU5DfqkI2HiIm6G9Z0O/vwGBcWRuEBqlYmaFexjNFEpz2LUKXhST
BI6RTq7+iPQDGeoaHsuIyhhLBT82xbUQtnGdoa/qr+csvkDIO4O1x7tWcYxtHTgw
RlKe5hflr8p8Ixvg4yw9FknZ6Me3R4WB80WhRRaFowWW1zaG6Dp/5XdQ8as1GiXG
wJ6kuP2uHh74Y/kHv+Q3XlUSKBWoyXMXBBXxGZjBOfPUQg9DYpcCagA+A0dsNTn0
vOu0fDEAexwa/nzXn+6T5S2MMWZlN4wBmeeRQC1KBjJePAvb9G7zv9fTt6gv3dOA
UhjYZJ50wP6f44S6RXkrhY6OioFV4l4WISstr4UpI6PTedUPEEP8s1uDcFiQxGVZ
Wt3Dg22FlCT1sCCqplxlHvbIQv5TlmsV1LIZJQ7HXDYWrhg9AXVjAgubmB8IU6dl
qX/yYbfICJzTws/NYZIhqALkQ11yL4Bc/npeOm7OwqXv6iwygl/LNc3FA6pttbqC
Yc0eeuKCPF1qVn5sqG8KlEX8J41BxBdc1oB4lL2lzyp23eoIzOu153TFmGSFLK4Q
8utydE8tZS5lZ5fK4wyNPRVM6r46RKYnSV2MSNJ/lDzjCsa1i//VIYrIjPa+bBZk
76hRtg6VzKmifdN51L+FmL6tB6whqe3UfM8QTVRZ1DYbPNJi9dUtk2tVbyzzn60Q
KakIbYcOuMDWBylesW6nneX4lQsQdd3eRDcVT28qAvSBDbygBlaJS8EHPc7VL6xD
DGzKGuO62MB9jlShjK0IXULDytTl75qIVgKEIq0Ho2sVWq+xp65o93zybX4zp9B6
W0ADb/e7d+8uWjBMtTfWXNmRVyfGMZ/CwgDlNOANAPTsRP8rN15JAGaU8kFP6YkR
5XrIikFFyMwAr9OZ4lujqTxVs1pk3G6I3/Zu7/Yn9PpsaTQPGknc3mCTaHmNPfH3
XRxBkFcyS4+gmxshPkotBDygYF1cyf+SaSjfhlpwkdXH5snbWb0eEloK2xjUxin2
GPc9gTCZXTfII/yKhG9GK4e96muItO+mnjm4sGny4yWHSCtGnwYCcIOE/S2wQqd9
c2L7DoG/ykBGFGeGbY3m95jMX0XFX311hQ5yb/RDGTf9zqdCgDu2sktfE2Cgo9eu
zSlb7ZfauYd1RmOhnHV+WJNh0cU0Ux/yNRCSwdrtVKisVYa3GAoGzU+t7cdx5s+T
A01W/etr1GcFasoW6/lp2QT2nLKkPmqv6WDpYpFDrLYzCNjwh2GwACJbwXl8By8R
E5z04EvttewkrG9KRMOBPZhbbiuG8iB9Br/8HgRyDaKIBu9OGLE6Aaidgf1tlJrs
sVCaLtxVrVZ7FwxJ4B1nMuTuAJX8gH+g0T7Rh+LbtwTCs+r98MLAO9OlF/F45ck7
YkQkWY49N/73+s0G3y7hDNd0pHkI0rAXIN1v8gGLAmSXTptdqH4X8GHgn+OHvmMk
7Ifdj8F83e+1IDNZcTuTeo4D5NQsWU/RVCFVfV67rIvLkNCI7CZdK6IT+CWKypWk
v6mYNOHR5+rF4f0DudE4u3hUl+VTY6UKM5wP64artff9E4cBbHDfQ0sL0y7hl4t/
dX0TL1WXkqnTQMjS132sCT7aMlGk6eH54ynOA9O5xOtRM/hjfzFJysiv4k9wik9e
9Ge8tN8ej2R0Io5zk/S8Ek/mvy7m/gw9i9KMnMFY6EzQbCtWuXhL+m6N1eu+WQMc
Weu5jzyQqmp3VxwA8MDz2DtdMrJHcAI/rPbm+QEooU9VdmgcE1jM+ZQ0GDNwT/QB
t5ofMx/XMonHAa3EaSSvrAqHsgqinuUZDI+12HSwgv4iqZje26wqlxNYH7n7tryl
Tvoou7siApgXvWKXipQlZXAiLXijIms1uCNZ3yWuPnMhUChAs6lxnXRVp2uZ/9Ks
BCBGCWAq/A+nwlr37WfqLV6BtN+Ro3QF5XzqhaXqGqLJh3iaAzNHYWZ2ebsdUc4y
YtKeOevQW+MqDu5cdoZu7lN804g5NYdi7xZVWofzZLgTl7MSDTSq7WlmUJd4QmHP
8LD5WGPrKTMjP22JuaJ8T00iYwOeRwdgC6A8npX3dIPizI29t6BHGcaFzwSxp19j
6Wu4M4lzGoneEDdKfyLJ9tpXfhQ0h5teYJMagwfdBskwgWyZqSynvGkXNWJ813om
yPSJU+53om8jnbnDF2TjJQ2Hdx+d58O0PTGH5DzoM8YYECvi/8E6QeK7CQ70bbo1
sKSoZHWNKBRA8vEWSi0vN/l7KKjrlFZYGpFM0aWB2r1ZlMtqVkpzNoST3y/+xA3n
M5vv0mioG+5uPVqQ+k1fUMBGHld3bpimOjecrBNtJtg0VN4AaOuWhGlGnLSD59Q3
cvh8e+l1jX8Vx5EnrUjsFtG+eYVaVSQOauGyxsylj/OSaqT/tHO7vWbJ4cnD+OxR
4Tz7Cm7fmeQ+8RPi+Q9g5psnUFO8w3k6xPqj+RKz3F7n7M3TBwuxUu86POu47dgg
CeWzWLcjbuSc+4afXMgrTAdTX14Pizm3CsFeTdtLMQVtRRXUSRgNE6Y2m1PtWMZu
qPt4LRqSRwD9OvW3cWmStx/LjKozGfPQ81mKs/xmfHk3PjpIBXls4WSmNlKhaWDs
9VQXDVFJ9wA+dYC8w0cgu4gg7mw4dOfc3lgLR8Fbei7q6lg0uNKdcOv/1vkX5VEp
8ffBZ5EKQYQaU+Bps2Wd8N2DPUJXpBj1GE/gozy9PPzr2ffwZq02nPRICOMHpEBk
+ZT5w4w+2K7+vX+oCBcbVRN6I/NE6ZX6ZtrqBngDtYyfXIo4Zww2wsdBO0PEBgAm
otBoGRmjd9QiKprHU1pxu8zMFiXCfkkZstEmh3aBRvw8/C0jMXcK9q9woKXyndNZ
K097XinFKoQzzZYa7V2Lrf9bSuDdbr18YS0KAVFY8ZDztTe17j4c9Z2cRV52Dxio
NCFqfUTgAsBUnTJOHMpH1VeTp58eR6lSlQQeWmj6bh4KJjOXRURPzovkcwohOs1D
917aN8vSPVvmxbd1rJRWHPQNj516GCeenuXutBDjfD5mByczFBZE92Mob+KKYCzv
URICs8Sozg+e5ivLNSdJRiaJVw5cL0vpI0MC3hGxyTUYrZ5JkQfJJjyA//IbiMav
fhqL6oLMVxtnCTrTgNwCZUScaLc0roPs0+kZyNFhxnAwmHs6t8DHd6feP8amW78r
akudvBEvV1vRzVlOSRxsKi8M4xfU6H/YGs0Lh89ZN04M8/ChIIson5xlicVKJqHJ
icb++CNKMWr+2CpZopaPFVDxlcHbMudr12hLVGehZcIGlt7aUtcw7FAz25FZTuLd
YLHk9oEdfXyVIUGhrZlMjUgu/v2tjZisz0VD3JNwN86NaVyACtzOWGjNm2gfJLsU
IrRwNRXHsHyLswVUAM5VGNSnVXhr0poYKoN6f0wwQE9UCf0ETHdcnpwayst030JP
5EU6dGyVIwRw/WYRd5ye5FlJDq9szBXb1NGRmZ6Er2Ld2R/w7gCJ8SSAGU7HZTRC
YqSMy8RuSvth/Kk8ahomZSaKAbk2bIBTO40bYPMiDXSuFgyR3ypc4T2CtuGrvs0m
fYIPHOlBXIZOvaRJcyPYNLL6S2uhbEcdneYVuULBOXS3xlVo3d+eKNO8jVo3Tck6
cyXZ+rsqceAfZKO7FQegjdYum43q3qHt+qnz4/F993dLC5yJ6Q+wGQ3nQTYuDNss
E0VgX6HvwlSAjg+tj+bCu7eZj3F3bNtIbUU0OgzdKNzjjjWRnIEN1ent1DLLqvBo
QAlf3MnY6asxdOla415b3NT+uLxcGbhysCHNkTodGuVmHkD4qMpMPBq24S8Jkfd8
XL6TlkBQe/dTjoM2LFZ1QJFWii5QSu0X6CuSmn7B5Mg7G2k9Tr0G/QjYQXtGkeYG
L5vgvvULpKLzAuaMVIeYuCx7GfYMY1XoYd8azp3gwkLEkrkYLT9u5v47YgkZAdPP
H2XxeC1MRUNyx5Vo3lZxyrIjvXr67SEZp1BbDe43zgjS94fk1tT3n9/VeMoZuqvn
ayh2LezYZ/tck89cOej5ZgkSUmv0XB/6yVV+x5cNA6BQd0ZdCQsbPhPrsfFffpkG
n/XGW+ZqlkhDFQRgt/LagsFhrHoRirWB4ILwwqCgXBFJdcHFGFIcwz0PjhZ+Y8hi
Lbem7Jv3+6R9JCZLhJQQbjCn2KBRsv0frhn+67+9UV/xlltSfNcINJ0Ngy6xONWe
cY0N/BVKEX0Xu0rjzeQJQvn2ZdTqkab2lTIHHWxvHojzCD+fbQec3ZgyFcHTr4an
SYt27wRFQ+LLlTxzm+39znXGzblbzxf0DgsfbCHzRZAlncFPKHN3uiez7LMEnWBg
DBGsy/pctBlyotLJfTRHLVaj6cEZN+X8tAI79NnPOgI8eUPE1syN6FQ/kjIq5+U0
gpY7UJI4MGqAn/k463aMWtThiJ8QrsOLmNSTr/QtorQ1a8u4IRna6lccY/3jlM0+
fZ0LJcFhEdfzEFPNcb9D6La4BWYSNmTcVN4LXkOnGafLV8aidSeLDhYSTchGZsBT
d1bQhTHBacF1x0RgRFU84w+okzAVIyJttVz3SWaooySGVxwjTk92JvQW6JKKe9rO
+h5Dj8sWkvOrP9V6n7Mz/mgsYIDk0/QkLOQPdWOJn6rNcggjqx5YAuKsL567E52Q
dahRR9K9fyZItc2a7gbLHm3+PLqYTTbnq1GNwoQ6xA7LL0/jFwUZQqln0GfN7ujJ
5UC7ZG54/8+oxZ7erXVnH/nEfYJqcwgkXe2Gw4Gev6eYGhI7V/KCOvsT7ELW+pHW
jWHMdBOptFH6fTT3B+TstUF8NTglFCznnHytP4c+IsAN9DKcDuKDW5B5M9wtTZZT
W/MHG9OWN4lB44gJ9Y5MBoaSa5D1026HpoyTSAcljRdgYV/Gm5mShPwm/t/Dwbbj
yYEUU12X+X2xYIwzyWx9ExfHyYiIwi6PuF1xqwS79XIziWevpp2DEcQZoFVd4WVe
luXaID6cPBc+5xYHtnLS17smck4JsTeVwFS+vQX49LS8Jz1Nx/mYi7yofgaabV6K
du6rbi30K12StOefrEQeSRZgnkIopx1fx6cTfR/XArBkO1kYTlevBKw/BewfKvUu
FP0GQ1UjhM8lt+My4yKTDNuyKfZLXyrL9RCRP1V2H8MmiTcBQn155SGdaq2gEG0w
3EyThaL296TjD3Qmvlr1efGpeD0TZN3ko+X61FV8M+bjXT19eCW2Xxv+m/L3WS9/
k9//YuMpOwtuOngyQ/yJ1l7gA+ll0lvMrJDeaKcSJLPHinfapr/D5gqKpyBkrP2T
QkU74FoISesDZUFLIXbIUfCqaikW7Tk7ICujmsxaQE2DHADCuzk+ZfutkqMC/8pk
SoTvJPVasZ0tkqjrE0/u1tf76JEaiEy21APr819G2WNLbJQCBMVWrCqBHeCR4ISs
0LKFJPuuZoqoPFBzdJDV2pfSQ4jfcLrI6RiJGBi/GzaugprT7gF0x0LRCNMTtvbx
eiEfiILEf7dUedaDjmkXDUA+cPwAZuPnICtgvd6DYav4jEPZLqTOCUFXu5jhwfh2
YVSwtjHtZl9j97kolwH1MDwX4w3kMdRdudbFh0mWxpAyQCaDvlt7AsypjCwqWLpf
6u9vIOYcBWmKfDykhMHvSe/Kd1wiNhrhn895jCTVBmsyPRlTI3T+82RBGPjn1Fce
4To0DxBFMWpjPQZXwsIGVCkLhxRds9EvivoiR7KxxYyps+cjc+SKyWtY1Lp65uYR
HmYjfAfQW0e0veW7laOHc+TebogZfHoiQIUhc0nzq9mLB6UB+FpiIZSoSfHXCiCv
C39spjRmQRoAPsoefJ964JfHcU+02s9zJXzTX6xPRvLIJQ0UU20f+P2mzIsSQa8d
eXZrpU6ebfFd5BZZoxqNFPjVHkPZUvDSZAJYYKHCeKdaRbKdDoLAAZyQvUFnezbE
crkuPQRDI7RsQcA89cWsihI6vi8hhJEJBA5T4VtPY1xUOJ1R0bIgqJ7+xKVcrM9z
4XKzQ6kqKpXx6h7hpFeoEgxFuTXG69+s5McU4q5AGmHZZzD96zjE7icjoq0ulZlp
WDXpZeECKzWQwK0bbpzTRTnfr/OmjKhC+l43N7fdjxKtBvHYGv6TdU+mWNmMsZEV
aSdfAebmrqZ6TkStmFaqAovA0QgSwgKKDV2n0ATiK38oYZW3/Gd/a9bRYycjKalU
pXYtDPaJ9Y4RockQ2SDleG9qglXcpnvUjzxQ6sioKk5ORm29enrQ/ReOQLHFGoGl
s6eANlO8GAcD3GUxXvXAIvxxDIrEJjNNpv6dBDQPTCViZpPMsOWjRckJxzuHQ7oO
CDjqV+P0XT5kYbsFJnPrF7o1z9O75b63LcTv7zH707PHG0q0gWN2olD34pZf1Rjw
iYdTJeUKLj0OpYEY53ihsVanADR72sfWUNmGan+X6Ov+2ffT51unwdgzpkogVLUx
EVfNMawPUBWfcdTS4skmYXqsNDQh9m6IyawppyPHrgXXCX+Zl7CYAu+GtG7351DY
gsZ+1j1tBgP7PGlxSM6lZSGvlAXA+i/zJ6tUXU6V1KOj4EZOyebUdJZbxnLHtgT9
aTxK6Z4KeLD1nNn/3LimFQPPxLjOY6IMahg1vrNzZ/DQeHArhLB6LE94zz4xYFn3
MngI6J52Y31baGRjpC1L9xQ+hB1sk9MJ8kNNySdnTCyA3wQsiP2ObzlsoU9eiwVi
ncTL4gX4e3RGpohqOnVKQM8o6/KNKe8zRvPOWPCMZKwTuzyZtD08NA9MquP23cmi
fVtz9hje3C6YEnjMRtDZRNdhRLLpitbscG53bow97LnvzXa4/U9pScVuvAzX+oMb
3iSgfs4nPJTCG9Smq4EcAadbE9dsPZhfVMQHFEZFupXjhC9K4Lwe2jzaHBQ5AXH/
qGYbbeRnSyMP/DXwF2n9/4yEQH2+TfQtLX+9P7IBGnBG66lt0oXTxoYTKeYZ+w9n
G5FwdYoJ2UlNvg4M4CmMv/BFWdclFd+pRsDYHhgEjKtbDN4yTQoxzDmxb60y8efD
HsNBXeZqlnCt87DILfnxWmlvc0rajh1PC484X0x6Jd0g6eRe4cBU1VMHRc1mVxNn
9JZGsE8+AJW6Oj0dkEG6vBPVdmmeeGQhfMvaUt9tRMYP7JS1CUQLjYkHoFF++lY8
uJE5b2JIomVB9O6f/kIvLO912qYjvkymYSQu8bNNwwnaFxn2Gg2vzaj5VxRD9pnO
pGMBZ1eGh7R35ZW+xx+5Ej5yf59K8p3WHZN39eDUmYXtpNoAIXyXN+YDb9uyV3Gn
lQsRZRdQuj2kwDpD84ePnWhVTCqe5c1cxhxKD2paiO2TUOsM6jX6l7OHMhU0t4fp
Wg2jQSnokG1BMNq713nayHLVwgE64oH5qTGPX0LctIiD7WfEa9STfTOXoZi/qdIN
qfnNb3D5OV97MheYXHlyELhM7QN/xQnMO8fRldpJ2tN+ambKh+md0BOx4BN5x+KH
e8J8JTOEt6A718a2pMWvtSsAIGVoVYEW8xbkGn+BKw4zLm2cteEvyEIgeEVmTipS
rSD6Z3+HiE8NBMbyVhy1AwkTjwCcGm46Ql9NyDbxCMn0kvrJYK1KmJb1G7TK0cw1
IF4fN6SggdyuxyajruVxLfHTZ80Cf7Z8Q1PIsXKOUm0IFMrX0RNwCHlsDcFewHEy
htHvxR0Vv5GPFCqs0iD+b7hNKHQVX7zUxWA0sjokd4uQrzt9KntN6uBoecd9xZyg
3Kw4Lk6hHhuSHGoO27vYohEXaRZdERPlT3Wh+dMA/uU+qYaUBTEJYgKoGkQkTVdw
ASV8gNhajWpu0+foYqo+wpA4PNjF3Lo/G8n1vib1nio629BG/cEOosC9O7TqI2U4
zDPFiVgSTRg5bN4wC/xVnGViGlz3nqkQ9Wg2w+ZkJV4tU4M36ArAM3L5QcHzyDye
5QpVbmN8pzsTiuCgum1OmsCuOAd8X57GznPsiQc4K2kl/5pY5jLew+5lu7+nh9kD
O84oQD1OtYlTyItrco21VTsHdRYkKHl4g8JInl6AWGpZxFzNI+grHBPJCTZDRaMi
2Yv8BnlPsK9V5cMzoj8/+KuGAkuD5J+wsaZJIINP5yurJcmAQpDqaLtLziDXuUrj
nXkp6W7ZJdJm+OaCcxR2GqzPIY4JL6WR56ojYjU0LCC4jeWGD1XVI6nE1xhMYPg8
BS2DxEBA6QXiQqpPk61spFWQQq38mhmCrYUxOaHzvV+GnLqfkkLTCsaysHdqpKa3
t/yfDjG2zYH0XyYVf/twZ5HD+rURds0vdd8ioXEt4bQpEvEiez0b/hWUFn1NSaqw
EA0uPYfEtbk4Qwp1Y1oSVIaP0TcdPxJnni2kI54/EEeJyMgOoJVv6kB1w1WpRE9d
5PqAdULgO0RyfjMGjuy81h9t4ZKPwfxm3hfVZmuT/WqLViOttrEr/uvSaSJjh4fX
lboOPzfEZkYcb7jY4uE7OooXlD9dRiEeF61tsbkopzlYc/id1xCbo+0VUtu3ugQi
h7xB59eSE3UxFXPJ2X30t4oQgOMQm4DB5IVb4mNHIGkEdRTd8pBsfz+u+Hd5oFga
L9mZinhfvqfsserXI6ddc/yhLQJnpxEW/qaYwJ1n2MRJekB66GTfPcWQ+oN0r4VC
tvxAx5t5X8O03BtO4NAH7jkz1nDBLvzwZv88ZE83d6P+tOfrSPoNWRn2XBCxE7ir
ZN1XAYC7rZmKSZrz++ER+t+VSak/XHxdV0Cc9Jml9hGt9bbTJjX1VeUEXWUyoGME
tE6OlDzpcT9eAx6xB9N4JEu0IEY2ZL+do4tzCpLmzra6XSwbNhmw8qOMWdmm0l4G
qYanIITgMXh/ILXZOJ4tDgdKGQZgCHjC0kBhXjPlov0qIlLtFAWUgD3Vn1HoFnHE
XADwLkwKADJTfX9cB3Vnrxuc9j0/9HTsjlfm5wLqrq/TCwxyx1kkPIEl9jym9C+v
XeQKl/UPaLS38f91JM5R2JZ9VI9dxKPdKjeL3HCBQuVnt1GIl0xyhajYOgLi2FCC
L/NfFsSYUINBNSb2KpeVYmQnObsorn4eHO4ozI/poXfXQbzRWX1WcNCh6CtYKkiN
5CiuVgybcy7wdKYVP4igB8DOhlf7Wb4jZJeJqD+FCX4zQJ4SdiLep6sv/X7qgdoi
k00ffVly3/V7mxuO0PJGTlxECtCLgB1+xzmXU7YRJQ3eu1XkoMh3XW8qZosC9QvH
bgHwIdcEpOv1ZXRl+pDa0p1weveNyI0Xi2OZDQjAI624TBk/PMWyTBwDxZNwhLEu
AlpcBzVmmZ5Ea9+IE6js5LnpjJPoOhKzfWkq7TDfuEVQq/BsJC4ngSpQiM0/DM8Q
iQg4cGsac8gtlZ0wZ+RjX2QHhnaSjFGm2Dc1vn0CKEa4ApMhyT5gY+pTbhPgY5Sy
a9jQWNOCe2j3KulUgDA1aNvMNIQCB/xPPcI+s3nowlwz9A/ZhBk8olLAI1pjo0lN
n7QQOVsCTDVj+B7RNL61EOojDO8NE1dCEZV4BJlohQrtzF1u/RNQZeRx85CfPOzU
j6YCIntQTW5TWaOAS80eKBFoikyGUmtcH5JrmJTyJKdPNwvUngJV9lLEfk/s0nSa
igVa9wZMr8ItbHeKiIturSbXH4CJ08tfwju08D2rIo4TaHY80I7rSKZQrA5hZrv7
GdATNxmB3f2YKfdjAXFT63n0wApdBaaMZ1M3u205Ukw3FU71+2BzHFkV4aI2O6pl
H1w74LT/XVNZNqvgl5lmtWYLNOAjC3aVqsGjVtLkP/3IhIBExwDP7tPetSwOq1vZ
0yZB63UT1mETJptA/OP2HvQstYX5ZFB/LU5RvKCsO27lEhQI33GdOpq/8fiJyzLJ
aAnxFQZkVndv7dQb9Xw8cPmPtdrJymAgvbf9/eyHwOZb+irJHzGkmMePTnX+S6SH
qC/JEHc2/xJm7urw1fIMhg8aMqGkNuo+oNy4EU/xaP7X6G9woPWsVii1l21TFTaN
79CJ0TbXBvw2+NilEOkL20f5UY0CiLvlAkKyI0Xwnw7vBJ4xj7BiYKqtkYb0tjA+
gkCRO3HKJTEZM5KW3OdVi5r6yJf3TIX5/vpDyDGDSCi1n1pLB42ZJNdxrtN+L+c1
jBOzMqmSmxl9hJVCsWGRDrdx/hMy3PmKMVbjmU+iN9AQagT7WKY5++8kU0Cd0ncc
mRCmFG/TTz74OBcKlhloxKKXR6sovIOtgPUmmjfJMZVAhSvTeDWVoJrmrkynI4t4
FGAyr23iiNcplksh35TUTZQMioDkSxV9O/BAW6y9OTfWPdqHCDQWQpUNN2BzO7o9
2+uMlGMQY4qc1+0GRFPxXi9EENn0gS3w3hOWRVJDB9u8imwTWp1dLpv/7VQqeXd/
CMuIpl4Lv3nR97ol+jQ1ab2Zf9tCRHhP6hjFbFCvjkVH/y5U+AYeruWlivcn/7R5
8rWVZaHW7ADM2WKI8FBVu+M8NZFt3lItNfmcZL/jH+jQHJKXx8f74vDXTprZOm+g
7Bv21WlFehs9dhh9BM6I/e290e3adsz7wy1c9sWKn/m8jQaM2Ka+YLze+Ymrusgp
FGbFPl01ljaiHr8EF1VjDZ5M99RMflOf/4mpz4adSOCZ5WEqCRQUVSw/3K+nGj+d
7ZWIIGoG3/bD9byOZsHzOxNubTvHJWdHfp6OHekwbspyJnqAwNmvErA97fYrFxB9
FFhRfw+bsEdLfaNWGQ2SyU4wFwBXbJYLf16omjQIR5zi1LN0C1TtfCI4hQEty+RC
GRRxob6RgkpBrAgJ5e024X1Wg8ZKPbHzlVk5JgZfjaIy3AuFnukjwPtaj1UbGbhd
19ui58oOTB+2wqpy4h6oZkYafX7MVdPkRV69SgZMIxmXBk3tkIrTZbELJOLGPXEe
nsugWf+hmiW6sSsBW6zInfE2zjdE4Xmn/liOl6Y7LeCA0QyoACdH+k4Cg7BdQHg/
F7KnskzZuFHL0KASTnWzYYRtZAkrYWcvEXp6Ekk2MAXpHBd9vypuZmDxrQryBuDb
bYC3nRZvlSoNn1HAKxTJNAYjAd6tf5YF2+5stuEg/XAqclzQprxQCu2WTr6ZvVzw
9clj0QSqk6Z5liqayfmNrkZe+ZPv62y2Tc1A+kO5wtLGycWQE3/TEvmDLKOesU2U
VaW2tRjVFO+aock76BRVruZZcJRWI244JB1nbkblw05zieaYVpU00ZzUoZ/PHTO7
8+VBYXHpJbXqT9dK2GNfZXvFgrBEXEyUlTBG6W7z1XIJyMkTh5Yp7DcGQY1Nd2Yd
WhVImov+PrNVvTwoVUo0ACTdtP285/1JCDYTTXSQOt4anydEr2yDoYWphx+myY+c
Te1+CV7ZMyEhI6HNs1xR2x3eyXBTZ/Uo9pqg8D3OGZyl+wwoi5bPy2Cek1r1MUD+
zzORXAFODptJtEDMPCsV5QWuWgro8VeK0uGgr7AAjDZRBNlJPxRMXlVASJeaRhvV
vSGcc62MFNxf+vYxZN0ZYnUvVpr81rVKCjha7pXI0rKXTjTNgc+p7EbP4p+3jyRb
dFB7RxNMLLdg2HL1xevgL9hbq791BRo2Z/CzrawhxJ4fYPIeKWG0h2BwMwR7+3gE
Y5sBXK9onRjPk7Z3W0+wSfPljnUNLGBhVD2cSM+iBHGJqf9+cgVGr/YkXOzPfVSU
RESVq1/zwfDijlugMbZS4/LNoZMf/7ibFo5hW36xh+GIuIrqUx0nObByF13S94kw
9GMXf8XhvC/wMxfI+7FWZFl5hzzew8T+uRxMtYvGxjEbEqUuA/xFZwHnQRqYdBtc
WuNnqwfgnbWVGAkn1TUqDfo4Jucwzt3LFavfVS3jjOR0LHxV5wS8N4gXPBxauRAY
aO3ySxvt0s5FPw1SCq12PQOMXB6dwShGkQh/nNF/zb83JHutrr4uFE2iYuvHg5Cm
XUVqTvjonDhweZNO4VU8FtnyQd0cswoOyy1W/PaqIKF/UYyo2A+QDOaGRw/MOGU/
rhhdvpgyUx0Ta5ZgFOwX6LGkxCcbCDGc+za0V2u0F6QFNA+CXBjxALSLrXjksCnT
Uv2/Au9q98Q8do05g3Q4YdmZj8TxcKb/8iiisnTImXxF4/wfMKOJovzFVzbx5Nw9
RFQo9c6BmxwTUX56KwSFohaYAyVI9kDQM0R85MyRFG9UI6u5SvIxPe1jq+wnX4ef
32X6D2hY+OStyWkNcAOsvxij7EZcHhi6DtViYFw19jJBee+zAW2OOTD4PHIfnXoC
E0Rz7Rgo0k3vk+7nGKUvWz9kwFUNah3pQMIFzmUThAHFHUWh89+kmbR317uiFTWy
g2w9YGt3An5BRVdYxflZ6WMY0qW3MT2EX1+bR/vnqSKstnJGP36+z6IX+LYkt6hJ
yTsEgmEiq0FLhSdebK5zJH7FFvD70CVpscpCCs6fn+rlcz3AigHCWdXqddkPavtA
7JCKI6aFSCumDp2DNNSVtUx1+lYEQCgw0ylWyqlMSfVOFDc841AlP/uFVaQu+VBA
kM26jHWi51ZSXPKh3i/tD1TZRqXZyrz6uIBgs/e/yZn534P1Nz1EjoWCKZ0toV9a
NTQOj85jiq1p4CWkhiY0rwc5KpgDD1bIAStPVI+OCnNhdQGwiBjG7jPcVTTUUtxv
ItHkL0yC2a4oW1MG/3SelfasEhF8I8fjaJal7UI4Rz9/nNIYTwF1DjdxkD/m+vIr
cLwuVFIK0SWF8vgQC6LFr4E/TNzQa7uFQXkPT8y7g/CYwW64/zJpSX9jzjsp+M4h
oxa8vpFUDehjnJW7ca4bQ6EKBUg9RkeSZPrhcIODnv2KmCr5gEG0rN0WKZIp8adt
YWaWQ90xtWQhE/+Ky9TCV7CjjjYm2EfTUGZTsycevr7fX0Umlimve3Vs+Jb3EZRS
nJP4UCW1NwI3kQ6ZN+LdjjX7Nnjn/90wIx6qGns8Yv6HoKHg5GTZjfJOpCxdxjoU
JQ22SrfvhGWH8qNURlMd2uPBN2ekigPReegIIrHpum7yKhPwfF9Jjtmd/PEYNdgV
qOzcgpuisqa30WNjFXMZ1xhSrU8hhCLNc+hcoAVjntlKWTZf2tDavGyAw4QDmOH5
epmi3nWZPbxMcI8oQstxLhpr0caxzE+P1JHfveejKvIIzm2HncoCKWiilNmRtn02
bDNshBdc1MQV8tAuquaOR/8unhZXMhfScomswwZg4+Iwq8ICAogNeIqE8lloaS+R
f101NGMMduOfjRwfTrjydMZZXhddV1jvfC9yoFMYqCDYT4nrgoj60ELDTZqg4kLJ
jKR91wVse3q9xjUjwH6dPPU9//DPkX2KkRWlv0oSKaJHpuCsbDTboi3/6GOHvj4S
8aOSflMm2Mi+LDYUiW7MLc6DH9nwDivvWXQk08fJDTUKAfqAt8stwAalbtIkfOTl
EuP5EKtJtpZr/EPNU9+pgxSaFiMr+RPF7GujsQd0TXH9UXelc9PyYSyxX06tFOFc
6g2EkMXoZqnqZs/bFpm7KjPvaNZ1ZuFtjqow7Vn30j1MTJjEcAxUGPOWLSZAkusT
MtKHHdBKqX7xbHmXwZw8p97NVLata+4nPGuSP8Cgz5tyraHS150Y9kQPRutlQ3Lh
BjVPy2mby6GwKgtypaQjoI9MJSfXUAVB+QX3zE8junqEEW/KSoZbUp/zqnixaswA
vI289birh2umduOza12++9lUm3JLUfMtkH8BDMT5mDtPyhGI0va8yvpP/ROMLoUv
rl+0QDBg/6vDtXFlaBcA9ldDZhvLc/7fNOMwKVntMlastojjsteM4TvH166PxUtz
JR/pwD70pCa9fJvZ6ad1mSmnRBUV062Fdursl0RtmvadK6xWhbS5Ku5zblVqHHGy
lgzQtKuY6RlAVPj+nFFXKlZmhXRCuZRoLfiz7DUIwZXV9H6/NMHtVZD63Mn1KVAg
gFotreqH0UoqdX+1SlErCHpqB8QNP5ta4uezteIers7lTl34R1PGMP71bk7koUKp
E5Xwr+HNGRYJCGI5OMAMFSBk7en1RqjWM5EteC/HiPNLLDBrkZEIAGoQzE+do60z
UL9+Xozgclwh+97Jz9VR+xnkOznpn8XgkZPhSwhvXBlu//tNom2Ti6BxXDsDeYPs
G9A9cHufzCaZYJfkYmVoFGVXXhAENpbq5Iv8U2SsIhx2pRAb1S0uq4VXbPvBuHes
ChVZbVllx+4pVEsZyEFA6EmiBBcUT5RAsSHXn7JY4PRIdiT4BZJuxys5tJ725vsT
maYbXSzzHrMygurMZKLwIUUXJsS7+1g83hB8Z/3Pmgph0Pu6Vuf6tjZ1tSIBOeSK
kziGjSbJ+i4bDjXziOZokooW6Md2dcXPJvQG0nROeb7snfjxSltFAD2rXeQ40mwK
gH9K+siUGl+lyNCMsZ9McLj6qdt6VgIAp5/OmzAc/pMRq8lnx+ytCaD1ZAr+rmdT
02U04MqhFHrvqNXy/Ch79Jc065cVtoCyg7ZtUwPfqcL5BINCIUZGXC5HUeqbqM5S
5yTeoK3aIA4l8cwIh6PAn7vtKT5r8nfGuXG48ZtVlo88ZlQG3jOEsXb4ZzWayOU1
jTNHJhOT/tWeixviEh2zzAnBCATxLDPOrn9Xu0TlxuSS2vqiQi4F2bJtXKasjLLr
xK4xtV6l+3X3boqFo5ImR4pkipHmiFYFuceHp4aZrhTF26HbQ0TuOYg857bi7vsP
wmKBqMQvFPf5Sqa7OWmBfVhnmrA9xiM/RQV05s0+hlmfSGH86lR91hbhEIDMuQxW
pWEJOQpDK9WR0WunSTZ9rmijrLaey09NNu68zh0Oz7Wboj5HrST4BVjarDWUmTqs
uTSKXiDPJK7MG2QxnFSWs+iVrKbOoZ7haFdX3T8xCnM+xbJ8ite6ZB6CPiEnf/1M
2NqUE7TmZRQAnHQZuX4jQRkB3GbC2QrOiI3egzPtQcue4RBBu2iMspmsWxGHQ4t9
HNsoMq2/dQFFoMz86XcOSljh40u343N8yDcGFhziUFv815dbHmMxET1wpUf4n9om
xoWBRvUBqrQodzBBW32LZ8d+LjHyaM8O3DdZnYNWNvvd3tm8j7QjU1jXCLVk2ZKo
xxWyFeLCDsZc+sAvl0T5X6ON452UZ9OkzfrfOEUM2q1wdSomIQ9A6s3rzUBS0DKI
0Z0zgD8nVPbbvIjGIbByqPWh1PE24N78UISbxDh1YWQrwHdDXBFp84myiUe++1rj
NHTYum26uNageQM+mNeSI5cQb9eOV7gVRqkaZ7zfxRmu4OudiZGU4EMJEv3Ief7k
bazfL5e8apm3yMYZEVpJ1lhBtrpFhwoKKDUaJj+5WkMVCuvWpX9DlHMiWusAVQXS
mT0oFvVoBy+5qGEFe0mpJ/cPl55Sa2kgT1m+pXb02Y9f15pft2aUNAr17BG/j4Rz
J6+B3zlxFkOmLN7Qu22Lt8P/fylnMQH0pgqyJHWl3aNYmuPUC06N6Oy1OB1FichB
9zMPpw8eynF0eDTU1032HSvlgznoFP1qfp8E6jsi0u+8DNMBojekxKKTvFRSMiKG
yBYgyAD/qI6IfNzR+DZb2aK+oyiHyazNDpLqV2DczGWOrF8YspJV1a31LpCWXiO8
Rq8uXZzsuAzGQ6jk2yq4MqXHnTAIP2rfmD8vFkjg/rL4tYd+ibNZLU4iMeYojM5D
ZdYAR+uLqk8/i80nw5CQo5AO7/nadQOdsEDGjzpjvCYifwJZgvdZjRtFJXRLu+tc
+zeNQwcY2U6EEfsY7jwELexqOQX9ZK4f66diz1G13+rXlwexUChudU1/Rvoczoxa
PO6lcSY5qOddvNJaXOzylSymy8IZiu8LkhPGl83DvBIld4lJGmGHzHeT7GIUe8Mi
HqwcmwmeztDBIkdvo2X1vR0bCv1oEb4ATY1StMSiQB7Hhii3SbDyz/XE85lXzGgV
s9VFg9XEOubBuaPnKVaoOEDqqZeD2mo9ESAZsNf5BDPuYwm7ty2p1eBaBnuhb7dH
Q/pLaetDxeOprmr9Eye0Eev+qETMPt4AHC3cEsTXC7QANioKR97EndY/8N918m2k
vrzO8BLbHWzqyqeZg1XagaM0xhaIeBNHKZefpUke2KUWXNOAVPI1riv3E3NnBYiM
BCtoVpPVo6dMbR9BVxCTWP/ORu15tvjQaxGDD0DK2+J2LUgQ7uDvv9loL2rpMDWk
sot/My7Fe4yQ6vmMvS4IbmDjo1kjXleLoV+l/DA69vNzI4owF1N+0kvxkbPK98n2
EUBLcIRhoToe+ZypZ2Rcx1j+Y1urjm+l6UGWwgLmF3fNZArDi4BOc12ZZMLUVIDX
x/c1Jrf+OZ39GJ1tUXvKH9Uzo7r/Hr1YWaKyUG43x5VL5vO3todrLaLGfDB3fQVW
ODR0hPT1FrrRlrli96ohTpk+S4jmSfeBb9zBWWJWLacooUOgo1jT5z2UG6CiIH/s
Asm7SVYm2/SPiVg9E/g+jd5k44BihO1JrcS8SQBBL1a3nAxMvdmAPmxeGdxuTQTO
Zr6csHNXJjSgxOMvDDDfXexh/8zaxVpgLawGGPjb2WC0mjPdRu3NzKJHXlzrOee1
hAPPcOA0AtQ330/FhpIdqff+qPZWWxjbQpV5lFoBl+/slhsTIMqVrxPJLUkuYTn9
7FiopZVCNkW3bxqetorJ/M+YQsZRTRe7xyk0uGEukkFVPx2JgMhsV1k/XC5V5kPq
wRgS8yZpErCvvOhcws3QDXAtzP9vMDLwMOIbk7J+W1faxcfomHDZCLbucfRnaGEZ
0/8Pa84+sgOPs+wQL2A3P/NB3yNRSGiXzf2LXo7FCKjkB8qqCFlieUaW5hrDtygg
MXGu/EcjA0+XIvAag8/sV4u9WFfD1uQSTK0TEczHGlkYvwyzUfUfyTLYf6v/wHia
Znescwwte8UUcvSvW9PTIIGSruFNfDiiyGCwFA3syXuklO84lDORoBk1xNOC259+
7E9NC4wfP/DVQG27iSawNI1xitMBePs0hKUyV97rJxDyfkQgKW1KJDjqzpw6GpIX
x6YiHCWj+qxBhRuPLjurOMHR4yhGTqwMScn6q2Z+Lokk+2z4EilHPnREf04KRf/W
EVy1Wwyhu4CamQufZ7zUsdQpMAa0Wde+OeCGXBGrUNpa78o/trPa1r9BTxLdSqDz
kd9vWYNyzC6CHgRXt9S7vT1WE5QPs/CmmpSkJzah+896j94N3NgqUw5pIMKPZ+ZP
ZD8I3YL7QQBjgMVEPu7SEGhVLjLiwqkGJ67gqhGgm/vYCAgN2wL8zBC+3WFX/ATo
jdLynj2quQGuWS3YnaxlEWvysArPjxbv5rLwqOY3jG9hGXbeoZmBZXuJng+uPDeW
1vjunmRWnb7etce4TSadEB+hYVDhBbMn30N0VGXVCYE2aAtXPc3BW0LQrfFxb24t
Lfy156POqGMfuEPotx2/rxmzq1k+aBJhwOMzeIXjpwTzn0kRDV10cbVZtUgzJ0N2
N1rI1UgSG5PCvFXDu89LI5tQhFr0krsGN1eUxO59h0JYuUUulRUL7nsZS/meRT20
vR9DP8F0z0dILuM8oHfbYxqzuNS5vZYCqrel0+rsXcioKb6WQ0H6vo2U6/nvIMBX
FvWSX8QUDCvUDg56OB2RZgBYUjh+60gKj6ZBUGoiGetk1z/pU8t8kN9YMpReOX8L
q10/E5BY0GRXeP/R9IXJCfNf5i1CKphi4O0oEZ1cNkC/N1cNNH0E/J7zlL862Wsp
mwdMAFZvbjtIG7fUUvDKDEcF4lK/M0xoideQn+souoRNRJ5/Rbys0ZrQYx5tuA3R
5uGbG3tNxsoOqienFcEYbnmBNm7lset+UetN9bvJttBiS4cDdLbVKgQEgsKJaFbP
h2/CRIZqvKnrbM0h7SKkHj7Sbitz+0CgUode9U9TOhUtoRYDbyCPDPLtEOVkakTm
exVbnEdbAZJYFXmVjmtA/Z/MFxX6E/5Sn5ZY0RBT5YbPz1WeeTZLEFNJ312EUYo7
CSgw4OOVgWsGYPKEzBXijJa1Q4oTMCnP2LlDRzZ6UQkvhXXN545+mJfnZ2aQ7jiI
wDAveBePqaDkLyoHER6QrRh/Tp8Rn06Y+wDXliYAJG6VZNEq0o5ZQKyr+xmbLlTw
4CkUjVRfT8an4uFoAw+nfLHcV9m9YDjtfClUkJKw7XcmnV00kSnoUHJUjQlfWGPD
RhyNN7qOfUbHgG9O2o2Q3g66ifocl/qBkeIgTSBbrcMf2ecemZfxO/z/LMLcngMz
zmaJ9nYVyjraNO8JD/w0q0EhCFUN4nL+rYKv4nKdPAGlE9n1aUNZ90G1kyuKzPp+
RGgvNZuShRtOxxbU0Nw7GiGA9k9SkiLJXSKMsl/bRNEvP8giJGzHHkbS+shMjsA7
1bJVHYpVU1JGhspXgdBxAd24t014q7YioXmWqgU7+36/mcOH856ITLaSW16dEMfV
ZHKZnfWyYqTLCj2OeJ8CMC/rwVd0oThv4m13nntaKDwDm4c50vkPPX7Pw7wDw2qH
Jn67q1bmsNV2HxbEOyCbgo7n9inHHgKEbqgEJmbZDGlOhP+6L06LohUc+jEhxKyl
UqQZ0TECwO+gYd9gjB8Ba/RWK+7zHfjIeWfveM2jpNLKgMMxUpk4MbqaQm8uUzC4
gtgHShgTaTiBI5a4CNOEjpsOcRKFs2uU+Yx8TNRRUv71D8XAHHsYvBqAgnweAqzB
gralt+xhPko7AihXcLblfzDmnOCsUvEOgxiW2Br2HdKBIop9fuRbjNSPR9zRXS/K
DRYTbLdrR7y6ppwb1hUsjtGtmc/sTxDZi1WhUgvXbs9b4lYYxQ74/120C81Ts60R
aHGlkK4IR+SMnwAMuO0NPU6bMNo7YhYjH31Js6fQ8GFLUOkypKgx6I0jeWul2xIo
UIq4Z8IYfJT+nPlU4s0tTs6sh07YkVcnWYgef3JHnCsRV/obyCxpHxd0ZCaN5Y4D
HbbXXHgxi3d0vzJyelJ3LJ24BgJP21sAWxgKRqjqecpGQYUKhhiArtn6MYurdSXp
pRNsbwkevn/z0A/RGNPH/6fdquMy6bi+zbr+M/xCh7HqE0N/1bT2meGaSY8SRIdc
QjAc2pnny9UukY+abGHqeyzR5AuztJGcZkLet74q/xHdtJTfS5Z6J03KgZOGSlHD
5TXI75PsjjMJi9qmMcCLSxiK5QC46Z3+kBFbePTLMC7gIJT3cqF7pIkSb7XfqSJP
t18dECGnwQUZxj4y98AtzTZIoUtHNryJZsvLn/jWorFS1dUhgfE6CD83TR8nZB1X
HEoQneb6vKli1r6aWsAqujrLkGZ7GH//Kg4K9tDh1CziV2LtpOqTte/EoqMpzshL
iwtWwJGCaKavM+nTkbAgpSh4SSlQtikkr64Av8D4hVQw843q/2R/G16wQ06cq0Tk
H6ZADgKZg/1YRtUz1+szfeaBXKPDQ6BwPrKRCUVsKYRS5HF6j0dXUZ9T63mHfvl8
NMyfqtJ2eom0V98VeEhO3gfgUp50LeHDzDZnKuQtLoRjFdmfeMQAiZbwG+MxHYJ/
La/qZup4qIW9wLDOUrnFyr9qe3ighrdkq01DQIVEcAbjJzckgoSu6VMQFvSaZiEk
XtWZZLc+wKj2pwQs8DXMRLTeqlh5DTaUb+bMU+uKmGf2cOV96B6ihFIRqPGwsrB+
2PA1/HrMHHaY+G/Ec8KsdGuuFcGtc0EtSBk08dCsSSmX2Nq407navmevR24xF/o8
XqfWpDvIviz2PxSyQyBmE65OL4ERHCgSv/RO60Af0mFBu8E1BWPilgdZFunz0mKe
XOxZpYdFzureCl9iZyFyYtTzkP/m6n9f/q09s85IqD6bCNciycf3wMMx1h9ku7Sr
s651I9fUcbqycTgSbw4Mq0N/ZOsXkgcfwUxAfjbVvGEcN3Lwlvc8A4tk8cOM/ygh
dSmYoFr+iUOTJwKwkyfSUBZllEPBTUaKZGxkCqh6V3V9+WopIr8i5u5Axh9mMmjq
gPV6xzK8kOuFOI0btar8Dd8ZLNzUQiF7aAfC9+1QYgjSR2MyRQRi+5HyCaFHIgpE
S4zZKJ6mi5YRU1s6ySCkC3qrQ15P84UsgshcHfr+KAjhIlKWxPmTwscAOV3aV82f
osqrSK0sQbE2T9zH8wGclrf3PPOUxEmBivj+82eruRw/hqg6npIKhrj9ZhHj6MWC
jshi3jJmYw6lAqHfm20aH7W0uhGFiETNWTFIwvHSfDfJLUKEmEAD6h3u0V5+Jniq
5CP+PYwpzE3ADtUVEG5dewSjYNhBkXYK74WecSPkAvdNt2FqX6HE7cmYVaP6zbO7
+RVen5+9485jvcyIfqGmjuGslgAsQLBPpVfx74GY12CJZ+r7TRFssKQnbCVoSzeG
aBmbeAro6uZ/7b2IJUI5myx0fUG/gtd5TkGgkNkva/CWVKCWGlbBjLIJT/NrgZJh
Yk+/1jD2apCoTKOFxu3D2oMS1YqOnQEBt3XISwyzRsw8cUaWULLl156koXQUVfl/
Vr+bB58+KND3/vNTGwjezUZrODnn7VYyxRg67d/TUdvI2o8HWFrP15kkgmpj25Zx
DCIxoMpY+TzCVoETRLOQ2MvAOzNNEPyJ17Eur41sLGKqLMSnZWlZ8K9zwMwemdHF
gSceGhvjizmN4XwtRMBnY8xHmYiJoD7tWDH3zsfjQ2bw1V4EzgTBx5QEuf3OZBZi
OfjgBsFgXN16gpzf6r424CPO285clFaQRevO4HQnSeHNpqty+kzGSW22NJm0/LEQ
tOyv6pFnpcYZW/kADkB5MTjid9UjXsvCxtGbnHE7IN1Q1ttAhhW43JpoaYC6RGIe
1wKTgfjZVueXFqJC7z8Rul0gIGw42maZibz8iTEdxbaI1/3yKBE9C6+phVW6POl4
JWLLTeT8PPBPHX4w0ESbveifXI6FICcBTIkEbjUgw+Lp1j3R8NHzu93kH7igI3gC
s2JyxtH0UVF/X1lewHp/x9LZMbTdGL6v+bJP3kNHbSMqnbAOmDq0cflcf6oGoG01
7arKmczAuusOWRGJmgtph5kmoXRS8aaz57r6l1LdQS9Msy0p30X37Dmb8vCtfNkq
UDl2IlhutZhNib2mzapDUVYYT1XSIF/uylDqsSUSnFl7nEvfETPSdl0g++r6Pf2i
EQV/U1WtQq4fdOLCWw4EITdob/s+qQqZYguPGGQsEaTplqDSvotzFcL++Dy5Z1CM
OJYE5F1u1RJRJWULbh8Bzywqrr51MxIytk+n2s8N4icSzKF1NXpIYg8yPNoMlpDA
lGtvJTg2f13BcOy5QLrekDOQ2zbsvH5o6i4ySctDRHlHT9clxaNOeeVN6/9hudHq
hnhNQWXk0MZlF8c6krK4Blfp+ldeno2v5cp22onp8QFeHWtQCckhWzQTOjlAT2Ka
EE2aD50Dgy5TAuGxiOSqCdEeS0OQOufBTfkQjcEhH5NmlqTZ6rwfsol532+bJqiT
FjyDDM7iXayPEahpNKaG/L4JJK9gLkL8QAwQuXJNifBrQ/czZI1bDi4MoBsHMcbB
WSKmlEUuuZZ4/ry3jDbfMvqg+P7FUlahyXmYYNr++2LLcOSlEgd0ONqAcEAhX2e3
Wqi1ZC2R/HjSIM6y0byzamK2ZMH1sSWiEIecC4D36DIreCpQvelhvI+aijCnR1ue
eHWKq01DuNWgSCwFwv5zS20UAq8y/66XpUrO9UeygdRkQCXtl8Nf/nAISOzwP0hq
UxPUDYbLoyBATuS6itwYlAG6KBT3WzwsYzscKULG15bt8zHjGaHq7Wy6y3jpag+3
XpUbYX33/XuhdPfp/lIidgSHwXeYPSEbkHMioTh4t+6M7aoZMETWL4zvh8vc8m6Z
JKQmq7G7Ss6aHJtffQsozNxONnG6m03KRk4hb+Txl1gZYgl+I06QgO0Q9CUbsaP3
LvjqFmrz1j1T4n1ZgzsRn/f6nlYE42rLnq+vnt2EW98hJYir2A8ecA39qOfQ08NH
/qDC6y/wf7qA7MasZUy8yEqPybGsLY8E+czh4E5pVuDD6aROaylL//yaqfVCP/+S
Fq40eZX9hkZSup4L6GPlfekiXVUHK6i5Sfq68ri2+dEzsKV1Xh6k7GD2UQ83GrrA
PkANdHte2116Uu1ZvMK+DcYN4twr3zZbsPN9RtNEmhmIgCHa5xyuxQt435sAKTFe
8BOCFMdC/wRed6Fa8/dlkjLHVZ1abMY85ZKzxfYzFSezJgLZ3bEyanG7UpAoaeiF
cZ3b/c+72xmcwzO441rkqJ6WOSStpM31oYrZHNp1MrQ9vOi+BH+yGYmb/lMyT3oY
gSOqu08Ln4TMO5or+xLCTNqWuN6sP2gMrh1KO3i+Ku2bMH18uSugyycEy8MlZ/t1
mp3Ox9rs/VAStUu2sJXy2Vnxx54rjZF4uBmyIfL7zBUPPM85Wff870rxX8UdnaoK
qmzWRsm9FMaGiOUTwW0/Ip8AiJ5xpLgtaqinfdv9AApxUVGeG5VnTIe7FyjnV26O
V0jvTRe06XMgpl8dDJ3f2u/8t9kW+3kfhuPRDWZXyyjlDi+9/DzFPpoXONlkzpky
0AlgJSqRwyOHOxphlyTh1XYHwe8alazFrF/P66SZPSivs5amJ/rx6XYtDJHu8387
RdpUrR/ixXTWdlw05TOBZ3YomGZe+Qmlg7Q/wWG86FmchehkTnGV9LaexezN2SOc
FTkGwB1iLUpX4ha7gf/DzzrNiId19fax+/D4GdcQAqdMvWtzFrzAcJHSpLxfntCD
lO+Pn6KzHI+rPt3nWd7P6Ln8Py/fAHGD3na5zGD5ukzRS//oslbKFlLkiY77Qa3l
Sx9gkUxcJglFC3SGJIXTq2vuRkFKV6BovrIyD4q9Svx8sfXBBROBoGNmvm/wFLvJ
rLnrmgZ0DZk/7aZmn2N728DrrfW2zr+W+XwCbJlrpWxR6uUCnE4uw/wjVWAQcwIt
VrsHTpeG8X+xB1uanC9J5ZBv1n4LVSqH09yGTLlGi5SxiMw5Ky2+6ooRrZ/3Rr3E
PM6k8LAsfS4fiYr2kBYcHPQ4fPFYwiIU+rTi2pcTrett7kK5wzDc1KkVDrNk8WFN
jVbtkdt6KLgJYntoeXxbmD5lMFRn7U/BCTLZS1Wot5kHqsIUQIjRENJO94h6cjTC
QfNc4CpVIkS4OUmKIuFksTyLsEDhlsPOeUjQque4pfsm7K0AQP3dV/4fMErjJM7C
x1ofEHGeumOA+hP3dZZGBb3I9ZDjtgPdSRvmJqQvq9EYCPdNnl6r7n5ekiNwOUJW
gR+hnkT4s9lZOq/0KwqQSawYrSj4IZtjVzGd7q+0LrTIhz6EoOePwUWYptF934pd
K3RP/hrXEGrpKNDUFA/BEN9TTGEdT0MGJ7c0kgltYmHt60+xMbZqSgZYjjk2JIyA
aklI52k/BZK1I9Fk3DCKaRlIe0LBPvSWsBmxpuTSi8rRnSI20E7viBX9ZlyqYIbf
mLfBT3ZRzzjOYTncdpAbIaifnIjksFyhlqxlMuMFtg00LpiYBLzdrghw2936iUVH
8xNd79R6nLcfI+IoJb0dXi2YsjlkX6W7x6q3vQ1ucUrJHMCf3ogerBU/W0tDFkEC
qXcsKSaAP7BV/u6vxIcQ8/GPpz1xOCBuj8AJSKCS0zeM4qLBOhj+X0ZSH7rCurCZ
YngKn3zGf6T62JFu+YmASu6/eyDJXRpJ00QVmKiuVX5FkcaI6XWT9TZ+3+YianV4
PInPmVukHTeDHa4mgVWcwTFR3AhQSSvIkRKa6ic98qfaGW/QNBAYfFoM0GaGfFt1
vnsAE/fSygnB2ZrQHBwTSK6obh4dFgz/YBtUIrFk7YeZhpaU3zhPnKTEwGLBdadq
jFVPHhU9/+JRXZqWiJ8KbxPYaVbhAdd86fXbK/EMQIJdcdOXIsTRu5fFkiu3QJ4U
vphjakkNCi8N+7FYuS+sg47uph7XBQ9rD/fhRL/zej0yZ+3VABscj0dir0U6/U4K
q75FWXr7IEiJHFH5gdEoyBAAMJ4oY5LZveR4bl5yT5hi3mM78uSuXABCbk2tjgNs
x3EkaUEcMe/9mtWPfEidHECD5rYRaJUIADwjgoRmngbYRAikEivAgngrMB2BgNlN
uH5pn9uFVWEw5vR8kFmMtkKipCeo3kLQXnHAYQuJ4kJukRQH8pYfRH2G9jxjjwHm
sMiloqbl+u3ShdWUEkeQWBYLArQT8LiUMYsnV8/UwP08o6ztql9ty5Phg/pDJMhn
reU2gQQUMZqh/3TTHin/nvR/HNBpoD0Z02D8LJ+SrWp9nC7aOH8OIRtZ15DieCCv
GbJnUILp6gjlxJwzyGgkPlY8KcbitjACXNMOiGreA8RE6vNovWnKmAkKIuWpKzVd
mpX0R5VyUcdodmLhAA84nT0R9AofX6akq9/dC96xmAjEsGN+1Sbr9DTqaIXgYz7j
fyvz7OGUg2Gfgs5ymgWp1bwACxcIMsJySCDiIz4gJGMZgFoXMw/Q3euHY6DvVucS
b8TUmxwlmMykb1nP19nvyOPRkKvFjkrpy+8jNrHOX8rSGJuxW+PaasvesgirABUS
qiHThjTnvmc0DyW3IAGMSZntz1N2J+DkxCLLtFrIMUrwyN4kae6OGz0gQgdqqjYE
nFnrmdL3vV6/P+fjvog+Syk2GIzyuSxQdUhcYdId5jJXmieab5FAM5zdbmynQISD
WOV0rttG1sftV/XN7NwRSyyKdxAcjliI7om2IzwbNR1RetYRieAyAO5LORY18s+i
gZ4NbjolmV6dRJzQ3QacxGwYSAnWn92FhI/m/nl8P7mYEgozrBVnhDFufsAyHc2o
EWSgWKXt5wCEwrwQ7o7AyKLCXFEHk3NA6eeLUGVptTDGTF/2QZIkETYW3wsLnfMG
MGFrtDZrK2LZ7rHXnjX6UpetTb+1nzDCUjinsio0Xok1IV/3gdZ2jbNeyhIqe5v1
a4/afHrNlwsNiqnC2afHfAkP5pS1gh9PGJ4uHEF/TzAPhYq70oOcPu7BOieV592K
uid2iNLOg7VerI2kMVVkETF35G3vaydbbkq2OErNbKDDfihm5fPNEyMPiHCykohK
7GX/kOK99wzv6prcamCOQIjkKdzV5F0enwTcBqjm9u1ISkuaOUZ9hnPrAa6mGuol
ZGHlg3lvoz4Md5jyZ2/XIp82IiQkhZjfhg/KsE+i5QeYZzfS4EzU60NJpBra35xd
m5hXY9isJiqtt9PoSqpso5LljPwqg33bMEUIHP8HjplWTXMeOI+vLq7ZXPWgR6eo
0GvG1OYRNoyzPZwPTUMd/YKvvV1Z2sQxQqwUFNu8hHxZp7dZ/8eXpW1vxxu6GPFD
Haa/+Y5k7P3eYO4SftGPbqvRzaM7OG3mMsy8DYi+NWWWlLatpepnUAHVTf/asU+W
PpG6v0YTn3Zdqu07b56yjzuoAJdqczMZUbCA0fY8Tsv0pvBw907ESyvxME1HD7UC
tG5ry+Lg7TADTQ+6zdSkIsxdx97P78FSAUtwad0gwqiMNWVVNCxlIZXlN3O2iV3C
8Hf5hnQ13zywtv1Zh4N9Rx1RGqCuPyNEctupD4J6+oxppGP48/l1yoc8XrfwR8Yv
gUgQR8IqyGRmCPo5dduK+6ABOZ+03vsAaOb+3Q+rWsYABsvO4yzSL5JHE/XuAojP
3JzXJpFBTWqY8495jRwHbIxISYilXA3ZpwKw5kMmJR/YATiiBsrF1WC568hOd3ph
e9D9TejD1ylBcQYzeeVf6MZRNDI6L7CLQEERj4jdGuqZveErMAAqK0PUzslNxI+C
dsUb0imd0IEDRqCoXNIC27Qm+lTVB3JFC1QfNnO+AVCz5/sE9JXlesPmzKSJaPIL
hzActblh/wwjdGkZkJCuuTKwWNv7GWC3+Uu15Mv8CHox/X5Xnp3LwxPPtqbNYqBA
y3aZQnFvfqbQWvrvBMszsVfO3YhYjin5/5D7dYXdcVwPhmmLotUtrhmiP+KsX9/u
MyM6BLWZ4al41WlTS/3KL42D16ISZnDvZcrGJ9hm3+8lIvl8wVf1bVoHrpsquw+e
GYwyQtjo2jS7pmlCDUr954My+9MGMOdd6ZYW80i0v7bRydJo0KM07Cfkxi3pjBfq
XUpi8Lv3YOhiE3E09e8EpSn1YBEAcUvCDMWxhyhVtkb2Z61CAWbftTbE5GMG+Kpg
Vk1nS1ovPXqUBljCSNnOXCFHYtYfNCBaHMivnO2c/5Bwc1fDYcry8GfLypKXF0iB
iR2CwjbQwv4nNNPv4MlnsaxkDA4micCISTlBT3vcOp1QDymnydSIHHsMg9IJR4IW
snn+VIvKHROeLTwVDpucdSIXdEpprZixt53BXzLWg+RrRY1Q45AwmJINgCzyK5OB
uMymePR9nWYpPP8qDhCsMGpUfyW4ACHNwtHBK6jQI6PTv9MRY9XnTreJyV0OrMFB
UZTNBCS4rbJy8uBGiNIDg9IZnBumO8olqRtEcGyC78iftwurMKW/pOJ5hevQe6Wq
G+sxHx7h8azmZgvMtYKYd7JIS4E47h+H5gmwg9CTDNTxMy6yXhB/nQwNtGsgb4mv
IUB+Q4+VVuk0wODH2Ehlki0OcfGrEq8UJ7U2d8E63RHiscuQwOfFS4iRHFxzSKhJ
zxmr+KAtQebzK8dFrtMgGCGowUjnSFtw5BBaR+N09j4SE5RcFjfSN9FTSGM2EHEn
FUWZxJbp6gDumcpsKlTqFwWV44cw6GcfTjgYlE9XftXj+2VcULZyITHHE6o+Mlro
ij06E0D+6+YcYBwpIvURFZImPZT9BLEVUw9KcK4QZ2AUbkn7X+cD6I/Bbq4ODrtf
3KiNoPiFrfIZaIE5F3B1RkNtmdJHm2JmArrOeO94IwEQ8WK1OiBNf44U8ul0niOM
h7o23THJSFnmaCQszCaulZu0xberGOoDC3n/Ujw+LklUtQuzXG9neU+e73ANZpXe
ZEzZk8plEPDpbgjRPyl7LS65obo8XBUUcFfqVLfCwqRe6Nhr+uvi3HYdbgJdi7YP
y8PF+bMAxSWU6cqenhql6N1NjEYotJzcJnz5o53OUsEPjfIs5jQ0toxIE65WYB+T
46s42Z889jbEQOAz7U7YWnelx7REWvdCELDGOQo/f8kKpwRh7sm+HJU1TyEOfUqy
X3xmsSX7155UaHrvD1hysUh5jbqHQSHOaOr9ly5SSNyLaAkpvHs4upP9HPwnDbTt
ww8HrO58QE3yan4ykSPTp90oddZgn7HFDK5rP6IiY4WmK9XAjr3mKoMsg9GQV7FL
FauhgoNhBElUW5tBNdTZGWts2JMHqjIoOxvgq6FnqTIwzbtxB/2aIdPTa/zs3xIB
n/vNZApN8OSMFlzga0UBpLY5HfLwDzsdYdIo0fFZIIumy/Wkbe64eMEs13mlMc9t
bbxA2T0hPUyaUGUzt2fR62YKvHeKw9yYVQXjV/RPYDxnMcqkpEGED+mBocAGQYYa
fFWyZZ51bkHbCo5EyS3YQL55ijxyuCT4FiX7zhJvkobcpKRKcqgHqtvg5dZCkYrs
zQiEt2H3v3KiXUB5inDBzDWzlpNm/7czdHLMFCmG1RsGSdG39dzD7tBOxQf0Z3pb
RrmikAgHk1HBykdM9a7yF5EeeRotPedPGzfl8lhWz2iCQ3dmC9rPF9HRLXEpjGiE
7CxYo0J5m2lLu51zgisSQ/TLtkfyiygDuHqsblM4K7YvuYCz0EZcQfx0x5pxmwW0
ltOhlniTTx16JZlMOa8VD4yUnFzRg+ttT1gwz+q/ULTFJQJi02dfDjGNTvxurFJ4
A7Cs/WxSVVR8pkWixwSFKYfdgzrG5R8gRg8O3yW5HR/pi1Y8d7nRkn6qRHXRi/Ux
vohqAb01DaJz0+HcovXgZcR9E+CWOu8/jdfx0M43z3RsReLs/rfskN9eUxNqYAA/
FFACO7KNIeyfznrza6oPjg3C/pFFLAXWNCaSCwG8FxU0S+U0YP6BsoNrPaZPh9cS
GZsdxJlJsrMSQ3iP/xjaLWplYTu2/Oc8A2fRTHAAE+hLDRAPhaOulQOP9SB9qxms
ij3RQ+UjWSNkyZuRsmxjhOcvSH3CXU/3kU2lGvO4zrLg9KNSluqgJXylvozrEVZS
LwJC1DuG+m3F/cEwsDguVNxYa2VRqrwxBAfBLu0QJm9fbqUjjJU5ZjY8GnSQ0W6b
p3b6fLGrSyytxd759j6vTrGeMECkECXRd0O4x9K1QLO9N675+4+ODbq0D1E3Al3r
a+XubpOb0W+qorI4JFNdYEebYLfKPZ13i7I70QlviU8n57GT3aBhTStU2Qk8bjlY
UcXHk41dh/pjMhUGaOilyMz2p8k6LDpRj5OHzBCW1D7RcHZelNaP9ucd6nKOQ3nq
QZRhPqrFVje5482Er7TGUUbP/u/Dq6fjCZ7bvcWn83miFRbueWAEDWdDSfp8twtb
h//uEOEoI2hcaZYTkQTYHhcn/DnkD7IKa6Mdr2FNcJ+ejMKz8l3Ww50VUhFrpxv8
Cks/3cdMG8nWIr5W8873pcrexTYilkpr00zJanakL1rQyDRPVX98l5tLcNCmd4nT
NuM3tqlXL1pZBPZI0vxS6zoFKnovRxmOS+gGkWpwd1MGlzbg+ojMzFEkp8qaPPeu
I5N+8Mx4sBJDy3vfZ1g8pR+C7dc2VWnEwjHrdeNjopWmJ74H77Ff0eXLmVGW9uP9
o4nVYSzMVg24N1NH/TVi/mamB5LGs4Gq8g2Tc1OYz9U8UA6AIMkjYFF9NMTzG5eb
1RhGYXv0r8wDFah2e3PbQL46cQpwwhcoG1AkLXZgG8EfNcd4MWUIGqDgESX2lUre
`protect END_PROTECTED
