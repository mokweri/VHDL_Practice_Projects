`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vc+4gbqFp2IMp7ZDKSah2RTRDzFfCCpJWgwJaeuYM1kn1NbyMLS1LgNhn7Pml+n
6jQeC3mrEHxV8FVXHsp7WTorbAB2SDKbW+tJxFXzyzQg24NIp9cq7nIzNcVVMCFZ
4bPP4jX/07mKhNvo6aH2pwx2fpgALWU0WFZDxc6zyDTFLSaGlVaV2dXhrF49YNb8
hRZhGBG6BlIGhMvLMWtpTUJA7wYje5mOd/xNiYlGUBxMISIYV5fMYOik0oBV+5oo
TwyJMwploClxXAnMQME4XHKjgXFEqebHf1wGeM6NKVs0BrUGMyHqMew6AhrwQPMy
xO7C2ZKprd8J1ch8UlgnDLbl/ucfqkQKy22aYq5pG0sJpGg+tf4eibVWA4rNWyHT
jqA098L3LGpCGhytecowzmg7UiGvUOyvDTa/XnhJWK0undSpcyrX00kMOcM1ccMU
SVuSsBS2oOd9xDxHYiylxTLFGF/B1hmZ7ixpNAIbqMIINy3TXWJfD5YXXxPL6ahx
VCTAGL7C+vbuIawwh85IPDCvRvPEBpeH6JyAGrrOq5MB9+X1tnPjhrNLWyTe9wYl
gHJMzkf2nfTUeaGqDzn8CW3DYBSgqQYFDLQKCiS6M0mBh5zSd5xVoBe5Ohq4AMm8
5tN22+hE9UpnPzrELrH7bl0zIgrHKjF1d29ZiYx39Hnz4jiY85OMrK1RiYDfdasD
dCdfXAQj913vE6yiRijkwWIQ7q5RT7mk6Nf71SXH5J8sC4Ns0sOcqQgsR23nvTmD
gROjYgkKADCgUdi8Ok2CaeChfQJAWSn6lcxhqyikOO5CcUrALd04b8Q9HvpWTEDg
2/yZwCViYQOXn+IDE062Vs8aAkmyQeAn2YU/DTu8POCe/AvP5cUZxW/W456IF0+p
`protect END_PROTECTED
