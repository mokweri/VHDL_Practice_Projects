`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mq2PdNCEM/y1IJOAdDrp4ws2IN2bIXn+B73jUzRloAPQm934dfm+xiM8QM5buS8a
TznftNN/sdRBp1kfaXHzzfIYhav5TMKGbONBIdjbY6B4fLDiUNymgB/RIZpKkmkk
uwf/wYqJR5ajpwrsDJ7OTYl7BsQnXxGa9EI2o67VaV/HRj1tZo7jVa5+RunjLyIs
y16XcClIibLhmlbZFlEhJe0X4X+WCZIS0hhmYi9++UMGm7VMesk3k/RlKXSRnyj1
SSI32mwsqf2jv2irA8Lk4iH8A3kPD3H9obIeIYjYVIGfmWdhQI+DYoY1xDW2xkPj
i7dEClpDoCgvYDjMsT2yoJZFemst9DD5n2FNaeOAwyoggBTP2OIpo4aoW4QSQD6P
+lbppsaUaANvtCfv+/cPBsMWvEvHk06XZtYmiL9KV+FeXROuSiQUj1VVVuy4157d
B/4YpeafUq12sY1uBUX5N83quOWeq7e9SM3g7HVEz/bW1mymptDcqaG1XMN1z5sv
ytGSU//4PyoRN516S0WLAFj1Q5hZtZj9+uEBOiBONUI8F492nFzf6K/64C8iL1lZ
NepMlN4QBmYmcMoY9ytkBHiR75iUSd1fLfKvGaOif0kjswWDmglB0sebMcaLZwRF
CTKCqGA5ZQA69JRTR0Nvc+Mn58t/Pc7o2wmLRMXKjn3spqsOpM3xsrRRWqjdJX2c
KdIdfFcWGR66YpNhaSVj4ApK4I4Zmw+1ZkAOoMeiAOSssuX2fQDqfuJalLUV1j4m
INUDbI/gdZjONuUnaQEIzK3Rv105YaY64DzNgj6eBJHFJ7Nh3Yy6mZplcDwofQYE
eOIRspmVij0daNuI0aqmOw==
`protect END_PROTECTED
