`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgF7uQhKv39KLE90rAS2sx1en7ypf/k4Qx7KSSjx2jGbaCtGbjHJ3wvI1HY+kG9o
hZNcXi5ROXUW2cWaGjMRfkANkoqDmlvvkYoWz7EHj/HOlhWMJEa7AAVpM7ZxmMoo
KVod0C24MgWu9vxz5vFJKkClhSHr5a8cGtjxNsjvZ+u5mTvXq2PJFWbtK9a1DJap
Zvz1O9mfeRUwJ/8urIGl1W4RzuY6C2OYyRoqXZVLStEO4CIOUMvm6fTUypO//sAU
t9MsIHp85zJFKK1A0SQ886Ymezr4OX0C6Q1HoRIAmusd5ElnAnJC4uy0ZJ7DAtM2
FZOmTHnx4pNvDE8O/5z7VSwiIhU3JfhDTgoKdb9T0iuWvoaauUIkRLzMwCbKKpKj
m0LOr+Gnff0JRpD+L09OSBRz0I//ysRlz4kSkXYFpWyb/H8xo2AdqhG90/8vQ5zX
gdF//T5TIOg6buAwbIb528adnyQpUdvjwsuZoSG+5ALWa2Kdhp0lDxhHIzRWGAvr
BBBG5Q0s5wQfeOYy8gpuVP7Pd5MbUJs6XbczBsS0arrORh0dwfkUAKwhQmyhoFjb
g+ltV5nnZLBn22t9MXgRH6SfJKMU+7rMmhDKYxlmaznA3E75YDo60O6qnGBe91zC
GNevZj7GSEOQEyRx1p3w26N6atoPYXq1aXLNr6CZi7rns61oioZpHTmJdIxweojg
e02mZxQjnSD+UTafqBNc32JXSpKZuqSocRD5rSqKLeaobjLltpMFuaSjc4KZDLaF
+eNjH+Omp5xLRzcbwURmO/0SlngK2fMS9ieSuLiaGhTgcUY+M6AcaQnutAxAh6I9
pg6TVPempUC7Z9Q3KPe1SFFE+mJBjPJKk/1n5ze78v0GwVyJ/C9gHBjeRMap9SLw
MzakpD81zaS66bc9uM+a8IT35RjmByZiB2I1Nl3cBjaBt5R/bHoyAWXt4yCIDzDL
u7VKj0SzbF1911e18bY2ovpP7T2bOH1uIaJqIlyfugurpdV5ThWoX2v0Jm0ocwRS
4B3q4te47qQwY1bZOsmB3rAwV0VuOxlJTGQislNq/apK1cefGpS1ic8/jV36N+k+
h86Evyzc6kPo/JGkhurGfr2DkAoDXDOUqKVDDyzRf1Ep70pSO6n9UL/Nrlm1TJQD
MpyIxo3MZyjoEsE5yb28AR49Reh6W8tBj0pOIbFkwNpWh0MZPoWbRYb4j4eKhxXT
gmFy8stgkxBRQiPgVLceCW9m3aCraPVBIEUBNGJFu6C3MGSkCxTLXVwplzfTaXVp
GXawpaFk7RHM6BdsPk8rt3CroFZR7sfnycUbHm70rrF9sFVCuKTDczwtkZTPePqE
KL4RI75COuZgU0nncFaLfrgxUpbyoLNKqP76WA6VVcGS3eDlvySGqOLYndd5y9Ap
9wn8OonD/mpn2G/TjCeR358V2Nf0F0yDo8HLM1KQR1RUHPI1ylVddCv6MYFRyBSc
6L2zEIXcBxsiSXwrecf/y1+TUxVxAvSAlK54Ra92os/auoVCiom+3KJXlvHGxlk5
4ZzwsY7OGE+DACVSHCi6BYKSt0jnd5tMDaHcOxGoGV003rDjcHBUN4iCurVGaCVZ
cuQNtuEMV4cN2veacNkXzs4j+VfKTYlQoNQW66GH+Qz733/JxgwHNJEcUx477wvS
CkpYsGlx9y77xtNPf33LrqVnw5HO8bJ4lR4kbNDrcFmjBuHnolNN0nRfAmx3HzKm
cJQfb/9rVvOWyhQib5MfkNGC8wzP7WGAB0Q5dwiuujD9sBMBBglD4R3ILARJTodE
cqqkEKye9lgcgQO/ZvUsZHsAHw4fip1LGeB5Sz7kAvG5OB/d0BItiMI7wLydC+5Z
2UVw1KMrOOKk1HINdel97gXhKa1727Jl1q2OSPqxyJdMCC7vJLbpaH9EhiXA4CAr
6Cv+LIzEDC8OTLUOLGpPd0hR3+W2DGER5bhJTu01Mt/TzUSLHuU4o6TTxDxxMcS9
VAZCPxSrQEcfRYdR/gBv5NEbCY5dSwX4IR3uTnOZnvHlRNPkERrqIEEYuQhk0Nhi
eam1NLue4PQl2ubRS4/yxG4KAxPZk1FERBV+NUORwa3mruvAmsiHmAgdfKsNgISc
BV0CODyGHqIIFn0EV8ghfRl4JeIx5giXWmDwOE2dEdQ=
`protect END_PROTECTED
