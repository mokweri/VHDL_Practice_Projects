`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rx5v8QDl8G+B4Ik5C+IAwCs7nTcADcNXNzvbNoU3GzJN2+2mmH8YeE0HIMrPpdip
zsovwpYLPZD5nWrmGO4r+u6J0BDBUsgq5l+tGnlz8xvwlK5HeY47K/xs/8SAG/bG
4dvDMqJqrhuXb8Shwd6+AFBHBGl2RGPM5G2qfAaBRVLoHTjjXI+N1faK6WVaTV0C
MfzcVhVjdM1X0aCfymAb66y46hQLlCDzmc11GdaLsPSqFlHfWLTjAGof5FsfeHzw
+wsMHS7Jg9H5ZQ+CYkhqhja9mM2IJBuvZdjS8dkgP7DcIjTALdNpb8igvKtSr6g7
8OP0A6BNTqnDxpxMepanTqWNyZsxBFMkYZsriFCzDTVRDCPwg4BlD35lfcowmF0U
LZ6wATMtkwPrVeoM2YfQYXBPsUknSc9Ni//l9lyBWIYYp+iIIvVux5HEvR81Ow58
+fyrpbN0H/qHNr8djx9h+nhniL9S5/RztSxqgEs6xzJUFaD25GYLB7EJOHGkIOdH
p4bEYyqxoxXUmH7FpH6ET9J5wOS7WEM9Lg2kqW6auolPURV8oxrGA0aC67PfGOcX
60OzMxAYmrm2v1FPAg7SpEJ1oRrlmwxP57Pqd4fPKnNYC7G/c0iNs6V0DfeEMHEL
8uGrsXFUJNw2U747zQP/Nme9oXETOt64+stqyiSSZ4ekVjQDHueKiNmr2tJMVnLn
YLi9F/rPzdMXcYIWdS71NrR/PaQhq8rmexsYHkO14DvYgtbbdN8yjyxmTX4DUhAE
wwYYtrQkxyVrxWcXvMGlfPJmAl0bqbsLUxDIhFxrjsqhtwKK/FIWLG3aOou1azX6
tRjmG268tp3H1x4x6oziv97cov5rGv5DyEpQ++XT+42GA9TLCKCPtIG7AE65/fby
+x+xdPs1SnXQwcVxFcWIuns5lYQC10CCam1KOXaQrddC+PaiBMP0FYhQo68rcEAN
+N2pl85K8YG+KDY/OZdTbNcymobVg3SmpSPWP7Pbr2aZRtkmbVBhXYZrjRG6dHDY
w8Sq9ld6qXwJgmFsV/Nc8A7v02DXnN2vDNmNL+Y2F3NhRAqWfCwQl42khiEDO/5w
x5w27sxygbIeNVMjzHvAc073Ng/Vq437X/q0+OJDJcyTjSFNXhhHttGL886wfjiP
`protect END_PROTECTED
