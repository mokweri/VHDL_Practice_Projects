`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTgSPsV8Dn7HlvKvuTbpr9s21XQa3RPBI7augCs+tI+YWOSaQtJVIey+jXCAbogi
4VaDz3o7y11f3/TsVevO9jS9przfXOWwD8Pv0tmqM/zazFG6zA4aX39tlMKWCT5A
74iz5RI6XJV6okFEwqS1cp8v0DZrsnOttIzaxS9idSvkXCiEpk5K2/T7gEEZqiId
0h81zkCCZZcPZvTHjklWM+BtIC1VVab3JGitp+DKfut3DXvU1HarS6hHgg+EYl9j
g4bPvuOEk+8HYIWpZ/oSdKJGMeWw6zsTnwoy9Gop6irsUaoO3ukgZYHHJQjKcRg5
XRHi8ZuWSW2Z5oXbSY+0XtxtLFnbLsAyBr5BzMwFY/yjjN9jVK77gU90t3xvYazR
MebMbkmG9zewas7nLuegr3zO0wIkDTVyXsVSXSNGcNdRLNlk98e4XwYVcXmytP5l
C3fpDgVus/5vGA8o5cygmPLFdVC9RYWLP+QV5ILK0sY=
`protect END_PROTECTED
