`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiKBK4LHdcg3MN6+t42BuW1YM6fbfesIyEtNRIQ99WO/cVDbnnx3cAOv+Ez7QjMp
STLC9Zduak4/Iu3NaqMhkA7fo0x1r2lunfFm5lUrXEKz5PslBV7TNP5t/JUtoF6k
3fKRv4MOOZw8QirdMdEeGyITufcYYlIQ9Xfo84mgIObqZeF8t7cqG9KCeBCC1kVi
BeSg2F2ZVctiAcq4Drpd9nblQrx71M4vSX4j+2WkeRYeb1+4mIyILnudZP+4qYKM
awh3y5bc576zwnWa1pZFASEG75/bwHX2tZiVtaV0QnqR/d5LD6NPwWHdQixgSUrr
I5BXfEl3Amy16sRr6OKRdimmCaSRHKX0uv34RF68OoKafkrQ9qrmcXfzdSTOU/8I
W+SqAwcJO2ylviX+67+oeTBdZI66ATawLmxmHV8otO7mpc7UtpllgacN+S5Po5WZ
fhur6aoKtYep4ghdB2fj4blWy7RrXOLukRxG99uKQWF0/0ltEAh0jEugxczyMx1c
`protect END_PROTECTED
