`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MRii2OvOSoQ+P1fsCOkNflgPUu3ETt3Slucw7/UzAJGDC1lu9gfBF6hHbRlrQ0F6
xxprcmeQd8QKHhLQMao/HkVJgssCSK+JFipKFq1/r+y3wRIC+XDNFbd+TvPDq+e1
ZHSCc4l5c7Yz6Rus/asuk1RIyFj34MZ0FNiibSsHieZ4lDl1lKrtvEdR1HX8Jd+O
NuufXxulAAXm5+CRnzzh5CcxcS7xGsAe5ZA9RpOp8xQsXh3mSUE8DX2PW58FO8KH
DzLwa8Pi1PZUUzEqJrdeb6QlMSOqksAbk3qOlftIWC/oLpygt3stA1Uk4IviRxjk
Vijbe96O0R5XQ4N0bI3GWKoN8Jjz1wF9ZiYVvzg+4kGO2ogtnNczQe0XUmpuqEyF
14VNTqtReEro9otxrgMCNUqV0n3Tzgt3wWLmNqTxUOqgmMXh3dTGZtXLT/RCG9Yz
phaZCcTtVRm8TMZzzyS152l1NL21ADVwz+6vTeNfejTC6zfC36+fGtKKCSz6N8dG
zFfMfCWE5vVaFeZqqE2+LqwmV0pvelsDxy3isRopWMG9X13EIN+5LIL1vADqd1pf
Jmlu3iS7ZDeoXi9PhYJQkLqp0vAgMzrXJVMbOXe83XRaGEdT6Lwd2OGCPpE3HxLd
/sXxMjj13AJf+5srxHJDC/K4qnp5JF6OwZHT3temIRhpVMhNxOKu7lfXX1fHsGhB
0svZjhLiDLvDt3U6LorBXC0LjmKGG4J/aLWCpHMC8XmS9WTe12PrETgdfAX8Yxv9
Wh0rx7Mf8Z64a7gAvbzZ85I7/Lg+mQiC+zSadAbUTkjQSjBlnsZ5+r9S+/DlFjYW
bAW4cQ4ZxaaFvVkGAJDAtA==
`protect END_PROTECTED
