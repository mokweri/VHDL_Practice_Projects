`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1zGbPVQ/uja3kyBrE+8FMKKWR3aYjgVrk624EDcAfk/SdbgsxIsRzTc5IkT+QJr
DkaXCdxtoV99nuMjyVTby8ffc9+EjmoGqwj/n+wDRrBOyuZCBxfzn69sseUOSHw7
GVY7iqhV0ntOUMrZ/pX08Zl7b2Q+tzaJnbbedUhbehsH3wvIv6AVFK8buOpgdObF
ATnh5pTsTj7r8w/Z6Q2OGnm48X7+nDd81rNez/nGiL88tEdFvuFqGs5opYgXZpfV
H28hAUz77fZt0JU4tKkXLwwdzlJ/xNP4CUObNO0w4n6tGNK1t8hNa7THMxmxvuM/
5Z0X+b/VA0vSJzH2T/cORMe9LCp6gME5SA4+yapv85UKQmGPlpI5rDpY0bun9/XJ
lBhZyrfDzSsXNm7Ji72/5oHrk0luFDQvdgatruV56U+t5QatpMRhK5UsTSO40Tsd
KjHMpKeACcIlsTXVkoKBB4pY0fKu08wOUzAxqykjjhjP1PB4HMSsh8Y8uVkkum5S
hzvt1AMcapuSoPIVLT4K3eOln6PeB6ofiqTsUsGTvF3a8SutsIdx76lnpE37MSF3
6qWXJ44gC6CVCRanqZPwdwntCiPG2c+ZGa2RQoYf51zU7w9LClHY5bRc25PxQcoP
6Hzk5C5KJ7N7Xu5u3PSodkz8kTfb+9SXaEA7vtusoRJYwyG8jFX+HHp67s7YlP1V
BYOktXEzybYJXYo7dDy1gYF0Zuof3h/nn3urSWaMhWT5SQWtpz9z7pJOk963el8x
MGM71CIbriCn/SdEBZoRhP6rZe6WRsWKDJR+Mfg9IpWoew1XrFwFHGuC9RPPyn8Z
sJBGdVM2uObGTRaMovaVPb+8VaXWFqQCWpLzWYmotBTeb9reQPIFcm6JmP1X1Jk6
6RiCxwtjacdiP/W6EP9MoGwt4WR7/wQNdL9OOyJ8ILXc+qFpyXDwjPvZ7q1UsWv0
JmcPbeDrRompt4tiQ8kwqFch6pZlEE2atL4PMVD0fgSHZgInpx9poYs6ZcLGzN++
2g0qBzyZKaimryugi6uoZbcIUwc1eo1fsSqHdIYv1cCPTanm7yWvF3030niYyKtD
6kMsH4n9GEFEIYE8CWRec4A6u7xHJM/AWHD4vN34JemyhFkrq1jLnoehaOAaLEo4
da5rhlJ/vJFnDmKENadwHh8UIHCVdCh1vD4ZBWJWBHVWgi0miJZ0TvG1MgzkqDW4
Siq7bLyMp+bVSLb8aUZYgHM0KpyiodcHYC49DIX0BfgbqE1ZLgEhjpYRKePwqRCz
6XdPFCdE4d5nD53YpKFYFZa17b3Are3o9/xOFeI9SNtbnahcmThwSW2O5CYas/WN
mrWNucoO8oWhoaz6tsEconAyGfils7+8BayaaVp1Av0rN5dXGoEPXaQ3iSGXsqpJ
hWAyidrEulkBGWgtnRJMhYOCGDset2uxfiLhlfS+kxsa2ia7Gbk6syVRgCfWhHwN
urdopFnirhumu3yxm/dge278Gg1fSdzoEfub2Z6jG50m4VTFHwAko7O5mLXwuhUp
ZNhmBCHt9fGYLa3VbbHIOkOicLiVZbUsZrDkKwXlU5JAWCoOpLUYRQeKtjow4YOE
njvRYmBCGmZuwM9m1EGkLdBB0cXyI06SsPZ4eyQHT8uE6VjcIK4zk/XAskFHO69g
jTmAzaFSuoItWkDvLXEe+hfdotSgaU8nLMSuxo1VZPy2enc4mH0UkhvgQ0xbaHzt
nAOADbaBOjc3L8qo8txgNHTRjEk2axsYGpWCBrz+hBRKoqAk2xALpWSF5gAGMPTR
v5tb34gIZKvM4uxU6s6HzuOrprsJ/RUJhER5/eaXktOmxfq1rgJjUEVw6BH99Mnx
6vCiir4TLogTzGnhJH4YKN3EgyQQYF8cmk2NDwYXi/mxjDgCLdgNIUXKrwr+IJ3c
4Ar0e/1SxA47kqRtGCXCBbMGfacPjQDL6YeBovlVZbk5pDuOqnIcVqaM5LDqvtiR
cKQUq8qTaZxz9Yr05M+j5h1w20vKdSaHzCyigtQESS2hQ19l9DqZ6hhjY1YJ/YhA
weesBDKNRntfZ9hi4wvQTZqS73AZAWZ5s/naTMBgpvbC4qBjwFg7CoSx/UiLOGHO
tE++CQionNLSNpjf1KOnoQZFOM+oO+Vg0mLbTZXSgAF9LYYQ0+Ytx7S6ASYYrf27
JrWDaB1Mq66qqivQ/gEkCqdih38+uvoPyueX/FBPDhzClNYY8iZKfsx2BusMES4L
4B0z32WQEDkREpwCI0KEuzdHRPjhNahe9PnVtxEEZe0sxspkoSBMe7cZKVYYEYI9
S31/oQ9Kfi22tMer5Y16yVgVAzo5lEqTImo+gVkh0m1ybuYNagKxJuX29/bBZTvz
12h+JNB4QKkPF0CSm1Co8Sf/x8HaWFUvrTZ/UV1kEc3nZEDPzAy+AYMDEk39IxqK
6Ayc51Idu5f47pKxBaQRFfHsFjoDYEf+Vgj2hwU7S1ZTro7zmUS29glB8AgSK7ij
v2nTLkANNRtOFDmar+WiSv56/tU7FRRmIbeWV5ObcPx9XVe5o+OS0RXtCmvxldsK
Y4CDT8w47u1yIQcGZ6cB5dYKiQ37p+m5PN3PW8WnRGgLdQGkLjYWFYzY2V+LGLHD
dtcfqpEJ3r+EzEuKCRL1TWO/oVxA7ndQdAVFvZgv2R9DM+3UEzNgUHrjzKwOeVke
gnBbMHv0SaqFAj+txQWqxlYA6mUxb5Cqz0LG60aLm0NWIkLYaWa3XG1XNNuRhau3
9Mjm2iavvDsa2VqTn3xR+bfWQYMF5HOpanU6RsuL5K2FaSXN5gbsY4IuOPqfLQoH
2HaeqdIKSdp/8bgzjFBTxC0G7y/JWirXP4dierf7+5J3uKIzyGGW3UvQzVvhWQRG
BopgJpcEIvycTMnc2lIJMy+f/Qp6hMFTQg1B3/mc64BRHLvBEZT18U8EAz45fMYF
VelgyD06ck8j00W6tkwj1O9Cn0TUrrNODNvD6WEIB7pLCJVNVijI5p4+HNX+gcBL
nwEE/jk6kBV8Zu3Pizste+xEPFEVBeJO3EKej1fwEBm6Tmly1PeE/kYRaephm+2z
4/xKy+97f4us5MWDyyY98xGPFpg2nCpKQRXn/rrZZWk0eX4kSnT5u2NXiM978Wbv
iXG1NIOa6mu9FrxKXwImQCYpqclURvMMS62WONJoQdEsDCstE2N64kZwbsJWlbmG
73B70EaSJu2VZVm9/lvWYcjTl/ZbJhHbVKkmVxyPRs6lrwsQmp5P2gFP+5PZYAQt
jRX/0g3a3VW0IvjbDKMUwblmAUPHVhAcLRs5N6exXTSaxIklRPRJvJZXqIKzTsTv
P+jrnfz5TptOyehpAA5lbCQ1vNyzNs7HzCw15xsFa2SOh1zR2iSerujwWtbH4WL/
GohyIwsPBlLh3jBo2VBgz0djqgnwg7nWcfeM/9deQcrEqrugwuOymgr3/fhhaTa1
pYGmbwy1Ehj5xVqVglJo3THFOkZlDuuTauAT9/y7SjlhVnS1ZwVLZMR9zat6ag3D
+sPvZwUxhNds3aqDyebONwKZQETLPjul2jdQdK9tikdVE8mNHkdPjKyGO9YzFe9O
2d0Jqpf1NX5bPkKuXkCh7/7azudPB8axfyqCTfAopup1wHNWn1Kgh0pBJrBhVPmx
A/B201kDnOuS4faAP4+SBfq+shBG8f+Iat74JfnjcNUZV8h/MEYT+fLFjIZ0SueL
xHNWCK/tXz+OJquqrMSI6AGHkx7wnplfjv+Pb/lhTyaDSe736ZkkiSVYXeBsrDU2
DJ3Shic15/DNiKpgXQshtmw4cCy7nZq83dm/DPwOU+sLdmKHH35CgPx/9YaCfWwu
tka4hUZomAILP1YFS+itnxeJCdQZ7E1rJb9OocuLR/vgwEGNusKVSA9inDXainsh
AVS5c61y3ftHFI67mkwkInVAu1f5qxteh8RhJ2YEHjkkLGrfqCK0EOiBl7sMkkWl
M76JM9oXimvJRMKm+jRlAo4FvXif5U1KWX3j8J/xiBlCjXkp0XC9kH1isihA1voB
J1N9F1kMl1PVNQP+gjOe9WGWmjHRy+ArQxnaCODJZawk3JHzz4vVUXkBHxTg9hPG
8G3zdCsfiDaKG6+rs5PYzfcgjZkbZYLr3j0RZ5kZJ2ccucKHhVUzWKy4yzdy/KAF
uLeVk71AGQq9mA+i3ZjEjsr0ThAsEI6q2zMuVSen7n3vV+XIbLt6MPaDZIBSQoRa
UvPtM1zXM2dZ7ary/D6VYTdI04yQ2dkmIgiVJqfWPVo=
`protect END_PROTECTED
