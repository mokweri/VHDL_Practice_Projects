`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMAhh5QlPJmU3gXBplQPDIybFWvOMY/v6PFcMopF9rlLolYUO4BlDkeR4tFqmg6g
JuDzBY5SqY0xPdjzf0+/fphMmy0v6QXesMKWknqdDfDl4zqINbNG4gLD7gtIQFpD
phQieFJID598tbrD3hD1m7LAh625pw5yaYGZlyknvktEwv1rQSdwp9xRYD30WqbU
e6o6/l/6GcOPDKu6vjgHB6XIVl87hIpySdlpFYCzYdJyA6+FUgqWgUIRTTiwwmUM
EqRIx31gc3RgLd3/CSfWj3F13lKNR2Cl0LpwP9Bl5xxe4IoiGUzoxbHqnKyXvY0E
+7iK+jCbBRCfHjooBxYxQ7WBCqVJS7LC9/UHMSsxL4VM1igN5xpeI6lIGNxkZ9db
RwoFWdkZZdhzXhWVcxghAaBCLSiYffVoDvIkOH86ONcoxZ5krlgg0cTtisTh9FEN
k79A/31KILwaalSkB9tnr3jrxXisnl6BcubwVbL2HbRT46tCEpyU7jbjYyyvk0RX
RpRSjlJauZIOGRu+cqYTkFW005nFxCyy9qZ5uGYeS/BccWVr+C0R1CZkK+jUkzca
IDg6tBO/O+FysBXJHrMiZWzSmu59tnPbyFFFbVpYCWcQIwIH4+iYzNGQAG3ccFGq
C6bNTDH+O2aQxA/jr5b9GmWNLv5DGiQ4/IyuM6M6Lbixp+oUsploOgsdsVgknJzL
ngbbF9D9cC2vh/lkpPUDrmGAxsHrrBkeewJwNP9fKgp4t/aNjxGSEau6oWck/fkU
8Mgsn7761Mw7OWqaf/Yac/32CXPm+ZglxLMn6lg9GhGY3r8qR9805jx8Sw1OFZxX
iNW4V94EPf4DLVvG2xnCIW//IbrOpKw9jYCshdo9t4SuXuAq5vCZSUXNoE/YsLBV
I8j/86GRWyvC7Vg/UrI0GSp4DV+eqxa9EfumPgbpxNfWI8HOatixIf6agro2cvFN
VeLipnOJJAZFtnVGqYepT62LNSDFK0b8OMe8nl/zOtw/AW224sBo0Nyir6ZlHcBz
a8w9hyoIehK5+X1LWj+YEbqzTJa4rb5d00DPBGX6VCoG447RgA+SMZGhnkATX10Z
EzbV0IYveJyFHAWzWk+SymA7uRR6wYLGXsyfL4vuLgBBuc2q0s2PtCOjqfnp1hZJ
r8fd9R5ARikxnVQJF5lBSdBb+j0fu1svmVtiL2+AF8/0vZqD1dXMvf/DQhHgPLNE
77CS1EqEhGKOapHnyd2EJ2TObQ+vc76V5xYEZ9E4exN3KhhFPU4L0TJalMPeOh6+
4StkFVMLFOeZOVE0v+0Oer7xG9uvtvClZT30sbnPxmo4/fF4Khm1SnmJvp/FsEdP
Hj0S3moPyW1M8Lwbf0t9/pc4NO/4XDxmKn9WsMuXr3s=
`protect END_PROTECTED
