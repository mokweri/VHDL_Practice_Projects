`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNEFmNNTg+Vp67EjebvFc7k04mDiLmY45qigVTkswiE4Ew2RMB8du+Bo/vV4g0PD
7+kEq6RVsJtYLJzPnQByxuNKs0/QYBcFnpIU1unzQ0KsThXGCusXwFbQYOafqysy
DBz5WX8bhEHzJ9wLjqAfWQopDiygRQobbWfBVtmfsnQri/5l8NCS4fqnoeRVPqUc
1KBFC6z+E3Bj0iHQlWTX8rZOqb4eQtjUKC+m6uLMG7PNjVN/RY/N/BN9aoBMYbei
DwRSE89DqUKtnblDSMPxRIjWDvRGRJ9wR2ZxezOCG/O/BVrFz9cHPeFNTaMzfJEL
thPTfRrvoMqO7EYd8BvLV67gy6Je6KaZ7NT30bquY8EOMiV36/6VET9za5h/9dHS
0zbhY4bA8Zvv9p3usZO25bGxE4ZSVuqae5N9x40X6U+1TQ0+3BVP0HZU5s5SBvN8
F2Pu82GuEJ0olLcVBbcqmTpTJm5X7kRJ8PqMo5CPfyYIGAc0och7pALVLnm/pU8d
+0yEy88kEHTVKivjN5kzJ6FKZOnrZPzB4LlN87VohGeCV+0s4W8/qfwd85fe/qCf
up3B8pU10SmCCQ5Fv78weLEdce5TH4oG/wjJhL7ylJ+lNnW4ZRbgq65+iHpdEoXf
`protect END_PROTECTED
