`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rhc+6RTr01jQ+iToWiLg4sDTQeLPxv9mMTeG428IFHk5vLa+ZFRMJfl1j32T+Ii
EhGC9nAhQy3Wa0nIQiLu64CBlhgy7+efNSgv717nL3Ys3XPPK0xdWO3rprJnXDir
KoTOQYE/K2W+6XtgEvr3Xh8pWRrpcp88CU3uFMVwFfjKVt/PKIodrG0tNQhZoUyP
aDajoUx52VDiSXsOp2LYP8Sq0fPPsM1KPVtnTVuOc5J4eetdkgy7sUTSLmvTiA3R
eZJVlu7SvEnzEN4zhJxbfUtHTSUUaTmubi7LSo1zz+ckGBT2iOXdEPS+7VzjPL+8
o//ow2qMYrA07jPMhKNXs8qjZvf09o2pYKXAHl3SQj6Z6V+/MT5NG8grdwgo6Oac
eeq77R5KyYl2PYP7IQcR7pfsbcN8uXCwMMMLxPOnBRVUscZ2EicrE903KEs0Ije6
xLI+kWlYkHG25gp+Qo3o30hzeQsa1eYNuoDqNp2UIOPuP4xMvSe3tBNGJGkjYbKa
qk/kDn7CD7Pk3TAMqM0d72PXs3m8MivjkbEcsRCBAYpPR+etBtiY934DQMjEzhHK
qdkfQ0kXhRy+e6rTy6LU5w==
`protect END_PROTECTED
