`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqNK9va+j5bE1CyzYfkJYBz7r0vDJv+b61rBgbj2YZAqLLxQU1WhwGovEuvy3n6J
pmk3qnRmWBNrrVl0Bu151uu28RVPmTcXd1Jk29neFTnHo7kSR827X4paRWPpba09
FyyGpVIEIvyJHjnKLAAWe6aZq7Xk/WycrJdGQNiha46lkxcjlWMnkhzHeneIanSp
aKmlhHqyG1eUTPidpDqqrRtj7HYGNZhTlG9YFCqytdH/8OqKvqDmZ/HsbWygmsEW
jdRj1PnM094iJQoRLDonIgU4Q8h//q2wimJarDPNpDHGfO4GyiNDsuSh8yCiijMU
kKJunPz1GeiU/GQ9aEOweKx2oI6gdewp/aVMTskPUShC4LZEVK78J0s7VhC+itFO
gPYd+TpY+Rh68EwPJ+Deqhe6c7/TW9ReYsHav6QPzzXe2ekNz8+vTYeR/dU2mjlw
GF/B+QczGOUGAXo1o3ecD2VkUBMywqHcAmu82x29WdnXVrovrdJ6mJZU9TwiOFdP
kqNKZntbV5dddqHfjXILni/5vyG+RgtrEY03cHK7UslXZ0senC59UtW0T86G6vZ0
JuzIJi8RHnYhnz5dERNLSltCiJWEAiWG7vjAVn+GTC3YMY+zyQnePdo/C1WO1kTc
KYWVhR9BboEVjnuEd7uqN6PiUuGPaj2SfN+IP9zvNmuVsBMQDSp2qgXVw6IjAX/M
uHtUBJKfIX6MoBWQDqpYc7Eoow+UAhVEBjmptdUeYUlA+dg4HTaFrEJLvWzC4XV6
OrIgdzi5xwiTPU09KD2yiTqhirC5fz3hq16CZW4BGGJtK+nVfNd2QYfUdF2J+cc1
ZtMPh+81LFEiKEVTaZHSvxEdAk/Zsai4W7zUOQjrw1ZprNNwaY8LsRfjVwytsAsn
LRvDTkvW7mwRT9ed6NtkO/RjN+uE7/SurnAGlTjgFmGK6S2oc+rhy/ZByTyYzfed
HJPfcqr6KH/lhMm3YoFWuax2hPXakYdhRbR7DOhnnJb0OLCK1JDWduj/xPw4TkeL
U97pvnKRwwwBXPa69Ph0KE4ZE3vr1kTDe0V5TYIgtumvSqhn0yCMdZ+cFd2VrPUR
472sSVrGSCh9WSTtNxzhiOsBl3S2Jm9jV8WvGJlmciWqjUt0O4sQYseQ3I31sIZT
68sUxLa44EWeso6hlbezq6ibvytSI0sPbk7T/t1HUu8NmJQaWWyNUqwIZ2ycJiZ0
x+mv451lU8+ofg+4miFUO0+1TbkDvA0ADkv8P6jDrnQ8dNLrJTYa5EUhgSESl3ij
IAOBgLSvrjNein1YXAH5BS8rfGTAIrIstlpZC9R6Ia7kleQjDQ3PEPmNAcHSk+5m
NaNgcXA5IH9DVy7wFQacaJiwLkOHR/UWBq62r56CFy+hm/ZFQxiqUuGRTbImh9vs
fMs8QtnS5ts4jDgrHP/SRfSga6LikZoTNri262A74HklYhPikw54zEzvSBwIWJ9R
FypcMd05BhaAMcVXzfWf0CCigWVTuE1BVK6Ps2KKxTIi/g+j9PBF//R3hOrNsHdF
PvJsrplX3/Nzbu3X2TNKgGIPRAHdY4zmGS2NXvyrGmrDd1+HwGE87Z9cKvpp+9w0
vKx5PlXilkm2lDul8AI2cvO1twC671KD0kS4m+4zotNkmDyNU7uwv6Vwq7gAEG1V
NUTwX3PeyygEdaiDndyAlgYpkYxid1hO678pXxGAYTJib6C9BPIXPZZp/0TbS7ZN
jDcOOMrBnl9H89gFuyWwwKWFeucqzBVDmZEHV+JuXwXdnvzLpmtjoZecFnTwKEmP
A86uX+iFBVV04DVETbqMrKzdzr2c9INQs851E2DQrBTptG+FFI+FPCS40S0UoCv5
mrfMNyNW2rga7yA+u9SQQSY9J56oCjbXO6RP9DlheY1mPWmPtKRj8ZQlHVb9gfmt
JEtql0zHsxKnWWya9pTQXGCce2SoMKlUwBJyuzJUU2Y=
`protect END_PROTECTED
