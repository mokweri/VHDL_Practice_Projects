`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OF64zvsjfpz7GR8LBhx2S9159OOiGQVq7fwOx3QpEMqBBVP8+AogIr5njW/jG2Dq
PU9fMYO6AuEcyINVRT2aO99q/MxR5abHPf9IHrgCWI7aBMjRu6goVk/uKE1zwjUj
3LyDXPFxJ5LuiWMqn6ycpYOYS3c85fZImXQ9Q0KKoTPNK1jUFOqIDx97mM+bLOwE
X/cv3vvQ16yDtRQsOUtq8FLu6DQJzr4MjEwsyYRXjHM0/rrs3gFFYk0ZodlQB+hu
yI8bxwVYcf8IWfb5UJqPpS3AQlQu6QU60N2hthAuuLyfd43w7qXIbcK6GxU8Ime2
lRgW5RWbFloQwYPZXXvu9Qp5PuSwOzYYmQG2BEQcjljad+YgevjuCoeA9Tb5+gSN
8GQJCPuwyqFPkclrXm4foUF+23GCpOCGLHr5ewUVhWwD+atGz6lZeG/+6i5vL9DN
rFLCoh5cPJG8uvY1hTpnv1fL2TF9sriqlBVbp8VUAqwBrJIqawWb53JUW3zLxXvl
UE7OJgXJ9Pv1Dsj6pRpoLaK/6PC7fttqKEvwiR0TRcX5Od8jsq67pnVekgu0R4qS
OpVIGXFHrTfXGCSMi+6FSQ==
`protect END_PROTECTED
