`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiuSOT7mrVYYTxebsMI38M1xUNTO/ApZxxGn7/sgh/ZGxK1M/EiJrn+OdJ7r4Thj
et7gR9HnEKunST7k3JJeT8w0LuyS9uOIgVf7Kt/zGsihzquO2/c4K15HZKODQGna
hf0nlvK0MXWgEY9/auVMUHkncQZaqTa/mCryQR2xAhgyYR7fCF+5g1Wu8MreBtwE
DabQaKq4NDTS80EgMBY/80w4InYyl9ZCDS19MFTJA8mq3T9aqISB8JWSgdeYQmLl
/YCV2+AUoHgu3ea2u1cLnWGe05ev6vtmPekjSoL/2clbkVDMg4XzPSDioYVrIWtV
gZi7xdWsrNzDAUxivINukVw+2S7+KK2khj1EqlRKQ7Z/ebqrnbQIpXMiLc8IM+aC
mmNc57Un0TF7uQ2WIdmC1fbLckCxliVDQf28PTRdmERMmL763IeJtYRwZ9Ps/oGW
Q1CwYVRczjShcv5I5IZd3YRK7m1GDzkT2v7olBfLQe/1QilA2XMFSTAyKLNR3QIu
EldTlpHtHVQm7LVV0k6xYfsQgRr/uwHUBNZu4CfSzzuMhBSEB35mr1SEKYH2JImo
xHFGlLstNLQ++vg0omGOjlVCCgmpwSl+49ANAICW4Io=
`protect END_PROTECTED
