`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUFnbH++DX9gqozog6LqEf/0XbDLiaOqHQ7DeZ46y/h969iPOMS/stpsbWNoSYGS
EG8LR1eDyBT+BML4ayDSFLTvTvanTEZ4//lLutmNYEQRcuLYPa1h7mReUOml3Flo
szmS/rXiyMPg9d7G0S8mCUJbe4sLgyno2hEN+KWmecvtKFgHNWN0JVmuQ+G8T8Ok
CVhXt5oyDv8gPPNPhh5uuMJsm5JpAblEp0wOc63ic6AlQ8waMDUBMZr0Tbf02QiU
xOrNmLToADK7aC7OHYlkRum+Aw6HWqF6X/+TZwm9yFKGpqvztFsdZ7hiuqzz5c59
NcvSFC7ef8OuXT6C70A91ZnGeiCSSbxAAWll/zItBWdUpdZhqqDiLcXTLZrkCxgl
vkLZoH89ABd0q85TU3KrOAyVEahlCiJjfAWw6Sq4z2h+xpcrUU85+WFBDsmujE/a
ra1kEjinbQEGuLzHP40E4cuyw9AS7HrkTz+nZFwxq+iXS6JH7cofY9lUexd4AJVW
Qr/gnIbpjCe4vo/Yff2xLkQnR4U6PMU59DaYf2lh1clAy18zMKeJGmblM7SQeZcf
/VwyeBbIX68le8+jJ3DYu+XfQOpnWRhxwVPWsZPzbyoCPYHmtKD55b7/cjAB2ZOD
5UX1bIAJkY0QM7zR+pZ//EnuJ0SBp8ySX14YS7cg4QqVz6qGz8GbOAkwvoL4H1jy
CHfLGHLJNoginoiIUlT1bZc2sx5N3eXg/CM96Cdsdek+s3g6g4mlmDMJsFWEDN7S
HPqWxGIbQrLkPXPlTp+ffnedwJleaMt7AOLHjNXJBdS62QVxm0QeH8QWCVFppVcp
j+cgftIfbY6mZu43OsJBo+Bz5GWrLwl2GVZqBi+ho657SLhvTmZ2ukhYpsGusIJf
wvAnPxrMIbcjR4sdS1XoacExfhGl2DQvHIcVlGLDofCiSevR9Mc2Xye5xaESyURc
hfVDuAJDAd+kZWbw3l8HfakwBDSjkqUAFoxFM+u5nthPLxdlYjAiarsAL0oXkEnW
gqp+k1J9Xaw78SGyKa7QHjbanyPt5s4qUzjZEtjUaP7tRmshuWUT5vO8Lf9QAOVd
G3IID1Wqq3B0mHyYLmfpzp0LPz/VO2nCbmgWR/7ciCJ1QHNzILyQjiw1yaRfJyXh
tcX4ZtGVN474TICdPlrwe9NN6uXse6NAqscO3VE01sx1FWF2aKxoEiboPBEnyRku
oAIAXqnIK4rwGOIZi+MbsQwQcO+Kb9EtLWZuZkyI3eY6oaRbbiNQ+hc8tiv4Y0zO
sWSl7BS33OFYIR+Oa+NfYzunKbRK/hfLbXEzoEPm8TCOvtzEovpDb4+pN4greCzp
dX2aqroFdLUlQ6r7V0YRpPyNudfTbgn76gwAzC9iT9mN3TOI5uTnuTxoNCMSaZmP
KU+RhyywJHdORRaUOvE/F2f/ZD9fMiXI2Sx0LYrz+AdatVhy/t5n1bHGUADT9eem
nA8GhYUJIy2MB1LVoByj4nB4yYuq9qhRE9yncmECwhcJVXYXfQABBtR/1qWQKZEQ
`protect END_PROTECTED
