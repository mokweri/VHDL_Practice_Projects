`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RYwnx94BUDfe7DucgLz16Y3UFFTb04kNmJ1XQtbaFkFOiwx1NEH8H6Vl3o794Od6
HqrOmjqHAnFoxI1KNVmaXCAR80ufJ9pRQ+9BltcdYJeWvtd8/YsSwGrcdmhqlD8E
4jvyEfKEPxcsQGjIc4sV/5LWpz6K1l8ziWLnZn0q1Za3k2PHzrldGaj3odw1nzN6
jQNlaWrbWdJSts8C37rRdVIffa9XzMrSEM+WUEyqdFd1tdrckv2avba2CX11EXVo
NEsTit5JKPMfpgwDydBxdTCpzAuuDJgK5hpv6Cn+/YXPIrUQGeBfDHwGA01A4Di3
JqZC9Pkv6uy4QxGvcTMyRKSuyHEQCs5ORhOkHNCbjkA+IT+zEcsRwCWhOgItsuC7
V13KBulZuHuqJf1se8zhO1YDFVNK7CUdS5EF8gcRLAaYO6hefgF4BcP7UqVgu/J2
xZxuknAZwfcTpPls3urSzHOyYJs8OKvJ69Su5mfB+HZejCsdmWafISXhd5og9Zno
gc3poLgFdt0SPDusNyAtjJKVfOk3YdCd6GI0bishDGwspHBCbZ96HL5XlT8004zU
K2DA/9a2/jBBzjEFKjHhLdIa/x1rCoZlFB2kZuwK26XeQ9nw5KnpIfAvYE66qKOd
ibdnUTIq+Lj/Z3oDz7CKbF4H8NPkImrkSH2Ux9BJNxorC17eSdqxvI3W/Hz7LxxH
CtnNyfOkuUbNv0ox05R34UMcQcmELUy1AJfJ341WbIN4AiIRY34SvadQypLaQQOt
f4qeXN0WK20yBi/caY55EbRxd3c0w6fViTEFMjgASZADppgJTYskjAiDt7QVFhhE
NEDpQrEsqJbSV/otR8wiIEBfv/ETRNfYfcaOLmcS3pwrPjTmo9jRrzlkzm6DiO3t
Nfe2hSD3b+6wWCKudlh/8dGyp3PO1iXdmfMISGjm7Bs1qIoLrBUFJa3iF6GjyNgN
PLcGCs3V2aJCXBHXo0p6GWtsM8Hsu5K5t9/FYK+R6bbS4O1GQOK4zYo2QvYO8fwe
OAAkYyZKtdEyHz8XUAmmLERgJWKA8cwjtJpJ7x7EkJBUMpgXkP1IZdNJ1LN3CUFc
2iC3FzRwyv+h2b9r8/u8te8B7/Ji2gDvXuKot2jgipQS4W99xclSl7kgDjYnfqSb
cvBDRn5MMy/x7i9fNV+Qm/K8F5GGA16lZVeUgYQRTvikAiwbyVJHwTv2ABBmt5oE
kzemyt0dgLDLVzvnzr4/ewFd4MLFFBq0okGbcogWF1OzHdNSS9s3cXjVV7jjt1mN
RhbLX1Wafnuz5UCflRe89hUm7rHmkeyvjlfzc72MofzLdENHXqUgdYbf4641VLaN
RJqgDBk/C1CFINminHn34UMczZmnSE/Qb8yBxfiuYs51wHexer1LoFbjvP48pEXs
vo+0Q7JVkpeaL8bknR4Pk81s3M2y8PRcO63qurITA7OOIR7uc652VJtfoOy57Um3
rzswvWJNi0Q+I6fsuhmX5K+85JNY2a/fK4ahe5b7HrDRwpt4/A8J+mQAT7r4U8+k
9g82H8J1w335MN/zn2/6tPVK9dhzHOE476+EYm93+Z/YJRQD7WLk/kHF+F/2N/EP
Ax+q5JtPQ+DdcPjCuxoG567bfar8ITRYtwt1Gp1qa1jj+M+kTU05WZ1J4BBvtd9m
DNL+YQVJxuAAaqBrfuBTpq3rplgwBUZ5ocNoe2533YKtPZrj07ac2X/StUPkjiq5
VMh/hsZLrz6PAeDbBwYSrJ3kxbhwjUoB5xOQgP6hHmGr06E7xB9JZxkBDW05UqRx
5N5rtP1MO4V/tkc5+7EF90K7UoZJvdEdwryLc5ihVtU8PqvqN01J6mz8BXgHYy/W
MOxgVWZAa2yLlEeH8y01Hw67MblpXXEsBYAJPN242oANa1gvKCIzOd+n8wVZtnEx
yuHgn/VDbJmmaILSUyFYyg3IBM2bDHPhni1xfBZBIAa4QoCCXNsjWfb3s3Swa9Pn
rP91GyiPhzwJN7/P2ifzRdxEeYOCmSCPv1EoccSDIlpqNuJPNVhd63t0wqjwU1Ks
R2knmkAr2K+DQtbDdAOaURVr3yIiVHSHksRxI2FwIW7oTwda3VjjxwzaeoZIOXX0
ZmUW4yRW4u7Y/nxX1ruccbMQVQS3qWo60/awE0vwxXFJ5PTqWYP0OQJHpNyBx+F8
Sf1KHkAIIGtBV0dhl2Orf3UYctWsyjojwTT8/1Qvxc/Mj+n+kRpt9UQMD4ikHX+0
ef9eTjXF7EZrpIIKqb5SQ9mZkVcgPFYbHuRfGXDhPwrHPM9orDSL10FFBxfsrGse
XVcfIZmtYdmKSDi/hYGy1+lEV4hn8LTca+N9bJ0j9VMuhNpuUnGxWCE5LN/Lat/l
62qcSukdrxJCjxW4DCRKx6lUQikU4c2PErgHpveZKDJxhtfdzhqM01buMyW7Ey/8
XroYGVRI5Ri+t8sM58sYIqXAQAybPEmSPohC2AIOc71vIh2r8N2NmjrhRoVGEo33
uQ2Rx39BzZXN4+bFdwBccrniBwPAf5pKrLoMJVfL8nueLBZ7sLlnMcantnnKi8YT
QRxGDtEPiuKF6tgsu6y2cZ/JV9Z38HBGpctIKBWpY79yf+H0vbLXIQZe2DnZxBrS
QhZy+7yPAzCDyIaoA9PUMtzJyq60QjhKh+zGP1OZvImwE6I/1Q5V7rali3h0w96O
+UOpviYvfXw3DH7lp4TLFJnaclctZ9hrTsD62+aGsx1R3rhfh0YQZr/y1tVoASM3
+jM2fhFV+Cnn78Txy0tKdW7+jgOJx6XPgFj6rGWEgeO/KbKyGd3hEYXLN8VZLbMF
vEN01NgqHyGuULgglExyhPDDGybtkeVBNeL3CCkdldhs/6V8NdXWGRUj+vv5QbRw
fcvccbyyoC6MfhmSr3ZQxY8UAEEMKc9gHuCHD1UKKNcr92ImKBxl4rN0gH86lbuK
625BWp8RzTIY5GTnb/JoyNRMPECFrmI0jgqt34vj++UsQZmahYr1cMj+GlTE2Urh
aKQxjETEM0OZckopSA4NIGA5Z0KFiJIeqWk9q7g4BZfanCLruSTBVyoKVFCqSaGH
2su8HLe7Fbef6hXlJgd5QRvadQ9+Xa5ZE9Wn0uSC+Wv2ky6IGypnvGxxf2uiSIFI
bMGxcX2nsgvUjc4NlOty5j5ufPVduRPz2vQhXhgKUmNXN6b+WoM52Gj30lYZuutc
zACkTGB6PklfaTCqZhsMn5DGzYp7HXJ369DDacvm4O2/U3K6Mna+X00MSXzgGARu
IILStddPa5DlgnETs0/ECtjq2YaNbPbcDFFEPOScSDGnvNElitNLesyuIz2ZOKd1
3Xyuz1OTrsyDKj6zBLOoVQAiQLHvDp+vabJ9hRyup/tXW7yZdhwqkPoyaD+kJ+ib
BPlcVTHyKS0zJv5AeOQ0ogdnm0H3vutv8lVaexjM5e1/3KndxoYQRf9pjx+mRXFE
7aHJ5Rg137cgsONgboJSY8f6jntdmRpRWKeaAz9iSFWEz5XqmdWJpp/MkA4z2ru5
gPdDnjp99dr46n6Wt83bggK3MYy/bsi2j7/NaLok/sF6wPj4mOy06wEKgZ6TdnAY
6Vwmbi3TZmnsrYhfNflOdLn49sIKwgNGX9eKeD45eLvwnKkL6DJZhKd0GG8/Lv/B
G6RK0mOXw6BlLCVQ3fl2ySLZOd5bcHxExI7TDI/L7IolU114Jt7m/gEoKyI5LQws
hhH68GOnNt1Z8EQHgpYrRepkLj4j293EDaOhksP+4W8ABA4Tq9PgYJXGXLAFXQ6j
lWTq4C9erT1GAothHerM/0oJHKbuu0dKcYy1fvOvgpa3hMq/99gAgOznPK20qqJy
pTiNWMYwST+kJn3Tw5XGkUJp7z/GgeQXBOkmPQjeM6BLi/rLts1tzQbFDhoFnyEd
upOD2mtPETBBuFXd5FnA9HraTqzUrWIotkGaPObgsNUSk7v7mrGyE+gg3DcwcbTR
1nCYffT7PMETYRpzW6C98RYx6tNULAMNqU3U8yZyF53tIrrHHQTHQ9+jfYxeMkau
wEplFOI4tLhuQLqNDfd7zE6mR5TdBfK08KdrBTm6zj7NdiHDKL+/VwckURW04GPa
AexovGNcGISD4kkONz3I+gfZfRc7RsA71OCaBRQ78nidb+zRpeAk1uyfD1rS3sNs
v5gTh50TF0jPFLTqwhzl3Hp9d0y0EUp8KOO6y+t/eSV5jjC2eCnEePl0fi62Ultm
zl56yxREvVVlOCJRAD0ptlIKclbhOtt0rSAKNjXwST3dlOSWTY2h7AmiYrqYYPVl
Tp86710H05Wz2GxhSH3umQ8evc8XsWoqrN/KryKZvDlYn23IdVn13F2K7duuCVfj
AzZPqzWdzLBG7hNShxSMJjzTVtfsvp+e5oRUO8zlG5c8aPvFiw0IEGt0g6W9lxx2
zIQH/oap9owBCSni0Xf1K8HDoipWq7AWfAxAyYK+9wp0Lk9hUEQd/g9QSAjwSClm
LX4BKY8rzvDQL4uVutul/MZJezErnpe/o1TQHgMxgXkkHHOwgho1eUtYm3dulyAZ
HAGS/d57YJ8SwnCMs8SsRXjvbBC8QtMbADlD1KdKhkubSa1sCBJlwljaksndnTAr
6ZLhyicc8/cct1HAUyPrPGcn55MRJHpOEVw7qUlZO838Dz8KD7wcUK9Ly29PgqRz
b6a46UxPSiW0rZVXmTdpOFPjCqWsLynudLXM/LfdU3eoKujrzg9MmtMXwY2Ccpzh
Yj6pN/LKk8yWZPfJQeVumg8JcVXcrHza8/sWPjcf/bRdnsLiV8z2/hNJvfOb+0/1
VPjDe0aOqpTWoP2sUEHpJ6QKZG7PpXGdx3JzwBiPCCiw8eUfXN/CjeUO5bKCYp/+
bDx4MXMfRItHjyLThAC/aeiKkSAYBzagTy582mzshl2js1Susuo6ymR6TgHechsp
XghmBqVTdPJhqqGLMp+RQ3iLioNl29ILNuyk9BGGqrUYaz6lQkLJtsjcb9EAYTMt
tWuRY96N6KJP0Rqay5oKNoxeJOkEwbV2UCLKe6n5lpVOuRZPAPOUsqDxzF7iUyzu
gg9XefqNoA2Yow83y4LGagIlQOhBvbSRpfCO3f9OggDdh3CzPP9eBa3kTvfBq0RQ
/+Gknw0wk7KZAJW/Mg/+ENdD0ok173f0SoqwzDvLQi/ALfr6lYXU4++aCjztF9/F
u2zWAVAtm94PAiSY4KIol2l0Hfbt4KAaEjDNy3z+hLRTlgI3k5/8WACjwgyE1cEA
8FW4u/1jDVfsymOpWHeORSjYp8NdbWX0Ag42LRd9xMPjhufrJlt6FO/SqFosOEMV
l9KVNe0ZxjxmUz5XC2YEB/hucyWs/UqemjoAgbvyGepHDQCjl6LALeBQRcw9ixKt
9GunwxvM04xJTfcJcPecwcY9N7HARWgvoRDQkkmm7mpr5bkZXnjfRGuJL1R6IrQx
Yj0eaQ4rKcT2GThIavicYgv1v0wDEGd1f3AVAraLWftlsrJkAfOe7D1s9kA6fKKR
SM/oi2kU/+6/UfxO3LeJXw+1WU/Kc1M4QqsXTd0+kx6GuHcwa+pwsUHpPNqFxR/B
XRIHTf93+0XviatdBi9xmaf6OFukpFyZG41qk0MAvPMJgHjgM9gnbD5j6axJQUGN
6X8LvU4bW+1KcRD/0INvALAikjN6B4M8QOzgzC9WKK8ldAX75819POjd7S5WvhwU
2vEJqwzUYy7VrJ1ZxouGs9L1DLe5XUNQO0U0ktuDCiXNGbPcIoaO10QZxSPw71fw
juADv/coHA1oZEef89IiT9fV0RuaZEbbPSMUwnsq9PBP5/6e9rp0f5R/vxUFxJss
cuWLQWzqxiFVcfOG5E4ExEWgdz/MMxKQZDb0SfCJgLl6RmrZVlcrwXqF6rPerDJW
uWAvYtsr2GY4DZ9J2YYoVw6o/nfHCIvIMh4+/wb1+z0yJDP30+N24hVsagR7aseo
lA6cYcoOC2EPZf8cEyNvubA+m8Pt8xwxcN1rgFDBHep0QFlLeNoqFuoH7MLTsYqs
ISbJsRlnrPcifRkXoO2rEwLVxhKgWkBvULLELGMQbwhwj8fVP7ID7kZNsDFGEFTa
SE7DPclXcoN92cS8eu/VCcqS1PbEsFyv/SDnpP9sDTVq6FsLgJQWVWjUQsDyJzeQ
PB5qzH+KE0TDnAgKLlDvLv/+ubEe0P1D0gnDkNcO8qW+zZtrxxtrRqlL0aRrAp2j
3PV4lQIKqbSvGcaZouTXnp9KWbZWK/lroL+eq3/29p8EW1RecJtF+DMPkEcGHtVG
FPWOOHTv/1p1SXkIz/p65ACU0DTcIgxrLzHshnu5giNGyNjkj2v6NkKJYDw4Bkm+
O3ztUUI8H3Vo/e9MNqUHdK38YX7B2/eSNsWxz59kRmIXj28QDBERRyUUHtBy7yCU
Xtxv6EpoD+/S8RlzwaUPXU6qLjbDLBn1B69d3BS0g9CSs8YYFZjKLhRaGDFntwI0
jFu+Yl4haw9KjtMJ4H0iEOATLWSiKDn/HG8K/YtgPaZE8f1q8EjHZOrVdJBu56kr
TWU/DY/aMQGRPfWkxlRLVstbNBBT8q7FAZK9V8FTq1FDhNhUeEEW+SMW78AfT7RN
etoklSYQJ+QvnyG2RpARMC3yInLjffSd7Yxd/brwjGQfxfBPE1w9kEuQvuKWrXag
HCdTG6XICMJDwao/rHFxKUtmjPzAqnTNjpq0iC/C1I3BcqjPJDl7zu0P9J+y3k3q
ObMgMyxHrmfk6Cr++Ikgp03iGJOC6c4pwo8CaOYbm392nsHRL3QL5lRFwkL+UhMs
CAmtwRTarpcj0CpQUH9gltFyGFSBZl1ovD8oOI/ynwOpZpFAk7WOKPt+c2tvwuHN
P1AkbRRkNSVZAUsROO/hOcVGa59wWV1JHBLP6KJ4RukyApg8PduAyEYeSLkpUcNM
k50yIqpMfD22888cV6iHONkW53o4Gi92hBlIPs0ILlO7UW67dqOUMXzBMNNREhWV
ufZ/HFJ0kA/f2gpPHcBTBDYyltNpRxokiNFv4XSXGDNP8hZ2+LQLx/2/e6lw5Riz
Rx2/S7jcBK0otnaORkPocbeyYOakiaSL1D7CaIVu01qHz32PS6pSqslvIG4O60qT
ldUlxBhqIAdA7JfkBk56Fl4FMyBfZc9JIf/Gho4CwuD1o9MZyiFW3S1AdzkhnGvP
y6kfPY40152FI7QJeF1e28hXB6UNlbc1zSQwz6Q+sV8ePwANSB8ChSxRd+xs1hoG
TNq4L04hYXPocKKxbY/5IEdL6Fh0G7wPcm8RIDXSxpY1fgQWkisVyuYdn3XA6F8b
ievCB8mQ550Cwox1TuLbBaxO2AR1soYfZw8CsUwdHdyHwnieJfmmvJC2vhzUIROE
lZyMAxLqpZHvKM0aAF+c7OQ0WqYp05CEX3wJo3TupNtq7eeCdg35UiqYNG/uBUgf
rhZs0gtmr+7luLem8SPYb1Zd2Snn1mq5AA0HdqXa9CTtRjG74ITnM0by8DHumopu
2iWMy+TSAshBt8oIXl6WfKxfnVVeRNGr51akylhjz6F04LxYAhInpEL2L4iHiO19
IPtkQHN+uPPdUHNZTtfKuJacDi+VhB0yyqHeZUZkZtr3UHbolOg02lu1nGakvSjA
4yDqbdqkpX2FyqPQIpg2zyDb13v3JdzX35GFXgPCrEiIf72sbSHG38dJ9Ow70/dk
7x7cJH+biKZMUhtnViQCVF6WCyJEO2KpI/o3NbIfBwPuCrIwO6ch4rO/WNlilbfg
vXeKKgaYuqikjCGnEuB4jcLFW75JZxBKLkzQkZTCBAVESbbWaVUEHbZiIJdUdY0C
nYtsR8yNvksxaZuGM4mg0+9ou24T+69kozBqtfxyFKx4T/sOj6CW947Bwn9dLE2b
OQYD0agRd8gmVzRpDYsjxh3CYqajSTpGZDkv9ueXe2YH5RCdh4F3qcxc9HZyuOLY
gW/zLS8jUDagH+yAHKprWWAiSNGSsEd4mf+oh5E8jVI02Y/DLtRsAHTVvTpW+Gjf
DPOOsqWZ6pV5fQA9HR8Y/WJB5Q85NcmGAE3t810PPCUG5n3aLbswTKenL4ej1Hzq
EX941bAVanki2/vVuZc19/nO0+RJaBEMH/e6drIrpHd8L0OMK+Rj18T31SfMs6+Y
RMpD85m/Y1FI7uXNYiB4E7jWGk49m0ty+eux8ewg7WsIphE/Kg0vFWaFkOZD1pZP
lWKr+wsINJN8ugIJ41CrgQOHJqEN5PwAfXYonViduVdxF/M1H1OTrc6tSsh3ktwh
qOpboqB6WnReDSqmAzL6042GJ5S58Nl4CGt0b5jKie92eYZJ6ehnwuxHOJIERsmV
J3lH9zvncLX1hLdQx2c+HuaVHeYrQRUVHKejLlUf5/6766lwaLFXr9fHhnah2uRe
n10zjrRkWkERN+XZ6si3O36XEr/qQQPosaIJkEP+TV2UTc94aYS3uTO422OBVSwE
1C86A2z/lWYLR5BM8zFMscyvJ/Gym5n/2mttntlG4DBCs/3K0KM/f7uKFL1jUNf7
2DCZJ0L6RekrRnJmJh+qAWBft/KfCgXf0ea5y0nCYQga9DEpWd3pJwx8LiV6vCnp
XoaoAuNBk5NC4ZckdrCACSPpi9dnh9DJpN4lta5tobzesIdYszO8VWELJXEeVe6V
dOSvw9uJRhGYBE+6uh0P9YqUa7NtO2o47yors+TYdSBLqhQqAYiJXSCjKFvoUYrj
/IDaQcmL7+2CT76kwiFtQB7Ofvmlgu762fIsibvwJ2g5adZMnKUK/iCZH//QUp6n
QJnSsyApDfOIGz1kSJmimkE+l5TEhXAxn0T0a/2FBLnLN63nNV7LBudE5cdW1i09
hpGgm13qO77a20gMmx54HKepjOk4BjLLHdUPsCCynkykV55CFfK7GE268bVfJk3l
UiuCwpSP9VXHiUyoc61Em7f/lFsVWvbBRCC1NpuUc1IIBujrRl8gAQyye+sUBgk6
R0WylJ3ZcrMriNsFKEnhWDvRDDS4GoF0Sq5q8gLt9vigxrzjLEBq9wLIvJQ3vQoz
hKbwGm10MQNwQdkuaXe/vk1T4d0meBfNvi6RYWOQjffYhc/Ry+WGh+HU+DapxkUU
88pnoUwg74YaV/1AfHIjlU/sMW9nEJSyJB31XlZHjWLNfPfuBogxM01zq8tGPusf
bgbvFRtB9acl+cLtW5SHDwyr0PTTAf9+HmHpP0IwYk53B+31vHCon1CX9o8MZq98
vgnTCdu4XwUf/Q8K02djOt8ahYMXc//gh0hvEI3ggbzf204hvbNF7YT/KedQmoSi
V9Ga2fYPMfiCBo4K09+0+il0onLJdbyBpnS+IsbisLANVWHx3Tgkao8d2j2B3g5S
H3s5STxbI+4TOXV1VrsFW4nZkE2wbbTq8v1Y+wccNFINGnTScoR81rW00XMl7XcF
MOZxFTHb2mvtVSxCHYxfqWeqfdzwhcZPEjaTpuzFVlJUu7hPnUgOzXxAKxvLg5Q5
7ELZsKZCLVpy5FPKlD/po7dL5iaSG7LGVub9Asy9oONYo+YnCoYXMx9iOK0QlUoK
DIBRGiH0bGodugdv8kqpt4raKRmq9/sHLL2+PBbpOvTQPMDDg+nsHm1uVefL3+e4
pAGjy7IkVKsZvW8IaVt20mDbLyOZPxZ49a6l6xs2Uh6fK0pn9UKn4LHAyX+fykZP
wRCgSSY0dXieYK5brHojAzqqZ2Tj7v9Jby5IRUmaB7OV257BiDU1rwvKF44ytwng
WfWgzTuz+sSebsSxqER4VaeHA1So8FoikuEGOvNAmiI04Ts1pgPsiVq/TFpgyASZ
ZgVhlDJxnvuW3nBbFvfBgDU8s2oEQ8VhduF13A4ksZf2mQifmzWG7ngaMRNKQxl9
L8GJzPnY9FTz33roWrPg62qiKh/rvipkEdMGCekWC2DHWzJQIYr30QJd0FAa0y2z
83mQFVi84d9RBu67WL19GdyELIXEmaHGMqafKvv+f2W67IevlX+UMC3P+qdXhlCg
qNOfZjYUDx1oICVvvoMDC4s8R+Ux3WkGfIdMEpqz4C4rbIfTTc4BYXloVP2BXUx9
l3B6FAOwUOGIfdAH+0m6Kpky1KI++8qPWDGOE5PrGT2cZsc0LPdLb7WPv/tKtgf+
XNADxDa3OLigMGzKdhObKrvsA57y/srvjY5CwRLCWEM9kW+T3nkEGpj0Rxfc31Em
gw4P4936zj0U58IOL4dHO92BVFrj0367wPZgunrZPjxXKnHrzRMQoA6vYOZcYUNV
HCs6CA4FqmT7LXpA6++mEh1x6i4a98zWyy89Pgs5VGbHxe2qs1KqzAsgSI5XSrfE
59FOWWiwIWrdb/mLmtjjSubXTXfBpZcUlCgnuner5ZtfveRCw4PlEudZ6tqUwQWO
il2U+q1JkBb45FQ1M82yiDcAO8aqIZqVaYAK6AkC+7E/Fgl0pQHS2WKeX+T/MePp
zpt5h9sQTp01YVeLNqKo3YliOR8tOcVV1s/Dx/YTUY1RfN6Jn36DPRd1eT7kUL5N
2kFjDjkcmC9PcBLqPXzbYoxeMAW0sZf0EBaqi96BrTNkaTlrsOUCZx9YEVkDjc9P
byEhUk6LQNl+hC0mNaWGUfxY148eKhkvlRC3eP2j+VeXmVTyxREiwhm3u/CD5hFs
bFZ0uwP2SemIhjFBRNyIGRaQsdI+tc6PZ1jy9omDxDBt9KMbLgViKrnMsSgx9Qxb
WFepZu9VDlNSA2hqv6ejhaU3yuLQ4F0zHXZ6FX0L6BZ0OdnIb+uRdeYSdbAQk27B
7NSfu2wAyVmYVhoLqPCqPhQnFMeXpVtPKI7dilemtNl93t/iWf4/DtV6ul+9fQEQ
w2xQW7u2m7DT1kUEhQdWfNRME8zT8hiOvgKlwhR2PI6RmX2hTmc/tqaIled/l26h
EFaseShXGYEyxSuSXiCKJzLhxM7r+S6tEqkRN9a1h9P9zMdwypE0VMW+yHZJmjDF
+VKWwNkf2+WrydDB/DOCFDECL47n1v8yLKbCRfowwZ0omcaxDAC9lmmdn5Cjzblw
MEsnXnWqH8WtNJHrg4YyO+CmvVXI0VDHR3GYWg1X6Y2Ty9FHRWXlDX/TbpsIe/IO
9UFoZc4QVkzptgvgeY3USCObkpPohcgfFB05rnx3vZaWaLkZ3IP9mIIAnxkVAkJU
TFxpXHL8rdTEVpt/ZLrL4qwv7vhPonpwzubqVzF8+D8v7mnLwt9U7rMN1XfVPA0l
CFqHuwAHXar8IUWlb7ZU5eb+Eftf47t0V2XZLqI9YCqfQL5v56yJpOxAlVKEVkZo
OrUqb1FxMN6lcE/vp1Ir2iAJar4DVRCr/ZIFFlnsPhmWhofDoj7csNIZRicOffs0
5Yeq5LMX9/o4XtY7rOTLC/hslM4fLkIWHqywFC7v32luuaPt3IcBQHWv1cb7zfEq
Cs8CBVRW98qSnhO02UkFXRQkwwxb9CP4TtAjWNqjXhl967Z1XoeLBwfjXtpjJgXz
fRhTAWWgpB1l+RM+O9GCBnC7ifz1jWuWQh25Y25KDNrkYbwoYss1lNDMF/2u0WHK
jWpAE3IYkYB1Q0h5UN8UX6rPEmsMD3In5artDlTMFPlQeOy9CW7aKnRrclz2ZX59
Qf4HnfYbQO/yWFPRUnCh3KdsC+wL6oTYoseVZuJrH0W1Bj467FYhRrVDpf7kjrAA
3nGCj6LuFGtU4U5ul2W64SmtqTcOUY8O9ce2WXv4I5iryKdfl0IBIuW8I4JMkxJb
XX9OHGkxJdW6OEm3jTdzwYIey6MnERBhWTkB19OScKPtkViUj3ri+fnuzSStPqgV
rAxjJPpz29ynUhcPnohWCQYjceuOrsmrWX+ZYiaM1YLTUMymUYKgrGZTpdX4gt1Q
+5rBDzbydzjS18xHZbAwZZchPA8QNxhz+nHGJcGdehQ2wY10fQx0+8K/1sG3dBer
X7r6W2IYuwYkgFRoUVE0hCB/zRcGE+EQb3pv6dGNlqc24w+GVqFcpByFJ6nvTBiS
6BQbgGwlDxhK77UVgIMuahnDyTBcHIB4gofFH4UC14/kJc/W/4Gx6KFUNQWq0AR3
ll2ttme6xKNM0kEHu5YvFtJrEr8QTBtKIwJZtycVjQRCOhh6WCA96UgYnnK7oqQB
n+qgHrldF3v8AMYUbtfxpxf8QVC7nU2ZaSvh2r1iwXGuOjDd8/GY2Nn+fdAUZSLg
EcZ/FYeaWyYgyS8F1DV4Z/tlRw+mbWDCTdigYqAZ7Rdm8haqwxjTyW//Wxt/o9rZ
I1t0/oXPxWnyw/xP7c0UPiio6BMPjubBYWnzkIdpBqbJaazzglE7YX8NgODg4mpj
yyTGqnQX/z2zSrGKwUSFBs7dMdM8dNhZxFRjzwordYdRSs6ixXjGhEZQzt/zBjVy
0NncR16+LpZOGI2u3nzkbOoP1oC2/8y+4regsLrbAiam249eMD3fi1C6qXXN166y
Saatm5LIm+8wK4ieEKccCdJ/Mk5vnylROZ/E2uv3jtOrgU48ZugmVI+B22F1BSsV
oIya8l+cPLXYzN8mhQsHzN/POW9fy1uSqsEsj6ySNrvfHeNvjgFiU3Tvxj65fSRq
iPp8XPVfGhJ/3iw1hgpm9H+Cc/1zKd8/fVj92eUjrqKm2bQXw+j2QYTlChyAbp02
dz6rBZz6VISfYZZ7WT/n5wu1leS1ClI0Hh29qCpQn8mKVSJ/PyOH8ROKB6XqGMZQ
4/Zr32P5su/qbQcoELc7GQC8Ejygy7bRmK5V67D2FRtcS6A9pRHNo8xvfOLt+baf
YAkppme7JGl61UAO3abrATQOGPVKE27RAOHAe9j34Fb4pc9WKYWE1slVsn+fMeQn
CeqmKsAnUiEJkuFnQuSbKRlpm/BqBVUVejFycYNsMXffBSr9FT5S3jiVIBq4jfBI
7CgV4VNNTHdK6nnuvkA86uAcju1ZCTKIne3QHdMR1FqoWuW2+92RAv1RN5Ejb3xo
qg6/u/3sovSW7UlAcLdflOQ7gh9Muq6DfMhnTG1A31WCwwc5N30VPkw9KRcq+qQo
Bf/uUJ/no3fLNG+y0ZySWFfi98QtORmEEnxjsk7NdZgC28y+uUaTCVfPd0Hcr5Mu
bNNtC0S6MH9X1xcq5KEgQ1tH/J1RL5MRhGagJJBg17QThcGiO51fdcnttF3W70gH
qym9nL2qsW+Dob6O6SjtEZraZxKBP7h2Y8esy8PBsYHH0uEkxZdqIR+tWaOIiEuQ
40dIRDHBqXkyP0JIVdgW0b+CMi9A/7MseE30DDiSvEWfp1hcnFHSvsQndKbPQPX0
yO3jiuKTmjt8QT4f1CPReRQrHzM1ytv8Y/G2g5QIjTDvcXDCZAmuyvFHMvb7Ygj2
5XTzNhuab+99qg4H19l1aql3RKQcNYuEIqJos55h4E7VjbC7sL0XIhRoNvvqFSaK
iRA7joBhU0/0Cf8rKyvEIoFu//6aekUP2DAWrJ+k0mYRQ9iC5u/n1Bm3Nvw5sQM5
CrtDhdBtv0uwD6BUpjzZPyIW1DQi23WXYKxtwYpODD4BVKPZFT6nar7yRz20Oi9I
ytupJve2YFR9OEoHJSSKLHz3ZwSw/qmQxWcSBpczHbaD+NMtI/KLmXxPmwsweZf4
vhXZYnY3cSMISZifhd50ozVMSdF6WG4sckc7ZGU+Z/Y24hh82r2aj8h4BDyU/5vs
B3xMEGEi8tN2nO74ctZXD2PXC2iZTjrWrVP4Yuk8DtgMCJpbbOrB21yUytdqw9IC
UMUlJesmm7g/en2pCjVZXAPunZSSLqsfzkT83kYj9tWF+9SJwcBA/tWCsJ9wIUw2
1xQnBz5nDj9EuliaeMUMfP7SfIOO3MX/MTSte9YEzSBQfw0WZGi76SwSrnF00uLC
PPYvvnGnbLJOdXkn3pYDoyZk6t1e4IlNmtRlALWrCSvWBJRlEMWXzEIW91IQaN2m
4RQ1m3UqKUXwlzKdmPdK30EeHfAMXalPP8vpXgli9IJRqAMBijEfKZKmoL+ap3OM
ry/6/HUz81VDCuNSc1f2eX8o0knsBhQVy3yOuLzrmIdcDs7+b6wB4xbJ5CsXAg5T
RxGGQzmV11SgbtXNvMgZHAghSUARiJIFlR8ZBWG2JpkkyataAANz8izMAyIi7unO
IdhFWkGHhwZwO5UcabRoR8SNMQ6IL1YK4G9uEsIQ3WZn9mnGbHR9seVK0+7wOiFE
xya422LdPPfEerfl5XStw8Y8o5nk3jILcv/XlnQXevZt2v1MXOGhWmmCjlogw3ms
T/+Vty3mTIoWKyaSDtiJpKE9FkdLjHkFbFauzHM59xqp5b9OYAYFNh8/0gpEOoBf
tpRJmR8Pp1073C6LKWFZ3tMYaZSxggrYyelVVdPLfhWOx1eybEtwbFWTvoVGxZZH
HzHYjnj0znE/n3w4xJphyyfiI3IK4Mn9o155kzrZJhcwMJQ0ITBuh0n7DQODkvZG
O0QGXlgNS5oBalFydf+D/umCPHp277U/lu7Pb7B/BRGYxvYarFV9FWoJdrM/ucNY
x8Ya33ShUYUHbBukgvZ5148B5cS37zUPUIqnsUBKHI5FJ2G5zyeEOqwzSomjAKxb
qeCJhRl450cXlql4dbk+8TvHJQvcLr+T5I5enOPSrDSq7dfoGNcJ1TaK3lvylnKq
/CuAo8NwBGf/Vl/S3yV1T8cHBE6XOEiDuPOHurrmcGFImbu8kOidIsXwBfl8lHKn
brz4S1YSW3GuJ1PU42fGGZrN0/6pr4kgjztm61c4CiGgiDr2m2dY8lgfj/Bu0SEa
nmpZF7WZUrWYx/Sp6s99zF1yErZZ2asZbV5YK3w+lb/HsdNG2wclXEpkIlFv9Ezy
fHY/0paIH5yC5yFHc/egjgIGaEjO+6DClIuCr3F2jT68xJZZmz2saijkEyWGKIoA
+fWqI6UFW/zgezWUqx5MZf8Jagr3KvDscPzfkcr+1z4L7N1R+Jwmuwq+3NXaR+ye
KbszolaLNut0zSBnx+hLcQ0F7MHjjJ9rtSAi/eLMwhijuSw+4TFUtXGvsm6bUjMR
EpO5abHvhcC+Ljbkfx2IClIUX/89ROBBhRxFtts4tyECrloBjIEEbjKytF62Umh8
iJXl5vPgqqez3AoP8Ri7ODTQ8o01x8CePVzJBzoncLJoAfDzT+tSwbFpfJio8OdB
oZXnQA8w5ETAiDavgbYwrYNRIT8WFPZic3ZZBLlMOllT2f4Ebk8KBhRamVtLNjcN
+KolaOezOBhLBGMoXVJjOI9SkbttbqUErbDkZiRBtF9AmJNOwOtb67eXgjP3vpvE
eFmRDRw3p/TS9XPrHHZW8fbLXaojWDKVOzEhikT72KN/oAOQ9Ku6nYviH+ykabYo
Lu9YXuxwOe8zAdQcWS465OT7GGFY+nu5Nddbbps5sJhjGboPReunUaRsTWfZOBBz
dvIZVFDvi9hWkTsdayYlmotNjtSjAk7kVxBayZ8lemywIMy2whRzGVzEm+59TE9W
lZygBBI11f8zq1Fzd2h5fJYyIS8aKX6T/3Z882vg9jSOWXZGmaj0QeX16pI4rZ4J
bX1GRkBUC7sHYQ6KiMeshtC7wNaGDmviHb/24k4sIlUwLmiFUeJbiEMxZJZSdUWn
m9mLDaXBj6ls1frP3eNJA7klvFET8fWz8ms13cLP3F6H49K46rhlOOTqXYnrJmrV
QZOazdpNxhrcr7ZOJgQ89R5mpZHvBpz0ePtLE7cRAbLJRf3XWogD59Q/jTuV9QBN
h+C8cW+ffA2av5/bRIzv1kRXpJOrCOEAyUiLZMZrDqlsWrB0oyihPdmYYc11UpW9
XP87jv1NJXto9m7ET3EeJrQhYI3Rpr3rVkKk/rcO1FliYn9zx28dwIQG1tWLOvj5
y6iOkkZAvkLVFWkNEI6iYzyXfz2yuOm/9RB+l/4QRwYwKV63JeUmb+1p9WJ2W/3T
lOggck/5TsQjyeboQRglgaY3/b/vanVWKbgIv5oAgiKFg1rBsP54Tk5doUB+9nnl
UsB+42HZfs8m23FXt4JOmwOrHWiA957Zxx8ikKAuAEsaShqTXN05jLLeSqLvHYAP
BTsP6103xR5t5Hwa3XcPARDbgkkhT7oBOy6NZZDd5S9Fmgqi3R2OGIGj7KG0YczW
DCqwfszaaungMz9BTkNOXYMqNKWt0981js+kv8ywwKBoIUqwFZmWapizqxuHhN+I
BqC4SfLDNXPUMlw/ZotfaHlchib47M54rEY4r8vH1f6M8miU0WWO5V5Aag1XoX9Y
msQz04cY7Zizq2lYfTbGsFUSXyJ8/DPHnn8uZK5TW+ghe6ydYDex1fPX08LWAZBa
JSwAM2aVsmlyH9x3Bf0l8Jiv5PmVUBBozKXCVeQBGLq/cFeI0dxNkHtIqAbZfzHu
Gnn3nuTKcOz13nFhvNeY93oh5O/tYp2JHwaSN9t2cu01qRV34NJ5YXdypJNyMdNX
qHP+tV9Q5exiXzEsiFYSmPu/4JMp3maAwXWY7Wjm1PMmA2HCztkeuc7UynInvnXS
uBNftiVOq1dKfa1VM7jMOWuK89PAabsLox8NZEpUkIzOVlsspbxxzq8lDaUfTEZ1
qTmZI+lYkA6hYiY41P60WSqBnvkGQEGsvWoYQrMeyMDei1epUZL1QPpyG/XatZVg
NLo9El9PhFIoevCHkDFdsho0aJvHxeJmLODtjV7oB+UiF5TSgtbI6Slr/w8wKWf8
ZrWLEtL88ta3fXFGDn3MDl7Vwe7kPF9O3Ua9RaPEgprfvX85gm2ODiIPz0WTSDff
WNzp78K7zvQbAfw5d+86GlXgTMTe2drFO01Xh/qqT/xeNhMIHWB5Kjo4cdt4eWNE
1PEXjbZafWMOeaHAk4fdxnEhH7RZZrGucuWv6pA8K2FmQEc3yhWXZ8sSbvCV+7KJ
rv34GD5RuTJW+HbHtuKYySqUpqM/pFqk0IUMA8wDQrDMAR9AlEK3OqvyBiYFswsq
BYSyOJurz0Dt6O+JwaVIAUlGqn8rnBdceVD8TrvUzcHlOhtpMpTEOk/Qu1f22WCQ
lIzoOgcD/SkX5TI7FCgQo6dRVjV5L19EEVNo6+C/kVtKRC8hUkUuW8cd2sTgWIoo
ZghLmAW75Hsk/4UR6mkGbLLEMrhVERDAaG5sdVfv8iT/96OSk1Ln/qBBYpwRzzDt
qXKtli69oTGO9NvuWtvXc0fWsQiE53zDBREX20TDOCbhXodV+qmfNxHCekyHUdqM
Qb2bLnAkCXubSt8NsyKz5rtZRoWGGnurulq9TC0IcmrE6y9gEIMnolD627MLznE0
YtZXDXWBxe2FkQd9adiV9NmQ6UL0omNycyk3kdAEDpoWRF3P0GNaklAM6T5iX4Ka
YreqSbT35t6lLs4P1gSCb1haJ2M/K36ZEJcVieFdOcxZ/SAfA2oA8H1usDKJDtof
iiP8bbtCaYTnjvvOg5SFJlVJx6BVBTKyKmvH1K5Dfw7dA+IJLpaBmIMzdZnPT7b9
Fp9hfSm0SVcRNNhPzXkBiGC7jGk92IQd3E0H//lmj4tTbZ6VVcZv8klh5z6AJlCd
m38HLg2Qny7rF6OvnaI6p/1SAHLvmYjq2EsyCf5oABVJFX+SKC9Tln7HRp9F4dRh
TCC1/UDqkC4z02+HdlqkmeGW/AXUFcmqVkOrRHwINOx2AEhsdeNbUMm403028aDx
i6GjAJXbuv8aL7ClZQasEnk+n1kPLKbhr/Zi7R8fM9pSbC7+2g4kdI7rsh/MXMOH
vXaXS+c9srNv4q5JgxQJ0ZFyjhchcpR2bLiX0gEFznmYZnvxdTfr75P+ga54svxd
c3Iykr0waEQhS5Z4ZLq5NJPyNigv5G2ELBfwoUDiN7DlP+AM5WmfereN/l1/MzUP
JoJsABrNDeYUsnMNvySu1vWhXRNLXhMHBwwu4cEMG7t+ZvMVhtuO/7KD/3R6P51i
r0kk9So1aW9azUY1NS91Dt53POTddjGm+Ry22SkbCf712zo8eZbZtg1IgmqYPes5
ke1PKZwRiqwGm0d9KW0eMLvPaOflhDnbTJJi3LLAhbhs16Qg9oJDxhxz5nG/SosM
q4NlCLkZWMIAib2FeKlRAvJRz/P3VnK99/KZhhfRUyuF+p/5M4LNVvIIuUMqGyxg
SBRPS6RRx7rE0+rJhoC0tvEeB73inJfnAqWHXJEqwqh6povUnqSERURp6qX9auMb
IcAlk/7g5xnzaaoQuh2V40apwGK56jvsSPWEJmbjWA5F8RNBv0XTX8C2zabhtQxB
OmgWZ1BIwq01ptwyGDwaBEOztZ2V6c/t3Rb5tnXf3RofEKYRAahi6Kwmso8/7Hj2
SV5a3MLe1h8s3UvR/yrgQwhxKNZ69Kv23zpCENkvtOa9vzafO0GnOrc2AIMjG7dY
C9ernMDhyFF62ZXu6W9NpP92zPcgYsudZIGhwhxKcrLcWDiyDpSDiCqNfIlUJWE4
P3jc+CGzCDKCyuLcXc4SaIWMyPl5Eo1PZ4mBdhslFkg1Mh2I/1fuvgMNAmociesj
5QMy6OsDQbnlA/F5txQJJ0G/IV9inPq+Fh57leHTxvtb9HL+B0zEyLIseB9hWfkg
2Vj1B9cCsSz5OuQ5h5tcuR2SiLIsaTDs5IbcAZBPciIHqJxWZfxG9pdxkBafdmco
MY/k7TDST+pOSGrsdsbgNEm0IYMxWX6CPjJ4gct4+WhAd8IWs+ZyYjGdyH/QQSPZ
puEI+LE+ZNp3/ZUYKL3NgmyY5AjPqzOcf9NPtKTaz+07ZT3jFybj56MXwTDw7RjT
c2EOA1VidnD/wHzShm+ETydlx0LRu63r2oV7RVc+EAOov+CCwz2YNzAWG54Vp3pF
vXsz5oPTb3YqSpwWIw1rg1cChqdGivDoHsbUDAlzZ/j+r8WwOw5WkaADBsVwFWeA
waFlQx/2do5GxvMDZ668ruFq4DS/1wOsUj2Gn72mUokUJo8UFpgW713nq5tICfuD
CimlIkGh4m5CT4gJkeYpa1neJgaXGqp80VAEtU0Nbdwc1Zzjji8S/mdg2+hGrMBP
5YgzJX/QUXIr9Ghs8DLZtkOTNjWNAzVyFx9JSRXD2/YwjSuHxNMck9A+4jN9LJPj
7+Hjbg0d8hkVMLhyGL8+YKF4qwR9nNWDZcdV3lzpEduE0wdppWCHOJDpyhMKIGiz
pf6BOp03XNX3U1ybwMRwpR51PmIvJUhwWAYrwDdDJonfkrYm7biPNLFOAwUexpOl
VctY020dsXXCfzTBa6imcD8eghEZvCV7AAN7xYaOqpVnXUlnFUa634bFOicyEK+Z
6Ev33hQpCbt4mpdGNyIEUcijPzV0o1YyX8O72NCf81ZaVEmvM6zsE1YdsXCyFEe9
dsiSw7fUpfm4ucAD3TcQHjz3im30sRABLKG/1aO1qcsssOT/2urXEoYdYrkRnoRs
9g/NthvPUoFno5dAFac1XKjNPqzQNdxqNjZluI+Oqwn0jE9LozrCjRjaE1R3kIFQ
YeU384vkQnoARKeNoZB39nil+2/sOSsdH+iNGHIYA/ta5KG1BNDhH6DDkxAZ0P2E
nG9UsQ+l1q94dkBrzQxG3fcJ/SjMxo81FaihFLefV5QVojS3yBQPboGx4SzOo5Ai
YYIArIi3ivgJxGGJq0+hPfrC+CtfN7xQWEM+t15Lgy35UOcfiY3nwjYAub2VQH8W
nVe13MMd3uet0HpsI6tbFk6Ap76tZA1dtIlqQCDxlVxZ4XrS+r8Y2Pna/dh0uCRG
q63mqdGiVWqPVnwFdUcWJtfIxBjTOO0nF+NcdjCblc1rQnZyrPqFaJKipFwrkTQ2
sn5VU5qqPkWxC8UksOzTB1ftixgl+QcTbWnNAeyyjPHE6cs7BDdsAzbYZlN7ClRk
SS/cFnpmYcNg9Masdxth4p87P0pFwr+//u1s1nM2nRfNvZMUVfiEKM4fn3jsTZOL
DGV20Ge2pquz5HNibuu1eWb94We1qVzAbCGv/KdKSCwkRVXX8vkH7uSVTo3GfzQI
2l4lhSAKBbqT5Nq+7hXYL+ibeeHM6tIsXRVqSCKxV6BJE/lgQTjK3OegLf/ivyY5
lKuJhQQQVBfkepdC4lL313Yj6kSFLUQWJQdRzq8Y7Rwf1VGx7lJSjgbbK/XypkB4
ngu06fQbSxje78mYuuPUaD/pr6DTyR5wUphKolKX+P+j3QRgeGLUd/+nrNPslj41
NbP8NUo1MsBAKYLWSl+LMU3gbocA2c2lZHB1/gnkhvcdmFuMzOuN8b4QZOOu1ZiM
tBXRBV31LeYBGc3BKEywWtR0djfeQqje57r1F4a9fTSSru6GptngymLC+549oYlV
LJA6wIyOHfgFUj48o3ZtFYxhxA2a7TcE8FgykVufwm17C8wNP5d1MdMt+qJbr3lr
9uXCoxfNgfoSMRO9wOS0jugw3YUra97Zktorzm7erjH9300zsCfCs3JGwr3tJVw3
3pHrVk0AlTbBzOC0GPFxR6l7lsYvDaPnM+lyNVFeawz79V5wNzwZxFrqrRssZjxy
TYEYbqwGwruijJdu67viStfR24aiv3MIGunxpXg8YPZrwds3mQ8cBXT5HnjaFiup
f5FIFaqLdmdJ2YuXOz5UC3okv7CF6JrtFxGQeCokgxubDD95QTVzOj20y0lsMjOF
GlyABr0lPsDpv9jy2GEbhp4nvNMr/T5T91Zh01x7Babvyj//9b6Dm6jr792KZrx2
/4s8JCKeaZTLHqIm1jCk9TIu0lWjZjHNaTFAgZzVZLnd11k4jQRj3ptxIVakxUDT
NtJPR8wd1F9wqyDzSnBfccLJ9g/DemPluEq+xczPxqCF61CBrHrDpkk1B41Oxxfo
o2oPg14KnxKliKTJuMHsrZ4pTM/GHehc9kV0dLwxwJSXb1FWksZNF+kKeLPJX5vt
X5EBCUOvaCO54NVFw9RCRNMIDQRYt5yN6rb0lxEimFh53gkUvqNlG3IDocLRZvl7
OUYid8v0H5HpfXkPzFzAB7/N33hjJmlVxK7sSEZivhv0T27cdOKjZ+iCPY4b4fAy
59+hGhjSj+2Rzw54puBXJ9zZBKHjbiycOOLE8LBxqlVj68l3Kr5RkvczEQYHuOmI
wz8zaAH9LTq4payrvrjQDNuY6ltDcvHtMQe2FEtbvqzP+VFSYwhicfuVWZv7AmKC
GawhjacU4XUPpZtN1/ZMUZlWK+Oq6ilcwZ+dDev7V6OLufhLp7vq2mDOwY7+2I+0
Tc8Kew+8Lsrj9qkb3Il0/+P35bGdLWKoCI3VAJrJFY4GhyjAMSIqFgbZf1EQKs7h
pCZFrycR0/in7StFtO4mA3Q/i8i9U0UDHZy6gwp8qnAOML95fnrBBbRwxDqHIMon
UgvNAe7wmqBQxfoB68V/LJyMtz3NBVEW6qiRCnroMBL+ARsHksrA5f4KIDLXp6Np
iBDbANttcIkB3P/Ghipf7DbKTFMCpQxcdqB2zhorC87B7vND9DzPWNjOHoheZg+9
J482ReuD8ts14tNIFcZNasdFLLAvfNi+OimZZEf6/42BuzFGrjE5IG6W/yEuZC3A
UfqzjiLiew66JlBUSgQtRKHnFFefWnPetssqlgwOnzCKzSibEeDWUcuEb0pgHUXa
9dGFdLeoAc6Ys1iqKlw6Zx+Q+E6tks+9KVPhWDMLr7iBEDa0jrNboUb7KkPl0LIe
rYimv5DsBvKNTYYxf4LYQFdDf1m1vQZLEj6b9VkQs1s8dN3IqUKvJhTBi8zWez2P
Cd2Jsze5iAB2xzXJjSENfv590ukyakV1tHH388caaq0FFPaxgoP2Rrzb7E5ki+iZ
82Zg254m6UOkgMk1rTnRVttJiGm2LIpJ94jxvjWff+/lOOQCV28m6CV+Efrp0cdR
VIwsivU3Di4gV6wNuU33V58NMkDUVZZ90gsR4AubnMiAJjsU/Wgs22McvjCXeqKx
jYj52BY+3BZk9itlFQFGTf/KGnpr6cVAhaYWwtyqf1nXTr1oVikxRZDfmESWPNGU
NuNoM91+17JsDxoidaw5bQRiF6Y8yqm3iJJnBkKoh5nD8glYBGMgQ6XnUzygozdb
nLoDxga9u9FpdiHwceSwdPz77vbjOd+MYrgQcbgsdWOz4urfavLHftRa5EPwuggj
vIDlv6ecNm0E23L5DnwAZKhTxdsOO3dmNHOGWQ7gua2S0fGp28czW8UKJbJl5iJa
BB78j1j5v3j+daarDCuTimZb4fXzorYPbTKdIYipmkAVQUQxcbFe/SoPNVF/6n0p
cJlgADWxX8QtmDb5DGo7IHLTPBeR1WjzJunn0ZAO4uc/9IGJjK+4xZtvbIDIsiyw
En6rCYZltNn0BBlmq0UPGX9O3CyvKWrLblAdIWV9olcCbUXTbGdJ/hHeC9pNDiyH
gEApwIEj3g8EjNeTJSrxcAMdlX/+z8sxFxZGeTfvc8hv17jFOO5/FK/aTWZKlAa1
aJLA5ioOslmwUwtx/JjmKWqE1BRmHLIsRSeUE3nUDerosBArT55h11/mqZrmM8JT
ykttCLptKmZykcJkNhmwl9uSLsGxVPiFk2h2JXm6zlTwTMqLNsHaSgNVMo71x3SV
ECSJ8s/V0j3VuiIhv2b9itHlEzOcYNkfS/R/DqWxN+Gkm+9w50XKHv2CUUYZkS92
uvb6BOfE6B8Uimmad9zup6CHkCdLmiLeF6pyxKVtj3CAFI/kIE6RkbejsKrVAAZY
BemItgbM4o/vJWHADBbr+ap4NIABvBHeWT6WMx8HPHfD8cWaBB7/SRmtDwNBv3rW
rSODyfBRaxsu2HFVfkjc9V/3RGXbv3S11PT6vYgpzGnBbRmFY0aWk27e0wlGlFea
EQQQwKLdlg0Gx67HtqCVu/JRlA1x1w+KFNYyiJ+rJ84jKH90VYjL9pffHB+xgXKe
yk/ToXxjaXtrmjnNesyxKjbxl0vGsXnp7NX5YxudC1RVneofNk08CKUM8W/f/ulV
AhZvYKb+3ZT8iTBCna4agU3KsVoIDPzZqcpxEa7XmoP6fcD9X/06xYZv47CvcbvV
cNVqEmaMHtKglTRn7lXwBfwb1QOZgzlK5eBppyvJzbHqq9cCqO/kLqx8atabPlNt
m8RSatilHA7yvumUEwLNe3ztvDKHS1a5s5ljIEM99Qz/HfuI9xhw8xcw0fBULhIO
2EUSMI5SEwjnHdQz4ff6R1a9yQoH6rebEjp8QPjEVqn/l+tYDN0BE/i0kwBNCArB
bCBLz6ofC9p/0IVZjPxwoc6Xv3zZIW0xyK/DCiUKFGPLZfqLKcbZjkhhXqKCyP5K
tRS7umLqkeqKbEIrmD1DPytCZ08gPwq0Az2As6JUI3Lo737atDeCt9U/BAyo5crE
Fvjc5tGNMZcfP+KzEcku7VF6Jl99AADZVB2ei4s1WvfzRhM4s00VUyOnK/1MjexL
/cMel8YZH4mAOn3wfAqPpz6CCD6BRnryTD0VmVpcx149EsGTBSi1z56orJ7bjwCf
eWpftj3G2BRF0ht5EDjPUYK+WsTLm1Vg4xjqbQVNVkiza2+G2+gLmHPue1+aPcYW
XAmca9DNimkaieLRK68HLy8vXjwfvwlrBOWZd/d+Bd8ikjVsCaS2S1jWvy0/RFVr
OyYF1LCNEDy7xkJtcymDGNgrMF9FnfFTehcsEquMWCDI9R3nVrQcAdmPkgYQOvi5
F/enFZrhCYrcn0EGPEIl49ypOGZij3E38OFWuxt4BqPtYpW8X7YLnVgNQ1Joj7i9
VY4qzERVeL0aT6NPA+94jm1Nn/RXjRmrnKKQEwPycFYGpzoVtNSwDWiPwP5pLjBC
PwqbmIcTOKS37rOrX7kyakPt8y6fimRb15TGKBx88QlDO849hYpWv08lBB3UiHRX
coxmiloLV8PtC7gIL8P+3Ak3N+7ADkBf/U7/dTQY9WdWCMI2Ln0s508qFNbQNzNH
EnszhEgExyP7SvUt8FguGu7hvZhZ+vgmdcU8W/qkmnZkSbjXA0cMo7vT6Fl2WtNO
lIqZN0VaVtxEhzTWYS4ReUAmaRg+zdSXrIsgtWnGZfE8RpEnZm6Kns1i3K6vgqwB
qEzwxEpdqdAdIu0BRndi6VkXm+VcDF6YjacG4y11bxCMJX0QkWg1wHlYTYc7UEOK
vTeoNPACES9NT4Y1+Qe146Zx19ps68pkEEuBw2wQ3F4=
`protect END_PROTECTED
