`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MM3bTwpfZktMmCpMjlfP4RcD9x2986Z61TR/T99U29/vL5Rmx5pRyHhpG7z8mJjg
ya7aVYD0rKFg9ouxHKYKFndgd9ahaI+kmhd4py9RmgA4LHgXifsM5hE0I6L28j8Y
h8I3TICoIYx8Y8y5HU4tBTX0GMpiYZsHH4uBvKd99gGq3SjORTILW1GX1++jnRMM
WWtDuvD5NmIJ2Alj9N8Rr6jCFKbwKDSF7Ut0pJFApqvSaWAoe0YHc405gWPbK/UT
QtX+KtUNAd+lPUdRwLI+B3nniQ0mBCxZNbYA9Gq7o2MWQ0aDMO6Y0jeBNe2FXCk+
Zry+DZpbefzPjmgU97VyyJdbXQnit8GpxViWB60ZbTE34YnMi5leCwPZjUpxClXq
kT9e+H0ik3ffH26sBAteq50YwNsuXZP6QmvxezvV1lhNo/tGL20ZEbzl3F14vV3T
PGWfXZ748vD4PT0GOSnHCnuPnXxF8XlhAiqeD8feFn7VcFrfOH2j5Sil/HdkaWpc
FJma+j4LOrKW3O8yU5Icjkpo8rD2+yn0TZhkHFdniq8ThJJvXSODM5RuJ5iwsuFB
hVo1+XCXsr9mtvI35ZFkB6ZeJjZ8C9roVPtc/wrrEMXW1YoFBJOaeEijgDsZZta/
bDY544N8LJ3J8UAGUK9sIGz8Yqd1Hu9CcjWPN9WXg6TclpsTipcwUln25D0QETwJ
ZOz0DI/Ws7Qbpk6u+QON3b7mhM1n7clf3fNAADhHFnjS2bft3E5BrxUAr2WT2Iav
Z1NK5VbCIla8hHbeaLB+oSEVoQ0wxoPIDUJpEwuPHZNCNdfIzlwbeQpw7saanLPw
7si7/P9Z9fNnDvcF60Qa8vPeiwVyFSeAX1rQkR2sf+w1+VkGQ6YEwGqujhXJ8get
GRRAkAA+e1Dfv/+RBdidJZ8aZoqTMb11/asGPFh67+qS0HffdAueKVyNqJWaoNuS
XNN0Wi3uyZhfXJ/3EF67BtanG9x6/AyRqhJ3O3GXx4XYaC9xFP6Fx/ZdUsfrwPrM
qNbGszejJekMBy5RFyO0J7N9sUuJXzSA0i9c8aSgP1Zm/1Nhjr8xgtpy6VmVq3+Z
0MVpz43cJie+mXHQAnIRF+qIgJ+L//PK7SUlmPN0AaQL0azc2hLanQXm7Qaoe1xg
5EZal5RLqbJT57yGOhPeM7y5uN7eS1AtKan04oNQ+r3AynkRbDj5O/7+qg8dmY0J
gulhoMj1D5NH87P3jNIzztrHnuraqIc1rGMhzQibyR0=
`protect END_PROTECTED
