`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTUqg1f0Tunr+5wn8urly4U+2/oN2kDg5H+nzGjf1cxdgbHznyR6EGXfcRdsOjEz
jTSEUkazojEnJFyjh524lT2+/gi65q0H6Vfd20JC81sNRtl2YjUoHLT2zR28PD2L
oUeJ34BirfxFvx5GQwtlgW9NMQqZK1Kz60dI+4a4mR30zp16e1UzXv3+o2+SXO/i
RDCZY9g/MyqYEGsr4dMEC12XrXo32U14C9kT+tqyX9H52131YEg2wBECGBaUNtid
1eh7eyxNREkfUyGes8fQ8QOfFh19wZAqogri8AU+DZg9RZK6tMBh87Z21JPiYkYw
HwlcTIPCHX8+jzvjgpeEQ8C0ARoa3dah/MYMQCkAcpyXxSHHqaXLarZnWEYXy5O/
Kh3rxeOUDlwUh++G/7K49o91WpdUQzLAWeJcApIeovaFNReVugYnG2HnC28kt1ka
d4ejHs3ZMMxgTSOqg8dM8DVBa8TvEJVLVxuMHjHkhg+4vf+4kiy73eSf9zPUQApT
Lh/ifMaIySThCJHdlLXbciYljnE3JNGXLiywMeu5UeOG9zUGeDfp9r+6aFh+nm9H
gLSgQCq2gv6WhGuLvLmxfMuW9HvrlL43zad3w3Ka1gEWD/yo1s2evKAdQY9JZ1J1
D2VgFHUibIWhVbW47r50YvaOEzVQt4gZvV7YhT4AXLvj0bXktnE55C0MMv+n/MDi
wJRLGfljCx2h+PgXHDWbspQgF81P4GXvfzZyDv/I0yoihNqTd+iAt66B+OoKNG1Q
fvXJ6BpzojicSxUIuOX7CzwwX0PFmBlHdYOaaT8nq8wERpScpsHnVl12m3KDkGJl
ZES4/C1tqux/5xCvXPDPvSQQXYEzaE9YEORsSgvEkj5hFQEiY9n6037/sZOtYouB
l5abXxVFTK+s9Anf8pNaHnfqQhulMKMI+5AdgHGRha6X7CS+BtT5Kw5tFkbqaQou
mMBSsEL5EIWie1tkFe5UX6yeutIul3dtxOtNKWuIhdAEtA8sRC1CzyNrwrcr+llr
CaBJRE+kcC09iFLXRupWDzueJ5ZewsOExIWwB5LYiaoNs3gofiUQe/YdSa20NDkL
fFDPLqOaslVGtXCWJpZL1Q==
`protect END_PROTECTED
