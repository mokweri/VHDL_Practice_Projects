`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t6yrt92bEl/XL+TPFjonbpttai73DHpw1q5MrmGg3P/TUFPiSLZTtYiMzAL09Vaa
rX8rM3Wz/Y/uqPtEW0FGHaIGwXDXv0vx4txUBafUpYeXq5npYY2jME6zG1VR7gPO
/duqCxamQIVmUhDXQJ7ZbIvrLJerZ3s8zpzjRDon8eSn32Y6c+iZ+0wofYQbCp25
+cM+ysV5WaKMZ/qYzyInyuUoMnEJ7iBdRx80wWjVI47AtpL8vC3pLYql4cWQ9s2M
CV+LVg2GbiyIuUieenT+CfK8yu+qxkff45M5AK64AbIvH4zPCh0bOxm4kD1edEKV
qnRi3UyELIzP/MIgz0ssqWro+9ouDqLeJgFpL+gYVss=
`protect END_PROTECTED
