`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lvSrkllXZoo0EQnRu1WgiHzb4rcfVOBNnn2vIpSrUXFjqBhnOl1JvHUFTQVryrma
Vz4ZaCnZ2KtPsrBkFg4PzOkb7SBh6UQDpAU/lKGhhabDwsSUkMU3BiI9rsmIuoIl
Qu7YuXR+b7LdaIL9FwMjYN4wxkuApOg26U4pTweWjQ+uTloJIL9slgx5WcXSsm9L
wvadZYaUionSMWQ0iaTnKibz3zLaiMgH3rzDfIZtjs/qbQjwrcVV33VcP+e0lbxg
MwSzGfgv9/jROnS9mCVK9JFJVQcDtKd+Jebsrpbetjp9fL5TvWyk0ozWhuR3u02+
VmL6ZnVi/GE3/J3w+cipV26UAibGUd0XBUKJ+3d+hqHcbGney8LbzJ4cYilF1CFN
Hlzlc7wI7fqtJHdDw7GQTkjD/s5rpNK09LeJz2n5D3N+32TpQPRZvuab+ueT/0We
5TR6Xo0htpK4UWZGxlWqGdehGE0rlA3dGwDYP/dosj7rPRPsBayTzLKNkrEVbt0l
0+Prh/MtOfPwX9ckK3JBFVfKDN+KuXHYSKoqEJR8Q6eS5OPW97NHmquYzIdcMuKj
fZIL6IYM0u4AfRBrmtPvcz2AIh8kEW7ox7JRPQUHzH5UDKQ+vBJWXU737w4QbR7V
ogU6cAspMSMDi9hqEj4YKauuM6Ne/13s6kT9lGWU/J2k/DwE3ZztSyAaTLKDL+1N
nlJq2OYSlckkXPsvCu9qh4gV8Z0TNq/ptM7ybrvzDZcOCVHZF09nQ7awKFDgAhJG
x3MWoOZ0aLSXEdn5iRBO13HdTD3kfEtWYLx7zwg57D59seCzl7eimLQ3jW1PRSiD
J/37gnZNAS/6/bjDIdYcaaR4VS0Xgu/TMTBcNjyHGywXW4BvywbVGw5/w5OwoJWe
`protect END_PROTECTED
