`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuNZyQd5CNXbI1g8DtBauvoBFo0tPkoUF0XGBE2JMf7LieBaXmbowObd9M7JNcoi
DL0Yd/BHK6da/ZHio7fiK/aUab8/brYSN0/TmFCGkadNPGIv/DxbK00FNMyOO2rV
kIhpU1iemekWsiC0TAL+m9ULxnblJGK8/WrfROU1DcB4nFicmgGYC2EKNE0dQj+w
7DGxkShTHYuQg2GwZeWCrufLAjR8a7rLTH3CORE/zMJiIaqC8E5J8qgkxlRF7G45
lOltDf/t7QfGmaENnYy3F5mgBUVLdL2DAWeOaY/ZGyqrf4QnTYEQNE4Z5IcSE18c
sq/hqOJM3+kydQAQNIMN3oZBlphNNC105fCLuDA37fNo/0ikz3skp1DUgZh36QBJ
EEDRduOCiW3Ez4vkFJCzniAQ3R8IMQ2r99hYjZyWbKNY4r6PQNXxUVxlYbCNe6/C
RtA9ED1ApgMggNyWxJd5AvWTT8exWSa4q8wWLq7J1NDNh+a63cACQVJ9NUWf3MnO
CpKo27yaiYeQ+V3ZI7ofK2C+S7ZHXfuAxEkCvCbXtUUQ3ihyy3HN+WSMtn/TOVuA
vyWc5NA8raLGd54H1u3D4/5zK0+M22Zee3+aU9gQdpdIWSIbuSJrQr9YpxVMw/8G
+l2mQN7dcPMpaJy8x1JuKVv8+Bre4oOnzkTLfJc0xPDOB4Cqs3ouNoVWBp41ytFb
Nxz/DCApCXPct9XzQiEGCb69hVbMtRS2+TDwfj8j9BCt6WyclMBTdvYIxW1DBi4n
dxeuSZWUGn72gnF51uXKWJQ+U1oL8odAH+MUMFs+pPEdYcrblGA6q/VOyrlS+iyk
ODV741UBtqKt/DncPhYhPNT/wTxkdW4IkzeOCrk+8SLeFzvU4+YBfD7m547L3EIw
AeeUC+PbjJu1WC2J7lvxp0miVKkrjSTT3fWMhF8cvRBL8Phvy0U68+SzJqMQiSC7
vDkWfPUc6n3A3ieauyyvyladBEd0jm9MiSjYRo+ejtyx3XMD+W4FuVRQ1uJmTx4k
lG0j+Q1ymVQwF3yA8TbzM2w7PFIMphOxzUnS6ajKgOh5OBIKVtvVEb2ltMSl8BEA
LEMz8h5mDlIuw4F97LWwbzW/HOvGDrO7Kdnx4YfpYkPEVty0ago5xWHbhwlVWFeP
93KYi71zLuVLl6YG0pr4GHDpdc2KQA2058+byo5RTtj+eLSB9S/UOeUCF8Z/l74d
gwNMuqt6653/RcxeKrSXS9vR3rLy98kUeXrpOEvdSokBk1gFYQOMZizZvNPLCqLV
bqBvkjSUGiJVexpEjeQXyouQPwTCRXN8MCS3QgHUjg5JC5NWAh19ehcPpkTjh4XU
F137zYmZcCQHNdNa4UAJ26JenE7iwQb6M1esaXbebBhCWu1d22UpyzrQb/mphoyQ
g5c1c+gU73XdUFK7hS9v98D/hd1tyQD46dD2E2Mnq2f1Bzlk6NOIcKWgGG0gD5EQ
`protect END_PROTECTED
