`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Da8uwDBv5M30sd8EK54eYd97Ss2Sjf/m2W3+9qpiGllZZlLrr08LERxVn/8OJ04q
hn/c0ZDQJawavk+qWlIHwS8mEUdYBhn1CUWei6YVDg2PEQfkmisMTq8h8vm49Qoa
HmpjCEo1t1he3r+3uDjQLsM9cz1INsMmMiC5lxRZhYCrpTTSlUiHYAmMus5IXU2a
dpuiXiC5YJ0Mu/Z4+7rIbX/E6rwDxltDNKGiM9c48TUEk8bg2w3Zbje1kheZGBe8
gxq49rcyxog+89mhBBo84EvvZJqBlpMOchjqsd35i3yNv6E1/SNTZAsdsD/A96Pf
Zx9SE72uIJLG4tKOq7u8Fn8w8LxK1PXYRptqFQZR8BNwF0X1gOfWEO6D3bkBGu4p
Vs5VPSWX/+mAikFys9bc7RrTOA61eWAl/2EBr/UFwNkHqli+frlUqCRS8M93rWbI
POwF6jtdvNn6FgmtcAga352FUZRiZMUj+BhhB1JvnZ7aDUYn31L6cZC5hb8EtSy6
t4BrGaBWKPEM61TFAe+U7Dmgh9CTJvzOTHNMwMZU2iB4wiMke8K1RjxgpN87bjom
HTtWg5vLQFLxPq9X6ICWRK+w2pQ/txyDO8z7K0rNXXWhwMSEsOJOhUQxVHpIpU/j
rlVUBAvdaeD2Crq3OyylMtFSwVWn9ziOvRgNywAqW1E4pd9w5r6zUPT8azvQp3nU
njuIMMrJeVrgzcW6FUH10SZ+1VX3l85lFItbeS3rUBwX9sR1W9T41A/gVOvlnZrH
UWPee87nbETgOnJc/6eVUCl61S+zE2ivPtyVSmxHF1SJEvTmNMH3nI5x7H11QhCa
v0MbzvmYU5mK4LKqvzWW6Hus2UFpOD3JBsR9Rhz3qjhPz/IPIKT9wOsnZW645N8s
D/+etURg8t4QCar1EFQ9gGf7PR+3vUGCsH0xMhEWsgzQUFa6hr88Rmd/9TvN5GJ9
8K3ApRjWfYDr+FkVBEOXYxKRz2iVP/pQoMlZ0T9UHSx4sxnwZ/O1JbXg5DINCxaw
vM3BVoUeriP6r/fukE701D7RmTX7EYULN1OOsZ5XKwkI8eq3/843D5hKsX4LNAQy
6d5ERZdnm/p7CpeJ4AJ7LBmv2INZNs0Pp4jZbn+uwtil34rG45tHctu3G5p2EZRf
1fmqQQixuiz3mpFu93NPJGkIjMkSizdCjtJrGzsKo1WdlbJV5O1vaB2p5hQJnezL
2XmfawWO5TQYGRXo7O0fJ6TzsPMa+Xmb2JO5YrrNJaGMbk7pZH4yW58exaujDB4v
DUqeiJhh2KTuPZaJH6JbFiu0yUmutO8HpIRmRhkde5etaYuuvw13F7qwsZpBz7fu
2kqIwnPu9KBebyE8BbiQ2EzqKK3T26tfTNFkSJilbdhPFuOpuTVmqHv8ClACtCe7
GOrjAcl3oSRzadjTBiMCKeket6t4WE4gQ0+dJkPgGXfGl8L4B97k8M6obvcaCn9/
jfeFjcNoXikAb8NC1PpMlfSmg1QXyvWw3LJrpb2qVseN8pPcZN1Zk1hvGSOJn0Av
HAqfKr/IPWQ61kVmFZbqAY/YQ+AuwDaZ10VFZqKMUPDS9+UzzkfGzTDoqCGjnM59
8ZgB6g0/OdtXiAwiRhVefpW2kCVgJjQHJosZ1o8rk4jfNNfI+j7d/gAuETh2kVeN
YFa9CMVmRn/ybZoDfYv5prwQITqZ49wJ2IM7yDWBZ3pYa9hs+P3PIuIutk5lH0u6
G/el5JPinOOVOEH70RlpO+6ABeIjI+DAjziRIcvltFecKRrprBc7mbXF66zC/XWs
`protect END_PROTECTED
