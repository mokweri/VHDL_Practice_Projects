`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbZ51Jz/WGXqn/WOviPxkrzVBcYUPd6Pn58esI7rYNaGEDc5GCWKaUzLRptu0ww9
0H98VX6cFuNYCdXv/KpHoTQ8RSDEtm+Dcy/r4iZqWLyMo7csFbh421T5jAnk5DKb
lqhYaxXZ9FISLbA5LbLwUg+wcv9ltsv4+/dBzp4tbIvTGtMil+8COIT3QezUpL6k
c9HgKLmdB6RINOyFl3T71fg2evRoIt79/IFvDtblHV8ytmrGKSznlTaFZDcl3rmB
YEar8ma3muzHoNAheogPKjKwoEYMzHyzj1rnqYBMVVwsDSuIT9vVWLrmWX5NXbvf
LXQXplwnS8uzS4cLi28yKTcSXed+/dfhs+kfRd2yq2PUJ88lxGZd2H10t5Lk5JJ+
CAuUuU84jLdPf66ssLAX/YJcWpZUmeNYExbv3iyLs5iwG0Ip2sO5LQlsgR2jQhT3
4jv4mJkb7xm/euOdMLlPQIlfb7LEG1KT1pfswgaxzBhcRFT67swPObbnVOuLadwi
+TCIaalhWOwzzdqxqEAIJvq0m29HvtAoTXPJpcDsvQ7/g7QYsvu/YxvNqSPYjHh7
QW0hhmPHQyhy37vYp+aY1oMQLbtgGJpODRqVE9Uvk2nFgMembl0KyR8tLWplcxPt
OEHb+iE1cQthgJCaRGpOFO4NY+OWP5KGJ+eRDWO4bK4so/1WD5/JQWfBL7KTj/dV
jmLXVmnPcEwMh7bSPzzYNu5Li6uN6FHCHLc1mbEeTHDlPV0fPEqAk4pQ0RerkVhF
SG+6CU0t8CU/p/VIUGEPUA==
`protect END_PROTECTED
