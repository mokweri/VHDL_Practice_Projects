`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUJ42ZXgRDpugLSr3lTONUKa9DlV3I6BEaop9nNEdSLqz5Ojzax7X++uQqhGKXt8
zr5jYYoa03ezfPqNMaPtRfnI0jIEtAPH0Gpi96EMCI0qgc5GZi/5UGU7rFUzuUs6
Rcu9tLJkIVM+xcSaNaDG5J9kLPqXNfU7Q9Fvoyfje17CBMoxGlhELDAfh0H2Zws3
`protect END_PROTECTED
