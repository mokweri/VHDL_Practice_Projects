`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjQDlov55QOKyfo5dqPqf6vTE9dXhd3eGbt4VNCsmOioh0x/K+f//t7wAUiyvKOh
GIUiG45pATWT/FeWfMCyUFcLU4dPc0tfnFFRJCSAnlrwLUL+NdPK+A2878zow22G
lxGwQUAYjWw+h4THV0iss15djh7wzlP70nOAOsF1fqix8PwpskjlhBhOdOQ9REDG
n4qJM2GMKj8oF4Mo1e351+ly2RjwHmDRqaJXpmCFmJxvYrEckrE62exVGs61dow6
KlybB/NlLuG0C2KzKuHDRWkQUm9uGDdI0CEoMTWQi5jkzSBugHpqFJeXAFieZjgT
vaLrWn5HcnmFbuXlPCzZzMAGE83Pfa1AIvQRfReLJ0yLv/wsGY6ckjUJk1wEKp8k
CfAnTk2y8i6JPditusJ/CR5aAHdQUpEZLe45iMUHrnDzVs86u7FEH6ypweolWlYh
hN5LCp/95s6rHRLJFYcsst20+YhY2RcT0WL1fBUUFlqRU/nYsOhK9WAkcQRrOQKF
HL/aUHDXn4QKwuhvGJNDYVUriCZNBObgtVOcC316F1I54ay2Sj8QIs6SKHB2K/IB
R+MhlB07TmMGiOpPMnxz9Kp/dSsDkZ+AFOB95Sgoo78=
`protect END_PROTECTED
