`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WJgN9q1wEWnCgvgEQuvsD0POUIgbsHgaxqFfsFhUVVecna1sSwM5mwLong3WSZZ
4s/Ou3ZBq3aifXbRw9I1AMHOaxpVB0BN8Isplh3/id+bLrqNvL7en8s77ZoQaGi5
BQPoFT+ECmN1awcdAXoAN6FvKeu9w06FMlHUTsMA5bDY3gbHr1h65oRLvOU5IbXn
2G+wDxTCVhhEiWE87Kn7c9/ZNYx0VqbaxNhqlVXOzuGx7/kK27Xjlwch19EHzv0v
YVD9zxjd8ZuvAU+E94Us1n66xLxEBYux2Fht4irf0Iq4ZbkElM60BcSgbX3LnL6J
zRByFmIg+6yarn+Iaqi/YHiulA23felLfeTMkFgP9kvEAYHp0rwok6rHeDmnYlwY
MDdPCA0AaO90kBES2t5Ea1eQ5+9FG4CAynXmg0T3lb6zGPdkSgKgPCG7VXo0/5c5
aO6GgGoJi0lxd4hJS/L2/e2+iTivmeeNNxoSvTB9R+vushU0X9Z8iwd4WCLH3fif
TTwWGAsciwwoH2b+rjpS4x8RCGhv/Yg2IZne9q5WE9wUqUzIuidmyPIrmZ5THx9O
gB52jiM6R5W/wr2rVm3vy/jogZrSqPK9Yom0OAl7S1eXlhbiTg6zL1AZdnqAYayC
1jsAe+WXTtgZiai0uN2g7g==
`protect END_PROTECTED
