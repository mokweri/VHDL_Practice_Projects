`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTTGL6G3XCAKh6gal05xbxthmwcoAjpGBvWVGcK0pv1ONLtdF6v+I8LJcetOKiNG
KalBDX1vY4H63EOCZWqCE0hUqjom23Xu9HpqPG/BOmLqYNsInshwpfebCb75KmOo
3PEN2o48pJ5QmAwscq2J6OATOlUyQtX3IDjWOEwTezGPvgHi9S4Uq6qNr3jFETes
z3BCFZI2Ckidlra4BwQcboOqB9LoG3I89u5TkIdsBnmfsjtH7ODh7xGp4rMqbZLv
ZJtXBY54/O1Hqa+eONEjkjCX3yNZGHgla8wRrTmxmM5puIgSVWZYIXzKTRgQcgl0
lrcpmRn+o+CEXo+tkTJyz3pIz4D/J/Yt1H8ynx8YpeMrkhFtkl53pPqE2ePF5HyF
XTcoRlUjaS9UpMvewQ3wdQ5JV4Ap5tUuY72p5udqC/4endAdYvRA+3CCjvEMjJ8e
k5QCIB6Jb9YT2kUZBiSFxLuUladUpJkP8xWjYUGCVbk=
`protect END_PROTECTED
