`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6JjFTdkojIt/yHtVKdAhSqOZAWhA31X4hqsZhDtPREz93SfmgTa3MKQ/86aM+YX
GOte4TwK7dY92YuuAipmCTGLyNK5Cd1075G/9K8uzwOoY6T0xhSXHB2hJlW4/10p
4KXFvOsD6ReMhEYhe2Cydiks2Q946liImXQh2jCdcPD0epnzlW9604+N4n9CNbl3
myAyxv37WyNundBz/42tbYTMKr1FVvgVTWYaXGDRjrhFJWUGC4y2CcIlzRpk3QY6
7i5TrR/HZOqKXYPb2SOlpGMJPW+5hJbDXuCyVvEsLW8Z0WPEE53UKhT2dcs8vSz7
jIf0o9zKrU68Sb5WY0RzZBMDJ5BHI0CqEdzoeZE0GhS2hoFK/CWM9bR0F4Lp+y7q
dV+bm21G16Ws3BYPNUa8YV0UN3sE0Zj+XwFkRQPOdBU6GiENCA6Xzf9fT7MtMkBB
rQG5Fw8l0KMv6/zNile5Rn10nz8zi/iuAmJYDu05HoO/xoPZmRFESgzRe0feMFC1
6/Q6up1eytKMA4W2aM/TsGNqKt+va/U3hirDfG7YQeq9iZLxZfL+XL5yNGcc8wzy
S2K7LtmyhonDRV6IIYzUNx7lNZXjitkwNng1KtNbzcYPJdVfxISAUIKlgifiEDhR
OvYecBr129LfpbpkIz6/aglrsddR1tE9Pw1nxNknUMtI7E43a+VR1MtgCx6z6/8w
6YzSTI8LVP7RNUuj2EWZt+2LF+ufj4cgQXODFjDFqjU0vyHAlVTdGJHBtN5sgMTd
9vJHlln+StpZjT1FIQjoOoIedsmDwbQBBd7QrpxBm+Rw+HNceNpI2JEXC+2BYmjw
ZD5P4y/S5/LFu7d3ydqWEtgf7p9m2YuSu3UVHmbwIQdsFiV2LXydUAYnNYM4w9Mf
/RGAL7yKpYasFy0RSqIQOj/HzUgJNACp5tYdyW8+GgPZ6jnAYkTAiXwhE8Yp6DLu
DVnHTU3pNAcmcMAUo+YDfEn4XK1Sb0/E3R2RaF3UivvAlbaROzI4r7pvROGh76Dg
FIiqrvy99tWhFBP9g0AR5cxdOJZkZIXn9GXfpgsBKOlP/W5PAMgc++SRZ+FcMrhf
+1RX+yH1DrZJnLPNTwLX9s9w5byRCkeaG6DP4s/GDne1OrnhksbTryKrEe2uMSS9
hjirrxAP5YQDdcSMq5ZspNCXuGFw7VcYou1AfDGrJLvvmy8rG3NbQS6tx3QrgVtn
4ae1Jlwlhkelr9M1Ia7MjqRZ17CjEvloQ7bnDT4n19zDXB90B50ZWvmMjeuDJIi5
q5sj9+lOktfJ5SieQhGruvqZXre53npdc7e4PwNKa9MwTNSza53cm6UROe9k0Z41
sipA92H07oONMDdO66+9O2d028o78RxpZd7Jl66yiMz5GHC6V/iiff+F+Sa71Ie1
Q4XVuCKVEBTMK8CjKeyV00VlcmrzlWNcxo30LHKHbmkOj0XDIdxDySgB2t1wGy5g
5TrzBBHXO2y9nIMZjWEnWz6C/ymNYPrGWKKWVBUZi8k36b36i6FUDTxx/Z5l5bi8
M25AL1bEQXnk/ynh31eE8tbLqhrhArJeTVX0aBa3d33yrf/GxOwAVBu5OKttliGS
3l6SAb4rMgURcFbEmVYciRqvDhCR/ynzffxGvorO3ApIvKcmCepLyP/wGF1VGvEg
3XzOsh2m4M4/VnpHJp9VVIIglZtGyVW+96ESnQFixq99H68vR9EBj9e5J5Hpnmmh
FRiQJPknWwS5z9iD+bjTRuuXhrBgAQosCOD6AXzioSi9gJZEWpp8BpzSSL3iYswF
S1CEmgQTjSEwkJr16VrkiuKfzRCjSVJi8ueQLxvBfssQZDWSQbs98z/lD99d4uOD
HNLr/KszY4D2XGgYkiBJRnTh0rzuKPATTMdVdQEei908rRYK6e9Z7pMV5pkaF70X
CbYCJ/IeKs0nhhvgigu1CqAgUo3kATGT1t/e+uYcf1u94ZWeb7SxZQCnIqqac4Is
uAoSdKRkybPT21KZWV/ZzrVTKZILuyMO86r5LGnr+5vfGCxZ6Tfu0tyOHRqKug9W
/N9xggIA4uPrrgzCMAkf8eCbDIZZPdaVHW9M6rZbHkb/W87RKtqUPH09y7dxvfEF
hSBR72ECVrJtHx6E+hKrJPBCgCYPf0R0TQEEQUyqIjiEknL2/AXR4GQSaOHy6Nh9
Phuwr3FvnKk02sDZRvTFxC+Qb6CT+jsgE7UKy5DLKFpKmHci7ojSaLkeSAbcy7DV
Ww1WNcWMhcZY/9gL32Is5eS7gG1wDFffwOCNoxTstQjqTMF4NYGE4QaeOSJr2jX3
kQiIDuITbnbmus+cAIxH3eZHkxHPOSp1kB3heBG6jgMzyPlhbAXqKF6mpKPbSu08
0UMlYp6TdOQsEFsnVXBH7dhmKJnEtHFesBMDUIDLVY1NSTsVBA4dub4QL6EqOf3X
7mK+osASST/yAVmbwrumlpCD3hDWSYQ1Q4IJty0Bgug/jlejfxiqEMulwzyr6ZpQ
8MJ6oLqos7GLw24omrLHHuOK9A1KO5x0EtR7P2VZD0hzQDwlU4LrlgRu/bnp2QHS
AsI0Lbi0ov923A6vX6uPi18A+y02K070YjD7QxT4HpLB2R83N3Z3KYgDrczO3NaL
Pm+ROVwNWC8e8w3lYMC6HoriABWydCHXm2jVs2jVD+XbHfw7eJBFL+m3ljJcvI8k
fnvyruKUHqIEyiNmpUmrvWjO027W2Mp9vGaizXdCSUFSshRRw1VOgzkGmd2T//uc
Z4PG/dSGGZufM5O6LzFLjtkhyf9R4WGgJABQmnbB+3QiAKWgGekYJ/gqAyHq/nuu
0yzBv3Cc19tZdTUuvyTsUdqLlcC14WHd5f/F9eedHa9kWnJbMHyE7s/PJEGHXK5A
`protect END_PROTECTED
