`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNQkZghkOXqvfCyW/j+OuqGEP208a5yw50afIZrwgSaql8MZSD+/wy3V3+fmNhIr
3JH81aVmGLACtupP0M9L+vvqnxC5vCwAEsQHbYYeZrSW+AnjZtqSFmFWJbYdH2Vy
VsSCrXmxov3eYcIp53dwtWLbeWi49eRwGj9vnwU+s9dAF8NCfXXtIq2STcmOVWbv
HTybD1CsjDfpqRB90gCEKIVAjefSOB40zdYuRBtqRPTDxV+Q0vOEy9ZDsDHNTg2d
RXR2nt08faV9Msbfb+CXUKFaTHjYj0bdSr9IApmvcFHOsnlsnXxBCcZZjmYDzsfJ
5UHFfaBMpOr6Soe45YsNwNlWPERJB1XuGoMmVDenkShEL0Nj0g9b0VkLn7b3oMOE
n4ovwaN7cBoLQVeryznHWhJfsTq7h0/LULiyiPUMQ3nbwd8s2bGMii0uI6DY9Q/H
H/P03vpGgkU36KVTRfNNNV9qEzfyVT6x2PfVA3xjQOmN/CjvFT+XX3Xi5kCNOZZm
AXXEDuNqrXP0PFc5R77gifnt9Yqz77UpZyt2bRrhDwyDJCH7eB5Uc7FUTvppuEG+
kpW2FaJ7BH4en3mObTGfHVPoxUp7Uvknz4YAZ6KMncTbAjkFFR0fOUFGBYP4OwnN
ElqPY2Y+TUDMhfZN+CcD6kGqGvrXykCjBhBt/u2lknDk4olgCXXr7n+szMTCB4DO
m6YvpLi0aro0xBNPhWZH3aXtGZfF7juNU46oCdpJrty+FBAw1lLFLi03oFvM9LCT
imSCwUzsAsIUlnvMgiHRvJbMij5PRp6L20VOhjUSQL1IM5e5u4RNwA4LB+Osallp
0x8IqvzUk4NH+CMaxxQjaDd0V+16W1MHqVxB3/TAGKBAE/PXjNa0BdgCLy7GDfvL
JCHodlp684hHN01I4MpdhP9gEvT6VRxJRy7PtydhGJ3gOS0hhZbKO2W1mEVRahC7
JaQ0dsVuv+Cf64HhwMBKNnr3aDDQseANpkaNLG3NErSDuEf5zgxsrnLQI439hsV4
tBlTY25fnqvOEkRokXCrtacqY3kgEgEqy9o5+GltZtlIm/zH9ZS7/oqexjAhjI1n
PiFzmjzZ47pS15sYF02d4BtJn86/zhk1Fn2L0YUKb1UsYzctsfOQcLhZwDROjc/M
6R8ViPnrqIJXg73hobqjw2HCPjvjgz/Kj24nH9+JE28wIs2swhsCHMnPcdPQ08D3
LlgCOK4uzLgOQqq9/lsyP6IDzqe/wwmJ+88AgVZvSmlynaW+4Bhy00YdvT4nryhy
WYmSu3tXOGswwxQM8SV6JrgB5ZCscjvF1OAXH+42GCTKdGVGFlyN12/eIpOMvzrW
AEDJzJ9tNZKGGb5Pnv1HCRmPePsitPlcjyNw1MzCygEKfa/XJPQ8ffSDiFHkDy4E
axtppWrY64441RAf2IYTmHFPqlhdoGWwgLqJ9mAvCtgHU5/2hJYDWeO16je4tjmP
swmiUkADaPOto9Osn66xZGeXNWJcDzkGYW1xwinVeJho8t0yTTBmBOR5WvSpMC2r
eIGDu+7QGocQMqJo1mzJSEssMpWUi4bgf+f9irtEkEvuRva/1OXC41bAQcdjlkp+
qzPscXXATwbidRyDqO5u3O45msk7FgWEO+JS8Lr+rNw0dAcHQsEgehvA+PNWCxaz
w/D21HNB3FxJSgAUrhfzq9a7E/5lKYu4I6FxEUIvrJYSOsh5pHqK2RE0/m6HAXod
lgekgp/l1DfGuWn4a6IpdJGy1FM98k+oGvi8gVIxfUQPjfkiPb4KK61i3FjJU0az
824Sa81Px8ucxQktbZmQYCqY3gQZSPwl3pAcH78yGTmQLKv8sumFZgLX05he/VXC
ptwTJ8MGRMxzNW+BzITt5sG1uxiVw66ReCg6e2TYPfFokXkePYLuSPWGCbqmefd7
fBZydQIBAt3eEm28D7QOBUzX6bTiS3d1YnRb1wP18Qoa95Tyi+7ToWc83LwcVaXL
L+lUxnCf9kwV9LtcPcFDJeK2a6/2faOYuxAiFCDree713ov1izxbcKsjOyaYj61u
6iB/FmiGo3guyIPr4gUssxdhCF8dL2VTPhZfLggRtLjSO1xtfqCVnKjYlf50tCpN
9S6kDRZUa2hSX+JnBpq3Bxsa4QKWPIoSUr6hUnyNX32gK7I4B/dk5fdZSh2AJgiR
rIZOzG9QFsitPVR3fOdKM92v+nh3sb1qjD40o3Q9fI4LcPPdlcCHICEjpLhcm5cN
hvZJQTPMDfx0f1BlGXi1lEb7YIYuCCOt1hjp9Glbl9mpLJqSfwTyCOvPkl7TgO/t
aKSzNTYHInAKkDx7wozTr/kDJ9sd2uYjTkGaYht9X9oF1HkyMULh94WOtp62tWWg
n2YnZBPXn4A1kQdpNcGqHyCbVbMA9NkoaBtj1Y53yvKHj7I5ygraWFQa9JrkMRES
J+0l300idzi+kOySgNTs1beWpICRLrnqXXhZ6khU6lcC5lmybVnSMJtwvy4/hUp2
2JM+oubyCFf3muQezwOpfHPiK8K9mCvu7h3QzASkM9zzHCAfAxo9COKT1cBWhhjA
qgKVTCC09/gAK2iBejrSIEBQwdmWB/19vX0WOqiH7U4Qrr+lZTeE2aKzaw2nT57g
XlDLARCl4FhDGpxJVS5bW9/XUd4Q2k3xO9WRQolW6IBqprA4euiwI5UZqEBQdsKJ
EFVXNe+DCfbWy0c8r/oJ6gDU0FY5ELTX+iGkmKG4Nr5fYZBoshyY2CLJu4Wknz7E
DE7X7eWTVIQcz3fts00DNomy+drn8jqdLlnsL5GaLTl7IQzNYv2gJkk4l6yKCWTh
LeJAtQ8NEgSmeq7Zj75H5O4o7idBoO9U1lBQOnYuN4wkw5OeVTcivxknkUtxQ0zb
YKRb2hRVhlVAzQhAfxrkbnThnlgxMedd8WUHz7y20L3PBYSyUoqzCNR5rpPfc9D0
merM8Kdh7hQ8hvPNlEE84LROiCU+LRXufiDTerOt3hYcANpfrJ8Wgv8nviK20rD9
t4DgfoHpxgzjnBW6FeTELIhZjJHu4wse+oOOM2Cfds7T18F1yg0urQEN5d3n3OzX
FTH6BFgDMKUYytMlJY29DSKV2pJRhf9YKYV/XoSBzsI0wfEp33gVlLH0G+0a6UlB
MlSmMnHcabW1wLRcJvtCWz5w2t2ZvWYXxczyWuOpSvdGYr3WEXLsf0npeu9HfNGF
f8jNsVwSnvi68apOA/3wezI+AUFa50/rb4NsIFFOqjnAZXrstcys7b3W2dpcCgYb
f5OpGRXJcIklnhNuR+iaxadUOXvY2MPqczZlVvel7OYq3We/N9jlS6emZF3kIoub
XaTWmvFZmrTAycdVQw0527ihzC+yIYabHXwVEHIUElhQdNfTr43dXsgYVjsWQJpD
KHHJLr1Va903epLZVXjR1+YuJJAh+q/4FGu6Aoho/7c1/5nmWxh1ahaZbRR6N+G5
tgXy3d7bQhlJlAryXUJPNB8A4l1wP+7CwlGpFkXXNRyep/dZ26eMmNeKO9HLukmZ
uQXBVbfww0tX4+JnpCOA9Wgdqlk5bIjf4VAlpIYyHP37/M8OOFwZmv+kixRsr7s0
nzTnmgk/L0ai1iilkZBtns7+FVzZwMeHo4B0BVjp65/yFgyfUs2GLsJYeKFOt9qb
TdfAVH29Lbv0o9sH2DpstDhOHPuk3wc9Z+vwaRRDnPgjo3JiQkCrYMJHz+MHIIX8
QnxdkmFtBfjRJ8ivNTf1/DZVMj1+VnW1hbiWl4dIgs4eJDkFKmwX1uRMirE6vSko
rS8sXvvhQGvJk8ZIpO1g9PUJPXOjhrRF5hwCCDqrZpju+1ZBTVyawrbT8ag9gh2A
DJO+5t2E2BgG29mECXTt2G/u1/FFA8x/xrXue3xfEiVjYyn/GIa8l7r9g0LVadd9
hqbJRJNsvcd47Nz5UIae+VTygXT5WhckzGYZqQLSs92jgKl/Xtt7mxMdReBxgWht
EkYGXk0dvlcp54ac1QOjZEvlp491fPV4Qs+D9aiFASAng8sXrprcMH6KgSXze84m
o52ZXzXSY/hZUz9fnd+Q5i2QxByJIw/lgl9Vx80ET0TEE+Hx111tdMPmiKquOdyS
a7YxqKLgBPldjzHo9TzUc2wnfrS7QXFn/sgfnSjlpbnncUggHahGev9G1eLAi4rL
hdSVsMB2hA9NYqA41nZHpqBKo+BAzWh4Jf+ZfNbV2oFJysHQcsqpZdzyEC0qCH/g
pQF11fPT8559nvFD55FYcvCAmulQGErA0T7R4oSbLVJ+cEthbd52MGFMVYgKEeJC
rXyo2/NhLoNUVEUWTwuY+L8JmbKgosH4qWyzXN5HYFwhoyAzzidqrRgmFAbsq42v
NKxp4KfTQAMUpfu7UvDS0H0is66VnvmkSqNR2HI62YxiIYuX07ZaRP0h1IR7qNZ2
W/CDNtdML3RfjCSS6VdI51wobheH8FwlW9s76QDMGWmB/u9LyusQZ/BQbTf8BC+S
3nqwU2nQJKaZ+hb5OWgSmwJ8cOBrrux4gjdKN+NzrhDnzsz7WDY+eMqnaJd4Qmo/
0ZzCMCKQgebL7vZSA4OXVMY+tfO+DKQ/+QZDIivLbU/4MHjiGFVG3r+a9efl+U8p
U+P0jrcymd7r1UdkLrA6PfqzSvp6q6yLCtRSSQ64kjoJjnozvo7/UtI+iWEqv3EE
4hjZtkEIDx4j3ZYLZpvs8JuuJBBsG5Iz9r+6xbL0StjvsgNd+tgt/HpvdJ1qohnp
7uKo8J56J/enEnua9/xILuBKpWIcxZUA4c16k4kOYu/M1wmAHn8D/Bn1SvjiGxZQ
i91Ah6G6zyykhtp2rAFDQB3kbLTLzwWXFwv9p/wt9g3wYJezHJ3cMu9MWZ/IDOc+
SctwOl1TQbWc8MvBqTIQvwLNUq494odksKJ0nWOefY0+FKXsFp3FTLcNODWijx7k
ayMnMgU259xRkY4lUhPA9th7mwgDcF84wvxfufrS3JyUj+S5K6QbCBxFDE0+UHgD
HBSXkqwX1E+cyCdFaR854Y4XleWjMTlbPx7nmUSxQCDM9dBFYUUPKFMP4LbBDG++
NGm//7+xT0S4akOifSLAe2Z5AVIHbYKlo42tEwBaSr3aprC6V+lxp1Ic+cz61FE0
PsnyGz9WDQaoUnCWt6MpbVve4FqZIf/9PFjGcuVOlTZdg7b1Y19B0ew+DFteEs96
YH8ApU78IT6pjfkUbuoz6FbG2ZiDa8MrJ6yxYGBfZWeKHhm4TPHmJmUtQbeCZW20
Dfs8XOOrJ+LU6R6/suBI6l2g56fWBWpLUDkXv95J0zPZKR9rePJvdVabOt32dCt6
wyQmeBRIp+k2xEQ9iHJAkQN5qNgNI57W+zqe1mzggjpM55JqhKg2by+1HdPORqUY
fDDQJpALfDa+S0ZlH7Urn2pySuhP86v2jQyegQZXjTwB1sfcCHRFfhvKWB6s26ki
iNRXhFtCbniorV0df9LqU+SOXuZL6qLivBeMQfUU+NeC5hXPm7FuEuWcpWuGeS9Z
CIew+ekj0GiUTJMk/NArV7VRgTzHxB9GLTKB46ZL3ZXJvDfVC72QWjLbqQ0iN31N
Kh4Bc3OrDbfD3SMMs/pcd/JiOX6tIGqa5ihGdLolgjhpUxvtyHigz1oWj6psXuaX
bL/V+wyF6S42Y1kTtaxo9BIcEgqqISevVABJmuPrGVhxnGnGi8hcyrcQ0RZ3yf/H
OxnUl6z+UXlv7MlOMCEQMOV7Uj5W7wiFaNoVwse3pK4YTIzcVFs+PIFFHRnK5TzB
aEML86X8oCLlBE8djrlAsvc1NswrEvygFRMu/xwMRlmEkufiN8oaVEdWUXdDj1Kn
BzdeVZYsJCH7M7OzRu8Uuqkc5osX1RNkSct1j5cjB8yzwK22jwzh33hq30zVLwUI
jCYXnSp6qKqKVLgpDtNjCFeYLg5tyUA4vEQKz/bOZvGmCLO8zaqOLKomrZDwmg46
Tbd3qxBL43u+5VHLyMgJcQPbg9SAhoanWhyczvEUZZiCE/BBQOnfQeSf8BnFEdBv
mZak+o9XpROgsvRYOJIaA72E2ruma6es7BajqqS5qzsEYMnDygLFHFB+zrQPhFur
wP5HYD95jS0Kgi+x0YxD0kxum9HDphKKxLvtywK9wYWMqdArQl1+iF3oA4chL4jC
jt9/HbBl6TAwA7wfsDAQx2d/Ob2EhUTOdj6GApzYSB7sMBBBTFWVUdi0WWBZHMeL
hhRw42auTut9x+iYAF5z0JeEBhQV7IYI9kBRb98iT3uQHZnA2YIPFiVizluPnM3X
+aLUnfVjl1bs9eoTmegRqQG8xgX6P5aARypHQd6C4ZfKhy6moznIzkXqBPbsN9w6
HmkK2inuOLMJvT15xgxmWkFC87CJdmx4YWX25rjjhDqnf1VzvvcCUgX4aItBlOYC
IjU5baEyMMajOWRaO8vyZdVcLsAAhvgxhXAgQNOBlL124I9ujb7jpYxMNDxtD3Gt
3+JbT81odkse9dNWhdjRI0iG4jVAYDy1mC9k5xuJCebuJSh/SMYc0vE6DnK6aT7x
t9gUcBNByE9SkVOaWG2K09cGHAGWXUDK52niafVAElkPYVFoxHMOlsdiBmBS4lLt
3ac/REgmaT59j02NYNecntTKHDB5chwnaxX5l2qOL3JkeAczaHa1NiHosC8vE3dp
t91DWF//Wj6o2h6POUFqivzZCJrzdx9PFIb8DavTHW/PJYW1SvViGSdR8n+v/NAT
w0m1tFM5k5MUqDLpskQecY6xVa/mgNDfi/Mq7yLKwMj3UB/jZnpN2FhQbbDchbxa
1QCWZ3HLaZmDN92rBVvXJofVXjmScZcDftMFp701sQWgR821ooszposGxyz8KCPc
wtTtxV/kFbiA3bHts9PcdexKcAqBBC8DeVIIYzduTpVZmyVQLOKauNpNJ1uEvaEi
nEErCMdvAZWCWJmABYI61ToUWOMwQh3tbqiW73dIK/w6U5g4lM/X0JDiFANRjF0K
F9CHval8qkwGaQaC9r8/LM+BaslLb28NEh2aJNutiRiq9Vqud6S2vFC73xvuh87F
81bQZSktKRag+4JxJ4Z6QyV25+/fyNpdJPUQ7TBxn98geGlcB6gJ3lueczbPyf8a
Oy7khpEnbVOdumkPEp0TQyXnCwNbKIkKhyZxUu0GDxRxeSuXQTOEY8LJLEwaqtfI
cHbwJGj3Ewr1GK2vvK0jbjBx0JueMZnh6eEb1Z2RhkIxbNyruYO3euzHbZp1Ix3L
f75/xwwZF4VlF1M4v4n3/XSG3p0yUqSGY2R1Nq4DVRfN9BJfnNmyY3wVCDKLHt9h
EYV8O8oAkDQzDIcb2WEkbdTKHDqR1ffx2ndqsu6CXflZwh8XmcXJcubQO9Rei8i1
IIDEo+bwW0MiX3B5+h19KGEid+hLjjb41FfdZi2PVaAi0C/2KlZUymyMURmph7d7
Ub6PK7hDhpnMIMsQHJL5H0quCsnk4tv3zgMovHl6M3xnPRFy69N18jqo1/p3O6Aa
MeqR7IiayAH+ptux5hue1NI3S4lZbWciN2BYLCx4/eXSfG/zvCvKXgYL4cGrxwjq
tGwqJ8QFhL6OY6El8RRQtc1pGb+UN5VLUfdHhhC7JSTC20CMOIbbfk2HN12sekW5
ojbpHADR+nhvwFjt2P6k+HuDaO3R0ONDdqBqUntz40ZYy7A6uqs++aF73mPpAGVs
fGXj99EBHBBEkh+gGzeiIULwI+BmOmb/3m/3aMtnKTvztJAsVAXwyciRCOlSj1Q2
WkiJxPou6FNirzUirUhu/XboMYEUg3Pl/OmSVA/zXkWdAuA3TmF/kcd/+EHAC1F3
nmjmDda9P/07ID5iWhiWXd/aZYBabG1jEnq8Hxoy2kx+XQBfCaIh1nT/O86vpr7Y
mKWdDS8LpVmHnHnWgIHnKWWRIQXDXf8iIpHVVK+pf5p6Uvl/W2iuNhPNxD7sVwKV
hdsH5Z0lCfq/RExfqcKwmIIx2YhGGR+IRukPvwM42/ZB0kv6Y8yHht8s3PqScptW
WVC8Vt/PG08V+kaKNXiG5pr12UuNxtkbXGzapLkiA5Zqd6t64ddmRTjmsDvOGGqX
endzQv95ijKrHFozwbQEdXmqhR7ufmf9DezFIQ0yovN5np9jnzJ33jwCNKrBXsNF
V3QdiJGZq6wsjIktosZzJtcrS0yV8zncEJ3JsUdDeKVwiGtpOdW9ZlVCmJA9tqfs
H1fo8Xc5SJMaTXBcaOoGgWdo7covAz63464y6WvXV6TqJqg63KEkq/X3vuwoL08Z
F94HtOPtZ/5meskpm/W9e1K9mtXRzeAZO6P4FSWxaaTIZPS/sdOA2QQw1kGyf60o
Flw1WY5BTD2DweZeyIjiXywideAi6d+A7WuWKCDRPpVsDKSEiVPrjviadO42/+Xx
P1Du6l2iJP3VV2CUtCbmogno2VuuvZr9sdbGPxEVPN8aIYyVRDptG8Dn6Kll5e5U
PullTWULVlYyjj4E8o+cDC0wznd7Yzk+zrylmTMTq6SgtdVAk/3697lFMLCzEwp0
OZarQebNr9hBUM6PgpHL7VN10vrTQmCfzxrYTc8AeU1Yh1AL/mKtIUb42HPSH9Cw
8XtllvGRtBJ2TxlwpJgaK4Qmg3DraPdg15lk/Cm0cff4sbpmXhKsfaoXbaBY5f6Q
EaYmGlND3uMvi0iG7hEiq5DZG5onZkQVvwS611UOjgp/tZFWbsukOO/WqPXqHxJL
0NclS7kWqyEokQsPPvilkDOI/YEznpTpUJH9eZhu4syypoCyugsNDsvwUV1IN79/
I5qS8gwM975nCdSCLPRLqopfawauBKRmPsQCZMZQTbQxKNkQNZ4h/KQBMoI5JBaN
gx5lo4h5/8g8L1Mxpzh+NjD9DsrvY5s1hfa6LdKK2qHt/0zx/PsjEz8zjVIQ5+TE
E8qshbMs/ZU/uwUbnorhvJ+F7EFZChqHGQvPtnHsS4hE+z4ewkzZS7dY/OvE9IMZ
ECbk9qCtsAtyqWq++xEWW2j84Bizg47FP9X5zX7/nvnCqpXcg5+s4rh5B8N+mQ36
EJ7Fa3cfcNsLH8xLGx5ZD427t232NeteXUptac1hJyzqMET0EIi8Q1GmQyQL0PRT
uEdgfYYF1rsGeBDKR9DirMvALes/MRSohFXfuaBY/42gVm99n5GzW8cGQsyYaGCn
RrZ5ZCmMjEbjD5rBiKuR+9Wgee7unkcRw4hmyZfYfwQBcZuy4hxhI0p1poMdXCgI
sg5CQ+eKIoxI9HBc+R/ZWhQxWut9IjA4JWvKEeobJCAH5vuA3MvewSlKjIRzHSH4
xLLv6T0Z/LrHqefe1S+Y4mSYGEgHWWEmLdxa7+T0jqAJL14jhPz3y8vmI+ZbXpSr
A2P/0VDzbVIOcMN5nCY01VLwgyH3dFiHiG/aMkVGqoNeaqEB5faaA8cKKMrNvV0g
NuLIkNgSIDr3GndDHMkTLtwJiy7jfsmUucUuYh6k4yRYOFnUvXc66uryf1dLTkKX
2eaUPuY9+zA1Bzo8dt3jsnZQGjpT+i3dAZKA/27xTldxVfMyy2VqsBxngCMHaQmh
GvWvgsKuAQuPVsFJi5HpuqBcgZ0sDYZ284U4adjJfhQMBGsNtSIRsPwsz8Ey5G0F
MEjKobo2+ycQWdM7XKuYVUFQqqpTF38TbWZj2ZNovlJHPYLbeBGYwB0DUzPMxJTB
rYwfYbkO29HX4o4C/M3tnRoigkxyQ8LeKM3PSZ1Hmb9RZgrBBF1Z9E2RujTnG3wS
P+7cN7v/EtRUaEFLQ2T2a27MKSJN6KMkI4XvzClYjie8lnftS2UPEaAfZklmPVQ5
plIzA6Gk9/i2nJw1UDtnW6EW1V6QQ7xQ3PD9NXljWyz0Sp2wy4F9zewoLMi8cwKD
AXZdeslnM8QGHiPYkrH1tG38b4625amHYsT4ZTLV2WJC7HdKcmK4lHBqqYF4YBAU
0B5tJaPkUMqupkifnWyQFFsdCrRPUgEYacYBX0QzvVDm3wwfNlNEn7gm6dD4KNny
XBhBOlwgwJCmOiOkIEIyrGBrBFVQWHrziC6v7x9w9LvjiCNswE6dmzqI59UoztOG
BaiZ8wNET3Mbe8PoQIiUkEv9xqeuQAXqr1bh7BWVH2nY1vReF032GbX77u2ACxon
c0ERzoLP4jQBHzTJ78m8CK6/wlMBvlDVW7WtzUyHQypyLAQFjzzW/Hf9gx7SZoqM
AZk+WoDQi68FP+xPD3TEcmt0nbafjSaHAl2k6dW19a56k3IygilcRpF8hBdS8m3t
HTYO4UJVoLoSXuUe64U3mkh2GoOdSNtH5AkOTYAdQVgDdhyCesAYNhEUs/sYWnbx
PpLE43/xw+/D8TRHPbNYMxTNJIuwIEMjDbvVlYAM+tTrj9M9T4yOhBqfqQ62ENpl
1UBaicAXJGDgDM55UbpaDhqKRBe6rXuiP7XKLXImKQ2bdVMS4exUFlz6y1h6cLUG
YLaqnUBz46x2c4rmko4b8qu/k4q1dTRr88e2eVjcu16fh4vyu0smoZ2UKt6/Vop1
vIlFqISu/w337A8liW81df+OF4zRskxA7cUMX4VxlHx3U/8MQU3ZoMGROjy3v3pw
UY2NtN5MydJDuurTbWn8OCv/Qx1jIg0FcFP+VwrZ+7UE0eEzavqLS/tcZPzRMTHX
9uYz4cPftI1gdq2ttMCZEoUAIOhFm6vjRXFTDfladCHv64kf7wit5LJpkXI01HMD
0Vbzj8BClIvlLoB1FEWcwlb/QHgwSeJiaAFS3gv5KDVIJilQk63e9fh3fTBmsqln
CYyJOktrDEIN3C05aVNKdbmw364fJ8k6H3pifhqKupyouS9CRuMS+Nzsc0of6y6B
/dAqSjoja4Uw7XfqwRkR7jrjm7/ATgVFIemgzAmLH0ov8FBjaqmi2P34lDgROzrK
4UobRvDfeRvx63cl1cJ3pGy0uRVlgs5hY1YV3VAW9yZIU3BdGAkt4YmRr6919IDY
j4/znGBvc72HujGdkrmS8kGY1yJvSr7E4JEv1XnGJ5lUJS69g8FXJ8cV9OzLVXVo
pVIKlUY9OutjWJDeVha5N0dzm7CfSLqwB1cyB3LOgKEyT78i22oL3XR3CMDMov34
kArDDtPSDH4EA9ke7vDYCngoyGIX3Lw7xOVLHvX5KtKK3TXL7fYLwtPFkTCYGmel
TKrMEujgfacW9+pG8AUhq+vbx35VfxAaVqw5k0h38nJfw4x2u9K0eG7yt8oU/jBo
mmSa/xXIxP45LI2KVsezJioyxD5F1b7DuU2R59qJhu1leOVGI1TF5EAmSuXt0MKY
7yeLgujEcS+dx1SyBxaEVrSbhQ6ukNJY+EbJEaeQhchUgBNXtEiTiHhjJ5pejYcg
4zUXr/5iFVBt21W9JJHqpzt35TingJXmu4C/8u1NLhMAwVXOSdx81Nf3ZNA/Ee6c
EN8eoIYUvWsuoC/+VK9bg33xzqZ+4MPzWsI/M6+meYNE/eE+81krXYmddLiZfmSe
ivHUAsAAuAJMr0ho28wHvZGKl3wvKg6zGLNHXHe93l8znNSjycqYTxwJ9Mq7oaUS
27W+rT3xuG8ODect6spZGSVIm2fvDpHrbBWqwC9GTs0DyxQHOpUSx3qw0Xl/7HwJ
KG1xZVal30/XTgAJ9WJHlpxDuwpL1cMWbp0gFpx4dAZ3X6LTsTYknlXBRZNjGK2W
Oxx5fcPCZeKMEIeZy0t/+z7dAqJLNMNxMq9JIPEBoVefmIlaIZto8s01ciBwHQUU
ArxlcfmzD3OgCGXUvd08x3f5SDWI+D+nLI2L/4Vp9tQCl2POd8Sg5TtAS0k42/bS
kSLcXFVGNmASHd+aofsdZf0nMOdZ1LMI6GP/JVYkRExlp6W//bvD8HZ8T+C3g6+O
ikJcDpZtfjiRbS0Fd/uBuQND8qcXiD9JmVK1l0geo1AYFv82b/lr3vzzyjzLCCJD
cXuMJqfrhFK52y7uQpFLCS6hJp2waZdH98SA67jXOOJuTrqSG7WcCdO8b6wrJbw0
bLRRIRpIVQB3npHxJzCTDUuxTZy5rZ9Wzo0i9+ic5Mtz9nw9IrNpfvT02DmvX6EP
RjFiyXEootW9g41D6DO2u48uKYv8PJcItqLUYbPL4u2IlNf90AIv/2GJdxjCcpYt
NCNi0bnbTmABU6M8ZLbcLQmUU1HGeWOU4Lkjzk8XvgjJNfYODYaIuQx+6C5v5svQ
Iy7E91mormbFzkS9jZwRSRi2Nu1p1yqCYoiMd6lacjaSlIDiAKY/sTzov7eu3NDI
zbWArrR/qJ4T3spnoiy5bJMopTw+7oXccFxKCPx3Dqmg4yfw9Fv1er6FKgqSju07
AuitFFgQgzyFk1rvr6GBg2aqreFQH04uLgRNwxDs+ImDaXlfFY+CjTE6o28KdD4u
8qCxbXFLzCpXzliwoJ4Jyh1rg+aWyZx6/TGdAa81O9ZXo4gznrH6ONa7Z2V7yFGg
5z5JljEbE95kX1/YVVX4LYmtDFZ1Fyq4nce4CIJzVfR+Zsb0nlImE9+O9GwJbQvX
VK2Ejy9WG9v2eOf+r3ftbKNZpFa6mtYW2K8kHburmpKfPZdYEVFz0eOwJM+SraWR
NhlNakG8Cwcm9FZqNHam+M7b1GlVzBfeWP+7VSFQ94BSAg1vHYOYYJ7UyQShOCrh
WjnZJFe8dG7iK7w6KGaNN8K7VEVA4LFVCdLX7CLgIQQ0ZNjzixnMvh2G0SoEEf9g
z2Wf8PqYXowvU7Ch5qNM5L9okowbIAr3dKJNw6aweuIFNd+xUFrT7j5R+/sxB4k/
2G7aqzkp6Y2WnBC/3hZfiSqNAKWn/k5TeE0uBSplbVLrFD8V3ZtzVwFQGsgXAMdO
5U3VHbIthmmd9Xept62ouqDMVaWZnv4IeBJYQTaEtQUw3yJoj7jf7gVoFVVejtMm
ci+xNnXu6hqGf0Raslq2sfY7NVzeJjdiFPWcQxtS6+QpfLPo6GCLi06O6CtFwpmT
98PMcTduIw0UyG1dVCPRw33+1xt/O1LnDmiGGRHpsAMweFpeCNv9fOviQD/kf9uv
Y2B/sUnOveZZLnc6tWm7N3ZFhkORmodpdKZV3dzFapQCoUzfOrBi1RjXuDkFTk1W
RrxDet5yg96MFsH4j69peM/RV5aaMM4URK3cmVGZMdehWZ+m4UiIO5AHRbjh4H28
MNUOwiG3yeT8gwz1nVPOrnMf7JrOS/zJ4FgUaOYPzpG0DdIeOLcwL9aHH1EpaDDl
6b3sSwyr8ukw4+5FQj9yYHV6So3QztjKvsRYPoOs4DWN7FDcAFDehQ2f6OzMBq2i
`protect END_PROTECTED
