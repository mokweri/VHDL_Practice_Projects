`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J8N3GmmTh8px/hDgA72vqT4yYolYyWDLyM99tszolFZFSkC2egxedPJSU3j/y5Tn
gFpEDmmNwWSoiXx20PleGrFU8p1S7XGJA36Cu67CArqkjGDSwKMjzf5A6Qr6QKRD
SS5k0Nq00jP1AYuiOM1eJHu+VB4UdoHJiUB1t8NlLz3eWUx1fFwzYrtralDdjd8J
tAwB3FX+XAbwRMfDrw/X7ELpwhgoUjNxJqOJm0+7T/UGgHYY+cFVRrJFhG4odrks
p687V7yJFIrYKOIE4SZ3sM1zUUzKsY6/Y/rJEdmtRJtd08fthKpf35thZywM1w8N
0LmF8dhJwMPvtFaNjMHc+nEmkD47ikgSk/XgzKoktmnGfcavRpNC6CGZkoIyzZi0
5yvIQ88YMdwYXLlmMuca5eP8O+t6Z0w2soACx2qRkkgHWl1gncfFAMYCF7P2b86l
dCPjxDojcagvdSjlFhH045K/9/icXLH4RTOYCc4b9KgegVA8+CUo2sOM6BlA97vw
N/jJhm+/OlpgzZqmhkDnGvr3QSQpXkIzQVQdhCNEwuOwFKlEh/Pp3YIwGwBwztGj
lDaItGhlIEfTtjg9aSxDtrzcChRhq7zqCAcC11sZyuJlqUHmbJzJEV6mBVTxUVwB
su1mn8mrbIpDzHZ/qIY9Fm0qDLp7RNU8u5V88Vkm4KiGNoMcRFkAct3kSVOiXiz8
Lyhor2OT91td0d+j6IRMzFkRyr37lOjZREMHo9/7fDTL3IGc+mQUxax+kfvygRg7
ynqXMdfmoErTBzcykF14/P0he1d3NA4vK9esuEIvOAJk9dU4S6LmFyrjdaV58E4l
FYth+Rfw+6bBONr438QNgn+me/N1ubc5Bw2Deix6ZNXNj7p+NNklGLVhfdTFZtq0
Vf/DTzBC4f7etnaSISeD+Q1QEC+G+AWXeExsUC0EFpuRK7tYqSp2MYmzvRvkBE0W
k8ucXN2KYWzJDp74lMXDnuBbiDtqhORhsfoTymg//HdDZh+1w/M8J42gGYYO4zXm
MUr4Tk9ys4tLFixth4bxPAo76aRQEylgiQe1CUH7h4U/JtmSyvVH48reCxbG6ro+
m7clW/5YwHeY1LhJhmTPCwtZzw0+2fqsi/iby3NT9a720QvqU1r2kf8DX+hP7597
blOAjCMXQ8zYipWrGBVKXjvmNhNWmHhwFRmQws8PpA8oKl5bS0kXnFPy8d29Hs1p
GOzp5fBsBVLlfYtpALCGEAC2MUAv4WstpIv4yuymjXg/ApAJ5gUpcIMWVGr2wvTh
fFs6K7i7pUH1uJKLnUlPoMJrYjbLeLo6bLPE4WV4S2xc/OsN5bkw95j+OUFRRKd/
ZGZ0U21RzpYUzV+5sNcNdG1pgpd7/JWtZJzWU7VG/HcPXHuhXJTNawG7jg4Kba6e
5XUY+j66rwg/z5IpkYDRwQn2j0ltOJsArLkCWxDRaX29tVJGKZDT3Rk71gRUWRaC
e+FNyvSceyRsExPD8IpHSVKMcjRIv+tpvohxs+WayPO0nUZG0nA4QR9a66HKYRLf
zuXzcxXaTUFCLS8IQmKrAF0sVnmaXKWVeSH4hgrAD8G8ydeTqRGpgIlkZnHSbmuS
TXem8+CFIuOzcYjd7bRc4v3xqMPFGAtxfLr08mK1rrlZ6t5xAejctf/KTqUmv4Dt
OZCnVYnvOTgjlgOl5PUTiILSsOMs9uaVyi4CevEPyejaq8pDCWIWn8Ejn5cdiTuI
n1QMpYCywvPPxkbIQu1hCg==
`protect END_PROTECTED
