`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xZVbjKKRZTqArlrd39IhJiXaogQrqhPXUQ2wFsQLRJyNz6iLxhwRHwnP9Kb+GPVw
GvxXkx9a2iUUIANMnRtIejmrCW/BE7YT4HjjcJqz9kzYrxSjdHRSY4UzOZmFhdjf
NEGiyuyWySiGfFT7EjvEPdTNZ0VIrxVkCJJRTDbu26vVIvt0im0tnGteHKeZGVK/
EeVMqsjd0kg0XOqAPEgDgN8Iem/02Gkh18+fdDlCPUHLwPeXySpXNC+kr1B1jGEg
v13jB2LdyLw1Z4Lzw5ZwZnpzjFu9n6aJ4nwJ/C+Ub7vU+nIe+Cka7fiOfvohS6wS
gBvzLsErnRiku0YRmzvoyoTjPUWXbF2d1jzufAOQf4ecjb3rQhwHDgphnbnkwWJo
NsDQkcKNBACf80uqdHTF24kRnSA611iw0mhWyPl3BTO7D1CdZOEneqihMXWOyA+a
dkoJ0qkpcXQOgbCl9rY1nNTHd81nTtgRUlvYLLvBr+0svecWolYiZNoaTJqurr5i
yDGbQWXlvFEp/nGISHU+JtQHZb4c8CfD3QW6SllwD+O/k8cmzNGneSyjaqbYQrbl
zc7rEVbnUKITrhoDKBhYkWfBJJxJzKtXo0qB37XtiicMON6YlHl/Vnr851W8xnqq
sskRnyNOwkAqa4I/xGUezCVb+L1sZIkwiSuPeFnYGCN8+CxSJdS54++mGtnfSMc3
ydOBHswuHY+WdN5Ot6vUbkIujx07AYGQBczVeoc0jaCzCejokKsNj1w73kOlnprL
CwtKjSk+CWbOI8wjohqIAMXqA0QOnz9IgH7ijtS4TuYy5tJoe706IDRrGTPC5VwZ
KhYLtJxYCpN5Ic7VfqNYzdpZkljuEQqlllDoRTYPkQAbofzEI5BM7GRM1bH5Zndg
1LZ1xM5XyymRuhkQURLPMayGxaoNJfU623roX4vPntEIK4OBjWFPYyZkh1tYK/3S
VCIUeq5W3nDsSRYnH0Hr2ZPVaOFQPvRJvB+rdfC7UMQVDJX//SIgbHz4NDDfg00S
P7QF8zURBcladOGOcBTGrWmpkhYWJMbI9kpEqueTFBYUtgAdNwhCStfQxcHk2WpK
gBMoH5fFJ+ypGKBID46ZFFi/ZHXvrGXpv4yOEd9Oai/aA1dbXw1s6/7mp8QqN3I1
kJtbx8Q+I5igzT135B4MAkVbscsG0MPGY99KnluvibtIbntsCJk8Tnpxzj595ZVZ
IBnP0279uOxxdpBYUwW5Q5hucDf0JKIZ7KUOEOEEyEs8RhdUVVw7/uFTy6VbVlhv
vwZAPQqJbluDIfHhb/qTsVAAF0th9asKByNS2hu9RkZEJwi2zYwf1lIBv4T/wPD2
V9DquslYLa4UnHxMwkU9dASDluF9y1vDzLryQL47BPm1i2gH14E1B3Oqq3IvqLLb
ZZfKHMielKG+SLmeTPNGep+kmdGdwqCchXJnoOY08KPV6EeGGgBCfq8CzS+rm2/P
GzBw9KXgNeYD7yZxkeFSs8bksVnE4F1uQ8ALXAZXMMs2I6sWBq3Rv/RyaEhiS/jp
+YnkMVISOuxyitxv5jDRiINUG7tBlSLDInSxmr4V2wyZtqtjYDJFtF4n6G89WSjI
9h7Vq/9m34NZxXbcoVhbZ8QpufPOT0efGuZhDfN3vDLLRZ6vuRnEo39JU5up6+vy
zA4xPFzuwGx+3/Gu0pAMt8CEgHNhg6AlFdzXFIM0ETKKabpsrg5l9gyJMHjchS22
rdbUXdnWBKhB9xEj6Z+LKuh/mdcO8zqg8fEnL5JAVWPcBH1+LAGmEREHkzTvssel
WSUbfN+J30v6a5osnItc2K9pgmzN7Vm/iUy64ZnDMR/HsLsjnq6XT3/6QhLo5Emg
ZfCRM9G6umKRJIm9kJ6IzJ1LHGvSrIl0t0q7jPnaC92QHMNSbB9oHYQ2e/+yMVjg
ym/lerxledB80LJtRLG56CVxNzHSskBj+/J9QDYqnX+miZVYkv2F8U+EVCVnZ26S
HQV/Gzq7JNRFPdorvAUYWXr1nBMIxVpEWIqFwglIdyVzKbxS8YA+9VtebZuV+jbD
vZQAD+jsson0ThF068ZMH6+keEE/wg4qrod+avjySvmICqlRqmuc8A/dlOgpwtMu
AHq1XkIWNgt3uH6hQLlqT3LKu1MTeTiSn13t3aawCP1zwUNQDKNgrLLb0zEcz17P
vkAy4bSJDWDlinz7wwQpZ05b8mAg4qD+pXEFp1Dyu4+RG1HRgVyQ/mr2X7dAtvPL
yg/ADd4F+bbKWVcZAsfUZe2gIVOaWgv9E5XuOXcyM6QksANsVLWEw28fgLDDxnYu
9WrD04RPrGvD7f20Y6lPuFAndN3D46SkiAIitoGkBF/0VfXjxVAjOLjOoXcm3jim
KnIxKq0aPQavxal/OMCs8C/n2bHKweF470HECiZzg/qaK7CKvYL+oSU1DHU/k2fn
WwChXXs4JXbUXNANEIqz8Jy2p2ya6j9u6N+3qL+B9CTRBtd+f8LOUvojDRUX2eE/
clQrCBNHcidtraAlm7DKbiBkhT/FSuS31W/RRnVx+LVCuQWCsnoiYiT8xgAczG0Z
J/4iGwZ6ol3wKF1PXrHL+HPWDVMHFt2Y2LAaae196GOH/HAi5VpZird1qvkYOvca
HczQW7cwJ7ob3OtCjoZgqjuyD2tkMvkj91MnKh/3Bt+fl3IVpH2xxw1bf1tX2HT6
X5nkGwcPIOAEpEZbqpk9QtGPTV2XTc7p40XxXL46uEwCpU2hWGb4qmBjqZUNejGY
Vo3ZVLRr1Dt8tTDMMY6x5+RQ/tyUbBLtiFX8GE14w5J85zgkBY5NfDKHFXu/6rRh
4YwuF7YjCKqJ0nGFqlqjogEogGZ9tD7ZZSrmmTrBVZSTVNraC77C9jadzjI990Sa
dL/iuqJ3df6RLEVtN2++yjIN4MHr8Tz+pq6PLTrasupz9qkvZRMCVt+wnQQ32Qf3
BRUhk0iLa6GJHYpvsyCVd/WC2cXrTA9B+RbxpdzmdU7JhpS+CyF1jkUmQNfVkjjd
IiBFQ53h4nt3A4IN4K2we+3DGThhuu8DT/3kch7e0vTIjjhgpNaO5njG9GygpKRR
daqbgyU0bSWRR+mGAXX5aMpUfunr7WOJS4C0ICsDvWwjR2TdqpfQCafLha40Qlbw
wyFUKiF23a8/Q+DkiBFb64rxgI3KXy8k+ViAVuo+QbN7Xa8O+/AeXxyAB2Jsnoof
M87oOUp8wPZFlY+SNrnpLj4OfJLLYNhPrOTsQELyk/JP6tI64tMniUw1toPlBaY4
/pUZ6FuNFsH/klvgH5PhRyH6t1kFFAXCm+lTsd0o1jYB3ewj39fss7+WHPGRWd2b
9kb1CwJmpO9G05LCPYbpWzTLyNnM9jaql6Y+786gHUp9r/9Nn9WllC1gordXimjU
J5osVkG7l8UG+pnAq3OSiIWsYsC4kryNyWkEo1mcOgs+oeLYwbLFqljtmPN+GthP
Luzoy8GqPOghZUpCLZA3+yfTTDpvRD+QUzViuOxjNYt9aTi2vdovCgwYX35oIOvO
2hsUKlmUl//CYUToPiv1xNPNLe2KFZ1VZV6bommzxtnMjcdCsqigJ9TqcczPtDVR
mNIv6qqtysKggGiw3FnLTjR4IjjmIviCz92yR/eu93G9EHTA0z7p7UGVx8JJeoz3
Raxh4Sr3FV9oJTBHqDQMByyfPATSZo9mokKUaXpr2qxodp6JMOSlKn8GkCn2rinr
hO6hqCPon30Dfy9LAtZbSioDeEDLmSeHX4MAIo8IA61bKu1Q9oFr9azX4tDtNkKE
kLeth9hFns68Z0x9alKagTqTU618v2++zewTtb+qkaS6kcARJL5j0KdpaLOcMvUH
2Ey+2K/fQIAreOIN76Aqs0CsMzcvqIpbP051Uq+RpgzONhH3PcSSWFw5/6y+H83b
HRWJxym3tqCdg4TzNlYOaFEECOgFV2mLMWHEAj6V451tydmHebad23UT9E+BljAw
nKBcdcEW9pDsy1st1nT7IZrEXExdl/Un3p8JVkeXZ9e5GY4p9+7f2L3Uk9IOk08L
fYK1zsQgAKckKUC7qB090ecuC9k6Wevgswv68iM1dBGqkMBuLUP+yu0PYRsW0aZl
2GAeLY59zCbtOykt678rRfnNeyAfu+fgeYU+rMX1GM/edAC1rxg0TAW3y7iiMV9w
YGHAex9xDylg7LneRVQ5Ao5lD96aZLNPuwNnMjTQL0ctONsq1m2N3sVn3A7rG4Ln
CsoqDs2E7WmFacFwMw0sjk+Iub6fAaRTGO54WEtnWP4azyHTSCEe5MnGRkGhljPx
2MZDbKSkpmdEf1rkOnhXA+C32DPgZrkVYoT1QWUB7uyaN6Yxow7wgb3DQ3YWdStQ
7INXtOfhnJby6CQlK+XFVfd0AnJbVlEvmVcrgu86sWYL2T6fSGzxZNChRIztClMM
QJuvh9QYZMXSPim6vQFuTfk8hwPcaNWd6zyo9cEpjQ0qOV6oJJh5oLwTiXPnXfRm
7c5Z2ieijQfmv7bGKq6aWx5dNFYMiVkF4kY8rdkfwQcy+GIj23k3cXI6pr8AAaU0
QKBsB/YfqJk6eWwANYoSXoEgvXUcCZCZ8JXhbfFnXBel6Bjl9C+F18kZkKHgLfcH
W69lq+wvzIHCDbmyR/6Bmfmc+xrZvJVtOQcHG0Fgz5Q3ypbBA1aZrdwIb7TZ/yAG
X8cWQlESAc8FrwIzcyG3H6l3a1JMNoH+FWF8RqvtyoDqwCsWLq/YLzTkyiA8GjNK
zp1K1/41JBTL2i2zuVbNXEKUr8wO04KESt/JNRKhhTGxR2QPBJl078CHmlKS6VqS
J4Y5yIzX/+DjYiUInelmRBNlZCM69BuFE5ZULltLUOxgkya6gJs3fp0r9kutpmP/
+mxWwnxz3LWnrE1c272Ps87cg42Y0P6lSVPzMCHb4GqfzZMLJjnp8o3JODApy5LI
pTCbt5WnUjZ/AGZkzaWQ3zDjG9i1X9ujC0OA66wfx+RbXVL8EteAZJDABmnjUwdj
`protect END_PROTECTED
