`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CtFCJTNn7+ygcEGmG6H5TwMOiunAb5qB06QeA8g3BD6bDcVp9Noun6MPGtyX9GY+
EPKcVXm0MiqaISKkXKlAdvgZoc5muI9+vLuHwnSZlaDwCec5ywD+G57Sbg0zTZOg
VUjo1LcQmA7U93kqDxcwSFXbqTULzBx0P3n3T+0guY9GdFMFI5nYwbm6Mh62K+6C
gpzCtWY/TW5kQMMwsidwABSeDxQNHUmbmKmxVbFIpIzmgpZBVkK/AudKeMUrpQ/n
/2+TpLxoIigm2ow9By2doAvHag0bTnluJIJ0rfQC11w2+7wq7J68AZmZpNk5pSYW
0nvRD66cGYgBFHmX0hPh5QZ46nIG0SktzxKT1JI88wGkhLC+Qt7jo2x8Xr9vM2jS
RsXnb3pgU0ZbUeCDegZQRsUUFgEQuII/+hjl3m9Q45Q6gzjIGHI5jzWl+Ktryrtk
laPGhMW61oWQLL5YR5BCQ/FkUXtWw7US5gXxWnWrl6saY8EguKkvF3NShEHVN9Xg
WFbN1iVvuiXAqQzUJWvptBq565KCB24PtO9Bkr8BpPBewQftXEGt+6UPSsHxvm4v
rBwf8FdVBafDB0d5avEAP/et8YV3XTI2w9sI8Sk8789bWEJBEHpStiWNpy3hrCvm
qIpGnfu547tzI2BAvlRIHVlS2svF4JTnNEBzYz2RKLEw43JSun7xoe/1sueBsDAe
vssc9jVhN4q11hY/mFo3mHkPC6AWI8B4ZcisjZjM9edzdZorDnVNTNuKx2A0Di8y
6HpAD7eQPsUeYON1cZ/Jc7VtrA5pQh6UOqJGQ6fWCvHqy2loJ8FHIYNIRCcmO9AM
vY+cKN5cZopb9sSNaM3luurQjjBq8K31oqgVmYk1ZSt/Oa83lDGrv3LZqwRNcEBN
r4Lco5p/m0kix3lV4uuJ15+qmRS/4R09jVK8c5lm3dNusB4ISj3+Z/YjgTdM9+fy
B7IVAo/Aq2sYchrUUSlseTnMa48sfPzC1gMZSwuvhxYpf7AI+2dNh1sSCPC1mCG1
ypIlHuwpWSjj8lzrLibwOwPRnNEuckQLeM3+RpQ8dmU5OORMuUVxv9urZNneq35n
lKJehMt6mpOYo2TaxM6KRLB+LZOwAky7ZoVWRsx+3Zz9GAtVb9HmnBtQM8Ks+kqx
5wbGl4LrgQHVcXTMpxo/8vkmIyugAG1uM434+uXVXJHYyLoX+OOGlj5tlmButN38
KHGJ8k417CWXNRlXH+IutJbeihwAxvbL1xkLd1zujQdhffTmri5iR8RG3B0Yd/we
tJf2WA7avTOfVNMjF8U1l+hjp7jPNU3ZWAFvylCX9SYN1aU7XVQRDlmJ1S4wOnGV
P+l/8h9TKAlF5JByRwKLFGjp+q8McCLGEtLmBmIwV+q+d0sms9/WLHQpVmMi+yNb
RriBuUK1NlMr4bdwiX8zY7LNVhCdlJxLAzi6fU1mthFjM/vhxOI2YqQGPwR1yFdX
fHfUc0w2ojNs12ImGhr9DayolGKvGQ13ckC9Z4JWb2egswyFz1ueFyUR2ZrHD23Q
ZosTu5rdCAofa12ZmujtxcUUvZj97zr/cT3GDPwBNDKQI++uEh1wtrNYrXnJEKzv
18P+wMb8FPWZZ+jdkU8UO79Oqs6vBMAiLnQQFTQ1F+YVhU9GyCkKWW6V5KX9Kn7+
jZ6d+bx4P99XrsTaIwcac4/DwFiNsTLqEVUKqvw3/wgp4GSW431nndBkkNN+XK7R
t3iktyiUaAvzsI1xend+ElTosdPUpoQbxLNdrh0CW1TUErBHuatkFksy5a8FQOHO
FoGvuNHK3S18MDgcAndKDIZ0ExQgXFUbYetEB3wKNkqo/tLZ6yVdbWTy/ugqz/GB
MXAAHAxD+0d7kCbFRgH4sonkOI2dDFv7vbW5W4HmQvIXto3oXtTwZXEGBpMoxfTl
2CCCM7L8vWiX9zNoTt79JoENndyJvyH0kB8aKm9nSZbXNjA64KhGX/JStdN1TKF7
TdBFtTj+NmMdGOXc57SsC8WRZnUFxPSY9KHkWLyQlWp1S3zXIU7depH0Cz3+M6Ss
VNVrHbH5U3Q0dJlemr/KM9aI8gyuIFErNh1wdBdxn7EZ7ArQ+kiifyXRRb+d+ZSg
qFxrjHobQq8Li9vJWAAHuYYXEvc6BspPaSxmqBz4IA2mmsC465J3DlYuH4WofdOl
XbahsRcFOSDUm4noWmvecHdQXqRr61DfAZHxCZnTkBbFAKSBv3HUxMjc0IFWqDlB
A4d1tjemnWBQZpgewBx/2I2JVtWmspUZAi/kpsVq6OQD3inrq9ACm7XRyj3D9tRf
8pYCo1E7xq+6fSGhRAEjdtMki9J5KXaIW4R2WnLFTJ9u1oOEQjpv0ztSBlMOTa4B
Ot7GUpIzY7K4iLvpM5uzmpl/Wl2UBazLftaEQ9KItpPt6tYFyBNomiC0uBAHyKnu
oF6oxJRe/PmHAbEJ1MSB9hbcZKm/sElcotFAMv+Qq/d0eNQTM3tQ/CyU6L26B7PM
mkM1Ae3VvflxHru6uIRVaSD42rRyCJzAOzZxFne8N95ueiUKoyFBV3tXFfq4xfMC
KtJD9xG+sIIE+a0yS+t81fRS68+VxJftwmaSOuw1JBi/I0qk4zrr9xlB37kiqbrl
5Hgt9iloiO+aLRt7VhiKw4UKJmeRvF1r6cY8iv0vhwHNslxqxTqdlbgdjnkNSgDW
UZ4Z3HkaNojvr7km9QfXr/JjUIPdEKTaZD93I1KH3X7d8lHNEgXheBsX9sPe3Lgm
TJs0qaV3J31VWrPOyDbzFNbIFa2hX6wsi5ZDQzoCMgA2IaXTTDUe9gtgXfd2v2um
n4czOah+LUQ8wgoDY/rz4n3EDvrcHp5nWnV+iWdVNAxIvtKOsnqDZim1nvxlpBDj
e6rZZC5rY/r81kMXH9r3OdwFLdLPM0O1WX64lZ2yf5yofmz6X4XqiuJ25vZklMIE
sUnZoBrKaZlDQAJrFTvc0IcHe5Qj0BmyYizhKNpThksxJEK/Y/KG34XUCJ/saa77
QsayqS/s8ZnPg1r0PhduSA7vNYckGfsmxU84MA/ebVZQLrw+aml65+ciTrOB2450
h6sKH+ZGWeXg5sbzjzwGCDUWJe0aa/BjHHo63I+TN36oAymZPAWW2/yKYV98VIWM
c8qPRqP6nRwMB5Zq9w8JRqYlQfAiXghJdNzKKMiKF0HQjVR1Ptis5qU0k3AWbbC+
9pov4JjzC4ez8lU9/WF0vf6P+wvBSlZRaoavbckMLcOa/g0RRYDer02NRWk/+hZn
mv4SJbRl5hMY/CHeARokO6smSV8kX5X/XvBMcuxp8Xx572nkjXobz9VyV4tU4hUu
KgUS8DwnDs4TSyw63S3udFMykQDo1nc2MR+FVS7LxrcJhJuP4G4QclbbBjrSyAGP
N6BL1e/WcGiRFrBxOl6Bl4U3a2E3GCWX8Ouf8T9TMK951whnEz/KMsTVJljLYh5u
P5ISZdrQdat/bAwlY1Q8TyDNQmS5QMFkIX8nh7XwkVbo4aQ68aoQ2Sw/E86NQ3gV
RbJ5GwqR9XysZSCmtTOViBi/pITviGjW7d3qaL0jfjvU7L+/SPYnWVtWmTK7TPJ+
nfyXTPaA/dmVlvIpyVBqc8+692UnuW5Q+5dwuJq8TEHXfBv9PJEwPh6HtVQbTcOq
iY36zUhu8lwksO37Ha4xgF9vWI+NzSZfPSSStGwOFiyfwRA6LdcbRMhjUIxX8LW/
tyfvc0wXgmMWhfFoZM99iecpF/tjE4MBo6BYw+O+r0aM+CKnuBM8UieGtNKUcHvI
3q7d23mchdXWd4OgyDeq9u9wi5DOv4U+aFz06ELzl1DCHxntpGs+kO92z11+miQC
i/eM2TXlisCHGjMPiz0kCBzUJYy2r3oAma50eY4Cd4MGD9OM/qaxABPkOP4xezeU
0K+XVlLcavVuyP4Ivp2Tml6tPcUBKiSwjHG0C2vD01nSN1VguIGdtUcYnGDcvLSB
/npzYUkgG0COsPIa+NV3EoG+ArR+mGQECKfQK3QhiyGiga3W1DJlHgB8bC0uWj6/
9ueNTdAJQR/v8uHngmQoPokn2Zvs2+SmfL70w1qCjD4ltWAJyTdCVm6GXudt7i2Y
T4W+TlHk7Vi7sicVNA5mWOQbOlTAI4GlFSDVpd5TTcbax80W/qsKmx9wjGyOjgC+
StHsw4DqH7R3OLBLgcnJbJZzTv9NUoZ5QcLiF9LpcxIhwGIdpIP3VP3PM4E8Y6J4
GPk9O00TXe7ksBax7Ug7l7I9q/VvJlpLSXvqvFSAxYn2/sETGgCulDN5CMEy2K0V
xZtJCQW+Qwgc9TrlDlddUK9emJ17+QO+kx/Y+CGwrIHmqq6nrCSRieLRq7mXG3Fb
IiAI7LdwcaQwbk7WYDwa4M8e6qw+/r2a+74RGv1thcsnfxaEMmnp9/6cc9joVkq8
6JdFTk39JmtUcsLAJIL3Oqfvhch8HMwJWlDL9NOYFcf0XyDHXOAfpEelAk+W6/9/
hdk2G3rewjD9jYjYQHghyZVdmQnzOeidBPp9kMhPE3pz1ISQwGrqqHBs7miR8Z2b
0NnSvY7PmHHgUOVfon69Bp2lstxx6nkfN/0cGfXY12MycEV8Zw3D/tPLBjuujS4B
4VMKt+dfC+yrIOF8cE+iBiGnH0KsenSQclj5oh+finXnTgt4fFJmZ743RRCXuvs9
jG74BE6jIJgKZYlvKNcJEf11udGF9NhsA/UAn7tSdIX6W+SyhIPxsjyDdxI6JNY1
TKjFlo/g4B4VM1SwPBcBr7USo52fvRKl8TYZ/3fSzyezcy1NbIcX33R3752nCQMK
XIMtkBFNezWNCexkiRo6lkIoNoXPBjkMViyK1TebkLbXoLmMoKxUNf3YNFgz/V00
6vYeixV5nt+tx5Uk6vlsTuro7xZmgxe5wtzCnxMqACm15d1fWV9Z47r6laBn9sj9
cNcm4dduXupXMPzOFoKrB+GbghXUHz7fz9MOr0Ox5CJaqKO+iG1wCIB70EwmM3MQ
4Hq+Hbrnx/N9uHx2bJ13n9K5h2y3sk0gGAMvVm/24E7KcDM7Vl+unyXKTMErGPNT
5rF0tKGWAyU5llG3PkXb6h0TOduoWXDkHCPLC+1lLWDl0MS2yxPW7G8pyx6KZHkz
d42jHOX/jzq33dA8ATfvaic/InFlqEK6nEM2lHkaKuGVrl22lniq0AZtmL23w0DF
9Llp1n33dW/zS1CIAkAK6q6QitvlMNJlAsg8Z53lBBgmJ26qlpbBdLFxlMhttjn7
iCD4OKN3bnjMhMPZ6y78zwL7AM130NEbY194+/Wv3Yi3LXL7Daqnj1RdnTlPtdzF
5XOKnGFTelPY0Bzyt9eime31ZCf8PuoySH4Ax5BtMVGQ6+/uPFnLLseHvS3PCJQv
FrunN95w6WAF8q00uo+4Ptki2YUEybkdutQq1K/0m8MWeiceQVbfODrvVkumwFZQ
aLEkR8OsC10PZ7ua3MS2zJAT4jThJyROtaR+POdbexBCDiva9JIJ4kX3rJGI5E0U
L05PFz3xYgXmgRN7gEHicg5DutR2WPTd18u8+YV17tmF5XkVjbyLy01bU+orwRJo
CI4fq6bzY51zqc9zuaQ7nRKlJMXgSRwaAGQf8e6TSqcuFGV6COgjbJcWYneXIv+O
pnewUJ8iKcrzFwwev3cX+XyiyBDZNvVwdExSRDHRSjePkcD25XVr+z7FmciDZrL4
xl3NdPk9JLlbAhASc1LDoh37s3S7RiLzz5CVQpI+ngcTIFrQNkQwb0ACpVa7uLpB
pNOxQb3ELJiHP7V0uZemdOnO/jaVrEqnvC6q9CVEbgoHiz6kGMWXhWbjj8CeAGC5
yfhB3yBLCIVUzSPa2Kn+HvbvAn8gUJzsjCkfkaI65weK8HWl1Ue6CmifC+WJ48N+
0409TCRtEvpYd6WvHBCqpL/NARHJoj46kV/9lfQza7a1Lch4Kw5XCCoyAeG9k3cg
wnp3dfGCXkf3C8E42PIbXeTTF0RpynXnyf8vkdQSBlNDPawuSNZ6V7aUNVHCkIsg
WR6tUPKvD1AYBGc7bDAUEkgtUrkl3xPArQHphtWnxnswVPMu6lOnQfck/cKfWVbE
WDxTFeQZy3HtJhOP/1himOWzLpu0LXAz2HezgpmkyRMGRfDSYOnV8BF4y/RrZvl9
j/pyE6JAor7HJG1tVnwMOpOTAm8amPegDrfEfrSN0OuqSVPzin/7ra9wjIex5LMb
lzEZNoCbYpHRGGqg78lDhcF/FTjPkmdsEnpFOJGv5uP8wZeUkHwEMgGyXZ1EDYLp
YD0Ieyh1Ukgic35UaPAhGofFDnNWWsg33QbJbxOMWbMtAoTc+hydNu2I5+lrRQzD
iL3rM4NWTg7/fnb777H4/MsaBQhrF+dTdj6Xnvp63AuucyImFdVzMxIQqdNmo19e
I2zU7ZsNrLWu1yQ3D3baVYEFFbGQ36h4xKE3UtpyYHe0c2ofdvwhTxbe5WHZjUZ9
pNq1ygkuKUJx8BKKEqRVmVHn72t45NYs+pzumA4c6/4u9KicJmNvpW/fhbEpO7sH
VbgYDf0dwDcjW6cnXfJRL0nMt6tNcc0b7T1fO+/D+e0fkPiTGweRsn7/I11aK+N4
6quBenGvxUdk78nHHUTLO06JPEj65M+0E7mpDZvnRkoqqjm7t0Wj8fVYM6fCLNf0
bp32vwqRxbFSdPbbcHzO92m0xxl4LXoSr7oWSWMxapsz2gIrvPyGITbN10Z5zp+w
IIsAQ6dldDDqUrDTRcX0Gyo4wSUXOSmaq5yLKfkT6ME1QeEXBjvVHm8P0wEHxUnN
3BU9WuEABkCdq5FbGy3BTrcoqy3JVEhgDYK3YVJIcqQ0/jEZuqo+3/mRjkqCf0VP
VLXzzf4WHAPFbRz9xaD5wZfWUJZxkz15yIJndQKvslZmRPbC6cJ0b5GDGzaP4xnb
i234npZJnvI+IzXZMw57pCa5Sm7IRc7mOesI1A2rziteK4ayiwcXoiin3SLBQGGK
z7WbLQ2ZrjM86ne0eoqWzvpstV8zXUUYCuPD+HNNjinFoZtshNmKShq8ykZvxsg7
C/eDiZMhnC65NPVB8ZDNzRxRsiQq/DHhMNTaQaM7Und70Cu7fG5rttKImclK7b0x
ZpwSiuKgQV/kUMGrPz6eCcBDH5/4L069M9GXzApNSnu0HzPpPgC7khFWGS3ffsdD
DxvsTdt/4NRycZDPUHRigglrb22CeaKqD6tXxZR8pzfvwLhaCnkg/+fWYCOUQkN7
IOdYDHEsQdWWgGLufB1xaLyVheijG/VD7p0yfE8XO3wmCGu7bPIJ78G1CCWKys+k
ejWKMfzqLJuk52VIDOETqw==
`protect END_PROTECTED
