`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5INEQiFa4rc7vNOCMFIcRkRZQ67BKg3oDMJP0g4csvTOt0Tgtm6cKbpRyu4MW6d
LWPWxag4Q+Q/AOfxiULaYYzgaAmUfwYIDOeNSCq+F6asXwSYCCSAyo8WO1rW1Y+j
tH4I9R/gou8vHpn5ba/kpTA/pFomJ4/I89yQ3Sk+AvZHJmvARh3lOjPKCFL0u55S
ZWaXUKEZel3sfTYhTyKdzYwWZcEiWB0mgFrGtiETRftz8EDa6NhX1Z6rXokRvji0
8H3yxsmlg4yW/E96YfKsUI52lAE0ZDhC8jW1KV+v7lxEpkBne2K17cMvnJo6yJYH
4yG6uYj+NDJXQjbTva4F1fgWfOw41D18wfYRfU8+KE9zL0L64bVsDJjy9+Anu1cn
D5ImH3enrH4ar+MWoFs5SqFs0bAj/7tU0Z1f3st4k7aWkUsuLHxrsTg8JRmw67Yh
tMfo6Dlx+9yKmrJDswOBxBHlm4Og+PqJ++9bWXT8fPWaB8DrWjecdq5sxyiqjCBV
mh/YPzFs7BVpVo0SrAbn1/6nay+uH7oKJVqITPpUq+CpPp07IrCYfMOORjdBs+L1
mXsAiO88AR/iKexKwc85VBE84PeQc0wOnQc/lsrKjiLuRhOIKHWKUgjz2/KGz62o
4KQwRgJJ1H24WqnL3A5XnzgNq5lpkvgphy1+y7Zrp+n6XRJS1Krt3LO9KZHHlcON
`protect END_PROTECTED
