`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dncLfCSdkb7z3prtS3jlZWVAhqBUnU7NeyFtHZ6ErxvkBX9/ZYdCdmBC4R4/vKVB
g2Hwot99tOonYKvijNHJ0fzZCKSmDr2Eu8ErMp6doyI9lor1435Mu6mOxsDrIgmS
43x2pKjPokhx6HaFl8UkMH5xtszKdmjhmhgdisBa5pN+ot1CB2zviqW3oM7DX/ka
M+vKgxJWRtaBkNTVW709vaU051KXRXTsA55C6haA8ztwbtLU7173pyoCEj1+9Fj9
HKEd9qEgdeC1IfOQ0dDFJBKZJj/aHsHLbpoJelU8A1pmovoYv9R03C3ZzbhR50vp
MXz3abUrCoJ02L2z1VM5Fte9ZRklceTIXymNTnyatIAPUaV/LPNQfPq5H9UQSRLM
bOqQDNPXr0vM81RaV3C8H7waHGXy2WedBdgvkEbSkSUB7vA+ayqmqMOZEwujEpeZ
3xwZ7R8xVUCCSa3f5CUZgShwmPy4b96to4w1j4lz/s2ryCOFWAXXFzxuIPqcP2CY
OqqGSM4rTS/0zadGbJ8ZjLYxbJUHFdekuk4o6rbmk7EZORYQuz+TDSXC+367R3qz
34CPmtnroLEDzUcXi7ihlcT9/6+g+qK2G/jFTfqvt+G45EcSeVjA0od/NTRGrCfp
aL8HoMIo7dtP9fvaJcgpxN4KOsdq5eWe2Q1W+tX+I2aojXKfs5C55K8TnYXV2YtC
HsA4eMouHgxtHLmkDy6xXszlZTftPZVuBs+yThF6hTmduQqsEg1rt+Lr3amOIgrS
jezXtEu7ouSeQ9g/UicLUebmJgSwGZfhRLOC6yCoax/Ta6vtKKEvUGT8KjZOYHpY
riVnAPw+baPxBeReMbmiZDZWfoVuFIAnfdqNtOjYVSs=
`protect END_PROTECTED
