`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOcXbJwiewMwZVvR/9yUg/oA0mrHBlkdmMNoVKzYlvm7AmaRc+ZljrtTZ/WQy6pP
/9g4OGsXCeBKyR0k8RBF5yQMwFiyPIUXssPs3s4Yp2IIVAaX1nvtwQVtzDyi3pGX
ieIRBduf9NjXA/dt2B/o1UXiA+P9Jmjv18380FFoFYYWfVUFP8g8Im6qkhX6bRjN
UM6dbJz8oDov6//Kfa7ZoeNgMI/vfmj6SxipWsSO7NFky83ZYmXNsta4u81tclMz
omgSYTQln2qepBySGljvMqnWcxX2qv5LLCo1YuJ/I10By/GSDz59PJlHClAg1k0p
rVec5Bi+Kee4qLq+ijCkrxf+xjIWaG8XL+FOKl5gI48DaJzWt1CSAWR49u9xi/uG
`protect END_PROTECTED
