`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tY51JLayRFU07uy6VTFeMTF/rAtGD6C1RNhMalwRtc0gAXEsjJLAN9p5EjkNLYjB
Hzq68fO6F+Drewh6BtlpwjCrFsyxqudjBwG30kHgrEnnxS3PmYJcBbcZ2KkyK92l
u3y3ykPyFa2s0cNY9w0ZC705PX7/QAccerEQ/t19wDaZDkqK6C8ntQgza3Makac0
22Hz5mtHm9/ZhtlutJq4czMcYZICh2bhs0OIEiwsWiclKrFGYPHC+cT3DAxtVJ7L
s3TSKLJx6lzIjWDzEAQs9D85tEyVT5DOkRLW9zmngKnybsq9Ouh5uFRohGzh07y4
Cms9RZq+FmTu3nNcf+wrhv9gKNYwZELE3kwVhsmvTPNeyOTzbF48D719uQ1K/88d
zq1pJcFITJXOtA5khtkS33+Zau+JZSlvVeOMzUuOsHDa48UFoDQ4p/YJIrO7lYx/
HMXUWKHgVFIkJvEYJCttPeg8LZ/VTfP50IfRcFqyN+RloiaMuYeOX+wLNB6ZqcRk
P2gdZQmUQBbcRZZRmLiaInfViddO0ks47DiKe8MM80ZSxAKrffhu9Els7FVO4Nhe
KcVV3+r2gjCvpVu+LoiBpWlJJnMcMQoV3xKK5oZJacq29+eM6u0ddLWeMm5kFvSC
Nat/gF0jAeYgthsWHKIBosUo9dZ0rQRUQqpxX6pc/oIk2GlKORvJil4a3ZDjk4ek
A50PLWZSsIvDUrMW0t1U0cZUQ6wUdFWsQLUd1X22jKrOZusgft++RhG2mxQtGEzF
WqUiwrk6JFb1Ize7UwRrVkCfR12iiQJLZy5TChUeqqmBJbfSma7peP/0bKPLxxqR
eGAfuTOXiU/CGlzjPlW7P0AQMhSxAoYAi7aVuhH8tHUz49hjwupy2UDZO0R0sHcn
f4G8yzVlKQux3bqXp5/W74esrotqk+aNzDQTSoLGXrp7kRd++QT1M9+Vz0z/QsRc
plzpoVe8EUkYkLmi8AOD5LDNyEfs7d0+3cEGy0RAfZwNWL95WomfuOMMUxwEi07N
MKRaCSz9Crj4adL5xPxCu0pkt60if97Qz0s1sOM/8O/d2SlFCS+zlPM57kAMJ99J
ZRmJAOb8nY9uQUkb6ve9mCKLGWy6tGHKTbrdH7fIIFMQ++4opQx29ZvSWnrm+FxZ
yHb8UEQV9Rv/7hIbqFH3h+zrbCWQrvNZ/2a1NL+dcoq7TINf4ePaZ9vqPPFGP63P
XRE6VW+6sbbYhDYaKZHbc4L2RP9mzcGBHmWzm26y6m/B32l6IcziEjsNsKKgVmsK
lfhxAYaxuAtPZOmYNp5E6cl2z/lm3RM577sa0ilGo1daK+E3rATvm4g8pvCuX+Z1
O4Fr3WgNST8esTqXYFyDPw==
`protect END_PROTECTED
