`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XXXR/xKEkRDji1TG9d389F+N7TLY/XqeLwwwCx9ppYHG2kJaZ9AvqfV7mYQk8sP
HynkJaZsQ8PSu4v9vIUfGX8db/Hrmhgy+0wscXNs6y1M0Z1vL1Sc9elhbaC5YYU2
2kgzMUv6vya/BmVWz4NqiS2PYDYVVYMD70sP/q2ssSrJGfnr0SVTlrFaNIR2MwcI
hoedyi8Ax9jtLFZ4kw2t5adI16SbB2MVpylhNjEbAYKXzXlTz42TN5XyoCzkqoir
mggEIoUeDGRaJ/kI69GUYa8kJ9d2MBfAG9ZLkwbE1DhfBBq4YXuYJpW//hNM/ov5
LrgcLs1ZawA6jkXbUpdJSFQJOqUY/ufvlV3ZAOTaqGx8LwsY1/pI7GN6Zt1TzybL
AlSV4gHSTPOW+iZf+B5l5WQ08buZjjpArfTx8MtemKlILmzNsDAkazUnV2/UHzNC
69RJOCG2s7GJmG0dL5loE1iVp/xAkBMQHf6cZ/UtuqR9/Wdv+W7h9wCYH0O3OkgX
xR8pzDlQS2BgTdsV4SlYM+E+9xFDXRECQ1/fXHDw/8IZIxSdiS+E5UpKTNUJ/WO3
8qvMS7y/2si1WH2wOIgbp7EiNuCJ3rhWl4o1XOhjZp6N43H+zcwC0YLTAD+b833N
K1VMDtTU6kWc9vveRpX655+/VQaUwo7m94oYbqApwtbk7XiItzFgCmGEYHF4HcP/
IQWo2HW4WmziV7JxuXEw5od7II6jy5cPumNE5HMOuD8=
`protect END_PROTECTED
