`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J1d3Vi2C1bJfsVyQyJRatYPEjyCjqPUfoZU7EG2OOIA3JhSxD+TuWWFGJVis6GUB
BcSxMdi1TvpkXTxPNf87foCo+MCGDpI20XUKcNqg28lnw5kILYMVthpdyDEenGOd
YhdAocmZhxWCaemd9XKa3gBDstVXL6VwKAlmpQV84qQ7Q/owjWpj2E3Fe3dcOBhQ
S9+kFy3XaTNwi21yqPww21e25fExhjYdkMe2RMO2bwhJtp1KMPuPL3+FLX3XtTLg
lpNSLCq0VINkS1W9VKsw5Je2vdeju0uPtJudNf33PlLoy+3h3urr/kSkzoPLj+Mp
tr6Z506aJNIOaffiaYdTELryDsiW/3FSFJt8z3sJgEvgCcZAXGGiU+wktu86CEok
Qz+a0Og4tsjDuDzvKnn/9WixEdnm1ShZoeVzviuTujBJ/5nnm2J6R9XDBRwelied
0r/QtnmYwIy4/jt+0yfe7ChoW+zweG9HPWWKJ7ls/9m6c/tzAcDwkJyJ9rfbQ5UM
0bntfYkx9CrWItbnY35OXdHEBMtWoWgLZXXVne97bzBUT67nf/F2c5qDQTNe7CZF
Je5+bi2mMFfVBLhA7nDVlV5iXw9BjL7xnaeWXLNZl8ZEy7Fmx4RSWaodZG2SFf37
3F6/A/PJhgMeo16mJFIkeBikvXYSiFB78Q/7C9kavqNIJTy5cQE4oz1L75Uu6OCs
V3OnCW+irzH+7ErJthMCOBCOaQQF70mJ+KzZ0pXT1G+dhDv3YknPdTxTWgv2T7Yt
9qzdZbOb6EPpJrun/iJDiZGjlW277I8CP1uiVECFAr+nz5Y5zG+WTh0iWWw9GsS6
ockMyKFKwv0qroKpBkxyXYuF/64nfZNWJqphV89NLVFUCWz8ofx0TzSJoWCVYyyT
WlVd+kJT/Z+7Xsp6ByGP+xycfOuxsCVocp93dw5hBvARLOcu9sgX34kYXBbscEKq
fSL+W92lIyCaZFhlLwNkl2tPRZ9Sfwopul1v3NQBZvpRnp82TQQ+9ilc8T7vdSbH
aBiWTy8/wzmxkypz4aeww4kuICXbN/tqlY2QDJWQssjSP2bz5PlRRotgMxu6JDuJ
ouT7uV4WA5O2T/5pAxM1jxWeReu9ETp4PwwQVpSKPMs7XC3td7DtjXBVUSSiHPbz
`protect END_PROTECTED
