`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sX8VDxdgW4hOuAquICBBzxZ73ZheG2ZxpKtSUBg4Jaq0fArJZWjssfbs4P5mBTG
/a1nsT/GWl6CunGjYUv4r/LaaiEmFAvyhrrYKmwkpmK7GpDcc7SNU/k1EzZNsM+u
prd3N/DcBWpxFo3ExxGTJCoplEuTZmIZskCJ32VCN35Qc5corJ0g2xNOxd1NR4OW
Dr42SZZyc412wh0hGN00JztyRvgZyY569su8eLfYgPU6fmJpTWoGH2K1+RjLgvWn
rfUG9HSH7pT1l+/cAS+yeRTMJrMSvlFSyHV7aSZ0xLWKpXHg6c9M6NMB6mTaDehX
7ScPk4eHnmj2V1Imdz52INBxjP6Va/72LuRI/LxA2uqt3ZtDKNI4NlezDBO1xxzt
hzO8b6Y+ellriYY2aW300H0GViKSRP/hPGlp15W3vlEMR9U3sv5ZXW+u4lWY/ZfY
sl6tPhEuXT0q9pwCY67wGH5cukL4mWRmd6KlihZLuIA5MsostIc0N7M7bmVEkxfZ
/9T1t//eG1UvJz4VUqiSSJkhsIzCmiWdd9gML+2Vo0jfRrYzavm9dfdRVlEBjOnb
wgZ29LRcF/IjMeNu67o/ltZkU8eJQ+rUgXg9X264ScoF8YUHW8S/vACxcMrUQRd3
bE27wu5BNXspUyiW4IsjCXeDxXK7VmK9/v50RhN0E+JndFZ//ODsggu/YHBo9fes
IiQZ+TI78fzO4VgWeh+PX50Sq1jBgt07gv7EdaiBs5PtqDla8T3ED4vyQZZsd5o4
89MBR7jxvzZIOmTfYsKujIhIUOE/SzlKc2mB/3VCjuDxAxu5ab7lPyha//xXMwxX
I9OqfpzCdx+8gO6s7LDpC1JR1PhXEUW1TWZexcav5Ecjva5GZ6DyY2AvcuZEGSfn
2kcyTuMD3hLZYjWgr7GO27izSOY/zbl18jOQkPwRX43pVJ3u8yBFxgBP+XyOaDQt
nFS81GLbeck1RiZ3sqi9iOlkDBBvcc489GEgc7Z41rA=
`protect END_PROTECTED
