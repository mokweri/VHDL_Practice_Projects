`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5jSI+RIKdNhbduDBCALHwbf2VRm8WT6jelYMsKwZlUzqDFkYWSMEh1F6tqG2Hh3t
b/Bmay92N8v8pI+C1XqRlMmpHdmoe2EO+NdORR5g5JoV4yEu1Kp5QLqToKm042Y+
uZcRCl5KtHLmyobQYAephOjGRqieQLZFN6AUrgde839Qt2rYI772aPPtJ3qKkotN
tYSS35kO6rwkKQCf7gRxPluNqberpGQMXJG1fgpuyO2IZMNfDlIdSHlZJkd+cdSj
u1EKdk6wSkUVwCWC97YX05n7Jq8CooGck+RuGsKq94FV10kNYGTllCDn0KBzMqTk
r9/Z14X/PM8cV3ndahmdd+VJiUjAum3B5E/fpwo1C7mP5ISpDXaCmaS7X7xbtfgw
N2QTBjY4cC1mYGcFNt6nGPNqHlWNm+1zRgS+EPHuG4HhCYf0EAx/TJKXJpXr03WL
vUUQNP+m6smsfX5CqtHi1Cu/u3O4Lcl2/FPYkQHtt3iL1oTMTMorPEJXctK23Gsz
ORFW2gptdYdv69HpMA4/Ta0epirR2NNYigQQDwlq9D3P4UZuPBODc1nXrTVGr/E0
zXKHJaOnUqSasdZl+gyWM9FJvlC8o10H2/TdycFsYnNtNKRU38EItaeYmuxRpnXh
1fRc8ePyvuwGNO2+T1zQLTbIZ4q6fbryXfo+bo01Mfeu1KFAgo9fm5fwTp77Ex+V
wBGzcHnqlMxuXwcxZyLhZI58ruVm63MwUq7Bi28+pd2OYCdL+lmWH3D16dfgSkmy
I+aMN+PoIsUOrfFLpkl87JlQNy86GXK6ih+BLZ8gQ/JVIEcoNPUasQDPb8Di2tiP
Dp9SqE5LScSPciAagOvowrbVRaKe7916NMcq08zmqqRljDG1hAkzSieLZKfPYkf/
PUyWL7AwNna3GO5dnc2ocABFTBAHFReLLn5jirvoS9tgLqu8HhN4s8qzpo7V6RQR
hFX9N6of1RRz0bD25DlQsrGGp8Wni1neLz42XY+YK1jcb3jk+ILx5BncEYJQBzaq
wd2VrYZmJ2lW3El+OXbw8i9IsSHoAcaTXVJVrTvPqabkJ9gMwhSg0FMh1Gq/VMi0
GWB1RNmwz+JLgrSSIoMSIZiV1zZ2ih5mepualjdnh8EW8tnjpelgtZ1I0MizcM8m
mprWXZ2/u4OOydjGnxH/AyN7jxzEY6mAsmxGM55YYftwVT0Dg+82PACKUwCtWP+y
dssOofK1e8Llx3WVRR/OLvD/iQzwSaVUXXfBcNSDG7p2Aqak5CVhtaDDzrnorGRY
Pq9jhpyN3fE1FEa/ujW33ukJji2hFnt2N3R1tN4HyObBsmIaqcrf5Avg7+34S1Sr
eH/+YQuxqDoEMqs/HC6sY8SyO4RTCJU9BMRNXgWHCdMZJ2ODUKkyV4CMLBWbXSD8
WwTBzJvPbWCUEcHntts1YA==
`protect END_PROTECTED
