`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9oMj1W6f+ht9mOoCt3po0aUc8w455kWyjoow8f7tffg+F3GMLbFWUzgqz9P9daxq
JR4P1pdT74OND4JvfWdP2+K9o2cnOCP94vcCiB21x/5Lb+lyfa2A2xbAyx2g1mCh
k/IbqxQfkL14ssEVw2Q7EjiHIP/dpewNSkiYSbPYI/7YoH9C2wg1sYtfXNtCdxDr
6oFiVNpWhPEeVAXdMH9377b6R8jT2S8X90wY/GAqCDMWtPq+7qT/z4vQNUeWMCLU
5mRqdhGWVVq9vzfleop7glhmUnytoizYqgoi818eg0QPGZeVy4ABRGd/8w6fa6uZ
zy+rGOVjKUL/jEqbwi1j+aVkX31oihuih50n86kQ9NfyeHoTjMvsllnfutD2MxGf
h1Q/CnDOeOpwRS7R2O9h0nx1zqJPPDHKWAsqW2B4+Jqjq43YvPW7QcMXbYTkeZDN
TNxhkLF35CalRXwPnyri+jz9jtArZrrYIE/dQaoR+2FO1UwlcC+5OE22jp4g3LWx
I7WpL93+fMF1uMBQ4VbVmC8C3NFvR7A+V5UF35tM2CCrPaFZnXxCgWwxrllH8gWs
/J1eV+YHFliP/f+hSWAMcMnECsWYuYAqC5Jna38zCaw9Vx/H81Nq0kn8hpo6SBPw
WiC592xsdMKZb9GtHRtDCmsEHx83BWq2v8uFQLj70MmjbZdoTkvEtc7g/o24bcAp
5AzZztPKh6p6ypKL7GfPnwFX+N8P6daiLm3mZSOAcwRLKNC03KE7/SKtj+0gqj0O
pJ0P/thOyiVVp/9En3OZoWbFutXhgVn5NRzlm6Kz6mbQWzhn4A6wzcIyY1ULt0K0
pmaLk8CkKPWA5otiBT5G5/B+YN7HS2gyFNqqSgKrffHAoDbvMkNcAGCOmoh4VApf
tWi0DvFtzWAgmDN8iy9aWr1k3JdHjJYF1hqEtetGNMwksA3tdpN2u+KPekHt7Drg
DVhVxDF6/XnCqyTuIDxDJ7BMRB6FlrbHOgpJ17vyXwrPUgA6Dd3Y0bHA+hNJ3NWP
okizakK455eVEMdyJyIML2HlN5UM8UCE6TYnfoMArlaUg9HSve7fDxceiqaDYavY
wMFVlAyzIdWUk/rhzmFccvB62abFbCeQOF6Md51GJMvl7m13lkecGGMuAn3GX0u4
CV9mnbEdJcg1EEhnOBICoKfB+yvHXtqpekAj5O0UOCBrplEmP17cDUgdmGTUCuji
lekYVZ3ERPk004vWF3NkRB3IxuPMsjXfg8+8ONQezvml9VGRnCnuVufbcvghSDS/
2TlfB80jJiBRXso5TuevFf9kddnxOGtZj34lk3YhLA0uR7KTS9Fq7pT2O1wPWfwJ
vwCcQdTMlGFEPb7VBTq9COyyqs5b1DsY24LGAMYE0fIOyd7gm+YbBLKoJ10TREM7
Acm7kGwIq+MVMHspmpnnh30iUFIvbT+BbHYqy2RrfoZev4hV4/263VhzhKo9YCNh
ZPfhNLYh5ihvIxYPJ1EMM7+TpWaqWV3AEmdcvlMnGJnmhdn3wlw0uJo7eii87GOU
RHzBBteDOen82Je3aWLjdwd+cxpCGpmxe4EtAGxyyhBEP9B5RKqcn8pGuh+Ydobd
Yluqr5eVdRkkBots5pbo10r8lHdY2vd2VSVNeJMchwZ2fsuCkHFfMEs8MESqgAvC
2SKqTnzb36z5DQIv/uJ6cop5qQQYJ8sHSESwxEpoaLi4R1lPqmiXN4mkCtGpWRsn
gpS+AUSAqFzLz0epxd8jsfKYOZyJatgTbKeigay+DMfTSaZVSp/Qk9bZ8EbIQ99/
ItDQX0iALWjmZqlnhNtDHcwk8+tfVDyb4sPGKExmx3qb9X/KbSWYZmD0L3xkXAuG
4BT8YG3wxZZtWkd9gWuvukVCB9o9h0BHs8YQvB16UxfogCQQqpRKaLAg/KQXxtn5
kKbJzsZEccgMPtm0bFA73vGbtQLA6VmUpGXyV45xgeuAGLmSRAuTLpfACrDxS475
0LornSkaVrXyhTEciLNxLfcURN2q8mniTwqxfQjUr2Q+xGOh3N7bW6CSKikHdHBB
jexqwrdaJnbHyn5u6zoXgtZkE3AqSG5AlnvOySwKMcJzZKH2S1lrMOnYLwmOP38e
QoRex59qDr6k9M+nOvvz62o9BEHk6mdB5rO8xOfX7humhD124/E+3Chj0UT2Fqrm
g0pVJnmJXocR8NI9A3BKYBVhSD+0SRpAJ2bEXAOE3BXCOzjcRoL4GZ9CuZO/hx+M
XPjuyKrT4DsHqVBCxDRpOivPPgj34h0pd1LOM7kEfw5QqobyhmfWQX4D/Y2j49bX
3z7QAbcyrIwKOLmULA9EtgQhU5j/b+HRskcyNpYg2f24jF867A2w6g31a0ie+yRS
oXyoaic2m6XjFe9n7lp026+gdP0PjsDlsYAGXQUBFxmwLj5RoJYrkobIeUWxz8uy
Nq/OZMnSsrRbZyvme65JBE0/lDR+3hexAcg6p9NaaEnbzQ4+hr/Vz4nrbAmQJR3K
8KCgNhxrDGb/EnY5TnjXniqHls5C5/CJsjE68YJRVOMxZhBAyQKQLgh/Gh+Mu6yp
58ou8wxtS6kAchXJhKxcfHvgaeMVUrS6x18+rphlPAiEwYMU3s4BVVvcCz3g6OB1
1kqdVTLmT5X1cTToYD6W/g4Oq6kIZ2/qjDH6kVJCgYF2tc/kPVu92PKGQTIe4+mF
ZzyZ7pJSYgzgkuzkA73Eszw+1eJ0U0U+6lCzVtpuXeg0KQKdBrAeA4NOh3rcvc9e
wVh+jHErDe9K2PGNuKedcg8vNkYY8jTFvT+ohrcsJrZBGxQrdfzr4e0vHU7HJ6S6
VEHvm7MMO4qGzbDTiPy3HWQIhrfB6Zaql7KKXTeGRNrnc8lMmHDbKuDB0lZQ0LZw
+30hL97SUniib4C5HcPRMZq2CkHpoVK7YiNUfcMd38aYcJOo5RpIun68xXdLM5ue
RLImOpzGHPgJG73ZoUd1/p92CHCMlAZdiw7WQWxNla0E0UkbeeDF/lERAsIYm2D+
dSlzejBQ+/LEdhZKDpFyOIz053+F+M3rXdgVkFaLa+bEj0+V6Uu+RkzNwZElkpW1
HMg8g9DnLxGJGcJpwrYldOEcOzXdq17mQz+Bo+wKPrHrpG50QgAN+JGI0o/+Pepp
E65uCcjolWTXss/iOvsYf0MK8kDi1LD5bUMKTYptfM+DyhSgTaMroh8erPmKx2/g
WULLMCViA9m2pg/1aTXFOJ9cq1DKLfrAq3IPpEBJVb0XUTZki1UfUNQTgyUTSfgZ
XVMcI2o7/Ml5jeMwZhVnhrQeyxJeVJXNyHv5IFt1TA1icYRCNVEoNUd5JHf65qey
IKlFXvWUpxA5UCugBv+8oVEpZoPpufJihI4R+o9gSFJ3ZJqitvhe4ShspZZjSar1
Fs37mRPeh3KaUr+Y3U5WZEI0LFUb0n5a/vPxgKRROEjFz5xbS7oQ9FWsNuQJOWCX
OWrEOk2hCUL8twDSiIwT+XCm4AUcY01xBrJHTym17pwCmgdIg6CvKsyIUrtVOthC
5/RDF6AbnVF5Nqdp7hf/z8j7aQUHzTGuKKhFHSVS7ChekHbZXHh3lTmuvPI3qWQt
4NA8FpXQrixiqw1VkflnyaLuAE+hDBx4LJ4Hfjb2UMqCdTdlk5iVgffPFRgEGH+/
Jzgd5eknluSHX34aHV0hj3DM+q+VmQp4pwwo9nqu4rZnu2WHKHFPf8ToVHUejYz7
33jjgK/Thmio83rS9zBzNP6CVJhZ37a7Tn69h6IgLP8035hGmR/7tljOq+JmXuP6
qyl5jgoerd3QuIrPYU6c2EGcFicXpAsQk1ARSC07SwrVKinPUbZzqc8Hl4AJfZiK
GDnb2FTVme3Yve2hAvRyezUFnnD6xXkOus1/3VCDKpSnRfWJzPHkE/1/PivjySQ0
DezsRy4cZScXLoSivOwTfaP7ZfL0c0hha/j1iA/wgAqvQudCRiCya1nxgiMDuF4j
RZoAmrly2QJXS1xlZ7O9LgSy0zzDdOhv6acYs4/TFmB2bjWwjYYk9pnEutiMgWBz
FfgmpqJSWFo5OIg6ORpSFwlBI8TYHIq4PeMWh4krDGhL85KjezTmY0nY0/WILTdB
+bQEqyOjGA/voymS0O48FcX3z3VuA4rGcgEoLvaSy/CwiSSvy93+z4gRs6C+QPLT
s7ylNi5EwuVbhzbhvkZqWzRzYiSivf4BPAeoJI5hAp81iDfyJ5HcpEzoGn2gMRTf
BxhGNxdaV7ZQjbjksFjZYtRgPHu86Z2hqWrS9OW2PHm2mSTpl9bQGit373m56U2U
SA/+le8jSD/7wtKumi1iU1XZXi9TqprwtLj+cvzZgt3V3W6phK+mdyt2NXWg9PA+
TBpCv7VePKpu8v/8XOq91CWJrBbWDRGHPPLgHz5pUb3Q9QT71jLHtpf116I+o8hq
w9dR4v35TCRfRjHSo4sdKJkU3PgZXrhYhTjhFQXOyCWu7XTEG5COSStYw8euxrJa
eN32na0Rvv6pWwAYsJVw1NNNMAXAwfSe7PC/xylxVhjVOgS47mu/9RucQhRXSux7
U9uVbRmbdLrySoau82lwxQfxQfNX0SiBPaQ4pmycyiOhoDS2aiwRt4a9fQCy8+7B
DLHCBKKlp7TwIcpUvZQHzS4bV+EWxfivyMEGAD2PtGADzqa+q/pFbQNiIfZ6xOdk
FpBYDg//TMKz3QP7FZmMdyBnZBgte8W3bSD2psbN/ZobA5ESEXfqBmmXPewfPXps
IJExzTW45jKiv/kxQaqvVZPEBvVYw18Rh9QLff4Xu6S4gn7o41Hv5fL7PMGSjbbE
3ld0S348cbZ552FRUcKUOZk8ide2SfKEmx2tm6A8u6F/5VIxgDWgR+uZCyPYPlBA
IhTBafQC96r/8W24D1eHeDzz8HBSdtPyiD3SlnLJsudHjBOeyW1pJDDzwQGAIWej
5kmVJeNzrtVjkB/QBZrk00S3b7eYG1A7621sHRXGlSoOTbYN58JEnHRXHxNAEW1d
x2PPGRx6XIr+FMHBhTo4wlNpaBQe8Z2Juq8jysOVBak+LsLikvK9SIANhY7anZ7X
WoLgXuE5tBxjRIexWpS5GaHqGBHdq4OZJ7m/gi1YM63gue2mgfy+stMg6fJConDF
fGSTfiSRDnULah8rAKw9tgkpuKESsp+g2H/W/7/Cbsr174ojZrh3qiW5T70pufuu
PG7rzMWt5Gyk+TuqSU0Vi4y0lNPlbH5rlBkga9HUNOlI57IQYbGsukaJqHgx8C22
woiHSUmd9kkE83kj1CwPyExt3PQq6lROIeArb4oa2PlH6AAZx95TCClK8NCQQWUs
2MoahizgU7pziHWFNXHzjnF32UzrgI/JmfR0YSLyOTHJ3dV6Tu1jCcFVpdqe3/Ig
ZPrM4QiPCUi1iGlk+N5KsPJdqf1JpT9Y22LRe9xtZ2SWB1fIdmnVXeHokhLV5Z0n
8ed/IhCHCCoKP9FoJq3tw6VojNrnHjBHILylVHHx/eT/ytE5DOwhjv8YMUjAURCG
A54wUv0oEdnTsyVOnIwG+geSMSqfq9L3zrUD366Si/Q=
`protect END_PROTECTED
