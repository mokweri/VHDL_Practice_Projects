`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xoA1mN9zrovsCX6COjnPYQfdSBwCWGmRiw+hk0Xf93iyRUrQnqWlFC/c1ryJHnaR
+a9Dkx2Is/YLpXZQcJJRskpFw2oew3doGQdoeMwIaAGD5jmRw0AEZhAOQ3pxU0vw
3yUqob+Hc0nkUpXZUlDbqIW4c5yyCg/2lI20NB6qyxVeqIU3r+dppKv6t9+4WsN+
F0BoAUTquh1Cwj9p8gtsQPEiR3Zab3zSy836c+H4BDPEYiqerMwKzJEGrrgvy1L7
BDf5PkLE2B4B+n3UfYoVuH3L6W9rWdbtFuL9GBrgkG4aALVYSs+YpoioPJ0f8Gay
Sszanw4pLbhhKgRqf3L50gdyGf/ThF1dcQJkCP3Rj9Fu+dDb/Xi8vYI0Fc/GyET+
/dSAp9wdq3E2f9Xr2QNA9enwx77p//NPCx2DRTysZTaUDePkNrkbIJpWYj4zL4RD
31oPM34PzeLqvNVcXsoZQt8tQDvnF04mwJUyz6RkNiNgqETb3FPmjKEW1iauJhBS
mcq7YXM3BWjBIlBDgJhpYBuOjoQqZGUvaopeFux7M2BCfmUozLcDAeKjoORi3M+p
aCklZ+FVqXEh3Yce5Ld+ClUmqRhWGxnuaNYhcX3PSrbUO4Q1d3z3EiOKcpkIxQcd
9zsguawWvehIbD9rStjfyYCb/XcOya+4ZrVayJ4Jdk2zBYHuiVBSVdamXUZXF8o9
jFY6K52Cxr8WrFFZFkE5EsG1pFRlQhZSYS1SCMubctZnI3vF9YgNnxwIddKJWJ/f
UeDdGRFLBCYRLAMnpNn6fVLXLOcYTG0fHYXngIDYHf58pzXT1/F55slxa5wQe0JM
fK7v5Tkvsb6PIdV7GNRkQMf+J8aiwey9TZE4PIYzD/plkwDJTjZ+EWOnukG4cYo2
x/yT4KHM47ZtyXBPlpuJJYviyPZGj5ueRrabGY7NL7jcv4MbMiaR/DWkKYE8/yyD
`protect END_PROTECTED
