`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpLx0IBiaCAoHGNHBh+4j3cn0b0i+M8f8vqjJ3oRGtWLh+jJEtdgtXXFx6vi/SKi
ukUKuZdsd+kiD6oxAWG7tUPbn+HYlyXOcyuVnZhqnnvRob16dO2Mm7EfyyYDoGwb
YvkMmNUDLX8by6DKg1fYtdCeQHTbkWiLtOL62gXcuVVtzZhsHpYxh2htFhItmiEC
/lEda5z24w9PXnuWspMFrkBpZhYyRqub/A+NsVBCOU7MvYFTi+6/FTjlzH6yEWxE
+4WtUWbTqc6FCgdRdBvsSNHJrgIZJ7EpoNRFPj4JvJp2SpGofov9+eQoTZdeX7Xi
EpZpnhvWP+hi+735BV4yX3eLOV0Hn5wIzh8EoLWFkbN1fhBeCroixEzLXrSrrxzA
AEMLpV3Vz2Y01/nIVuHc7Ljf8hzbnIoOU1NcQLgeBVaXBKnGvT1BRatGsmA+nqWp
TPl7Ml8tnAMvOcjqSD/H/wZsLqrkgBmcMuAIJXnu6vYg2Q6NS8TkEp4OV6asCtsX
LHTW0oHoTACK6oW+wdaI6dqDoXDnwxnjEyXnIDapiaK5zO2MFr176Si0/lc5RSXL
vamxztFCMdUieZKEWCrRbWHU3ReqbCzkcVyNAz8vrBH8VPtwR89iXl8Lskb1FMMO
vGDUm/hbumzi0Rn55eye7VRtEj6VVQsDyjkO2T6PoYJwvZI9rtrR6BpqN3SNQDb/
29zKLLCFPVQHLGHYmIrN2LleWbFzGY0d6zh3yS2lH1JcrZ9jNAQ2SxswV5+DH0sv
b1PgKHA7DGh2tfPKL8qQB8goB5TtpuM4xKQWecam2XZANtyIEFAlr7bzq8kaOWMu
DmOHJg9hO8chDxqn81+buD9YjS492k4hlJfVIAscUw8=
`protect END_PROTECTED
