`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WG0i+70Mb8iwuSumhtGvznQEfjt651WIPMF3vJcmBr18UYn3w/yGRL1S/ep6kdyO
c2TJDW5NfMvs89fti7GDX2Y1OlAryQnJqP/qDUieeFa86BE4Y79VRtgkoYFhR2w9
Kl8np83/6oTKAdqIiJJP4i40hSWA8TKMA3715NFJy5oEBsGr+4DSnfDCLcGvDf+c
dZ8b6zeAGv18q8aSIRGknsavM3L5dNT5Wz8fmbwdREF33I2UJH7q2tLwOcoUy96/
+lEe9M/wBCNIz6wu96JxohlIlkSR3OmPqLvlF/hgFMjh4l4EAPE4Cqw/Emw1S/+q
KYMflILCg5DuRwbYFZEtvP6sWNSb630v1Ccy7r4QA5WNk8DJgbUJIw6dtsydLY6S
ktIRXzfuu3cq8dfinoVXTHNTmTG4FvzrBVKcTStci3fHj7IceVG7XLMywNSIKcyO
n4x1rGjzPgW/2UQYFEGhv51Qd81Tvu82zoQTe2sQdtLSTNUbYSgP2cJO5Xqrs24m
mLQEYd8WxarSHAh31k4T6zvOyuGO2bL8kiOwePSPFmPKvrmZ5BmRGi6aN8YAHhmc
NUFZLq22JL+C79Q7WzX3DkZia3/CiFeE4zEhezzXSPKqWUof4jcIGxaZYVOv6N29
idXVaTq5q9c+m+Yf3ptuBsVM9VB0e7os8yBvLu7T8dXtBTSojGzskJuLR0pIU0m7
9VI/RWfIrBjg+iWpQ+bEKxkNm5UI+hr0+YEwDFgeGKshsYfsUELSTxlQWtnknK4w
XlfQpJbwmFgYKQG1/S7nPl9rRATMl9p9og1qXA2mMZPTUiNjcDC/4pu6s4ny7dKp
/0CShKi7iJZh0n8Z5icx7Ex4fj4n2mSJip6gsF5jeDxiQbW3FCgLEcPRNehce1yP
EfJpSYqm9MX/w01FXIZgSL3dvTCKrFzEeahY82qhzdVkJTBzt/p6nrzbcBxVWe3P
2HruFolaO/9ZTDILIsX1CAY23+HpxRn8f9FG60HDbGDx2itodQ/ZxoWr57PZn1Y/
kbdxppQTzGw4kwsTtRvSXJQOMd9uwt4mEVtZIvvwv3jGHO7hNMx2yWF334S+WgNw
rdQkLAsHaBZy7b8pP/wG+byzZBipKLt2KdYS/S3yD/TIj2t994CDG/oIhSUjSD+s
2ZMpTXq+g1TkKiqI/5dbpfDhfvwodaFCtDpLnw/LPYPTwZHVFYQmmrQH0PaSi305
mUlmZqdL81VfAHHyyGHNUaaLsXv8Ju1vbPnjB09gKTvyqHY8tPKjgR+/1SYTXbbb
HXhqHY6AkLAQbhI+WvCLNOOxy9AVVKfLV+hGoQBv0Lsok4HU9cnB+reZuS8DJGPU
iNkRgnn0nMZf16x73IiLfxcehiupVBKGKwLExVUxDanU11byJ38TSovJ2eCNay3r
mq6IyVafnpZVy4yjTWU0clmEiyO3ssSBMJ7V5/BugtQ7iz79nu19bvC8/qNmTjlK
3wZ2ZlaFzP5q/vEXZxFvIUA6p1fqOzBHELWl1p9u4mCK05F+2fJQkH/Wvn+TOqVV
Ck/43IA28NjHUve/WTFHZpD4cHNV2Fl6a45VK1SamD33UTi6lI7r54Ia+a5+hsm2
AtgDF6XKZaDDk8agu+FFbZjci4yv9wX1IVTMjC2egsE5idLFMuFFPo6xOFgjavei
w4zIzgnHL4m6DgeUhnMJTfOKIWsd7CMaX2RRhLugMSpk7EpNW3G25Gpi0XCrs75B
uqFMa+rmhxsvNcpYFPYM6DKNd899HiK4FTcrpTPKvUEi4cE0vZn91bPmc2BP2PiG
7SafkK4/xUUSwk57jCH6WbzEXupRdHfCx7zZfkWG6p/e1gzmSRYCpg2vQOMyL2U3
80l2pwKTRf6xX/ScR8dC1v6L+J6ZBqB/NFSuSczQ8FME+Ly97Dvt2MTGQDNTvCRN
thWhU//b26nNDccwJM4GP6Fx9laqCYAkEWmXdmQIvtSJgQn1gfUup2Or4fIHJAPx
nS+5CFmv0Z/KuwsaOieKXTlcCfT6WC2JohlB8einPDE4lv1zsg0xndYruRasfUJr
5ecRYUmGXeOadi7+qoT6n4V0wUfJBGdhyCxu3O38xlmyxpN/2eSp9LF1YD++cEEF
Rh9MBH1tyNTJ39ZVXzA4SUl3Sj1S7d6HG1i9bV4QBUtNdttZWHNKuCouetCzrz3q
7t89EjmWvmIokWDJkRd6sU1GhdM92/wUfirtn4CNXvycPb2rkbjmkGg4iDPT8hqo
VnIL2iTBrt18PTmsNZvSOyqNW1mIQsjimykfxTVuZxxMJbFoxWoiW9oNfUjp7p7g
rfHjcaj1r0hgsGQR4nNhHzBYA+8igETWjhOxPAjoJEbT9aRGK/WPEHYhXAGADAfQ
tTuys/pXWBOFXBCgfHFyZ1dTFnRxS/vT1PfmFtM7N7TM2lj5s/uY4ZXDLwnSxH+u
R74MGOOpeWdsAFdYOqlevzqQ9OBJNPV7k9L0llPUdxgZIyosoWGKucbAisymntQ8
ZvSRP8fPatXn3rhdQn1pbI0oMdbQyRC1z/Zye3b1y15axR3YA4dho1otX1QrNn8s
uXObuC9yUtoiibjdUkNwporlvu1uFmGyRB/rVDIy/sg6xRS+hoqxIBf6s8I+fQWZ
3jKfMjKpfPKVhx3SJ8G3e4mmuI0c2JV/RRErYnDf+0TwcrgZLIgobaihlwmYxzzG
4RqBjMVO8T9S5tPMkcDVEvkVL73Gb5Y2xxs85S0Nn84jWqGvM26zOf61BnGVfZ5q
fTzGETGOfut1NPsq47TPQM1/hozpIqMoP0WUe/Ar/5gD1X1t3rTPplIMYr59TpR5
wyHORiGkR3FfM4lk8DdiFE0WntvQt1Zg+ztVvbkamoLOajERf1cuvZ8zSWiWrB8E
2ORTn8Tu2H5ErWyZc0K1xrqMfgp58kVxjxjl3XMGDDIFHbP4eA6EhgkXU7iEkxU0
oyzhhpMSJ/g+8ZC9q1AyPbC/8MKkvd+hPKi0atZjf/fJzUxetjvO7MDwhxUA9qlf
ROJ7tI8DtfdTaLP94tb1LXSI3kUhmq0nFEVc20kNtfkXUsyEKKz9EIbzRCN+lcQ0
kou/bs5FOZT6rjsGuevjxtIWddAr6tP7KbBoOP50RwRrD5Wcj+dBidmeQNt+Qn/b
jyAjUORVH1jkb7OvMMy/cagkkFFEVoxmfXcQFZOlv7uP0UN1B2za5noEwUhAL2+a
ao10IOgORUDEOu8qSLdaHb+Oh2ezvVeW/s0PqAxdnadAE6lXWzCh3veg3HhhFaLU
hoKIVAEFliOkImu3hzFNiMC+C0YATqPGwLmNyyF3qOr/orjQ0Jm755VXMO7lXxXI
yJXo2+kQbdn2OkyhkvPOoUMg10zbPHdRNEnf1pe6E4+q1Tke7qtVUKvnR2JrHa+C
l8Jvv0/2vY+7fKUnBtmyIYNoncAeaTRHj3E1fXS5oPdCCzJMzFf+ypQmo3Y8Q/Ac
0n8AnXYSf8lcZcou37WEh6KrUqZ71QOGKvEuSLHjDt3pxlZzQpdzngU5I6+oGP77
3qgM8NU4b5eAKUBIdllhYazQl++YRRJX/3apB68xvYeyGqI6p6djNI8WlLuWfbni
9DylnM+N7dcU+JXA7XxW+mbbE4yalIjos4BM0jBIvwvg+5YP6wOR8Eah877ywyQe
xGiHIiKviP79evIrGH7i9zQnVMOgD2JI0SuEEiHJBvxzqKcK/BT4nQsrZzkAfDv+
wr8XwbZ338496sOt0FKMuqrvqPgQg+RdHzj6eYvqxjKvUqFbn2N69tXwoXQaQ+CR
NebIjRICi74b42S+J3tUgnjhn1rNxbUwk/FBCwCV6boLS+31Nll5q/dKQ9av+fCM
ehJ/eq+iWiGxu7ZIU2WrA6eit0KmGYkxRZN+VCQWoiaTp4JXimtwEJb5zGk97QmV
NZZiqeqnH8dcwhHgADRic0zxZ/Ojx36J/My27jesFRSqAVqwH7Cms2oUEZlm76TV
p+kSljXWO8N1IGkDJY4hBLqDS5lrWa8TKE6xJQm8voc90aKIS4wc64SH9IUdXrZb
BTNnKJjhx6T+ceA4YvSDP7TUsY/dBJgPVXx7oAHxX5Uo2WXu8ts8fW730kNaW1YP
tDnXRYUrcVfu6skp4I3E6pjkb0b0+TyowNF4BZB/rObWBzljoOd04ODXMCg5vLAc
`protect END_PROTECTED
