`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jHBM+eT2qja+Aa7RADx4MCvT//FrSmKlwfwHkLvr0bXQNdL5TGR1k+1/EtDFqcRa
ij1V7adxOLbLoh6UGO/KKwQ75YpOVnKfPt/AqTfKHb4fnva5h3w3x5YdQ5zXeyio
OX/xqbYGloH8W9w9p+penYWlJOhiakOf77hGccAbZCg+tx55wU7ArvsIEOihRAps
yAl1QrA4Sue+7iSqo53oTjRanYSlFOTMjptX0PkHV6Kjz/lR8xg/X/nui+FBmaJM
LTZ36m6hwQbqP3oomrRg74UHXpHLJWngsb77LU5mKflDhvQrGeSK4rRo2h/TcPtw
JZyCP9+CArn+6THkEc4gx7Y7W4xc9JfsSjP2M8KhhHFlhKH7P8cJlJDLOT1vzD4X
33P26OLG/SHHldYzK66bfeC23ljSdgpyD5qQXZhxggD2zVubOMSoYvepBgUztK15
MHxARhTfaWcXrfsC2uXFLCxyAkJpW2CRjM0tBDTG5X4av4+FLQlLgpy64fw+kuoc
0OeUyVC0I0JLDmC7IjUWmK/BOGOJ415zQbwqfH9QEFxTS9G16lxCTXlduiP7SPrl
c/L3cLvfRTm71uEU3acXtJSgx9C+DYZaxft1/ly2Fy40fwOolBNVcfiMoKBGU9l8
IQBQi2TuM8lyo7RGa0yatX8S78PN00p0JDRkj7eZdPeMwZSci1Y0hzT5HMrMkiSP
4SVBfFU39Kvw/O793xCQeVE9/K3jZbMkhylAWJDOIgflXna3axD0lrdpKvPbQUpj
cljwi/s0KiD5+YwVtPnMUvPOSvGVFcJYhHSAdD9DxM4ni9KqLar5EP9XmPO02ZAl
XNK08NUJdahUumh2cuQMY2XPHOw3sMI99/k6r+7e/4SqL8eoD2rDJXxVjN3hOC57
K9BBnpHfSTfsQvn5XB8iOolGMy4mfvg72mMmMAFwgkrExnpL4aSmsMBRLoMB2Khq
bn7iatvTZFt0chKklnvbGUfGZSrLq+iRKV3eX2j7dsCcRgOUXA9z3tlvEzHlYrjl
2K65paMCcFHFCrd/H8qzRAH7nFHFVRdq9u+4O0YIThQBcaV9CUXiIyVOAj0YGfV8
QzpdCYocNweruk5wmvIpz44yEnfG1sNryMPE7c2QpQLKpebF8F43SA+UF5cq/qnU
2VMdr/h3Kv9KZcU0+pXw8ux+PD0wjlDiPQCWZJLmG/Ff3/EyuHRXGKknRYy9+v6i
+//3lQbQGpZdXFsk2itSssIFn301a8w9lrbGnqil2Qyys7fih0I72QgZrUM/zFHm
Z/Yfq/2t2HUnX3t71gaBY3HdxUet3VkPEo1QSeYRlXtXMI8cZJq4zz5IXrG6hsuV
uoqR3K3BTxukOpEFgTTxrQSrpOnGG6EzoEhsDY/LP2d0zRYvYzzYMCsyviEmj6Io
MUF+dHQYQd4ylMXY35V63ZHLP7NxoxzWPmqRKpf/8GKm265WQJBA29uQLeEwTDsF
a1hFuZWiPFLw0LaSr8TpcAUxhmYZwO6ofaU5sE92wA9hAOIt8roBF5gJPeOW7R7l
/DtXT4LxWe2zE/+K1UBhgd+pyyhaIKFaA1k5kC8TohsqQwEESnRWqob/rmy3KLXl
N2xzE9JQOIB3ivqJSSzMhar/dcszHRzmxVek0e0FGgJ8clXwN32A3IvL5SgLYKKG
K6fWoXIWb9rXR5AUvBUpKp0SIVHGoziVLg7Dys+NPgUHAEePskaCJWuPMG6s6TOZ
478ZnZttpEjMUSuJ16x6yjqyWYz27J6yWaNYLwNtoVKOZ4HlmmtQkeCdsqMbefPJ
Sb0U0j4Pwt/BTWl05hPl4MfLRywdsFMf9l8YlG2Xn68vg9ATp/ldVAH2MZxyHUDW
g3K2VTEMtqsmfgKFi1v70T84HAkULVMtMcBQAyufEnirvYZLcf/9iS8xycE5f/ih
qdaACxMWDzXF605sQBC/HA==
`protect END_PROTECTED
