`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2RVNbvXUG0PWQuz51xpiUOe5+A7h7vEuFgbslCCL+daa0jUztNftuVYCf6UpS8uu
s2f4/kZzqT1GcWngeTUQFWllsAlkgKyNrqwVPWjtatdcTiGqJPOUm4NI+EbRudpg
K3NWVUJKk1WHW1+nYcXbhWJkZ1YA7kKDXuglIG3YOZOahSBU9O9UKHD5ju3dsc4x
tLYHkzzICRkIqZOyNK8ta8S+zLrKn0cNA2uGuHy3MZSC9XO5GFYb8gwP841tAEXc
5K4LbQua6i0Hh0byREzYdZwf3CJcHJ66A+nuDiucN2gitTeZGkq/iuZhx1B7RoXn
+eCZ6Gco7+cnwuYpfDFw57Qn+3vYyAZRbULrmnuBAZWQpC8oElt8hMxTZnV3qlyE
yN+GiZTi2VBERilg6Qwm15ltLfxx4Jygc3CNRZvofw0wcBa64DFRVIP3QuqIxa5k
IMoP78P4N8E1xhOae7/7lIPLgC64D59/sc0SCPBPFnFYdVwUQ1UYP3aiMSSVrDEI
E5xnvMEQfe1Ez0bQZ6cP+GFWkMvVGxFPVj16hH8EwWxm842JVOuvtB4yk80TDZDb
n8buuiRDVTzjqNQqEoZzhvjUXxUQxLhsiweoBPdc2h2zUsv1jJoPrHNH5B0Jx+6u
F/mq1p6BpEIFOb8Gyk/vxePXXu1yBjaFqs+CjLPACTYJ8dS4Vb3HsDdi/JUP4V/u
xgyRgwNvWibzsnAnRv/lazV+B1nDrPhVZ6Y4Eyy48t9BPOMpiS+xkrtLRkerza4J
Bge9y37oD+dhAb38pcrmEUllsxm7O9hbCdb0BlnnZq+CwpK1z+2WappOx8/RLIwy
VfCBKPb51nuf7ffV7tF6gKKe1jrYQdLbNpgppfgXU0jKgD5AiJfbb5Zkg7fx9t1b
H6k5wzKJwLpv1HBUDN6mA5U+9MDTjybXYLnhqfLoZcZT0g4+TiiLlHlaQYhO4oI5
5lOQ9rCjKsOTufdQG13q84Hgui+dlZ0xxydxrOS87vVB4cghLYyDS9rFPH4LAVj/
`protect END_PROTECTED
