`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9zkIRCSJ6Ya23U7aWANv0JLtQUYfa+As9bMCFZZRQFVJdT0jBCWJ2WAs9EEbyXx
ci0wX/7WGRwU9JFAnCSGWdkBxGbEDd8hrmnnGaAUKfwRouYiZ4kIFfFMvsHVtrDg
yoNY5vh8PGauB2FBXGj7fD2R/ChD618KsjEE/v6/jlDOLwXS7/wOFQ1kEffaUR3y
uISC7haLk5DwDVU8aJa/s21Qqk3r0JbXLoO2sxIFt6As1iFEm7iTV6amhZ2vjnPc
gS/97j6r6YOkJKRwXBRXBniakmD1p9yaLxFNR8gxNixRYi4DpNiOgAobqk5iXAk2
Nj0hkppRdo+0kxHADnlxJIrcuUgcRwV39Qh/05ctK51vd7G8Yd3V3hycfBFWbwGF
jbM+mfoOnRDfzdwoBH8WC7vLjeTkBJS2q64xlPyd6o1EEv5pwafpkK5+rhTbkf58
LmeX71aO2t4rMWqTNmuFM/+RQHlpnGbOmSRY/xoPVIpmNkXTphlXvRxPBkGLmxK1
gQnYe+gkhcja36vDOsoGBmZLUoi9mFWwrpk09zn+mhKRScrK3Boz3PPjWaLe6nOS
OOlXGDMD8mEvIFoFZ22lvYMPs9VMRK0stEeZ9hH101F9+lRSt10GX1pxSvrUMdpq
KqLblgZqN/8BdWuZWPYPk9kNRluuIPsEnmOw/CC3uOkrXdNzT+sbA7h9wfowpy0w
QDZ0YfYt5jMn7q5NipLQJA2V4R61Gn4RICOArMSLpSz+I9ec/53PKpldOZ7CBq6u
NrtwFB/NGOfDccbSg4zxVmXbSXRgLUKDxtQ6duvpxfoF2f+MqC4Gd/TaM6NPX9c0
FwCKmc6L00BdwDBc68Nq6liSiQiO0HP+1pxWzWn6bOcf464zXaKdLflP+JAYPgZl
taA2Q+i7CFIzMvKMNynGEUsS+iDlilDbUV89CaGu+kNhUX+qlWHQFAGR0kK5Pjwi
PFK3N8OZJ6BIZlYJvAdamvQLTUTGUV0FGLVXHQFRonMXiVQLHr7m317HXHgDX87M
UsLglb7K3FO7piMbY6nl50rKimhR3pIOH+NUX5kH/Tu0aQlxs0gMdQzihvp5BrlB
bsDitkLGQX+dR6g9VXgpD0RjIAOdo4HWV1RCRbWv72y8/hbOFChsG9qE9n4mvgIO
BNOPI1vNcAFxpN41phJw4qSG5+OatphYjCCcivix81Pgk4MeTi+KQudJiMo1S9vU
6HFYT6Gx/4pXYS4eC1TZ0GNJZ7ixDpXpwd9EBUwUCfGDlEFqacSvDHIdeuIwvsJl
Z0zOWT8UBR8l0eL2eOhGCxtt25AZVJ7tMw5CVZNfS/fbUI/Zb9lQf/mEnpP5olVG
3utolFf8JXtLDCmsGOg+W0UnmXzVEuPkH3ILS24Bp89MlIzGvj1BsPBdJGw4DNBd
nVKTeJka0XflhugAe42qJ0BEMusVnP725+tmPlXFyiY=
`protect END_PROTECTED
