`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9RmHOz4UeMftILaaZvcVR3xgdflrGJLK0DCJ+lrrumYlAIJMWzGAcoNC6b/JblTG
4di2F4xjh0rGSVZZ8WmhRuHo4luvkZJY+eJlcILiZPFnyBoDDILK3MTcDy0fVe5s
iEp2wmMGt+gJ/xUQDtzlN8SC+r5ZAlLqjRiWh1njMvAbuKWtP0ID3pIOXZW6f/bM
LS6aF+0sUH4vkWddrvERTGaypHqM1tfRGxHhHvPJAul5pgUR/DFoaJnypp3wVcPP
RUmyCVAQDoEMuhpBYx6bcf7AiejVT+9UsaEsBe/EzgECTZLYvGDjCNFcKMsdoAAB
+yP8oqP1fAOtYElOQp6LoZ3caiatJTUst+eRUf64ES7O6NvPjfkYP0SmgRfD9D2j
jdSam77dwOjm6RwtSQehZsdImE32ZKAxACOwPVaGMfQW8nm6SxsIzzT4iO8ZDyBD
XZ9werhdrbwqu5qh5nmAgXe+Y7q2y6hZj3TNaqJo2+COZzkQxDtiZqeTI7Gu99ts
o/nN3zyg9Rn0OvvJRie43MEfqdmHO7ntTeQBKPZDaTMfZtAB8CqlsUpO+2vZb+2X
W25FqLPNt5/7/nENfZ0d0Ch4BAjbMzJUzU0k/DJEopoyC10FeMVnoKioYBX8kCi7
hL7BWQKaaWX5Jj7bE9JTWXomXdlD6hpEO8EKR2A003R4s4ybFmzBtdhb7Vbts0rI
/Pn8ahaCQsm2pF75EdyKN7dLUdZnWmTM1B6pVzZvolifWN+qqctLWkDXCv8ekoXl
69hMtNLMNplrMNC6j2wU/aX5aK2homnUU/2Tc5MSzC+BD938R5Hfnclc4r8hovpS
bnOS0gDI4l2/Qm78IJRVas/Sms3H/nAZgOxF2r8IJoJnmAqqCBsQdGC+R5g2k2zd
x5WVBEoMB3NhVwan0gF2A4ZatcLueVm9+75zk5RBKFGg0TF8Q5uVO06pBmuCp1sR
GvcchtM61SvNERTb+/Hm3P13iboTF4XPZCuvG5UdSmJEINHLtjdE+nIQhzw1TGMC
7AAiG882zyfYXPEfNbMscDzNXft8ygvD8OfD4GbQLDPuuKamUBrRCvBXx1RneZK4
7nYBWllIhgc/voYcpmv1SqKd9GXGNi2Gdqrl6BN6c7/bb9fpuHM+3tu69qY9YPy2
es9ygUUyJozjQJOXx6pkhJYS0rVxY91SxrkEektla6Zhwv9RNFzBoP6uu+lUppUk
LO341uz74S577jIj1nFLOqa/6jVER2JqYY7wurzYutS1mJKfyKFmFqeGN1LNqtlK
KW88F4BCgIZmqXMeHyq8Ih3qjjYIwnZwMkN7Xm5MiAt+Jz9DdzK5gTe1jjaXAdvY
DgZnYG5Cxq3tqN6oUNC09/ezk+XRvEVKjD0YL9ozb2Em7UAwfUe4ls+sItcZ0XNF
OiVQCjPi0kTUUkVC8+HzgTtdWc475NmgE8ZeBgAvxWqiKAPOwWDkAm3I4bM8I+sb
rPYVsVC6bE0de0X8ds0ZJvJQl40EH0JRGBzADqtwb6KteWw1QcftNbKCAV80FNhd
chKqxBYbU8CCuK4Hgt46MtcXPvgfdo0uNV8qSq3BOLksGMMooQx2Jb4j+5pRA631
aJPxWIYTdpCdefO6353sxGAQjx94JA+cjLcMXVxe+u2ZW74Ngr2LAoDDHHPrRzS/
cPhWG+Y4zueIJSabTwrljJZDSzOCx3UOjOnkVnNq97Q1wek9cbc0as/A+vSOT5lU
QMvRtdcidByz4/Z3GaiAEdlOznzJQlkFXIrj4WO+edSBysfaeUkqPmwNRA1JvPmM
ExHg0rzzQTsEPpGRk8gHPgApNtI569xKVCNF9GF4SsicawEWGLGax3YWSoWY2cBq
7g3VfaBVTkh8zQT5NoZFrzWSH5ynTdLC08eAaV0d7TU1mE5094Oov6olQuR/73tq
T7fIJjOPLyM86my7LMhWNhZIWr7eM1LZnWGbhCfvZ4qPcWLMbWEB8Kaq8ElpQerE
XPwRoAtUHejVDPC3nHSjjil6qc5ZFrlqf2gcsPR9biXuJMTH6dh9gANPBbYjVUlv
Do/29qE9O7UuEek9me4X0Cw/aVHPw0qOlVxcJ1efZ/kJ9DPszDCxz08R2nfNPkS3
VjeJTcCsoYv9uxcLyRpXo8IlY3NPAr5F3Rd3SrPMC6jvdQ8dPs4bHyvm41fBJxPR
xyzyY9QBjMnKX/7BcoD11c5g2dnZyLZbzfNhBNpwEgAFPyDY95UfEA+YETcPE1Qg
zBwSclkGrzQrb7dO0+0oqUXTmdGfZv4mtW7JvpU/tLcQUFjxVvvI0fMkbyPebev3
nFr37meLiARjpMsBLRNdvbMyTQlmbA8FI80K99dAhn+YSvafG2QSwzm0Fo9SAark
LRrNu5c0rTfwynBRT/rJZBXF0M5F+XyuEn+CMq0Q5NKAsnsc1rki/IxK2M9x1fAu
f3+Cfzwm894tUUk9WtHLa/PJ9FbQI5nAXZV9Ru29Ywh0vNBmQ6w1euBGp3Dp5MxD
C5wKxd/Im+tXHGxg/BnEewau3Lgzkstl9u5Yumz/w7MtbdT90kPJNNBuMa9zMgHS
lz+z1SZ4H+Cu/quIwhp00PwQJW4Y5Y0byz82i6fR1AQIjR07obcCVtcVe9E6tZuG
i64Am5H9cGNmfsFNiwwFjGCTfhSeTRJrlGs/V1V1xOGgYcjoM823ieMAZ+BThPhw
BOdCNs22BZJL0aFotWBb/IWQ4lD6YeCCShHL1W6FKs736yMKXeMaaxJXNebDo4Aq
9JFAXKXrZhHgUzQqGl1RQb//maDNuHXfUHpPFjhTBaxzQG7eauvbusiZdmhT7XBk
gAqJCkhaNtciCA4sfapzhihFNpvmy8ILDPGdO5nbp1AN9esjF0qpfRHlb4xoUpQ8
tH7KEpUed9J2rCX0DWUfPIODouGHM0cTn9sSUi81J86km5o1KGxry3UX/2NvYLEJ
uHhX3Q2L1HxBKhc6S/PYIVn9xPxR8QrP7eklqWDzOPs2UVG2q4osLR/qEa14ppVw
yAEGc2iquhClxb4dKWdaQDSEG3pW1vkjZD/ekAOTai4i7oO4u1MxyHjfhttoCiyn
BETMXX3IZAZ7pngMNTfUFidnSR0gxymE8SygNoaI20CQAMXSuCqekWTygoUIuV2v
Sihxq/bBUZz2PyePB3uketSXR8q6K6O9f5QWz9pr+W4aejL94odP4xUEZEIdt+Zh
0crDLySbQqhiYw6DscZhQDcWJUTCExItw2vzbwOxF5EO7XJ3hzg2fqNCWIf0XfU8
3A6y/Kr9O13BqVE7MUGVH1zyelNgKxU0rwSKgoA8oUGc/AEYYwk9/hs+PRfUJ0vZ
uIwBCw4N5LsQcR664q4xJOLQZPr7RpHuUg6vxe+93bQgnUL/BjCkEfIw/9upsjLp
d4632wdD3GFAvrKIWx5Z9qCSFOwncUUdxMs6NrfvlL05HXOrQ18WErXowGkJM/t1
AW6IS6i0NyhZv2kpxc8RSy1z4aAcS5QMk6NdnkTMMIYY7JMQEwesbEyUxVDtAVUE
tned94ZSDBE3AYpjv1/Qty/RSixs6Qwp+nwb9A/NiV28WsG1XA186qG7a9GdAKOZ
jUvXlTYJXGifDR+n0w33A14/3qexLgbx7fnBxxPyRxZBEYVF/LVw4wfZTXW6yjB6
z6yxGxZQCaGlvEdG6ihxG7kNc3tx5Vm+rzR4WlgMoD0ldza0iQoHMNUnZGD1Hx2O
GoUl3xQ4HMkIskHbf2KPEyqKwO9TO66MdU92e1rYdYxU7eRPFUMQy/RsO+E3l7w1
hgPfpXH6CchEGP3wTpOxd63LvtacmhJ/bSF9HzVbxG3P16IIFt8Mywf+piUGiwlt
zmPJucI/RBUJkNrOxilJ/it0NFA+QWrSGjp3G3x0daGXz8BMIeK+/XeJ1hr9XUyW
1lY58bcfYoZGdRYfouHh6V5azq+TCEHkPxmMjdTFAN8YMYChPr+OHTACy8MLbjdv
3RnLo8qPby289slfsauRvMfbb5eZ4329o2uunSodCUM3vZvYJIr0IgG/vpNbAjJ2
V4T8/pBR096LBR5RhG8CYu9YEvbGrGyVmEbx+I4GrPLh/AhX2naAvQe3MgmWR2K6
wG+qPkTMT4GNygTmfomeIHGXmN2WBNkixp0iGOjBtYefEKJB55hkJvOb7q0qBA+R
`protect END_PROTECTED
