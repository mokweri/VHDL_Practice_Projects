`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xLgRpoBZv2jxvJvlq/K8DZXbNY7Ux5nFhq8/TM6pjmcrQPOqnlfF3Ez+cZORC5Cn
cDSIRT827/7bpG1MzsZU27FiynPiX4KUWxnMSQAi9Jxnfad0j2zWP1MSmE4cXUOz
vCCpEpAVlcytkAU1R8Y9GjEwvDZ112ho5LpVcZ99Bmr5X1pV2OdaDMGQ0vByaChP
9wdLVtmTnl3SQSaeGM/UfZEaLO2KpmijKr8XSiP8YTHPYLrOiyEL8lQJ44UcegzN
++dVvpTOR8dUPvtwMgt/IVc9UmuMV+ovNqmVnwfJkoPkPfhYrsgnJghKGC1978CV
R7wjhwl6di/yDfJM9yc6jILtyUX5MBs7Vb02Im7P4errhUpr5VJnAFDBL0dxCAMG
0et164A4eOAId4biaufKQHxY0mufJ2u+BdUuL9JyWAwTzzBoS7aVmjoSJHjesVSE
mMVk2MWRg8weA6GzeT1d2kjkHqApeLmcTzyrrcSo1J4qtNPs4J9y+lmHa5pKNXB3
1xsuieGBG5k4eD2HGB4sIAYT4Dm8Q7q+Ht8yPAhGe079kmYoPN16B/WKHvejQvZI
ReGL3zjso0jore64uAgNxBGJ6TnCA91llAg1kOEP8nXywOqT+tQoPUj1Sup43cY5
L2FniH81kiXQFoD9eURxzzl1h1g8KX8PHOLl/9rioIlILFYTcz17f4B+WR9WeF8U
iTSXv2z0utXBJzQWtcyXuLTED/vk/f766XtQlIW3sMdGKrcrTbfwDYoqBBEZ01xi
jON+9eW0sF0ANpN9Ul+SeV2MPBHRuWG/9QqYAokFP9s0Iz2uTTKOKKDbNFvw6NbX
GODeyvHYNLKzOgRPi5ckgfMxvjUoFvF+9qjfpVCfUBVYF/2HQPTk6RRYqw/BxHQ8
7YS2v5nCNFGJiAvScKfO9JUhZLn+jVKxIpkgHl+ZPK/ongRk2kz3BUyb+IptYR6j
aYecVcYQ0StSG322xxY7ZAn4BYKEEjlw69h4yMtRG+RwXjb3T1E9u/Vy5cfBhoVf
SJ7DpDBTjM2EjeomfBUpKsNd9qJDsiG2hd+d72qyAwGnZfg+Z5614/FM8mkD3XXl
XaCtlgfDB1GfljJ2sX+qvJqpso5T0mpZcHmkI5Wj77fc+C5xxXpvqHcFEPyTQ12l
JUtfWIGX8fWvhQ7HcdalRt0BV30ybmepylvSi2Z0TTlHpeghFvhUth58VOHG6yE/
3I7K6uIu2rIT26CVP5XmO89H0zoFwLkZsSgRONd9SD2GfBCxUJ/ykWhdbAR6TSB3
xg93yJ/ZZ5NZXCnfANsbo16f4HWRamQT9Mq40Svs++HMj+BvUYHuEQYu2jMIv89e
8P6V9kwJPZWESX2xjKwkQOoV6ZmOmFgGDg1hs8JXDvAl9783Zn6j2MWafOWTwRwP
1+YR8aDfn0OMHpeDTedjLGFD0+5pXuig8NX2sjT7OlSkFsLiWaOsq0pYxLDZHF/G
LNlKRfgbHk2TBjvCvoPEfYc1KgdN6FTEOMA2uIyu0SD2KDThnIqRQTjtpDuQJzEK
kNlb7z4MRF6av6K80ngE+mJm7zaUzw8ivRUDV94Fp3BsEi0MNdz38MuMnjsDnZDO
2JQVrV2Zn1lyx7XfaXA5v/ZPSM5Da+0qCVcE8VB5+XeIS6lSbE+jlFhLa1V9Umpb
p7hlV0fwvysZgwNdmkBz4s/RBuEKtb7fE0NP6ZPizOjCvAEy7GT4ZS52krZUu5nt
1v0OXw9FDgZ5IGhR80hy8WxOzshP73ai7baHH7sAaQt2hsZIQSQfUr2POhzIECb0
cPnNy3djrTUIxW3EksGCMakHa9wcSXZJ3o7Oopq5lcege2g9anugRWQqJu36hJJL
pSdZn/ngyP8cnJxZPFbvqQUnuPdq90Rt1LMtM5cp+zWjLFE8oO6MKM+kfAjfqijY
olmNryqJuWHtHJdzv/uiEUG6K1OfmV9Y7aKgQ2LAMER3/3Z/x7xmNQTsLuuTI4p3
XvwK4w+wKajUhGtf1prmTCr8Y+LYkN2ldSbL55V+eoiSU7GiHRI1G64ayUiOI90F
1tZZbpJiBHQ6twXzGtKk7ne7on1+WsRmgtIRsdqfI+Q0MYEx4I8+uJF486nKwuro
bTny+UT6JdT7H5aAcRaIcQ7/gdt7izhnHfWu1NppAEGOrSOQaHLg7NR63Med7Jm8
dxXs+6sjCREEDmHQDqlP74eJBv8b/Ppe3x14qiv65805edC1ITwJsBf99LWJJz6Q
F3Bj83mWN1aIxWPQKKmlCrRo3qmmieNgnSjlOzmCvdU+3Bz05mhMiiPbaYJre1j3
Ka4rqNic3pEKZhplf5/dgDimWuvnzcBTPgsV0YvH5Dkjp9k4WTqAV9ZtjFIh3NbM
OczD0PsBUnHXAVs79wtiDnaBUwBbWjgwcRU4AsLeC8fPmXNmqzWPCjQnD4fVvrut
2Ji38wte9HVp3rIxf5Y7mdhugfkzd4yrQGqPLJmQ0Yl6e/ZMlV+7HCmkMobnJVwd
3VfsdszxdqM8w6mpuazJHUIpGDSQ1I3nJrNj7bEkmlrupDUvLAZ8zy8h1h8meD3l
CS8L0NJrV4ITHmpQLWhxbld+wHEc6mkDxABcuTO6XPficUsrMduf6XG2G3aQZJCH
7Vogbfy9W5ALobCchNKjU5z0COhx3rosnWfjAaj4i8OfH9dDfmGExAoINA4PuX6F
3Ua6g7jkOYXaey8AyXD41BW/czqV+/iGr28q3eUbjvEtbbk9a5mV2FetjqWa/XkF
QtbACWvSYnzt5/cq5QAUdAnJdDLH1XiWCDx9XtmF0qpGfnkL/SdRPacBY0nJ4BcS
Q/ZE06KYhb9ZofhhdJPbVZcakMw3cdw0t2i1akncQoHewQN8PnPvKCrtm6+tq2as
Lv11wN4IjwC9X4yu8ANmtfrPN1sSU1+CBbNDgr7I8eAOdwUGcoUiFsgh26bFapui
JouQN6b3uHlR//+NVBMHqs/W0GXn1frzTkJG62DwZ8Dq8risiepUv8DWfbA+scJV
iG3M7nwf1G/g12wutm937kOT/YdJWVvrxBx/7hVp3m+/KIWE8pXSMhCK8kukggdc
RDx5FFOdO36WsPPQe0wDnW6P5Dnj+5h5wJ1yHp2y8J0OuEVXI6V3ELZ1JjOEm4YK
RelKG6vNQfJxuOCYHzVLzfc/kP4+0M0G0XVaSwx9Qu4/iv7mvlO+kL1x+Z7qpVXr
GSl4Zb9e+Rrr7LTr/m/mMdfghPo/t1rezHfOOAlhNqEVO+rJDQalLufIfOTgInrh
ryUfgS8yGQOP+rmEA+vB2fuJsMymWzAIbNtA2l76unIB8/owZeKaIzxKsBB4iarl
D52Mc5b4dcw+ypR4iig/yhQp2UdupfSW2apci/5oYSh91uQrYTJtMypHTYcUBTyv
`protect END_PROTECTED
