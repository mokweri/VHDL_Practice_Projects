`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28COj0hpIpr0Z4E/9Czt0xKxqIZFJExSzxc6UIxBY8jYXCGsVYqWmyCrTx+yz6f/
/c+DoELfaEBpTPWJWgUbWgL6c6rrAwPUnYGbrWHumBM+KSNY3LdKKUh5bz0KsGZW
dBBbebDZqAaWM4pJi9ZAWt0ZkQIUhk44UjGH/I3mkpvKFyyjYvMqIWNp3ASR8zVp
vHn4BwLHVt/6g77dDbs8jnvmM/Fbn0cBBYCudtfq9a7s9Dvownxqao6oLb4otw4I
Vw6LREP3svKxQrsDkzFgMpWQvSJMig7fqDTt5IO+7xj6Px/BCOIgkV2AkVXjQG5H
q6hTYEBrtkYsSQf6wU1OBs2pox6+kgU+cRcr41MVJlgRkRwleyMadfM/CLdMf8Hj
RHOws0JeUxm4eMqsRnAjmbBLY/4r4wshceBAC8qs9YX2YCnV3PKZ2tB9ZjdUoHDK
VMu8h8qyeemucRD5YKMc+Ywc8X3r71ikKvO4/j7quzk12OvBW/CDFTmG/7L9MEsS
5oCGOGb4sVwuN8eDUfg3238y1KGgVKA4D8JKmuBxA54MXlWsdrwR76lR929zR6au
TT29EBuHeug/GJtPaoyk78/4jHn02ujBT1yyRXkjfw9uUfrb8PcO4uB9csrSbb0I
t32ZYmGxgCr9xR/GsEG9LebxbXiSL4MlPjwmcZ0HxkIXEw4exL5vLi3/dH152gsg
SKmMNKH8vY3dOxN+hA6M8+P7Abf8D0L8lm2o/R8dsh4xF1uCSlARBTbnssrLuNP2
Oc1ClXX+rYr4W9cplMWe81IGfVg69bOYfA5dj9eZuJYO5cm9X35SW7CQKYs2/V9N
OhpxmLJMFCXzUvCu0oXYUj1BYK4WswYKF3eLpAFz8FhfyM76K0+maU98QLwsU+Sg
1tpPX03hv1wwjmZpXuz3ylOn6zJkHIW3DpsbN+bZ1DqjmBL3ENq5af0Rymq/KqKk
bA29dEmSLjOa3ImDAkT75Qe+J1a+/8E3pP99RqHW0cQ2P+LGT0YGcfHpM5aRmYPy
nIyzWyhl0bXhQvrDM7fmPWlVvJf4NBvHzx+Kre2Kz8SYz+oY4cGJackvNiLxrucn
NvvJ+jTUuZPoc/p5WOGtLp1+PgciMZr7h7+5cu2CLnJeLw2kD7GcNDCT3aSdRIdO
0e2ySQRW2YwPXNmVp90ZxgZL7Svsxbq2KeuShaORBP2/BR1gfaIdBEDRvaiCsdxB
ntv1FuTG21+qezDWUALvUAkLGBPq4CveVHY1fRJnFFW5fOx5EHG+6T3UmZVu8ZyW
WSNKAJu9jwCNmHrgniAPv3mhxtCtUyX+KsQr0cCHX+3Ivo59mxfJkyppsedguW0T
bPUbLmyPwkZ9pilMy+wYQ54smkgJf5cfL/ttKr0PV+I+TzgCsdsbQydfsx+BE3kF
BXvBmnBYTATDjeY+QzXjsBk6SfdpjDBrY+SpEbY8CwZjCXBKOxK3hKsHsLmN/D6J
aZN557vWUVDBWVWlCZM3f9fnA4zX58O9LACKrImMjJOYz+TOBqCTwWorx0FsOR4Z
59kvDiSOPs7yLkqDmPFFS3DO9KJIyRDliQ5c0QnxMAPFgHkKxkccRiLBPfUZ0JHs
lFiwYk8BYjubpqST809QeSr1VqF3/zElaf6CNnJfUw3aekl9fX0ch0Mp2hnjRozw
JyteVJaEHAzSMSDpiR+iW5P+BADujR3icbavqyVaG/VKFqH6zuA5Czk6eubFC51N
pfhFc3bqH5edbwlPB1/Qz5UMUxNyimLmfCNmK2KeGpfuN5P6gdhm8F7GdsvhuiTi
Jjh5m/xnA7LAN85BmCmnDgmmT0WutsYAqxieEFafZH545gdJ0fnQ6A/D3Vhqhars
bqzfEuD9BiFSHPhYzLNOLxEP+Q9uFylMbe45sM3KqbceO/L9K501g1axZxo/L+w0
p1F2hiWK6KZU6wQflQNzV0oXILjZx/MRvAzE+v1Z5mJOv2KMDa3ZG0rRIhEmVfEv
xf5aCJNBCT2bOnudyc4PIYD6vsnbhmRvwrka6aDk113fZ1lqtQLTGgoZSiLmwkjF
7CFUZAAubrwrmuXki6iaqq2WMi5K01MRbjnBMMa01vJg1V70dgj2P8UaCOp52Uv5
/CG7HIDOJtyjcnM6b1HZXmAoYdPe4168qjF9OTS/rnOKEJBkagOiYGsSIjgm3VbM
UrOq4uCf9Rkcp+rhUsaBPeAxx5shfXFWnQxCfYRqAdIKOvw8ht9Z79j+8FpWVqOS
gKsilF32+npWH02jl99MjlG6pSgkUjf6B97e0YnC9lyaOIuj7IcUMmEDwcd85Nor
nbsElyX2kAZS3LwbbhTIspFKZFV/UTzBzbWIitLjMCtgaD3/a8h/AAViypZCppYs
LRQReVg98/VEUsABGBQjP9AYIuj/ueGf1i4gp0rSeznDuIjhkhWH78bfSIpOKA2o
RHyKtRtp1qhmlQg4o0CR4IJAbQlVwMcarrTBHVUel3GRdh+9MAPdj2yKsMdk5jK1
mJLTBCZZ4w/AMg5sRAKlBcYLrHAo9jdxFy1l6SFAtVseb1asqTRDg4cCGiHDMI1w
zSvdHpfc32XIbbClT8uAoAbn+xuJfDYfLowifXcDjRTTA3RpgJp64ZDboLkTS+nW
AvLogRZcGQX2Z9/Y62V5ewvOYmh1H4KISY7jdnJbZcs8QF50qrA57SiT4wupanMx
Xc5pGC72A4sfN3T35NKxLI0f8C/XBZ0t5KFeD16j5nuogT/FuYEtLdPgJDvluOtD
jgAQaHjlRae0KSt+wGFTKNelZ3mDdwhwf89pvoO6jfJ5fIJhihQ8KqlNYohDCtrk
a452UzKb9Q3ssvdFexA+DftnosdC/vUJwX9jHQOs9M/Vj4xgZLF6EtUescmhanPN
bdgAn6iXtXQI59ro5lne3XzDl7zp9eVIAr1qtTOwzlYPj+a6nE96MO9h/iOlgLxr
/yiMpom95wlbYGmD+se7vPXKaDOdxx4K44hWXtufDjpSuAx7gsXVPwTO+bSqi1i5
S9MPdtKxnBQoRZ7mgsJAsLf0lhF5J9K3bQZsJn6O3RPt/Mthzx7ghWY7e5QnsD9+
bgNsa0KH4L1pGJn+qXykjPDhGZHkTupquCKZCSdJ7vChyw49JfO+OQDGt9mAfHRZ
PPIPxDzPmZqmkTEcsDUVXc20e5w0tG6I50Z00HS8J5J95D0EjGJFxkCaf3vk0zcQ
Gtq8la3dH14vexOPbjGTVbnS85oszCIfF3gq6qggjbS4yV9/Y7NcJ/djMFIr8qcJ
AzWwe9vtBIPG7MQAs+Qzqw==
`protect END_PROTECTED
