`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tTIqYfJT/JEEg4Ok1JYR0lSohr+NCiuzSF4aNazIkIFDXnrDx4cq+qHua/W5ANLr
11/ozj2LS1p3UsUegmAqUOp84FThwAI2n5s+XutRbAxgdelSpHOpPK/HKqe9XKgY
PkXa2XDQ/2nuUxtEGIpRar4kHYMzVOlWu3bx+SjLxuuSd7CvIJNQ95gsswaYg/gk
OQ95rEP8vk2Qpg+R1IFeWDOZ1RpqB264Z8xFApidLgmo3fZajvYjw0qXxAKo3ia0
8UtP72qVpTZGOx/xB5e3GRja7PC2Zce7q57wKdMkLbr9tbIdWIWMMJNA5v5Zf+u7
w+v29jUpNJd1IH89CF8n0Awg6qOqXVlNQPnm1koLe23pNYFIQvMm3LXSFMEsiNsV
qbs2Wc2PCHq91MjYyyvaeKKAdH8RG2djmQYTpJCxBhVNfvLsxATqY5Y1ZhW81P4I
94Q7BFF6L0sfhVqCUXOQx3Zx5GwqalXZ9n7Uy8r2s5AiuVeEr2IhSgGDZMS4z2dR
gEaMyBh6hExpAk2ZGvmFy0cK+1QE7ZO8Z9OnWU0ouq6BISQcNt0iwhxx6ueNi+5d
jAQiD3dLGZgVFBD9ckY0YzLnyufDQksozPHOcw84dKe3NUWzoaWgmW6424OwWvrv
LIdPXObCnKsNnrUY67CL4owScK7q61Zu+n7LE/7BovU=
`protect END_PROTECTED
