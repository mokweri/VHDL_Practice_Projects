`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+UHOAXvOKf6C5pCoJOQI0OMnrNJn8g1ZvAIMFGjyNusfE7rWrD+PJiMmmzF6cum
6+nIg1sVhdEGyBIwxNK+SxamBT+fcX70awcAXX695av1nfGgj3CXRqRoBiNUG5/d
Mnxbj9/N1q2FQWTTtXLpWlhSH4XpVRGFNVBggAX2aX8eZknHCTlhEbuk9kSxpwTZ
GUo0txNUCtkNJw9XPjcYVV2UH+SfLhCi9AZTS8hJ/FL/oYgRjaCrhpcBZtLrDIlc
KsKZjFMCol+X5Joj29fb2m71+n4KondlTDGHthxF/oeRiFLDNyfp6ZF5eMuQhfqF
pjDFtyU/cmiQJB7HAZKm0+dhKjdhk0huwooZi7sMqGEtTvaTv5B6IusYAHgSniTA
4dZLQdLmgYZ4sYrG1Jh9hanXAYGzHJF9D4sPdRQ+ykYdxNVyG2eGbqss2g6tiA2m
ziZkuUbcPsq9Fenx3PE1harOkltMmBQ9AvFNY5bjHRjiy7DrR1T+jQ0/8JKqELTq
tHVEVgHFckYY4mSK85o+uA85iv6wKIjgcP8QQDuSdicax+vrLoA7h2Dp44r6Sdx2
PV90/nxWtH/OaesF+WAEqWHorHjcHG1nZf57DNavDCSDlbfa4Y5VsWc2y56wDKiC
WsOrRAy/PPR7HFhHpp3yHSFiaP7PoFjFLivuMN1FFbGoQuMaozs6XvDcqFZv1AxL
YJlm88O/Ce9ZKd3CLrq6Bmr0cBZ+umqozzF/7EPZfWLurBLhf8j3OBa8rG8ueWOJ
TikeRhsqHJIAr2ZAg72KZ7Sv1pCxRIkdqRdkPEbg/Mrj1v/TPoOJBsWAL83TJfty
a3FNd56cG2n1kAFfm7XCQnfehRwMjeCP8NySi7nnGumsJPbCyA2bY/L1lUwacTrw
8qO8T7KShD1j3D3M0BhdHl+GBiOUAlBd9LGBblnGbmd+CfpUwMlDo5ikYnDMQF8r
IYgFVSCYhPdfPGWhmtFxctfz4qeQyXCDueHk2swRm34epItWrVrBhZD07mn332Iz
xNTxzhg7b0dkzrZxcFSQaJZ+fO7QO4GSagr8KttqfNfZp2qCJwF2i0whd3YWpPcq
4fDkgacBIpHhVAl9/7dMFcU3/j+BKX/kxjZyGAOLo4BshW+OBgwj+z6DSxWwF27T
lQNeya+nr3Z/92OQO/u7jJSD4Zbx1ItoGCRyuJLa0pz17dRAhVKgWQBeZRsvLeBy
J0Ly6F8pDALhoPkPrRcl6bWr9THKN6FfC3WHzMXE9R8wWkd2Ih8MXVOjSPaxkzNy
gfTNmH6NQJJCHTgKSaoabTMJP0VknqhZ427+RshDzSqKXGFB8qqGYOFBsg4G4soD
jWSM8UYLPJpFEg4UtwrA2C7/2VSvMms96NI/T9vSDq7mMD8UqHDH1VXHVTtm3avV
mCJjFOs00K8pMVw2y1sQabdnUK8Ey4I85lir47LulXYfCWmcbdqCleua4vKqG+98
0f2qp1vJK1nxWQwrNAian0mp47Iyp9w1pYdLBOwz8SrocXb1zTu+xAKfHrDTLrpv
mKHe0wspGx+LqDkio3VydiZTGLu7X14mxZinAAs0HhJmlRLAmQrn0vSJwZrnwHZD
SkoI1W0oFSBmSe+Uc7l5UZOAECTa1BCVQuI4k6PxnBal9rmu7uJFH8pvEg2MrkTM
Rw+pY0YOAo7yf9kFXBt3FChg3hAGZVX2LNY1zOdoiJdCA0tN+wtS1Z9mkmDDINaQ
tix4/oX6C+CtHaSs0CTqTCQDKJoLH607zPRS4Ofk+gBzH7oM2SE25+LQ7SkaZzzJ
NIH18mv5LpiF81vi3PkiozXuXj8L1d3GfXY5U9H8T9mpsG0WrCRoNcKiTGLo9dj+
f6zKl5UrZqvzOcAcSJRf2sT0p3vddrDVcevpgSSFQfq5EKGGvcmH3blw1jsC1m8G
GMnlPJhUhXKDnQPWaZ+6zvpzhKng93DPYgNVNwKPJTL24oyRvRFmU/iDN5P9KFqY
gKW9vnM+PaTuSXavDwAdzDNwSekb4idNfFd8H1iVm+AkjZJTwNVfTf5ijTc1iiGl
qIM9mQFfR9oNwgv+iIYp3exXnOKHEZ+4enLwx9seYSgyffyiCIUD9S5tfKTP//fc
E1fGGEtfq0BTXPuTMWvsymYSESeyzvF5VDIbqCcGfBjUKRT6jcCu2Co7MWIJEHEa
YCTpgZIsfRat5W/wxZ03rzr3J2xikgYITuK7o2folYv/7rM3vgghrnzfcbGl1XtJ
T514epJuUDSfa5G220IxPtCdb13r3wgIcZUSCOJ8JZFgOdblEsPWRgV4602CnBrC
dYPSZDlGVnDXuUS7L2ITkWcEjNVUrfqdMz5M25i2E4xRCXC9lv8p1PgyqGXByByS
uDDuekovl01hL8TRQPlh0KAytUGjh0VJXyyetNfSvvLK/TkQEKFBfa0gU3SrHBNr
fCysv7yZb9nby+9DLwEIhYxMXfhjaZoZMPYPNNhCjvcq0qvWruhXAMclwyBrzsns
/uCTINkDqfBOYlWLPM5o2We11AeigJ0z0tMBxlDZJqJbotbnDQ6ONrXXdofK3QPr
dOdQ/+8GtMSCc/NomoXUo37aYAc1dsOoHDYQG+gJTHJ5Myjru4GUi4jWHNjOPk0y
bro+b52Olth1il3Xlsq0R0PmgKEQpTl6N9Z0IQIE5nqVS+TcJZktsP9pJ9qtytmf
KpsZsnZs5nYpTvc4ISz5izu8unOH7pnT1M/MNMft32dlnkVR9dTSlDk3FPgzaDoK
7OyTbXI0pi6DSKIHBYKQGP4JI3cCvL2WuSnJnDwACI2Y5IPCO7bMxpn2jR/LN6Ah
D2uF9oupzTlTRg9lSvWiY9t8hrjNf+psI3CWNG0O+QfVj3kbp4XLIjEApaPFhQbM
hLxHRACVX/6YV7u7kw/GWaLe90hYyQPmKhDVDM9YsCBYj99OWFXZKMX+NFfmy6HZ
DqqEN1Fw/YrtHHj9MObsy1d11l7aKB/sczB61rR4ONw=
`protect END_PROTECTED
