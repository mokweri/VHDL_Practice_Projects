`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y7qmXy14Q1z0m/vMChOF537knuMnx7X73ninfd5m7Gk0jGPJHjnLbhdX4qSzShQk
KgLtIw5kHYXE0EgI/mp2JyZnQ7JloQhOpJxLe89aWvgu4rW/3nFAnU7Q3koSGn9U
Z+FUPU+fn3Bb4TEBR8TBwkmPqUcqcjbtoUd1vPyOg3gndWmzMsvW5BRQe/9WRgf0
tKIMIEiLZwlVPJnnVJ5PCmYeT2ALNnIzIwHo5csa4JoLKy5PJcpqNrUOTXtiCjbM
vxg+GZ/cVObXcqUDYVQBDJ4arKvn44BiFpl5sjA/qJRGtip+zhlLSHTjWk6hc9Yn
giYFjGYm5KsfmL16A+uz1KL3FSmH2Vp2UFEx7SbnRMXOLDlrsXRuurOEVfBbQqSF
a1/ucHUHQi3uVULDceuQJqV2/g8HTEOiQPRt0zI/32+qYZK5RazmtctD6wiUyaWS
WA6vTPHPgPPLdy9Yiqk/QSSCgeTQ+6RfHfN4JY0BIRpmPkJwrEdHms2+GLLSGip0
lUIwRHE9UrHXfhrN0/JAoNerDdCBZqGQCLxPu0hj+jhcv6Yz/ax+n0X6zS0xQokY
IZnUSTMrqShMaLFsDEGHCZb0cO/3vVRNMKHBSjukkUONna1jHyVHyUcWx/XR8RzH
Tu9BwXhb4QVUgI7PFtI4mkuAeohcp7FCOAqPLdzw5AqFa9Ayd0PDKEaZwl28dXr5
MQQJKYQ36FKm+Vs6PxgQLWrYj80mWgjbgiX9MsgvCVOopiOn+1zQWp0/WKdKCxVk
26JwxAhmizVJwpyGgOpDbhP1bNyldd6Yo33HUlzWlIOhXD/yXrQtq+kC0lTOy53g
vWlU9X8JI0XEar7tDdq9kvqyoAA74c7QMbcyANvtl0AiuVJPGWoYbczcCtbuGYgg
qiEEUWaScSrE7H2s9frUgglF/Ex/ed0/KOf2iOutp3C37OyjLf0bellCltWQYkOg
oAtsMqa+J9+RA+kEj+3GApqe7KMl5bK5DkVMdPuGCo2Hgbguul8d8WKvgN4ctqPH
sCfApBoH3/qj40LXCyRtqHbXOREYq867iucOE+CmYI8sd0PXKIc9dGEjG0+MtrXO
MQr3jgaobQ9PPOEOC6pqUe0LC1I4x4geo4XJe5JXTs9z6nDSqXK9atbxak4b+NQo
czBmBzEVR+mM3XPQRVposxzUQM97/bTGxQr5c1WQ2TtjIYNM3SrZOnyiOY9flkC4
ev7WqvXzejdWg3EwWkGg1w==
`protect END_PROTECTED
