`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rSf1PRfQ78oam8sbAMTshAu8Y8vpg6PNXmMTCbZs8zXLHor7XX466Nsyd8927vw
zRquScUk5UFEEEAsDKzjqHjOVW/3DTZHC9ms77ivY6y/o76LbEumPmzWb46dVkQo
87yVX+IIDbwR8As0tWycdZfZj2XHM8jCoXZ29TsORa3tYFeglepz5MpXA9/NAzUU
Kvlkr2VikAWrzoy0l3+csbQwAZnQlBAgHQDhERWZQBgu8b2hy9UEgor+2O+ITgJ1
UL7EAkClwhiA27+fu8Etp8tNCrBYaUIowQs0YU28B8K7yZs6IfDZFvD96njOvpIG
a+FbFg31OaTHocvfSKJF7jp2GK12NHwgIi697mpCjYcGnf4opfH1MyuqInskssK2
dXaVANhF4KtZwsfTMCsHU98WbBCr36/3pu5vu2GwLzXlbnYeb0myW8fGNmBtCpc2
ehw/BNZe1uanH3u9M31u3M3SGsJ8NTypJbItPFuzVHT6yxI2ouN3hDER9qUTwM0u
`protect END_PROTECTED
