`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UvAKylPPPLwTQbKbg3U2TnPMqjF+OkQhOa5/UD+UJdoyXdBqMwRThVUvwJunK09P
0z4ZlfPU2tDBl9zdR4FckwkWGhouEMCHB1bsC8naNZxKcUiA7A6TGMxpmQj22VFY
BcPL+F14tEZyZ1HgeW4Vw9bU752j+DIkW21HBz5UkC84sRgzK/XXi2+T9WsJLN3p
gaD3eC1Riimc6tub+J4BEMQXNRl19p8rBolYH7ERPr0B1T8SJDYE5oatY84cT+x3
y3I3RQIl2ZTeQ2M+RKrylO5FwQCW2a4Y8ShQMCezE4vI3Ea2JOx3arH1zjWXu1db
Z5sb/eqtLEDk1uuIh16HpDKP9818RvRNAPKdOr9kabE2Nkf5oSwkDobdz98OSLXT
ksuFI25lUvUKTP49WN2vn18Hi+pGizd6gfWJjfGri4tRTYhD6W/QVs1X36/JDYfg
hfVR/0q050f+jSC0Jxg+DCww8dRNtnT8cdsa2fjA00aaamyvnakqMIUbbVgg2k7u
eJ3lqxULlaiIwwgOFxyz7HfOdtSf6HxNp02yej9K5DZJ+fVjy4ochr4RRe8uwsbp
r7Jcb83gLOuNd0RhpZnwaPvs9q621vi5NL3hRippZUWCRdOBsmiqo3ULOAWt3jWT
yEK7Iui9aBBMPvyywRWqK6GwvXgBfdWIKqlB84SdhNp2trQ+CgMg0pZ9pAECENQ4
YXbTRsp3YdHWTJNjmoztKr8V0pkJGaZLXeYWv8eeSyf6WsLroGS58vfeBq6sOsSQ
+i3zLBWSXxeadTEGsXV1sU0U3R+MDKxtQ1EBbVleFnuo+ZIpEEDAHLHyfR+7Itjm
f0VAiVBphVeRhsv7wV3KbjQbvtBXvhbR/1/+vw53kDfT3+dhUaHV2JN9mQegPONi
EM6yvnBVs+U4g4PzAOUJK/F2YtP46dUP2/qVCANTC1DXbiu5oCNoEFJItMktq9dF
/mplerNopFaPOhUaaLb6qKe6klgV22/RLXd878GQn9PWulGu7mjNr+0nYFIiH1rz
PQl1Q1Sxkhii51TGWb19WjtuGOI6egncHypBoHIQXYqVP0Ea7M555S/BxC2GWh88
GL8WTYqOG99fxEt1Vg9kKPeNneH3k9xbqyvNiNadNzPx0Nbjhu8mhIG1vx9rg06t
82MEh949nv1898RnrAE3BTsfZaomIOtI32HlgH55fPN21oThaJ5kE1w12VxY+vrE
s84fMYqeVIbGR8GLpzXB+JwpCb1l9/U6uTzGZ5M6XgM+V7RnsTQIAC5QMp9UOn8D
u+Lq3kmfeb+YY7V+rtyi/k7RnPHQwmPVNmRaEJIJWh+I0KXla5I05GZgsZMbuihz
TLQTzeBDnruD5ao93i2h+au2Eebo3IlMIuwf+dDAKCq8AQAuKCgnRnYxG0oRS9lG
b0cUSzhxLVU5tJo3FX2nV3fCpFfb1TzxL8PNxMzTHgSAV+wB+Te1hqcAQ1S70c0z
qI8N8umSwDSOsL8S9eza5yDkSnB58RpRPq2Md+qNn0ScbdsHPkDlQPUAjkS1yPG7
QIWHiqNcm+LvmDqw8L1VVttvhgh+TmBp81tC2t5jQFIVCvOPt4wyHopTueCyMJ2i
+AXbLDY4CR3KT8qLitbd1sv2otg2f/Olwlfn8bX70Wc/xbJ9TRTrLDKVyXWw/BF3
ciXXctNJSZ8TepmpWAgWwCtnknMaU1l5ZOneXkM6ve0foON4jd+OhrZxYo9SBKyS
3tOpJibV5akyKONo8niAQg1hD8BzF9MXmnGeMYKKJyvab93fOFhk2Np036LLVrhf
hOiF6qL7VW+tyDpl3pgIWpfDRQ3eld14yj4o3iEAWdXx5bJqGvXK+OE8sOKvM8ft
gLdbcV00/Q/GhXGA9HxweVqd9tUxZsM3htbrdfLw/fAZNBN6WqQzVcwKgO3c96+S
RacSAiOksc406+PJPbCzVjklXn8knaGGhH4obaNhXBdQj9TZ+AFtHr4XkJExDHnQ
LO4+6zy5BRAzQ3z3dsMaMj0POG6tgpDt4kNl4MKR4nGyE/wbV0gglTctmhyYVMY0
KQjCeDfOGU1gUm7pjrZpK+3lKAy3SaJkebNbLGUk+BKH5tQmzQ+YMewfN4gluHzs
fKbLTDsU55iZYlHdK09vo+bam36mhZMy2lfYUO3meQM8wVlpT/spRj1mRJo7ZKFz
tgX5ii1DUTSL1AEIbuL6/4orM/RcNu8//QF+QLkzpd7jJR6QaZ8byc7+CBOAVOEj
umwjx1ixxC/oK1950mhvaU+7ER2MbNFqglq8BSTuaW9g6DuBWZ4/JfUF/6DrlTdj
P6W0g88D2b+qWNGkkY5mfFkiq/CCTY+F+nLin4/mHmLJIJcDAhQEh/dMx0aLTd9w
csjSUhcrDz1kxPKFhoW8DOO6jWSnv87WXyqLQv6tkJj1b2EjF/yDJR2tZqm+JwJ1
9871tsecv48CcVZqFbkioZ6mb6x5sCH0GZjgRE6J+8bxRTvqinjJOtM+ObYStSzG
fgpSUMn2MGQKxWGUgCx64fH0E6kgKj6r92zRB10oOVU1BpEUP9t2o2DXMgdRcWmA
J528baEOToeu92Hm7+NpiPd1rIzqYym1LSaZM7mxr1RizBOAvmjmnSjVTUy+16bx
CSG8TBGm1mWv2CkmC9bC4A==
`protect END_PROTECTED
