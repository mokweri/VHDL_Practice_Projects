`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hNXX9R6pmloLqKXG109B+6rXBrQE5CYHgJzF5AsQ96cIYIb0iAXmlF0Js9WayaAp
VqtJJPUoQW9+dcdfGfP7arncfSwKF+shcCqREQuwpYDSagjB3A6Oh9wZvHft/gUy
C4RY28NeH6tEcsDKZ56BGQbLMyfmGG5QlxMNYJ7sfeuXOi8F3raAzO5sZMH6dJR2
u8b5+qw2MWdvLHI62smiKqdNZzVFwLvQBhqnqD0OisQv/mw+nPDvszByTmfErXf8
RZ7XJnGy+WcCA0HstztyUJagg4XNZB2l1wnTIMEFvEnluB8nmWECtXxaIxk2PJLP
/crZbbDFvdOPrDOgzlkpUIzDUoOImxbWqlClYsojHPWiQK4dVvYr/G2QTQPYpQcJ
OoWvXEUQzvgi2IpmR/V2oWM1WKg7A/b240UZC5SihOxOvPuRdlF9oSQxMNegElDm
znqUCLbMy/CFT8zAGM2N13OnanOmx1VkBFfV3FsmKlQ5mw9nZX6ZSQ1fderixPx9
cH6wsQHZ9q/aqQ60Uo0h3FljDEa/EUjfyEX/KUkJg+TLl33LFFYHwzGSRk/f3/Rp
JPyeMCAhvwE0+f0VVy/4ANCih7Hw4Mm8n+eIYzqxU9lXUOPbb/u7ygVTMa5YDEeD
v81sBokKAj8VhYZm+UFwe1q9nD1MW5QZxbGHyxoxr6YE8UyOch+TFJXXlQDzMh8z
CKzdnmSEDe8f2bScTZCzxWEB3m6Sy211nctFWf4ZfLa8UUtB/jGR10jzC/KHydRo
wG83Zkix4yfurNDZVMvocjNPEf/1GCSoyfsCNdDryk4dfiivRLGd7koVmDvRQQiN
vN1TcQx+nlg6rRmFhnChiu+lg3ioi2gWaYLXvbUCSweRUj/Fk8CCRSavbdoBDcHb
kDHV0WIeUCwEvTDXI/R9p8mq8i3FZhbzA5gt705LmkExtR1eNEPbH5vH5QpLvnxv
3zlk/GQJLAQCvOSa446Fxky2pnEj91k7nmgNRqigMWLL7po/1tws+mrBG8RTATo8
0QCt4/Tmagh0CPcUI3UGc3Gj73YS48+Gr4vm8MGImjsuAYHoFSQhg0muEN37cnsf
3qCBzedYe717+yq/XnXnxs/P5E3PCJRKPWHqr+ihC+IR3qDJ+4xEQ59cPoLUxCJV
712eLhIvlceHbJirQQDFuJEffqgVz0n8OAtsqqxzJyJlaSNlusQyteyEUmOo17Xf
JdhmeDbkamYBJLeOOTd7SXiQnZKYHgCxPNHu15EKvUad5N1HLYh5EmMNGITu1YRn
llsCgoFe2sRiC1DvaNh812G+hjCZYJveHGt57SSIuUk0YTcyCtk2yFLT3NlBi7Qf
AQmy+QWdff+y0fHh89uCZ/ZLumUVT3MFVMhIymFKUzGNtSmuc34Ws/UwKUOjVJ5n
G8fUuTxYzMdfbImAAB6F5rs8uSIleclJ6u1pyeFKaTBMZbdibbyoO6oydYnFld6f
iztKQgSKkkeut8cwBAvaXYSBEJCdi7noZ/BCMvAGHnnvqOJEVvrlOImGKAQE8Qbu
U26SycCHTDm0tZugJVK1GfYC95GTIyNa356aRSrYo4zdcmVM5Af41NIOIyLslxkK
A8+3ojMxHW/2EUE8u8hLm/QiaRs27w8i4wFktPGxGsfACFUKVbJeWC4caDEmIKBp
1eM43cNkC90TlpKZCJ6WjT+zR/AdKMOmHcEsS5Mnt9m/QIu8bUtGcumKALlFiZAb
LLIMrD46nQZhSp2oxtQulc11GaC4rhNRJvtLR6qn41rwYF3we0Tru24DVP+KYmhD
AkaikkGfBimtWcoi9PiNF5ff3v6tSuVVc2mCc5cgTbfaYebVXP3wj5E4epUdh+3E
m6lJa7TOuzBVkXBjD03y2ddyA+6fwgBEP6X3mqjHlz/6hnPGj6G0/9WfnUMocQ5w
c518DNMSkIJwCqpRPL1VXsjPsX//P6PAmc5tj9MupcR3kgxt1r5JlS398zG6TiYZ
3N81k7xVRJyAs82WynXL9KB8yAchDcLgGNVNm9FUUHOZRoXH2HT8lYFGs66VyoLM
fUaGCatZSjIUgCgCLAnp3f7uNkHi2WsbHNVarvA4eeJmOSWZDlV4aleLwHW7dKmH
o7yFlmORcU27J6c3YpwmrBhFbDjqvrKu84/GKIsOlQho00Eop8juX+2dYLqEUUDp
AF68vtlZnK7fN/7jakz682BCZ/SXkK/EcOpG0zCZpLuuhz76whXc0RC/DRdNEKZs
uuT6XUH3GIHiKZYsuaeFemA7tYhcPMUi5Gp7rUazjUtAatOAlWCc63RGkrisoGlI
diU7VAu5uEXfcF7FTfjo+ChCakvyLAA9692Sz9ddzPnqq1NGO0nlIBjn+ihVQpXD
W70iCEagdMrBczCnXe+wAJ11YIr9BIuCX7N/VcSg4Y4ZqCsuP+3sq2dfc5+LUJ7S
Tc5Tav+JQ8rqOAFocvMl85JUN+treK0XU5+kFGo4Cbk/zxrLT9zT8I+PXEdStViM
DVY1ulmJv0SBLtvboHJ1sI+XfLJhiv1kBUUnu3y8x0AYhNjMjvnDTqEQFEjDde/0
z/k9suj32VDiga9O3btlvWLdCAj/kMhZhkE0q4le30Mf04i9MVfohO4Qfx8Ha9ER
RBxeyMsUMuCcyHXxEFD000q7vlIKRCwi0cCYP3hP3ro/cTw6JOlfpdpn9YYbHbdK
AiViC1bQnJZq04TKrgrvmghEfvjEb6595rdcoHLR9Gn4Es52slfEZwbM2su5VVNj
cFhsMv9xjlrmkjSHLn4kHcsWgH1CnSIED2GJktiQcIMULmO7vyGXiaE5hHgPpV/L
k69qFEgLgO/gb1oLkK7IM6Kfse8DQT4PAnPmKEdETgRD841fEyT8cAWlRQ8KMlje
2+9341YDGo2i1c+8DjumwP1+znlNhyJJFZ2NBsuXwQ2tArneOq3HD6UprEWgVv5+
1lTdQN3zjfIvKOPYpfRObRJiEnWTzeVJID0J0k6P/Kd20vavfc89pyv+riFpqWPq
PHFwLcZlus+SWzESFt0eVQaOrwsIlzIg3ibwR0qqwLrSAYe5BWfB1HK0+IC73VpZ
z6CNgAI71i9QSX5CISSg31mCD7K6iQv3O40xwUsLqyy83qCJuk0VkKhfHJAx9WLU
SA25QXWCATwEO8GRQQ2V0t3HDawW9OkLZS6B6AnLGbH6iEh9Aj46gU7xQE7QQ1mm
jn6ecQvg92XPFaNrXBBt7GKp+OekPjFKXwMyKG16hx1NulbdkBIXfK9z7JGrS355
GCFymv5g6hvA8SGrnDtOgTMgh46dpNshbBKKZlU+2oZghlHcrOzO/wJTO7M/dXok
N716HMOqrz65bi9oYGCuhneHlMn5bK80uMdTZU75F8THhfik8jp5wPG9fFmWsIK2
yfv324V4H2jJNkRGwUlXxBwVa583X9jyvzHIZYaYvKUGo9VHTHb5IEDrUGhDV8RY
HOiPBYRs0tEZr6WoDK63diDxcSXUwfSun9Ap6HXGSDqvNBND1UeuodunI+ZcZLYO
FyTl6BgXkamYACcLXvf7FTcAgGev/C2KLJJnEuKoFi5zCjaTlhQxLKdFN3X81Axc
4xX3NqWVDclz8KLphBKmEB+cc1tTbbvRnN9hcgh1xmq87hITMt7acq1Ej++HUd+9
8/Vhom7fkyk/Iw3dV8YJpktQ30iYc6p+nmwtQg7AnvNlFlGxfssQs3ltxi8csaI/
w2WqBMmFu4ma3nbdcy+KJXSohc01aqLsBvIRe4R/Z2qaOZmMTFcjRoHAI4NXKt1f
WvbyyJMYu3bJYfRtg61w6RjG27y39Zxpr22OJhfYN2Yj2JKrTDzowjoq2rkwaazW
Ac7MJz1kjik63Fdf2xB2Hqk/0rwXE0OMbwN5m7B8SajvU3vXIv9LjK8MGd7ZK1Bf
5dQqzmfzLGnlQM5jC1ck+NmgD4OuwEk7Yz0YjJC6DnpQOYt9iG1UPzZD7P/FL0sx
VYkF4yiN7QSQLDHE5qAsHctqt+x9t5HyjyNzdxqmM/pQ9q/xG7iny/T3o+8THaul
u0MglDmjWR1I4wQrIp9sT2h3WDYJyLLN8j8jmg1SaJZ59ZDBd8EG3SDJu0HuCN4h
acsbsRf+t7Etg7VshU/+VVuhMFYZfcCuwP/wXNS/ur8KbyUzwyT/gDnPuH41Ehk+
PBfhz7o6KXi9IY9NXOJu6IZhtOXKRHwwa9ipULLWhwF0aWMxE5TJCR5ktif49mS6
NJhnPZBw3NKmbak/1IShQ6zDgMlyNgZ1B4/JNPhDzVrcPFkEKU80DwdrILQlUmAF
bmd/NAYBNxImy4/GMv/0WBh9ETEWkBgvpf50SGZqCzf0rATN26gAQukhk4NQdbfa
q85CPBjEqHbclc/vFLLq+AIjE/lwLLF9BVSGtS2rS4zfc+QwN9mNclrOEe6LcFsU
MLoib75el8RSUjwiVRecCiBasRLIK35CFP4h2s052dnIZa8Qt155HgtAN+tZkc5p
Dt87/IDQqMDKZBeH4m/M3qZ8l/UOG2ScGdViE+Zp0LbgIyaNSAmX9Ob+IkujHFDY
av8wSDNJxVWIUPyWtWMdiMlejVtzMzXA6kyK8DSIWU6QTJH2EKgQwxEAmeBnwwi0
K9ocJsueuAfkj/+Kdx1kkobrgj5Co4Q5ndDRRP3FH2BqENAtF4ixic8lMobTRIqQ
DIViICUDPf8Tq2np55/OXjeWmAMRC4q2gNXZ2RJ/v5eAOG+37IcuZFd0CtIIZ99/
8htrFt1HosMRvXqiYe23puIKvxh5xA/NS73kxb5r5gPsNeFVrw9bi1iOEVIPbkIP
TMCWVcWI46a92e4bkcIrDWLTfFdYqehgIAPHwI4IS2/lQ/OHSEoyyeLfxQc77Azz
IUn+eLuptSHm3yqKnc6RLP3e/KjiTbRJ8VOQ7LduUym0I/R3WmJ8IQEp6WBYymNJ
ghMsQEmKZctqZ1CP8N9HzpQ/0LXBSHEntxsMSctKbiL6fECDEbwl8sKsJO814p5p
eMNgOjqu77EzLNtC/9xVAX2m4Z8qbYyngPX0IFfwGWn5vbnKjk569pt7Ibsbcea+
bIODxNjbq3dCczWmiOJ3mOKO8jPcpjG7nJ2otnInbyYTOxCSblmS6meRcUkfq1A/
tHmu24gA4DrMGdeJLXIqzucC81eh2cm57649r1kQd44n028asNJwWDWCWG6T0UBZ
6uroCxtfVIAlyA1qgPPHZnKHAAMibXOE4+nt7q4DqjoJmY64EroXWHXO+/WDY5gc
EqkbZZxmKt4cIelVCYt/Fs9YKO8LLlzdW99ZTFF+gwYQ5vZAxrhfwwWjCZfntV8R
tvvEJaDG+lts/y/CZYnSUvBviogTh1nIzW5GPQKvL3OwjAjU/W68tb1i6aahZWse
DOLHWPx2/zPdQJ+YQ1+jFMbRS5L6Jzc+rZahIBSu/H1PVgr2SbWwfMFhMzvkkfBB
SlbAmERv9Y0D6BRO9FYyyZGWZxb0fq4wrQ0Lgfbte+nuZcUJ+xC0c5H6mH0ETXgP
kW902pXuk8H5E/dBMhEgBuUIBieSG44wIYmIc+jzYlrmwabJniptpOuz4K7GkKYt
J1q+N04qG4P1bx64d2dRN3wgRgP7K+YtVvGplrhbi4YvQS0tQXPNih3KGrMjVn+9
VoKomoUcVoazDDdOTgEXZkPjAqWZbWQIwcq5KMbkFSD1noZAlRl5mxLQHfHfFCsH
She6LFk1dvsxbeROMC1okW9XB11HCFQ8hk9Rv3LTyEvR+8M4CJT6gl2DbDfP8PmC
r1Lqfr2yTqnvUTAkgM3zDfMOk6bePjBVVWXA97WAByjtU//wVSkzo5bo8WR+Ichq
DPHj0SZSUMlECPLQFMoJtH1kdyVFlElxjL70Jnzj9x+5upjjAMzcex+4Mc/GYeFv
4JsocCGlBCSlJLmjBfTM1rOInx1o+aPbeh/JBZsycUgNuJqwHhLcYpBf0RhjFZ7D
X4M9UkVTouVJXRjWAlWJuKHbjrIryvRyd+oY6KYDw+iBaK34hwj41h0DJzZzoUPZ
4iuKJqp8CTDP9vHzMriNmPmbquk1Z0a77SNsHCYjmATCPhQq0x81/LkK9LrqUwjT
fAftiPUo8v61YIp4tqlUMEp53GklYUs7ekMkKxIL7lapxij9gifIk0X1K0h8UGsB
pHFWM6ETnwyaAwX2Wli/bWr980/PTJ7kLPSEvnb67l6xZD2l4OqCZ3FaNafyMQSL
apUm3QSr9jEoiy/6h2L1o7F/mVEZWJ+RGIsUO97jafS2PtyZJinEIWZgbWM8HHJF
7ttCUZwNMNy5BvZUoubNQmbncjJLObzm1tIpG8BSi2qnNkDbv2B86ZvyPXua3Vk3
gYUAIJYHXLBrqW7WBWhvEx9+w7u9iiaC3Iw0E9eTqCUPWklcwUejMxdTYT6E/p/W
UYX+fZx58A1XmJBZovhU3jpqvzTFTeuCn7+hYgLQROMBQY0yPAq1yKpkq+U5kp/8
zys9U3Q4eM2MW8WBHz4/660q05fcvWtaKd6qopUO8/DZCBECa3RDxGAu+0fEQ7yy
lCZnZ48CZrPrcP8aeYR1piSJPlg+g73uY4qHQXuxtNB44hDqPlnIWhIv3UC1aUHE
f4WQCTG4LFRUQAa/soAfiodu3lsZEmVWSz8lA+Rsnvw32hLCAg5m7DFSrkTcLC0r
N57E1njSnA4T0LkPVNPXU2gjOHgzWs9JqkBZ5B1cdefHDS5yfi8DxEv78tFYJcru
9d2RQBtlVmJyOB8YGOvqYNNmLL3e4H+bjezIQGwZqUKEHc7AlE6x6QhBTpVdwKeg
yrtl5G5elQF0ngV+e9cfotDU5a9vD9+dKExpAmnCPGaWG65NogORXJ+tgx4QVm+K
hU4XSTBlipdlFjj76wT2BNJlhlQNzvMVulFjOzw83DMM3TEnZWo+4/oOAMhPcmhH
TQ6eoTvxpcWE2WASU4bD+TvGqDJKkYL2u8mqZnxf7zIItNrUG8Y8FEt2buyezLiH
EsEZJTKfj1eA7HOZjsCvGx0UoQe6dZCMQQsHlBxOa3p8SYqG2tHp4EfwtKxP//vx
maVLRQWPmjSSLf/DDII4jiddNIkX3G0OipuWyNoPXsfi9X1XNpGSzLJQBvaah6t1
Ioa91xr3oExh/+2Z88tGUhE0cOAfL/+3ZNIyU6lzMLyajKftWhv1KJsNOXBzQlzJ
Sc/xky8JXbTFarJ4nVqD5YTTM7FGpjU02TDxt8rbUV0NXUxlKKgK6YTqdzRugTLL
piq1FkZ0PeIf1CxmFIfRYHfw/Ucoe5iW/VZa6zoe8ciEhY6nTJ9e7iICENXRbM4G
ooJWsoG2d2umiPRYjcpQaZuaU9f8eRLAOHYjKIk/AxOs5YYAlypTLtsT6g3tMscx
CeeU7IlGm8+9HbHHBvhpCBPutXDYCzdXxCiQWRIRQMDfeG1tIuB5bg1GkrsFBLGW
5rOr8mLJDBEJNDfGGbHysO9RLbcrhTAV/mSxTxaKUz4SZY0Pq7wgfaAKBgEzmLXQ
mL6f/+vdtp7Noa2/q/C4pzZwEEJF5GvoCEx75WhsQhGaDXciSGvR6r0Gn/S0uXM+
JhbgNzpUT/734FqjzKo0qF11m2olw13PlKdvpmOix1nviofrvNvq4DZPxj8cbFgl
Ctg/nr80uj1NXzFoQwEGnDBkZb/cOCT0qUFSLEjvABYEc11pu2K2fM5U4NMQcCfy
u6LN+JWVrmBeJt7VLnhCI0gQms8bKPLlrb1IDfDD8tO232+jfufqoNFTNj5UyLNm
mfK7kXKq3MtSQhpesXuLExSMeMIPMKWuDI7zA0Z8nTblmKjrNIZNTitc6633zGlt
1zYEvwMJ5E7eOwaZjRkEI3OLTv5NtSaIKH0eEuGrOQT8e2j/yfPzDIhv5I0c68sZ
Ymi/AtuOaIfSH/iDZ7wur16QrIqjkOgb1em1AA57+XZG9SRXX7F2dS9XB+oASS6P
Kv6kVWy0F0D8WZ27akpqlBYaM6+dMpqtivVCRXx4m95KgPQRtloCjt7aCsJRe6yl
DDR0WiDqGREfzrsCMywI5TQ0kGlbjT1g8s1Svjc7ScHxZfeeIvTsSIecQQVPKQq2
PiMJ5Tq/ceDf8sN6fyqwTARy5V7TeBfB2ogzDIyaW+RNQ+umrQYk30gceK0Ybo7H
w8Jhubb2PfGppdkmyCMISjuhjWhAhqe1Nwwrk0vRuaJ1WZuRVeqrBGXCJ2b+d2nL
sd4Srwg7+Jj+IagVCM6ZIqfh4Rkua4hPrVLyR8ENmN54TaLxVpDsebUv5jbHJBH+
aDPWqa6vcAECAosNsm+3OKZB+6vfGz/yUfGXJ/iDniM9xTVwbF20bA9vsuyIIRPy
paNLCSlwUtjU7vQSLu0LHMY8jPExRAkHd1VqKhQjpVtHRwfKj4FBKvfpYG37Qw/q
eYVJT3lLzBfFTM005soNWABP+TceEHzBjgM+XqF71wO1VgZRyNDNpfh5cYG3pPN8
VNPqsW3xm8157mHUQNoCYM1/wKkI+Eto1Vq//7CAtNCWewP1gG7LISvxqivFh2Bk
Ie4Cq1J5Txkm7v4wT79NdciFOAMaRLYLyzMKpb9+VJ6z+M6Aym5l+swIjlo50rZk
/HUNN06d+H8XVm4kQO41LtZXEUIIfl1mLGfL8fOCySmTiF0/n2TztIJ/85SzT0Fx
+uee8WvDdM0vnJgIjbwxEgT+W0hpqnUrlr3cTirUTzMfen3ObJJZrViEl+be9v9V
d3d51ZDeCNt/W2iivbZiA2X2C3CU3rarHhRYDkDjNDueAP650nQ74pC9HOlUCUJx
MtJU4G7d7BUvb6OKyEEhf8/YlyedAI3c7sh6p0pC3vP+a/VvTdsCJQ2eA5De4XSr
7LQNTbAn+B43faBOKtBQ2nGxGOrOvBsKy6ufuGMCBmF1w9fTRkgvd9j9s9/C70c4
9GdOcFyubJvF8wTtGQD5drnRaxCSdyTGCyXBR+SDpdRv9OhdVvPm0Okm93PMD2cL
ST9Ky38+Dt1BfWN21mfUuDpFhDstyDnhWzZT59AoKT8siMV6LDd/wHAkif7HtTR9
JvGrvmERZtk7Dm1D0sUMe38h4xGdCmSNgjOoGaiT/Kpj6YoO3j3X4WsV50CrYNcw
i3sBJnePDB6u9RzRHOQctphAH6p/3nTW9B7fje9HPoBe3UyNGEjg8PL3mJYZsngE
5L6yrm2mGgPRuTfEphSCOZU8MDMVv2ZJY8r5WYCKRYeFlJLDOEx5aNIWDYkmr486
WZUhNRJj4363bzMnlg2HPDESXkWuHT1Om1KJkPB2HWfTELz5ovVYp4areRBa58vU
xG6hQJ7RYVvxQq1N4IBvZsCRh9Gqjs7xYxmhW4rIi6+SZwvgUlzEzd0TVXCN9Oqu
mVs/yonVzHRmB7s2mtF+2/XeCxlYNtH+qM4uLgPuyySvcyMBkdvAWqDR4IBKDqUZ
AXPilESN0MfzlMF70rGsSi1+NkJCPXJ/dqtED/f1Z+4VAhhtR6cvwIPP5WsRNn0D
rgHeq6M1TjRgcrE4EV9rIkug6cNAcIJdag3q/nd/aumVI3dEYjgDXviWf7guO1Pe
sYmQFB1WKr4e113YTbchzC/y1FddW1EzErbkYV0YidPchGCiBBuZnU4uJDAo5tOR
7vtxICAReAWnWjEyCQCyJO0rTNWxYfPfzNDAfy88JOrdXrL90Qixqzxxs9Amffre
IoKOW7GZ7LYDnpMFNNVS9PO13xUsM/sg0cXgWANTUg7Wt05QkFYngujmy9h4YvJr
DBFj56QFLl2X5h20Mp/1QX3qsPef+tMLKyB4pKXF8t5Y2TCjAuqkNggkLgYN4E8P
2ibGNGjOVMnqcYH5r1PWILVYbkMCRp5i49SqUgFHyiSLvF+VwqvPs3/KU9cRYfph
Hs2ik++YNRPM/KWKpC/ICa32lKokIbO5cG+BB0eEG50XLoetn3MMYntsClR+bul5
fyY0mJB4nTSAjjSa/QLOOTNaFRKW69r9Q8xPv8IrYZmbzSywkjM3Vpvb/4anOw1R
CHunMurHLn3A2WICcRrtHn8ipSafMzzeM9JyTCzv/y3VCJ5KuMMXIvi3fPq486jX
uIpgBrr3Fs6iFW47zJuI4AeDMKsdjJaQwNgwKFVZskCQ+N1tQqPn3B+L9HUjAibZ
RejvkGpNiPzg24gCjWzko8qnmxMrBD89wfqG7HHSFT3SArvu4AOYDOizyKSwe+yO
ynyizhzxgRZWqR+eOA9fnYBoghUTZHYUPFHpI+skTebERcYU3OBVYP0RJZ7SHJB6
kR4JYpQCCZ9etZPfH8Q6nj6IBe/gHNonX8eHDRJpT+u26QOQnxSFhulrdBsAMcHu
x12sjtLpD75pKziNuovBKYBg33b0SKRnVdP24zPT2VUbVGR5HqmbarTn4iXRsuz+
tqHzaW0BJqHiXP3IW9Tvh30CnxrPsFaAyXVxvfxLMD4J+488Do+XjK2JI8LpUcYp
ASbpN9n2FYTYWiPTBp/DhUavuyifwqzN/2LU3zRvUXtWcRQ7ciFiUHiY+GXbEXmK
m6+F/U2PkV5gVH0/q4HFBr2NtdQ5hnvK1KMcwlcE2bnTo5bbJ4qGPfywlBXCyuz6
8EuHorG8Rz5lsyPNKDkyAGSkpEorFFbQwl3ppB02dA7019UmSTaJ6rn6dKCD+5IH
zNJ7MJEtvYu3TqyWwYicThTmYW4ANtOIgIkQ57xvXj5qF9toGnSm8ftrImxol3zN
a4InCfyYHBbcEzIjukkmHryr+SVZ4PpsVZQDud0xK14brohS3bcKduopnEaQS2r9
/pyqj0fob8+Hnin0Xx87+NqyHYCNag7e8usuZKsmtutU0L4j7JsLDFQXsoeVNGnE
ngMzpl+SOQfbmVKI6YoLrCjQUaUhMoGtRieDEykXIGJWMqjNx2bp0jG/W5lT3EPc
1mai1B8Rlw3HfIcPpbOPNl4XbDdsstKlB1ebvEf/pGlzDf6Ez/t0QBxyBcKHw5Dn
MkO2iREq/MYTUKQ+vOkBRqi12Y6fk/VTvHOvF0bcpk1w0G4BrRXWbKqrGbVOcmDz
1W9EX8DAttkTwGG1Hrj9W7ipmXT0Dh9sKas3FGFf2zscjtYaV3CooF3Ej6DkvoUo
sX/3eYg957t9Y2oX2Ufrmu0br5qEAWTPa2qd8dI4hrUD/vf85XJQoJ1Lr/BbvXdP
PUG0tQNT//4Cb8rk+HMUEU6rI+OgN8tlrT2itWcqNbTa5qTiyLB0+rDkVj/etgn4
PErYFPsdApyyQTcmKzBYWzy8C7p6GXzjGCdB+cFmlISskC475XTnJ4SLpzP1HIW1
pbLARVDaMSO3Msh6qJlXtom76xTH0+PigTO4QXrymGvNNY5x9yTFCTmuwcnPzrhL
soP3yK+Fns3z2kAu4ay0Uv6vj4dmP6ZCzH+x8iJ7FDxC4bmT8V0Ky8P1MffRMVkg
PJQ4rrOapv4NwLzM9GQ4DKUBlznKMRCT7XcDJfbGeKSmjAkMPtNMkVk6mm3p1IsG
ZGMmuaGW/OagSb8muFgA5gBhdJ/Rx7vvmFercB+zrQryeMMDZPMbOJprzJ0cE8lS
WvNbUYkH8ZzJ2fjkUxAR2pG3WVubvoecRx0Z3c2ZLTISxnCXIzdIB47Ig80GMA/T
FjZZVuCOjbayPsBxUFhqRjgeV+7ES8h0ujJuGGAd/GgQWtqWuVIeArpTPo1Sdl1M
pjsmV+2mm+z4HvASSCVIuqMBHuTFzgC4wpYKP8PJhZEhdC76wM4NqvjE+B6kZU8Z
g5yR66gXGjLNqtTCQoZSiEn9w/RJW0XUhs1X7nawW+ZjgND3h8Cs8OVVJqF+++kL
L98EKCutJIMhbUF+qzDLBwAnbg1AUIX7GWZJfu2NpEpfKu8ckODMc17bHQJBNEeU
0UQj1veB+fZKuGiRoT79JKHqhLB7EdNBR+H/oOBE6X8ZZRcWoLKvjqYk3j0I+KMM
+4OiKTiNsBCSBnIWvmQCj9dERECuPWa97agv4fyCsh2kOxXYI0SC9Es/l85wPmwu
Uv1OtEVhYl8G7mak7WEJrm9MrkJ5IhPMbnIQHQ6SNTxHNTtj/+YOmsG5wFd5WKEL
gpVjCzB60GSFzLRXonBFvoEInko9QFaCev14DjLn33OEewI6dh1Sg71OyhXJaWzn
OCdbx5r4L1NX2PkdFt3REIu5jkwbKX2SMADYWMPIqNkwVrKomjml29JrTT/B+ndU
5nNYEdHM7uOioOmdtKC4B/t0o1A/gOljZDl4E0nhp43fgIZywSaX4JYCDcZlu2bz
ytm/zMQBNl+9/dQ0VwVdC+b2x42q6lrbg/DPnCnZwbAZr6h7GLOIVHQDQBuqcX7a
nnRf5cw1zOpr+O7Ie97J7B513jyN1TUhOMS1RQJzSuzVKf1TUbZub+ka/QuLXRkT
6uJFMLX0Rl16DyHilMzW0wcfFqIS+P5AHRnbjgFqGahZD+ltoqaKJfnCaPaTR6AD
h6ftajU/kHaL5X91STCCJd8ZAMUCkK1mO3UHBBb8eKbopP07YWmxTIHMCQNLhQPn
ICnwZYufNx21Z0RvbV1xRfDF1kZhMAwrpbfjzoMQwqvT7B1uZ8EmOsCxmug2vXex
EOWf0AYjuQL87ZcMNKW/AxEjDkeZmcvzV51QnVL2Xrq2leebwm/ELUlCiy2ZBsp4
W/6Zia/eyuJZ38cTstxK/eJ4HfSjiYvgxgI7Bi0C5xknpTmQWeDWoquUakXay0IY
fmObwmQfVsybBD88E7K6FYIN79jTNnM0DgYRU6VoHLONO0UGw3ndMIlkvPUeLwPA
LVNjRTY+JZe9cqZ2GEJTgLMi0njs3f2PCR6Nod8wZPrgnw7OsiKFh5vw5nSY2B4X
O1V31XRwCwfbDWXNXMjmPBq8JuULjvH+pZzOPG7QMuBBasn/knOgkvbBmPmHJiU8
/H8f6D1DQ77Z/urPCYrptkWnT9HYiiFS8dMu0riMRkfgFaU9sJm+83NFX1avTkHZ
yodsK8eB4D9jXnzhGqVkmuqA03UtROMRA1JIsMuICymh03CA2MaykxJdurt9AKc7
b+GmWhvB6olvh7oCxhBtRyWoecxr/hqFZteSvQfx2bBYcT01kgzsP7Fg1rDRhfEK
GSGW3CMlbC699zN5CN0V3CgIpF7a62xkgQOHQBTWfIiNSbz7qjperT5ZTZzl60TQ
ZavXpi7snrnz77g6d9tBT8Z2D100sZQ4HC1FSJEcQHaUwUHXYpH1ZotASYNAg1vH
rTDb+PvqD81smklMenmHl/WJLzwdaUwtJvtEeRmXIzvOJ5d2dtw5MnEiaCzD3K21
28Twh8f8ak1WSKV27B5KWCHvB/u9UrNr/zJYFITRf+jM3LJtvgBsyErr0mZLg5Ia
WhDVjetIQ04h3Z3hySXqMLQd4KL+Pga2AcMyAA45N0GrqrVLRpRuGHrbrwF/w8vZ
vQumv2oJom+OqfccAZK/Zuu1XB9hXT1q8iTJKwLbl132a05SdqTPjnfNwnKy3Ayc
nikJuIGZz8zpYF8fgiVmq1c+lgnaTk0imcl/rZs28LBVeWT+6gN3qPy9jwHot/Nd
wZFqElHaL9MSV/7OT384MTtUaCsS+IdIJYW1lfCjo+MWH+P0Wme6cVJWXRBUjSCg
igES4Qgpw5ArtJxn3XGPLJ0cax2jQ1a+tmVBYlRWblKFnKOzzXcOh75hgJgdA812
ZuyIUkq72g4EH7/puUzjcWiiXOBztQVTzelPZnupAoBnk/zZWIzGCHtNVmRyTMDE
qrkF0YuGEVCA7HTEtXErwJsmAIhNlkCvBDan6UHUso9+NqapRQ5RN8ottRMBZvsx
nKVZqkFUip66xClKrQA9gpltPRFy82dJq0+fofiweScX2ZEHrH+ARLndzTx4u31d
AXX30Dooou+IyzpQnxd3FYmyQD4r90aXT3pfcbmUcsdS6afVoj3faOIsVVIJwOkJ
mFVYHtFMJGxs+/H1L0XDCCrtrSvPKfO7IDJnefv5KVKNIH6saMZxqluHDwoytkAo
x2IyZF9Ha0r8KAVbiiG1oIBNHpM91fGVeweKHJu1nEvuor+3TB5hLAH+0cdlfCdi
0xhmllwAKwvS232z8EY4bjLYvewHBvrOxSi+Y47+zOBX+h9Lb4/zmzwLRMA1mnrm
q3wBT/C7WdsQ81/4CZNt/qQU/4X1cHcJQBMF2cHp0o1sLH88u0Jjh6C+wO2bIkxa
BmregOmliEdd6FAn8hD49nrsoaucij35X8gheYKnsz2STg8neRUVjxgyKslmMmE3
8JMMyfnMwXzab69PI+3ClC7MXIWz98foA513lmkAb0U2oK6+2ezXVaygYWh4/xAQ
dgwGZFBcLBe1Accw+feLs102iITI2oe3VFqFb6qwmRbzVTrUj6Vkay7/VLaYVFdT
ArbQqWP0Scw+X318Db0pOE+JWvr+Trv96yU6B90SjpHGnObs0rOq7exPEwZ/eZTZ
dJyXpmVkksjnzb8cw86Km/VtpIBqu4aFE4RI/qiPkl7uqoVa/X8wC+mNsJdd7vZ+
GypagTHqDCPjuJ8coOYoEluc9UhQzMD0nloDB6H+rMo/oU+bAdsPFFuc8sa5MPbr
xLL6DAsb9dNhwWsYkz2j3f26MSStbFWL9dDohSQG9jIvOc0sG43OhmEt+l4Sn6YZ
BHjFRpEdUQtyBGGuYpxQw62X1Md3ma0lwpPm7NVxp40rO8DACVIcR6FNGSigcG7L
G7n+32P1nFxSNehqCf0+Ptl5OLkU6nK/RA42AkK6jIC+VBkSAB/kjpfHGvF2SZde
UpJDhLRxkyhavw0Yosa8YPuWjy8bQH2lXinFfwWY5wTG+lD9b1w4e6eKGGO5HidM
S+fbcpFsvf7lqBnjANHCsKfmfm/UyMH9FClxX2ZkIDLJuPxFU/lE4NxSHtP7jlcK
hQkvEIC/HQs8vZBpV/J7HVbp3oxLf5MtDHuIKDKvb0z5AMJg9EBuxzbR2rz6Vhjw
/WPX32+txqNZHzoMhVdPdDhyhoJYDV9bwAJwX6xyMHHHydXflrPnZBzAEcy+x1aH
JbXWGiNWOkc/8nN2arOv5AmtpiXU9Z1bqZQOS17qyPBq6k9n7SuwiIj+DBG4tkyd
IdC9PJfDnP6TnGk5xodpM6aHPJ+crfvb45QPX2+io5XfnjRPQZw2rpMX2N9Ip8Z9
LwgZpFh9eHJX5hePjN2cmD7sslcRMsEIWbTMF5i4raGvNeL8jIYSn7DMr0VEl1Gb
rrkg4QjIUaYq5nokWBQRWwljDDgbaLwBosBK8Fk+vQljnQubYSDwjrpzTyxbd8EG
lW0fot1DKWDmMslhesO9L648sIDiIXRWQjKE/A0ZZz9JbMNQlDySSUTGfad56Yox
wzI7MPvfouGXf+G1I+/qU91rrHynS8Hnxw4Qgcxu55T7EBbnVJPSQDz9abbQOjPd
cVxTVUINZOW1s2JNwe/qUuv/7AFxO3uA5WuPH6GxWiYknDkq6qXXvuWBFzGuIEZ+
pGcx/iU/Uwxl7qoedWQaLGID3KYX8uAT9BwL8vLoCE5rJJlEcKUranBWlOzXedLI
otwsG7VnKBHhCgTfo2d29y/ACr2jh3v1cBOac3rgWFkB0IODy1lD0aPlpSSPZ0Wk
L9VQUMoeWLDt7vDzlucFsb08mMuBuKjh0kpn2gpXTSqknOS7R0SDeOoMKeHrha6c
cN+IGkWe6uZNiSxXi+S2tmNGLNMbAMEl706PQrGixuOeyGEenJ9nTM1H9Q7cd+9Z
Dg0oHhhfdsO+kp5GNFWZQ7sQF98qg40AGJfFLNuMjOaSiG0dvBrXtzlcEeiV3/hi
+PLWgIdeZ2njFKQ+oJdqNTvQFJ0SRr/jzO/Rc24wOQiBxERqCsu1hepAYz1FS/cH
PF7LxzKRwMPTUhjE+CsEARhDr9b0mpn7uAukejWzjV4uxgvR1qg2gGiGmmFucVqa
Nt+6Va4rtwFSM2EecBJGztX4nCEGTHa8yjaxV5gSeog0VBs+/ei+8fxEWspV3BXP
z6SBvavvlEFoNEmSbQ3MacmMVcoaxKs5UpxsZUqP31QBipdJ3K2oERhi5CdXwLig
E4woz+c2kevOdZkbMB/tqdIx23zESXLbsynttwSovzJ09m1IvZd6Q9ZxTyYJizDQ
KsU8R7GHfftvC71QEPejwLUpXWtBF/sNjjFj69uVEPm0PAbqIfGlX2nAJ8qjNjQs
92uoRHz/2c0ociKLN7D1eGJgTZVJgD5APnmxrCDQYfi3P28DwEclY+royqSeZtFj
54pqsuipZva5DieGPB0SzZQolEgFYi7yIKBl0LAlcMGLeAV46FBTv8u3dHtgDhPZ
G5izs9L6nJjRp+eCfcImVCHxTiQ8oOGGwpwEN8Op2HZMK7o2ECsJSZX2DzklJHnC
0cUf6y4oDY3NN8feNps/tSBGaKM4ASWTdwUtH+mpJxaplrIP/kOCw50odEEJ9Wcj
Z7HCLvm2XqVcuHtOT9haHtn94VwsoI9qXVEQjk7M6my51fJc6RyYB9tFm6WqSY42
lw7P8NEURTYYETRPUvzVAnI4U796+IH5dFE+wfNTlGtQ7uvM5iDz2i/txasSdTrJ
R+5aRHfDJ860xGOnXQZJnEIXjQMZduroVKCcpDQudi78uHm7IhsFN5Er38fo3ULO
kMuuTNCNSdI+E51Xbut3rFbtgIEc6KBD4KIx3V+DVAHifudBOIln/bxfX3+gibHa
C6dqDNqrc1XtIr8Zr5VASvAUDHgCtxZAz1Dliw+E9koTZLRXkDK6QIl53Tqr2HoH
td6xh31B7G3SqejOPbpjf/FOZ0Z0iQ4UsDnU+r3A3fKqBNB6mQssamaaoakHAAm5
ZoPBGVsyFpUAtAuaSQPxv5UvfVT+SzJmnZZnhhfxLT3FbYAg6ngwAdCNBt0RA797
5w1DEWNEAeb/VSlugJPtUZBHzifbAPZW544ltRipZ0F0DuniAkXPyKOwYVdb5R/m
P8zQVfskmyRdSFmlfKvNCdB3Q1e3R6JLGPk+XzbyhCMY2UDQ+m+ElaQGmKYnZNAS
q/GNp1GU0qrfBVKyOHidXw5e6LnfJwo/juEJQedqpbCMK3KUtp0e9tZ97sXqkT7X
Ujym5cmDd25wEs+ZQxUl7cb6/RGV4rRFCPRigsfKapgAywgyyyQnyjhK1BSSuks1
VP5OYMAKuz45ySRMqbTaS1QsLT5bWdBdIMKFm7uPWnchlq2mv6kpQDHlO4xmLZLT
Ne1FDAuqzgkqHe2gD/WvxaEnYIe0F/j+DMB+2TtFpD8PJZeprZpPgwPSy8VfyHPj
ZaU2nwGImjszd+tZjuxX4II1L/6H4QO86uVyxDpdzduqrmWT87Y2eA8Q3BjH6F92
HPW101ciXs5A4NavhUdbaUpxT/qG84EH3d7mtCeMddfnIkaQYw6/O8Nxpl+MH8AQ
T79QP5idd4M4e/1QOnvEVXzCSaSXIW23px4ybVPkeucJMvUc1ewkXNcFp88WXz2e
T59MufXeCzHBz1ht4fprztUh7hhi/c+w34bPidX/Ph38BIln9ElACUaVN5tgAg5o
19mYeK8mTf8e/9LemxH79TpR5dTNqhl03BTqFZpe+JdQQB1qUQZFjiRjDrNW+Idb
wCqiybFuGezdwzi1oDX19YLCW1jhb1EVw3H6P0s02mb/Zh9PXM0FyypBoNU9piaL
9gNONy0Novitggdy8akqpFIDF1lHu90o+PE6Uo2j69Ltq8HU2MWeTXutW5hoTTpn
+jLpqj8VKsmFEfG5lJ7Wx+Rl+6Rve/pV5bYZ/SVmONTpwqJZrNSszA4lIv+H3P64
Ddba4ErgkJWTwWBOvvDscgAmQ0D5HmUxwsL0U80be2NLlBULPMt0FDdGGAL01dbi
fr66m3e5u5dUZGcRDWISmKEJ6xiwnyY5a6i9a6dUJi4edUpnaXtkPk8OXwCAUe6f
YPbA//tMtFL8PvTLzkwoV9C2rVZ5ZEFTZo3nZqHfX89W7GlnFzftLnNpKMGo6RPC
7GiH8GZasfR3nCCCu0QHXsK2Ec4DlFi9sDKTqJO+yWqVcnjBR2UWrFQswyqgqu98
e+KTuBZJXH/3pp1KIOgYZcZMw+0k7172/JDpga9XPS6uK/gHxj+omqM4qCRUp2m4
jGNGvzZfZZWw4XNcljIglIHG4PDbEUrEl8z/mL8DocWWlKjcygr3KLIbpKpOQU+W
GursAjXdWzFCHxr9pTUsUC4bYfYdUskzZ+ruy1dk8EWU5sXlhIC/lXsBp+saW5xb
Y8Pdfw3ycb7dGYr95h4uBxdNwhv4Dc6t1Xm2YQQJ+j4v3O0KMxivEboXn/PorePG
/5t+8ECx+STRf0neK+glT8oET6Ebti8ylVqbve+GNQYnuLlojGvWoo0LiaLXXh+j
RQ9XiGtOAQQ2z23gVrMBmVSnYe333gK3XD4f9J+B0psMpVmM/6c2+SX4gKI/nh+w
Jk9yAO5rnImlaC4yJJ439S59AOmFeLRu9nHOjQeSXTE2nM08lOOBVJc13VZBSmYw
p5FSWU8LVFKMkPohjBCt6bwB+JVIlyakM3rZBRdHkvLKua9X1mxN2jhKBtgZTIwt
/1SAxLIVrbtKHukv9HdwNtr4L6bYNFrVz6Ho98+cWbxe2lDCSlCj7TNm1rL3jxL5
/Ucl1lhbpsS53Kz4w6LKhq/o9geMXNNMClHpdR5ox5FSw7CgpWR0A2BcqOlElN8Z
ycJ5nkIlE/cejz/XokHJjZTHLNJw9/7+JZRDdZ4v+asygrZBL5hN4Bhn8bibt42O
VHZNXzWee70gIUz/9rTgt5SdX3vq6ptoMcdT3KBy2yat76RqefISr0hihp8yRQh2
ribunYcfXNRHv6bVvQkI56NAbUozmYBMASQTMwuAZVZ+5Pp/fMvRcjQnB4uphM2S
pm3IyyHNGIKfBAfODBe9zF+KW6wWz+YsQPhKAFINn5QP6GREb5P5F/lDHXHaxmUM
I6V5irHWBdIO7grxxHlalLcB5ytjVde99m3G43jz+gV8whcIKyKSawKFw0sZGksO
SWpegquDwrYZGzUp6LmWANlviZN7OJI6PhRh19xz9coNORwp4QM414obsL1YmqdH
cUNfmoV3DnITwKhsfBs1kIzOMAyw1Lg3LCnJdwBHbj9UyjbRH7/ykuf0sPj5ue/Y
7Mpu3aGsJT0TxbjF+lpIgrLWq/I3FuRv4OZlff4SEVrdVYWN01rkC9S53unIkFJR
70Gjhhq1/h0o5ajFLzVsq0aknv//ifn5G1sv6yee7OrPs4RBMHYp9ThLSNeUKu8G
LOpuKeRWpXUZV8INKZkHRGiRELkP/TpI39wigLfeSy0C2DCU7m3Fs/HS0t2/fmqz
GetpakujhOUIQ7V0knrajZpoDgvToXRzAVj261gx58Gf+IVBm7D3+qEqgVN3zRbg
NNoROFeJHtmoDhTPZhEr9lfTjzgTjk+lUcog8Cmo2+LJo6dR6i/mvBG4X/0/L38d
zMDO/lxTNiWWg8pOZ8/Yj5KshJJ1DLnpNSoLqXbsGbo0l8H3uGaXM2D/rDPD9VmZ
rSsbPlQyMna1eHXhPSwvsDhzBnglDMptD21HqxZbagf1+Uab/ZEcr03ZM9JVaG8p
65JGUBZDgRknCCdpsyzyB7QfNv9NWRi3SEUlEm7g7bYoxe1iCIqZM+ZVt5wbk/Uo
tObL73eRfuIM+VX8ubtyLpsbUD5n44aO9PAk3L21N0KVP5hPox8lq0+3xY3+19z8
cawTutTqQX6bNG1tRGfYx2L8PRvj8uU3XQcp+sGBMXSz9J9/dYaULoFOXTXBUsR+
V83irxHEcOLlZzjIVy6MMSsAENvaeQ8GGFSJ7B70FA+yG8wREOv5b9M+u34lz5XS
V+2Q+bXjr9OEPcN7HDzMBVd+82AbUJxGXgEp8pHt/FvW3/uuNwvAiaUaAB/k3HHS
kIVkJkkhOfXbDsPkWp5Hzl0alPbX71VJl/LG5zxCAH/EY+QdRyQNJSke9CbblXaU
IamlDJw1KHd6QoBFAXUBTYDtogW0nbUWeUTQ5y4opPizYNvCyeI2docHSeELuZyz
RyO2cv4oRCqjEpr/ccdxZ+MJb4/oOzoue2UKaK7L9bzhbBIAyZ6UIf6TPBINf5Cm
7TYllrIWfyllDE7ZXii1C6vdpn//BBdnd2XaCh42sRugaRhVyMBA06CTUhCeVQd2
i48hmv21AexCzjASbRvSybU6mbifWZW8RrdfyLzNvnYdfRpI39Kh+lNSgnJhjhHY
oaAWvmhGRSbgtjHhsOkTfCCsVWQETaTS7xjHxtcLS328ABIzhZ4xQsD6/31T5EJt
OjO9hPYq5loFq7/F7eaqIF+3x46Q6/MElQ6CdwdG/qH/ndP6ZiPm59eBXWvqnVIQ
J6kFbH9sWw3KXp2WdJNgVfpLVI9BAD8BzeXn8876IwuNNeLr5Gr1sfyflV7amyA4
qmQeelzA1sVFBIggiO25KTbWbasm1VYQ013r2ZU+CxSbZkogkTH++KYVy6qz0eUP
fnPFMS4A/SYgak4atQt+fWT+90YhjDGlL+hV4ucj7DezwzOOItkPTJVV7g6HA64C
zjEWNMDEs0YFImz2Q1YJT120fgPaXNYeKMnidJi4mWKQxyWhhcv4O+31sZ2jHFxa
ug6r7Qlu+bcuWNOPnzmXNF7zwdEuw9rfuy5HVN0XXYwVMYfdQXiDv9imrvXIT6Sb
ayx/1F5rcUUSrQHaFhrZ0tr3wr4r7ydJAXX2KgIpqLoecp3u2dydgCMHVJUz7stw
fhTUH05x1L0cRko7NF3lLncPsNQZ+Dv2eo4Ran9Scm4eVomb4oH3UUYLUkWbY5SR
QZ0CvaV7k3JT+idOMrMHvtqNPDh/BaLyaPYGCflB887uTR8yDgsZt7R36SpBlRtZ
DFeiKJyiQi5muXxNGErYEqs9oCAYiwg/wZ0xhbSLNWIc5oiyPYOG8+1uBFwe0bNV
7zJvzERhXEgHt8293nap+F1wN1X9gjnIs7+oooh/hfJq2IPgRS+7gJbr5rjGtDHG
P7WIjtHzLNnN/d5pNoKxAFGvIjW69wlar4gcgIwveN27k27GWwcrutIdVTj/6PKx
iRszJ/I0NTPaBfSE+6OfrnOaKBXKM0KPm1SrdbUhIBxzAd5Men4offp937R5xK0a
s2V/Kd3tdvL8/wVCmd6xHtuns0LIbUVH7in7jJx0cro/VP5bM6VLId+0y56EW0Ft
SzGGF6BBtQDdOL2fc5cYSEfVA0jpWOdeJZp4WUcv7RftF/P7oDJJ6E5OxzvP5zGo
iOKnXi5VzvXThF0K0OH0YE7O5hSDSkSR94GHRklUMf3TvzrMp8yfChXccttGzAq1
mSrzIuExup6apjqPqmgFFDEXLp/fNHn0a6cP0dGTOav4UN4POrtAi/9XdlEslKD6
nHbMJDk3GOZdqmtg033O4qBXtYSJKe1Co3w48rJLhPmLRMkztHnZCABnlPAfU2nA
zPHuq+X9i20ceoKwWKCjXNZ19FfZ6azF23l7ARm+bZ/5/3UzRSY9eWna8zyPs936
uGBhoDC+uPgAaMg3gvvxYBM++nYGq2pSyRkDAsyuo7uSR2BBviSqoLnghrfmJQjX
Hq9gZPKyCctgNldlVNUwyo1Brb3A+QWZftpxOJ64NAgkExVtDHUGDn94lkYWxG7B
V4eVWEHTX4ek1L3KlSWUc0wOA87pHTU88ex6zd0pELW1k4brrXZj5OwtuMZvTWH3
4vFOIz4By9h0FPVVnvp8tVnjBQLSJvA07M7D9hVFPQAqRrIEWqc0lvFFlsvvDzCS
/cnkafjykFHZqyPfXWeHU4ZDTcLeLOQ2+La86TobHJbq04kEWX/RPdtXgdNxUIpG
EzPS1gWLMVJcPK6sl2c3Lo1rMMyqfQC80j53DhJS3VkD6gVwkNsgmf2th8IvePZc
cWIllr7qHnCShg0zt/eF/SFlYjfndk4UewNBXDB/njVeEwbmk54z/vPtZ6mT24u/
i3rCmfoXzJVeWrIo1HY5w1wkOC8SVeBBOH+A5GP+OuLx/wo3YuETQlx7OqbK9p6c
5wIm9Qj6oIvcwBV15pNIBT5LcCpPaVERGhVtaCzcNgOlgcYJk/z4UJiZo/iCDjDI
iPd+GtkQgmYNmlctNx1fb0DkiIexnmb0wDaHBg8aWY1bgx9XzvZlH3V/wU6dVDEV
3EYdsowSM5UAY77FFF+SJcgd3zA7ij+sdd/VQrVAkdKytzruFsEqlKSQe3075YMU
1OyrAnGYdTlvp7ha5MSC5AERqlDNoBtCAD+23tU0Jq6yFZsLNn+kBP6BOaKT8Lpk
dcLo2OBnLeUCiDlZak/eidfhyIRwurGXID9uqDxT2wFtO0PasQhtvLvfj+t1ReAX
wbNaZyt7mBkBAWDtm/1xShTGToMAp6JJqh/SmUbQr5f1PjfY0n8jLUyuw4OWRmho
mO6Z3wcTruZ4W5GNz2745JEDWc4HXUTrnNYnKpT8dlTp+PsSHW3Dhqzl2XLWwy/2
OmnMwAjb9AigxKveYQ5V9JuYVAfXDkHP3QOOP8Yx4SecZcFASTLBniHgANQlk9J8
JxFs0ElXNKps6Cee2x11ZH5YW1HqfZMuEdO3aaTp1mzDRZTNFSZD/cMdBgClJSa8
eU1wkp+o2EfHIAaWviV8EpqW3/KXoaJTO0AXoDmNgWT7voU/fgi/Aywcal2KIj/U
9VJ3ZEPfK5sLAxxCbySVWSMd6EWaNxHeBtHAIx6SasLUHu2XwGB1z86QmUvfJnUU
TbSw1zsxuY+BFdEubiW+YEovQ8boQwQjxU4ES3LMzME1zsw8K/SaaSe2PG9/QPcB
onrUjxO/3iXpwvQyBVnPA0KjQsnQZN3w7KwH0uMgRUooaVc9RLhSQkGj6vmltRnh
gmsiEMdSq8na2o/YvWF5tSGmoZn8std9FKazhe9VfoNop+FzQyBTTSn62/WAgUlT
BUMR5cOFXsScRRlxBqQSiMv9cSK5BATRPajtF4Rm1i5aE2kOZNq/SuBVvTj29k3S
MJDBPc+p8/FClUwCNOtkXvqS9B7vo23I6oV04yHM5DIbf5ZGD3flF9Rnj/O2V8g7
sGefa5HpPw4AImoQeU9REZ8Y43iTn7jnpkaGkS4zBPONtMA+0yLOXGpqi3Qt6g8r
wWSP3ClPdOHhXiO7nL9dFLSSpgoi1z/VXat8/H0oWqYeXigdcHBWcWjwhfFQBtRN
/2stm7wG2DYYd5XWa0I8X2+dUGO10cTngo7s+3GjgvY4qIUhkzRHxO6pIdD2pjqC
CZ+NOlDr8UjhxyU8izxjX9bFFXjEnwM9h9qfLYEOlWqZHOIlgdznCVSwuG4gVXyi
y8k/PAdRPLFlc37ZinMzJzehDmpZQJt4/HGvEWBkWm/cmaPpvZwKZFjUZ98eTLGL
XhfJyRp7OEhILcUeTLmTCkF4vAKWysGVDYV1I6/GGWtY6m+wU92HJVfMKTrnj+5T
FV9WCNG8fOwKbaxB2zY2+Gh55lDvKgeOdvOWIL5a0TN9ocKIgEU7u43ZfRhGsr7q
e+NU1QpXYfni8Bk6RrJyefN90Ju4bB+dqYXWRs0RBhZ0NS/MzCd6vT9N1qIkFY/x
aUiIs9S8U7iaJqQEVyBv+iMp29UG4oUW4BoPmKGW4jUauTzPEdVosGmEKidpaJ7q
RSytFSBBXNqRuBXVjTp7EXh1u9LmoY7L5GsY0hVBhKV/roIbdjnxB5UqGcfpKkG4
OBAet50UAPViDzkBjBPL2ChC/E4xvCOvQ7UP/O5+s3xE6+sjKyK/OVJtPW76bV52
Y+l4HOkJOvAYwUJI4Nfg4td4ji6norICmUzxjjdsi7GFOvwaN95KRSTZNhUXRyM6
HEaLudagubmRtw66gqGfyqVPUCFbfN0n9IfOnz4T6LIXQuBfI3RMerZcenq2FPJk
ooVZi7nYUvOk8+pJ3JP2qz/7cnUKUigvoxk6NVo2GyzXQPdFcJ6UpXqhiChH/ry1
aqdtsvNPEdbTVgQhPN/XZKiqxkLkyvglOEizEguRTvyT+5cpNBY2/XHh5HoU8KpI
cJM8a5CfYEB3skEwUgLIoGOGPwIp0X1eym7NbuV9eGzlspPi2wDygW7AD5q10UMX
VOADPiVWcqTuXQfpDHI5T18W5uTZUO9M8eeVNFU/bbeR6JQuRcKpL/N1cG7JYD5m
/VM1nMEe09fUxMMLLFkSB9ut0/gonHOqNqYg2unuKK534TU9WPl1W8nGMvyHPUxr
XHdM/U+JQlLqnhW4CEBcaQJz86ITe7Cxsd6Ud+nVRc4eAYLrBcN8CHAtpNTIDjl5
goGZgifGwDQQ8wvM4rYknUoipGI9ACGWkDRLpoJMVFKWIHa0pjkfY2RVnf2S1Fhf
ei7REKG4IYyKYhdXCrB1n9wEZCUMTf/uYuNzPS/eP6jROPgtEEihpy9R+I1n++8S
wr6UT3aPKAGMXrhtkfokfkwjQYrTT/IKoodFEGsMTxtypONOSIToR2fado1Er6cP
s1aDd/1Fg0SpAPVn9vknSmvQUb8oyQvu6yCJRSWbw/hTpjjcPXjcK85u8iFQb+GW
BHbgQtNIfONS9zshdEDjJs3gDgskiVXpH8jGBtqM80YEWtjFwvj7geKmktW+zPju
eujb+CHxV3Ja/79MtEvO55mJ/188Ek4Nza5upisDNq9F6mqoEXM7IWgukP+BRVkt
GIA6R9sC69uDgxyHQioZsgkpY6O+omzT1JfJyGOq/D4SHNKYuguPn3/sQgm0AopL
lgLh/wzGEw3RDqoubYhYce1EncUH7W67Lit88Nasw1RjSbYIS3IMx+3QvBBQcAKE
pNfVDdKKY4lrlHAW88MJLcEfQW6BWIcJU9arF9PeY1ymjOUe2PJE6gLBT2MB+VFi
jVbLGLMnHEn/CwjesNVogDpb5RmQ9JD16isDE3bFtqBZEdJzq5ABlWpZXJM0jqFN
lEqXXStqhjA3vSQmSsoU23qaJ9YMeffD96MMila6OJyZL0/1Mm2tlKE8X6rWuAhY
le/CuG/ewmhDWlsygqaZvy3wlCjBCHlDmzm6HLC+Gs9djnLPJUhYnpI5okOlF+oD
4mg9OcJjqEoS6qegb5pMYCmNbhkK232quT+jq/V0T5GIWu9vAc84QIEgcadKPYVj
4lL9M/55evR+dYxvP1pEb3BHW/C6bqe/l0FLYfdXJdKuf5ubsfMDJBOvo0c///oq
DTwiZtUxjPACYBmXzHaAK9emsmcxBcf0TuhjFdmnvB1Vc5BLckB5Pr4KjQ+L6YuS
utF2XblbNVabfEY8dafK1SaZuz+GpEKZCPnvqOY/75tB7YzwVzuKBxjBt1HMfFPd
1al2oVHbMsG8Y0X7haMua+xnekYLVS0TyfNPqjD239toiThXLG/D/Yz3dYVVnHSI
NbAA9PFQBIVjKZacsjnWnu+wCSRrKlBd8NKlzzi3n1bijEYdcYZ35pdD+DCuudow
faRkFWPbk1zWilydJNIF6yu9eOcerx21z80WKbPebAlJ3lz4UqBkgRS6LbpsVWV/
EM5Ulg5F3Qcvwobi3sOG9mnKsWNP8+Cu0SxapNwzvFUyhALKgtj7PnaXcE9YCeBI
qrJtf9jqMgjnH/Qfx8ms5DEZRms0MXkLx8nHkXHlevWBrvonOnn4rE/zeV1xGNPM
qAbZRxA+DM19ylyR71GQ24HvSl8nhQObYDS5plr9QzSxFLgwMj9LzQFk/3XJ/IRd
2tQMpWHFqKb63bwgdgRfoVsDOKTGXe9aYRhxkRdp0o4uJUqqSbJ3ngWYDoyKPvKa
CqkRpra1UPiolgmroc5Jnd6QnbAP8FSEkAraWLMY6i/KiG76F7smgAD9V8hruXfT
04PubHsMpX/k0BPXHPASE8ORFxud9kSWu439EnZZZfiV9xNy36JIQuM2wrW+vVEE
QHkCFtDLtBT5/OOK/eq1uqLD8gJ4vi6AIgBHUa7ny+fP+N8+f1yUYcJ98wPdSINv
jfHA55qSvy5oBOZjoU6XM7v0WNIqlgY9GvC2ROiCW19OTuvBUDWxqJqW3Kcs0E85
uDyJvqK9hgD+C/Gaxro0Ahtkpg/ZXfY7YsqslzaXgAlizC1MkBfouQTxH7RE4wAJ
CItHz4kMJ6VsBrHSv3Xo1W79p0QXJZY5ZXNwtG+MbrewlS+BjW8yajg3/Kjr+Ldp
jU30BsBBFBTbrWZj0EQciLijtPZgzwTIRhn/ITtavzSg3fBIbre+naaTgae39wB9
x9fqcDWA6VMkXs0AEq8Z54jynm0R1+z3ip9/w3zamRlgN4TOyqbrULqwRfQvAr25
izHFf6n0NBpOP/7I5LOVV+AmxFrvbXdinkGsLaTuweMijyjSyTgRCpBVaK3LITr+
648hkHpmlmigZ/Xdxa4Te0fAKdnfhlK3b/BCM7br2w0WYDuAyLS+dxfc3rT25ABt
LBCkCjOTDytSOuyZI9MvX+2EYXmGEg3BQ/GwAhNRKfCbcHTAcO5cN1Iasy3tLXEJ
4L+KnzKpheoFDgkUAqUNKxA/xbrW8c44ddCxm7tQkwaIJ3byUUDOJosohsoixWho
Ji4d+rkb1itRyqpbi1cKNctgZsjzBetfJVO/xJYO5ciWIoaK1/yJfZe8ZH1/coWD
SYLUI+UBRz5AFu4XjEq36o3pjrveIXGu5l+OcUYdNxruJEQ4OadFa4lCR9rg5g5z
gn+eS3lCQEidxbDY6TgO4sQZc6NadROntwul0I4hhhlufzmFu2gdnEYRvOWANBe4
EMpp3rvtENtb/v4wk2AtMKqx4N0uArZDqMLZmRf9L06atRlKdGvB7TnLcQX+Iexj
8hxHA6FCoWi7VKEZAg67MZ8srLOjHkW6gk7+W5wrP2V+K7kLgADe3bvc+w8kkDiJ
Wx8mPvJa/RYXazIo/RUzUAe4idZxXyPCe2om30PGXelt7E3t97XmxnlXE+raAF+U
pxrpWrH00GS9xPBvfjbV+Uhh26SuQn3Z2A1qzVFyf+csD/16kDEg03JI5hJbV2h4
tWdl6sutExfUUfrSg2PDaKCUQk/4U2c/iEKe68BlYJH/IeKeZWeKFUfthVyd8rIS
P6TBi/5v2s2ZhjJKq/+anKDKcA/5zuhkKloneZi/XiYwCdrngRMnuW/GMEj/25Wk
Sh8XJuXszX4R/OypmuEHIHt+QcNx35p89btMK9f/STb2VsHOpvYacy+dfUYlXLr/
cDz8Y6wvHNMw2cJXo2CkfjWVc7kqA8DcaZs/qoAakcU3leGXi5brYh4B84d+11Lt
Odk32rCwtFVJFN6CTdgCzGkFuDeo3LOZpJSP55Hk030RaKxGw0+dZO+CAQlo9iGb
/4Ey5+23YWXUGF7pm/nHkvrdEemrhgtb69g7BJC94zMK3LA+44ekgGd1cXpqkq7z
JTYCYEAb7TlZ704Sxf3O/6Umf14gyPWXpuSKA3Yg10izn8ebPSBE9aCWJ9pKX1uB
+caOZk0xhUd4E3AQtD1+goEZlHf7EOTYCJ8PS1LRjvhIzm99/xLv2sYeHIe9v9mN
Zby6WPtvEtiNL2OoVwvbHoC/N70gMKymEa+OTy2aWrFeCf+7P/DqtARhV7mWmdem
ps2OPPYDWXmV4Jy3EZ8xuDlVs/KTcNupNrouPyKvZQvAPFjr2BPa6UtQo2irP/sC
PHOFrwo1Zp3gNgg/wHJXaFMWbsjYgJ7EbUpkwoDc5jc02Y11kbcvbxhq87mkG0f1
Tdl0lkSjmG6GH16U5TVCu2Tgfxi0nt6O1O3N70IIxuBwcnDI7wW/eNexwicJSoKB
l7QnUas3g+lwTYm66+EzTYkp4kjM8ui/NqN1HorPoWrodBrJekjja9pffWmyt5NA
obN52cCQsdKaco0Y4k1G2jiVgQ3YjasmuRevHTweVXcGr1gXZM8q0i6iBgyUBHLy
1kVmEN8mFSZhTYy1akTCQyHWR9HeASkVQ+oNS7llWp/4kyf8Puj/NIAf3otel27+
Nqo8+vL/9JJSCOJFfyRuBOdVfuv5CY4pz7OnPm8WVqCV+MH8mjdRudvbkbsXA+AP
SLprxbdWNR2gGLT6PJmy2dMWzFFAS6HDeSjenyAHccgmZG0XNIIzq2rZRznRSkpI
FKQqdz+N0QSmEeq9THkKdsl/C32+ltSlLic9f4iIU9Nm0nwvP9o3hCYA5DbveLlR
lex2cca9hxSolbwukYMiGKtgZEnehdWKh7Lr2ziezPtR0t1UnnDNUksWCQPiNiE2
3gf4KYYVSpO2MMBFlHckB4UjRiRQaAeIf+rO/bWf2wuJI5qaZcABHCoUMzDxA3kr
nEEdlxPdIRNM6exAFoMuy4w/ANAPDksaA/UAcA0CIBSRPen6Sq0IqkTl6EIzMQoo
ia9TiUwXteNYtJC/IwukmiZpnO5iWE+4hBVvDDeQixV56lUyADLiziWKlPauyhIw
kwFFGWk3Ru9AeHcKXTiUpMEqdnlvj74ZlW9ewwV45nssoGyrDrgegZqwNeI+8j6G
x/sL6Na3UCe+14iwMIFuXSqfJuC0ojGXe407RSPSAFXTGvnDNg6va24c3md5N9P9
u1UXyvbCK6Y1QkEoYvbM3ZJmxsWQngBIuYaOE00GtipV0LYOcAlkdgjDjqmVH17q
fUo5HuBs7fpMUpVx4ZnVYRLEx12vUxlBNZwx5FNTI+bppFfOtD7ztSRGB9qOI0Yr
ldqqtLIwcmP39WmKIx7JiCrhUK8hKN6/1k60NLiLZYSMP2DVKkKhwLfbOdPZWHD1
0OEAWvQ0KYcJMscW9VBsYjm6GN4g/6Qn7plmq4U8j6PXnRuCfQOLYdC9pxlBI2iI
y3UL6iZGJNI+zOp7uBOZ4oFeUbHiaGAzxThWWqbSWVoB8qgE4xoTZlq6XdBuEgZo
Ok0k1DDkM+9WK0PlM/AfXR3Wmi4fbcMdz8wKPuWR1ER0HjCcfDg3Bz8oHIHTjRZD
EZsR5N21C3It9ppLsQfA79p+THJPfTQ0hnrWXj/B2es/vFibfM0Yg+pyxh9ro537
LDjjZmtEPAyInpZtkJHYlZb1F2D2tnY+y5Rw7nQI8u2oaiVJ+NJc56gTB/uy6C0k
LBvrhL7GMNp+rg8xPHvfsnKvZb+s0K3M9DgJHoUVVtAhy15Je9wLGdaOncjYzeg1
jhSb5FWZZD5vYGMWY45wJfX+OEBPUS+2sQtaoaCw7tMyo07KHjIryJFhQud4u4Nj
9nJCtZjCA907u9HJPqOiTviaXAVuLngYzwA2wMLa2+45XmKzlnMcbkXpQbBNbpVM
wWXnpgl/sJ5+5BQCinTXYKjRNvD3XqvwPZu04MursS0H0XazBEGSjOD3fScO1TyF
UGtkCDmuO1Btfyh2aExrd9u6QOpmX/70WcIZd4a19goya49I/EN0ptX8r6QjnrBU
F6/21c1LYJOMpIkAMKs1trpY2FNtBY+Am84BGZHyHcGmEOSiFhPnCpXmyTd5o/TC
qKK9LTRIQmsAqa0+PHpXpW6W890/Zfj5hjrN+sTE+xuwnV8QM+LRk7LTLbF7OHrn
DzdAiz0DLNNyyjMqXsWHKKEeMdc676h3AsR+KPCI6zma/0/eWTHlbDYkudvmbuhD
Ry7xW4qd2iBre3ZWOnEu6KqVcyCnhxsJkQECQBGboGZPCXf5bCIjSv1kFE+1xcEI
buaOOL0NDhc5OlBI9+TyNO9qo65ZON6sF6WxFFgNs7ekywgIpBuv3nm59w0nWXfq
q4FXlIku0g35Q87Kj9Frqm2QmFtK8NJ2EqVKRrlFUFK71J/ZnK9QdrFYtosiaWPL
hVeor2pKmJ0+q7sUM4rKMdncDTW19Ndibdwbf3aCiDV+S2Ru0HyLg35op7eprzHP
ONEEGkv/yZR81ntG7q5omjcRx88ZnWw1eOpuAOsU0D2EbJg+dQjnv7MV12fMy/2U
R1IWUCnymaQQ4NocIK5W8tQ2ckOCJRxM8mCYRxVeqN4U4X9LEonct6aaAW5noz7a
tQxPPnAa0sckhReWhCKg/kfcETbN9igS3EK223GbrOmzO3qGJjv+M5rP/+6JeBsd
4PXoghDHzuNlKHtYMfZgdOEFZObOGWWbZl8mrtkV8t/6Mw4LS4OTasLzP8kZHZpg
J620CHuPp8oFWVvlClknI78h9+JfHN84WglqEZveAwKsne5nswogeVysQsjy5ClB
KqxpxO4NLSL42KlUxuvL7XJ7Bsm4KkrB/pu+NRaAZmNZOmuOHLhl6c7rqOdGzrDW
TTZGuzYx7k91niiwkCHq/oPbNg+ahG0mA8TIWsdZoVOInKhZk1XmU2sgoORXPLF7
6KulaK7SGFTk1VKeI082IC+GG5T/NL8RjJuuksWP3EOrbpgvQLQ1zsNVVW8ayeTm
fPKcQneRjaDyTTfcls1Nijd5jlxHmi+c8AXgHazfaFevT0Afh2l5wHFUHmwF4TK1
PeNI/6+l6+DKNhrGptnnXxJbNGaRsqYBDH4aLCRovPGcUiteb/1MwP22RFyhuHuY
EUPmrNHrnK2PYQLOA3McfM5XZdghDzeX3rhazibO2afhg6InMubiv6i+Zzxl4jnQ
Jj86rC+pX9i96XVKxv9shHP2J4/R9I2LmcJQ/ttxJTYnTGePdc0OhaGcqbnWwgmd
7+Tm+8LyDEMUo7CyzCy2XiMqV4GwiiQ1+zyarpieXlaJasEJp8ZBigvujQZa8qxe
OdgqEBMxr92zk6WFWFpQ+44ZpPrlz8yQdcPmMxPXJSTgmyc7x/UIGnA8nOFWb5zT
en8BvItlHyP9vHQAnGH510GGZDvDri6ZhF/0102tVrdVBbsc/4QzaNf+WHsqq2Wo
bwDMt5xnpJEJrlVQ6gB8/XADdIUSfXbLkCpsKEFvypQFe/8gQUY8C6mvdlB1bWrU
ZPN5KoWXqUuBwv1zTJnIaqDDQs94pZCsF42u7s1pLMRxftIv4/VcM1qSXOze5yZC
yHVO+2zJKC1Ow1jZSSnqlkWM46uj5HugvDglwZu5jsmIke8Gy9jQG6fFQu52U6bQ
VFArU9NLiFL/e22zwbPR9QlLSUxPM8MS5ZX0WwOkI6Qyw9e10asYLeqb8ZDRUCI2
0BVmzW46yiFVafrIzyWoU1oMkOmqiTkicgLS9JkzLDV0F0dQrM1jEPFOZ3y8qdB4
xvbZbLXl6+FJ0SCvAA238pkpCkSgU62ctASJndo5Hbv1iaxARbKpVAjPE7unA2kQ
uiE5xgEtyzyjaW0oZBUjRefx3Nz9YkzbAWk0gBt2ktw6zVdO9Mg0yCD6FW6vBNHN
SX5Pve1c4i5VQiee0taXSVI38A5srPTn1Y5kfmKgM9J+4Y/gGZKfr5svJ8Q1cFnZ
aGfG8vyKNOx/p+HFgbFBZwEImG6opmUCR+/3CYEUi2oqENhX0mGOW8A4abIEP2Hk
rHEVL6lYd7MI9wLpwKcTX6TS05o/3a6caPUTl7sGG7aX5iE60WrlPATkMFQhQcGd
XhFWA1Lvh9239KHABRXQUxQdooCEPq39+ixf6pQLBYZ1qvY/2rwCQCfeZAsMzQsh
ghWMKVSbguh1vCEN48kRB+E88QU1W7+vfR4Y5bX95072ukhppQzEGmvgjTtqBCxx
TTwmFm9EB0TvHq89pTRzDFDFP7YcWJfOUMwNZbpP/mdhYy3/Exwd7n05jgwZCtCq
odJos4vF2Eqygmo2WCzhFngfypWCQRojiSM7lrOtHgAozMEq41s9env2qwzsUNzV
iEF9NY/V9ircwSW0bo/cpmLWzLCc5IDCH4LUuOYdM9ir4tzjftJCg5++2vy+nFRR
1c/hQqaHaTWJ2WWLFlM1SXyID1f1lusPpwM7AWM/+ypp72GyCCXcOKoHRFYznP8n
ez5CzTGQ8u+5Qfw7cj6vIqV5tAbV3tVoR1YQ34D8pBC+A/wMdubguqQLvwZDvz2l
T7vEoOo9SrZngHHgVgwdfg3rYORbu4VGEHNyIMww5qI/KsqNJxGRpjBavs+IsHCl
sWCUlQJ7XQBQM36TJO0XRzTzzfdUc9WmR4mht0gb6ka7GtMwcNr5+CRrLtVxGRUE
VzECceBx7/wWyuoV09bxREAr9d0DE1y6+xcRyHb45f5wc+2A9Mtk/6xNyhBbPuGS
h6jXfkouh492+hju4w6AMogpbWJ+rsmpSARO5Fowf9nXz7GTlL2I7OpafS2DhMuQ
CWc8zVPEXVOmC3kC0YZtbLJGGk6AQ8dTgXLqle3QFwXp5VCDlDiEf3zsL8+tc21i
7SgBwGm9Ur6jsu1CM9o/ALZ+vKCYv4O7IulK/67MlaXNZcLkkl8Jpb61iHngXFeo
xcmq/SiVeVarzHokXg5kXzpEDnRhkToy+U9JWGqfh+Q770/aekBlHrCE3ZNCQleW
fXvD+Myp+xwTv5oL8uRfE/YlHWWO9f3FMYtwIskMH9dWWQmDZO0tcauwKjdfnbR4
Rg8t/tBpFaHZMrSsQQKNTcZ0naW+WTOmBXkBhe8qT0vucmAQSUb9k5/LtJU/8w7O
IwCDAR0lofc0bYSbcPSzfY+ZYpwjzS4832PHLXr0ph38eHV86TK6kAx9tDsGzms4
YdgvuT0AXOfWfcQJqZ8aQiAESS1cWNV6J05590CEUSR1V86fot9d4u+CFwnAIRU0
FphBqAJfKDuF/3Xpbxu6jSqqKItF7liy0pjwb0+Y/NZrQZvKXJJT7YDiakCFTNB5
jbESO4IJT3krTlTXeZRE01E2WsxNI6tDCjjkc/5yocYRyMNLBqXZexFlHQG+OKIX
7+pPXH1HilelxUdR2/nyxlvLKbTR6lIMPouNSrMwnzvUTa3OWaWlr7mPIs5QxuM4
ZcBIYViOb5NlzeWk8scsvFHxLdpFHwafLwp5iXP48EU1De7TO4OwKo5w4huRpdki
ezY9o7HWe1nWhuoQaE06Tht1wQdCGHlFbef+E2dSo9OGh+F5aqCQcHx9RQe2GxP7
mseiGyYrmMF0MDwcslUopX62ZDo3zfl/IyhPJoqh5mywt3SiGz5r+d9mKH9yXSWR
LUaNmk/sbfYR9O9pek8t0sU+8IvxJ7Hze8TJea8hQuGLBMnsBuH8KA1+bDWeqSyy
EDpEsPlA+taeySGJdcviKk0WFAP/CRCYj2fTwRg/FfqLfshPzi20G86zOBLfDCIy
sV5oeMWgKdCS0M45QXnLw1igePi2zk/kAFlj7oxTNxJIOXqxFIZZz7sob/m/V3pt
FB5P73ERWCdlPuiZcqbJsKV6aMjoUFa3n+bHEcPP2tHPiQxtXe7cHkMGIcBGXKut
xSUThy0/3z20U0MJhIYgJdchGg1oNy44ykAgBTKBVYINYlhB6gN3dXcvjwZo0bO/
oqpZiWduQaTX7UDHAR7B9HwVXPIDeZlyBgftJGm+IVcfPLHj7iLH59XEu2rMHsIn
ymn5wR5rim6TAlNvX5H1sBYOEmK7cJ3rqo5LXCRr/gXiOSRyHrDP6dwUTy2c3tiq
LEWSkeyRqwGqX2qMZh9mZ2IcTnzqbgjUVYxAsuLC83AP1ZQ8ZtY7HB82MMYpLzLl
Y1/si7rdmC8zLFMKhZazA13NrHs9lDuWHt9w0yNhlqhvOel7/tCmpCa17OxLX40i
6lxq9hGOXs8SgOiuM4hht2J4j6xel+Lo+y08QWw0lv5oP9EklkvJHbeUQzl3i3jU
yGXqvWyUtAFTX00T0VpoRtgvXHjNLbuPOuS7Cmxygd1OqeOibvKRArcdKJwKw3mb
iqN0Obe84+PE6K83JT4kPvICMcHEkHKgCxeBOOIsOOcKZ184SGxmbdC90lYdlp54
hU8eg3Wo+FHjShTd1tBA4L+xsIuRMCoajgGUiUi7vei8hAvcVlj+lm463IDKKFHC
Ty9TNLmekV0ESc3qKUX2k+AKEhMcIb2QSOP0G0iBch+6lp0l5LnVkAXkBK9zn0Gg
1xiVQQ4Na/c/Bh6JkpSkM8hJ4j7HpAwsjF3ahl6eA4Dw8F811qmGqIqMEJCHY/rG
qoFCIMMzMwddr265dccwOtxlQNJd9l3dWRqGp4C+PscAP3+I6BUA3E/wGKGNacTt
UflxuYwNgh7390kwtYhN+X8IAiQXkwtg59MskoDfultyHgwgIc4yFa5VoEOd/cUV
XIgfR6UV/U1pO4oy/RkLcJ25L7JLuw0OmX5nc7ujHNfp8SQjR4W94vStfX/pKD0q
RAZzawD+RoFH0Y4w4j/Ibao//GZnFK4gi59lbxxEOKIce0qsIvRWu9mbrfvIJIiv
WpBXmtwyfnX7m5Vrw8ReSkKEdHul7KVYExo+4lHi68XC6exdzfWew4iq4rm7E/NP
aB+02ZQJoVjBjYQ09SuyaB9tyX9e60QX+CxHC9H2Ens9veB9TWV/FdqAyAvKZdPI
gqP6w+Zf/cPfiQ+e2BCpkFol1FZ1txHYaEQgJYZhNCyDAS6Id9sGks1lPv7rWNEl
9J54R6xf3uznpmOO8Ec+YV9fi6x2MVw9sXl85njZzX3zkV7xCKX1FmLZzRYPTSDq
qHYowy01/XSzIh336YY3lm5/jrrbm3oEu0GuvkbkfIn32Xeg6xH/SXH9kJLeB2l3
90Mc3OG+WtV1YfYyVG5CKzTjnsMEzPpv8xHy4BoLQFnsVcc21zNvByyugifxrBeh
fjJVCSHB9DiEfxGnhlSDdmaFycnxlbKLy+WEBFx11gFaE37mEbD46SlKMfsycIjl
yvbmnKnFGyhgtztBzc1hj14h+NkoP4OgrQni2YM5Gd7p4MHBkDs3qBWjoppzYx2E
FJwsaLohJ2Pvcz9qhNOUDmf2BtGSvZu3aO/DtrvwifLYiuGbfxPjdU+lyolgzgvy
PRTfRAo1dfDrdrAapA/82P6upTnb80hl/pS8dnLeRlye3x3aFGZenUvljJwY3JPG
Dhg9m+jkB5Vl2Y1YYqXTaUNPDdXAnbr5w7I6WKTtY577+ZtH/9ikfbVAO5YZQyV/
mwN2ho8OmS85ORMbqt1Im5MohEGM/yFS31MSn8HOmId0zM5um4FsUQrRCwywMEZl
gCCzPHbwsvsAgwcvnpcgF/XDq+G/micYLEtcJwLP3wKMKdQKDwUSg1TVeVj3HWWb
pq0YK05+jmxBdy1FHVgzKzAUnh4VRbTJBu+ewn1v1Wk97TQhbHp5TBP1dhcuctkJ
yTNSiXOagVAgVuMM6qE9CEOLCqZRS/sCzrKq3R0aYGFRZJKXVBxorNIazaHdxK0S
yrcUETYa72jtCm8z4iCR613BPGN3hoBLwbmb/5tVClkxastF7E5PJ1v56CP8XjPF
X177BelZ7l2EBYKpYEshPeOizgkQaB3LvueeI3RZD2bwz8hN9PP6qNjgFfid9hDM
8Wbjax4DmASB4M3hz/HQIf9PWy/lWvh6YaunuZOJ3uE+DvvZTCFmQDnNU7RdYRTA
Tyi3zhW8WXaTkX85Oow/fcmp+LF8kxfXMgDFe7qlrTv5qWGxarrE8+8/9qcYhhjb
Rv9HzlLUV1qkfQedU7jOWqB7B0sIGpsNSar1UJlXCURFyEiSaSIYuk8MfTgD25Hg
nSyw4KKHXunF3Yqqx4mzdbMgmZ4FigQWfmAztJZpnIUjpLvcsv9MqWqQCp/Xx+96
t/iYQir6jqMBu4ExZyNnw1WasZBDTSj50OSSoYmNc7BorERnIsqmeI+uM5mpPjF1
LuSpCEgbTgcyl29N/rEe8PUOwm3j5LRt/J+KgRE4LNzWK5aVY4BUEMC5a0Zlzv4L
L9/Q348/JbB8Uv4O5+l07Q9iEEDekouWe1gXr+SRSN04a1tDr/j9IklTDgfZaDCW
id7oSLXVTka61ryPUeThJZ8KR2Qi8jwN8aq91ONVz6GPqmKsKOrqEbHyQLbVqvk5
rv46xcD4kmTq+HBd0UrC3KWHydjz1h2QjI0UIIf1NAl3bZIFWlQDgNMTnur/hlK6
IpitcbdAxM1x6gAH7NKeSk/tKx04nlVEWIGP3JV+3+NBqzgD4khvjCWFvLe3moG5
2gmSPQoJst9PlkV36q5UcLobGWG/teepVNz4x0MRff1Sxhq2UbtWQYYr83n7PK6H
l7WZXLsogWgqTftfUKKPrYL9ZY+jJ8ut49rrzOPr+GrorjIPgc+25B2VF7zftxBC
/pUIOBj1ux8cKS9bTIc0KAuQI3KpY6NUsyFY7v2SgBaQsIEI8UqvfhpY5bzVu3N6
E1TDS9SeiF1+okchzRVZPu2X2tHDYXm4PhZcLi6MRIhw+l0d1EJuySyutZseTk0d
vRQibsjVgc6Ws2qc7ioM22sF5HCUNNd4pB3jYyl7RbmMM731zYLEDlS6PtOqjVI/
ZHCiCZDtO+XifFO8/+koEI2o9QtdfOMbHoFGOrODv+3fFIOsY+w1FlO8MMGFtGUq
k0aJNzUKIOu3tR4t//imjd+X4zoMJEZJfqCVBypgODoII+Vop0Lugm/mo6FYxvpL
vIDQ/poaJn7ErGL/Mmrcz7SJJ8I07X4xoCgEtHj2JdYZPpPb62Wkh5KzzxButbVX
StucasrkNfsO49mJS+W7w+bO6kI9CDJQnPZqSxZ5Bi6WGj3bZGGJs5JGLZDE0wSl
WnmmxVrhA/3Xb9+EoMyGl+bECLiOz/4yzz9fJWcurr8+WYB7MuAX5sCpDyZoyzb3
4KounicPtxiEkRB4PuIPn+hk7f0a/W7juOUl6KWRH8Mk7QUH7ARXdQB8d5fVNL3b
Serse632zVQZDPkqeVsRk2mxcv37a1JSlaNKl8RYwh5sMEc53/hvNcLPGWoKim/X
7VnYijBF1s3NUxDaU/F1Wf0SNFuiDTfJU+Yf07Wr3BPHPTmBXlRBbDrmbs83bw00
+jMdAK+feIM+76sLX6yeqgw7XHd1Ybm3uoE+cGk5ujz31RPIAf/KN1VrziI0rl66
EefiLCAuXNu0TzEWEYv7YW47YuFK+UGpYvayyC3AQgiOsALGlUfdWqdph7wETa+O
xvTbC+G+aFU+/L0fiH/wFXbMggaDbPI6hCtciOAWkNrHxU9NIWh1yVdYS1pivRiQ
CBeW2twe+YgyCwGE4DwIkpq7kuFjU7OxjygaAVTcOeYUqoRUTetz26GYecYk8TFR
XImafJ5vUah3oNc2ofYXei1W0tewMfvNrMYf62Bb/5yQApTa92i4D2JH7fUFsMOS
sP9YtXspTO76zow6rzNvihTM+6Mn+Tc1G1ovQbOzwo86n0x55IXiQqTQ/ZsdpROQ
c93A+Yxg02EkSxt6MNRAZKFSACFpYMIGP/J6eh8rTbFFPPTT8n4I4gyzQ4PYSoUN
xR6C5n9RjNMwLswPiVM7mdIs28W+GIKWsl8173y5vHTVx30D+/YR6MfSLHIIpL3T
uy871T4ZTRcOBITyyYXwLqZIyjGFiS2gJmX2/U1RWdtvlCUixFbSrzSdXxNvNUhB
0KHqRyabT4ZVdaiy7RIHfETPFWW7f88WJrWiYhVjbUc8gMjnCr8SwfCrfT9pg+Af
RkQXwr5SupgM3qLX4zdii5ybFPimiG16ZRCVNV6p6S0lyOkKQm2Z2RDPESCQM0Vu
xY19usd3/o383VdK6UYmCVKqcHPdH57TGR/kiZODJofsuj1wTyQCP9DBAFbYBDbx
Evmg9qyu8Rp3dB4PXu34iCe8U1ot33k1SPtdRBx6i47n5x3lMjI6XPyjEI3c7anZ
H6HB/uqZ5nlVjOHp31lQ2lra+EHpS/8XXR/Bj3kyOUGOzIEUZma5193/U6Ut6cZs
nMUTOxxK8b4S3dg4mnyeYljtTlFmfSxfJMqcgyyNeFdkmB394kAhlwa/JNhZuZYf
Se7cythx7crEBFmaH/Ece7fijDeQ8v/pxZoIxz0Fc19UMfW7+l6tO0C3cG3Q3jeC
LgrLvomJk2z8LIXdSAz4nVGXTliIOzVJkPGeaApYKEN3VpXKEVGfq9M6VYQqbBPI
5ZF1neiQxC4AfVM8yVdXS6BA/TJ8cjPQRuVYpgTyPl5I5vBECXlYiq3h8NaADH8L
LTAfhr8Dv73h7tTV3ffJggJgykb1EL+KLznDEE+U0crkognRjI+Pmy0J6GJxvKvg
gC35jSzKjEDe5jjp+lJgQAY22pczsTpc797P8lCK4cnLqJeEKiX8h91a9JgnPX9V
nNx8Gkgem2BTYL+1mn6OVmiE4apyrQnYit7EfNYu4Nl4JwDGDvBmgYwAbdDU+5K5
He9E4AQJeXR4NdRGxg/0KuLex9d555JVj4BmNuX3scFuVxCrmcw4E1nFlGe5FXmJ
PQwLw3ogb3j7loAqbjtkFOl5h00QrQF9W3v4hZfylnuywOT2+DitF4FRfNVy6x6G
ZMwf+VudnGkXSCOK7AcvxDFWVBds0t3Z7huyB5oClWxYpYX6xFO520NLuIVKEPfK
5iQ+e/D3uUzbFCSu6VzLWrmEoa5h8G6lasgeo2kYoY18411y42lIMcsjgyWjeqXu
gKiWGoPh593hnkVT0vZdGOLO0sOITgekd2D6LQshIFUKaP9xhSFrocBptYOxnGnR
f/LzxgukzN6eRaWhz7P544FhnLglT08vrBvowy4qPKAQqa6HPqYOGpah/oGZ4AOp
LMQPPK74DH37yEcjd3QRDO2JR0UG4ibdsv6k8V1Rzw/eQSN6lyxwVtMJnWRJSUYH
0vmt05bOWxCyzoDD/CnCY7qQBtzf9+ntfMLpVfYP45oaQDECX/XzzYvkm56yfCRS
5DuIjN7CyTZFTCUABrjMicg8t9U4x0CNhZDNIuOqOfjf8f4cIZXUn9qbV9a9Mfbh
Z4ojr7pZKAKs0oxDM9osXIMEMRbxNOCuSaGHyekc1Nw6pidTK04SqGJQCh6bWr8B
zK3w7jR33/wd7ge/5PCgWqPXhpXRLKLycbqcmLQ0q1XUV/AG+N3UKZFDYNbjQ8pq
NI6ZUl3u6XSSEa2ualSwGF/BMQLIiLV9avSsK79+SZ/RXh48o0gS7MKYhX+KMy67
LYXu+/0uVtyBg2Z/67aoSavrorrZsezx7+CaPGf0xfY3wM5+3hApqXHEHlZXeifd
pnpUz9qGLdlbOLLFSl1out78daLZ5yEjHMbsjBaocsHaMeBsc6DSnr4RZ5Se9Jwx
KcoOmgT5hchRAq+UqIli7BZrgvtQ3JZE8jUUP9FLfqgIqwlu41sFoYiTWxhMCCej
bzdKxfZRbNhn7RW7x/xyj75iEU1waZ/Xs+B6s7LG5gsbhHHTCsWCJ6L9njjkPZlD
57Cf6sl/tCy/t5cbQEuXavM0gUA7BHsZrSOzrWUO9wlgrU8SmP0CADCYGNeJbZiw
8k+YDpFKdIkGmw15vqlvVEeV/Rpjlf+JqE8oB5uO73FTPLCxXb1c4LwM7ozrNN9q
AxZLyITKjOaTQnHsIJ3Mui/9RFF8G7EdktSJVELulvBFa09yy2DWVt7cx5TPesYt
/u4GrRBCaUL8u64vL/EBQ0O52ro6w4OXkIhfs1O4/Wvk4Cw+QFNiEgNQK07R5NoY
NLwvOZ/qHU/IC+tW8XGSgl3Unm3DDM3i5H50ZQ31z8ZS1zzEo7wvYSM19swvpPtW
s1VaVZxrw+30bTreLdpzMCwHnIexXufrdI02lr4Eemd3X3nksKYzbrxszVHQRZr8
9KSFuRDcGtfU8wyoJmlbWayLK5xMZkzPJr1aFqo/GjhXBvnwv7jZAxoobRM8Q17e
8zhcK8T8paA/dxbRqfSinMfCU78NBMoNhQeatcmEDqasdrcQziSM/JYWlY9wMnen
15v/JnDvRkZm3p/KKcRX7aTrVdTGKMdVWYFqABfYwdesJTH9J0SSHsp4VXfnhWP2
SQ+VrfO+HI4lC7JTAJdmz1gMHYw8x60s18EavTH5i+SzY+uX361aaNe2JSPGlfB1
vZPJ1dxF6neYD2+9KYfunbWEhB8o74atM5olD46bajUOUECZqAouV0kJHEyX8/1k
NHAprhrxeMwqL24JbF6grK7cw6bT33wjHKVl+p9E/B9s+h+5kmsGwyfwatDdrLAj
d/lIQE9pSV2jM0vX85k2B0a/+1T/aRKe0MicXrqd/PoJURIM6RlzOKnkGBswB1v9
psE7j6qWyzsKlaaRDxWAkNnPFtqzk+pfkN19BYADH3zYI/ig22vwPBLY92NPR1wu
/Fz2KXH+ARSjrvrOfZu5Fg4GgM29+EBfRT/IRWLRLIiV//qhffHbuJ3e9QGbWkmk
ias8q+uVvLj/o0QhQQLrHDstCsdQ+MhlIA6y3pXFW7/Lni44WZ/g2N6D5x5nI1P9
HES2a1NZdj1mQRJc/vXqkkhBcUl23FRXs+waoeT4y3AzX+C1hD3AcMd/Z1aGgqQb
jM3JxxqibOVHnsGungd6HcUYrewuSskBlfBFvhHm2330HkofSn5URjEEidMNmipm
l8IAgld9BFvjyl7N2bU0H+Sh7EOj5Thq/iOJ8X8DCZN8q+cXX30Jf+YsG4ITT9zf
qWHfYFIi9paHvqnme1UFWcCiRbF6SUsipL5w3RifqnaWbd4AZTSExak7dMWzqyZY
bGHVK2v03gyNd5UqkOUZi4w7mxkqhkReB++xPgQenfyJigfgKRqOtJfZ/92F1UPO
b5BuF1RWYJUiPSP6hzv/zj6nGy5zI21seVAPHlw/ryt5w9776NPczsrXSLLRhSQx
QPhpuFVSiCqCp7aCC3+Jj1lUr9KW+kqxT7jnIHQNMKsdR1YeJQxpXmfYZZX+mtzx
pA5xpL5RtG0Ivi6VnMhmj8TR2dnSf1RcTA0YO7O9Gbj0EgggQQ6EjAWMzRNtcjYA
LOoWR9NMikEChOrKiHi0ARBcfOZcNSc8oCd3uJdbNCcVYskBFiHPXHcadrc/Scd/
5TInH76d/w3LLa4aQjjmFoLdHq+W/4ezUZk/xsOEj+fyWqqo6wMjM+EXwgIrEvBZ
AGb0c2/nCeqVPxxK8GTywA8lS8Td45wjNE5a90ld0cWSiR7Cx34TvfXpKk8u3Vha
oXl8wNcQPT0yquBYrXUbSBtI4a1xX3+zLCPoEva626w1W5gkmCbbggBKgWuEnaV9
RVk4oUn0VLcbwg4Hf8otVPglVKYsacy7Tq4pmr9JP7rLKF1QjJFKpx1RtkmGRwJ/
S1G7X89cte+4TjwoIvm8QrBmD1P/Iprgm7JUU2GIKfNYEydQFdkoixuGqyKNASXN
mSXHDwa6FCIsZbiZ1/K2Uwkqaq7Xs32QGapcvkJqy9KRL8hiGn0wfMlZJenSbxdX
iO3zIe3oV/kxwLbvMmcCIxy1StH2qfdwSWjQGxZuNtM2wYpPV+3XH2ms6sVgBa1C
GcLgNoUGKJ7x9+zrs2T30F1SgtsXryLZtAL9sE5/o16SgsEisAeXceFWAYHbclBO
CNI5rDq/X/Azn9LAnwC5yWGebn2bEMU73tvl5/FS5v5X5E1FWuTAXQaj2kKPReCG
fQyQHNUat238L98w/9XS9EyTkSoC7YXfJSZxmVFRG8F5ZWFzq5LaxTukREcaRpph
NZlKCiiF+Ep0HrelbcXPypTogIK9gESDXb4w0Yy277l1ZqLZtaXh/E+Tv0nKQVqw
dMqCicfy1GIikhNEHKOx0HR0+0aK9g8pBU7RzeN7R+tD3yrgGJw7d8x7nzJfR9hU
HKjgVkGnX0ceXD0lEiGuPVCWiUls0RxGxeGzMWwdKJiAgL54PBLS5kDS1ODOFUNL
pMDprtFD4FXWbIUHAmwJR7h1xopogm4SW1PN1qedHwjm9X1r4pL74w2lB/6PIcM+
9Zg+sOzy9E2YkK4ROHBSYx+uGrdxyP6aNdDcayPoZIpU0XbR1hQ/4+eZUCbydn5c
ZIAK0ISEdq3pcjaUK+X+FAIyIyUl9kMOIVrE7UsjE69JdMa2kvU094at6mri9H/z
OAgEccwjUtOh0mFvJ8LICaXmhu0gogWY7Erd6MPgP0Ct53k3n8Vs8ifVa2Eaj0GT
M2ueJpjsH/VJOJXf0/W158bmXJgMmAAGGtOVEAVx6U8J+TG8f96v6TyP0D+W7QgZ
svtD5gKdKkE5B9KvGP68EDYgRe1zvAElfd4jhiJ6AeFc9PxTt2lm77PU96/3AwFp
u2ARd/cjNVEIbEh41/kkpdImOMfriVxvHo9JMjcf1HNS3042KV1PWefaG0ux3V7w
PgUEf/urrHOcO5dROKSpJYEdR6Q77OxQkifdBAs3IjFrbESVGZOroMJws32OVOdp
nbnZj5J9uUAYDHt4DSRUuCU4RkQv2tyHCgrv5VmFviigBC/zRIbDtGw1EGs7UTxc
JML7gqum8N/+rKxaWQeZxFqyzeqKObI1gJuPJFM+lD1RGmChBVhHvtq/pxe8HxHR
3Khn4LtROsjLi+AGQKlkNb6MtRql69FrqgSpjq9l3oHMImNS7uElnJ5LfaIUMisC
bq5D9I43JQ6UNXeEhrIpHTw4DfxAzIz5WU3tzXm5bVOt2y/hOTFSdxG80N7Uw/i/
02/EwKRPJdfCTZ3X8uSC12iJijj5PDPb/nbyw5XnfIDRfZU6jm3cUD/8nlC227zl
T3i9oQ2LwJKQH/MQiXYAljX3eFKqB/ms8wY8VoIulG19Q13dVO0/7UmH+rzASqjE
Qzb98pbT5TxPeBd0bObe/oOfAqAC+PPyv5cLQJ2FC7JlhYHEkSe+MTF1sDqqkM3f
k8RNqJYbOaDz97peqXdxktpV+BS9UB7LoIzE958JUgZn2ImM6ltwuIKWIpeLV0EE
RfXtElcV5Kc9ygxy4bkVLAFC8OIj9xrPBDjyJUl+spJ/rfBpWx91eWLhQwFXoCbD
JB88uhncuniWaJFJaLY2/mtUsggjiw7guZsDaDoRqtJjiyhPXNzSGUrUsghDe5Ug
1mJnEcQw8C8T9SC3VfE6ni64sk7aHOMZON01UM1fpGMr08s3eyusn08zKb4z9HOq
r5JtIafVmhLVS11myWZvenPrDRE2bszDb02jujs6696rmorP1izW/ZjYzFMIXX2X
8+pdN4XyukaVQmjQM3QLstnoanilayEny/AOERpHVpCdM8FEoy9Z5flkLlvEdnj9
CgbJUCL6Gy4Ok2R50QKg4jq+I0hW+NnRH78jb5ydnhy5NwGpldoPipBG8G5NbD/P
2EB5My7vXtDgfPYEh6MaHhdDi8eBF81XO22v5EpCooeu+8LwF1JkrP+nEFo8bps/
IijuPxzgDDizO5luadACbI4M2iSUq1WjASLUG9RzyazSEyt3kwfd5FtwcwVWiEXe
Lsq+GCo/RSsGxyO/qo34G/3Lgk9ULPBXQmaeR9COfOd2R+apDTg7PFrZdTVERaUh
6kNFE88Uj9wqoWX2w0lxTE7Gfn1n94elrrENST17tsWlXML32IHRCvFn/A6JbPub
/v9kvXsgMZEwdKK3Df/9A793ZLXAcFtlb/Z6F3VEtox7zQothpeSL06RFVVz9I+V
Q93Brnkgl9fmM73qaFsytpYScBTV4W/wLt6wbaMnF39bvrzuzXLriZKOrznUz+9r
/o5M3fhiJrVKVgZQqVqsyZ+hvGsZx1Z7xtyaGv3XHztfZLX1+Qs3VIHbua4QNVsb
rvQcRA4a0LrPys/oThjahH2GZGJJDpoc0HuC2PRsB1ldRyBnjzg0e3J0J1Ygy84K
TBxE+zEejJwXB34vLvbM6h0o6gdL9ypabowa8nG1eUoJ/F7A7+KaNbpXWvenS17L
BoDiQhDoddMiMaI1rqLb4EYVoYCSQei2ZelUyS6v48R/NjWgPbrvF27ONMGTvtwb
+9o47wj9QntvF4dtAK7lJv4+0yq0xqhvln6MM50me0rVqGDucuq42ci3CfxJk9c2
RRSGXuwJ8KlfkNNP41a4m2cnOmpQgTBtBFZ7bcrdo+IRaIkzchiBazifkjpH63Yi
g4dBslprq/z99Q0ap+0kK4xynDmkR6BwwjxoXXMlsSG8rRrYdax2Ggz6xagwgOzU
bN5XUi87OJYDCPLo/cIERbLBmk1/4LEwwyZU2dnW20tlw6f492f4UqOzI2RhH2F5
4Y0IF0ONc5MCNGE/tKoaj9/rphNNxhbFsaaoxQQVFE8CN0QBUk2yR/gKYrDd/z6K
f5HpjY+aS2Yiq7Ws0dDHj7XzCihCgRziGlzjyGRQf79LTxRfQ+eAqRrH110xBITV
lvsn/RpZZkERFWDkwL19rekcbYfn/jfN7ZdsURNGN66jQy4dW4Rm3b5cn/nOddsn
t0eYfGwpNHsne/a0cl/G3GiTDXMh9bJjxP7iJu5xfyWf5Ahlpwhv2yTcc7ZBcFh4
Hh7RZTuOPuD0gc0jNVCiBn2ydktlJrSgUbMvdIEr1sRPBjIiHbaQe3aGauFXgJjX
kZsEy8vtKjq05TDeT5ObUn6Qig8wZrbCWHDPCbogx/kDKHhYvaEBIfgnkPpWTSfE
B1FRK6MYoQyuwll94/ClwcVFsg1SlkKEdIVZtNJw+ltsMXkexSSNUD2prtkA4/aX
D4zMf8H6yWDIkhHj0olDjob0LijA3mavd22Fhbt3NHa1lU82vQw2KA5Aeu1b9hdW
j4aJByCV75HBAdw5++P6POL/KXx8cGDWXKab4rc/mRV4w7/tyfnm1TVfV41HnWVj
XVpI0jQMM2dZ1n5Q4lXgG0rgLGIJGv+6mO83l8KG1G/aaaRnxe7SOwGnnEoAHYzX
CFdOXuYmGl6fKbiaIDDDI+mnTkyHPDieoIKC4yTSROX5HKJ+BOHOQW3Txk6aNIQM
GMU47dKDcGdeXDd5tOwSkI31KHqRNdemmW2ZNhrrmkHxxxMqTTEJ9RdofQYIetjF
WbmSWHj/oLMP73uVMWBN4uo38BZmgLKX4EwYsxUm9G/ObyTN98iRdnGEhPanaeV0
KB/BuvUa9iLf+Wb9FCcEaNtYRwhi1Bs8Cy0zlHxs1BHnkK/wU0eUoygP+vBNhdWQ
g4tVfmxYq3F7iIjxqeyf0qXJCsF+YCiCVVYFEiL+De+T1pF18sdWqs3SjQ5k/zVR
cv1N5CDyleV6FW9ig539jK7itRl24L1Loaa5Mvv9zDxxZBS2VK/W6Al6M0zZbhMB
+SAhK2K2uxJtfqoi5+e4EFViRfEfh9HaxxIbUZGEuhGKls8bkzMfHcKihrwU+LN1
raHvc7G61ufduYTN3aMJS8iXlT1bTKBUQUq9ZT6PZJ0Z1Wr+e8xO1AOBl3IAriHa
1AYBCat8R9C+RoHeGzFiSVnKcTB7ryMuq2UoJHZKy3qEnYalMz3uGtO/YT6j4j+/
fEJTM4z4QSplYXaB9OKEpazc4iFAFDmAbbOhcNBjstBeuJtGgYvveRc94PI5QWBn
XmvZouOB4hzoP758AAHOsLUzBniuZQYCmKr/j0an1fNKT7ndPvEynEh70App3klK
fj+UikUJG/o9WHRnGZHQ5fW1Ayons02wluInk6G9UW8kbFOW+vKMF/9NetJeStXs
vamynUK7+ffgPVDx99665lKzbtXGWnHFu5eWrB1MmQprl7AJCMv6Blfyk/Ng7vku
ckLCBew62zzdFOUW1f0Yohr4dKTJkevOQltUY+B2tC6jdZc8GD6ezjI74dnRI68k
JCGLLAOfcNvTXVLTSMofLCSqPQZVWcR7Y1Y1KFrsajGbCRVNtS0J38Z3Z0OjeM4q
SJjU0LDzzXa/oxOy0128AcakILF+aBP/fbjN0dj2NYWi/vedE4ua7dnVG3YeLHlh
2Pa+UiuoYxrAOp9CdzBzn9zcl33KMGb55wdrsHA4RsZ/HFnDM9RfkHoC22ioMWhR
sC/Si6cpCOHKkvlwbUX1x6I/tLflxvhReDY/l2g22S27JW0j2g+QWku1CHUp8kld
abNL6ztMGNpwl/piyunTZLcXOv9nqj+Q3+9/h2o+I530gbMU6qOJb4TXQh2hCWKK
FceokB0BrwJRStblKxAvYXO7KEFEhauYTpEaZN62uDTR3QtQK51Iz9EQ7U5OnHvi
L/uTljO7lJhb+pYm7UjDzrxz6pOp5A4wV4ihbZ1BMWd5cbHwU7pVyO3gPb3ZDjbq
gEapIji50fE0qVFJSUNTxPZSUQRip/WnXI+Xn86ntQaiJEWXQkcr8gUcRdyDExfv
LZym9VSsR8oTqbmS7eYzzabtETKv2NrPMlLm71IIfInYZxBMxDT/YOgcHNk2MM4r
f/J9TnwZ64Mh4DVX22O+QmCms1tJ3PNEgchUEuBxZRO/r29YIc9PecwlenrR6i+k
oe1xAH3w7MpfgzUC19jpEOWVdgCIXrst5e3I8HnVIac8SbhypNNUUCwe4N1MgmRu
58z0ZVpgMqWm9NBxbMNr/RfZ/5PZDEiVcMJJxIYtTkMNdv8w8F0k1f5SphWYIOZ3
bGaix7GKh6Wn8+iqFd1lZVCGBp+ig+PMPir8FggGSlbypfKoWItjv6hLd1hd/1sD
dyLSoZFncCydP+Uum9+O/d7+HkaK6p6bb9hHsfSJZSR5WqfIdw7nGnHSO6pLK6xv
d721E1DHrwOYNK44NCDCdHZIN+FtmUUKzJ4wGZmtcht9efdE9Ew+iwkowrQxZtWx
jUtbsMFoqepVrbSngTx9MoHUiI0mdj/rmn9XXJvoUFAvBOi2wfhM1bUC3dJX8ffj
OewN3AHJSWORyOA4byhn+xz7l7g8pzQxZhAKUIzOnSkEi+K70hu9NL8NsJKpS+wm
5bPg0BpNw+TLTrzZVBFid+CRJTGdB+yUaJCtkrWi/aOWHwWtE5/Q62W9WQlPbRdX
/16TwuuGbnXZPCFAZOBtCCS3wFzbb3Uu1lzVX1zXxWKA0schQYt8X1fRp5UKI/fw
qyw+EIgMPEl4HVG1RZiLP/wz1Tymt3km/CoCmz1trEKE+cJyy1mX8vaG9SDDCR0G
P0Rs/QKB1YritOhkdE/wGue90T8+aYaSEfQVKXGrYkNx5kH8Jv6e6Boy+l0BuBX2
GjvsoRs2c3p43bNp0B4sycCpzbJMPhHBcsG1yMWQVCoZzy+JtqZeJImBLxKS9Bcx
PGGArfKMtkw4PatB7avM2MbUiVif8xkzHJSq/ApMnr22+VcS84GgNBnk30IUsaMH
tnWuxAZnXFlX8PwcwSMoK3Qxi1LoslGQ79SONaaJ5TZRDSvHwVeYrLxopQ3/DXp3
uqKYF6SVGCUSDcrg53A87SG9kIzuviis5WMobJtIlUmGsWDdX9IX97acpGUdNdpI
BTVxeu2PZQ88YQr6KPw0nFQsS1LIkCSE8AAeNWEMpTCL+YhX+SaAk9X174eJlxA0
EmlQMJOMuZDepi3VzHjiSip9VhO46A2DcmcG1xinfvT6feTydh2HDstIEWwk34b1
/NU/KREPJl01Qk9sj/CiBzoBxYOTdBP2Gwk/3YPxiY38CjUvQdtZUKCImSHC6Opg
XmTZGi5J9YBPi90g8ikEH2cr83Ab6dFBJUFoq5zUCxDM/hf1nxWKcpoDpNFI22ss
HI81113b4eRYmYr+iAVxkvkR688bI12ug9EiOStFjsU062wq63kdTMci0bfTFlBa
izAAtfkgtUADcWKNho8FlHMJl8QBUirTNAujGKxTo1WrT69wpYIDpaQgsFbrw+Uk
gBvSfrgSHBJoxP60v0PfbTfhJhObFbfzQ/NAVv5zecD8vfnwkOPBONv0CN8dEOvv
batoJLn8j1J8LgL4IBTb5yCv9Z6ojxyiEr/wJ9EMyMVkNNgdLjnkySgOViESlZSn
s1ABEWUmsrZzCzircKZiv8wSLXBJQFzD1rcigw21gdAl6UpDyG3xNCF96wff2eqS
RSj4vgs3YurPaE5VuTzUrVLmv/2K2CAhsmHfl8Q9eYqPeGpo0/vzjv03jvJh2jHd
A9soxl44XmXWxh4k1mgnobwS0mk5gnzgYeQf3fmLJAv4sm/vXZ6d3m+tWhMIuxLX
Wa4x3nQb19gzwoyP9r+rjf1pijM204jtKVcXtFamQ98su1cUljpI2AcRh5aGXcft
1fGcfgymcroVIRLl/x0Gi86rBwhF12lv39xTfZd+dlp1lxhXbqkb0JGEiyzgUUD1
5wmloFRD0//IhRpQu+wzs+b4Z5lE607CAgxgRkKaakDcst3NNHegLI0xBdhgqPR+
yG9zTwfp3hf2bdyIZIBVfzYRqyua8pJf5XtuIM29T3Ko2w/CaXDMXKEzXRVWQ+fI
YHLqRotMTnEby2LOgEQtCLCf5eAASJlGbMF96SmsAXTYOVwIuu+aVYWMFanD16oO
7TW1hb2MLmoE4i4p/S64GRpp5WBCsb335iFhvbtenDKkj0tCfNoSSC7Cbng48eft
LWuEjgibOYQVMzMGLB2YtzXsDIEHZuRquelPewvWJzSirWnK6PLigE5avIqD4zgx
GO19n4zkLH3IceeRDCbo3z0abjNfGoUpq7Td7lqt5Q7V/1yktsKum2WJAueexcMg
YpOFKCa0XofBVIaz5U5+32ob54DKNNOImTml9RbA3s/CN7nyG+yqch13rJXAT1wE
EwMVsWvJLk63jXvK207+0WEcjsnXm9l9Tc5V25vFdpgUHS5FX1p8xA7QtryBjIe4
1UTTKInsSlzNCZgO+34+Pld6zCfICuYoNP+AcxpYC6CZLyrj+y42++Ta4c1YQFFe
S7A33yM9Bo1x1/6QWejekXB7gSzbkpyFj+5RpBzTZtz5QgpzerfpIPRjT5ECcxHt
AW3KecXoNGnpRD8wiVwxE2cKghaYsiQW+/vgXhdP3qj/tj7vYRCU1m1XZUVvy0rd
16vpHbL21vln0g2qxWkYaDIsCo5oqKRo1HB122ecapUH6DtrrCYO5Fjr3ngH+MOF
cqogHy2Qzek+cByY9wA1nGmxy1MXpkZbND73L2sIKXTuGdzAaAli/GJQ1oQ6XF6o
VKkUKF7vrANHgKNSVruPjwh+G0t2RhvYY7PMLvtH9O9LL+cWQAcLlZ9bwpXx2Zwf
e8cgzqUrJov8tG/QiwVIpolgWg9rXI9oAbDJ2iLqpbAtw+q2uc558grHx62IhQSx
9FJMglohXOgEEK8Q2m/C8G+3InfGt7YlO6tfZgXrwUA9TK7boMxNEXnGDhnxtznn
DrWyD8jfDlmtPsdc/MaDJ25mEZ6kRtJSWwHtRj4NvyfPR8Gu9IN2bqCLYYBb4hME
etvd0XpWQGiW6FATIWb84wxdwGD85nh8znqoOLBO0kn1Sc3egyDCpFBrO2L7FVyp
rLGJAYHcNB7euf85CJkc/q7uTI92Zjva7MvDgbbpt1T/xTMamextkJCyWK1JrVTX
XWVq8nmEyf51nbc5u0AHSWheSoxLHH9lPdOMoiWLKDuwi3I6wl1gvYtEb2nnoaHx
Yu/eqK1ByMDnManbfXUDM1jVM99jfO85BYPtPYELiFFlbBHfn7uFEUxBm4mS9rxs
T/QtFgtUOv4Idd4dE6EeN/yqftzsmHH5yx9dD6QoaZ7c5tgcptZ9ayTPjOvAAqJ4
swnpuB8RyVxDRP16LbERgOzpSA/oEATNjG+OBt0pwBW+IVTBw5Al5i3HMnG2iPB9
bWl113pOl4wVzPeTzAvYSkHUyC/4kmtlS6/suG6lg0VpSlY2ZkzRT1lcG920Hcdl
zDHPRidI/j7hmnxudqCrEnz0dm3y03NuuiKKyYiozhGyap4PUNQt3fMdYfLa8YfT
TeLlQy7CFuHlZLGND1ON4TSC7gJxIIfV0vpra3eBZtMP97D4otixUOgRAxuKQC+O
dtICXDwG1BU6ltNaoYekJ6y6g5w8vrM9a2Tu27kQ7hTdxEBsHoDyP0G7hupoyBva
5jQWhw+XAjJowTRIskVC8tvmxf+9ZnSBtt5t+5TUm76ja2Z1uTw8NnarcZZQj7yT
JTAABh4x/QkVbVw7ULeBYNTXX5UfO6ilrrMXk+G0nB55betmSBPkpSTiHXLb8LJa
RDP/IYqiVHONr411acAckCQ2QZc4raT47+9SoUeFA6CnAMkEJ+1ocQeTuux8i4om
SMfHTWg6/yoTke02Fv/ZIz54QYhdrKfYxKFV8/KP4lZ1lFmhR0tO9WRhEXybuUbp
DtMZAMisbNdAzbnMIlbzPTASHPjAeX+XCUvVaBAZsigOIqyxsDkczQxAaG9WNVoM
2jiUMVUXJTGxweEEmNcBww4kPZeZnaPmU+etDMu2EcVv+l+GUuslMxwd6loGFo0i
e6RN3byamomC/J+v+D5cAJgmV/juq7YaOKBPfcd6oqJOIMD8OPbD8q5zx/9e8L4Y
ji2z/Cc1j4TbRHDH6GIZS4jEJ+cFFeBL2oEjZEluxpMJrE7/knqTWqpGQHNfeZVB
WaLxZEZL066T4npNRp/PbY5PlgODsPeaHi3/6t4smdQ3hOIpCOOR7ck9zeJ+9ubc
mh+cz07CTQLwuAp67TcGLY5e+mvfIe8pnF4uAR+fesVvcJtg3Wpsoa81vZ5Q+EcB
kY8CmwB/OIGEUtf5ee3OGTeDLsf34OQXHqSSm4AwgK+xugp2kYxvjL55YrBzbT1j
tl1y4WOxFzI6jh0TcUqLWoI1HQCcu6yxyUVqcpzQNBquKvT4TkEwwi0L2tcM/bdG
Xc7n+NfPshPj5MWjlTH/F1RZFTICc8eS+3pQkPGkSWGBWwqzDVZ6FGP4GQ5OCV88
lmZvIzPreE553QXDO/kB+eRsHh/zuIY5MtgeN3FbbmW9EVXDYWy4zpAkmXQ6I4WX
`protect END_PROTECTED
