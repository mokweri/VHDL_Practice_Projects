`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7TLa/O+pajFlZNt8dHucdfGxgc/usEpxgbOcXJSoCqE3BBOnkmvTfVKU09rD+e7
DhFPlzBvfvTVVGxbb8skdB/6qQ0qdKF4iyFVsikCeNRXqedRg/nLTQ/xgtBHgUys
Y3DedM5B8C8Efjprd0wWLeA7DB7V9qjl5l0Q2ddkPQUFBxrp9Ukc4gtr+rv5OfAi
irr7eKNYh5nX4iwUvfQKZ542QuX8ZNwroj5H6vCe2GIPjJmrgZelmu5CIrlPh8sn
ypkwmsUR7D05zZ0V8ad5XZbMZWb7O0XOVij4pI9g/dcrb4scRihjuR5rroTAqjVw
i4ot+W8++HI8+jJ+KzL46Atb67rATDBft2KEpScQXgLhwnIVibM5JHK82rzUkBro
gROm3H6L0DSVhRAe68HnnwD5lp2uOuJVsv6fUmOHzznDAbZwo0IGHtB3l38djMCS
MQOkoEevxFf3wF9lvIAB0G8VyeW4e8FhV9FH1oQpmlran0Y3Z8vE/23hyLWRXLEO
iWzyfh2Iu3bd2PywHpfKPSRWmJiyKCdsudliwE5mka8DvM/TeHOSivprx+8Y12jj
QSqynctdolJh7A5vPbLxF1i2UlOglUeU0ORzML1TUuPZWdE5bXHDAOzyWbwczjJt
3T33o8slj18+zyv6JD6BS3H4d5xh/colCmJYw0pNfzpXwqhNmKpi9W8Q50fWOU3i
9MCOwHM9im4k0VTqi+nrUxZ16y4bTT2kR6EvB300WGWjrjOFb++vWNgLlFAA/xP/
o2eBj6qPgWeDFTgNzTlQp5ffwOOUDQCIHsq9wfoE07fXdXIM66vOoMxy3hlzQr1o
F3/9FZ3PGyY/hiXwISKE530gU15nqag8tfHXh4FbX0Sip4KaBptcz78fYeTwiLhX
`protect END_PROTECTED
