`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/XBkRnx6i4HDULTGvUE2EHZjBCtRqFl8m2jEJhlpDzky4FrdOWSLixzo8DudMva
fRoPnelRVwjuOQzbpQiiNgL27zEoMhpuQxD3mXkfCKHHUsBIzaJ+bgH3qqYfzc9e
UXYOB2ATQB9qDwya+EAsxQHo5CGwZQ0IBScy610CN3DlUFe+n2cOachsBZLg7aqJ
Xu81BTHDhoPwF7l/kccFVBqK2oPPwKPkBP5ckwZAd0K3+GxccYebmYDuPlldl3Q3
MUngiIoPWwizPSfGxIAuVqyvoxfX7CdCdvmVoziMGPaiqmmVND8dSXZFG9jSYE9/
0uF/iJSL9QIu7wTfAYsMS6VlGb9j1bidkfudJGrnl8m1Zn/lCqO27IoLIkBBqOrh
P1bVsl6/+TDIYvXn43A2te1ryLKo5VcP6osygQbtnmN0tokS7pAqEKyTqzToOSL1
Mk9GKvVAXjv2wXh3rQl79hdpCWE3uPYsGG8pJMSzxiLazB2SdiGy+Q6ea9cjGCPm
ePdAeP2vj+jFxKXtz1mJwS4TxCkfiNEaDLRkIm+Txq7u0H9KXCFs39mPPOjtLCl+
znsteH9W29Vxc696e0b0eZ2Aay8JHPiUCcCeQJYEcTBBksOFaG2bZL320gtVG2Zt
f4f3c6pYCmzw6Y3DcNa0xX5DbM/lEGerlcpYgovq5OonmcrdL4Lpu+xShXtDyDv6
LPsiN4m/UAZ1xDA1QCK7LZSA9FyKi6fRTrjJm2NY2EvNIv4q8nY4jLEKfgH6xkh+
k6KDZTzXn05hm+EJrho1Nr1IPpWFosaKMfcu1+abLbUozWb2A67KkkJlv2uyPUAk
AnsK6nHkrw9/Upc8CQBhvxZM/P2xJRdsRvcGE8E0le8FiJDATc9Kw4+JVM/+zjMU
ASQq17Pp9TgTQ+V55T1O3azxSOXTcu9OJcT9bh36WbqxC+HJwMH662+VgX+Vvj2U
0hvt0PpUD9pOX8IKfUhCow9BbwqxNQqtjW79FELSYPOCr5LYM5qsF3fJFpobYK+n
bpB3Gsm1nfur479GlCxB2/NIu1gAWbapFqdiAMvg7iD63CG7JtrgivYz4Zhldkw/
RE2Pn26VFEG7z/rRKEc0IHpg+e0X9pOCX14qSzmW7ad5ZuCuZp0dkZj2RuTjxVsz
SzucyiZg+Si63xdlbCa9r4W9ZW5NNCjeDM5OxFK+BtwhOaAixFm9ZJXXhIufLfMT
zSCx9hXtT6xLGu1VeH0BvW6mNzdmbZsrr2dPd0Z3dIqHjJIjzegBBM1WKyBsrU7l
oSCux1saMFMSISEJtQwKc2k6J2Hk2XAtAVzqz1eSuBveZTA25MMOgWpaNFxRkTS5
vm73Kduf5mzonuNCkgD4yaa6T7aWx01Yiokq+ZxDjvF+dKVPm+lYmwLaQfWnhG0N
o+Vwoi9snMGq2FuI+4QZ58P6w1OBH+56drsBAt/MyEBfAspn6pTlh5Qofo+piIX7
XkMw86cr4cxG4aOiBpuSEQEII0RUGpYxwDSpPJhJtfkdx+6iccoZpy110pwnyBGI
5u6kFWyltCskbeH80YMhb+GfwApqgtWVYDbh88dATJlkPK5MkXaQhUBnyfFqPwfm
0rz1Ow3nOehYj+7NCwVhf2Men1W4VcqtrbfSXVHuDPpOEo5k9s9ZWRWgvztua6Ht
wonCeIpTPj72FnBVZF8kYlYXZAdL9ddJmN/CAm468gbyNmcd/ATN9nPgilqbnDsf
oRVMns1J9sR7Fp5ux2o9sivAbQSDP6yW2/WwoVF66rQ/tgEi9ZA7F//qvCshE96G
GrZvDO/Li14QOb/ZJ/oVfP3PxCT15qkBJwp/2uqmmzaQaCVxAJvjeR1b47Wsg49J
q8Jjz2zlVgWeerBFGxONwmjwpB7HYxZYNqVm8N1panFNraWNqDwf8PNVTkDrhNmv
paraot9TqIbFmvpelqRF1xHQuJoQfIjofRfEGVzg8YTNI02TyiNnz+vFa0YS0p3F
BXa50Zn7tSFA6GJfAx41bcsP0m3qxF2gKedg3qaXmTP3BFuxHRXG5dotzGiJfbV8
0DOY/AYNn80QzuWyNoR0hjrVdARPuOkb8nSqXwhglIR6b/+I2mwgux0G7DQeWCtR
YqGckpHaN3m2MRW3TYjqYfjVqzTqf3U5WvPYEgMd2fK0dbczenIFxxDVemm/nkV0
6MBguHIuS0GuAkbZNyg77cM7ojHYUPa8xkEIp/Cdb8B3DmHEKJ0Va4wheFfEoIvo
07UWdeOEaFidA6uRCA4ezDq2xLbUomw8s/jb0BUp/FNLvnDOQxEEkIvHzNR/kOCo
nPcm9QAKMd3B/3ka2kA57Yk82CvgLspsOjPtb3vJGBVTIsqeEPpAgBawPiJ/hV4q
5Z8j2QA4hDTNVxsrHnVNLM4MhJ5URrtVQkGlYPrK+mjcw4siUo7oCuS7AYaiIvrF
0LEYzF75I4XXdhnd+2qX7VulGtgWSb3GATKIP/ZBmi4lfBd9T3PiPIQU7bEykUP1
iV/8mzWpkEihhbwQ1/lXTX0rIjEHvxV/SUksy+3FBz9aecFKLd9QlYbl8pWZSngc
9Zai2/B0BOqDYnSNskTzL+4+kLzYOiZQeE5DKaDBkreh0O3N5MvEm5ZddYA1d2CP
a5qQjyV4pOtMpeamUp6JBf8mJ2w56nt/KknzE7sOTV4ybMpSE1+52WhfQ4UCxlSY
YTc+1iSvBPw4+mLxwxGfH3nx+3LO2gEyXib7lGEAPwV7P7ld4nGubueVjYVcSdPs
cev4xZfPlHvY3ZcCVH14EOmnwUfT1CbZewlS4fDEFJUFY6KEfFVA1yttg6ilpazZ
Uhjs9BhzBsL+jiSC4imPntglFLJwRkT6Dqf7WI2GyBTaRF+OEpkGnu2tptgmhcLZ
dyx4weg9UNN9bqajpbFKs74ni7QLhwzDOQhB0P+zfbIaeJt22HkzlkKDeOZK61Lm
49k5TnlP+Sj+vfAXbCav3GgTNTwJjdXfX2qxS3F4SY4vKCulecmdux1SvRU2JB7v
CRNK2Em+KUNg4gMgVuB9/SGr5EvBBwpa6WMQQawmn1pZXnNmYQdZG7OHoSM0nwTx
oVt/r5q3h8RaTKjd3/cw+qn9ir3y0gXGqfTZ8ZWIrPZcfBNL7ZZh2BT6XTh3NcPW
xhZhr3spXFUZk5YrRv+bGOa1qWS6ZH0spypB1UlwOOd4sCNbsO76V8TMn+wrs3HL
v1NWZba1wHJcdTd4ft5tialzG8JK1S1uYiOfeQLRQHyLowaWhmw9X9XOrzParswP
fWSFxo1jXhy2ivacRfa2cYrHWH2iJp2f+ciM8qtoh/XwDeteL9TdsLUjQl3Su5ZQ
7Z3DCV1YmTSAsbRIyIzITXHOWLboMsZUe5wOR6yVXL3HlvWaWr5UFVPOrjzSmAPX
beUY56L9q3nWD2ttjTsgRjXImUbRiZH/Piu80dGYaK7D1P0RCXPgKcalfTVfVeUI
CJq75yiU3An1ANPdhpzVL15/aDdCpzhhgwHddxiVaY/Pa7Tq2ABBnOmfg7UitTLt
qs6fkJb1T0P2YRWezUljKTs2b+CYJRzY/108xQRAg6hWWq7Nv8fBOa8+n0uKVsci
mJce59/L9nSIcm2Vb9zaLQ5olit2wdjsVzrNMYkQcqK/DUb06b5vhNw0lcNNliGa
I+Ml9FNgTAS9GSItLBZ/6Sx60Hd63shHTu8AlJ7cQ2ZWIcdYrOUr7Pau9eyMoEOY
B93QjtD6i5I1yEsXvXsUURTtC0Bln4dKNkvibYDmtepzyI3h/fa0n4+HzK2ILS9J
8/IEJiZhELE4vzKBM4PIwHo8/015FvcwvIo9NGIjiUb9t35tXvu+W1Nt83DMfljb
hIG6bvdvJiWQNKvxVI2eP2RaRV7b4QbjRIGoKZPDyeeaUXPdgFCSMqCSMmciBcxW
sw0dhqv0LCdk+dRvxnXA5yY7IRbwiWk4SoTtNIz5B16aNGfQ57TbpHaxJWpLpm4i
nMVCoDMTuW6rfmFUDXBYllmeOZ7U7vKdiT5khPD/N2VV5f+DcsoGWgwAfFYUzkDA
E2nh3xVH2HcFgLr6Hb5VF9nnp4JsLSLwqxqwezKqgezsw+UP1Aj1B8/4ku4hoOMG
o4TkJinKst2EmxQ1OqRdQKpBSNxyD7VysIZZjomAW+h/sj1Ph3CKkNaDrYhi97UF
1hfkHHvOBFCM1R93Phi/ohLV2yZXibtw11tqYavWr35e/noO0ZgYk5m/fKveoll4
HMAUWWrXwyDpW0JNvvDZ99oEy93PLGCDc0qYN4JbuDfkv0/TUbfvv2iriXBw9wWd
Fg4OvMIQWVPOjNXChbyDbiAZhWJhtCsEuTanWRGF78YJxEvHCT8dIYQWERvUisV2
SWmEZQUWSuYnm7FPzykoCfFLsRo00kPPCC6SAI/oSQsZBAlb0rM5n4wPTHzWzTrA
bPdRFaw1wZh5acGF0qSgDjOYauMF0foUnZLPG7AFFzRBq7UldcoxbV4X3EqnWus6
pLCbqscdVNBpCRyYMP5x+aXhGJQC6tkdftJYTGY6CnXyWzvCyO5wheUm5XMyFvmC
DJZVYIAW3+E1y/RLSprfSktzaxYH/Y2cz0hocMy3TfipvqvanMEF8pjqf9+Xs6MO
qSrwTjAhtTUtZNUXvLnf2xMj4k9uIo4ajXrCJ1OLBNvC3HLOyRajTzodEhlbV/Xu
XSv8e4g5dZ8tcavHL7vpElWO7IMwQH05XHg3qU8Er48fqV1OT4updgk0Z1jaxbNB
b+0Z+zXVeiDsJ2yXDOtj7OG542ef2ELjrdz+PrtpNsJ61SCGS+dF3DBudDklcbD2
4MjXqwmikVFRbfbJ3XFFBE+mUDJGvYeR8nCfwwZ3EVOTYniPUIuFnu/hRvEG6wjl
Gw8xhnbAqm34bqlyv6QBESjUaX5ss+ovzOcUAnGiyznZLJDkhL6BRfySwTnsiBXo
DXh4IhTzLRmbe5t9Ktgjxv5hYXzWmY1R6ZJOzcoLMLFHwhjMrbAxPWgTxe6vlF+U
9Lbs6mSbeg1uFBSAZ63K4wr/iCFbR9oHvb/6izqCJW3XAzhKCcRGmibOHCE5r5Th
28l1wzzpT44cQAzhjhHGvNKgp1AZtK/fA+RXHPrHYXGzZmaVBJRH2v0wPZaSgFGD
UTR4eKnRj74fcTmDe0a8MWNPrlid1rahBNtcKH4AJ0werBhAk7y1mjjTqr90Oojk
LIhnh6Y8JuvD18ctQoVVs7zf3q5CUnQRn7GIE3ZyGDYys6lrlOu/d7LS2yEF5ndt
x7j6FUY1fDVnpb7wfzynI/iFDfjnjHymuAdGAFKS78mz1/KhXmXzpvG9YR0jYCYz
GgnNI89QHMWpYAncWlMVgi0BMzqkIyjWQemXyUh8rtSwPnkl0Os6AmDiGnB6Hi0C
Zyvq1EcsiBtwPgj3WXa0/KPsLmJXBixnPU4GcgzuS8Nw2XctukmhfIjWC15aU99G
4cikVf+fWO15ULMPA23URRwA9d53c/LF2/pIvLAbj/E0/VN1X5NIAuCb85VvpiY0
thKzuJdF8UXS3OLP8hqk2Cik79Cu7fBUCpBMtQppsPOVwJXn2RIEC+4z8zdp/N2/
mU19nxZTksIFKgUtbaMnOabRpHcxK/cnx82omYevrzvLSStP2jnRrqyn71A9djrQ
6QLqQycUszN7u7K2uwS82rm5eC57fvjrO91IZAUFvv8nBV19o/3D4WJMqt9bylzs
S+ZT6UuMOsHKSrBLcj5nsYV8D/WVC4urANpEx9JEKREpqeThKF/FrcPUdHl1XDTw
0oGuwXoZzqKZc8NkaTxC7HNAYYQAgT7zQzAUcMK7svJp+0lea4LTRSiUMLZAR0UN
0bcCWUHLA+mROnGEU6ZJ7PQDatgtoNPRJ2k+7Qo0LKICwgCqa3JKnjXhJp9oiQ3f
ya3CrsS1eYzlEUrbM2OyGcAoEj1TnITQ/MgI+eIyzYU8i+7d6wooaJGcXjGrNb9x
8881dSbdvMzRWbFfmzfAnmmWmXRmOvPb2nOezEappMZgS3uZS90LsmHTK1fCaStP
DEBaCkPILzYU7u7I2tjhVg5Rkj73Q+0IzV0Xjte3mmpfJGP/zL+0hXN+MS9473oO
R0RLFEDul3Le15f+xOab3w37lUwpIUL8/j8H5TpxLgIhGXMcfLUdAao2aJeCm9JT
ynD2cchPSXf3ayVOuZe4xHu0qSZHqr8T+ZLx8dTDQF0/NXGuzXBxcd5jgDiLAMC3
xbkUY7aAubLSLyMenUiStpKGR8A6kJ3KoQdY/bB8iwOajMSNjVBHA0oa7PodCrDW
Huc4fXpsQrssjpi0A/b4bLySCNqMUwkDh1vdn4MbXuKUhkvsjZf9w8Dp5d3FlDn+
nZWdYlmRXCapcH5+RwyaiJrg9ucshsKyoY2E7RM5lEhvQXgOpgNN/xP4vsdXIlOn
nforc+4/7V4pznpCtAHOh6WVG8Lurgn7GQaGrVytIKyaLQnaaxmkyj9hWB3c3Dyi
+x96pIP6HdRCGChgmVDKWt7z2wHhndwMXy5o5qgf2EEveJof/6YtQlt9zsAB11Zf
H0WZOnfOfHeGSd7y4bAPSCn0z5aYXbA2IVsN/d6WaRrIPzFy5SPIAEgG/cOenRQb
dvFOCqCwVeCTZXBXUZTge/uQCvb6LVQYSBwLpeo7Sd/Se5ER78AuGA9TK9h9mjia
de5y2ry6uOLzn3JcRUgPBDGwOTbEuEGmvVKFLC4B+pI9sEYaMQimJGY6eqQND89t
y1vCZtfzygcIekZ0+0ssniineNDEXlfadAMJiUFQublbGU8LJBE5UX3DeFXLJFvb
Fob85V66w1nd0QXHQHuhnXaPQoLa9xWkorD7SyOKKZqxyqcweaRjOmRNG1g77wph
TepzY3UoF6aj3BOOCGinl1+jlWGnU6gXEy8f260JVTCHpwaxp8ZEn6cP/PQdKW+v
rr/GwMSDO0zxMg1l+cdEQtRs5xODf6Y0gFy6s6GfbXSdMCr5c4ZSzzCv+IEmkT8f
cGO5p01we+Cmkp+xviZtfAd4j40AJHFyQTWWliqYH9Rp5MEASpV5z1fgk8M24arm
4n10ohOOO4AlYmGRCtqHG7TFVvsiPLb7VpGy644NGl3g2TeSij6mHHAVy7jcf08d
RHgzutONIlQSwm99q9d3DptwnkeEoF4I1YvxuEOTFvVNFseTdhpg01+WCzlxs6RV
uEwxDiz0H8TbqszdYHLPM1C+Rav3hV4ORXhj3zrl22bTVqhJSHnuuWyTJXEX+ZvH
EJiobIRH7sGu1vZYAj1WWPssxnfu+s8qTCWtJ2dzEOnwCKFBXTJQ7PC5tdIua4Hq
k6B/lku1D0e9RlQr/pFbluxODQ0xAqTOHISda98sJdlxGxrakcSnQ3WwMR5bvR21
s57aTTG0C+SSsn0JK6nEqScYlcKIezuf7kCI87uxtNUWlH2hKmD3MtDeJVWR3gKg
pviuFBhukFCmViS793LeU5iX4WNdRMd2tKpJC3KMgEoMXXpBwmH1CR458Px7uRZU
5ZuzJYpD9f7+s9AFNzS1/RL9JctY17jPEQuBNopDsdqtuuUzj9Z3HiwNrvgaVRjq
2XEKmCqqUcx05KgCns0KE6YRfqAn7DzIlqKj7MY2/MOXxtjl6R068S6a4rBPQWua
KmbjHCQb1s1+8qt3cWHu6xRy8peJNIfZ2U+hy3VKGHPXmeJvpBJAfXGdG+uEwvFH
f5kP7S9ED0WvXyFzJno6GErRGo36C95kZrOMVjl7FMsM1YPt/mmf4xpslXomXYhg
3yk+kebY/YhmjNcHcLJUUCXJngtxU0ixXfJUtxrJ1OvjbTzhaY1fcouosTiemcXp
PaF8DwnlQZ0mtuUFN1nU1vDojhdn0FaudvUueaHq4tY6874eyFtq+tDwPkrgzoD1
jlDdfyufw32MDQi85QUBpHdWCyl/3+t1wbhVgnegRMqJYtjsumfLrb1CW2YuCJAz
oktCoqA2c7tk7iTBGpTzaO9YC1ViyyhT/5UfmIhUY4P+3wlJz/jPurpNreernMjY
WxiLTjyZzzBfKlU0gkX5QGTTGYj9FpV33/LWo1LIFnec0t6nBIiB9azsFgnmp7BH
btOq4FZRLJm+tqkHuDseaf56ardi6pj03IWhM99bBbUf6fSf2VRAlr4cMfV+5Z2C
QDdVLC9gMRx6gxhvYYZJFIdSLg5BH7YG9yNxcI3w1UnqO+p3XcanU4HKgKMhverh
hqCrAp1JP2FQHbB23f5PSnojXc33mqcBI/4lCLk/+HNMIgYeG3edW+VYpuIiogcA
AbhgWajcQQvv1vgfrGZUSoOKj6i4uTNCO7QoMVDfWkuf0Wn3+EasgfPB6dqpeeu4
Kdl94c9f0OJk2wkxvUPh52EsfdExvFRlrb258sRBPfO8+/cysT4Jaew+si7CBMHz
7VXWkckXIUmGU0+R1XqHZ5ymDn3XEex+kb2NBFDhqUXYIbYHBYIiatXefIuYjyHV
Ok4EG7u/qC4CwJ2os8Eooe3gNEnh6NuZwUKw4ZUN9BVywEXP5m1t193L5+yI8M0b
YxuwEsrbUfHbH3roUMAros9aE3R756VI7iPDxlmOz0KpC5cbMgC1dJWG9MBFeGi3
IKY10WE9obA58XgzLpmEewSjwfmWCWvYAMXVp6mmv4t+My03INO3IDKQtKKz4QWE
BrYLTE0RVMlfWayRLuMFAWhiN5DsSPMkIYPAv6hNmKwFZfPBFa7FnEN9Q7gUSumU
U+TwEsMNZdE0b23VNVMUZOubXQTtH6EkPNu/z6t9028X2pmXNevds0yjh9oMx6sr
PM9pfhppvowVr6HR4SxgkidLbaKKg+5GZRSVXJInKC9xKL/0L3P9AbAyFxr7rLWJ
9j31K600IR6N1HJJh8aszMD7lWEoJSt1x+InNzlBAN0LS3ewYjvCKyjs7j5/unTV
FmggnDuiyUEBfqqbUG8kguzFgpMDuwYnvuoOvrfHP97rlB+X4FzTd/VjVnJ9lg1S
mWSCY8MUJMQ0bQ/jXpX5hYuT/L9+r/nIyNiEsFupII8kSb9S+wsuDNYugwZtZqKb
2OwuzmKAqbfCJ3xZ92UGe8D5+p/p1yWQIuhDPXu1veZpt3vv8aDh9SFp7AgFAfD1
S6PQz1LT7OtckkYvLJAFqAqvVKTGj0xUr9SRq3z1b3YqR4VnC/5/l7lhh7Nc00x5
arTVm2TqGbbY47clEjxw6Xmqr9ZjnyP+px095agL2UpsuJLZ3sqCc1zpSH3/PiuN
DAzarY8NsCpnYv0aVc4g14WMNfuoOrip4iBtovAZaC31GxWpSG9DlMbhiOJ90XFv
7QQ+ToPT3fSs/jVbLx/cxbA5GltG3rY65wwEm3ewSvaSaiZ4eTykI7SHrAeIVR/F
Czv+5jdyzRyLlY+zUKhW6EpMrghJ+UQA+hPE495MRR9WzklcwJBq54d2r0/uPgjf
`protect END_PROTECTED
