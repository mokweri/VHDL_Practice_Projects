`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdHi+Oxlww8px5dZf8cpX1oHvakre6RSYoNOoDUsx3DVrALrsvjgYtG0N25LcvNe
TH2yA4CPXhmxHnDqLDgMTxga4wQSGipWr5ZzuSMKI6AfdkVnLaOol8glsNmTPT8q
b9OKOA9hGI+BnduP/ovioSRdjxzLvJeApQcsMRHkV2rRnTXWLq3rdKRTt6MhDB0L
tONak4PeCJh8M4dfhR38kK5nPne5wjOZZNBquyFLvdwuWk2i68hMb8DONVZ84qhp
Ikksxh5I8Geb8Deu7FDbEpbMR+1Vmz3ZqPOwsqAMN1mhmA7VOnbasPJSuBzECQXg
TSDXodCVB9+2ARduL87QqYPBMs/QjEgqCjwMxkjcJjXQCWMmryfzCB2xhUjWNGaC
EPe0tjEfywxuYYvrnfWAxY7X6oF3H5XXanNapg1C6F5UbyO/cmyuI2AlKUhyZC1L
GWm2H9Hy2gfQbuyPJdIizU5sVioo4SE/jv+hPrGgzoIxyWjK5gBLT6kHmPPPXfQY
OdcH5Z4gZTMlZZs4qAHtP3p5KxVmpFnJgctXGNuIYd+Ko7ehhkrx0hyrbpRcXygV
GWLyTMkTphLXwz9LSED6vm64PDr29pnKpohC1aZj1wmEBVePdJGgxpv0YIG8rVjn
PbGjrwRnVagx9iNeq9Z97kGTK7W6IAgscROuktQl+9OlOwibnEPBQopeVJzaDc3s
1PJnYn++Uqre2R3mvwDuTpf1Mxd0CwE6TA9L8iLF2a8Qm01sjzYhDzVeQN86zfba
QLv1zlDkMHq5XgT9jKwXy8JwSwihJCP3ebY59YzkE8r2DVymvschL12SSyBlk4Vr
EoiFtAS5C9rrfIsJWK2yEi/kU/mwFLCx6DTh5YGNTa5gIAoe+BU5f6gJHgoqYm9g
6cy7aZEw3JCCIVbZCp/TwYf16lAG/fwvJI3JNM1J1Qy7+zIQYhMciH3/rWatdzYB
4aIxbDcwK2gmB+oZJT9at54u0aXUPUFU76XOInUovs1oRSWzXOLufG4g5EYYH9cH
cMFI0NaEK+50LVq12/plJJfhUYzViclVRK1f8oVO5oe/u3vhg/RR56RnblfA3ZiV
4OsqtkoYQe5/h07bnzXXkhBrYoijBfgxeoBm2NtiA8LMYHzdhzuM67G6FkD1nOxg
/Kl5LDGeaeESg9rztMryOASUFzh6SY+JIRPfmdGamzSwRpPGP2AqO5K0BSVHl3db
mRg3Tw7ik1ZtSHanOP4hZgonPJAL4WR5YWV6YuhdfCvzc+5fby1x6r63J887piPv
XbbG0XJoh6930my1h+dt70qV2Ap9iHDjbHdAdGMmhlAUzMIGyH3oOUWPSXSDP/il
NDbXYyn6TJ8JAYWxRyDXMUvlAIimeAleuOVdkjl4G43bidBXIgrcjWL6nwfJnUWu
LU47bSLebM4d3R6o8IT6Ww==
`protect END_PROTECTED
