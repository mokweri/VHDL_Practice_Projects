`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZqR+gW5hexc233xAx0Mq6TaXSZg2/ztD0dbjj6vDFkNthBHcEXyhmUkodgA3YC6
yt8pwvdILJU/Bc1LafIUlHUw8fGsaX8JMILoWyb0NZ+gndTSFgbPirsB1aWyHrgp
Xrp+IVrTyRumN2zFXNIWF/twIUaDWv623MmCyPUmEneONjsFWlaH161Z40je3M+o
45pO7fEK4mz0LeWNHzrZ0SCLUcSRSurIBIk/HUO1jKthy85pd175aGKMdAKzbUrp
RnntOuPlpzP6i71FJWMoDgBmgOVPdabKQUgjDB6Ie+OfPq5+wi4eGpoqMY8xqyTb
QJuft/pSSwzp+uo6a3X8rOWpBmzv/3EiOy5eFkvaAgIFScUE3cIpJxPPJb486E6u
7B72nVxv456IgHrTDEIc/nJttkPoTiJ8DaD4WiD9qmf2QYIk0HTv1aFOme07Qv9Z
z09Jhb4i8+QUcdP4Og2z7sGOZrP1NUKkYmDSkVZI/Spk7m5d+qOeMxEOmXw24IC9
SLSHYMEgBc+qlZBQNrruk8G3mCk6AETngfx0P8uBOZsxAUFN4GMs16/Fyofd+E1w
Ah3RTnuApu2bKukTUtdmEGwDCu0OH9NVjhFpjUYvSucT9kxE2qutbFIwvuM3J6Wt
6cxyVGVl033iP8AGcQtN3Rr1emazeyT1TL9Wtrp0swVSc8NNdMHfzwi2wWBC79oS
0N+1dzN1cnfe8q2kxYVo7FNXvZ467HhDuq1sPxUBXtmgi0uMHTLM+pr4tjQHke5l
Jg5GfnSSXSgBFY6wzxUu2Lxk8oZrEGONE4d06vpujg3Klw8ZEMklp3NAbk49F0zs
`protect END_PROTECTED
