`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LQv3rNz7WrghjQc5xH0JGHoMwcwb14Yuq5KLVwV/3IzdqesaJCOHoxx3iUVpzBQs
RvRoUUnVjUXz2uHSnDHMtBFNBny/ay010gf8lNpELGDlFFNk5bSOc+ELngPVVqyH
SAs4qNNVPmPtLsGDd5mvYjNCUX8+54oK8lIvRHIRerabSL/y+xM0P7olcfEKvVb2
+L11eQtoPVem//nla5f69oFAZX/CO3FpCQR73IM21GjmmI/e5k3hyRhwhnJ6xywo
fXgLd6Ngg6VrWBUrpNVoMNPOPHDwq3kKxSYc7qvx76G85YE7e3Un2kKVhMKiW4jE
4L0YCw8UAEQsFuO5oIHQR0NQen/vkwXgN6MkEmTYK435aqmxSsEXeUN6xvrk6xza
iPGT+pFVI8VQ+k4Jn3DD5cWiP66x7vQOvssekMlaJWqaejQWc3eFdHCyO2E8v0Fw
mAKnhsgR4YjAihvy4rJxecM0AD+IdfJst/3L4RU6hGRT37hr6Clsj7353mG37UB/
aOym8FRk4StPax5Aj2v/H+874v123cj79W1tiR9q3vXC6D+GqsaBPWCGjiwGNlVl
AgQBSX1il2660pNuqyyuq2NEbafq/lsKoIxSL5V3EPKWKR4Bj5wTz2VmWwSaOpi9
0kWa34N7xpWs/69KXHgXwzjSmeEQRzghXvPOGxcx64eEoSvTy6yC2SFgTRHQHJcu
0IzCn4D9FIpB/e00Bjy25QKwKpOWoZYaBeNkE9P4Qda9KcC9ZiqGpyYP50Uogmr0
oZFDGreToIKRcNrDVVTIgUXcsfJtLQvGlWvO5qqeyvqn/v6y4S0UCt9XYHRBDowC
GTMZNbs8mxYfN9PE4lJwNUAMu92QN/FrIg4t0HQr557EEz5hOlP+qQDbUeBNuShc
EXV0wi6mAUDhHuicXhsMAV9O4zKOtMt9qgLSsRGmSNSp6My6UIbz6dauFStDqbEU
O/5iCzXV6tHozJXAHdefbyC3Sm68Z81EyNvV2By67aTrsBmdAOJBp1TkJKsp1FgC
MRn2LsBUWqSios60uwEkO29SDxetROOe1PYiJneoUANCWFQzayjcd28yrdYPo7iH
37a4dgGMWQ7mVB9M3V0WnW2DLsynP++10XY5gvAOoF9AlVKFY5dTkOD4goLtJRBz
9Pe19sem24XVdkMmBDAbqkltd6NizPBWSZ+G510vI8IU41oh8hhc52saWlBDyU1+
gij/tQ4/K4oWL78YpfP4K3Tj3vvQIjTOmfiFOtQfu4arPz2Zn7mReZsrojdFjRRF
zbrbtEuhadBK91Po2wLx5xbs4bCbU5fMvo/1aSslZOImjP+h7hxRPxg24hW7qo2k
VoD5cbI2muscb0KRqx/UjjmFvO/dRGJi3UBiBmjLc5TOipKMb8qmW/7KgvaxPPlS
WnQYmUsePRdGmrGEsj4po26rBSyNQCDKpesC8FXS7MTUQNScKJGhMEuYDnxqLwoI
JQ+IXcDi2pw4vbJHCUHLgAxwQ7aweN4lK7VY1BW8LwzHxwlgco/Se8aNs+1UOJ/j
cLl2/ioiPK38AXQTBbw8bvJFVqN8TSpUt8zovvZXeOHbMtBJUQ/Y2zdFzK5c+GIz
CbJkBgW7KvzC7VB5BkSxB18nHadxY156IaLluF+KzsiLs7YkqTrajGlb6L9mHZXR
ubtSt1xiTqmp0fZ7IjKXD4OOTE1yk/DCGhpXSNRjR0W0IhUN5+m2CkcT91VoYqrK
4888ZJCBGF3F9ubO4lcJeGwKwkylKQ4hh1ng3dPoMy5OuL0UQVRtTu4ir+CS9kM6
KS3Szsc3P29FqALo94Nym31rqWWuJRCExBElXFMsMWUEo9KusRaxl6NCKPd1YSLA
Zhki66FsMBljdr1OZY2noOEg7EqXiYXUDwO1CdmmHk81tL8eeR68hu9gMD/yF6x+
`protect END_PROTECTED
