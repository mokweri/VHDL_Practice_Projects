`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kLRby0zOptld9jJ7Y2rt3FsF4yBd42nrUON4HjU25+0NuolRlAe83crLujvMlhQI
/YM4K58mh2OTDhbRrPgLKYLisYpAV+tO7HyDeuXq3lsdmYLi7QB/tawtt/hOTtKw
qyPSSs2pjlYSD+U5sRb+Yq9QTPCLqFpKevn4QY0AJdr7BIW+P0NLPqaIiJrMmjAN
vRKDhZw539Yqil+LCCdlpjFWYHIqV37XoEWNsDAIMW6wpTZ6Ki3r0lrSxQrGiiZt
RwIs0FFZ1RW6AE0TjoEqb9jtd6+PeBvrLmKaXXRV4G7OOVvwsb8L61FSUhDp14I3
juXv+kU/cfUVIO4LtpRxVQTUSpO7OQEkE/M5AuAqNfNOy6fFUUK6Zjq2RbNp7hLB
WUmQc/7bvSf/t6KBUwlwX7mxAGtp/geiU5vpa88MILgetM5+rdr4Y1FBMnCLOHL1
0oc6mVhgMbKWYtLdIlqzupq8+nDRZLNBkaztIt/dnMGPvxhYejQvjxOg8ZoufzMq
LJfy7FVChDX6tSbUWktRhHd6IeQ0sUpnrB0dHWGScLGvNiISsL78ZjOLIV4KzeK2
gQP8Dokx8444E4eQ8I8YMGRl7Facw2qfafdpJaOhdL7jdhNN/giNhio6Kz4HwTUn
evgSTG0CWodx4Fi1M1X3hCMZyZHESkjctFL11cw3bqLIkQP5LnHVRROvvQpqReJx
3Itm0QPoRWqNeD+9JUarGd4+X60Nku9ibt0VpqEXt5motXlhlHhzb9PkdKU8XTVt
Sb/adqFrT84SDuHwau9Hup9KZVVn7Prrckcd/AjAj71iVZJXhNVJEPCLBBGmOTDq
DgzHxZqA+Jxdpn6fUTK2C6q6lGUZdN65g/m7+0NfMORpZZizi4e60PXbMoDW5iud
lumB649HLvy0NGrXM9uSsej4tsHoCtftT9fShk2QeTyKE91/Y2lbORNPSuLlqy1K
LfNFJAWNqah1WIF1agfi5WF57wieSVR2y6C5u9+CcZ3sUZmxRSZGnP6Tv2vS4Yh1
/293+P8CjNe3qKQ7AZ4F32ibiCqokPNoVvJSJOEod2fOvrCa+2bxZf9FzZjgOhB1
4oeUHFsHpN7CcfbOP9GbeHAOVqlRArDAIM99MT1LckQFHzozNezS3u5LNg+h8Tpk
zmZlHAC2EUxUkQm/K00bQc+xL1/JApzVqru/xggPNCkE1/8DXigov5hLaKyir/eR
blPxh9BYq6PqdcIZ2kMT26b0FAA8Pn0U1B9SoVUou6yvODEjnWT05Ql4UcTusKy6
LJHUo9gYGE60eEnsKm+JJGpqWSxy8PXmE5viRQe35ZnU/v6wK0ot3IQUe11k1pGO
XrYxb/r0Fq+XSbT859Ut6w==
`protect END_PROTECTED
