`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i6v82BsscDiM18rrjZAML9NPo9KYJze8pMyCzdPk9339iEabKm8SRArITlX0SEjO
woyI65vwJmDy5E525KyKfBUF/30erNKkRo1ev0tdrLkWdURxGhkLOrxHVmCvZZv3
oRMmKj0i15/bl5q2YyVBnq3Hut6BgrrnyHI6ZPbTIur+2nvaHhsgzkPyCpN/CTYZ
kVKD0mpM2ARHA+6o7u++Eoj4d4ZWBcR6WiS3C1Vq1JUoC+6ePSL7VzQcx6cVc1/b
OVFIlAmVPqNFTMP6naukxhKt/c4dwn3azLUWmjsWSZ73cGQRJqjCFfQQHkrw2ocJ
yiF6C9tYD2vN/ACu7iYPitLhW3Sx2IHUfM8wK03MZ72x80Z8d34WygYHQNiAuDK6
CWcovc8uxawk+WVY22APyBzmP8cEfSIifNYNyoDsCrwrqibTk36zGUSkpVZV3tr9
feusnZy43CXe2bgrl29JK08pdlP/Hm0rZzI0fh2dB9x/72bu/xSrCKD2BZX3IdoM
xxCPCppbp1v2lNtFznDuhA==
`protect END_PROTECTED
