`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtQGVXdcIm5VehBONukaAlgTs5qvg0Vt1TehJL+BNjVWfxKxOuaUm9XWTR2oLYSo
lNztM9mpcZ2fSyR730yVBYcYacoWm+2Mzf/s36ecWtLEfuZ+SiiHkwYCKcAxauow
T6onmFGOE0RON4456WAjTOgFFxWaTa4n/g4Ri1QDI4nQcVapT0OlCs77W8gEWDxl
7c+Nz8Jk19Eg4vVLOBl7N/pJh8I20MHhxVgFm8nYYNwGPN6v/MYAEUUwzo0AIlqq
tMXSXqtyz+ghqV4uV7fY11CUfNvjjpXJ+7zWl13fo7B+dyMxDXsXS5la/03fHa36
J62XnVXf84xqnWv7gqEBsGYsDtFFP+GFhSv20M5ObZNx49sepzwxDnZf+dBD2tLi
Z6XrdQw5VSwGdI7nJ1Vy71c/4udz52h/Mpi0VujMtbVjshyGaQt7Y1vk/NI1qZeU
i82wG9hBiG3TLa7sDmTs3AfeE9ATUjcL5i4SXMVY442cm5QsvEM7OqgBMXL28Pi9
rPCBtAey/smSJUEIQaGnlop6qOXSI9utFpNV0/1pEUdYvouAD7ODysQCLDB7kxsG
oJPaFbl8fSeXWNtSF0uANXzNRJH9KlteYIq+CcAh8B6Hq1ivtRgiKrH63zPQTABb
6q6w0csB7HdC0kGIeh0f6RN2kMQBNRrw6s40qBs1g7bYFjlxalzP/UjIUzeIFfWI
LKrLfj+zt6NRdWppxsAXnuLtuuxrKENaJejkczYvWEx9feBn/yZ/431FDiBvBLoi
gC9UGW8vjJR9/BT6TnCtjME5wF/D+nY0ba3gqFuZKmLu3gxO2qdjzWlQ2mdOoX9C
qipnwm+Alp6AVmMrV0LcQLaFrFTXwYYC7l3MutvdKkiDe/EELG+7Mrav79Ws5kf9
H8A2nTaQkzJP540wJdXJI/47QKZ1uPwJB41NgNen/06XVj5aBmaz5SAM25+Vqc0G
yRr531CjivgpTLQGmdW/nniHR/lYeN9gAdDOiMcAdAOXftB3HSRCIzJ0ewea/oGO
Ha8IztR8NGlpdZjJxuNxB1MmMyumDBy3Erde8mqDrtbxJ5097DkSiDBdlM/0kfpn
zG1po0cj42r+hbtQYxtTbtYdV5BS9opWApfCE7DJf9J4xG4Emuotoxd8WdXGgKMz
iF9Ov9dhlwByQA5A+iAia7wLHWsI3UZtNgru+0REQGAZZ51W0+4ouot/eBa5qFgE
/VFzecGFeYzy3XLneQ1JzDmkr2R7XOv/JXV3VySdbz4vwGBHCdsaiutIwaKy/SMJ
ytVQnWjr66cCF0E9uCu6ykRnXUYD8XG5zKFgbC2f6lU=
`protect END_PROTECTED
