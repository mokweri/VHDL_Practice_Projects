`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQXYup0yHA9WultxcXTCv4hT+pWKlp/f3JPUoZ0gbvyRnVmJleERU86aUqoqxuji
m9H85vthrKxMsHw/RDRE9/LmY8lLApIe1HzqxrXiGJJ2llVNjdnLL96vIjr+8hx9
dSiCXDIHxKippJPzyJNpFOcr5G8wEMfP6zABxZVA4MWlXjbqId3V2QZkxAQZrKNd
oNJJFRm8HtZsQAfp7E8ngmjAC0ytOwqOuwzhk0Pmmlizu9trdxACMJQJFjOBuxUp
V0PWSwKLiiRpRdFtAaXVnoGR23OQFnE7OgnsHlhDkh1+9rDPigFanpfSifUp63ip
inL0yopZPq0T99pYf8le4qR0Rb3IFaT4hisusjVd025CwwMn2dD4op+ThgpXvxD5
EAyIJHS+nrABo6/z4tPGhVpjHXWwQGBUbIkkQFtB3yWFzLOo8xnEMucYX6qleesZ
C8QQ6YFMsfOyY6PUuSgGNERrqLHuZlyU9CMxKNYzam3pLBPj282GSBpchNrJZPC6
pU2e7D9UUPLV9uFSxc2YkK+hEel0D04Unma5/6VmU9WZRgOvAJ+NdhFMslou1WWX
D525dc4jUyJPWhf8BjyaJDfVslkg9rkxbtT06I4Tvdu9HttpqCG5u2km1nOZh9kT
b6uoMApppMlBsn6HFhxPvv3P9klqJc2ivtv1PbeX9Hs87R8ut8NdiYO6FOKnT8AF
Y4om0Tumbrz94gCaQDy2kV9AtKPus0dQsGCaWGPn3dg0yOVbxUiOALzW/wohGseX
nS7sKNSumzmqVvItMv+lGtmp3LeO6mGtnpPA2x1KgMQZxZvBce21z9NlJBZ1cY5p
vMLnvnFokaHd20jMEH89MjCZZ6Dm5FO+Q1OgOUd79CQeY8Vq30yPKZypr0WuZwWO
g0QZF4DmqoFbQK/ZrIeK0khC15PwFBWGku2osmuTHoU4ql/9UKnrFvtkXwOcN+qn
/+16wZj4CN9cPtg0EtJL19rsXD536UG2i0MljQRtxYJSIfZAWuKVt5BoLeAT4wU9
XqTKeBHBFid1jhU9VsEdvlCS7sEP82jAwdASKegS8Gg=
`protect END_PROTECTED
