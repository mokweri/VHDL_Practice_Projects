`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWxRy8M46boJjMXxTrrqhS8HGyvW/rPT+ZzfusPEn5AulJTfWth8g++4u5h4Ct/Q
0bt/SuYRiYu/yyOxCGgSDdBiqVyZmNjmUgKJE64ETFGeeBRAJ3hlSEVRoixfB3vH
vEK5w3dvWfn/3JUmyz4LtMA9TnAp4Mn1OxLNkV+y0ESswXn1VNORLSuZBLWMz9Ta
yS5FGstGQRU9LSezo9QC7QmM6CgI6cdd8FifuPJnM7IzsQqb3mVyrFpZCW3HUus5
jZF8pUpTG+r//RXWxV2M8kCVaCZhQzWLlCr4WBqCTpu4Ysndlek9G0J/5BpM6S0v
LJ5lmXmPiflBpf73Fmz9E1VXMZhnP8zxMDZKYWsshmN5q3YXuSI4YR3SO74EojUr
n90l+oCmWVLnDwPxRtrgkLzEMDlhCF2tXPLURFFLOtjBrybU30ohtcqWVod4ZhJ0
il+l9dOt0+ABIQ8CyB3CkVZPmYaq0iK60sRgY2IaRI6Q/e/J2bHB6YuyLSeu7W79
jjiCj7bxEQJ3gixICi3bgs5RE/L0vDC4piFLk+j7o4p5Zd0dKGDq0ZCcjDOYqsfF
11VJvS4NSekc9ntRoNsPYjmuxkhMpvv2M5+N+K8LkCsPCB+5DIEfZC+32lwyq7Sq
V4Bbgk10YYRa3cxEf5Uqsntq7v3pnvJRjidgov/HGq0l87Djl2yLm6mBHPG3ooa7
z8agVw+sebV9WWjilf1XTxbbvAn02zd52GpLstlybTPijBVsBz97AdKYzmjfrDSf
Z5tYfN6IwR4I1sPVyG2iK/PuVNPFSbB3coZINvm3xFqhCceNxWUhbcqQ8QBT32cX
Tv/Gtc0iOtjY+3PjhMcZoP3PGZazLUHNSGM1Al3yfcxRkcBgRdyrUlBnhhMBJ3k2
fzwjpbIG1bCmTzmf0d5xdI63ihjUptu9y57LnTJYBGxXeMgzSRETnza7HGqBy4V0
6xA1rjxMHXmyEpbbuacYBuGtq081KysmDdK6XAj9gc+K4gIQvUYQmTexTYnHOwU7
RdtZLLvwGkRqEAAt5jrZ0VZoC29u1QDhuR38CoPVLYj4IAisbNaDID5uWd6BKmgA
/2AaxOQlln7E5X7WVnJCs3MxMUMB8zJl6QXtAluwk7qbNeYgBcQjjD+yOb4WXwgJ
nUrrFzKUObVf4DAwLIYyr1DJ5AH/DB2WpB7VBu5LoJogfnTXTLDOz5J/C4FPxETb
QIlkCinZP5c0+5umv/Hfwk1kDRZQgcufPBneyUMvHwvrEjnxZZ/cEMQLLq6JgnQW
r0WxmZwFYKjuRB1c/6Xu5u29f77UCl6UZNWzpKOOBpFMguGGwtHi0A9VxC31e1bR
7aspXwLEvkWxBAElt8JP57YlXMykZIdNYVWz2p52sZ4pHHozpMT4+uddJNyaFr2l
b2jpfoHybs/soTovfvva8wuKNPQPWxcqN5S0KoYRVeNs6esvXVeIvTg/A7q8wlzG
qawHMebzhLApKVtHz+QcMCsX3T4pHwkSCWBTGFiqeBY+TxotBnvc1hfABTnaGqnR
3u+jwJDclFRlqV8EHiHDWnW8geExkPpWqlfCY0ahFLFhmOmSm1KCRar4pYwc8BPN
YQYqJxxu/kk4Cbr9Uj1B6DzucGkpa3F+YxiVYNdyHz1LMcma9GMf+Zcqv/NEJ+w+
Pwo6gNmi5M8TqRJX0lKR3DxIdxh4ld7ZLkkvgqwcI71/9xRSYclfKeB12tZez1wb
EuBXRNHvhAKgEEwAZqg4lRnU83gJFqXdPqxqODg6om6dWwu+MvJpBxXF8RkdWkJB
F/RgNgLPxWyjLGOYqtcPa7irx14BivqY+jhVQy0HYNsNI420xj5P0rwsVjmGmQ3s
9SpfOc4bQEZkcNuR8hSYgJcHQvyF241oo9PBiV30GsaFbkZFH0nf2ohtpnggKj+Z
L0Aj2ixCW6PHDrXUb6M+K8TrggDfL6IaikbwH1LgJ9n/o4FLvgbmU+rVpXp2tarw
f8vkPlfmcY0nMaB3eIJpINeyUdW8nfpUvvYllBxcl/byXZuN8IHaXq5wZYMUctDI
jBhohrKtoh/z3jZPr5Di3xByTIHjt+2LDNYcTb1qA1YwmFXMwjP0LTqKzc/gfARa
RlnaGfE//HSKVwuixmhZCwfoIQiFaPpEsmFj6GraYo8nBryi7lPHz5qfHvNh/vQN
2PbsDFV95UEEEFYNvcKAAlTPbHivVqoiJPkApmOUGEQhztz8ESJR/skrlwAOsk2Y
8D7Z0GR22zeoZjbY6ODBhe1w0jOySEE7Wh+l5Yntz1FdpWhS5UBRWCxb2qgOmHPP
2FFo+48oYGw5O/brnon09dOVWXdUfg1BDO6n4lyfU8xNmAhup86ey6HLWr1RqUyF
1wV25f0wV0jPF1F5J2yHl0V54K9tliHZQggcTnHVbSCNlHsJYhv10O2m2yvpEzjf
BcBex9YJzwnveT1dgaUumiTkN5ezgXnnWAFghvcs3uy4f4027iO6SSU7Pc+a/mKR
oI/7g1C+YwvNu5TgQYU3u17nBtfzCSzRTL5cqA4bfQDzsDyCIITvScNZ+6RXbCR6
AQ9ys+elHlr5l5a3U55r8Z3VC3+U0RyZtYOoaQJDuseEX2r3eeZAeeFPkpGXajaU
Fn/rnjIl5ISffToT8o/7v6aJxGGilzw5HNQxVUHZbJY2UfW5WnbjX2KhGIii4jgf
ID/OF+36lWpsbNA8rkp+AtSC8Co67wsBRslsbXkK+maIvMAOg4KnEFN3sXvjZBLy
Uv2EwSEAtVfF5rTqO6oU2jYNBQVikxe7kmYgXU+ozfAYFOWoHZ9gXD+P/rWyRXK5
nT0t2VMDblKZdpy/y4gjVWHJUBs6vm43Az9xypTwvaHQuTWbLMeKWHu46tepwicN
Kv+sNqf7av7evdzSN9DHuDcHnKujqXwojhihM7+sezuZ2VudqfqjvcZWCRQ7u8Gu
IVNbGJzYcySRX2FrzySVfgs3drfW/elr5UdjnvBDvS2mdVh8OSmG8rwnoQfP4ZK2
RydpRwf+4aWW29S7LoGhWVNRYRUSXdnJJSE6oInxWEJhaYMmHgJATRQLboFyYb/k
wlgIknqBtTmtTeAodlzZcySETDpWEEtvXiyyjB5+0coPuriLAaGiabZqKA3r4ulb
4wq6BSwdv1DHYs0IlvT95VN6CjoBYjeOBWHbDBQggwkpipsA0Cn41a4pBLCZlf2V
ilYJ2bArcxOwhqQlDPuBm4rO91u1OxXtr9gDcXYHwswbssZn0xI+4R+2bfB5ZAMc
UGd39JbJnu82EUFOwJ/qTPOcJKnDl3ORhCJTJuIi8A25yraeHgrpOVpV2r6OAhga
WiuMHxS0Wo09Udj2KAsLoZ32lm98LfXeIEzuDWCT2lKdDp41oCkNHB3fnpd28GAa
d0NLxLiRQ/Thg0EqQ3SFKrIffMnBoD8k9vbQ+Pchw8XS+cu8PKDjUE2mFQJjg3qB
/hM1m4J5f8v7fgJda4QJ5JH3A7WTnn33vwhTCN542x3zyXNTIicAsdYC6PjhHYcc
bFFbQWV1vr00fKW/rvXImA7WFTuRH96nlevhgJ2wtXyTrCQDbkUWGYSnm7kyIGjw
+53fj0jY1311Qds1wZjQYQzA13q1qIqbFOCmYF+6lTz36jxdfep/x0VyHdeUvu6I
tSKtb08UpRT/u2xjHJlwgt6k/3mpqw96dcnYorkNy1gUiga8GUFC4iOfThpGu82S
b+y5QnVTse5U/5B5ygQwtfmrpvLXUcRtyDCnFUfUvaa8qnf8QOJT49riMXj4ehge
Up53FdkmUiD2mCRRW4hhU4JdMzbEsuGpg8N4FyOCK5Ag3KWkDhBoePkUf6kZYszO
Mo1Vd9tPuIj0w29mxiQM1TXwSl+jCHc/vKIFQLsDBOOSNQzgCtdYYkTZ45NjVHIZ
UzIDg0FNFX2T8Qn1asjjZ23GrwFssa84EDJzGMg9ufPWNyPdyg4UVoKOqji5ABY3
YYvJ+1dKnS+jXMbN8rmkWK9ZAyKhQ5WSWSz0goa6m1SfjH1khiqWM+x54YbYv2fp
IuTJyky4/kWKaOivy66z7EnyzgumZ+n+Qc4JdsMuGlymlNb3am8geP4J7m0VLETP
objSP/fboarNm3f6PLo6ShFoPTapPbW0duN8gahZggVnKSRkXxjUQmT+OETYebdI
Fjbhz8/wHqgXosw5DgrJRv/lOmnLdqVD71jtrL+KKn3r32b9XRGPdA/nh55iatSL
eGhMk7THACcOHgSNUhA+kn2ql2em7FGR80SJ5tXfM/FVQEXahdp4m3wmn3h9/At4
NNcrgVN12GcaKcaMD/+HQdxUx3pOwvNEp3gDhwq1gLqJpLd+CdE1PXVayNY+60/3
BSRDDTgAVpQHxR44GPVaHi6AZBshgnHmMKTLbJ68m6q8uOIuCC7bRdjhliYd4EAP
nBR9cgCmAsQQgUBbnfYyT3aQ4bfmV0ld90HLWnGzrPAFcMdirEXmwQt99Ecx63Cw
nxdbeJ4vN23gAVyTmd0t0/hjWuwKDrG5WjQOyAsT9EqAFLQV0xrxSEpzS6lF5gD0
7eeszznAFtZiKbSbiA5H388AoVO1v7xQlRAo+4r38hLz7/bJqwPLHU7HNlcKuxUB
uuVDgj2buJ+7tHMqBZdRbvOP7mlxq8FOVZd3WIkA+d7HhqpnBTTy+H2ZyPFcL1EN
GV/ngOLzLr0yOqxiW8KOogDtNI5Pc5h9ugb2Lw0iKMW4WglObvWhvHe6jinALW2f
Dz8/GtJb7EP4AQA6noclWkwhr5vDsOzQo8HNOOSsoGdrbTA+XES0ZSB2KQ7bgN7E
OtWzM4dsD3UkYAfLUQnhQOr5UNaEgrzwdHzmlquvlpURxA9PyXA8qLvVIbyUoJWU
2d8d+QP6VIsx0iLQI2HqlOQJY5qW+T3As55S+8AF045GZgKRoQ0fb7LUkpTdI5p1
/QF7VGRVgixIpwJq6gZmLJWw/CKhpr476fAXUy/YNqcZxTH16hLi04LkuzgZWr2j
Mt2Mmqhmdv/yLLyBRXCFscSy9vpbmqVKv5d1aSaW/r7NITroQK9b+fbZUwDRuGYw
VEjIFE5U2yuqwWh3m494kuzt2xwZ9/5xFnpGLTvzNKIYvVfnMl+XHD2u67m+BkSp
M6606f5Nm5HaV2idkFfzTm/CS6xyqdFfevfVsOSfGDaYbf/+v6RgrtHUh22kxqJ6
lQJ+Itdv83TN0RFbTGLqyUm28ZfnuW8lnANO37YE5W07PTB5BHl+QSc0MeezLFsR
dF1GkgCQBUqDX5Pl8uEHnn9T8tK4zdGDWRXvuhBVluBhE28Pg3lUJA2FK93yatA+
chTCM4K39SfjmVvAi/1YJ6p5A0rEknL6TU7k3kajX8HdfR9zN6DaFt+eN3ll9nwA
7mBFd1bsWgYV/Igo8+KsIjDX5xGea16BCuxNPo1EFLvNmCD7UDW0pH2MxHyQYdtb
4ANbms1G4tZssbJT9QNETzyGzHzz+jgin4zczldgO8jOjyDDVP1vlaOTtiUvEcsO
1uQ3cQnDcR7LpMbG6aTbgG66G0zoYyZkC2q9y9o7WxdudS8JExn38Xb2vGom/N7Y
oeo5SZov5LDS7LOP/bH7C0g8l/lnURQ++kDUoHC3oc4MXqx93s0GOVgLKg9Phizr
inm4TsjajP58ZXeUpIIfSPwkHWnMPeOn3iEFDDU0+zB+zpkTn7c9vLdI9pN9YCMC
T3Mdpi4Ir6QPGHu1JSe4V/M5BmUUl+IST+bomAhbjaJxIUe/rfc9r3wSJJi1X+3C
GxO5VxlAmz8tO5wUBWgr+eeuab7HEuLhztrWP4CCufoUrxLAvsOcCTBFjaJqewYJ
i0j1xMdttyakX/Lmd6tnMl9iQ5ImGqj/cFuBVFqCv8JyHA6FXKRifJwapds36OZ4
ca+rwW1HOdiNNMp7L2eHdxEuTjdh/BcOwyL2wEuebVNEBNvSvY4Fo5LiSG5dXWnH
Sl2en/6SeHDxLIo1CSCG7EKajUMCR0ctzHpvccH0+Wx81+vMJAJIQC34/9wEnkRT
cl0kOdFOF08InJkEUl/OoU7EcEn31DTIZFN8CmSF6Ne6+xIz436FDI4posnyZM3k
lUn9XrYkY6zwQKuxEIQ+bL4Xp5cqBeg3cTM6942GHv+/mFQtM/p7aK4vb2Gag/rl
vyonoM7L4vUbmL5AU3qm6Q==
`protect END_PROTECTED
