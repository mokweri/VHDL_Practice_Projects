`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjAi0HyyhQAovYxOphIIuzBWqrdwW56stqKLXnkThwyr/Ok5poUabOolqpBh/JRw
+KbIblx5k+2niUEFJo772pboTV1il5LgNOGqlUa1va/Tjpj3Z5yKUxC9PlLAxZsc
eNeMTrx8O6h9pMOuFDqEyuxS0+YePS1vK86XOdg/wSzf+3bC8pkzRgRcfYyzlM0y
i3cRCljUpMjvfRh7cklQZln/pg/AjkwfNlK6/DoFuZcBmGRV0nx9G+q4HvXUfaOF
/kwDoPafvGMydLXIgm3WpuyF+EK8tX7y8EieeS/n0HzJp3FLiXXAX17MEBm4/qsD
dD7Cytv37ib1BYF722w63hWwPcqRv6mWMsbcgI/Qn/wbsi2KGnoyPTLGECsU4AJP
FykLuH2EBpeYUiz36A73m13c5+l6uN+JZSg8y1eqVzrtODNywRtDKk5wy/SizlAQ
TFGIVjytTl6hZsVBmfVBgjXbId415WM5dltRdCGhr/zcdTRZf1sCwwInX98+PrSm
bMv7E+VcMlkv4HU0nYzeKpPfLAV3NRkoch2EQ9IsTkzJNdZ53SJoI6X05aio24cZ
yUBI1GESySEal9aPPZz64HovELFxrk821JrwsFxON9H8EcnSPhCJcb/S1LrSYyRU
gvf+1y5CbYJvh9ed/klIOQkK0NQQm5a9Wh93xBjo6t8a1Dr6SthM7peWGGU0xHbU
0PyIwP5a2kaC1Dlx0tkwQus1npgwx2Gyp8C3DiEo9aFxtcC9NMi565lO1OiE9R7h
usRrMYCtUGUQJxIgN4l8jCYjulNJxNZheE1kRqRTJ9EMqJ8r1sX5K6C5OtzZn5pS
mS0bl6vD5C0ANNjIQ8NVrqKn7IX7RCOQ9yzDTbck4SIgVrtlqFeHbtRvhG+6J2g9
JnyBgAhIyJ6IylsORxR7IK1t5XuzQoW9tNQkvrveHyp60sU7HPuEk5hR38Mcbf4C
TNp/y28uUmaccEpCFOeHmIoguOeGFotF2cfy4bZAgoY4pZPseTp1NobMLHxqsyTN
hcbMFol3tjO0pG47UlvIdYlSPm916WzMx0aEB5gilbHDtabF/D0GENgTqesLpa/7
XwnLljyLcMSrtczwn6sindJ9/ou+hJJiQwToRppsafR7SqNRjboRAXHQ4o9P06Eu
zZaCa36bkkj110aBrJPWreZRHncqd7DAt+TuGM6wuia2IxWnpDdIOWWC5QuVqDFw
kx7UnhEJzib83JiSfto6wGUH0kpBoC0x68LAsbvZx2yK8s+AoOijGrXdwBQ9tlr/
VyL42J6x+rPMuOFElV51D/hXNGVCLgsMJ/CrDY74yumdSK6iFvQkza75hi8twCEp
iK+6AR4bAwmRSDoF77+flsV7UY5q6eT5fDZ6jKBUpVT6yB5Eo0lQKZZnygiE/AoW
OIkLnOKd15cEppB9RJXvth8OGtQTQ/NYcMrJgY5mdecM5ZHQjPKCzDcCXOmCE1zG
AyR/N5M3TnIdOhAgA9SLQIhWP2exwuxncfPUpg6WAqvio1vFx5nsC07kCUvC8DQp
EhCcee3E5T64593Sx8UmTWvUSW7I54n9w25XEMB3pgSsM5TFL2FSwlduIdeVf+rs
hE4QtqWBhKCqyby1NZccGms6M9/SQekmEYuaDw/cidYWEfywH4lVrDOLjDVrVK5N
VGHiJ3A32xqkpbvslJE0ADmja36BAF1PYi/4q/Lo+rsmqYw0aot4RomoVfwnHJoF
Y3Irx1MaS+14QeGmU3giwedSavWpTiMYLytkHs75khG2wJClAjPa0lLbvMxQlmb5
EDKuSoPmxHcNHeEZwZJSCAU+ou64NlCTMl18M5NsIjsdSNr0L0J3NfwXdUDtiaF3
x+a9Lk+7pOZUFYT1ZxiPYHmOMh4kB71M29rTfT+fvbx9QJ9dvApmM2CbmK2YKBxM
/XKKv/qdp6+kt3uVnCSqc1zjJTgggysilHms6+8LfUFDIx3rV5CCm6NXwnc0maRC
loeAWctJkP0HbL5d2jIupx+b3zbNdHw5I821gXnLr/FctEY8JhQ0YNgPn3ecaMZv
5knevX2ufN5V8vT4OJ5DxCpa0DFik3O58kx7RvmhSVS1imW71Q3KC9qHdXG7acHY
aUmBFvdivm9cJ+GPba2gzXyBS01ph3elz8Oh2g4vuGeAETWz0XCX3NwwW3uQSxlz
j7CoCUAcpx8xBSHmzT51xKArcDkoMbqOSh2NU7fVeJb07SmlCXUaTWrYbt4JCqFb
rHm/hg9bsZSdTpJHC5utjmQeHzDvlhWJsn6Y5CI9PfrZ8kjJBN1RRhea2uT6KB3U
ysD9HdIFIfezD1Ao52GQHCh+fg76GDHZPzUAiPazRkFTs0Wp+X6LtEj2Cgc8kkYr
rKZZacPKkeoAXdVSKY0Mpco9ec8Opum69ynSM0FWZZxdf/ukv1kLLDO3o6+HQ3Ua
hinpUGHflkuF3Yhl2Pq6sBuzJWh0ugZH09ShdR8UrxuVMwUh8LhJ8n4cBlUcg1Vf
5uWwCOEZ1JQE8lVE+NwObQ==
`protect END_PROTECTED
