`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nIylLIdYMYi3KDY/iZ0016TD9Uo8koZ2DBt+MT9a1vGkwdoBR+3en0ETksFJkygd
0siVRn1fjMLDKsGecYt02/kUzMLaY89uRhuAiANVzp7UmE4WfIrcpPIGpQviwm17
AdiF33k+757yhLXFN3bCTxvoq5MMuVL6KGKZdPifqbr+dB4xfQPVHn78NZOvZk4f
7lXRickRahibc63Dxgt4gnCM0ExXsND1H1dZTL1niVwk8nqAfhPW9TyMnPC8EQYg
pUdXEZM7T6MonbrPSPg1l3KYG0Pgp3M+LQWJ02ZJRXRTanB1479kV16ovsGt/rdV
rR9mojT6bxH9GiVfoEJlh58FDMWC5nMAeoJgNXx3WEUGOF2MvfmnJE8/Qkx0BcW/
eKImPMFnBX1iHAXOA2Dtn+u2/pilDi7QzG3uBwtx+nhjd8Gncv3fZ1afC3UXznhC
26DpbeZiiwJtZsYJo+MfiEMJU0VQWuf7Crdm+kB9IU2hgNhqzBw4gnJXFws92Fq/
gemeMU3kchXYXYIsd7xcV/dtVtIlXyQZ9bVwccv9hB5/s+p8GSh2Nond2vMID3BV
FaAT7HWjWaEW9p+odzMU9ky8FimVFSAGhPSsRWcb4R8WA6fYOgHimqwbofUOwNoA
bKS5ETRLms3k8iIABJ+MjDKNA4SpqkH6Qq6D+XQM0gXB0V6VzJsob0HH0fzUOSpE
pPuQ53Fr+P8HdL6OYSG8sUuoOKDf/B3RweP/8aW0sOnUw6tANUE3qDUWEMts/K+g
4r9tScMMaWxnkuYGYV+RwIKfYenPJhET0RCvDKLEz26bUDSOP0nsnAEqoQNtuFS6
`protect END_PROTECTED
