`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dX2dP6ANFlnHq2cv13KIIBmlM0VtFi3FZycA12wZjTFtr2xd3szQ+VK0AuZLaPf+
Er2Q/McnHMoV2R7swJDnpi6SY/CpYMklANu71ZqGVFmOAX8ubKcc6Thy9/fVP1nz
Oelbe3CaTcn8rWwks7A6n3IMLOf4/Oqr2kYYyfi6CiaevYw9LsOFOC1EbLmDOUtb
2OLsSFndIVi/IIR/0SGbCQFJRZ2v1d9R8ZlmnzLZ6zP6ergO5q52Eg7n80qab9ng
PV3KaJzso3zaP9b5eY3UNLqRKJrC5dcVXn9bC9xX9A6Ekr2QYD7Y7+bLK7bku73v
0VsL78c1z1KViruKLSsAb15XGUKSaZzuMSRMuMnwt45xqBa1Az6k0aRsvhH/EzyQ
TYIKHrEKmygmMxJgQ4zLBWr98z6k5QyKr1PRWPR9vqX8mok+yZyr04z138ojmxn6
wjhnDhW47f/JhdfmYh0A3HxcG9hNutpuUG/uPmrmgEKDLNaPgy9kvjnLMxBmalkm
37lxO0G5Hh6fDbUU/LPiyWgrX2zix7TEQIOXqSzUZiGFovD5VMrIV7zTgg6lpPI5
q3YBVrt6/k5VIa5XSRUcTrabENQMr1Y6OmgmduvhQpUxR8frAlhFgbl8pRke7b70
Cy6VTltcfbqYCPsHg62ash28DDE8797CCSHrElxgvH6bqJPnxH63yqu2K7MdRAw2
F2ccBnbGaOj8r2oHgWlAyWMnn2tD2y/9oVQaYqC+nb6gU4Q6x81eEkuuKAKkmdkS
KxTlNjx8RGs5XraO5vPJkwUa62aV2+GGwso2EsueNPmitioMfngkQKWsminKPst/
bNY1JXxi5ojchbwtXWzQxVBGGg5ahP1ni1gHQPFQkPYQKXl0TfM4OH0mjbExc/ui
f93yDBG8Oe35NMu8yvOOBaP4AKFvsil6PJdkc+3+zj4Ztf+O4Nvz7wvxXmLtLxpF
v0GE9+VkMc8rwZmWkHx80otLnzmBzFqun6uLGF/K2e8lFani8/9K//3aplU2RRnT
q1oN8B3QRr6vYbe+uDtRTVPOZie+7X9AZIIQrbpCyufY5j3b5t97+GigucdjiQIr
de5n/8dIUX8B+Nppjovls9sbxAF51UU6Y3jLTytKaxgoXrJHAnlx8FBKEIKH/54J
yNJQVtljcACYkKWt5lmR5VyyhAB8FOO7wzmiVPsj567Lyg24X8sCMITdaydabVYl
5aVgxe3ZoOmw9mw5oGTJZDggmeNi+xdJnEkOGpqIULw/dVxrmywLhWaIAKkuAsov
GWrxXD49rYzzH4DBluj2L3rNPc0/r61JQL2mrZUALdTBUiILDdKXVSCpS5ns9Y1x
W2Np32ozpcTheiNja685QlTqFJ+Bt0R4tFdZ7FI38BKqMYaOMASOGtPoVrvzQY+P
iLzF8kOLuc/FwdWVXj68IyGumNbkEtTfYUb+0PAaf1TveW701wlpBCehNycFWmsS
Iyy2plxFztEOttxJL8cmspJUviF6vaHQqQwJpOx4KPYAi+QZXqY6ex5epwNKdX8R
G3qOpwAFYHbaXMGYl9z/+g==
`protect END_PROTECTED
