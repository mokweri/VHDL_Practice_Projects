`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jJ2ZDU8lR+GGVO9tvSbgQntXMna9jQVH2kCXlI3UnpCLpIkC9xk2SwHzcsPTsEgK
1pSoAJejNFTxnmsjKm9ZjuXZYCEzQGzCjixnWS1VNuv2/EYLz323RE5VIh3Yycaa
FcILS6n6G4Fw9dwpaNB0gAHjmQCiOzPIg9rCmTkXOe0+PlbQjDUAQkOlgfG71ZhW
Dcega+ObqL9ELPJD4qzRe4d71tNu/2wj0ebatnpkLZkZPdAQzi8+/2Mj127AH5Wm
8NQeROqpY2KurcSG/Y73SFIlhtMB/RzLFRe88MxLDvcz7sw4mTg4+L3iBoRD4Td+
0pR3be7NgSlXrAgFLLGSupUW1S++6ScjBtVy3Ns5FIzWbYTSZNbQLRSdFOkK4VdN
k4V8V8qy029JbGkMC5vclXzR5FI6p9rr+FGMRulmQlUlocHkKlbTVZBm3rTmK7w3
OcolgimoXgqlHxDafPVMB02Iv4HF8ofG6kYyhF7QITseLV/PuKL8ZRRaDczzFibI
4fn+gVmnp+Y4Z0YjXEmBf139dHTwhRSdsA3ABJYvxdlWJl6IpgJCrJEPZUfwWktS
`protect END_PROTECTED
