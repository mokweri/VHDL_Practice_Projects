`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80KCv0iYg2zV0mlqFi5/eJ6Y0WLJOyfXZl/UdzDaecsUKLHkO/wwshqozqy89jLa
A5OCQ6IRaFZbtNaUQFqQ1qqr9yy8TRGaIWi3R+9xKyepQsunhK6TR+09fC1TO4wT
7lpDU/btBOtPFy3/uLmPnq0yfyH3/6lUL1g9QodITA39MjW2QsVGHbV/fHkM47Og
1U2SDY/+8Cddf/3KIbiin6hSvzH29Qkz7Zd08hJpz2PxEHM63lP/TgsYN3/YYfqC
s06wZiv4kZ8q0z/E1yNQ9V4eNXihXGbbP4cGYdjU558TbUfHNMKUdOlk7r3T+Zxg
Y3D/DTE2vNuOJSqqOcVLQ9pOYay/2052Y6xw93nzUfh+hge1G7OP4uEZAAHALPmC
19Iuoo5r3ueIZD3yfJ16+bYwe4W36w8+Hk9372mLUEOzvT2vM/ppyKjFzPBXXfa9
GISsiEm25QShjmegd97xHyNLlBPnP30H1qiixyglSzpL+CiWvawvQ2Fzn2QXH3Qf
9dx5jGLsZDY6mw4aSJv3WjoEUQJ8ujDECRaFZnsNw8SJB/p+TqxM0TZ9n8j2KL3G
cauF47AfQBdsqToIbEXkeOTyfcrx/yYCMewTc/+RAT9sTkzkwaU6cdy0SKh0LI4B
iaw3MWUF/hFMGQbtYzSbU8b+hTIAMrWLJHYK0MfnFF7lmvl4B9a42gUVwOyQ2jlG
Ya2t/QI0XpDLWIK6LjAaxsjVWf350tvGuDqcPKoM/5Q=
`protect END_PROTECTED
