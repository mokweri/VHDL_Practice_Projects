`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEUhf0ssYAJ05gXOVuBNHV481ij2593cclRFxwkcX2KH6KOa1C9k3kqErkn8rv2R
LXegde/MCVX3Rf78r5JaxdRlKLtz1SM9odNglJHXqvvAh2V09zeYVAdsmvNqBVQw
uwShPln/QqrPdaoJsIVfnIqGo14HNutV+Y6fhbMZ2189wLZCaq4tMFl4y5HRfyeN
wsy6/MLHmsXc5bkjgimWy47Q+DN27YcvY8KwwjudPDAdwBvMRO3ukZ4U1pchqMTE
E/sM2ZBg9sWA02KJF1wO8htMfp7a24aTwLeehpX2cPvJtsYb4EyPqe5tRveA3FUN
dzbH/F8kkv95Bm4Rs7Le57TzrRbhrGfOCz+0gb/moKcd9UGyHfzXAviLshSXHpaY
KLDO+phTZPS5/B2nCuwPqXuq6J4dmJM/6VvWj6fZjcxrEEzZV7UnZcQk6xpZ16Sa
P3T5g8QWPAdE3pwO6XgytWDRfv4hfJXVpvivw46MwvQmrEBKjqoyoMTyRW1eNvOZ
gzWjVFy3Iuke/XWlqEvlj/Si/S5VI6PCvle1WvyIp9J+6G3e1FVbHTMn7/HZEInB
/n8kM5KTwzNNAlxYbm3RhSIhs0GHj/oWo3BozUmWRjRRBPkrNSmuWpjZqgrD1Yl3
+lnHae21t5j0B5ShJnjJ4JvKFkAF+2xguC4NPQXowswVzDIdd7PLDMz3nVsqATBo
q5+2rOXviOMUq8DMoa0Ly+hTSq7lBKaS39qTgu2sV4SDSTpvuNQs5aPs95VyDbm6
p7WNQ5ym1B77LzK0g4vNrnitG0s3qlvi4yr+F1xz/Y9q10RZWZUu3OITj+ZBnqlU
3VN1G4i3YsxjCqlrp01UKyDfvscFS/rdSCJmS9zFGcPim79NUIVE/c1dSKFsJuzC
JIW8nKT3Z6pmHTqrjST6EShGW+sb/8eQ4YC3B6hNA3Jq/a2ZVThvEChmYHaC/MWY
15HngvLk8mvjJrwty1oS9r67G+wNr5QQ8T6H8pt4Hftm2B8PDoZW9KxBWZh148OF
0K2vPBISXDQhHxYamXO1SO7GZEegwQFRfbXNHMmxs5OPbJZmDvlYSLt8xtc9Pvwp
fgqdf9Vw9MveHWGPVZJgwEroCuiLt6eKY9k8R79lYx317PfnKhC0fQc7TXvrsKzG
84wU/eraZeCOGiAO0u0JQbZKuRIiwwZzWHnR4bNkdfb4UfckOgLdrEyx8N8rWsSB
b2TOGIZ9BA1BnSeWcrhLnyV3j8fnYUr2AFNSnLn+3SZy40877vshH5IHp6TKcztr
ITeILCT6s4L6DXlwc677UtngZpPAKFD3XGf7j15ejZdD19u4PywlSIec38k7Uf/x
pvRMz6BpkbmRBsF4v1sPy2aYb5PS9P0EABuouuXC3NwHeIzUJOwnSZlyJohV0GoK
KrccO4PM3FTepvPdV7jSAeNNzR6xxmYuEMP6KHYwVzb6Mx2rafYtsupIxUeZPIHS
UTnBAB7s9tvoEkl27H350IaLjEqjahyMLAmDKRrOfLrQYOkJkosdxunX1VlaYnfp
v4lVwHLHBizZKvEWlfXdF9QE4EYbRDoIqjKvkdwjFL+rFo6wg9ivD8M1tQKf2I2N
UeM7z2YhOB1B5i1+8n8TIrrdSZz/+U5yLzwjgH0T2zAAM0PhXKdyAMQeYRX//o7t
1cfbC/X0qTmjs7QlbwjH7waxnoiZqKZ4ysJTNbD+sRA44rca7hlGA89GK/GDqBe1
+fVQGno0BYezKZ2l6jVXyVAA+ICUSfNcD3lk/g2vufsbx8KQV02MyyzmSKWqatet
eABByM5uY6q3w0br/17PY0UM4t68XiR4YtAga0rB1R5Q+hoNw6tzS7Tc/UkDwHaa
7JZeAiM9IV2F6g22E383twaYivV0dcNCjexp+eXBTbJo+h8bkSitwCBUW6khAoE5
`protect END_PROTECTED
