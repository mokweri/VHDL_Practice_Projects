`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoV64ogOA/vTPGjAFA0E8kozeJOmW/JOcM6DVicUcrHOtWj2nett2iyXxrliqr4C
I1V/VKk+ojVYBJbf7aMg+U4KMM5jEoDa/dQ5XVEpfImUq1yHVttfU1Fybbe1TJaA
AWqe2t85oxp7pEYam7YoGeM3Ed+/lphL+5+mAd3EL0UYXEOycubLTzpyu87bxrV7
cqF4EKc6QIFMDZLye4MZ+8zcFkujPKDqsG6tfHAlgT3/jE7O1gxqfRi0AL3d4MFZ
RfTgh6mylN1dGGV0v9KEo+WJyUkFqr0c4p8rAJRSqUzVz3gIPwCP8VOsK24Xnx9W
6jFwQhmwjlo+4B7NRtIJqsWK5NrysWzzdTN12+lH/U2iwlAnuKtoGxG385eSmRnf
V228Yh8FnON0jDiFhDn3he127VmR/0JSBl3Etco/9uzuWTr+51hrymXV1yBO8WxI
h07fQ6fmto/48LtEFpRZI3yBcm+FE5w7ufAd9Cj8rV3DOEh/aqjARISICACkYMLQ
CSxAG5tOYo4UotSNXXxRiemcBAdNbqopjdmi9M3Be9oWQUaq4s3x6V7BhBAIjnGD
ooDjTU8L1334yVBduTK3FThdtZRuH3+0DSYqNm/eeNuQFTdwBOq9J12NSGuyE7N9
FC8FZjgmjXr95aDFYI2LySe96I5hrFlwTRMsgyhNK05Bw4SSDE7M2MqopjLtWpkL
ygq4cilBRnv+kGyXbKxsEbDuG/7nFJ+4N6HBluoMUM8FPQ/FwC+pOLIjZRz66hE4
GUaNVS/y6HjeAfcpOvKdAkkwbnOaw4NafFh/PDWi1/gA/2Dv/U150E7KwFWCru9H
OeSL0dme6mdNDA/SD5/kH907UyUhA8IuN/fpP98KqyoMqiaFZNj11mXF2FEKl7D8
EJBGC4IilZqdb3B1WZr5t4UD4RwH9WDHNQEpvEHpEzzSdf92tJStofoqHU2LhKpL
CN0sRP1isNHmGkWTrWBQkykwTWBQGQcCDLx5Oz4Z4PWc0ganVaLBbyh+TZy+FIi1
jJWvUehr5sCaAW7VgpBAMG3X1UD9WTsNSRnOPCjyu8T3OmsJz7cMsh0K4CUSkW2F
vYzk2y7+8zFsO0LY1clRL6ucZaBZhSLS+7BpAvFI773Uk+WEhae+6dT/b4Zsatyu
rl5ByQtQQWyr009pkFB9sAaxwrN+lU7iPBJILBgls3JU5m3sLILJQ4qn0oKw9pBC
2elj7yABiaSYKIp+LdzUr1BOJqtiY3UK34dcI1q87uhX0TXpOgsjEIfflPYg3Pxg
pPmeQzflpp+9DYRq5i1j1nky3qrsXdWqgWK1KCy30Slo1IfyzNHIz+aIX+ATbJ+5
B3oZ9gdwshhi1utikv3Inn8z3MB6GU8KIgMAHdolR12rS2eCyKZOurzAfdnhXRc1
`protect END_PROTECTED
