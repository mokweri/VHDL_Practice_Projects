`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8ZQRZuwVH3FXqjDUq7dVjKM/AO7fSfaLn7NfMA4pOIGRKX0jmkKuLdegD9eyhf4
HStScjfDyFN62YIa6Xxbbkc6ylFnquK7Yue/vxKQL/ywXmR5RPKvnHeebrP5pLzw
J2imwRwocqbn1JAtpX6U/bqUN9CIQ7EYtSC38cSXsrggezKawB76aqhJ9GExmffm
gqf0qTOU5Ldu8/LbIJhhbBB1mzgFJbm6L+MSvo12zFTKW5GVeH35jqUl+Ca4XPiQ
Nt48FQxg8LYdBjDRhVCNkDGjRSl6m27L0nLv2G9EOtwXZpthyxdDwQhbaPn0L7xj
0HqtZZK/Q5Nk2jbU9e1VZsx4kkyVSIVb5G/FKLuxnDOhA1yeD+SY6OEz6tEuY8Xl
OXwZ+fYxZPlBSMjM83NrE0n6KQGm8TSzqrtmrblH3r5lPj79fEO4Kx62uUfrXqO1
09W28wgDMzobx8PoWA1fmz/qzijr7V6cvVia2cJl7j90S/5J8t3RC2xckpnHGD1N
jgYBN/Di48XsQ1Mr0X6I6XmLTMGYgPYbnynTflFAfFSWuqf0sWhGcoMQ095UbK/4
9x/g0Fpm78LkbbYZjupn5T7j2sCy5RkrCvMvXxWJzoScnlVesLPnQM+H88JYCpTc
K/LpF8cRv84NxcJcPkOGM6dZTzVCK80jIdS16uP/ahjIKM5z16np5SJQiRL+03ZD
jJy6xI8fGz6Jr1TzfjCciov0VUbMp+lAHwd5OHCic27o0S4WsicLRrpCRXfQ2gA0
wicDM1MIWh6uBnx9ZNOvaDicYNNOImzFoXDge94Ha0S7X/+tFR8HqZMLKyjiKh41
zW5PUEj+LRjaVVnRMBUTmjCS7GXP+uGw2/fabyrsdUE3HqXy2ALyozkz7w47+qVR
yN6DFPnjHxBKK/Pwibk8HuSN7OqfCMUk3Lf4WLSDauC68GoIHcUWfgjSILwCPUQO
/+J8/3ifduDmTUJp4fv7Xse/vluXyIp8RdJb8k5mr9xPcunTLU/D8Cd1vT10oDxH
uhG4tibsQvWhifOV43qq7tuYNi8A/yKMVH4y6auWunEVShGfDc5QGoaP3TnOx2mF
vTk6co97KmoP/RWj7TeN84/+Q/A4xGy5Ci8KZPYAKoTQpOVZNwJ6HCP1a3yqNGe2
bEApEWGrlhhXBi7TvUr1mUdXf0p+ls8/GrRmeQf7J5hihyTyiWaK281xqaMGGDGZ
BgyfaeB5sGC2Mgy4O/I7otO1W2TwTHTpfDptmBje6ZNbzjs/XfacibdGeg6h/UrR
AcEiSrxPT4x+smn8fKeZ5sFPjDGwJL8Nu2ZXGjkmmBmk2zs/Ziu42HgpimA6f3TZ
O7WtRl8L1h9M0AJJXcvI7iGbXJ+lgGdJL/JbDB6he7xWqAsjLsW4pChBSEGkxbkD
J+9xcOlrp3sks/W36Q8jwmO9iJJBx+cKxQ4LoUVJb11c9Z1gQb/kpJr/UooCd2qH
KdqGUy8y3yITGvjh3twt0mmFtRUGG4XHlw/36TJDmiel86UUjUNf+5sWaw71BnLG
P/FsEYkIzbYknwWE0PGr5CKiBLbeuct+zyizRHHc3AL1zI74L4xYEuGWvQPOCmwc
fXkq7DNY2WTjtmtY20LLZ7R9wWxGwFvPUJiT6NsYsEgZiAkNR+WlmOqynS5qF9Uq
aXz2d+I98HFcXU/6wrzG1e+EGPOomMz1iLERzqXRaYlzUZL4SaWD9cLQ8t4o3ihT
hkyPTmlXnuWu3Xa8pgfbq8ioyEiea8ppqaIz6pGODUPe8IMiQ5tApIXKoLzHtkGd
yC2Bz2DRkeHHVZxz43OitQ91mGXFs4aLD4cKLclvDnHyMBPAu+M0PlMvNh4rcY4J
p+pXs74D+o9oxlTEKXNuMC4JHEp2PLggFh61bVFm3HszWOfjPRKEnW1A+L+/ZG4f
`protect END_PROTECTED
