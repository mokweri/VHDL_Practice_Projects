`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6f79rsUIuin/KVav5X2FxlpQXWT4723ADRyOqpjbOIjXDlH86V9PNk0NLPOrmRs9
5GI2bUrlG9ikiZKBMaDCwthqNLkRRpcCyLM7XT1jqVuaZZBVRBpZ2iiMxlWdHHhG
tspOdoRKnfqDIfEuZu4bD3aL1jbtlZFQwj0gHGX7HKkD4BslUJXYGx7YAjp1Yf2m
cPJONxS0DcRvr/pssMK32XeRROF8M097eMpuRmA32yytNzjy8+l7GiKBHKt4zQ63
emrAidBePCvICyu/wFvgUCo4vRyWKY6V74Y3Qkf7h/kg1hdIBnRn6pc03q3IMIEI
SKCUUyijPb04eU7ZiZTv55ASTLMOoDaA1Eynr89SsYQWZJh3xLfIr3EiAn7CZBxY
cvd5UzR29ofLxjsA7PXD2zGBGKEiEEBO3P9b8TWOyr2wYu6hqGF/WmzFdbujXFZ+
vkHFmFWyPJoyRpH94CluwWaDt9G1PEkZBsF3GxIt0cm11JVKyiV7tR4IQIuKIgfY
/vXtUVjWcNzT1dzc6C9wE8TezGWzzYY1ylOrlV7gdz3rbTk2WzQf2nBshwEKpVC1
ly7Z9679qeKSC2PtZTOkqFXhvWBVc46QhmVWONFlz48W+01qa3EnY3pys/+N/2n7
+JIUQWke55dzSt58ELzY10ijVw4kW5r/ReQsYphztrGKajR/WfG85yve+9AUg65c
GPaeme1qW6VQSfW92SGEK0RuWYtfznLokGLI7c7vnrV2Z4AlZ7pDx/hzhYSTO+b4
wDna7LUkYl9RbgmqfuF1aj+VDq44lkLigHXBilTi/RKq0sBR3QdIbHVhe9RexCKd
zVjTl/dBHTsNfztBdtevigINbzyAqC57iV8DjxR+9nE7+8PxeGmJsQ9Q+PhxL6UG
hC2JnSlVfaqzSOnyuku/czvSFDeRes/t6zGp/zHfIGLHCaXgmAN3vcqCrCt+SblO
qxbCsVUd2ZCBs3obCAW2Sx1PvkOghvnNUyc9OyBv8Jc8W4hoq7hpP5r0XLfEWTK4
r9IhQgVRNKtt6HeNi4SHdn18fjBYG7Qtwwk1RD06yXszkUAfdBnpOvOTndaUkYwy
4Hbvgkf/mgQjBBVtzttidCjKkBfNPHh6xQYwbhvPuF/grPK0KGgHARRQKXvGRas8
vV7MWUtVdzSveVGVy+hf8t12Tm6zntLub17g9AEzIceucbxr9fR7IW8s2Nyq5Bme
7mJtyZrh5TELuBNtFpfg8qfmPx4XdOnRurupQl/IiJXE9+v3/6Z1p9nkufP1Pd5s
cvb0bWr+jp4iX/Xh3OvpfvI71OS8oZZGJtgmc9cqiUAbJiraV5S1v85724dW3X6D
JtxAOq5AiM97kYlX8lARV/R9u6lPj5yN/DnWmo7JvL1cLBTIqSeJeUlmQo5N4NYD
ByZkW7HDHjNZE8qn2c7yuYtiAUhHBbUgc38zdTZSoACrz6YBfsm3H5NI/CA0eU8Z
W4Heph3Z+oAxNYN7UhGicF5+BPmmPbbljqxNVsBkR2UJPK2XMowXOPut2JRWg942
HYtHLhGBM4U5lEArB0+d8w==
`protect END_PROTECTED
