`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ss7DQ55ooa1JicdCARXO8tmTrAx4ebdUgfySZlLc0Uwei1tNRp740ED70E6HdZKp
CI8WaHqjW5xzbSkcwPqnJuZ0j82Or9+Ec1zoKFW5Vo5KLBngEse58R2DMEXELgKv
cAG7seadC6rLv5Mehip3Xs9bF53vAniOIzvtaXCiLI2T2WQY7Gv4dMDZA5IIeKAw
Q33z78JCY6XUw2+STDyaDp1oSPibFJLcuqml7n/Cl3XjH+vubuvChcxviFyIZ1z4
nO4AYYN2J6QXZty6TCTbxmpRyW+BI0ZnC4oZPLf8XnuGNYOo+yOeDD4jJM8KaKvd
9VFfY2gYS+/obj1zzLn56I2i51En1Iar+CIOFfv+uuUrNBQDEoEqq+j3rMKEm8Zh
C9BPKSzGJsl3etA4TKFi21jkUVlsk1tAlY6RvTDvNUiKxfCN7JmbaMp/yHdnDT9t
hyn9VDl/WyDKeHO0PidEh/pTRnO/d5/ABpAIrUcAJEFVcdNB8CwQurFFXKoNEDH+
luVDsM2y1SZDvkWhww3jPkyhacCN+PjsX1W7+nJ0POb0Iow0KQCJ29fiwpA/0CiT
e3oIT6fwXlBGvaNyIEercImwKMuunTPMDC96EVUquGI/NcbZQWf4LpaBvhysq2Re
Z4xIwCSekl1iQPqhOVpn2PjXTXeSH6oIJxj9DAehM4I+gS2kbDSAt6/gDw5AGdr5
xnnfUC0+IKykKw/512cnLGoaKMahycEYxo0iIrq58eedtBH9BAl2c2PMh5y57REU
lKXWJTwthuCbJ2O2ZXCqenIG6z8Wm6o/XyeUic5uRuELg843/1zkCFt9tOR206C7
hBrWf9wqoBfn+ot0+MZ/RyTCrv0GPiFxUoFWtCIWGgkeyuNzNvr4U42mw+uzPSBT
`protect END_PROTECTED
