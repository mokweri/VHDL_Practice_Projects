`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aOuPWtusKfmyoM8XvfwK8H9oRoOKQThbHcvB0JwnxtndhmYobxz1OM6OY28VbAUo
n1uTwTMVMQ0geF/8r4N+WcdbrQg3YZ3MsCf3K9M5KAdN7a7ODzvvnOUPtDWRGwNS
6yw9wnY8NbezKUY9slyOFDdVrloSx/hk19inZKZNn4FqSHGw+0p1Leg0WXM/idv+
xucbXZ5ocNdW6mUujhQeo8nY9pQrrBTYrzxsRnsH4Par519U3Uyr6DFqRyzwUd2B
4QpGEvJemXgCnCOKaPlKddH37B9fVIA4v/ZCZNoFI3cF88PWqPKFDm6hdf6ldW5i
gKmbo0SiITa38JfSHdd9OVkiSq3zWhj/F3UXATryqiwFTD+5KhsIrr5HZB01UWxc
3ls0QjxnlPWeORRNERN/Xgbu+Zh0QWIfrzShs6CiHqoosaf03W8fdZtufbAhA0m2
+/oxcU/oa0ycP78th6WSXQ==
`protect END_PROTECTED
