`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfcLzd9nGxnB9gyOWf8am/CI/j/kwXbyDmilT0DGE33N7ZeUTQT4aIaoje1L+IF3
rNeKUErqpj9FEFwEq0OMVKPtAhuy1XPOLN1kbxm0C49MU83yJJCZ2YnD78qPAK7T
nMuUz+UXRTA9t7yU9ENpyREYI5Gze+tkG+dNIvLsxh5k3wEyOiQOJ9TL4H6bDapc
6dm+IO2pNzQ3zOSgJ/rVbUmC4aK57gDNZ6g+dgPU7E9ofE27n2IVOUd/L/ROjt48
HZpM8EYq2JqinACHbbpqGFYBwEciQSt6P82E1HzyYG3h+VviB7BeJSknhX8P0H4V
9XqllC+p4srhpjgoFc2ZoRoXKq93cG+BLOPyK3NQk1DsFaywckV+RPVQ0TAXOznC
+nPRaqhFzfXc0Xp5SokopaPiTYYKUxJ/CC/0oXCTJwpq7LCLPDStDXgJ0Al85o4/
TCgHo6zQ4HTrsYFaVii+kIi8yBBcnwqMFWFRl9rueG9kPb9DqtS76jXXhE0z1vUL
hIInoeS1SpXSbrPKv9vc1jSIiI+I7o1gnSJpGB9pYBlKZQDFCgeo8QDakbDuC4VY
uxzsQSrWwcB/njVjRwZrZvJVFGGYoV7fcy4oJWySDKLk2AauKaQHVZvmt7dV9RES
TUmBWW3pPjhpjqwbA/bnRuYxLH0bHk6SudAnmPjO0v9YUBrkDgPmW1BX/YyF/r4P
maZKwQtDoE0XG7JZu4dlG3xglfUCvFAg43M6a+vhthGFZxc4AXI1GdiaBIhHKDaI
A0ZnEhgTrSUYOsrS8LKTF0Z44+nxhCB7VLpEGfGur2819iwQ9WJZByqcBeF6tI+P
8mhYWq/Nmkf6wCdZWJxYxAs6M2TYtK3XCy5y3En/NC/V7yTZjw0tfKyc2abvXyLQ
v1DUOwNWR8Bouw0KIPY+LpNWqQ4ghR9uOfHsR1RsnWyfRRafo6P1AsxVdZJ6ThBZ
k5ED74ekGG2qwTes8YuUxcYyWn4zk5VeMYKhN7YW0yUie3GG7Gwn2I8mBahbuIK9
N9gDXLAyQScOzjgPubu6FxjEHEM70J2S81XwgnsljY9wLK5QCxw/HS7zueEtG9wj
cGzC00Y1YyvRA7msrGd4FJshuUZQzhxKK0nh8p2knBZR4zEjEUMue3gG/SBMAeAh
UpBWNBOZrzHYEEiQ4qZfziF6f4sBBvo1uXEOorwBwnzoh7bS7C/ACl5GY952MwSz
4bLLU0NFTg1npT67jfWz5w==
`protect END_PROTECTED
