`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RklzotPTrVe8ZkvTUKmpGsfY/EZoOj3Su1qTwyCKTLjPH2EwLGXZc+IW5bHWiDiV
wxxzViIhRWMNsL9kwieZRSbrU3Mok+EsE1ati8eLFPK31rO1GTdnA4zdZcgGNeQh
W69n5M2dJGL8mrsvaTsBkXhhC3wtDSbX7VKJ2xKiHX/wrflZsYNp8v9DxHsIAMab
5LSkuf+XbsJsHnjWapucufcRaRI3BDjmNJhm0y4w8xgUov0bCXYWvN+HAauPxRVn
LZx7WGI6UCkfUtTMGDA0cyPX7Zj08TsE9zyw0gnCo3b/ZDpKZ/b02KxkIYwRk72n
W46A2+O8/sq8pPO6KDzz3mAjBFxKnu6oJ/gQa26/ycB0YfeG8S2pGvmVEKnHV8rI
HdCT69Kf6bkqXkb8FsB4uA==
`protect END_PROTECTED
