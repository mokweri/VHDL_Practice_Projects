`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1EFblc68uLD6SynutTSHrtqP1w2ujbeKqcADQdbDkrmcwKzgfM0aMCrNSmX0ocp
c6S48ojXQIdYVCkI/hFYiplXhyBKIUremqZEADXZlp7q1AEGdkf9CPSSN5ndPAh0
HT9aVpz/4GzzjTXGDbrXituH2nZdPgN6gqUErbv2M2/FfZx1w6ByQij8ioNC3us4
5kKAZxOHK3qcjy3BFkkV652LLeYsijQozmCB7l73iZ9UoSh4Z+USAQ6A74GVgvy3
w0k7Ys+jgpLElgLrNplBVMoE1A6sHZjN5ITAiiBS5kHxUiSA35SanX6jxADLL3oC
Nr4D3mvQZpbFxiiix5uH2eHRZYGKf8USIwfGFhiScALs+gzmZU4cl9vjBH4MC3Vq
Z97pfSpf9If4niIuuJJUN3mT+XOGqCz27+x4D/l4CYeQeeWSAY8KwuPWvAVn96qk
3IPNp21V1nODeHiXtl7sfKeEC2Lk8iB8Nnlj99lU2bbPd6cWWWMgLsqYoaha7W8N
zp/ow62xPdFelsIDFA62QY3J7X1u6Uc4ITptwUTmkBuP7X2jfECyVsrX8X9VWbhK
fhRf+X8S45ldYNaLdptUB+8ho0UFVy4xGSoRZS5O/PVMTw6LhwYS9ySkPL0RYrph
bcUKSlsSiaKWWnTQncI2ZCJCpnIJtFAMIsVW5Ud8pJDT6xgs9jiyS0qMunJ7bAn3
opZ1hIm6cR4D8dCqUyeinRqGM0aK7OJ72tWR4Ydw6RS1x/ceGmmb1jGt9QqSZBq0
lagftbEaUhl6hnsJeNhws4vJcjOvXQmZh1i61AYylulUO2PV9HxnBcD5IPWkA5iL
Yk9mhf81qKIyUjzMF35ITcjiWT1+sfbiiegQMZbqcFYcJWx7zzyOz1v+OKj5kkG1
towwz6JrpnTGwCREdXbZUBAgHCLOLOjRtY4B64LzzSUNvl4FrcvOEuGPhhs0fVCk
J5EDeegHclUlxQW6cXJ6k8T0WjvAmujy0ezOxpwBDDGGqBB0T8xro6zi3sRDViEn
WhKYwTXv8m7axhZfC3KrQ336M6b09KYzBNBP5dNlzTm7HLoOQpD1MN50QgkL3TFX
mEPnq4Mf/h883S+aX/69eOHmAfnL7xiPf7SMufmYx0yIulhCBxZqD77lEFv5VnT5
Yiomg+On+XETVbvNbZB/OGgdsDXD+jAErRjSSTCe7M6vF9IAaIiDX7YJNeCjNAk+
+8HIiqV8ChoGtVvQ0XrL/mnizst5bROsbmQb8l0lV6h0VKzibkh2mnUae4LeqaDY
QnTXY7Vg1rHQMAO8DuD3kiVn6RA7aod4qr7Dv5XtOcw20XEilUbxKH0ycplVkbKP
RT8Ljrl35CzyHPD1BqJ8eodzC+8r/8fv882qwF5F81w4AmZYN1NfZ/9brYsK7zLM
uXyN92RKQ18qAUFY9xaT/Lcl9bXw4h/9dgnyjNb5K7PPoFwW8PxeHooJTSOylHhv
Vpkldx2GBWwf0zwjXtkuW7yQT99VNYwPW7Vd2x7B/RQ9YcFeji85Iznk8zs+4KLB
dW3XnqTRLXa8IvjXfRW4jzYdiLQ6yFYEZDOhObAqVrUWkj+P3Vi6UV2yJ0csBj2T
wszccwS+1hPTW9Rh0rylaWbpWZItWR2T0hK1CV0nWiMNZASa5dZ9GLbcysExUf/3
vkHa2poP6ahqCFWwl5uIrOwuc/Get0qo9NWa59WMhJS9xOocZjn5CJ5pRXDwhcMJ
RsD89z1T1fpp/Fkv+g8UX8U52fxlKRty7b5HfbPOLtjlVJM7f9Q43uKwnUJLwzff
HEWoCtqhYJhYPlxo3HJ64QxKxsh+EtzIeKWeAP8m1ax3AbTCumw5V/GF6hEemoCV
9t8Xq2F/Z2i6qcOYT/aPfyDQ+cNA6Qhnt2jhII8ZqbwwVsH2pNW2S+XA/nYWGd3/
44G4U6Mo3j7BAFFgbC4Kje1bFVKPn9WwFjMYddf6TEox8YufdES4l6j6Eec2PlRI
8YwNwjnj4f562J++AdBAyhsW1GYTiTqRZ9c1eAcYIAhzl4vPtJxz2h50cjvGqSui
ppn0iFoy+25a4phVn3G63gkglkLUuLmVlc0HaMEpkiee1pg6Q0n7ZI6iJEJph/KH
ib6XwwKExciyhKmymp75AHNJLwyuiExXsZ4xrL0WtdvQr196/ZX4W7nMVkCDcVAr
WlatfX6ovvbdc/6w3vc8Lxqr0Gze0FzLwtWNoJx/1i9Hpx0BslCUX0/mAqL9SgCq
8h2D46+IGZ9oa5nbUT0pkXu34BJRSVFpzlrkUkFG5XjXyXUkAKFp1UKBcLCUAte7
aAEdX2sAOjhkbIg4q5li8H4jwjHrvwf7NSKSWXd2ljSeyFQHtQ4P8kzwWJUPJ91m
LW1S7N6zyZ7jPBkgUP/koKYxIfGdVl7GUEYS3PIJ/07xTFjrn2T+ogi+xzNdZosp
4iVpMMF1+qhFyiEFaElKREv0TYBC+TjpxXmtygZzNyzGJ5Eyono04LU1SNjy66ya
UE4M2OF8Ibmr5RoJwu+63kS+hmRq/UvxeThFiZ4CAzEqsWAu9R08zQHfU3HH7F3X
odjMzWfRGlca8zVR6TXM+lCBBVl9IYCe/rlPa6wCQk5mizaPw9MZWSasch0np2DB
Mv4mCMypoobyqtZfx5Pe+4t41ly6nPSn/zqa1mCBWHPteABlFd77oQ7v1tJDLdMg
bHklyigTyAMlfcs84lEqONjJ7NyTXm+qxVwa57vjoJaw63QeGnRVFQWqBq/JnfIK
C7QoE1GyoCBgNTPAJGXxOZiYGpfyaG8+t0zDylwU661HvZ4Hdw5AkJRDPFjfK9yS
ERMFubX531XYSGCO+JHV4oErvurMNMje2ezWBnFmKwl82/ABkkcAA9auls483Yt6
vNcSsWWGn3GwFbz//4G8aHJ8UmsjU3y2B6ih5iwOkoDYb/QyUyv8ooiXD5p7YvHm
Acll5ZRr0XJDAzN0+sm6CiNKITLEMgAJPI52u2sqxiTDrs/z3K9EUfsEVKYUL4Vy
+bgmMXPgLqG+N99SaaFzGZi+MAfeVreBlofSWDGs1OhwOsoJUqVCmoVnZoMMmqJz
RG/PR1l8GqjTHeICA/Zo8oUO2WBFQW1XOYw1/oYlxAamlA/fyb2yOA8/OH5BfEbQ
yVr9U7ewNibXjnD08BKeLM4W0wL2hWBqKYXX0Es7iLZ0G/bjOsWin1QrBWLzWeFa
APf5mjVtmo48W3E26qAVHx8bmqtaGB8W5WsUJyP2xmunl4P3kVg8ccrOLkUF0e0v
wenWOgMOdufU3doz2Me3V/gcL8x7nfkvq2QGgVPzIXnYXrXsx6pAV+gjxRy80tDX
NWHyMR1uQXGy0ChZZeGI7SQWDIrRCPn3A7lDTd07dljdo4R+cB8IwJ47yk79uaYl
i/SeA51BvknwcW2N4gp/oUVYxT4bEAAxNlIjlh5iOfdqAA06gQkfh4omNL/kezSj
ZCRnzkdGlv6Zf1D/VltkPi0PffGOhj03wdN4e9jn/6wRbiksf9H2fIDEVFsxfOv3
RJYd/+KmHzw5gNgF3Cv8JvtTfY/bVtkaXKOajtNBRiG00r3XF3JOa9rvZoglkzcl
iK0ScH7SHt4HQaopkpk/0J6HjAB6vBOzI/qqEYb+Sya+KXtTuScre9fvVwiQS2Fv
rSgQ9Gqy7pLqt63R44PrjNGC6Ngd9JUuv/fYF7p0UcFF7vfD3OZZoBuCGF6QWvIf
dudpPcTo+ECZau7Yf1bNygud68NIW72K9MFJ+ckH8yiwuaJcNAt5DbHOJfoygiSg
ES48K4y+H2F5z+PJq1uXOZ+eJE2NSFPMAFdDXfwm2GSWFO641bp8b0bnNB6Xo4mc
H2ph7ASHV+T089C0Qun9i9h8h3NHv5uEtBqf/LQor9WKly8m4dxiNXTB72ag20ta
3w1c/2syaXEdZzIxlRzv0s70I2IvDx43GkJwz3BGc/zCIHpG7OpfEuiQ2gQcz9yR
6X7b74PgWZeny0QOtuCZanFur33tN7c5aVqM6UdsSJse2+7xOpiQ1NV9p0zGoECk
KoKWQoh5bwDxl/Qi78X7jXc0VQ3w52cbYrPtzIC5zPgOsVY8tELN241FAxqrZa2V
ogL61ySUAbNOLS93Dwhi56RNDLLL/oJMd/OEA0izR58Q93w+YbCbWE8v8VzKUx8p
dUsgaBY9fm3mXS4x/KKxRkDlm4sE20xQIKRg1pKVgoI9BXqSC4dM12zjX8RLbl4F
BjyS7POnQAlovWCi6qLORwpByv97SCMQJa/fu0QXWVhainpDJt+auXO/bVIPOH70
U4InBxndLFxpxeFFUk9jNJXbHvdWd7xC0+fsBGyzo0hm9ITHLDBX74LFpPolZfmZ
oKfJdM6g6kqqPO0mK04geXuzwToSMC8kM6AiSSK+VHJtr1yVjNjbZtFlWcF9JN+u
AcyAT57rfDP4Gvd319rzOccXX9NRnuiEGWV9ydD3Er5i5noiz6Q8nwU8VU155LEX
e1I3A/MQ49rynoQVOiv06z3fC4J2fbKx04bKCu8FMuFmermgELvXSOlKyJbyzg49
32fGds6e2rwteyGbPUC478v6eGYsCslcwW8WmN0Ed50bsJnxjp5q0Nsstf33fEvJ
NjgVCnwWi7jINADCe5c2GtE/2C6IRqtmA6BNkRKOg5iTfrloEonLbgEur0S/mJ3w
N5fUD8vZGcFuxlg8M2OklQ0yKEj5bqHj6guQueBiid19yviYiKZjtgWM62nTsRoL
XIlAP+VITgO8n3SlY1OwZMacAkNBUxF1SbqoIb6M/KK1iOsCpaq67FLQyB0azu4X
orghgWhWH4hA71485FFG2muuSEE9nKHGNoFaSGXnyG/uujBoP8RNHXknKWXuSsdY
9j7SWjrATe4eDndqaj59xrxuzNHoFuUND+HQmQ9r9tFni4E1l6xJTUr1uk0RhLK6
UTvqHBkga5HN71jIW2bbB1snfHUGK0HfRAB/DUsWDdN7bdc/HP11rDpficolK7fC
tl+DO+KhUO0ApMPcuO45GNCSUfFvR57TXuAojpmI8rPYkGb6F+phXFbSohHjgwlN
7UJl8uXsuTlGM+mvvd3hm7vPWO0cPTjJfJDDRsVu8T8od/4LBM+YpTVZzoLPkhQu
LUXpQoFhvfM/E51hBU1P/dJzbpoEMNd1N5Bo7RvbCfaxGga5mn/QeJAfXK4v+cf2
o0cddMn4o8aelWU+X/kjFFH4hHbjVonEjnsjf8QdfJWtsKDs0KWw+ug6VMSE03kv
k7QwT8EcMCzU+uKjCOI/7OppRyaAJuxzzZXj6qVXMzMVL1uRjezRJfEqmCx++F9R
0j1R5WdFaMMsacA+SrSx8Y5mMD60ApEdJK+AP1c6t7HHAxu4JTgmnrAqPtCl3OCa
k31Mn9+XmNA0nl6RFPuhBLFjddW/zapd9wm4gRnTvn3/Niflt3fYvMQpxfTCVFxi
ipdd1NCf6A+1BmX+fl6tLtP7qg4Pnw5ey0MTJsYFHnNPmw71EThqjhSZ5gTQYAIm
XfoC0MYRZawPsutiQNVPDor7SrQmUoZIRJhxejGCWOI6wWkV9X4GjNKiN7oaONNF
o+poYswthWnajhwUjIlxRQ5O2OgyrYX01n2xSJSs2GuaWQiO7BQnVbeYIPvOEOZf
Pu4olcykchRkTDL6OnurDrqtga2BrYQAZ6o9O6EwNmD6JNm8QacapKFF+PpR5c7B
4cx5AJYN1S8brpjBdpI3DtzAyF4vgdwBvNmJeegGBjDjKGyi+Bx5xcE8eomQTdyj
a18vGcWQ/lPCE38V/lkt/aElRYG7LHoWWnVbJ3IeyZiafwrHiyedrxBVKH2PvGoV
MsovQpWgwUbR3MDoDUL+axsWxZuk3ZV9ZpB7JEPK8yDFcWagi92vA7s6rT9wzHeX
0w70823gt9HX/8ITi38MHG0mOUgVJYvhPccXFt6VSGEJkwbjsYKFYYdUXdAQ1fNe
/DCISlDSboSJSTCKJNHjob1M2eYaH4Jq3+Pd7rUrxfEaJS5cRbMUDNllse0LvtXL
yelFhSncIBytNe/Bw0kEapn1fdxq1ce0JCeDp14mHiFu1Zzs4SEXwTIAt75pan9B
RF/IJp7OfP1ZKhRKjOXhOh+rk0fYjyHJ+f2h4bM79Lk9wIqTpu5KaMGlY4i8l1F9
76YZxFqD82b5l23fKN+jnVliZSWzEjQ/x12+PzAqF+kjRg5DZboS/+mb1xYQhOKZ
ctb0x/hVBi39H1/a2hK8O4AU0Eb6aYnEo0/a0HhkrayecnUfheNeV71MB2ejKPtr
lXY+oZrwxekFGDjChSCgWsnsgqwtG/xxyUUq3ktaALCHYDMqWlIHW9rn/3v2PB1/
UgtXJc/zff0DWePx0cm9S43k/Dg0lPqu2OU4H9qAEdHppz4LqMJUwSsY7Fo/9mLk
IHDMKENsoSqBQdSdu2lp/q9ogVrNJn81IIMABZHJI4aLhoX2x8QO6+8fX5UjlPGj
JvxTPkv9dn2Kl+gxRCgiM/S/8yAjAL4wVHCt+9uT25NWpQeI8ZFGTzpyr0mHvwPR
hiZFOoHl+bwwDVlNz/97Fj1yXkUkAq4wPnVqG9QbuiiRfp1PE/Rd1aBTRgP7kvO1
IdMDBEztumanFn+X8czGusk+5GYJxww1ZskriL9wQZSQMWRa8LE/bL+H0DvwPSxt
CPsFrs4V/G/SvvdRWxiPLSM8nrHU5gpP0mPi2ql8sQaHQyaBq2DNBM8VsA1vasUL
RDlEIK4lOALzbIpMKcXR4K/2ZBYGvbmsL1zKuLfERv7SOVo3dkOhQ6oq29gBu1rx
M/zBG9jJnUFAaO2MD1EK2KWbvSkFvJ3/M3sAkIC77RdMsIOil5NPemIrOQmiGS0q
vUjCax4jsatIEZcSXfJQ1IO6Au9QoXEE97qPpE3YfznFqgxnxeyHOAEWVorqR8Id
D4bZ5QzmZp2IZR+jP4iQH0A6OscmOKYuzFf2ImDCmdJ3R3yw8gdiAvrW2LN9tpnw
06YZb0syyCA/3g76FakDGTDpYvYadxBOeyR9KSg0PnJqR/KNooNIPVRwzpCG/cWe
x0aud8CVlPcW1JbEaIwFpP7pzba+BPyiJqJWZBAbsaT/PyN0v0UQ6mzv/iZ/zMmf
e1srKgYG9sYL+m0NsFI5W0g5k3FRmfxm9JanA5jmi8OzN9kXyHyS+ao+Las24jM0
s1ZVkqUODwwHC9llsP8ZnaFFHcacGgWDkkdwjJWt09MzBRFLktbJMgkbwMl3MNPh
PwOLwhPmnH9+y79Kf9kbRtksp/SqLQbkjDBDOfFQMluHrbTK8DmlnFaUKV14oopS
S30O52GJYw3xUCuArDE65/T9vI8AnW/isjZQrKBu83EyicWXpVyyEzKYgXcRmfnh
giZiggBHJ96UsAweVoBtypqix5h9KAl/36+hWFTDxmGJ1r4mm1xML6fq9q+ao6gO
6B7ZHLUHuQ7K+6VM1oKFsEcD78pMX8c9OVpgIB7WKY9iIIy2Hi+xRcFZDr/uT+4U
wPjHsR6J+nxxbS6I1TaL7ET9bRKib5mr7sMScbhvKuadMt8abGKA2CEQoVPcif9g
uyhB31yvmK0hr0gghz95321wylYUbl0qIRbmPo5ITcJ5HfC4/6Uai9hfQbZrtupJ
/OxU6iYPkvlv+XVa1zGkx5V+qoIg5hsmOn8AG9eaiOavqA9IwT1uUO0CH1s2QWYr
lVxeNkwBuYWSjOqwlauA/0tk0ZIxIzZ3E+Eq26FDcGpPDfjlOU2kmMShFDNlvuhs
MODbPyzNirsqA3fpJfFYyg5KUTmBqO32J8+w/J0CFpv9lTyIdlcymag3GUjaXb9C
FG23bfSYUG2YJgWyQabXuwHIEDWyn7LUiZ4yaHrmy7sL5xFcbFlzPghvXnmASpwt
IDGL6Grm5uirMkSYpxqYv4lw4LkTgAeS0kzI4Kw/0kdikuxnPU3IbAY9s0cfShJm
rlvraXbYdCfqktjKVvFuG18U7ovC0z6qg7Ap+Q+Qn2PQrGEikPvn7CQU9P6+/ozs
ceEiNGvyRSvI5N1GPMbxAKLgxJxYVgBltqcGeCdJUgJsZrKCjlRvJ/eGRHk4heCn
84OBPJWU0LwPjN1zXdNA5L5ftsuuYVuS9vQ8S7p1r/kPuM1Po6eutFvJS2WwP8uJ
I8BpQqkrFuzqVOlQl9L9NwLDiakvnDAsFFgo8CanbpIAO6ms6/JsGXg559vGcFc+
Z5SfjsOVH5thO3RB8Gnd973heJ8E0IRGwSJgEuMo/F5gWHc/ultmaCCCi4zS1ilz
htsQGgfGL736a7tW8KoK3xMmobwjMawJUvY55LjhM5JxVvvqEiCbklnDSXuCrZsc
NJcIFrSYLUi+HOm9xDVB6l2WHoL+uU9Jr5YaZbe/+CXXTGg0BjPNrcm5ELCLYBzL
SjKxIHsHPqUmSA2Dt3AQw/tFK6SXN/FyJe8po2o6MRvS+4FrfrrvHt0PnEjxx4dK
UNyv5BtyCZBYPtMx1o569G/WneJjIYRQ297EEoe5ILGr9K0QG7Fzd8AoLjNyGtpM
DP1giPQQkba74LBWUPTAjaf3Vws7xBjlC9YEE2qNxL1MCoM/LU9de5T4tHeWqfVl
ncyV1PnDpXMB9o7qEnZqu+RumSVC4vXljcW7Kvhs/ZhTwwHnYIoJR5ISVj2fmQjx
ob3YPqKsCJxP/Bev3XcXLpWZRgz0DK4d7MqYusfGFwUnX7rDhqSdzxvJq2fuWS7D
HS47qEhjvdB7LToC8EvkFmlHg9GkAHzxYxywdCJStsXf7jV9h4mxdvCrVKolnblW
KuAkP6amQgGH4gk12XlJbZcgyh3dwjw19Da8talcwgdNFSE7TgfmnremQ0UZoBcK
V6W0HTYlLJglED6YKVeGJTk2o7Eoq+PJ0IlrS9fl3UnuQf58PBpoX43mUTMY2BtU
Pg9I7H4WsaqlvYXs+hSpWEdXK4ylxX58Sz4Y26yJHvSrfExmAwUiFMEny3PqeV3y
29p9fw4Q/LWoUcW0iZHincN5lT+Ca0X3siDFne1EBf10Y5OXbVMElCZ772qIpshr
yxnwJ8dlTFqVQ6489hex/FcRFSNwaZZwrxY+gwmCsBqlHbWVnnghgyHexCiTZVSB
RMVuGFzIfmiImgBYncj1BEYHvK5fCLSE3OxTV5+BoYVUtklvrRETFhagXuE8+ON/
3iQdfmyHsZl15228Ltk/+R/4SmcoPkcy1zL3KLQfzuHjHK4E7tcu+bpsNdy+5dGm
dSBMeTq+9BvJjQR4B0oXo6M/4HTQRE5OF2IDGA9wCLDZAllmnjP/RNjFGAS3iSb1
GZtdXsZi6wS5Rmjx1iJyiEwS6b7Z8oYIqTAqj0sJpty4C3xl70ifvdeV4SfnKWMs
x6LAPSikO50OmoCVK2QJKYSBFi6GpKlK/QFF2OWShqg4Fstq3FSzZATwrD5rJmvH
DNqOr8Imk9yb0ap/82f9KnWTJZF2WmuiEgTzLNqfyvL1VhZWT1wl3BBgBl8AQ47p
/IbhFbignBWv30EI8Z8jAOnqZPgiqgNRziXllo0gjQgAjE1WUAToO6G9Yk2t8gRC
IF+ecyLx3kOeAJyV0MA1aTj4Uf8mgtanIHAYuZa5//bxLuaXLwtu7VtmHyCrxTdN
KxUM/E/UJDHHp08exSZnvW+AJf+qnKigfqe7m7X68p7htX/zSlQFOZ9xwc5fJNlY
9xFL7cn60tbhmJmkYvvdLiPe1Au3KmnhpEZJXGpXSwxv1DToctU0PiH7Qi+gQOtA
i/h87/VZAe/bq6rWFS5MuRDrOfAXXLvyh8eIM4DXO6YN7H8e3P+zNMqn3Ri+kOOc
jYmf2F1DxBUHTB9x4h4D5ru9EFa4ghBRTQPmNfR3Dg7JOtrqe92mE16KLp/dzNh3
3A9BR0BRNOQ1X50k1lJ+iC6QQ3Jt5j7ff3QDAZxK++nGlgry2VvWqRjVrKjugSJj
5EyqWj/YIIX9dDFL3h7OgBTNRJdpfP/uyjYWhgCzd159a/H6BtGdVYdSIt9o5wcO
2USjUYcgF1eYX/9AFPz1tuLJ1PWh15PAF6ToBKmoj0DkfQEqWKgus/n+8M+fLzVC
g0BImRYngOQ+nvQiS5wuBhKbXVx0gMcy8NOam2HFWQ6ezAysV9fGKQdXrkh3+56a
EGVOnP8oXWwxh0ayB6kx0HByZEb50EgCo81Wp98zslT+UiwJ40hbzt0vsmrhA3gQ
Pv0dQgZPQFC5o992okDhawK2nNZrmYlP7MynXYkihEBIULKPi8M3cDxg+em5rQOU
YbV6vZsjTh+Ud10RHeDuG3iNebKGpdhoyNBhLdTDEbdNyYJMAULVhlmVgnBHLlfE
Ge0sAXSzH/Lai6L+kfH/SV4zXwvRmNxPTbNvlJAPVDmQw5KrWQ6tB+SPFq1rLpRp
5cgvDqtr85CjquAOcBa4U3tWBEMXb1AFuA0gfg0g+K/fwbxiu9PMW6/kG338/YRt
pwaDoa/TrUqDC6A0BdR2qj8RFQk2ugSUoK+QQJRFi4NH4zX6RA+OzcL74gRDYit5
JT2HFk1Ybyw7CZVMN62w4QvVDkieVjipN1GzZARUJq1vmoFJGBrRpwTtQ3QUj8YM
Mq8ScwtfRPPI/Bc0729txKPrH2ixqmbnpAwIv2GV2xrT5eM5DSdvaW8QIpmpsrRg
NYo0kYnqrBQOKFNPym98cWAaGHurACaR15IxhMNiS9HqKWZsBNkJD2/UMwITUimO
e8CvAV9UF1m+b2Hs1oAP+HCLD+wQLj0RWsbMs7qPVj11047y/v13LjZkyC6W9M+R
kCJxN/vNt1f1vCCyhDeiD4dILpmLa/7dqrRRPnw5uS+ssB6GJPYM2fMlL8MHU7J6
TAX1LRrlWCmVOC2h4PaFmQT36g+wKt8jrXj8TecFXsCp9pwXAw6SomEsfI9JCwdj
sVjdbYg1hHYr+uZituYPt7d/xpdiX0zUwDqfkzytyXIhHzMHWkv5rjyp4SDjQJhU
MlDED+pnyUneViXVUJ9uKZCt/msdM1y1E76XTxp6UTrzRxMHhPFN4njOWoyihwTj
5Kk9HXVnb9m3tYOhKTjK7EJ1+e3LwwraptjcnBRKli7HExw+HF3HNtIlrkwyyzuy
Qdula1hBZJa2WBdeWO8o3uVCi39pE17j9cRYhRLpYxUCpz/t8YDru42UGK8LHKZi
CovxmRUogkKssVoCU9VPe7vC/G1VKxz2tCV9bH5r69pcvcpNeXvZibeOKknPOmsk
fpi7heNU0INRV8sq3c2awKJhKKL6agtKSnJJBWMYcW1/pacj7v/tqKuTeB0C/mt6
tuvFSHtOvP1neOkW9nLiGAsd5Lx0FN7CGsMk9FJJQZ1HCzKGh2uqnppKLRElH63z
GRj3IEmXUwp6B9V0Ant3tw+VULIsmIdgcCn0xyQvlIHhPhbCNWNSU6l26GWTpz0z
8FmlHT0Fu7EzIoaW93zP2IzlwK02ZHrkzn4hwfKT5CB/l0o9yOqHzAK6yVRJS9sX
/8t1mJ3nWgpJ2Rgwi8FVznU3AErukVoT086dSbfe7OD/GZ0y0EtRVvEGziFX/Dhq
SpSkym8Ot+GsB3DhWyPHcQZetRG3pFf5G5B6/GXbRIfvXGGBg5eeF9SQSg0bdFB/
saReEH4ecHVK5uywqnAHS/D0lGjJy5aGWGnDxkMsUsBSxo0kMtxB57XrbGLhRW0D
JduvETxZlvolg5jvlD+l1WornxvgJJifBa7tM+uA1r5mM192nPI3VgjSfdX98Xsz
9upQKC/Y0/RubgHy/F2g9ttqcJMamOJ4iT9lMZH42sKXdR/Q0z3utwc/NlydLkw2
2msedT1PW4pw7ydLKV4xFjU00ZD1Dp1MlVT0/PqKADGCA0S+5FtVQwx7o07anpjT
B1pd9+wOqbpI5nmHNhjAGAjD0WYlSqqTTomI1fvGX7eKahBcvgFPDS+SJXJAyYYS
bT6RTdsKSt64Kn/fDYFhK7uxHb58TUqyIXmfuztqK8H2LOhEgJOZYcYc6KEeNoai
X5AEYlx0XjYTesgHaQG9427iBGs9WQhh2uTcW6rk7psCsXhs3rni8MIaDYpyKvbM
jFSfTe5U8S/Wjum17+x1L4WQt0Q1Og8oNoDu6V3mnj8yeCVLgI35223fH13AKNjk
uRsmEDFNOwChksEDayHgOvBxyFm743cRqw8kRhWvLOT67FinC5+aZuykZHzDxPOt
r+cC+PKo7M/GQydTpDplSnA6kgs50tFD002bua8mwiX/mD6T4BZsWupv4HScD56S
0MvDKpAdRsokj2qpsK8wgtMmJ2y4VLZGV/FZ+TyXMvM+kMspFdrvJgfMQEGyKq0A
fjfYsJN4h2oNzDWfJmLhjhzpbISeFjN1DpAlsCzY4+vg4ePspGyASQYSp35ZPzmC
2OxsJcHPdJZpaoJcUiBKQZqqYazkmzwr2X1PqFVuVIHxWnqJAaVUza9ltspd5a1N
evQNnhIw5X6Ib9CU8EgqAOI/aKWfkNvhflAT43mFt/NPwxmclNVd3wohJOUh+Pcd
/OPkoFfqY6XdFKYgZbgUo5q9qBLk/e9q60fq67pl7DgaFP9mwOvYortQujwHAPcm
APHF5dN/wwg3hYURaAsoRUQ3uNUJ4odj+nKjjdWqJykWB5Lh9ZR1UvjEPy6etxnF
r6HjI6smgxFqWL268ZZnclTMyLYCBSW6bJS0D8zPV0VMCB/MW6WTlBsbnG6Un23y
kHt8uMLimlBj5shVie4r+z02Z+Zhou+WgUnpgXzSjCKZMt6tZzXInkp7xndTu4qw
G6tN2umwajmodDxZ8EjqHQZHdYogtiA/1nC+/ZrczdQmus/8TEhNMeSg3R5z03DF
waQ3y9H8/+T1MOPunWpgOfC6XIr53hfm1xm3z/N8KfuyTCtGzxLtjLjhlamHHQ+v
07jSkN92dBEtpB8+BvZE9cC03e5A825PHoi3MtdHTL3LeSGj8G2z91MVXlPyUZ5m
e5ew1BaxDbJnh5d0pf6PExRNtLdIoc2FHVsR8G51533lAeqVtfRoBUvuBxt4l/rU
WuB/cGYjkDGeSjCrCf/5c2MevW8VMLE7nm9SpWguxXjHgejrR41cM+UT4de9g6s9
5YxkfT5svKnChrOhXfei4Y5K0rFFaPniwMwxSZHDseqMsQoOsuT/TUaQNdvsu+dt
rBSPejG568ey/G/U6H8P8uhcecULurARa3LLzDobZQW7IMWO17/hOB9UEJoazny/
aZ425+opUmFbgrDuPSGEZ92wlul9mTYJlDMae8PrQF6ef3MAxeHe1tBI06o5aHXj
Jtym2ZvyioZhQU1xIXrVCmlpa1t7Tdn7Bx50AslmMnqCZnq/Bh6wxiYri0t3+Vkf
+cq2/tRu2dRIw3NeP1KGnujNmcaCfQxdTVeChvf2sMXHTZVCj07yx/n1FY7RFF61
GgSm3esc60RA8V+/QM3x7Ctecekv389tSh2+eBqN4/e1j+LJMXJn36JIWXzzz2My
lgGzbRDxSw1/uds7/AcPMiCpBZVoIxa1uUGbDBJiFxOkXWMCcwwjCKCRFkcipDvw
+frrsWh0YfXw/I+b6c/yc0JKjtVn+oUaEFyfMtS0gy9dSNqqrtsnFIZnidVBzoB6
zZ/Ihk/omeUpYx+EqqLlQ6GYYFUsxg+Jq8ii3za1tvypFBZ5OturLWCf66lSGwKp
poA918qReZ7+uI2p+L7mCiXG6t7/KzZdlMzjqoxejxiNvEKsbvxKlT7xZX4n06QS
3BjTfCLDJZwY/4Fzm8LU4GBxSSUiZPOB8UDRBZhFdd1P6/H1kpahM1oAOFjgfKRu
Ul60/cgVccIKWW0lbWeXfDVV7nYSR53Gd+HUYqPncFLSmifF7RH6PP9qGFTyTLic
U/yFyPxUukIUzpj6X8Xtlj32UzykP7fOmIpxy/CAvpFA/uCI1fremHsjGaHiOp6C
sZ9Qv/dxssx7PhyrbG+aoyTRMkrdF/ihbMYCNxbvac9ZP5ZG98cUR/i1Ys9QqIMf
Ph2cBdYVtnYw0RAOMwKnFTW/mnCoW+9tbqUDXAq8Y4z03MCXiNGR4QMHIkV07Mfn
9zLlgk+VvUnDWFRfsQiyOuJn1VsSgW/HPe1LSr7+DH70v5ZsHB37yRFk0/e3ichc
X0VYo0QbAnDC1zKSK/noB/hdJwF1qH514FPAYL2snb8dfaWm309k7QcLoM8HnVu+
rMn7h14j8xHsZcCOIoKj6f4pQqPEEXeeEiUNYaM3m4w0LY4B/NYkFwy1y9QbRAXk
RgpENI1F8pNo+RR15IefAjpZ86zm1HT1QXb12UUaHnZQEHpmXD223Caqv7gKqite
CcjiuQBpv0WA4HmRCAIT6AV/iZp1ymvS8ekdY/OfVNDey3lOScaLpl36F1No/kP5
uRwnuAHYsu2F4++JtZJOJXSVIewC7eGFOEtUfdwR6TXJfeQ6oENzRqhCwbeHKAAF
8VidGjh32Trhm26XVFiRrjv36t5BgnybKkUgAjexWRqSGBmR2NL2GyB4oiZOAVhy
YF8OYCDnhO9tsovwcSZr5n7z5fKg9ume3TNtAC+OuGY77yKDpWLPTgb8KkyZcLac
NvcQ8ZeWZ783knBqyyagmOhYqTn7D1TOfEw19S2g11H/p2TahPfCqETHyKdrHYVa
cOKguI+aXqYqXbOMgXaKf87Jb/DOkns2L0//iV6G8qVnipUlZ8GY0lpP0Y4jLTDL
m6eMARk9Dh7WE1ToTDZF8+fVX00ELgWQCvM8ctXmfeyX1tnL6IXDq2CRbSx+p5B+
Mz6ICWOasWF0uN++7cIFrFh62Rygw/MxUT2qoJiSaL9vcGQ62inz6zYQwcWWyWld
AP3CAQGeOqR4JpZTZTLMBE8ChiCjlQz7jOPQxUeRa1DPIx/APmwbyvid/JMFfe+k
MnZieV5jYKOskrM5wLva5ks6BBxIBVKR8T9WAXD1G6kOyPpKg6RAVkXSBkYggINx
KEqDM7WRNU80kkjzJ3alNnFeVQ42/Sx+uooVWMAnABL4RMU+Wyw4eTt4a+BoXj/p
8NSpldCEazfpcyVNFQxegzsGYJJzQvgVjn2p7IHf8yQCFeLkjOl4aNFIXuNH07xJ
fT21YolnuHThlGmTrn7yPD0KAKt78VoS7bCpiIo4glgPJe2h1QkGVgoWUatTOzeA
7EsQrph4K5HPwZz4ArdSIQrrDJ1CyRVDUh3GkV7/fWiuFhbBmSqvR2hh4bDLYtwo
LfPOQV4iEZIrG/6IjmWY0re+aqTmhhmOkobd/l06vYXDYAsjooKQI4d6J4cdKoBA
HEg0ZwDxtab3IMHmPxv6QqUJUwe928vjVlDynweGT+a9+i3qYYB3ES5TGak1CvU4
SuRMmF/Xu7XExvT1oLnN8RImiUGX/gTvwwv80a26nXm7B0+pfmLWjIwf72iK9utz
NL6P1PVT+RDUngaj6xz5sxJTQmReysSZbdkpRG5ZMqASQCsFE7skXXee2rB4DFJa
+WHbBF4X0TBUvwdgFN/UfKmF33MvjDJaMj2TQK3/4yQhnzXpPp+CliGSUxbAYtHl
e9G8toXgbtAbXakKbMnkEM9ZXJaRS9ooQynVSB9dzx05cKD2DhkdrV3aYv1d0d4G
dYnBP9buvx3rEj45nYPyuECroq4K/rulBzQCablSk1UjYyOeBGqsKtS/mvSsdb6J
9FCelzPaHK02Kv7GOTXYRSbp45h5qDI2enN5yMAH2rj576qlADVP6d3kG/FnkmCC
rrK9R4EetTRUstiAbKkKRWo50jL2e35arpupcFhFuhozdxbEFMJvZpLo6Wl8TX/A
IrChD3d9PEkF0VaTsL7OQYod+9264G0b9B00OsQinzIbaKl2eHVzbENvAcdqYuX5
sp0SZi73mnimOWD09AWAj50IHozXECoZxgb6naW+VzuQcHA71R6Vhu9LsstTafn3
KYKjVO4Okw8zuijT+ss44Iha0ejWD7C2pqN+idXycAYvBifKB69WBYnMRDtSOv+g
QUtw8hUm4f13s6t55B96lHtbZZo2hnXFWt8fCo3oQdoYnALokYEwjWk2qs0B/tTJ
g9ye98spEZdUAXYQB+bqYtreLA//glDPylJ2XrJYh4hehtDacMQ//rk8o1AHIQTP
BjcuLFRfKWCQcI3wp/IBl5hvJTT9DzIWAyV3bHHQdYXmCyXmMPLz1gicYjGpMOC3
Ez4dBPEYQJkgF7XQTDeUV6RpwQBNBA3MbDqNCnpIOSBwxEFSNqAVVNeUnLvwywY6
5mUpR9SWF0pAhJr+H5DzAHmLWCkr20xevlq1zSk1bZs/bq1h9El+zYhrXNsa3Ux7
5AMb26/28QkHSSAayu5E1TkIOloE7UJXN4b69XRLwEeW+ypIWuvIRMBQETrrLkWD
O6M6cjjn+sZroTQNVNQluDMPM3vDrJrxf8oJD1pwlUU/786WRaNb8ccB/DJdOsvh
797prqg7lIXyWtPZPWLuAbewFX4rh771ynH5D/WQkCRZH6JxCfpKOunRH2YMfekq
RXGsqzRYmThz+95AGXY4ixR/rMUHYV7K+nc1ZEcsm3G7o8bz7c66kMDqW0PAOtmp
YXuVnOnk+UZk4LFvgKgY1Mi56VCaTDaiaiBQYn0r0aQmdoIb1kgyZ0y6Ctripbu3
9bZt9MCjV+aeAtpT1OKxsUy+LLbb5ZjFA8Ng914xl7lKWBG96w4vR8wEXdclmXbj
6iIHzbhR0Ss9vDt8QTFZH5EZgziPc5oJH0yEp90WOm46AlB+JZwD4oZPPJBlPr4J
HF4v5X0LdevXB2ljcqMJbxLyDEtrc+70QHsQ1bi8Q1+NcED3s9ITe1ANFMQRnJbe
JOnGByNJEAiqBVgXu7NToMI6z2RwN2/DxEFWJuSrSBpfE0TgcgtaAOOgmse+JNnT
hoytPWtmeIQE0L9033wWUdL448+r1anE7sTPamdDx22lA9uXiPEXZQERNXY6Iire
hJgBFLLFor/g3rGg+aPiGdhR9Vi+Muul2nBEWEkLN1eRwjAc77+0Jl1am1e3wNyE
4Dl4amNq907kXstDPno40L803GEnt3F1RGUbcfmDEV88G2+0LHqa64jbc7SdZ3hl
7Oc5y0K/M0RhkqC+Wo8hiWNVcP+L4u3JEBgdH3hpVZj+yi4CEV8yTiU+PQtmXMZ2
++lprFhVWGds7YKQSns7FBtnGbY8K3JQLB+Ex3itV2AbFSrhnXCbH1SY5VxqmBBR
Oh1vb65Qp72Ej7I0WQatJOOeb/3tcBiX75pazCe/9cxsk8IhKzBClU+PSqnRVUuQ
DhLttxvNyZ6j5yzux6YnXo3D87kQxbJ07ZY26iBEa6PRzq2pq13bD51CNzAoO101
iRbRsj2RZ2TvSvq9ISF1w9mssAptEDQAcl4WZ6Zoxcdxhixpq/8pefx/7BKMMadR
F+i0gbk6WRjgd0KO8wn+a24ryIlAcsi2vzEP3hOJ5EzSVrRiOvRU/3vSYfSXWCCU
dGeQoPltql5eG7aG7oS5VxvdFZDzDgOjJ8m+OTvM+gGGSppLNhGpmBFzmCsR+38Y
bSlXTD3KySGSq8gY6VaH5rRZ5DOc5SwkxMQuIlwCRB0m0rWal+UIFx9JhxKuMByC
D5LYLzt/Schj2wLQ/rFp6zEzUVAlIj4OiNE+ffalQisXSTpifUx/fS9ESramdsZC
HpNXqNA7G50MOdZJPBNt/jAd9sN82m1BG+XDOfWwedvoqYfj8vdJvIWxIApC1P1c
DtsVTW9n/rdGZopz05nuOe93BrJLEpigBjc/SumOeTVWo0i0cHjNo7w+1Tseum4U
8j+1LBg1XX5v+rc8upHpvMLTaDGmMZ0dkjZgwpp+RBBFcOdrmjh2Eo/b6tZB74KI
NwhovawRD+RKErGM0piS1vau0hsUR7FxvW9ZLyn9a+BX7tMwNOZPSls/JBHNs3OH
Td//m/jV/mL+GIXbBHkXLZS6KnbsHsbCGP4fYG27uNmvwm5+UGwoxTHbV80F3qCP
n3bJ1W9LA+uXX2+ekXEb2ILy6I8ogdlT4i9IqQxgWTp2JJd/EwGkt+jNUrupgysO
QaS/J8Gz3lOpGP2q1SKkPzYs58WWFyV9PcOontRBPBFtC52CKrI2xPXjjUDOlfHx
1r9oZpjIBTGYSfKGlsKyZBqDJ/rsT2St8YS2EbnklPmikufB3IGeMu+9D69kWNoO
X7sxrlXXGFKOF9ptC386uTcA8/mH+BPc6bf03BLHgdkLZynUydWr+ed1el6WFVeT
MWj7jeJ3NR8E5I7LXodSe76R7kYeVBtp7Zwb7XalYoRuyoW8aTRrQDlgGM1zwq/5
LWXlEE6TBtLr45SoTXyiaj8rNix745ZNJTl9JFZRtXycIm87kPsuUvmhy0uF2G+5
3UEx4+zxxCnH+75ymqJ38G9GsFXyTgqpg+YbPbf2GV8kxgjujP+dplogvJzhyp9o
MAHFuLl+Ip6bFJ1MGt3rum52vVTveHxyme9EBb0XliQmlz1VPhh1JPg7fUM0LrOu
vwhcYE06pazcppHBVc/TlbmNv5imEDc36tLPtSZvWnEzgFt+5wa8Hc9ujcokhj+7
VYIjlo2MFmfH7tQ5/o9qcrkasQviDJkTvZNjqI0MIalSusvmEGjQoZd6Ql2roJbu
RGxlcVqLamPjHQxY1r/ehIBpVfWLB+cmFAMsoRM7j4/Hf4RMYFFlLOPw3A7JhHPC
tf8CGMKQ/sGEBlVokubmspGNcNef22CW8lHB/aQxEIrFn/X02xP3bZeTJqz3e+88
BjcevXK8oF98Q6HOi9Vog0hDT+qbGFBfXd1ls96Ts1NlmEMKVb9MdEn/d25MnIK0
d+ixSL2M5uEoLCgWGEbPFBBsDHKdtIT59JGY/vZryhsVM5ocHYNIF82DaMRw/IiE
WL2EFz4fjD3DOmQkUOY8nA9R4SkEVbfVOh+GyUy5kWKYYsEhukB/HbJ97DFuRfUS
rlizyy0bSG9uxf0iwglTi0tnogGwNnxAH3ghvO0v20WZqRmhQHfx8NoRSutg4fPq
MX/PJZ9BTVHknYfwIuhpLKCKnm8WvQ4QG0+NJkkKEfYk3vXXVuUb/hVGsvZUI0r/
Xtu1PU/uQDbs2R7f0GrFns6Oi/+sWZ4AkWwDr44x8ZHY/PbSMdC6uo9pQU3GeID7
JHP6OIelz4mjngqrxWu7jFPQoyL/ByGyP6Q2CtJv8p00VisVagW6oAhw2jSGTWPy
mdz5E7njce2cRqwSTMdGgV8AljjIy7HqHlXdCVPQPKkIr3S1AVBelf07dqiHck4F
I2koO5SxjYd+A28uwBSp93I7UVRPJmvHnZxfO9bZ5MMAn6/tBefoDeWdGJHQBPfM
MR9uCvu1uSlgHQBcO6Gt9IC5LaNBq+1+Hp/T7CH+LpKO1PcN8sB7RFvcWyd2Dd1D
f4wH/SOy0WCbKEwXay9kSWgs9bVx9Gjf0yUfH8z4R6idm90c7y2RT5aZaV0kuPan
QEII6FPSiLZXY8ufhp2ax1v8B4HPv4DuJmiPFrmOXkFpLgI6Ye4OL9OMjlhP2/qq
WN6eIPGmUeUA7mhM/vTLwkz8WMOS2cqLBuAR26T7E3sGLp3CfAKFqSoenR5wQ+b8
MvMN2f1b9+TNxN4wGdRP/QyaWeK4H48VsZUIYW1crNBvPxFrtoWAjGYqgzvMv2eC
KymcPwu90cTUVeyLRQ6YFE5oKMc6p51hHvYTt6KpFE1Ugj198aiJQRBpTACQzy8G
LOxJDm7QFUTPVUsrnuZq+n+OZsahKSWN6MECdt5q5JAQN2j73GVcMNgGIyjQMPrY
SAcYU/5ubuq4AiY3MaF/zqriXQdlcFDfGY/E9M5WbUyRtnaPyhu9WTye/LSkrUyV
T7+k6jteivv+v6AxgYnVYAoDTfQANCe4/YVIRyABeRBxmL1HuOZmc2zFarY224zS
5jC7Cv/dYvhBY943hz0bSEWmAh96gF7H52cNNtx2rtnB0U1RfIQhyJXZHlvHMdIJ
9x4kjOIGyXf7nVOx5TJp+NCnWFPoQBtUYmt81/VzmuDD/uoCjhW7tiSqDESuftHC
simRAoVtBE55vyu2EHJbQOFXmEl33LBtkbLm7GB/ppalA/V5J/ELOmrRrJhQ2+iq
yA/SaDRHRtSE7DRuOE1h9RuT/uIBOl51AmWlzBrfVS09UQbUjhwOj7p1xUORaMN0
l5VD/NxyN/bHLPKit6aVHiyxvVeneztrDTgQmIFVnu/eSdhxshk9ETiBcMhE1ajb
i2BsHCitJDpdHE8sFxu0QUQxw7cSI0YsOWCj0VPBa7pXg/FyCrc09is3E/oIrii3
vODtYu0sxw2uVP6OSvI0F0ZbfTs5TfN/agZ+YVrss01goTQJnpAzxJQNVN0TLJS5
BA6keJd/4qCl4ZxcfL3bK46ijNzHOig1uW+nM+c/EIDfLQgJ35CKTdvdb7GTZqxA
9RCP6H/p7kDylVs73QrAXeBIcWNSXuAZllBA6MJ8QVrTz1fAyagDvdI2yfjA7M7v
/tM66lmchhAOS2Qh69z4evJFWv+8lMIJGn+b2te78rOyvI8JgM7sxFGeYv9t7hTy
09aerJ7tTraqucJJO1pr+mZgl4y53vQ8b20Ejfyv08Oq7fqXP9vl5nwSCo0VEzIh
XLyaa9m42rhuSAcpBQyugM8RT7LcDZT8Je2JLN+/4KTAqGvRouzeanQpvuyJFRUR
t5rTKh6yaM7XdPIxgfAAUmXgszVCFypssHARD6/+RIowffS3e1IEeL8vXzhNf2RK
LGaOrDWiFDzywmES8TVLm/vwPrFTb5tvw+gheLfkBZUfjtkcczt4Yjiln4A7eglS
Ow5WTzODZjP/hB3WByJDxCI2PLwYzKr1F52h+2Pkf8mwuvUjzSr/UY6cpJfFYUmM
yoMy1RZMkUyUNeheBhlYJKaXpceWWuYM3ZcpzJHUdAyJ0N6iOEgmW1EGM/2r5aav
0WebUxD8XT8rqwQBEcl8ePbGdy7SDd9HXIBjpeET0TbHN62dyuMrhy40FZJXVohX
piWCMMk8f63M38vYhI7RmZaz6U3nn3FclGvr/V8OiHsScF9UDZVEK71LR5/wJD6a
331fX9GDt5XHA09K19GuSHfV/+BnOoxNaH47wkXB6RQ10r5J8ppCSAY3UyTKCn29
9mCdqpmiZGxPaGWmSo4OuRKcwcso4l5RxecyUBoUVOj0hlhrOm/Teujv1hEe3B9U
7cGaB6ZOR5icYoyVVVsUMPS52aIgov6Tf0ToyT7b+wg+Hy3Xn0ISrlnXmbmTEq4u
/EAYkrwcX0hUC/4sX6it/b4eCIPypju7F2T6FSsTHhoUZ0yIpKOKyHw1hUeDsIuz
tCZ9M5gwVxQShUKsegDscoGbZtSg+FeZSF3doYXbhiA=
`protect END_PROTECTED
