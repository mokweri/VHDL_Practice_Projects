`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1GC6jrK94LKHZ52bBpewPyOcfcCUA0iEaZHtcT5zTQvt/HUp/0PfMfY5ki9Z7J2
wIgZbowY36GDWz2otQp7nU6gX9bW/ZmEO46WiPWZl134rXcEsDj47Pi1LZryehiQ
12kDOpZZaFq58DmgCfRM9lmDcjcnUTNhKxRWxGZeQg/gMWJiRni8ybba3J19hALv
T6Fr/HFF7X2zdIevx/55eCsOAqM3t0MkggDi7ljDZHPOjSl6axPtzsEYxuJt3e0c
Cpd9VcqHPkEtgeyWnb5hSNY/lFVIl8DA/RU2T1GWvzeZmMGWfqUBefjtiVpZlu0O
Z5NfK9fjUfRc0RzF9/IW7nKmexz7ykGMNF7dYdBbDiKP7Mpi4mubFdx3ZBsp/pkF
B+fHr5AbHXa3mNHdJTmDTqcLkXeIOmRKFa89bo//6FUe5m1E6YF0/rNFMevQslbN
aQ/Jiy5QjcVGvMPoUVFBaA==
`protect END_PROTECTED
