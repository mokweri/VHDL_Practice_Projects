`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xkMeCU+nYC2D6ZBchrjznKYSrxYaah1DiRFzveC4zsHm+IA7EFYRvtO5LGjgWOLo
xYFt9k02H7I6Loky/9Exv7Pq/CV1P6kfolByJiJAgdaHv7TzWlvR3Mpnu1PyqVH9
5cB053CHjOEec2QGtiLDdO1/vPfq+jkp2rVSTy5GKNBKPglNl6UjdptHHAdZGzXt
cyY4X4Hu+v/dHhrRoSdi745u20EVUjPAIepdta7qgcUr7dfrEU0xlyRdFCfv/ABx
6lckReQklJnwFVhVhbxrE63td1wCESvuwz96ag0GJNVq1N/HgtmSp8WegK7l+waL
uTd++wIuSou3G5eP3fOvHWzGBFfZVKasVXM/X0VydoeiG+TD4JUkhk078d1f70qo
xgv2tyWykgF8nZhP/Boym6kKcWznvoZH1XJylz4Eo8C1XFB/whpERMQOoh6nAVVv
dQdl5hlxtK+ocP2/GH0GRF7SpioAuBOGlwrgFhdM9wCOtR5oinEKV7exraHVuRUw
9TvJ6GFrb5yrkEBVGly31/hv1W8LPNbj+t7Z3qGfFWhxA6zBqCm1Zd+V7+XbzS1J
pe2QpSjC5j1fdYaYzdkC+8HFpKXS80QNZ3zEXYbrg/824/U+tb1aXXiCfAhOhG27
XWbIrPSzCKymu5gz20+FUWdZaRTKat0uri3HV7sK08lA1jTuZE3mu0PZPd0uYLSY
lbor5sIKAEMBT65LLhO++Ie/UEaJJPGsSuzJh7ALzjMPW9oY3H+THtpz5YPLoxSO
p3g6mLGTN00jxMQSqDDwtW17eWW74QGcDU5nvdHPjKnh02sabfxDoRqJJet87c5m
TZ94SyWJ32PlQPtToTAbG8wyuGntoqokbrMjuoTbE3H9BdRRJqrOR94RWIQwtcmY
i/C9+wo1zH6PlWL16J4y8l+DfTYOxxrcxehfL8Nrj7uc882x9ojA23zyFyVlYN23
6P6uHVG+PUpPHculw/UuQMj6ftIi0dyeDrTMRAqwCpRgZOijnaxB1Tp5vFE0QRc3
Cxab2M2waXQiVZqnPQb7e9sZ7XmtNdjIADQXromFp6WPwg6oUKccgJI50bj7Lkdq
nVaJLUwxzJ1OuDmzpSv2ILKe8r/xHDXUG2KFoA+Fj9MukX8RpPgnCt0eZ5utrJu5
U+COe6gHE/bm0Pbo4mQyo9vBBAxM8p2qQYASOz3ugPx6eE6RluTTIMXffh+PLNp0
vffyUa1bUmFkY1CBbdIclJBLWakhgnmXBdfFgmm8PQLV/H9SuUjdOu00D+tUqdnk
c/l+Uvs8jdUiy6UDJLVCtpY3vObcyAxDa7DlFZ7qeP2r4Z74WwvgQIlYiisDbj/s
i7l7xi2C3YQurEs168wHDqmzocla9wIOHyzGuPH4sbVU6HbkF5pZ6dNreODvmGF2
xdDUKxpwNTolZpW2cnoml58PS/btauIp7U0EoOWH2grquG6iojN/lsjOQY+ZEweD
ck32nRtbiJZo6fU7ywZ/l0IERh9FAJSqNa6EvDMv+42x17fGdczd71qkV3wBwGbl
AfQD8ghdBDEmFuYVSMPWmLcabPELG8GT/UvHROc2R12bPVC/uxAzKt5VrONd4qyE
vWJFEbOYGsKhx3PGj0EW77hPUeXSTRPBlJtJbdnVdgR/Lw1bkVZBarP9Ue0cs2KL
EUVfUMfdwZ11damAiWwcCxbcK455gJWsJbJkyxGDUXb7H2gLguiPtewWW4P6qCHY
oNKDzT1dphr8IeTPnxjkfKoBJdlD1r9S8YgFTiXLGxWmBY5vNHhUgCGnSUlTcFm9
LLPDFN4LqA9S44KIch5F1A5vFwDP2WCJ+scfhX4xWWJ8EdydKyPDZNAYYDtDO4h1
K7QaRvkqh0jVuk35s+XJMs+pTAQYh2qUPZUXg72e/fLZBFpx/IGpQBfQXFkGnkdu
U3UjVGGSYDrKW/wNDsA3mD4rIQXc9jvfpMrKF5t3lxVLFBF0O7zBy5tz/9wVsl6M
utEj2iVLqVPgDMM9UMK37lauwH0YVrMZ1GDTfB3eg2TL1DwT2wqnfQ9CbWoRUub/
wsLF2l0rnbMslp1e8EpEB57jQ1Qgr8RKsdLKkhrhOxjUg7jQhLHIslLJ/rcxV0nj
hDmThYbYXf56cPlj/zRNtBl+N/cr3mEfGYM8tmmCJBhPnx/UHGf824cAI0StlLXs
E+GhdFBYfnmKzvDIdWwxnD41ubD2RQBdYDQ32rHSiDsXTGEM88NuA9koynlJztPF
x2xXZSEQU7K2tiKsQqv/BY8Vgk0de5xFa4Ljhu8ym7uFlX1KsOb+vSAuHNKhQiTS
LADcpLaqxgTqywOMAp+FRZvANZDxe6oQo0PJZ5VDukQJ7fVuAGOXcf7/zjM3PhwF
t/qfU6PSUt3EyXouu+d4tUSJkgB9CMEvpqEPiKr7BnnpSdWn2kLJB/1TG2gEZOP7
rXcjgj6EfEeqWvlBPd7izIKo1rNUV8QGGjX5kefEStI8Ap8TOu0Vh3i0aecfmdtv
SAzkIeW4V3QkXRJagihLqcv0o6nJ30P9nItsajmjol63mGj8cJxc0QGODIoH950A
TjOpXvwctZp2jFS04GMfyzVgL1Xmm0QU0DdOgNVRPhGwkIC90yzYdVkyvyjTJe2k
3stzYKOGC6+NIDLZbZkOjOWnU7Ofadljf6ijQb8AmK8oeItSEyKOCQWt/Sb4Lnm+
z2WSCLboqkYD56BQNT/LRQru6CvJ3alA5PfMFHsQPxqTcvouFIR6HATtkjTB68xv
p/YYCK78MVtVXTvzKIM2t2j6cVLPXoHwwgwo4zHsHdt8TVwirsvXpJxOyp9D5imP
QP/W056QYoTcPR1SelXDwgSNR57zeZbpnahDfLhBKnUJkEKtRV3fPGJdsO4tQhH9
32SO31vDnnxhIY2G67FGgw9+lk/qZrwsRW9GhnXCBU3MUDNakKMkoWSSfkXw3TgK
K1BWQ3FEreMLtgMFjypYAeTbelZNG9/vmdyhbScccRWaMobWb1pVssaNF7SpGaK1
Psc8zCb4YTwIKw4qt6LSkVolQDLL+vaPXQK3HQ93VUcBFVMynRriTBTNl7DebJS8
Ryq6Qh7svU406UjjpTWWxUcqOCNSIE/MLV2m6IsG2FRB5rqFyrSvAZDVPOp2Qigd
m+vfgMZeM2NwPXYhPAByvfD8PyglcD+MZ4vzBaKx77vooSiiH7822E/d3F4uRgbe
tmtP3r+RZFR31nbd7zNf5fW3asArJTWPIl5HfXgfuQnxMZOIIbfNezfR5dlkcq/C
Q6hfCj38TePkU1dzJcWQ3bPMe0/hBDq9BZaBNAGPVX26sFlqrOlyrTSHcOLjs3G5
gCd1DGDnATe2pcoGbMWR3rbKHjv1E0/GDkf3IDJv5PDjzIUiznsV8yPhdAQyAqHc
CSXfQ6WP68b59hOLTtYSdNxwfnilZToONi/+/Z9/ST7C4qT0MZj6gldAsCHYJMRj
1KyPtagctwQP6Qfc64jRaol4q4iseaqdJqnhN1f6gtByKKL+GCrijl2bmgXJs1mm
ajPIbqFxxMYJ91zacBOrRsK3i2z8B43V7GU+s5+5bJul1vWJUFXxqUUzJN/4F9tF
Sjzn+Tgyds9mQUf6DVJloGdmr+qpf19RTk7dAjtwmWRRbY9BCvvpew+PsCjAxrCK
TaOLpGFcVcBugKxe0pTugiaH2P4JEwyt/8bkatin2XjAxWpfz89gboXOl8MFKpCf
Vi4vSQJhW+ULqExHmX1vIkcMRChEYEimrGg2UYVXEZzKnwfS2LeFNt5EDXcFSyje
l18899Dex+R2UVbX7HHlwXw+6HyYCj5nMaNM7CneuyAw+9J9JlP0rK5nuG4GjPq4
zsib6AWBSX2aXfSWY04ktlUi/6Nc8icqaPBLWeUZCVKMZvy9YKV/hT/mRjQjJ/DP
HgoIxT5APH4RGHMvDQPMeWkbAfDrKNztUEYpHe24HMUWO4M0datVr0WiM/tiAQua
r2JFQSuL7Vb5m12EA7eiIBxSqROFY9B+Cl04UzkgZDw9QiCW3F6e5JjeytBM/O26
D9TeBeN9oULPq428ujvqaQhqySp2DlGGEYaBkn1/9Z86K1I/JKftdErV3Sxn3HB2
XSm+N7TZt5RKPyw1C3SP0SZQ1ovk5u3/wMyGDpLwnHa2tKxh2m9Kgkr0IqGKek6w
`protect END_PROTECTED
