`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lU+j4DeJnlfCEfk/azAENYoOgN/O8DzjWxJfwJX7mOO/j4MBe1fAE3I6L3+So1SZ
wVEJaAxUEct7xRfNDlidV6IXEDvDN2gxAmV+rsyEOpCFsuDTQCaThtn+rflUazWe
ty1zJKuMDIA/EqfO6tG4r1EfoAmmMZEXJumMU8KZWHIA2jt1Se//rs5+3mdWtuLB
b+1lML6VQGlOhDeNj184ONMXfxGqMClGIdVrjzsqoOAz9f8DbIrAe/DGgj++lM1f
Mgrs1d8+LZxsFIKRFGOUksjal62fsamEAWzWRgTfk+GjnTirJylMmtnB7nyQP5Ch
J1AchmH+NRSdslsXht7Jf5n7Tvp2kJU96Judb+50xAUrrOEBoUXqdJb0/2ws59XK
`protect END_PROTECTED
