`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LXaQ0PqJoIL7LchYN3/VLSbgNNE4Ph8oHJIR34EYtfG6OBItt1TddphZHw6UKsg
aDFzzwIH8gEBAObxooVpd3muhguvVi37P/gpU+5/e4yBvrY2Z6FnRwVqz5C/QVGZ
WHpgOZ+6t1KHEFIdmwFelSR5yOWRlHueM3XjFBA7ONZW64eHnpQp6AwJRU1c2/dN
UqKuM+xSRD3hjp3ZnpXIjPzrFga6xfzMjqopC7bBdjeNjN+5m4yN65l5fbBqVNPM
/FOE67GWAw6kcRzgQc8DiPZoiwzW44fw1hTGU3giKv+YiN+sP4crcQEVpDSXyk3T
s9obQl7m63GZ7hTMSFJ6DhMoV2xPwmQLxBev0MsLbnKldOQ0aJzB7isrhxU+kFCe
BP5gEfR6RpG9qS5oBrWlx5KVqsRYp//c65LPKh8uV9/ihvC/YpxYZWv9PZJyMvgn
YXK4sC5WkkP8gK3v3gTN8VNJ8MFJCoyBWZKbYEw8uqae6sdfuXnz8KptBxR3bJMS
Y9UFJYktx+IVsSXWW7j2TpmBDvDCKQCDo7vGDCeALjkE7fehwvwYbfqTUy2Od59D
TZdnqQS7+qSZs0p6u268pdTY3hxbPoXwyDXbDCrYw28Cm0VgV5tpRKgvIGmvCb6D
gzUe8SET+1grcoMvw/kGyJZGkRtxF2H7uW+SpHqZP+s5otz6Vp8UwJo/+iTicPqx
uDPxNn5e7qVxErOkuL/IAkSq63+dd4S8S6EZWiOs7RfqL+rCyNj2hKhwLq3jEEcC
poyzmYXoTT9QbJukNG8Ztnd/t6X0yP3vTmiQn8hhACnsyEwkclymz4TZmPa+/BAF
45COhGXCUsaUwDZpr6MAV9JFgFt2ZLwDrypKuJtHKIOEpKC183YUN26Fd5tXZ30S
ixa4TYQhuv2bfaRu29wS72rU/uB9eox8RvufW4A2f4+cAUIovkDmBtSuW/fdSbOr
vFl/Crl+uwQgRlavl2sebrxL3xGHkmtV9VmXmLzH5TGz4wpR2l/5O/Z/XnRs1tsA
JkeQgQDmIieGOFMvrbxz5CLxErZvtUPKQTt5lUybbc/0ZZqJCfXJkCagtFYIAAok
rEHHDBWcUsJrE97/DujuAFn5oG9D9vSAyV4Zty2UGB3oK4Q5kpU8cYMrrrBIdvqQ
TEoAJ3lT14ZIy1QtgBLx+fR7tG8bPKDhTEV1iCkKG8BNIF5Sr41ZA+0F2SCnG3CW
PONpt/h+IxZ7gK4D3ROTP8dukF79xR1UT/mUxaEKodoNhkAXo7u4Hiy6LJiZFJRh
wL7lr/ynVVcqAfG5JKr6IjUzvjligmG0+J+UD31A8kTI1E4HpqOmVgKvPjtGDMVk
kowz/ut4AoTHi6/gzTdvlIcu+wS63wOenDKzwE+mHmbfWA3yuDFEsvbDnAOp2Jng
4Zfr0qVNqAiKqF9gzb0/Xhf08MWgHLIpgioNR4dT/5yf3eNA7uM9VnRKTftSLT0j
e/j7KvRSdPdv+JTz0u6hhnzTeQ5/MW75o8MOMhUJK3o8qvGq0ljjG1xF1KBqL8iz
i9FfB92Doq5+52bvnXmbv8xa3FRGxShgbGVElf4+La5SNMyQfxEO104za7sIkbVY
5DFeqehT/TncuIqBejIobKvXe+VucOFEI0I0mPgKYbiJlh4cB5cVXy3POcnngZUi
PDOjEeKZTYqOftFpKMn4CKMZTjpeQDZRSVUSMrGuExNw/pCyHQU5xfn2HkZC3eb5
ZszwAC1KhTciLBXLqQUvdkRP2ySgYZZsAwXX1CexbZAn3kwOv1D3uzGFdPsomr+r
2tfr3ZEnoPExOUiTo5dwtMEqwUiVZYAuGLp4Er1853R+4JsVaWCc88CAN57VET2j
7uxWyPrfNl6ZdeNoTByPKiRx4nBbQTHGR3nmA55Nyj1vMX9AQZzIZU704XEhKj95
mSGRCG0++7PdK211T1WUWFR6rsQIRzilgsnDnfGvDPej/sgSmdqhfOv/RYMWaLbl
nZSPKou7A8PD/xz3WCZCC+kZ/UvZ4I4IBbKlb2wBpgm2kUU89wsYePO2wUqm4Ofs
`protect END_PROTECTED
