`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7VhiHWg6lUGv9Q1ZWDmjdk3kva2FjoBINBJ1lQsCIOm48pq+vvzJ4GsfdU0JXlYN
tQ5gOm4NMIIJiVKmzoId9PUqh6UOOHQriGC6Ohkrh/TMDoI6TWrWT7iyx1iKWtqG
1dCRP8O8WzB3AsxYcV44rmKulv1s/A+SDpS55YcpyvkfuKm/i6+GtEwvRrt5mIzr
5oJiQMMjYFXq2Q68BSfU0gK4hkPMBwnDPnS4BqjnMbd6FsD+kkvCbqXbHEsoE1+v
KOXfR+3cN1lAqFWMnaPeijhHP9mOJ/E1t+4N5qSFFCmNARqVTFTDPiH+04E0kjCk
je4LIxe8soGK8Atovd8OiME32Tt/m5XWrEgiSidKKhjDu24F28oMDYDB/Jf/NWFX
ZJqMUJzCimlhqe/QPCuvMVTgc0DUNSl9+PzEdtWMYJTrgOutCRCG/mwRbvWcYGmA
S8Ba1jjWC2WZqRnQWPg8cpJxH8EtWSlBjoMIzG0avG6a3ho54jCQs6FBmT0vNSqO
0lzN9N9QLgRHawBsTCsaGVn8VNM5UpWpn/glqzN2KTj3awkB3smo2KZy0DJenJB1
ks7j/KYlZh1LIoLwxMJsqpg9Akmk/ZiQ8rvRzrB3I5GKGGEc/801Y1fidQNRYmnF
OZjUHwOCd2uFkO7s8Tk9wz8SbxbAGjvWNSprEgEnhdPw9nOy8EcQSAlf9Wx0zuyx
jIvJqOdYlBSUXLXHWTOTbspntDkyyNdIoU4XyXZToUgrSZeVtrBQRr1D6zdIUgry
9ePoR0TbLX/WEt1oh2Nd2eRcRbfFKC3zfpqs6x60PHBkWdai9m1iuHe2+FM/9Wbn
KyceWDkuBKfByr5bcC/i3SLJQKz4tAAQGGeC4YYMtaJz0pj++g6LYkrTb7dA4vUy
V2/CmZNmDX5q6a1VSBOcXgaPE6omRRE+91RK3QiNeIrTlsmgoq4G3CxadrBQdOmL
zSNi/VWbNGKXgww3Q/S1QRus5eFuTfh5FaNCmxgk7R1uJEliEX1xKJ4eIa1mToXJ
wbiODx40w5FbuMqu6PEalxxG+sBRFmTVfa+cYLmW2OXTxUk1lktMK8teCPILGYUB
UHR9q0au63xhul2Pdr4drzXYBXMWv6scYMCKs/2yhJrDA7fcg+avfwLirRKiPgSs
hO7OfN0i+DIDgtC9RW81QGTSw07ssiWlzbvFKr5YZ6cXMa7Ui41DbySUlh728qPL
qfYoo+dGtXt343M6+ddYxEuCCK1wlqPMyRKqKFTTVgMid4gZCrAlzWVaH2E3pet0
zXBZWrSxU6hjhyAWPXBxYmBp2JZUgSguL48uJyJixNyR1KIKLeRveXJk3F+IxSy8
2x/rHEyBxGKsme+Xp+/s2qjQZLKOO45BrMDyf2slbIQLglOEjIZ8u4Id+CIWDiVX
Ptx6fvZGzzPIPiYsrA8Fw1dUAw81iQXHxHtb8F0qw9vnxH0J8jhExUUN9YEtgL0Q
Hhi13hEz/G1IIkrIHxXJjIJdByF8z33EdUVXLx1L+Fo0cEhMihcvqiHNHZD1PGZ0
`protect END_PROTECTED
