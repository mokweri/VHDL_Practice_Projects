`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5JJZNYHyMMfivTXv7uVgbU8S3WphL+7r73O+usRxmnFJescEXve0qT9UvuRNIRa
8abeGo17h6VKM+C9bAVhADDlytxmCjh+uv9uUi4Z11iLBcGe9yGg6HrPlBPwuCuz
Oy04V+eCrrr8YXFQH/jJRXsaMHnGSNMBpddboHbWVhZBJIFyhY5IvIwUW9FmQ48a
4MJ9BOWhMCrLsVcdTW8OBLGcCO4MeTSI5IfUbRcDyvueBkwSvrnntXR2Rf8WKGMA
lsEOCjaVhyMvXGl9mlz37E5NmHZCXmaCsSLUJI/SRIpmih5p06FMHz2brNLfynU9
VvZGZP2cYLLggm+iIvGL69QS5kjG/uQ2StV7zB7gPFpjtDJPiVntJeq0IlVrTqYd
Lv8omobmAeT+Vxcpwkwii2/16WrZssEY4MmVPv3+CryVVj21BtS53qnDJFGl+nJv
KruXDqEQgwayUUF4d+oyj0voA5+gtDNAusRO/jwNKR9uvdTXSGw4LPBjXq/m6fm3
IRFDqkdN7I0fbgsVwad6HigeU6zxbzuChVbYgq7oG7pwSfmwcDxc/J9BKgyF+ZEA
aoHtzDhOElyAsg5aFz42qDhs+qBXhY8vra4GZmAeHfzs/US0WQTwsxy0zMbbWQnX
gzYYEXg8BYAFGpD1PaMttTHE5majSvCFBjwDL2Hdxw7dS/neRWaRGTDmOMNdhrT1
WrF9mML/aXT3EFJMAvCZa9aWQa0qn9domj439IcC5RrowtRQ0Ilw9a/pU+24ivrz
haumw0d1t/oU87XbUl985NzfhiwoIMzS8uuglH2g3A8cKYPovXHVEtubD06Uap3O
qlBOZT1u1YTkLjPNfHs3O4JZ887qKdd2b8VWWZqQEsD9bZuMzbOFiy+NH5KV1wrO
Fq0PzulBy8L4aTatxYAOze5UGCD0s8/Ou2mleJ2aGp88YIjFBheqpG825nUhyrV1
8ox7clGI+oB7kY7m8EWcnEbBxgAAMhoegmL+3YSiIyeImNxllKfiQ7w4ltsIIFl4
R6Np2c4FuehFCmSS9yxHVdE/dRwz4aoFNKMLO8jdY8k3GAlizWb+vRKycNFmI7Dm
rI1Q3qZI0NbYLEZRFO4U2kHjyGGjCutBJKk5+unllIplERZOo0osdQcH+m3BUi+W
6Gd0KiDDuBsFHDT2mlfRkpCtl2Vr336snflSAtl7z2L0LPGgLBLiIs8QtqyOiYJL
N6GDIXhfslq5EXRS0ctIVsDzt6CwwMe+FppQAs3IPHDSlFyj+rhNoFcQtH5aaRjJ
Lb6iA6fZ9nzNCEuJgzO5Gvo3QvXvZeNXhwDSKyWzg/XMDDIjA+m8TIER8v6rWPVp
Fpg9tjwYPJ6Fo/9X/jmK/IiAwm44lRfsDfwswpfiDtIC8OhNE16fVcVmXsRLLYC1
XWDLDAyzdCVTQrAUgKlIUS5nkcCvDaX+bwQfbVeWB2Z6RWP1oNlPwZCOhshykY/M
3V6EJBWuTzD5e2w9kfnnHMuy/bPzq+vv7EK7mvZZpqq5TuP+R1ilUNKXjgK71SRp
W7viNb64ZuN65/+EoCqzsATYK9k2i14lJhAybZSYxCZ/LiqGNcV7xuBreA9KRaU6
5n2VRHkzGaj08xYF9NvecwnGSYDy/I+KN9BykLx5es4s+UWLx+up7CgDdyo2bWH8
8jYopMgDSJSCQMF5qMaI+KxAkRa54YxZ07MB5g2q6S2aobBznnKo2yWgtxBdrFh2
+5uVpPdZOjolPQjX9rt0p6YJcnV6jDuqEsbRRn5OVpjDq9Wni5K5gAjwXyEvoc+s
hbQAvU7TRJMQzqEKSpFkbjXU9nOkpZWt15PNmJ5HFy6AEVw1nd6KhPN6WhTDJAH7
gYSgGU80/FesXMVh9qHqUf3jHcNIS5tnTBMZjzwmnQhFW8XuMUy3MEU/NicTUuyi
Wx97/TAUrcI0UDmgywsWw+y+YiJ4EG39J62+1z2sHgbDixdcStJ/5BJ66HmXV44r
F6N41gq7WUTZuazym1/MzpRq/LzDP45YtjylhRbXbCIjjOJLgpW4MVBm2jk7WLqa
K5Z4fJj9BC+bsEU5JHLWnVDO8+2XpCVP6/Z6qqGBdPBqRl56W5AQOlrLntuVDtMk
tpiuQCyBh5CG6S3Awbl6FO3BLrAmwPk5Cax4LC1sNxExAY/uiQIvMg1N7s5Xhuf6
OYKAmsn5AyRng2ixL4qL4kUjNxcUQBX0ouUcsjp9V6De95X4prV+eJEEcvHuzSXX
9HF5noy/EPx3ODg0D+mOCJDSkyUyVJZeVEhu8wJlEpZWlvcb3sSfeJjIAWk/32nb
i2b89jrq0itHg+NJIXTx9mCRZD9CZyvxEOjj1bEc8uxwzuqxUHj6E7ne+FimPOu+
EYatkcA4wbSUbtjg4e/q8tXxnwZztuSn7Fs6nc7v2SnmGD4mBfy25I0XXz+B8A3J
fQfvk+Z1PFSgTJmFvWdTdTX1Obgm33eMYd/hESMPli18z4J3QFqCdnWMcIMHp+v3
NbEW2bXGm2n9F99yqUl72R+EZ8ZO6Zr8kYz+NRoTeeYZdf/tBhli6llYXU/4+7Di
7I9OfUDLLtwG8OfLQ9m6ReoleAkklRUu/q4lgB+p6WSO11RrCyyxoZm8p4W3vdT2
rcV79kTCF1KOP3xNDBdLKPqgRoV918A5305YxtcmD24jF2Ihh636KvtrJ2smd1j0
cSziUedQmXoFTDX6EQZqjoniKfby1Owg6u0AKKnbj+sAn9dF/OOGGts74Pbpp302
IA28/JUfiCRMca0izT1vxz9LKmwVrzZTalelLfl2aDX+urK1FDCAeOf6v7v839eU
spF1OJ3ztbTUcKo03exJzC99stfw3Udru03h/M3aJz3a0KQANKLQqunG90bc81+J
CP6AuHrHrq2vO5I0VlHsy98hKEYvRS07NT55upCeUzTN9sCAEnXtrChJtPdUt+aj
kogmM4Yj7D05WQJBAw1gTwA227+VSYyp1aYe68ZK3rMRrmFz2WGi98WL9MFO3KlC
+4DfvYIxJ9PXnjZjmMv518lV6KL0W/QOacefLIZoBFHpCpi+8iVJsdoXiAhtER59
46BuXqqy+6Un8mIJAdmgTnvz1yi2JZx7egpDgO93729QwlcLp6ZOgDS01SzQskmO
dcOYRMys6z/3YGMmQs7rZ2c+k8bU1IrE7o43FXLo5eu0yPOOyTeQDriNBaDXapzV
9f9GFIqw9VcOj4x/m/V/AquugV6xrPKwdx+fxd1H9w2htaTizQ+JFD8Mc8F7vXq8
ScrCYX7CGMSlwuzQaidBia9OobyVB5y5PHffCLJbaX76mWGZ2Oia/Ja8cXXR+kGb
TZ41Cb4iD+QvZcYMZ8KBiq6kTwEmbzvdbx/bOyWRccqGuA6XJDKWqo295SGp2Y6s
pw8bD+dhfkr4MDwiEMt7Tbd6NSPWZg+sga0okNDcHUW6LhP8J0cizqajyZQ3Xw5h
GzjGqwl9WgnlNcJY9iCzNWA+4ezg2MgrQxrOV18vC8wAd6NP6GBRjWTttlvpQzo9
RCKTT/bla0khhL9N0eiLSc8791lxZLM05DDnBxRDZ4Ev6oAfQzQnPE7pDDE9JdgG
iazvXXrXHRzy7ajFTS0/BF/1iUmwNAJiSLSV+u4XgypZmAWIZaWbRi/+DNtkJ3cg
SgEro7SHNb0uD1lQaqsqKnibHO7885fp4oOEz5uPZPKECPARgXSZSXxuNSt8qCkp
1YHGSeNpT92+hGcOqHhMLNpMS6gfcTIwzQgadxhBiPr3l4ghOIoxAHc3F8ynKQbU
wMMTq+gHzKLUJvaYMFyftatuaMc6Qnt3sZDxfWP5i0ksOAcOZUUzQc1mGQ/2KJqG
Hi9xYNtqeCS+oawiI1VMuyVNwQdNGTzatxpUAuWI3dTvZt5x7JOd3VjwRXHAtn6y
4TrjD0dpnuykkrkSzHEnvoseHeWBgxBT3pWCbBiC7PFCMU/dNQLAQij+I6anIdOT
RyZJa47lmitKLzTqOLt3dQm148hdIJFdkQNXYqVOC3GWaWESEBeZDc+0JJTdXfCy
MinBXbV30Kqv1oM2HjYoHyE+FPNu2HGCtzwBukQcCJQMzn33MjX+fBOSddhop4YO
f6QkIgepbYNBBBvNH/FTxGhzYyNNDzVnBlx6jJjwxpep4SvvW1FvsJsu+MSQhdSq
FJvSWv3R/BiaXsa2FemjtUiLZCLIMsYedIZx3Xj279kxofsLtZxWOBv2ExncFNcI
NYvUCRRnTRRywjCaZYiw/KvYUItBknrpQRvehdX9PsZJllgCSK7n3c39FsTg/hal
ubWm3OpEUlLAAEbimajw/Eg8Hzvwfblx1PiJsHKxwdtF+SVjnwIxa7HA/Y9UVIMh
hFAtTxvZzWtBrPkF8mxUBjxWhWh0vS0wVBE7Y6O4WZzB1Wcp4FWswxhCL8hrX6d8
IkZQhYQsc1r63uQDXEgHJc9PtagABULtTukK0YRCJqydMwnyV5mdJjyi3vXiBkzz
n7In1VxZXmgjxOX3iNi8HvZGLlLxWV99xcPEZT3fcPuRHhYsLBLU3TmpYSyESmLJ
9SnVL59YImUTp4UFKJxys6xtB/NFQe5mWKfcyOlKpBFQscAX1Zl+Qx720/uDBmth
MbfxB+BDxmfq3bLOymqNWHjA1G/d6UC2cQIPhxk6e7gnIuY/+wO4xGat/ON2pld9
PUaw4snuCOHlOI6pVn5VxWc9I5t4c5Uv629oUbQ2MMYkQh4tkXVfbGQjmfKvBH8L
2l4qEdkgk8yltv5FHjd3HlhhOkab02deLYCpMb8Zti+kSjoc1bgdQgHnZIokj3gx
NPPG30q42IyfUzUgRYjUs7hEHOHyf20JT53MYF7QwYnUjChVfN00KbpL7NbnNc+x
hl75jEy3iNmjHWtxm0VGmiq58/oJFU0eA3H7yt0vUH9Zr9WtBhcovG0WrM2MCIFl
+SZEdvqH6COFSQpN2ZA7CP/5bDkQaLcMxE/0K/6vCAI/oqJdIfE11+hpO4+f59Eo
semSjwsHgoDUqYUXI79qs3/gL8BYxpY1AF5E36pwa77xII7UHk3IVlCu3qyLUmjx
rsDfBOksYYTqEuX5+cH7Ttxl6781DgTZw89bHJJtLEnfMgu3Gl1/bBK11eJEta3S
wKqNcdvGNWD2EYn882yCkLxW1N8CSWOHzFiTGbsog5L0dz4p7z/97iZD2ZkPbSTz
yCHOkRh/aZG0RkSNmLdJ/IxTJnMqIuvCunDqy7jLLWanceXlwbK7Ic0M9DpXgMlW
wl2vX1BROrhR65jbmTGOuZxdMtG2mudXmJ+f6xdWSnKiH5+qKCXTkwTkPynw/tx5
M3Os7XhMLD1F3olW//Fa3lWSwxYKCo7uOACC00yhKgtLdPUdyTjVh0DwYFiK7vkk
b38Wug184Yufxhc3cCzumBTkI717WnF2hgmn7MGVhJbgKRi3oGKxs+bZi9BxMGg1
TJCGdw+MGK4ALZZVpvgooO+aCgQjaO5LocKAJ178w0N40sMi6M/6J78cWX0XvpAo
L8gCsnk4pRSiCbJAhYnmFwolIi1sB3FRFmzY5nAFEMs2sA5W/1KbeQrF5dvoBy0D
Tnp7rkE/Pg5jBoEiv47xdKFdNdGgnOUu3wHBSH8t+cgn2NEYAqKrvTEtozzTQq6r
QpMvnfU+2YwEYwEpORnYCyiUgbt6czEZSY3xNE+ILDhe2pxO1FqTbjiFRKQR47GF
N/OpR08BckkOqh39J7UzsYU5DGO33lkjOzrHhYtxhZOfRUjAaPgT7v/HuCLjxDCK
JgPn/uWYuKmPpNvMl5pULSk8GBbKjwFEPuNr3GR25RcfbgyAnfhP9qkZHqa4WD1s
z8t/crxC1HLOTAPNUEMIiORU97pJoFLaQ+WtPf6Fd9SQ231n5kEJOa8xsMi/UaRg
XmxNKgJhTmUM7isL+mzIda+R+uDdQp2yImup/1wvlbfzt2GrMR1P67FXh2wKksuQ
1CcaJlaXHjRM3Jj5dGEB0R7Gv7k7J3XGwsvKq+aPdOxwjNMCZEsjM3Q9WgzNIwE2
e0l9Yomqk+8BaG6cTAu2SeNuOTyfI/vWGSDxXAqeahQ821vJSMq9EEnrzL/UuHxb
KfSUi31YirqTWfXkHFw1nNn4iR6JWuP0JUpLZEjVXeXvCIU1UJRXSqOH9kEoAyi1
1ggUrhP/IiQerJPpRnDAmvjhojVu9I+fMlO3cya1edVGjGn/JhKnmeHhizmOSVk2
V45T0rBbP0NKdRdgMihz7LTJ0SM94Di/+3wDKeB+ZioojwI2Qanq9TEU4H+gbUpe
APGddmF6FzVJx9T0zzcgmeOgNblUk3MLJc8fdqEMvezo3h6ZTIVupNz/xWKbt62u
VNG4wmHvmRkAj3GQUdEyk8KuqP6WgoGogAq7B7Y2kB0h5fPXhZUuYSSrJvP9fVga
16PlW4hWpnVr2N7nbZv09dI6TUSE5TEnTUPwe5K5mzX2r5mwEizd5yWD5tX2jb+X
FI4E1ScR2dXEglq0O6jXvEanKSu8wfBvKH2w/v2gtdJie6YZKA5ldVxKxzCZfA9z
jF9l1i2flkWMl06PwLlBQj/st7a1Rd+EUZuxTeAxxNZ8T5GJd+qZregnERmCA3IS
jn0a7tx4jIFK5aTGTtofb+MhLnSLkiv8i0u3qPkxOgIphoi9a/mhXSFtr/VDYyHu
TWuw6w1AH5rJke/TzJ8EEsXP/6OPhD3sn8QiRljy/Qhfw3XfptvBt5+sV2KkqxfD
Jddh37hPKLy4jHDjD9AMYOr6LbBoC5C4e7CIlqNS+vDWD9hlWvULKwBprj6za/iw
y7yjI7hNaJR2BBy60KpEG4UhRagFdE9W7e2fwC0dR3zvLTT+WcZBPqW0YIlPm60w
zKfNgc1GfDeGbMGw4rKPVZpkiecW1wGvAE9K1gBB7+/dhw1fZIJy8qhCf2PJ2udL
cUmtrY+Jd1nEKjS3Wfb7LSHJHaZORrarcLB1r5Iqe7vzHsy9ZUJmZ1GUfpwBmeyl
tGJahf9u+/pxa7IUBnDPT3PwBAuw3JYR5AFBMd1vs8ycpwKndtP+R2j7gKi5GJYU
UA4I9BqLezU/cU6DPeLTYdzWM6Kvwc1hCtCRUyT8CBvXau5VnfgtH9sZ/u9a13Ro
wVQPGxJEs6w37U164qAAoaSzw7OCZr6WGNzK3LVrmJUL0iTUReBkW5KPlLT3bWWw
Y5Mb63zU0HONetpTLTzLgYftFi8uSwlO4s2sx0IzvkyipkP6js7Zhu213QeQsdYn
FLcejJdG/HR0fey6BeJqDmSxyN/i4kNcE+ra4tgThxNTTPjjLQE//81Ffofo5yC/
DONAPEM6bQeMUG62SnEjTZsJzMxojlhX8W4Ry6moKMaYMo/j6CV2uLixWrXE1GQD
wl4hGhTzY1ZvjdVVnSxEne4l5UY0LdIT7jn+IDcSA5vcmfG+Qeb/vENUGMEx5Aoh
4CIMbFvVWEK+zriJPmSYr2oAu3hdREVOvowSVhsxbKRKUbuRvRliZvaCLQPjtpgr
H9iuDDlIkdqlfgvRQl1zqWHicB/onrjMB6tUQUNlBfxDfAG6XEtTN5ZO29+EvhDR
SZGk1sJCY9BS/PLXOP14SCC5Rtj1ptvgLH8ewPFCrt9RUqfLK7JDHIPN1zhWLX6x
DpJd7Wi8E/l1HOrqm6g57e+moSTDc0HHKMYkLv0PTdUko1wj20ytCe+wqNqZrNDh
c5ikiM+eAnhZGHzbAuMze+ignWYm5vrrsgzuZDamh6Gs+uSH3Oq7tMBjGaQf4ETB
JwjCkjYBThoUD06MQ+jPXpPykEcpuiWoINJ9lbNNiBjm7mfHuT5s7l9Oxjy5SwvT
L3z9Bd4XJtQC3q+FPPpj8Nf02Q7ES6wUBNoXGv1DUiI/b1q0wD535mm9E/9ZVBUv
JvWVB1KQID+j/2oETvhRfAojNF9k+7ekDEW8OnORgM+h106PjP32aBQijEgLutCt
Jgt0BI2ppuDHLJoVkFdL5Cz7tolLYl6Ol30mG87lrwvySft8jVzlZtImeAbL+RN5
cfN0vewLhhqvZPR2xZnjO0/Q0WGgYdeUiMyZtlT9aopThMkHgC2jZdyQ1Dh1ip6G
sJ0rGrtkcKxUlNk7/D9iBDBoKlbvIghMrIy5vKyA7h3PqgBYN5uoLN5eTbLgFk9U
x9wfH8Rt8rNRFyYc9YVOPQY/T9ZgoDFaLQmBHilXGcIVSP2sno8RsGBAVaesB4PF
z6f972JBZlkDxLzl3gRpRBdh5LD5CKbYcYVJX5Yl4VCgwHZ9QSG7vsZ50PBpIZLw
ApPpZsP1gDFqSQvt61EUmqKpwE4wAiWwCl5bCE8xZKHpKcTsD4g1wFjfP7yq4E/G
PkQuKCdYr4/WikoPN4/4NxmAUELqudlLJlg0H8OmGaEvPlptJ3UvcS52KKtyNfC4
755/0ju6fNiNnRwW/7FLTnc4GAfCCpJdTkfPli9h1oGuaFU46q7PMVqAyxPPS/pr
xs7QaHY/eUPlbbAoc/v9PtNTGyfZxibjtTXvFptCNRDrxWxvHNjTo9oT/aOihy7E
Ar/NvK0CdnT60aJ/L6Bfgv/wEvjvkauSaCnG25q47tAe2Bt77JWHq6nic4JhZ7+d
mhjPCgaKFUPjmtKcuNP+Ot1pUFRtLqBgvQzOKkZbRf2ja4PfX/oNJJ/BU4tflsPJ
ms6IGhebYJBhZm6kZuMiTVZO/tfEI2fWV1RTz0X3r16rDQjOo5TlDbqCpUjtvaPi
4INw466qzg4oXqzXOJkUf12LYXJXeKKf/MEuET8P/P6S/JBvaWRPXGDVeJlSw3t6
cpOs7mHD0O+qa5di+/+0MVbC/S0GQY8GQKAQaLVyJpMDCSgPGQw3qcYedpxK1tFo
9exN6HW+yyi/Z0h4eZIfG5fiStWPqqCl2YOcwgNKyk8De+p/XM4io87MpJL/uYYp
OU6wm4khJtp9TnnRYS6EiwFDn7WfWyKJUAU2lbTzefOY8uErmPOtoADKZfX565d5
eIDToY6DH9Fc8KSmR4oa36s8HfvmusYswh6DIadewakK2uG0XLqLEFGHO2sKC6Kf
wmPJQFmx92SywqBFuu+ccJ8ZgY1/xwSoDFlayXc9GU77zGrnXMRk3t2ab5h7ifr7
y3/wY7rhcytdqePcBJ/a0hfy/r8f4zeJeBT/vfBKEXeHl2FVz9cZ95M8y72QBh1f
cFgywTo0gi01vqGjL8BZsIGeioA7pzdpUUJZ2Twi1PK2zlpeOvBEcb+HXG7LyyLQ
K1+/PeLsyUHxaJRbmwZvPDZn5bA7EElgBCRWE8XJE0AiZYpTxAj5jMh8SpN27BO5
OEMbJVUx4AA2r1vo+NJOkJvnT/m6Sx8eFxr5clfTmzrCpwNf2M9MJ0HGZ5MlDa6i
x1LrrnKU3/zvMqljnFBrngcAm1OWDgmCSanZuJSrapqRKP0Tr6mYKG3pagOBSe8B
sI4xAQAy0Fnao1kSMdYw62vgoQavsTUHfQyHYsMxZOTRE4nP8M9LdtQ0w/0ElgrU
XzJwIZnomnwZK9xR/alooTkal3uCbksmZT3tPWKQWmY4u/H6TKoTatjt9Mtu9/5U
93PTxVC7II1NbBJJLnczDmh+Qcodzu4lNBrHXW+tdB1I//30W0CwgGhFvzpsibDi
6ImdDgjg8ksw8EGexXNdVmfuJ0hSOX4HbebH4YRROOZwOTfx0/pUlS1M3w46B9hH
`protect END_PROTECTED
