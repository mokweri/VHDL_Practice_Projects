`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqz5whN3f16ipBNCu2fSjd1T5/rat3IeJHqxAjaz6rF/VlAZ41GJHQEhc+U9ekSA
ropf8z6P6RCO7wJYV6tQmRqiR6YrZg3gH8r5yP+BMADoAYqHl0hlRWB/Hw35HpDp
MdMo0EC66dtocrBgakZAaZTLQgh8zyX3mEy2PKGndXeKo01yasT7A6Pnxz9qlJA6
yVAON6ELg3N6mWHpdcsEz7vDwAgmgiGRw2w73J4qa+xL2ZZ6CQ6wZgQ+B4KB1ZYW
NuFY6LXy+DwzjNOOtaN587yZJVXZRKr9ud5SLRHpSQzirGtlg02RCd/suYHtq+ii
/WHGxZdv1WfgbyyjjQCqCiwDR+l5gweKucNCre/90As7cZXgpo6uctesHeAzvb6n
eXiDA9kZCdfGp9hPIYD/6BnMHYHJb6Pby5vzUGBVTSHPRa4vUX30WKhbOaFcqRVx
T89ZoXPYzHQ6bkbfWIpxEVMTk55l/hm4E6vI04Bdr+2HTDAjXx6vHzS7WLGC8Wvp
/wxtj5tK73F+o3pp47eHnK1M3yu2UB9FCw9+ueg7o74fmYFG9ggy4L1MFeSW8w2H
474luFQ8lDJp4owk7bNScn2KYssv63UDd/0gQTND/s2f7CiZ4+saGwAy17nmHaMi
21f3I1D1WMVfudx9DFt1t1nz41HbqlFtIEAtjTVK6j0mRC1VGe9W+eqg46ogMnbr
+gnGEGg4e7qdP9o0SrzOb9JOCfZqoDbOnfeQ+5HybSBLjnLzMZb8vEXhNCyz2APo
vxhNwRdtxADQc+X7pFwYhLm6Yjuk09Zht88rw1EmtpGaPSYIX/iqC/uUMrHn3KmT
nkQ8R+S+XnApK4XrA+HwpCbKaBd+1B3GVoEcXiKgWrBRR48ZqU8beQkzjHcwVcSn
9V7daePswTTn748v58PzYW4xeXQ9nN1dun/B6JxyZUmTP5h9SApV17HqWNGh3vsa
hqRfWcEtJMTAkPBVWp6IoR/yNLniNxM2eYqLHEokKydnNLSJGO6lwAwZKqaqdWuu
Sh5dS2G17bMoHArEhe3h1NmDfrdmWIjNrhNpGNTZzxXpTTUDdNzHoTJ4f6UnJvpj
Ja2jdMKn1ywIB41KH449pKzhYRI3r/8zZnmht8eAbbTk/giTzSso6xYavd4EWXun
at/vadnZnqntSE/Qz1o2Ib7MN8cCoYsfU6BmcZ9uYiobfL91090zDvERESoAbAK6
OaEVqPK2cM3ghVwQFufYwZvehVvIuT9siyrq8f4CBNa1ezMsq+FKbIzCaNuxzVU4
3kXAsx2GTF79wKhGzVGm3ph8tnQ1IbQOAAuqvW6AQ4MVtkXvEA25kq88l5jCD8Sw
XYGDwmLFtdhdn9xYfH/BmvfSSKWIZMNgb/Mr7Pv8/nw2hge8dQ+Jayh1ivGc6btF
jWfIhBfwCLYkjxcw3zC4tor+Z1ljAwlf1aPs7kEoBnmovMOdz4gD6n8bpVkuU0d9
L5Hz0ZIWoPZrWah2pawXiY9ZxRElQplc8JpBrB+zK+/xiZWLgblG0qOcvgSUFue9
iEa2fPcA9TfP3yg98D93qT51FhBb0VasABxYI98LufrT8gQD9X2jyl3kwmK4az8r
aUCY+v3pz/wFVS934shfQwZ3X4oFAT7HZWMgk8cYfnqv4SfDvcdM3GqDYxgkQ8Os
HhPF0DMddirYh/+GmK+fySievQBbFSeh/3ThlV4WQ/+JXOL+AcmNSbUC7qkExzVe
mn4BcgYWUSOi0giSIKSpKHdJWjyCsiSt7QUff6cnuMiCHj2OwxZYMUNzvq4eRVgz
ILtjjT5+gcTUutkrU89gTGp6QEcyYqUhFwCCCSRH0K3SVwlVHzYqePE2klqqSHuZ
EQt880dw3N8R0iJBa/47LN1VwbANxD4eCM9RdWS5gHYXJgy7uEmINXZzJx6Xi7hq
/J+U7aCmGDWonJH5hT3jcrA2vSmie84R/sVnz2WlMGbzPmEYeGe/KL6JXXd96x+y
V1so7Jsjht6pxIYOiBRkpM9YseywyFCmk/FHcZ4pxxS43pI2js3Lc2sr+XrkHUHv
H0c/aGFtPv6fgJJJNEWWT+GN+t1OoVX/PYHCByC4RcNeTAYgj4i2bn0lu1dyQiU2
QtVXgflNwMjycPfmlGrpYh1IoDnaQC8EK9Wcz4roCh68YtO7/XC06UeWrP5uCAiK
3HxU95stnSJSCZoPFTIo2MWNFBlAGMBDzLURWQAilzQG+EhMzo2c2vyhHPnW40zc
Fq/nYW8eRne4o2EqlgTXHL9iIs47kVQQhTnrRQD0xfc01yAobqI9SZIGgqayVNe2
HoR5BbDXLL2Me2m3MlnPYvQpnEefp73VWmjishJ5DTUURGDImWZCr7rk+aly7EXn
lmfZIJuXtxsdKVgp4FiwkBdSVIMzJfMO2ULr3JtecwU=
`protect END_PROTECTED
