`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GFZ8V11iqZW12UvKYcGrAz5AXsRv9qEidn6Opk1oXpsRXTmZ+sPMsGGQXiMR0w+
Ws8hobmuTNpSspHQRzu8F/RdJoVeITRTJdP6PvXJdxq6eOiL5WX084fjR7b+h+dv
FO90eWs0fltd0pbnX+J6Zpvy0dcvQjWmincGy+aMc1g0uM9+L1IcLfmNxwxE2vpx
vuOVySyRVn3tusxuXq6a6g7L1r4SlanzqVumGd7Ek7Fbo6N5nfd2/ORy262wLyta
tcIyvdaQqRNb0sO2W39Fx/uVxQDHTBCJXo65EivzLoB/IZYwMtrucnvP+IynHg28
l8zBZGnlxFiIvJF5hOwvy1bk3yPtzJYy9xG+O7Rh67HsDqf8pPVt++rXvMo3p4hR
t2q8NqFB73JHDj24SylKS5lUL2tPUHyElNCm/utkvpKw9z0JfslWz4EiNIjZWrWu
61x3MT+hcSWVu5TlTgKGTj++gNaqrXitiTTXst9/tNQiF5XEESa5bo0ZgCZgRPfB
gSg4QOWwtXce4Ff08b2x5UczOJuN6SaLSQzUnbPTcZaMcW8tLk+ACI5KvZcIpwb5
xEvrLJC3bK1q999veKbn/8FIH+gCcWJTLT7IvndKxIM7j4gyhrrgpsibCA88XWVp
LHr096qLkS6jqJGy7k06IA==
`protect END_PROTECTED
