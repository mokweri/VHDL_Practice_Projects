`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R85EpIV4z2o7UIz3+ajBznfZCAHxlwEpVuVTw2kbXMhs76/T8xntfAXOgVpHYSTw
8xQ7N/xaN2SpkDU2elOIQ8J0//unwdkDbhWWItO6Q+xbkRXvBFF4xpe2STvT9PX6
eIsfwNFo/ULIjII2TA7lMbYloPZzddte+r1hZ/ykeCEwF4vpIjpWySg/NLlBPZlc
HhbjA4ZAL/0vh40leVXYNNZFVYqCnJ787RJkpmziHmsgENbDYQMKmJNYj9BC9mnr
ILJNIkE5N4DVErLpUR/UPI93fAYTN5ALwU64tNq1ny6gqVBmmPCFLB/0qpjxqz2b
DKu0siLFz97i5fDt0QByDVLssxQkwbKVqKGDKSdUWrluk36GFF3IQsH24bhkKG3k
S7isjzGDEE8rht7+3y3NJvT/QMeFB4FoFO8N/URMdMzv3uaAxxnYTtGxx9kGa+sm
1bEdjRpF+Z2nUyOvXT628AhgGdJ2xAilvvXUnw6MMw/TVIjJONw8ajTXAXIZiA4V
SNPzgxRGg/fXOyKDt1RVylB/ys+IDMNvDaIsk6JmZHsp/zun8IztTwUyvgKBnk9B
h/d4nXQ5NN6Oi3FkxdvODb0XdozkwJR+SYY/oy7ILmtGhu48K7gEHtC05Rr/X5qj
rsRf93PUG87oykCRoJ1xaVxVEvJKKqxGgSyHHwTFk9JTZ+/CGD5eyUcSQ4+ayrxc
FINnx+RorK49PBdL9WdRzn7nssBfft6W1hLsw4s6JTwo613sjd0bDrAmnWP/Uezt
oTCiPJhpfr4tEeRGbZWY9VGxZXwEMQbkmTWtmxGMHDP8cF+TSm1xwWeqReOaOUvI
4ZuDEYaH3aa78mqgA3iSEIKIaXzgks5SjKZ6xhxxeayEXp8n/gSzKm0+tgJI7AAW
udfLQnHGAeDKWzdtnMD/K1QTrr5lt4EXXaJCwvkAxmeIdSeSMbMQrRkaysjlS6Oc
bwdoRIluV5F4oRGDvJ3pQ6nzoUkV0VsgKtdMAv85T2oZi6N26I/xI8glPUVWq8K5
js58kM/vLPCeMmbNfRIdL+qFxejfcBcVUglLDbYCwG5rjKjV4/DBvaJ/zuKNv9hz
VK43AVeF9czWzAwbLq0NxZKmeQXpsy/VArnb66RElBspiOy2nTORWvMa6LQHtaMJ
1jp0yeDNYyhzwR/uYjoEBlVwdrcFdWNS/y/mOTjQciPsv0GASKx2pLBLuEjuZzrh
927m0wdJ3UWxrsra5TKiP7E7FnHFfRfpBNLP9p2aORAYS5/N64t3ar3A3hEu1gfQ
oFW7JKW4LqTK8XTTTMe2b/2JAX2wsArzEOtFC/71RfwPc+BixPo8rQR7pIiTJ2mE
LozT6e3Q3ih9JatwHm5Vwu9euuQ7f/AWUO2QBU0LTkuZ2wzXLC91Ba9+1RPJdzZK
KRT1GDBsJBKeVgrOdGrfbjtt1PiWszTQrSFgzyJG+MVuLGKeX4NPVot+Oe2z99En
K7tpzdBRiK/19SkZ+7EpUhafN+5sYVl5bvFLw9akT8nYDZQQ03TGqCZ7f0hbqoLT
Teen30Q7MJ2q67rcXuAf803Xlq0LESL+R5uLG8kXaHTWk/SbBhuQgaWBwNuPQ21j
W8sh+ACEPOL5pHU4VOvfTi/0Xey3tBFQUI6ZbvxlVXltJ8CWDvjUTIOhH4crBoRY
uSOJ7T/KzXH1B09/FjGYChshMPoy1GbmxXh4rc8i9V9bv7++ivtVRHN3GveuKx4O
RlRSAGT3e49vQyxZz5PhF5UoD0ngyPyaEOa5s0PNF156aFbA6oJ4DowqbJshTmGf
nZc48PLalubpwPTjYUhDHV9RDboVkgotOvZQ02l8uxDWHAqBXlKggR1uJFP1eauX
kmgvvVeh6YIlVo98I+LZH7svyA4wAYIaG8mYsmyl29kzljsi9LApn3ug7TkJXfL3
dz9J/2VMzNdIUtKuFB3NHoBefL6mi7JpyVGo5LY5STCwe5jG1sgKGnTxOuh/jdSo
rJtCckUTBAJKnpDRGShfzd9ZEY8Wee4m5AooqyMLfc7HsvGWNy0u9khnP0xrHiXw
/zw5/Z9SmfXFzx6/uAC6wKTn6oHK+OqHuiiM5LcUlEeFXRhXdw4na/IDVIl2rP69
SkV0avpdjzs4yIQqVKVgezHdA1hvTp907ZCZwp6AhM5hD+iSrKkqstP/D7ta6X7c
0bwavIbdPEZliB+Rl7zvE1dpNMVU7ltMdZUIV+if5t2PqWAr7HafjfDRiJZMrbCz
N+M1vvKOg1miivPo8kAfjAnpL41E8Q3ht5XmpcSAS90AOM4s+8/dIua1Oz8BctwQ
VGG89dh9DyNT0k67G6IicLHYNyuPhsaopH0yFHvi4etGFzmHOc2Dzh8s69NBPN7u
eLCp+Elh+nTxmqOpHVaPPvPxRNoHfd9hTfw1OzY7Daa+a3dTghWqn9hH/y/mFe+5
KW6zq4pKTcGHWj2l1wGq1qCAxoMywb2M0oelOQhTnt+TDJG2zsWmLBkrdguzi3zv
7OJTy98HkkVkOr/GaPbxJFyND3ORCjBIyyyLXamESo1Xmb+kRAnVNPQDxi4dNJc2
bMRVtj4mdfJpiByUH+DoA2REoE92fQHRPwFt0MU2xAD44eLdvyCL/0kAXtD9Bvgs
jSuCnPNqztK825CPurGa/qFBpoolgEja2Bec9GCd66Isi4IhsXAmDbfbxbSXzq+w
vyDAPOED6uKIxjTlDTMIfJ3xuY0JzgT11tIRHAXXOsS1SS+u3PCEugKpBGkwgOoh
NGpJgU+ZR72wSi7AxeZm2oQRRUgderwlrGvaleRV5Gps/2m4A1eULaAeZG6Y3bON
ROCEZe2Bi/YIo1vcGFinmoTI6upLCvv764GUrZVTvKIIFe5mzUdkZXVriOi7lvZl
qrWRFHmzDA8S16ErTeEexgzOMw7N3Vr9J2+N3E+v43kuWGFfN2tatFDd5Z1ecokC
y5msdg7/2E4Rwnwk6sre3yXUTOAlLmOaUpscWgQFQyfj8c2vcw/I+WMJdk77sWa0
0S/dMnFvaC+BMBo+S0Q04iERZkwjLZvCcmGCJgQaI3TkIqpDbMPoxp0RIAWr/p7p
QkMfSp+6WI3l4O/EcNfUfxM2Qzz+nLBlRMonilZT6GQ3tyoNCXwmueWIO/DcymD1
AwXrREsWqkXrUSRg7h2mQuGze8b33Jh4hCSREw+gn7mL5YwEU8liq3B51QLd7QIg
OmQ7AsNuoZwH5cBAUoCgTwkDU0XMCPKBxyUEeQgqAWDgHF5h91dgQdu5HyXZrC2O
wSz569iGiJNATzhcZ7nxtikvo8t/1DC4IOwJ/0P3kBwKescMXrtGVsu+ik2FDRRs
Wr90xqflFJo4dyyk4dfurhw8DNwMGwglWqL50kk+vCtxnnYhs6Cl1z6kZAiHZV7v
g8l2dr1/oTW2TatVAGbG92zfH/gIfnbVJ/eb3UqoN98YTUi/z4NP3fuBApDrpDWA
IeKvrIStx85EbPetyDUzZnfUu/9VuxOayVqYAtuhTO1t5Cun9DpQJ/oHVaSxzCc+
9FbLb2F56bqlyZ2tYv/bRvOZIOfgyhNQl68n3a0QowxxaCYu90k25P5liZPoFw+J
c2nq19XclMeUp/uArxq8wnD4HR6kJMZEPwPKW7H4OGF5Dc8Ulh8gbcMhqcbb6m4X
T8aXosg/LuESfB1LLKaSevFWSshfpebuWT3OBlbL8QKPZibr+JcGMnfIOp/whCt8
D6jmY3smYMaS/m3kY7cz8pqniPE2CDJDyv55b2k5gRmtFfHlfd9tDXONFL7urU7x
pqFsbJx81RX2nblGLRCl4i0NbKYSNkav10epArNI7ixiK/Y1/dp6eLqIHigIOdWJ
+WZJkSffWI0+/GamKTHdksUS6YD85MTsMnSzm8nLolFDG6ixVXSrk2Ry8q7HjKOs
/oDByaKIhCwUHAF4yULTvwi7GQzF2HXwf17O5hTsAuWU08LYd7nVybu+0GTXQHOq
dTd9Rfvhx0AC4BAqeQIudjPsOYN0FI0Z5zh6YdVMN2VshSkzbbwBOFhdFuqaHLyR
7XHAbuk5fxx2d+5/CxhsuUuxGnicrbgtbX0lpD2EkHPDERibqNaF3b41QzWpUece
Kek3b6V6nLne4sC2u2ZP8UYfekdR4k3xO/Orxl2wbrGr2B45x6IOCOP2EE0zPH0p
9kRYciv06/kwV0/k4E3xnO4B3piwamlX/1aS14vnEl4Ep9awnCW6FDKvLPJaLqXc
`protect END_PROTECTED
