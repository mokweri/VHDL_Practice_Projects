`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Zv9AqGO2PlYPkIwO9eWly8caBXy7SRy4N8KmayJgP3UhPuBI/vMWhbmNrY7trAz
ebpEU6FvdmGlsFR8hMPyfFpbwVJpjAynS0v5d6PzeprLWmuYow4loLo276eIwnSH
hz4H1ZmW98hTAQSvTfXR7k+LusONjkLwxmkGM13KNpjWcOWmUypG9xBtIEJRRQY4
kGN46mdJiyGacX5PEwEzMgoF9kKDBGqUArZO6I21bK4CbEss8lo0T5c95wmbU0by
JXVuKAMGl7sUwIxwUojBqFmh5E53JC+XklFdRgLet4ipUq+ZA5TvNVfFuutrfRAG
2DOLfusGQ/L78c1irCGVJBKhVbTM3Wy0DUQ+0B1rL9Ocn+n0ZD+wOOfHZDV3HJU/
j+rvwLjgLzk69VhuWczQjHeX3QAgpvVcIFoNWaxAa6PEQGurdz5/vhLR7pzDrYsL
NtKCeZHVrYbXfIO1hbTqmiVl7sUpp3VUxCcWPMaFd2dn8nurmS+03G+Jb+XnUNrF
QRi/lrW0KRd1ts7+6OJPKG241vJB/OTvc6qZq9pSwasHjZn8jLzweqsqS65X71kh
DVVK8IAiWacUDEKqckdvGZT5cKFBvtkz1Uc6ueEl35iIKAiDdLjRpkdrIxaSka0i
k42vC30qtQkEW+SymgBOlvD6fEEJbho15gHYzFKoIt3L9Nyv4zLL9daMtWleTL7A
Nsqw6oxy6YJECHm2IRKyPWaQX2tikspfPtXgdNDGNpwB0HWKneeABxNEGBVwVXI6
GSTJgbLvXmUzpJ5HE9LwrAZyHHlENgjXHaoBWIVDf4FLBeCIx5uprF7OQxBiswSh
darBBF3ZDin9YV/yTSd9yOYIjhFrJfZiRzlvKt3RChrMt30uw5bBA2Ti6PufujYM
cP3ek4JaBKnR4D8ni8ZetvHeOi54gj0oJvbicR1WJuiUXptlcaq3bpU/MGG0lLdC
B4/xb5Bx0456/jxeDPmsHSfODN8dTnXVo6163+aoYJKoPZrOoREwrIwpP4T3uOmq
ieYw0vNcI9iMSyCOpIuu3lGvzcS+V99hAVlO2nbX5ID62YXs05FfxtuFs52wVQbh
FK6qjF5tmMX6bX72hibS9dbg6bttsSf3IGm7RKu30J6GMRVLnTRjk469wLJrXC02
pP7SGN1OypXToTIJJV9FCtdrJQTZnk8tk5xdnsxW0/sQVUAuGQdsd0AbFFZ1zkLm
Bfh7kC2oqQmwQHFVTMng3jlXZvMof8TpFVDGP93BxaCBdX7VGDvF8Vydk/TlOG4r
WegjjWclnwaosZIPCXSaJtyJlFdv4OpWDW17OkMCY0uWnxp3Mtmt4s66X4lbwyoQ
MsBJ979MOZ2YnJ7LkIKB1QZfOkbrw/vsYjqpOzAu2nUC+XhaXxuPbwv16Pjv7E3n
JxtTyCHGShEhD8scgXX/K67k0Mr7vKI/CISwQp7Tr36EAhK9kOxsYwGOFBJ1C2L3
/eWWtkuIKhG4qM84FsFCQkGppJPXEmJs5cx3KSxvWRWwWsr9ahtauyjM4NwO9tHc
MUN04syVMDoDNMdgEmUZn6R4SIMBOLsNnuHSbYzcxAEvdZZ0FrUnGBS7hNz+an8R
ytHMfVoQH1iDVJanikB2XSICBJ3ltwc9tqz92re2V3/jVfVnCCHqExTT28me5vYj
ZZvjRU0BQzq/BOUYIgaxpb/j9bqk+xApfsesNCWqYRPox0VFEj8l++1UGwlWh465
PALww8TtA9tvKJyFt0t4sO4LFvQimattVPxXExzlA5TzRTvMBNN/kZhP5Js7bXQa
WWKYAQevoyNjFYQwKhEmf8h13JNeKawU7RbnBQZ5LodoBLGArmtqRqDfNCstjy+U
I0NbkTTAAWmo0CJ9uAKSha2svdF/FBtfhNw37AIcG0DbbSalSVmcOshshXHJSxp6
ma/h/DTfBGPkftJ0sUQJbBT+H40zUVQv1nM75JRuwjACFjeWhKyBxx3sIEqQGDqH
G7rBFTP1YhSq0JFi+FOLgLlHRXXMk+sxz8RLse2pzLuIQWe87EQPN63NVkJSiy5Z
ySxP3N8PWoVGV14SFuoJGOaO6EYwCFGcBGStQDDahyIe3g5LEOsowaZel0tm+NHt
F5oloZNbGnI4XLf7W9UIkG2YNcGtfggcA4dhkdaBN1lf4KEQ/YpQRYXBlIosXGKQ
PhDmy2imeTRcryvnjr3w21T/TjNSIB9BNgTyYSQ7jLXa48NxHlrn/V6fTjcOQ/pY
mB8qrVQolgLf2FILtf6MO8GtgIvN31574kYyzvUTYJBnvhdOzcdPGxjn5gpMNctn
f6eAoVVNwbopYAtPEgH1kQQavOp+ZSwi2qoe27f0vlBZ/ecV/B3Uya918++gekUX
h2proKMN1ldFwlaGlRwJjqvsqeGZooejurSlLNk5Q+eddiCaYQuMHy7JciNuk/g8
e7Q3eWLVjHSYWqUuJmFIg195McSoSh+8+z0AmDmjZ7gpHwcZPI+2dYeQjUjKHPsO
MT7lnvRJVZL+CX5ga419tbtcrKpqHRVHNFDOQ76iwAs5HkcWj/MWL0OSZ0wRBxaM
LJYLQvSa9u2O8fjPSOHqc+OKBxGYnyGr6+QtrYQL39Z2SukaYS5a1iL+VcV4622O
EtekvkcKsnCXcCzDB7lZJEaP9C3ZWla5QXhk5ksGfp6cty4Q1oEA3UgaLQrIrOPE
OxOXQfNMz0ilvf9dVZenhK/Bv8N2TklBPrDvtAHbCj3KDiAKNOHTTp0Xf0HkkrSe
+hBm/acQ4HSvt/2LRo1LMzfmJrjq+FSGufSoeI1XligKzbO3WwA2JN+HKVD160Fd
CtEOh4VMLF6N0dtrwdfGIxHD4a/GjnjqQpRVZqVN9GJd3Tm7wCt2crUPMgUzWqUA
fkqXEd0aYMoRygW50262lBYVHeVyZ/GoqyAyfvTBlYKRkypjsiZCRRJ+ThdBHK+m
wiAy/Bd/HyxLXqsOFZflr8wzGbMgH5LlUjfat7rtB4PsD59w6m+N36JSBbR4fssH
4Pa3Asc+7yEeu9TpRoZixE7WT9WEXVBGCI5iwtS2EB62OrvarTsBxeSFFnVtgWMj
+9WptQIzifsOaJ4V9knufODyyas4HkWpqkGbugEZ9YAOuJoC5C1sQTbKwBtHuoq9
6bWBwIg8Pm95o8KCrs3OEGb2bPulH3l7ZS2bi7hAXDQAu+NdDPIlsgrjEdGSOB8O
YqBbLh7M5muN/TDyQyKu7e1MGFoHpIDsnnnt+UiKhpJ82DKfHtMiRtPuar0DpSb9
S00hVB2rV9E4Itb7b9WtTRMCWTQya1sPJ5w8o6s0VXemFV+wOMJ/2oo3txP49cKN
t+zDOL9VTrwB48lPg/yPOlnp/TLTJgnjxDVJs9Vvm8eBnvunPCmbc9+0APXaO35v
GFzvtftpuhzZHqkCpHp96MgI7AWxf9U8z0hskRu0kCoTO+o9QJWBkWDVw9Fku2HY
fs4OFX4mtTXKRRYh6sdb6rv8XCHubV8o686GAO+j8tnuzSM2VylMIPh8943UkQ8R
/0fogxFgWJ8L5D+g8T5jrSDQKDxGr4bNPu5EN7kT+ZF67euH3JhuWv4xmAJFp7EB
mYrEpy+Pfs1FItUh9+cGzfm4EeG8cjZZko2bp5hUFuYAOFD4t338OGs4BHpifc+E
uJkIoWbZedj7D9Iw0jRHbE+qy1nwFE4aWCo040g9BiHei9cCGd1hxF+RzYQ1x4Ex
`protect END_PROTECTED
