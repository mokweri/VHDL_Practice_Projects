`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vH0lWrwj94OYEqwSIr91JQtkBu7964RhVFUycTMKACgqk+NhV8u3Zn6vASAHPHN
AKpSImQsk7qDC0j6kipDv1E+5F+RFA7f98Ul3V49HklspBvUNPr5+1XaKtLIKA3q
3hBSrKxvtLP3aw/pELPwiNzJXa2uAbjM86HSOsyCuiWy7vbqpVnAgCYdZYS2q78N
J3Pfc0hT/7aNj1ljPI2GRw3mSELYaL1pIgn8x3yTibSttNQXMEiqbOmpR7VQU2aP
UDhlD1zmA+uXmfusBf637uYpKB56kE2UDua3145LprxoSQn40ymjlRrSQSA7Fxol
0V96ZjV27uCFEZcb92yql6doAUCYJ/N2fHZeA1egG2Ond1CR7qmeeEM47+73/FxL
PaiSk5Dtl3Zq8iZjLEay/mVjI6Ag8YGsJdSDWP+lzAX/squxbfeezSrXSNzTwnKz
2eCr3hzAVCjaCIaw1elre2vEqsBAWDBXuPhDw/Ub3lRL7pXNKy//8JtDuedgkUf1
Tre890bGmOLNYH3QgoLeY/LEF0R5gKwZse3AzoegBUaMI1GYQ+ktC2ECBfKQdcAK
u1XQGJpTDwfQP6x/kCq64EJoVTpPS2/CbIkTv3ll8COmgaKtf9VbhxBMupZWGPGg
a3fbfyICJEq0D+ZJy4UYbMhrFsJMpYT77BVGH1zuS4lRJOq9eEpO5hI0ylNm1zbu
0MhqacrrHLn+U/foyEl/0rxrC9x6+npTNp+tcLcFvCIRBPJzJBnlTgRAK2du3cS9
ZpdzehUj4FwPL9zOynPpngogEnDwxEboQxeKzCypiLHlIUSjSjzjtrStwJNV6Qxq
7OwzL6v8++z8HW4PeySIAPFb9KzEq9Hhgv7qPQBBWZ8wYCXpo2gsiJ8B+zxWmeA9
2/7H29oCzne9DJchXu58hzYX73cnapyQiJNzM8rpAUpv3pAXQ/H4uqeQpKuXDlwu
ZdITqOiR1nIHJ0qu3UssvG/0gtBznGOoOqs/SuesRLhEijyuK8NWojNxt5HSC79Q
4G8Y+naR7ymq1xvtsOq7RUK7RwFz/r4M5EGAL90S/29pXLAamBsP5ozxMlzM2rVB
ISp5VSirFQ8jCR6RXXuPrOwbelM/7WornUajfRAnUV10N9VeKw+77kJcJaGTjQwt
JguU0Q3jGS7LLlrNW8oq8fi1UASo309A8x0ncqB6UpvySHtZltdqdOOftBrMZK0/
vWOFZrm+B7C50i/PZuZ4U4Nw78dXc/djSNsPvMt1g2LVg8p9vppfNCtwl0Nh5sFP
+4LahrT7RnKKx3ulWwKg1ZYO1gBZ7zD2p4haX6QZDD/QN63IC3Iw6N2BoXdEk/Lc
4VJedRE1HiYC8vkSQWHzwh6+zLvr23urwZZ8nJiD7Zi4H8YNfOrAtCWpeR15CWh3
RXoSOMzstUH9Aae4lS3TjMSyk2ybNrF1ZZUli2GXmfceBWtN8Fnums4j+IQAtVUZ
PueCYsnDCqBhl4WVM+UIIRYcfOKDSWYWeDOWqXXDQBXiH+NElc+GsgP5zAxT0FQx
3rr0vJWxs0elLlJym+YumE1dm+4mVV2g/ENZa0NOEaK56jYSYogz0ANY4B/+RSxr
FC/oXLtCPE/4S6+RKDM5EW7BtOO1psGVSF0mzC1k+as=
`protect END_PROTECTED
