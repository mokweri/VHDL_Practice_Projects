`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4w2zi0mHov670GQz+n1KQhxIv7YdJfhBBqTihxScSQJSXvjPcAD+Dt0be82MU20V
Enpk3nmln63kq74u/G78Z3hkoQGh+rFqgN6Nraf0Ptog57M7/EfZdZAu1ehxxbQp
83AqO4WpQ9pPSkibHyLBWJZkcPr0pNjsW9EH+at28tM8GIIRkJt2eXQewtgvWVR3
LNkbTX/dg0x7BEdzEKt/yO+itMBBggyKOO74ElOIhLpC2AlR0sYP3jDm5riFnJq0
OUpmPSZG6UWVcS9bDZE9JQXvFxKkBDqUAFxBEHVrsgZbey5vke9BaTL+gOyKwEmZ
U0ZjSz+FhzgE0nOXyHD5+VVNkHWBxLTG4ZbmeIlhu1xfli0r6VXnV6msD4fCjqPF
7CMKn0onqSppAsmGfCMzlIm+sgkPlHAUiItKJbj6uFWx0flhZ38c/1svSZl4s0CV
b6gq+WlIwQgWQjBZTYdNgFieCb4/BggjKQORGELe58cbXp88DhOQTuOg9qCHweJ/
8NTw+UQoBG+Jajxvw/1iHGQwxbAkQTKvWUaZy54RkbblHc8zx3IIhBMgZY1nvMj5
hq8l0oLLbVhUps7ieuJ0ssubJcm8cp2O8suTDWjVC6l0bdSES9nyM/C7HKOOqw0P
SIIdPwfhGVfiVa8FWyBi5wtlXSbguvlkOm6CRt7UZGuCOdg4LJM5v8QX+WxYPpAs
Sxj+PVmGaIbJFvs12yHjwb79bMDlAAIsq4F6O6LwSJz3f/jMc5CeXk4BkZbefzfv
AHo++lCYo3gzB0n+MTXoi3NVUpnelKyHPEc3Bih0wfcBUOhKKIXWlgT3U9gYiyGC
/SMAIHnTY91GMQDLQ6fqpoPwmx2k2sVWNO7yAw3WjcUqYNi0v3DrMDa2Cm5v8e0z
2ihkC7IGT1PkvcDv5Tn4hvNMj/4qZHvGH7VxbpZ6j/nZQwgeVGmbnyTMhyfAk730
ueqxf1Qt29XOyg2JOcAk1gzXgUovQwwutSzuA0jljX6aO20hTwKsjYRTiQknLOAP
lNSxODE36mUIFwzg9YlM5Fc2OPhLnOeW9Ha7VZSTRJmsqa+tNQiFOwaSkH/b+Zy9
XQ3FX70mfNGq3UFfEN7alliWhRIJnM5CsEWvRMbUTOEe7NTmlV1szRPVtvuqZOkr
9Men/YjFP8ssSK9XrEXy+kB20LO1mwEadNopEXRMYuQbL763w56EaaqCAw5ShBwy
FIOhayQOMY20begFtG3vB3jy7LWW44JtMf3qfjRwr8/TXcnuRPgR6oRhSQz6Sg67
qcGExL5GjTrXfbJC3QFlbeTRzDV1Bz7IlctfGaHH2dkUSZKpmKhb9i3uK4NmbcSt
Pogcoo4Q5pK/KdUi1YhLrji6HTQZNyjNRbacjBOyL+CzZsed6fF5bvIu89cua1WX
J536/jQZnM8b+aRQtTBTqEAeAIMcrbkKhoe7eLZqKTKkQr6hiFh+Hhy+t/ko+G0h
tDGAEqkJBOSn+XeN2xDGXAhCo/RF4m6Z48LWJdxHSe71EuMke/Tnltln1SWiSFb6
XImoLAbn68JJSVnE7U3/1NK5Du0R3QllEFMnD6Fa3/G1NGiPhn2hWp9XM0QJh25I
lnGjsvh6xuxIU5uniMknQV+NcoHYHMp444SsvjGLM9j9mTHJPwkopBKhA7bXHuvq
uN9hLLuVp0Eo78sdz1rWMrEu7rTeO1kdtBOpsYmaXljr/XdddZwH0E7QUK8B/HUA
juQZE4Ms3u8UonMIlot290KwQ/RG5FkiZXpr/AetyRgd2K4wOxkSCdEM3fV39qNZ
DFLpURLyrCWDSNekf9h9NPf++rQcVmFUEhCG1vZgM+0SiQ8+cm83ux4CMLRNPwds
lasJlXgbgCh+2Qn3M+IeYfatpCtrcmi30Qcz3T7C+XYrSOl85FBV2N6k7eHKddLy
7OaqxL5Y0yrHxZ0j32P5cmnpSL98Ezi+WxzMewLh1XFEaxVyv+bADxCJEB1Ba/qf
b/iNkK/xxwO7mtTyDYTgAPZXgi6CjfcqaS+ObfEQ40oC3ak3ACuhA67zVQ0T6Wj8
WLMcHEYMtt40T+D5iIhHr+EXJiWP5toAKkLQImkYSeoTWEcIKz3S35oyDlOTnU58
8qHHkPCTavvCM84MHHnE2hGUIHyMINJLAJPsY05BJFIFC/GthDpHkFpsCGgDG7nY
dO7qv1JkoMCNF7N8JEO5NLOm+GTuNeOZm5y2MMWDNNtB9l6GL4cBQeFz2tXDmRrp
w/u5/bH5yHt6N201BrlQs26gqI85xcjNd97k2MMvcX4mSpo+GupPE81zjBQiWuBR
2bBSZD28DFgQpE03EoqQ2c8SiD96nZuSsWYTFDG1FtKIYH7zHm7ih6i8CzH6Lb/N
cyQ9GVbFqTjSTvCh4/MvK2X5p5tAAoyDmaUBCFLraWZse6QcDV7CRZK4xdfzU00a
sIO8SUSxfLNBL17NQ4q8W6Ogs1YRMaMEN7MOBJQYdsf2lijrX/baNls/9x8kukET
cuKz92D5znd98ridlZ7GIOjP3Me+P4gtVh4Ol6ratYMN1+/j9fzQVzSycTavcGt4
xdRX2E4Di8bAU1FHsk+0AeVQlpAId/Rb2SNCrKRJG41XNKDhh5jlasnXCZsxwKmO
7C7Bazlg71TmLiWa3+2ZZTBHLMnjqEgItFWpttIUubCmQEXVubxE0ughoh/R4mWH
LayGFDx2I6G0Udxft41JAPudeW2Ef7AQ9QItKY5qXejgGZT77ro+06GoBCSgIZBX
q1nODr5H73HXa/VjSwrfksqCiVgYktG1YLjCVtnacT9RmBIu5c85vqtf3dpTtIwm
zt2D/4fE2uS6TWGRE/Pkmp0St8k6DodIQh1DX61SMsBZ1DunME7xm/bKeL+jIvqw
/9liyUKtBHI5zCM3VtrezwFtmF+gdGW+zY91NTm9lYdUPUZbWkzQCIzuWe9fczG8
A7dEWjAi70USifHjQofD65j0crvrZAlMvIdug7TVL1alXo4eIsYC4ePfCw3V73FW
xffvCgcaoEebXuOWuXZFzvMDtZ3kuTk0buxSlfJ3jr5pbBRTjgiefmw2x3s6ifMq
cSqFeCWPe3xGsCJ21ndY8d6ArUhFQ84FAvkVpmOpVfpWV0XJOO+sXfMoqt2XL1gU
GXowH8FDalDEb9yyD79xAE6HNg/TdYHSOA4H0M6f2s0uUFIZlltGcpiflqXZLiuR
xAziDVrF+Sq7tLQEezuITSyR1mfujBTKlYbwjJp4ggVT6r7H6bHX4vS7l7Ne1DAe
8EblN18zElE2AoS6VNy8GRLtyGtGxUp6fE9piILH09HWhj9U9Bz15u/qHmaE6HVz
vbF1pfjEFsvpSoW9zrUn7odlDIX+H88B7pUAoBpd8GuJTljn2AJX3ZyO6tZnCeEU
RtkjhL42l+ZsPTFxV2UdquYvAmcGiVl/H4/mIsDAzbNBa/ii7+MNEn3rXhhVZrgH
Q/EqBdfg6b2lmpTxmX3ArhJdyHvU+I2fIuHE0gbALMP17etitnlVemrtP6b/hB9k
QePgN3Z4fGTWzF/oABPwUIATJsEA+LBBcHHfK3JJEr7fWJdv+Q2uDWRvnAUftwLZ
byK9l3W6DPC0mtzwKMMkqBsD8iBgRvgU1ciBCuegmds3DZMCLYxbbDaoUZ37Ytpp
H1YqG2IFDsDUyglRQHNLJT95079GUhFSEACEiYv1242en7Fx9Z+ARzDd9SXbyySC
s/PNZu2iayZnmNFJsdZ6o2lLDvI9+WN59ddH8hatsmNxzknOtkfgZb+5JryIPBrU
CWddHvlfX8XIP1lBXbrXfgrb/HwOkY9Ucufy5UE3eqYVDuf4SVg8G7KphUkS/enA
N1wnJBLh1a4CbqJw5ihoIThPBzeUqI+0eTkE7wI6O/zPCb3No1aqeSbsFwo4soAm
vuKFYlEtHUGzS9P06HMq7TOv4KSRCPMhhUY0zD2jznEDcRmKNrsuVomWlfyatnLQ
7A8Mq0/2LMBRt8iwMF86LgZSPmCPSQGAiGF68j9L+WKcqR38cTeEe8prvH99FkFw
anoDl/j6wEp/afqaj9jrmd5/iN4NfZxd5exUAh+3KnEhu38EJuKefUiZD7iLvef5
kCoUkeKajbJTrSj/75ILhvzYpAH2rCeqdmhjfJ/EPmDmBmYEa1J4OSjdGCXjW0h9
4IgrF4CCPDZnR15+/ovFUb10cqzUjc4f6x7PL5GyPTTY3jnPNM7NmJ2MPRjd1SzC
4W3BghvT4OscfQgTncOAn5WmPX8/QKWJnycFkjf+XWV6q1fC8Omk3cjgdB/p8ZFD
MF+A9LTADaPxb7ZHykEpHDCYIjVvLkjlO7RHw4n0HrMT3Dov4zr44RkYaFBo9nlW
60/MXCZrEgFnt2gj/b1mTrFXpCgU4PlugOkAQSd/7PFAU2uQ/vPssFWcz3lmS4nV
sv/V8wL2QzWXop2oKUxPGukRIkXA9pfSuZkPbYIjWDfFEN8NoA1SAA3vvMGKPhhy
Hzm5Z0S992oDWbOSyaeZMjbyyHr165e6ZjiwPkdyUGHqN7+/Fj7ErW20/bEVy5Y1
hQlQS0OBsLoSHtbmHIoc41t5lE0OIhcTTvcoMBKAuQMBg/SB7WmuvET0wgoNQ7wT
kqAYWyfoQJXjR3n/Hr7FM/f3gBmjsuTham3w1KuGerTs8xA0i4FzZmtjbl0BJxJ5
x+8113lojfffvApzfwaH8doHDO7qAGyYBOMrZqCJ+b7v0fQVm0tG2oDhksvMewf5
BN+yDerc+5Bl0QNsaStGXS4RNCtsd4V1bFRw1ARTS8Rp+9dORh/sm4JjQfKEA3Ui
P9Ifo9qPZ9uASv/cGHwKEkJRcTkn5vmBMYgtkGLicKm5l7PuIkE/dEQH7KEARavx
eQm0SXpz4vXgFlJtO3OOXNStjpXDWCWPllhGmITbjejzB5pUoNuEW23JzenSDmOs
HdweH5dU4yMs1R8Dp5Cm4q8keXhnerUDzaUCYmQ3taUwDMgtWu5nFUmIIrlG+f94
68PIsN99JqtJO2HSxdDOlPniQCrYmKp2Yi5o+Re0mBLvQLs/d5ex72l47mWAuGHn
Zwu5W6FuhSfIYRRl7pXK5YxomywEScp+JTN6sb9f6sdGS5oJJDwPQLq+FqOlx1ME
jmHswAYmgQxxksUa6zWKkPUYZEk1VvZzj4+o4yrLU/UWdH6jFXfBD12Zg06XNf9S
pTQBBouOCRZRpC7+4z50DmyswFHK8W0ouOLlSK2F1/ayAG3zJSZW6PBRNvGyB/fo
6AF9VsE9xhaACmRy32PaAXnK01h08R0aJCIsmWpXViNSLTRYtU+6GjZUxXwT8alX
RGBOln7sJmsY10ugk0lVlLNqRfNTJPm+Q8wH7dve81N4qkrL3Zo35/DPaM/3Bbb+
IBD9Oxf0tIS/bsG0p6Uz6H4UMENUlpKDnvzLWVcm8mrK3Qip3dTw7DeLlsRyaRWB
eKGkvwIH55GhsW+P1S8LMEdLfqHMrzG2Lt7ueg2vMFzZgxvo4Oa0Oj+mh93sayXD
nR6fIaXQ9XQI8AyOBgyI4CzBpprdRHmJ39+FLGc+zFlIFgTgT4ugGD7HinFFWITQ
aq6/L9K1PlYyIV9+7PQd2gtBwwZe4hpDZ+3HZyhK2q6dp/jjbTgI2TrC8OUquICf
FTTVUXY92k2MMNnRj6EAmPtijrIIXcIRczO7omj00DeE9YQCEeDuVx+o0iZ68w3y
zC9ppOQgy2rDqN0fbJYnV7dBEOrfwKEAg6AEaHqp3o9I/ayOj35MkdImpzqN3+VE
YT+E6pVeboaswKK9T9NkTgL7jdgHZ/v3UTsZscKOCBrK8sDzF1AWgL/dPxlXVdrc
XYbAiwc5Bk07GifRuhv/RZhCYOAhiG9RnGd512SpcPRQAWnmyTDtVS5QPKLG9Dqd
p47RpLV2zFy52m0y+gRPKJMKa+T2cFsXohAXWN958k2zQoD20rko5xRdeXwv4yW5
HbaILl77AUnq4Ebyt6rdRMXYdM2J3yDQLkZEfu1aCa7ttIbtmKPGw82wp/Ad/YkM
UHdhoHC8otTebX8dbPIP0pnJ5/2ZQ++7LCmbqM7SFBgkLhKVDp9TNfy9Z26xqZVj
26J/ykNCFQwgaHAT2HQ8LPt3vGJ5KLeqqYehs0ahgLfW1K1y4yp2E14vpKxPGuIC
CZlU30jVE6pR7xXLPCAFpaMRTUYqL+oaMSUkUz5GWVcVnl1homHd3THfZSscPeua
eeyyJlWpH+5nH74F39IwXFg3QtkfHcy7K7CmUUAuHUrGP0Y+JiLxtI/CyzVeQlkz
4AAOqidyg1GezzMOBR1WfUunmsjGrjB5SF/EwZemtjwXRNRcYIypcizKmJe3q0eL
6cYxf7Xm+bdkq85xQLF8s+H6eyaX53J0NTcODTYkYST+WltK82OZd+1i600BCsC9
i6P92GUe1EFKRWg7yKfb2RwJJo6xUkVXTWFdQ7V6y53cEPPGCrcAVJNdfrZnKt2T
DpqcrEE59V7+gHrTmRk0r7KLjPBi8/NUW0I1fze29ihFST8nw5GGudg139YQE3Uy
Da68i6mlLM6RHdvmnb7SXZJZ9KG2J8l7L8ba0MJRxWyKPrvunI02Ct2v447GECGL
A77EfN+4QeNdiYV1jOPPjeSs0xj7e1qz7OQfdw+NHrmUJcayNepjXmpT85oQOKsD
kX2KDVIKAbw050pFT8PFaUOLCGDIuxcEMPp7xEGSCKsTfBxvH5HXMO50QU0nYzEE
0eiTYBSGVT3GRARbuHkgMRhV8K0JuyF2oXOq7HJqKvnvxzCKcE+1megW7gCnrfnT
qjr8eyFPZHvX1iZzNZ3Gxdy7eUF9xnTuquSr2QJtgb12tbKsSFtf1q9mAeg4d70P
pgxV5M+mwzUV+0QxMuJvmIdW//QG5/zrG2SQ9B3wIxYiKFaErCTL400D4cNB5wf5
OUi/0wnOS1Z2P92Wpz78+UZotDRQE+zC6Makdgw1mGKcu/l8z6iKZ/yYHw10ytSa
fKnt1KZvNd/dQ6FocFKIXZBUMIms3Xygo2qSodbj4o6IatAXrD8fu95Afjg8IOz6
K9Ci8NkYCieoA7S1ktmfeCJ5oDJSLd3wlBJCG/UF8hJkitXPmI1zwztLAaiXlG9D
eWLE7Qfzub7NnV0wRCARG1rpffaS/YfQZGLtfQ1bCvwhsM3eyiOJ7zgl20Tnl7/T
Ni4vkT7kgDeo1FfSAJL/eViZu4zPafpWCQqULfpjF58bgBz+M4gkR7D/JG1wYgyu
oLW46znmy9Belkh9pQXGn7IZJPbNAk8svIMidKNLfMuU2W2KpuxPFwc/Kh98vFZK
SofURLydrVp6jUYTN/YA8TDjro1Af7pJKSjKRnvFHDi01djPxmUoPAz4Xvq3hOhI
Vk7PMAb5MPNlzSFzgQgWJus1X7n9bpzKk9k/8eOLvFMNJDjo+iDDNONWza9nnYF6
D1ZUN39OOjcDnQwJUwpHm9Jl1CkVEvXkeOMdYf04W9plkl6qTYyQePJ0Xybwhe3t
YIbw5qrNm8f0wF8Ep2NKb4IZ+PbsDN7afQCALDaGy3k8tbMc7qdggy4qVlTFseST
vNMXcvK0n5gLsbF5syb/1Db8zeItl/XQ37f/+5e1UFgSNjyt7tcr2Kw9uLbVoFy9
D62undW9Vi01gAubZM7O6RICAuRaTdUZsNtGSvNa11SetQPqnqAalViP7gmUxtv+
wK/J+isboRU4v8Kzk40gSiYWhZBv3sNUpkbhvvy6PBuG7rPbWlfgjkd28pDrURlu
fq+am2ewA1UMyE0ao0aD6Aym8wdhfveTTmgkno0Y4vH7xUsO7PNA0xhp5X94Yipu
j82Y3g3DmqgLPDwNPxkXWoU6Nf6pC/RXEASZci4dXftBHG9mS/NtSQ/ClDZ7m1mu
efuNgEuTvvWD+RFl87DiO37cARb44lxoKhuwhGvNACCogEoxImarrGv6z6iUSDMn
P7O7zrsRhWA3B5HNXmePYb1bseidUjVIE6YnBrQ18N9JsNcj6wrD7qYmFTXWyCzR
RcI/CGhSf6U7GFm/i3n3tpMXGk4Koh+M5CoSokQYdiFsSC/RnzBQawigfNEpUzXh
Ox9SS6PVxjAPyTtAsOX3CuGe04DQpCek/cN7owDGEWTn6PzjNn+3U/DFmjA2Pgtk
FLHG0FyAikKxvb9kAmV2WOV3AqIPYJ0UG3go20j4lFB94Ev63jbRuGXo5uX1ubwJ
2nto5uHZY7vNOYKhBPo9anddc49i4d3Wd1fpLX6kQcMe5U9sAHmSmn9r0pr3KYta
GKVq8vXB0txBzyfple50Fe8xZWASCOUmDCu+S7EFuWlW8wJSd3NaNTEMEctbdZt7
XHGmxyco4CkeuW26cqOaHIajDoLenoei0gYU+/z6OYguQNkQkYEPuBduJyTbyUag
xv8OmiaofLWXp8bbIX3g28/L5ahU8QdNFWsLgFf0iSyv16eEQ35uOXLycBEYKw7+
3P6xgSl0OvtQhFcGTvOTujWmsggnEYJ+SdzA6klVVK3znRLNM91/jrajftVAe8XZ
TFfltGirgHwBR2neB9NzxgtexlZk8r79+4pYS06xd3HgWp8vgTOJk7HM+TJD5QFz
n010dDVy2+J+VwbGXaLj5zhPEC/YUnf5ty0awkx8jRB9/YBYWNhXo30HavK6qJFl
LT9ui9nFLSONGD/T1ODCHW8J/CcHZcEj2f8+u8gEyLGJioIxFhxltRxq26MwpgMQ
tRIUVltV7VaRejvXdDmuJy4RWCHVi1ow3gKUDWSx4ciJ1Z6TkxWUAl7EbnoGqx4/
AJAdF8KExyNkTAXw/qi6sxJ4SM5wnoGhuYeglEz4Tgf2W+N6WhH3X6WEIqtQkEk+
875RA19rJJ5M7soe+Vlgf1NAWdeG5dDVOErQs+s8SArXXBQpwXahX6Eig8lhp9Me
f8uddZ9fwGSOO7qlggk7krcnwx8ndO/6Fh1w/LWqgQp6++vyj9BijXi3kEAXkNWO
fvUe0Sex/DRT1/xCGJHWp4eTLfrJLLFrjVVVAmZ9k9NUgUsTopG3jNZlMc/nm9uE
DKElZneC9padm/fs5ziYJ166Y9BqdAM2UjcubOnOB42vnnjNLfgsaNlBIrBWOEQf
6SXCqZmcwKUCJClkvDLlNtR908G9GGL4yIHH4xddPq+oIeMgBqhbMAs45L2KIdVt
rqR7jwcRTufx6rjs76SAmND2Y1CZedVOT44i1gg9eCbABJaYcSQz4LV00DqPCSVa
1eSUE4ziCtjWCFkvNtOV30rgY6aRtHsIpdEDc1RT18NdoLVe43BckUhROrcfABXr
hY9Dq+UIxVqJIraOszinu1J+U6A6d17lGTCl1z+NQ/2T5n3PeKzf5WPrYRiROABM
2765/9nDk9g8aGtQI2qFyFx2mwdzH1YupnqHERMoRwHm6rM2NCG50WKBsR0wXAZn
NklsOcGJLJ+h7e5mqKQRWnxLF+WvWXBzjFmvaQN2jlLl5JKWJRBDpBBygvvQkLFc
HWD8tGtrhj76A3Trh0k5MzCeyotoxUs8S5sem2up7Z4iQ6SGuG8zxHJuoehNZEBi
pmNBrWwE2U9tEXtxeh02DCGxcB8fp9jTor4umfCsPhsZJyBNK/8eKWtc4/rukaU9
0EkobarvQHU/eT2e2RuI9ZGQokid1Oeoeqz0gn7MtKuTvAJaQROd7Y7l7cTxcqrH
Qx6MOuQJtTrvEXB6eFrkfi9AhGthO5lPgcLKDtfNrb54tA0f1ZI8PhmDRtFzrgyj
dpNLQsoTIHG4/y8PGQYl2fqDZtW4rqJzDxjw0o8k1mStoS1/yVL27qTsCgILjXs8
ZpC8wajgXFKT/3BD1iHoxBOu2POw5kjyntnGdJ5MCLwx1+Zx3lP4OkCC7o6tBqxw
eahSWbbBYYrhuakMSaGaMrOMCaWD04QasIEgZn4j66AcAGvgBdTcFm/OnoAQgHR9
4x5FUBGPqy/RJuqqBcUQW+mg00PMkuxUnH9jVc+lNcpu2E0E80Carr5ES6SmXBRm
PAuaSX3izoHv3E+SMkzT20cNJj3Z2V8G8c8iSIoZJm0iarRv179vSiivAkquib/c
9Fj+Bue7e7p/nwDVOqsYcOb58bpTCdzIL0M1tNP1UM6OecnwzILjvR+s6+OuBzVq
v9yrMtpiSo3WnB1u9RQ7jwdvOJ4omMxWtCsOgOSC+9XT0okqfdWCY1rpmYrB8+pf
NTGmYCcxhYaBqiqzqGa2pmNQY/frO6K8z6QWMY9l5FSmrEQnO1ebloGgDCoIAuhR
g3PvQncj9a6ELAS4IWGhF1Y3nAw1GR1bU1M667sg+5UdQVX8jtu2cdWWuekozHEV
NPRoggC0e2TIepPGqmZd4Wwg9c79B0BlZ+hlvlXTu4JUzu+tR1E9fT/ZZBHmCP7m
v20AAmqnR2gUF3giJNmyDGYPEaTAV78zpa/aUFTubsPFs1nhHKe7jNyW15aroU0a
MyismNE3/JdzcBGaaKD5WJsuE3wAeBH8UbZp9dZ4N+WIisGhi1TVvPpZ59Ftvdif
AhQr1dGuIgM1JfuemkXLhjVp8Z0a0IgmF3cGeGu7VEWBvNknszl5A34J50ASPkv3
UEGkLNkd5OSsuKlV22nE/ybnfUd9F0HBNXH+E2u1PMuVEvmMBIdfsuz3SsJcyZcY
GvAJFa/H04U1naj78MrgH65c5qOzkpH2SyoE/Qa+bjHxX69+Qc3AbKdYBvzhGuOf
ysSTHqRz+49CLE1/WtKf4GEbykbH894CASKMmD+TWJwV985DnfmOrD01gEa1aaJk
/AAVzNf3opic67OL49qB2UHAOX/3U0j/tAQHCY2knRHZ/pRDpQrchXh9ekOTBz3K
8daqoJYw/jsLZT4UV+lVTz5D5nPssYcqmt35zLfZud22NJ5n7R12VoJzW3vO23Ac
m1znl82Nf2iPNgGD1b1Ou+A7aPtw9ZZxMG72lLw3y5/UaaGdb33WO5FAA0DFzLQ3
TmRqQS+SWFSlZYZbMZqtC4GFjsNSMepMhu8V9+7+iQ3zg71fpcMwS4AxzSAHnrcd
NjsxHkSFM1P6s5FY/O3fvb0UJN+UvZxSbADM9thtVm7sM2WkaafEWulbEIHDF6ya
iACYaw3BlbTUZYNTBoJay46gae2xH+5wHKGmNkToL60JcLGkIb0q269Xo+Gby8Ng
uQLGS/ACRazE7QLVt+RJ/X/PHXunPNqukEt3DQ1x36S2G7AgdWmMgjgDAPAK5KuS
PLTOPoxNkD96lUMv19Ermkd+K4H48O01o0NdWJcWeP8L6I/gj+jIiQ4R1iL4DUXa
la6cQ26TACT1bhQpZ2aKE/Ac8I1koJFLiFOH1s4tKXOXMDcgdSLztj5ncObTOx8N
qMV00hDjJvn87YnDJTbNsZ9GKlgoaDMmjEG8L/n1X4MrjgzZWzLEIqx6jkK0uhiU
K+O3k+HBZx3mQlsBTNMpxmzLBecuyTpfECMyMDJMSy5YpQ1YqFxqRh7605UhrUHW
g1P6PWV7A7YlCe9/NaXiQ9Mq6v6Yb/HNqe6HZgT64lShu02PWILRrJFKHpwgqX8p
VfqTzzW0btt9EHFZA1WzeIOW1lU3BCDXeDjC9CjKVcSiBqNu4vafoVivV/wxzO8a
idMXZOyTqOAuwcxHjXGyZlChM81bJqAn6rWyZ8xD3KUMzAm13Pal3sIzJBVpvQIl
8xUp1Xa6RpcdsZ05YBp25dnZYSBiO6Cb+hVB7Nlv89tznC5uoF0InyU8jrvlDPIr
3TO4qdNGew7K11NVmWuTfrTgR9fQBZn9uYuS1xRAuaNbLV+HVazsSi3zI2A2xQhN
sKtbFApX95rkShsKKawDxOIqARNrbDAXhxUd2C57K7EV83LYR9uAPCNbc6DnWsvF
bb767a06Zl2damyXqd/eyajeMfKYm4gM2nQXkwDU5OO2yoavT4WKnC10kDzPREt3
q015w15pKTStW9dkb7xiFyBEThsyLDhMuIK/d46BXQ46XODBjlUGskAY2gP8dzPi
KzLy4l30BsOBcJsbpuQhlcAicQoeRuCKodnwKthlf1bXg3Kr9jIAmtuH01uq+XBT
lkcteJ8HVelI7c7Zww7di7jxqz53xmKm5PRtW4KBiUb66i0LovBQYWkfPN+XEJAz
Py84M8RT9Co0daIh4tj0aofwLzMFlBX3QmYNeLAmlG1R40zEvf+xxJ11E/hy0XJo
2Jl/WzOub29iKzT4BC1K0onoGv9NHbK8xb+BYxYVMgtG3M5rnkvqYYs/hn8mu8NK
G+1sWyJu4d3H1be4oKBGHfD749ThOqJTfTROz5hoa+BwCn2MMXLl5yUfcU/e6o+/
ftvl4OgI4/LiWgR078YMSIeLpweHdIkcI35u7E/pgNHeYuOuCHQ0pSG0o4mJbOFe
l7C8izvqkSX6TAooRtj5GxtwD5Zv+VxJtYkkAY6/Uto7hXoJidx+Dms/0oIIlNJs
TrPupxfmp3zN+Cl4DXfVrHVO2tz8S/g7qd88m4C/id28za6+btdEWY9ykkrSnB8m
c2Y0AfdnfFk5zP1oL80BOjgPXDa5sJcMDb8W9cgJHiFi/8CoWOWJ9p49cn8Vy5Ev
yn0tN/kGYxFE5a1QQ6/wSUDUK1G5zh/mBYCBXGHFimsg1Ot06fh484TP7g1Ul9Xp
w+q9qyXXaEhTMH9djwdCl+7XjK0mnxn2KZRCJDaH3US9fzs8nnClv/0GJoG2Zecs
NrLA9gTTXg0vKj02R1ekHWSFfHkQaUXnIPpW27spopgCHpIPyWV8FGb1Od4930G8
ZS0bfdNNA77ITDibTA90NWh86ko7i/Q7hZok8Ih7gJsSAP9xL7P92kNnGu3ookcm
uEmCHuPi2AC6WE+DqIILMvB/gZx6Z3UYyvTDR1kHC0e2zeK9kfXMzWgMTZC6dWRK
8cPVTK6tMw+ZsWCV62/uSOZd1TM3lnKS3oGzuffYoBkmip4/GCxP77OUdoAPvklz
vYfgBikbCEeMeiayBTuK0ygCoLIyU8wKClBl/BpBp0XcWsX9V6I3Z6JsSt5wnWsH
nZ5ULOtNjgv5t8xzGIE6Q+qlgQAtozB/udPtSTkZ3f0JXnfWwlhXgvAJiwvlJVwt
QjQOx75TfVFROHrY5/EJPy9Drzgky/GmXy5zbG3yX3OMg10zm6TSfQL/cyJCzHVQ
7HmnWM9xL+JWs23LPjylUdl5tgz9u3tSuocrJYGqwv36mXcPJ1wLLPB3eaIglUyl
6jgHcY05HwqCqY6LeQsXP7jKl6LZtPZoi69y6oUI5uo=
`protect END_PROTECTED
