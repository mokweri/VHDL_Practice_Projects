`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+o9ikohVd7Jby49d7J0q/aZXdRxlXBL7RlK/bzAONXG7eInci7UZBncBsU531ky
xEotSXxSauDZ10nlgXyzczuCVWLrhsya2T2vMCCjAL0I9YraoNPnYVOLWeRm36Hl
puhrqBWucoa5rzEHK6v42snq5sUn1lSxEVNlwd2gtdgt2GbIP9DfzW0xUC+MRxy+
NaDVQejcuR9Ygfjhi8vCkjYXQ8TtV158kkRdFmHGWrSfIEfnbsERlECKBfSSUx2Z
vT+/fp9GIwkc928TScaDANPxefbbpark/G21A7Lh63T5MZEyG3VEosnSRP26Ajol
Ry7chzugLTelu2I2qgka4AHjNRWzKZzlhn2oiKHKHphJ6+kvgmkNTuQ7j4ttgLie
VcE+2hbiJxAc/yLIg9y1tQQ2YV4K9yHQr92zWGW8MoLjDQobXEDIJpcaVZG3XsnC
IJTCkL4bxTfU8iBgDXEE4OTef/gp+dbwstnEW30Dt5zbkFpe5amzAOh6ACRLLPQ6
PRZKdfIOaZLYZB/p7jLDt9fhagBB7FMJGvkjAndgZHjqWUUhMfe0avHJagJmTIn4
mWTTtVR5CFwRgCpNQslshv1Bv5SDZh4RjbA1oBgToBHqpRyOY4BNkA4l00iQi4ht
rBqPJcGkVQK/IOP8aMb6gJ2dIzOLw3fnRfglmYMb0TRsQgPiP+4EsszRpFwkJ+xu
QARcu165vNkAQUJH2iWOApu7FC2Jj0T1sKoZYnDGcKU4gbIJ+2owa5EukKm6ws7F
PXqfIsUBb/1vDqg44ZytjpWvwY4lEvAQHlbks4pQLnqyw436We70HGILm0YxeChL
HSu3O+VA4+1A5CDtyFQ/k+BvpjVfWZv/pCeAgkVdMzyZbnVZCTd5mD8LlrjiFWN+
6JRRPDISzp6yilXx2Mt48uJykAvi46TLUGFh4BRIhDtoGVJ8zEKNeDQPOUf3rhPj
/PkIc9/wIn9x2gyylqRrjG8SV/agfu2tZuqArNNCUP5y0/gbVC6hFTxYjrjgwztb
sM6EAP4YD0Z/1PMLh5Ys+LEyLU3hRTNyzZLYdymYpzbCGYiTexrd935rz4at47cL
2+e+pu4oMzDwyp7iN7AgtmBkJqrzCyAE8BT3MGbQGwx99BIzx+fCRC4hQBbPDRqF
7wof9YS4fZRiw0HmQBLVmod1ctnRqzCl6WtZ7h0mx6vjbb19BxZslcJZnTnL13vK
Fwc4KANVLeafsr4gps7Yxw==
`protect END_PROTECTED
