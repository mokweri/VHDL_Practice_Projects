`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OMZiiy4AUzKN7OmHK1cHyFOUEDjQZ/dN0Cx5prx34CsHhqJqojP0K9GcDQh+3MEX
37wABE33ZuMsTrj0mjOiNYM+YUXVARCvsCSqKfWPNrCGdgLpnu2RAIXbkqRw6gTH
iOeevcVQ+tXIihCfN2p3cNt2QPK6pBmOmqZJgvFTMb4FWmi1tAKrR4Rg6F4TOvJW
7J2N4G6aIxwtqWwT/jgMjnKwu3mpZCx9bzasbMUyfktX9cfxnOeqUW1zCq5UpUxP
pbJSTdKsuYoy4/8BjFz+NfljBJzTYrHKu6xCnOvf5M2S+TQu8idWjE0IhWiLzMZC
bCD7iMW9M3qgtG6/RJozkkec6nsAL9F1WIU6683Ii4++sxMsbVG1bmJR0zI7+Zf7
gkA8axillH4qT0/RLtGElrFcHhgxIG/8bLRcyAeIXF06Bo9K5610y5qvP8SDZrUC
7cokT29EseUy7ooLN7GyCvdECOHunHK5eEt9mocZPoswzsxOdbBT/r0BJ7MUD4m3
lFtekmSSsYstfBDSI9x4fQ==
`protect END_PROTECTED
