`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AfR9BnLA2jX4EerGINmtbSSyXZzUa6AX5X2AG2Lc2zSXRcDlxFlA3hKXJ1hUJ5AJ
/vc62cJHYxKnpfimEbuPhY07fuUwfLF1XVGvXHkmGWsPn0Rmc5l0QStLCwrdcZjK
wVlB7PRBtidPy/dVmtpi29N8WqcG3DcqhF9T+DQ264bp9gvARo7LAI7FgcXlyS55
Epk3qN2c//5ilv/MVJBrgaQWNCWmQVHPWNCIC8kyxwtrXAuuClQlKjxICTP2MgDv
bFerqhz44HSmBCXaZm5CCQdqaozVWiz1RTNc8iInB36uXXfpJxN2ILLkOZ5OgOsQ
VsxOslILrVD1q4mdR4q36gbWIoUp0DooQtADHItPnb6TOCEWz/M8xuV8sNJBrIqK
8vJd/H/E1nvuw7UY75WmSioAXwkPDcfLnWhcBjVwCgEDfWP5AxnSRfLEolc2nM1H
fbqvmloJkGPUdDyNFvl8QU7y3wtuOBNtnujSIbao4wA=
`protect END_PROTECTED
