`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hv5OnvZFFBKAne7WFpdbaYh/veinhj9On6Ol9ZdxeCu7Eaw86IGnoWfRtwE2kHl6
97+C1UsGqneXaOq+1j+LRudkvT1+yWN3KZj8p+W1naShlGsNsd5NUDX2uTFAwQU3
K0LfruQh4uCDqPSqoToIVe0USdl9ebT5zKtowX8ZkuDi1AYJ0Kxr2c3b/P43qJfR
BoTgzvF12uB72ZLEi1gei8eTPQma8u5rORqNxSx7rtzTHYDad7Icg8TPsW8psWc1
94GERtqDXNMpGYJCT0lxcRJkTweTYSlNIjNZM3vbwJZYt86e8zQKx1hsN6YHfQpc
c28MI5NW6mySshM01ms1ateX1RyTQYXnF0Q+O0RifrsPlAjkcSyA4rf1hi0i0onK
+6kCFgCDVLbaNMJ1CKHiJzkrbpHP4aqzQcPFTQIdTHcvPERv571wOz1ktLVeP6oG
fkyjbdTGEUVj+DtUxAdxI7FF+Bv2+qnpv8UcZRFKxsDoN/AajcRFbgdsBiQnkPAI
2sCZNK53CdlzBsQvND3LLGRZYq649UPPC/sSxJjJgHAkaJJm31TjFa6wFUXx6eOp
kcwUoSMJRQXFb/opVwTWNBmwuogV5ERkbRfR8iRm+BZ1i+X6YT3K9hz7XDBqbuyQ
KIQOXuZnvyF+jk8fGr4J+PntKBaL9VSPL1DzppBVrHS+H3MdyqdyQXRJpFU1z74Y
+9mlZdYf58Bz7wme2q0oSqT4zs2TP6RCsbXllZkNnPW68YuvZsrajzVUaQv6jnwG
OS+FLpH/tknXN40SM2CejOeVSxwGsYJFhjG8ZM2DW8tfxZuNfs4k0/56JLjdZNOp
KwwQFRBGm80iXb78r8YF+eT6h/ERHq9D2YkmN2Q1PFIWELyKlSqiWhFU9/qFeh6m
1ldmWYosQ7pNzzyzaU9/aGmKWmslBtn9z76ZVCTatvdETPpVzkoOY4zUNBtEWBfy
smOnQlt/wtONHS7VZryIcGEjXkUFh27Xj8aKjJFavtE6CTtlNRiEu8n5j/j5falI
QysjgSLKF0n1coR9pimuORdzMZE7+c+EAfoZVl/NnAn5iReqfuMXcbpa0SQ3T8vt
jdQoZVZZxeEnqGUi/dPpv+avxHNJDxeJdTHvfmv78igEs5DW9hqV3DuVevivmqoE
WhVKZadOe4ZPXl9h+5+09BDjVMDTASqR0OcHzhJHum+9xCujhEAVeCEsVQxpjtNO
`protect END_PROTECTED
