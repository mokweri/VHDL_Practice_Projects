`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oIwiMb0EDJGGbfbbRKWSedVuseZSndM70xoPTfXfI+ApiN2QShy+kBJcIXMmtvBa
bPvF5pE217wxjO61iY8EbgJkfGxBX5MU1BOQfShj3yfoE7fLpZpZ7OPswFVwQ+ZN
Rnd433AC8fJVVosViAuBR/XaS5bbYq8ZrnGCLAbGkmrQW5xr5zMg+JQn8o1M7Kq4
`protect END_PROTECTED
