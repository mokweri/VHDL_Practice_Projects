`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAWJpbxdnDsQrrhCwOlCiIUTQ0+WJ0nk8PJmvSJLuWksLG7OufMuDhiHnD5P94Ci
GehSyul3LlaQ3u3udENYXzFmd23iFOKi62ibRPvjPlKI8l3o5/YDB656VPhrQ4w2
/TxMKobvEaSWD31Eqhly5k6cCnvEx56yVY1UYNufNoqcndTPxifmbiuS6jLxWsOQ
Rxrf1P5Yf0mE2WIeTJ1DThhZZGIuq/YKIn+Lkvy+IZO56uqx6V52xpcWQnMQ9DO1
EFuwwi3rlreosCuuhU2Zve5EgPxmYKWxVChj+RTXGzwTLLh8DJIJIP6cqE8rY5mO
AecTmY64oJR8gaaxSoQ0adn6C1B3bikxBDoLMbqrFX0ddrNW+uoZGuOCpTi9VHV1
EiVSfwxlCPbB/7fLv95Xa/F/22GSixK+F/7H+vT0PBaSPblXNXQqpybfMLlFJJHX
3N28jFL0yCmUmEnc8qmb1p9iL1IRX0A+RD4F+8ZCr+T/tmQxW0zoaqGt6LKVs0Uy
9T6JdGaFYxdY+/BILH9NYUahf5j9bZi64vNdHIXiEkATAsyMTRvQDQbDAiSrhho1
ezkwd9xorWKpInJAhKp8Ezfmr5DhR+iR1VaXyBUeYnC4Wr/sFps9VpX92VVO3cjU
ghA7CwRt90QetLie83kXcOUwc8V1SxuJ/4xEJyE+Da02jNfnhxju8ohi2DLcGAui
M7Mj14hzoMFVw08y3r9a/iAR8gspxoCER18X9l7YDOAsq+Kw5iWtufmQr80FvKNv
ZzTEz7SVhl3zUf/9BQf8olZdcKJoPVqjv20xzhTzlz6ZWmjzM/r1C7Bt6RmRRl5i
BSPeJvr4nTA841Px0A0jvtiFSkO1gwDwHerytc8k2gupXCPdQNYdKsS9h6jjXob2
CbAX751yvSH9WseEOEEVY6RBJqAF9l7lYydJnyHAof4daLE+9gyTQuOwHttMOCk0
l9OylUR0ay9OxjwKWRRMMa2O4tdfFKWyR1j+ljXPzah13x6Ddg2GtCoDPJ+M+TTe
GkXIKYzMWFWR90RJogq/DDWxt42Lfa5Tapew0FQ42m3C2b4LvNPzstURbq3asC4C
BS1vaegzm/9qnL2mJDGzGNgMJYBci19G+qkUwaanGjMDqqqu5puEbAWdLSPA1DqG
fJQ+IZQNGh1yEryDGrurR7qPKerRjMc6lUCgATPiXJE3JRFxUksFOOfy/C7QZnnS
0FREz+5FHgw2q0hUmWATsPeAnSydHoAACM2yvg2ZDvfkXq3eQvOswJ1XlAVsXzLV
Uumdwnkk4KBYMyITMT2cQYpbEYiwLgRwPT+VRNSPl1GeN09b4j8pLTd4TDLRzCuG
fOd3PJ166FfrLR0eKeQR5ejFzEc9DiI9K6cvljSliMXqhm4HRwKn0Q/kPRxkmL99
p0WmQ031wXAETaut1VKgQqKtpdnhKri9MFhKnCd1mYaMBJB+/Mzy62bc5rtd0YU/
9sZI9BSRjlD1PToXuuh24Jfw9Xzg1aXdENVY37cgXLlG8UgqHe1Q2lAmsRvxC8yX
OOMG3sQxFAX7gK0ZBqyMiNBQYpGhUcZUaG5yHR5kvicJTj0Wfg2xul129+Ac/+kS
s+gVU6bATzazxfwsKMAzdasi1ETspdN9FKvqFOJh3qOT1dFHtQKz7drvN2J0wgRZ
b8sDUIEEl3ZdOT7XMcxYSrR34u9au++AIrj9dslKoPF5603j2CiOUz+6GHIi4WBp
Dzx3VkNyWqWjzYc4zQol2wA97gNFjnXX18wLarL6Is2dOM86JOlJIbYnBUKl9s5G
PzPxpZrCCx9Wh4tzNbRn62f9wQCT/DnVDYDIzvyMNejHHqq+34Ak05b5gE43a+11
twZkdupiIx4BziVonyIcFeJ1ZnfwQMOmZAKan3lTfKDyvMiMwYKzxTlyOYDBCnUv
e6xkUpG3PlP6umZ1ahd3kfRBaE12hJSbWLvJzSO/NJKvVpERm05CKYt9XujDcNr2
Gv0Z8w+lqh1DbSSmdYsXxwngt2z5tBA5gwTGEG3Ag04QGilP3BblHCbYWnthyupy
1TZ0m6mlOfHEOwVoLHXe2H4E5iINMjh8/jUgUElMWXSDFPW09+eo4z/2PATK/swC
rMujb00IqnbGaLBbgp0gsWvPbooxpOEvP/NHYzpweXhxHn2lnKjcJVaaz2MD7dTy
fORpStrjYjfy8/NerJ5vjsoMhAlO+SzbB45khWb7ccud2za5eIJTlLJoJcLe2Qes
uFwYgQFpsNcohJVeZQERUMaw6nugEaAgmd6PGXhOHnM=
`protect END_PROTECTED
