`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcydBqnSxXmB9VF6DUa0UsfbdECJxZgNxcxfeq3Ulwrktp29S6nmxQzyWlN2g6NR
BVqKnSnAHlZgA5gCkyNvE4jfctgtl4afqgYAhZ4apfvOEQ8oTcZqflZ/Rycwbig9
slXHak8P6pRYlr6UNoIyzq48OBS3ncS6dWovqcPvr1Ie4LLbH2fhLJ3aOt87e+xI
VhtUot1yZBIO3o2HBSyeWP8/RHRJALvoG4l/yzkj/3liFo5ZQtNG7cV/YDiWYfrh
hUxGlo8ZQGdNQJv83UvxTPT1fbtxeh0WFJ13zTTyi6cZ221UIrUgCZr9z9f9SxjO
lW9JGm8V0lj3A28Fiax8iQ==
`protect END_PROTECTED
