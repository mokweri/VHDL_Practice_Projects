`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rp4+UD6kDUU5Skrg3Qa1gfcaj+nrLtOXM9/P1BXNTis8TxZXeVmsM73jE8k1q8Zb
1TQIqPXVp2ob5ReWGP9MNmGT3ZZTVzM7sF1YiEOoc3sohEuThtKwfHkyLBgSraxL
oDlg85yFauRwTryaQv8x0tVaTsRxYvXAjtiM7lNcbrq6yPTLelQzsac7QOHS7JeB
GamtXlSFx0CIEPbfnicJaPdQIw+XwXMX4yyhTRJHq9UTlFqk+3drbwzsoEmeq3OH
YzKMSeGsi/0h0vLCOJ+XYc4Vvs0cnOze8LeGP4xuGSH3Px2H4ETrnjb6T6y7Pysf
ARGEtdJJyzRmNIQ215ZChK3QxxRBRq7Kxhg9bpFOCAtIwyTWj2/cQxz552vwdkcB
01VwSKD7DS7YtRyOxB1qjNyLqjCJsVdM3SQhDqEgDCXQJffqNBL77cmRAGNv5Pfj
li8cEae3BhdHdY1p/trB5lApyiodxS0eDdGWBzbLRbev111maYS0lKujGHS3NjlI
xcxAnpI+tB2oZ+abrfxELLMhQRFZiAClFZQaA74/ZVBXOybRUgS7cmKua9O+QvWO
UEsU2Hsy9nNVRF1PoSp/2PY7MZMhGSeyDCaUinl1Q6E0xZWywxBarWtow7TTRQ2B
CUa7ePJGDZJhnkyEKeJGMrvJzO1ICMiPGMwYLXRAq9AjvtLQvxlvTlOOKkRIBaAA
HMnAz6M4Se0QufvjjgoJqEV0+GA1Q5kAToQwKRdwSPqpKI4aw61U40SfUYOHlUSu
Iy3FSDvMVDOGG3qNg0eefxPETBzRqZLdeXyLuvBTO9WG8hWuNJuRufgKVyq0l8c8
Z8dKFu/mRCBcC8g0Ok80360IxZsSB1aVqTmpYiu1d53Q6j6uj5UboEThROoxNssu
3j0BMV09Rk9kbJXrLNevlaWBu1wTCqQy820wn9Nexw8ZlmHSkol9+9jMIqeB22o3
fInhs0McEbW+MKg7AJfwn0zya3kpZU2yKXaeHT0ItqbArVGcCX5c8cxdlHzLtaOY
yeT4EfKKC11L6TOHw9AkA+OzDqePGTDHXPljB3hhyIZUP93qP8FLjUlGWPanb+lT
zzxUjUX3L41xDLrZeju+U5J9S0AJrlvi/auQtrM35zEle7nrLnu6xG6yPs/Gozfc
9PvqDfml5FeF7T3ZJdk6uiWY3p0800DnBFbe0qEGigYn3s/4ZRIZ4H2VSyjZHiDm
OA2dpzFfhV4B9jlBhor8nPBnOsVBmoROip8jKzP86AaBPgq1dxvbv6h68DaHIpdx
`protect END_PROTECTED
