`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3NYFVp0kVEaQHI0Rt8xiL3iJlfXxoXk7ad6NuGZcWaeqNWy0mlOvD5ET0opI0iA
fJYKDNAYHs99IIWAo/M7O4dfZ4BOjEyr2fmZtAwN7KnhznL/eU3Wp1lt30q0Zj1C
3/YIDfQ9IyJoc1o7WJkq44Cfg8MBzlg77NwbvEH98jzJ21J9PtcUbXXFhzoJRsWc
xuUuYT33F/4IXowXKzejrqpauD/cSpkS4xjTObC8hXYDL1VTdlTJkWuILLqCE6tX
h7AI/3NbtyDIBKxMiqSNCIX/Z6017qGe+PwgEtOyBhRVmdxEuXf+RrhQvxQAlEGW
YtlbWJQG35v02vjzTv1bJw75okpgg5qX1ludL/lCsMhfHFvMmAmsdyxvxTE+6zBS
UHPrRLcnDiC3tiNgWcGsDsQKfXh2o+hQTG0KNB+DxkJM4vjD/zxfHk3TI/VZimTe
kJwqpCiRiIGZdiFqyXctYv7eFa4np69hoDCzGqPwyODhVQS60bGE7APYbB00ZK1K
F4gCRymlPw3xOV2y63lR5MVOvEBhSbv3VZdRhz67RhqsPWXBwgqdTmdojQckVpq+
iUubUQ1CSnK2PattEYUpuq1vdNW7ETI2gNaPZUun4vA04PfkOo9edQOSOGeL/5F8
RNWhh+LUXs5x+IjGyhLhKto1wJT1eQjqnElOdvb5eor6A4kvRbF4yCzJQwTz35gr
/+W5KxWxg94CXDu5rbmryB109LcooCDSkGFRl5eSHb+FMhwJ39Tq6e0ALvAwRJiH
yMKRHFrdapKfz34Uj1O12b7/pC9RjWIF4LxLjoRv4jV+bLxuMnGQrLNV8e4a/29B
wQ4zToqSc6KVGQLXvoeOz97hmwPPxrw3dpNsniYvC4Ek0hrAUuT+jEjxGtYItk/w
UUjN61LeQGJ1EEY/uHp8F6E6C6isW/ol83apaJykSESlBxYJyiBewnw6YCXu+Kqa
7lYoehj5KaZc3RpgCI/LBtZ73SLoOhbMJiDHj3JEAcR+PovJJao4/VLW6N8UQ12G
ggixGJT4In8UAaHdTKRO/Yq1T0J/XWt3DPKaATCtK/Ru4GBk0Xtlo4BoO902dPSy
6QQK3o34FQyZ1gjK0pNUisEs64obEvHXSJ/rDIVXfUdWp6XTrvP6UwYDBrFQyS1j
WIGW1cEchGS0UBjJZHOIRcl/KqmyrRuYdQHXBMVgONQt4KfyUV+ynVJtWg8tcp3c
mW5+6jRwFf9qYkIcpCyi5c8svUcLJNlZdb9tRwQIXXf1zlzg3HC14nQDMbuNK+wK
UInSGo8oCadciqDKwSbk8YwRtzFOVGKLVwuUceIQRfCQQRHJQDwLPkgoynzsByHC
LCIzm3fsNbR9AqCOT32xOeD419pJRiiF/k/Ysy8T3tTcDQM6xipFPy6lHhkfa+9g
tbNKm1pvahByvqorRSIO0eiZ5xma2h5GMHZo0ha13JnsVR6/GJMrJLqzMIiAGuTm
3QWnqXUx+ddBYfCBMrMLVQUwTvhzKJvBdp/MeDEmyhBE0MMIS8dS1WLgviHIMLj2
w2qhf+pJZ0wKJKY1KEpkZAkq8b1Hp3MlTTMtkX1jFT7tX19CpdH0Gihf2OFJmR4+
j4MgwOSO3R8lC2u+uBiB25dwX4mdD3ZFdnzecn4LxgxATa/d9Llz9TuJFRFkRWX/
3MOn1RreykwezHF/deNYZ5kWu/icahLx2G1PA2NmmHb2nubpgJjH3RHL06RGbTuR
QI8/Hh1ffyfkULmVfcLkV/teJYUyRL2v3ik6MNqr8KjWe5F07ZPIZKD23svvaeTI
24T+b1HRGhFz6pVmn2tYqsBvl3Z/YE36uCFgCasJn8vP75o7znTKmiVfS1JbZCjD
kyzD3ZSwH8Jtg6Vt5VvSdAIwxfZtYk64jTQIDCIhq4ewYx1u931Onh/IpFmeqM07
lNVF3Zzz/3i9j6pfdVgliKIL2uy9MmZDf/I02EGhGuO7VUad/wo+VgONh20Xjf1y
QH3BTDYSUK8zbLAfhxut/Ld5EABVjRMWEqugce1R40hwUpDRX8rb52E7zebEp+7Z
GvErf2C5CwQMmiIJDrPbW6FQw0v1wome11DQGJ4VP/JJwJpD9QOAi7SF/gssGV08
lrjCqsS8rWqeWD6Jg2NPdE7BhDSma4b5kkdwUobtjrEg7ZYQcET0f5ahtTQgtAEO
Jed3rG1nHOHi81rRNT0y0DUg6aGyyE6KKx6scddL8/N986m9XetPw10wjY/1v990
qsBkrmCoyT5ephN+BkE/tybgQJiAk16iQASymwyubPFBjgfJJteC6/NCP6zLFC2v
8O7//IqzQn23t0MHQ4fCo/XHfH38ijZ+eni3Rdw6LhHefpHeCWH8MydmY5CZEc4k
zAhyKdLj+a6j/1kyJ4kBb2ozXEbZ+iBU3lbSJ6hwDnrTt6Gfdij+Icdeh6Or+owd
CVyoiEKnAk8lNCvcykVnr880aUtMV0d0upzXTb4WJlkFgcbBagoDwpExSMgM29kf
3Ii8KKnPycJoGv4L7f+4PPJCdtZTX8naWPCy89qsa5oHuvu9MX9fmB+qAaUd5ci1
Zbl+i8Z1d+2w/BEfnAo3brefS8d9UO6g9va0lKIzUoM1L6MVbZfBV2ysfS82keEu
85s9FX0aeRmgyRYQNt7WkzlwHhNfNWAmvu6Vi303/cUsOrnEcGI+VAtJhMC5JqIe
ht3dj8wdKM7UhKPCrjo+9eN7ez/0qHi6Mva0e6Ewt2FhDYqyC3cnuCQBIZlmWMkx
mJCDTjp4bphkz/fRSx2V8sDe2/+rMgZfbwJCMRLa4h5rqCKSvKcxyIzj45qypinE
VHDUP3uSLt9aAfImZ2DcJoNixyzHdPRAUSuihbFY8+ifjOIiwVjjgf2pGKX0nwnf
I0HgzxkeQV4IsYDJDDcdaZi3TGNgebAXWJ/kaDAK1O9Onai02eNp5DhI9mTJAcjm
LfEQ2LYVpImxppEZKIWNfHfniEMNWuB11b5ZIONJTxDWEaYV9U8vNO/xzqgBjv2z
gLVR6FW3/56gw8K9RwCTysSnUcTSLs78ltIspdhULr/ztnXH6IRfIH5eSC6fuKUT
M+ziMokH0/XNe21LmY9/N37ZKboz4kojPeGUG7ScpR15sbgpd/rtbg08GnW15CWu
GOAGaQmg6v6l5lJJGchRp7UZ2sn7HAUNBZ1DAtD8LAKtSI9IPyAeDcqS0nwGoIHH
TDUH/kiCRUjcpykIFgBdsNV8sd+tho7QmW8vAJqp09S/zpZ02tm2JTMUTINCIx7q
cEMFntHXE4sZ0jV58V1w7amfzxyn04LeD8TygfMwG+791EO2uwtw5z5WJvZcltdr
VrRaDAqM3cuapFbTX57Dr9sb4wmA3+4ZLDO7gpyvSe3BrtfR9o2I8ieyLG7B0qwB
QUivBi9UDPaZzcwV3IwCWvtlb3T0cI3Ov/YKSRotnFT3eacrq+OOoqm7BybpA3Wh
3ZPU1xFaQZ59ixUwOJw4Ozyhmbt/7pNIWhZ3RowPQTU+R0HN8YvLVw/tYZfQrZnx
0MRCQ4rWx7WNktbFnAYVrybsSnti1js6KJskHjWrVwEOkQMQQU0xBjrYNulNrhNj
C1tfPqgH3sky7qZkpU/nBmBE5f/sUFQhCxNZ8adCUhcdKsdCZdE5mrMfICjqBfuZ
9IgCKQQVnLqVFrlavC1J2KIfYqE+U2XURT75wwLg7Hk87dtFbcbjEs3lHiBbUm1i
rx5gJ0N2vXmtKoWcg+zL7clwZxjLfvDcgR6OvoY8kBqkiy8ACoQdCfAUVUZjTGtz
8/BejbXEMrNiXXwsr3kAPgBQ9pkUwSRtEcy7IA01Bit2x0OYQI3RQi64iwmjGOuO
2kcQ+6FAnJrdzAivIHJXRakVq38IsVbriLVPC17dU3Xg8FvxTtgvOngrhXz0gNHM
G7V5fMLRD8LFlBfYpt8gl0jvwgIicRXf+NdiuTTDKC+W37D4O1ANaeJ+GYFh23vV
aLdup+6q6kvHSHQnzfagImMdwl+jmdbL6kKO1TfukWRqMprT7rnchUQJ9xYTRyrl
qO7Ha1HuEmPVnxSiqUxurb5CnVqpE8fRUgvzXocrXVMs152BgRuk8jep8J92n7VS
OBrsBSXOBk5ayYYBamKaR5mEtYZVs4ExZ/6gobLZxOVEprWp/U1z7CII2TO4bgQ2
xGPKakIXrvZQ3hxBtlg1hILDZzR7P8mUbMHyMfYvEMHqxovZaOYgxqHVSe6MdGHE
wnzFPV13gk4ByzEvbyf6vq80JeR6wa3QZqaDf6HPFOui0U5kLdjFb0HPbfRkskEG
JylFyR2wAvevFss+OBzeuNDSYXQT2X+t0jwGPbUvuaxU/8H3xBznbHLQVPQn4MQt
SSNUFyZevtogDqUGtf+ikYXwas2vge4HTExr/H+g6sWBLc+iAdOtkiZ4MJwqa2sQ
vOZuM3Oe+qmj91MnsvMMcNbWAP+CCb2gJzUyflqW2/2W0CB1iWqQ01KKl/4noEo+
BfKWGgy0nkWCGF1EXOzLz9XKyjcCUdlwDtXvEzdjGivIWy4laBb4RDrDvHiuNsyw
R2MotT0lSDk5aPGsaYi+ffOTWsnVt3d8gpyAwe+UA89ZE0KRtnAqiMjqO05IyO0V
ZV78wXiWxH0P63Osy/Jc0v2tSgDXh/xEi9K/B8Y9iDgMdNvV1R58lDB2kNNViJfY
Lj8ejRRY5+cH6/gK+IqoLJ4ZFNNhUEkfbyo9nZQRzeKPwhwLIwtuVCCxpOTNEvTT
wo7EGJOFZRidplPMqP6qnJ0pFYxZNOMMuywTGz3s3hUlXjBye7xoqhBuJTio4vvg
6V/xvzn0rsmJjNpJ8cq7tLn6KVvcQWPEdbX5kZI3OwyouxhtZTp9Jj1QTQmwtdC4
JIEcJ/aCQlU9Z7QY0Q2jxbH7uRx1+XJbqzl/jEnUxPOj/zcurc/dHUuXrOBANfBx
Ssh9IppSrHJXfvBlZy/UnJG87x3KcCTrt9a+/pKN3WWqW5+rAqElBwgixqGw0XiP
hVDvX8X9IovCJMyVGXBHKY59apYIXkKG4J8mEIlLPo5wtanRY0hNlECQ/gcrfYmj
SBMS8IcECkIz1qc7AEHPKbW53L60HHaNZNWJrcZH/PFSc+Wq2FsZqsSEfV8QAJQ3
DbVHjtzibtw/SUUmzvi8Mxv6EZfnmOpTcaQUc49yvL7HggHwTvL1rHfuJGJLL9R9
HHLJzlCMZ7gwRfzPl603uhqjZox1mR5qLmCA3IN75qVhJYBfGIJ9LvlNZ122sr8G
KAMfF0KOSR4r8lor4fJgsUi3XeMdNDJm/mex17lCsnoPrN0pj0zLzXwlrXEcOZJ1
56OGClnccwmBn8PdYCoj9h2oZrkJXzj/daisAMYrXYi9KwvZ79gjxKu3OJlGAAIZ
CW1k4U1JaQMiAWVm/n1N2Tbd/0jg6oVkEdD2Hez/TJOdbFSzB12kpOKyz6s7Y/st
Q+76jlWPQUg8gTkuZee5lYE7xq1Rkwz1wVGGU5BZwqA/j6IFSblYt+d3Cc8uorhj
2FHZGjKyG4bxBhjMXFuMeYqhA7HCJYGZU1TImXv9/O+Onn6GmQ0WYtvd2OAIOAaZ
pPjHdZEc6m8xBgY7g50Cy6bUOw+j93MolVqcDOJoRR/nTtVC1pJ8WU9ahqIhQOl0
uuSI/aSfurZ5YgHCxF7bUmrfe24juDoiQyYgywBZVZLaQB8KqZYa0GAeVnHJv19W
yb2j2YoYG2jJMfOpbhs95JN+cXBNjjFlVBnGSq9BqAz2RVhuD2O79vzmLEl7Twz1
W2hjr/4WerdhusCsNfMtxaVrRzZoXinwKPmzQvNBUqL9sb40fF4Sm2V8gRONLCAM
rXNMi+fx84QGVRswhHa8WkSj5KAjrYw9sR3rIRWQ9k9eJlSy8LeBN5b9/XMsvRC2
sv04Tb10jKaBEQHQaVa3B+2wq+GUOZFZnCAloC9gWqGaDgqgpQl3jkLVrGnaRgvV
CmfusnPJ1nUDIMgPz6/lpLEkiwxflF5n2rKKzrno57wJ+7ZwHokoO1QFsN3/dAeb
LkhsCD7A5eXJUIo4TUTG3ptPobJMwnq9Eps8gb9/fE6hHXpRKrBgSD7hs3xjxOGQ
0FqKKSB+IkpWtmAN0oDGavtfjzPQqU6RDgxQmZMGJPjYL+glBonsCmjRmPwg8rHH
N8ul6pCDrpPl6VOTT5iTj93RAUW3zgzf0lxE0BxxG4swaumgWQRnPP9ohnFmmMqS
STif1qIKCb29SUrmFNOMIw5DLqd6jxrx03q/X6u+OWNB2K9Iw80v+vV8AQIB72dL
gcTmULiBOMs2M46+z+9tHUj8cF7pYChEe37gkuLAgTndBFQqyYJwD1C+OSrKkoUb
2Ro393uxtsk0i1+z8reo2Sg4uinKXw9yKM75KD8ubxa+mGEmde9aXTYwKZJlFkiy
5IghPG2U6k2bPxPOX0F2xLGX3c0Sc5S7Oclj4XGJ0rXvLGnSTDbLUQ+pWb0Jm9rl
8EfEDH2GIjiwisDrhU0e3VvfMT8Sq4AN9NcHtwhqDZi8rdft/HSBX2W1vpflSoQ1
nfvGMQqSXes3o0XpgwYbBxKfh/cjRSjMf7ZOoWuTQRV3S62/vUHSri/FJ6j22xKe
vTgPnU2TkBrfcbrH0UORA0Omzj9PJYXfM7RG+btzfRIksQJmvQVn9+In2TI96dj8
eIx74RBtDaTJmmwDi+yc0XjKeCwRlIzUlqyWy3yW27oYiqqa4/cfQa/aSRgJF8Nh
zzO3JzS/2RAkr40qmcLPgJbpPexdt4xMvCRSsmy9uIFUmPrBiF8uJ/QTc370VA3r
oPndQDD8BYffTxxzz1w5/39+xFa7ZrSIB6r0xg1Mp2KIVnRjBMlhweB+Wzha2SGP
zOUThag7brUUDyjDxgg58m1u0Fu8/DEGAoWkCUP6BxSZZDuaTpft0y6dsbA/LrSl
5xOCoGkQzU4E6uh1qQkSO9Jc1SUYmx8QYhatxF0l5x9+fIhy0T3mhHVfo4PFa86+
DfF9JKNHmkZhVUjiVDDLRG6dqF6j1DGqha4vDx+MJd9cOUocdPAOJxnTBxhKMdUd
XafkuLmrRniozsm1aIsSwOAJwtjCCQ1vUdvL59SFCz+pM7CYnNQnSjJSQUsgKfMK
XbMtShfz5ifJVhgNxrglIeADZLuzUd14K6vUYceRjtyG2B6ovzeUmRKeBO6+HwaN
7Kpud1VSPS8HoQ63kWCcNir4ZvoDFRVhu+UDIoBIm/09E8SHqRIoZUVlx65n2axv
WRVDovHZJtcl5DOEiYG3M5EVR7VsJWJcuET/RsBwhG1f8DPtcVeG1MjId6xzH8uJ
GwnGP+SEHvjqlnlCb1b4gIwmUOtU2/W7uwhoXzq1oHhqu2fgUVuxQ7ecpz28zSlR
ttFqbyxmp0jMk5Okk6bSMAjAOCijZosDqMoJhcwZg2N25yETBMXFf+EzhuKN2UuJ
BABMCRfp3JaVTxQ1qaQoLGih0lrRL3gSgsqRptAeLwzB+I9pIItIkNMChRID/N1M
K5kjjn2TK5JTJpYFHUhdOCOS40hXwjuWhTlnHj47BjXPKmMTK76vbjsU2yhcXbEd
BGEYHbdwrA8qCGaYnzqJrsPePkvIumwyqxWUV4b6NFc/tAR6GIh3+9n3n32goX+M
2HOnCPn0QRhFl+L2G1ovBe8E0TsJzXcZgZD467/Y+SRpr0K2ZDy/4iRN2mcsDmcg
amyZO3ufOD/3PHelXY9X7UsH393mp/pfOwsUqioqz1OnoWaLwiFoAg0NS4+Gz13c
fS2+c1nL5Q6QJmHwSDcLmPO9tW7l10UqvCf6Qv6DswTfKNDET1fgr7r2v/yc3ZWI
62yU7Lsruk9a3dKToWEHA+pqmlyLtTW+lTDXmbdJ32+eptCyTHiflee+BF2J1T25
s37VzWg1TBJfTVNvFk1AIpySfUgpMgPvqnLQnqUCKiH9hqsw6uuIw31NNcru7mjC
NovFkfQMzuilyWE631ty6TTv0R44rwzbgHgFgNbU3WgQg+MypGBr0h/9Bdjv/INz
gz4fKQatgOCPEgYFaCPbyKb+Bj1lCgvABVUMdogP4qduXzWbn8eZzp2xM7eTensT
MqhgxW68kQrcfVc+jwNLRxQ2xfk/EiQK+u8mjb3VaoXSI7+6Sztt0FRaKmY+gYP0
jT09HxnpXhnz9/TrMfZG8Qf/TVZN+jtpJf4A+W1222tay8uM6Pa01ZxzE5Ky3YgD
NKuPhFnATFGXU2de97M/hfkHUH73RiThbaL4J7w/HSYzqtWAuewuXCUVha74yk3n
8bA4XqpgMxbX3FH3A75q9FBwhsKb2ltqZ+zEAvLryA9/6VVr+m5n+kUrQocW6Ha7
vQZlgXH/WXnZQ/f3LsqllzcGjYLXofVQTdpHsTTI9yQgcYanGFUg/HHkWEULiaKN
N6MxgG9w8zyftGXOauTyfgZi/MyLg7bYibX8lOuqk3woiPu+eUjp+IYWpo83HbzD
jgsGrsrmV6xvqw31Sc1XwkccN/mQCR6WW7Kma+F+q0n91nyeQkcmLkfWgqO6U2Md
CGlBw3jZJ+gYXirWj+H5zN0sGDdYnhcS6UEKDx/EMQcAI9YMuUZbCxfGEFTX8HlX
63VeAsYnaOgzVh7bYE+Gr9LNSZAVS4/E6OczTlkZ4P/3YlqI1AnHvoRVBOtfmxsd
y3khaMc5ilUnBbmkILOh6ekwzQOQQmPrrEab9AAobRsRdNKASK168YIE3CdH/NPC
w8x5CI8Y5s0+G6aY9Dc6vuLIc2NKVjp9wzv6fUoqzP992Edvt2QzEJuj53o5Gn4t
W62VilVCnQMhE87dbLgRj9zo1QuvExr6o9d9FfWZzMvws2ktb41FBGkDh9ruoWFl
sEIQw1ChTwuzgW9NCvcD3hZUbrTzTc8nIG6Rw4NN0/wtkM5LUj0C8PgzcUaVmm+f
swzVaeK4qab50TlfbNvGQ7hTC6Yo7+Tlqri3n3nKOfYxvCuM8uZLRz4BEUmRcjp8
02C1ESZtHS4PxPmGz6BadaCq/Y/HMrQbp+BGBtfpqPjcMZfvTzKA/k5MEg7HCs/a
3S5/eRYXd9vyNO4Qiw8SlN2o0X87bJjI+8MngIt38yU49X34XizJyiQcEHLPO8h0
+KvnTipr1pW5UeduI7vdMGEBzvtpo1XYCtDOeLym7u51wlu151sfyK8Nvb++Y5QI
srCyTiRoIM6pZ8Ecf3ACqZPtbEifLYrdMgJRVKOZJ2TsYykh8WCWD9yBrVdV8D63
Gc1aZE2l1UCD65hdPYL/2x5gZZ6QV1MxgTke6J8XipTCTEig8IurLCXdFLuMZaCj
8z8CimAHN9/Gc7j9T26XsyIEuB4TNhWsiitEzSMh6VOFCzyWrfDMVLEuQKt5SayH
fQE7bKW271d9YLVeZoRtdl3fJzClIQDzx3lua/DTrt5LVRJzfO0QdRrVT33D/7Rs
2Ua/53LRtJcRea+2mQdYK/dARvafqqFLdgCZQwWK64sCuqQN5ajbb6S3JLIxCqFB
grQelM1MGFB+ENy1NtyVTZElkSihg0XfGPnT1RDWjlT8LC03mbedLBWdztgFWVcl
oj81CRarfYlEiA4qqE9Hz78Ot/QXiEe1LMw6vxCs99vtMIkL7d3uZ0OBOXg6R2Jp
nuNDKIOJJpNSdwEWdmTLY8aWysRlpn/Kx/tsZVPmhJx2GhERWH0l5h8RymVM9Hgt
Fxi5AikRKbRf85k2nhajqcDKuDYtjONa6ZQiaxcQwLtR4NFdVhrfo2E9SpBQjQUy
lx2hEJLADcYyQvokEeK7/qnm/jgHver0nE2cvdEcz4My8xoL1rZK/06LjR0XtinN
nXMxQIIX2H7ahiUnlG+hhdTeF2J8wxgEnwHcV+KdrgedR34MdECE8b1Qc6q4Mpro
PnSouEwOKYFB32vDSOkqamr9iT5iurJ9KIbk7mPpXMzq0vWPZ+CHJgnosHni2qiw
iEiH72rHxK8nDJ1fmJHTzZXbEwaNjiEDT0iCUC3BzEQw7z9UIPOlZj8juvVPKCuq
SEPShRfTK5rdqwjmfqQ1jg2tij08rUkvLO2vFY93f46l8QbnKBi9AhMnYId7V6hG
Djjy5V4TMa3TI9sX983kd5pBPW393PvBNYkituELuy4y+8u5KE/jYYfHE6A/Sycp
ZNw1q3eYcAEmH1ZI0Y6gAnbcCQ6FNU2nEbY/ICMRhnBVHo2/KLTLIjB8vLLiD/zG
QNx6TXMJ4/R6dPETXfbqDCMEHHvY3AYqdq5ERz5KscjsbmILpHSQD+oYV1AFMWnO
pc4f1p46QuCslDjfABPbfWz/aybA96zg6m9FsazL303yMYmfypNAYwO881AwCc+9
HDsLFA/bjW+//1rsdnyxutwjZcAxJ+HTLGYTDK7sESc0U3TUi7gj6BVc8MUBdf2c
67rE2JCnbh/QQlVFW0Gg1z3ALRvxOzTb71VEsqPIzPbF6N4NTj171zd/IX9owv3d
pg6Cjl7btBohBAPyIoQa9WxphQp0Qnnsp+pDGEjeLfQiNLri1St/1AivJ65z+E2G
igAH6XyNmVtBYFw+sPsT9pOWl8wLcOEh2EGCs8MIJH1ATTIYWCfi4wUGcmQnK5JX
u2jY24RIZftWMo+ubw0Pfb3ziL1tz8zRIQx4QuJ0tJoWeXvf9N7qGwQZ3ZbXqN2C
uSItaSn1YGT4MGglGNNEocyYk4/0qq0yzOSbogoLtsfOsHZcT4VCVyka5I6iSxCW
HURvsWPGLFr2KI4eCHIz4jQtA6lUcJAEWCauE3wtYwi8JU0BcuVvFBdWBA4W4Suj
KbQ1omDRxDZtxhptnUNMyewcA3G7EUqGyGvchXcwaOPE7MPo5PMmgN+1wIq9Yx8n
Y/IKAdwq7SrH2IdRMyNcqrI8RFW3b5lJxX8fP/S8u279BnvZ2ptYqSb3ybwLBWB3
2YZu522l24Cxrg2jU6lSc4jxiiVjjVejtloChtuNFAsRTmH3SFq+CjMu2YhL28aB
f8qHmSdM8+KV1JjRBdt8xF3SXHzk4/cUkerjCTEW2XQak+HIcTL0dlrsjZG5k2y1
DcKccRfHERecIz4La/TnB/18dp2JLaPJGFALtZTzWih6liwodhkkwgp3/PLybz50
8ckq1yNHpUKwp8Q8oh4PRMoRXOVLOvmIqX5N9r9y7td9oUa3ANosnCNYBtck4ktf
iH69PCpt0odnUGOwf6YuEhYCwnBUuE4L5eNAguAm5PhnfH32tV9meYOcGIw/1BrE
AUrY1/d52Bnt4WzkfZAC5OErlsZrGD/AWElIi+gNeoyz9BWF91iZEJG67s4K8Tbq
HhBUvlLqYIhuU5xXb4thwEOmtJSgP4pyW1/zRXM7qeUPOlmW1KGSJCC6r5/Vjc23
datscjcrIK2kzvCX+OuYwvhvn5xEcQAZKQsJty8Lc2BiHnhrcYbMK9kAoZAC6YtV
Xp//QxHbvzFH9bw2DLJy73o4dR/sBhKmq37vKfi7dr9+1dtRf4w21xrYbMekf2o5
N9gXO+e0RqoFQ7Hgu/u3/NzMaPnm/BQU2htfdj7qwco6mxj7OWJx10qJEal1+5JM
27wEO36Vr32BCioJH8fNO8pYAQiIPKKVmLXlGTP8Sq9xFrQUxxovqZ6h7WkjhJkS
RVWLccMSjW7OEfFS2+4UFKasa4WmTjdxyU3d4xQmS34D22nrybyJg2QTenfrcsvz
XJ5r01w5c78a4WhQAfC+2RQiIFge9NGrSHk7lfeSRGGQSm6OQhjwBwbs9ZF18wlJ
2yFpGQ9k+EDWzZZw9Y2zYQ3zMV8hS+K3na+QydUMfA+hDbTPXzM/1jim6ui3BxQp
FFSp1VEGrhE3kvDDJntrsLqeqxRmiYoEIi25BBBLtT1A9pTh+RUiGWe7Kq2T5fQk
/WZW9lk4vBFN4duGxEjQ6vnqWPBaRzJK3aMr1Pra6fVQ/++szm1aAkqxWC2E5Q2o
8apb93HpnmoMS3NYGwnp/LfhgZp6Km01G0zdC7/qfl5YpR/4un/SthaksQPeNw6X
2hFhRcTDHpibkFEkHO7uTMDKybH9yg1YQ005Zp8dVi1rwWaTmjRMcl+caB0567/h
A/67SIvt3KSFfiGkExP4Hox5+2oxPXqosV2l9lOl2h88eBW9Iir6S5wqoT5zlRIy
0qO1fMBp98vS4rBpQgxNL0Wg+f6PTSbHFfYbszV1nceOX2dlHrhDWoN3PmQBYh+a
j+JDVCK3WeVfkl/K6z7NebjQzdiktQOlYT9B5ZWvHlHwVbm5ClJnN9ttbSj8iFsf
lxOamIzEdShcUV6LYnLrioMmmDXETZ5Grb1NQ/nAMzPnLvFJ4HeaJECte7fq3OxF
xeQmGFfeX/yzLwmVDImQCHND/wLiNHzYzRNKpxt5C7JCWWkbfrKhkm4OlHwPsH6F
SZXaOHOGU1VrmMrBDAA7MObV9YDI+ZRoOt0zYoMakiCfEHo950HQDBuDMs7NkgBS
JLWLYEBPTdy+D2KEtGl4jULK0Ty//ZwRMd4CqJcRfNgNrsthdoucUEFEFtV/aU7h
qzXaaXcb7U0KQCvi3GyhlLnbUDwx1oTE7f+UBS2uIDL5Tdt0+UjMxuu4ytE3T6eL
D8LaNNLf23L1BuQZW3aJCw1Q31bPAAEgPZ1JK1jc5BsOG5Ls8UXfw8EZhizkVn12
385FhYD26Vy36qNf+icnY11UPVhNdklXe9uI1xbDqG5e6BKY9mxqauLTa51cEgX+
Gl2+fZ+X7aKP+Q1qhhCCY3fHKhDdetzQXZwqBbzDNntPbL+qOtDSJfxu2jAYqM6Q
4Cc6LmNrUZGD6gKc0uNVweORyYFT0pmWelkmAl/IbHElM2AzfaCDFAkS05eeSqdM
bQStvveT+mAWL/waPpsxzmV3K6ctgZasB3EET3jNmsNzEiF4sC12FfnVa9VFlvwc
8bzAKIfZ+BOwkln3R/X84YQrjiDQf2V5/9AGbzXjDzb4uM1p/jazI3LjZqs+gMxl
m96+Zdza+kRk9Ol4MjRTVhaBORuu4a9W0hDGL5nSqKzwyn2H1L2mkmINpp2ykx4t
V4p3ZE2apeRJmRzWtLyZDyQNbJdFxFdTcM9wob7hALcA/tnAzkNmdcuy9eGQ2A3L
8uYdNdoRkqfTFQjiurI6MLJlFxNsVV9E04sImJQKrzPmt23vkBNtH4u1VFkmhRgv
fJY1btKT26KwK0wbouhRh+5Xd9Cne6XOnPpyHibMn59ZScGV2R0bctZayt3XvMmJ
lkWhqTqOLBP1Y0MdaegeiriLWLoPk/2Z/hnsRc8j4qWqYzwg2Bg6Ge2QrPI31jF9
jWfHAQ7QGuzdDA9Lx1BtidSMzQrUwQQYvEVijC/9fqNM8Iy1UMavGqtRYXlZ5iBG
hgPU0SDB2MRgf20xmokA7Pw56smM6BXLLz3/fBKqys56rl633dVlpZzrJqlHUKLb
oy35hIMBQS6wTy6+IKQ1In5ZhdSBJa+QVzRhiNk5rcjvj9wQhcK1YDhkiD4+l2JI
BbDvANc7eh69iYc058yigic9ZtAtu4LhNxl7Nm1OnlOcyfNY6O9JfW+YZWmWlTzY
9swaq8U6MY6IJaas0+PyXhvsqu3xeIqf5CBPa3skbZCacSdiIcD3wUcYcyfo40a3
iNcqHW4EQMj0l9P6nJDPmEp4/Rh/iQeW/NdX4CEE66zWb4qVP/rIfynNJ56YZQz7
E0DlSfbZdqXaPdXMJfRRdbivf0zMDQlYUFeOfj8FcB7WKMMxdrypkKX6iTHtIwd9
uqKLLkSdYq1E9nldCRKpsGPVjkyS/sfb4gzTYXUIzlbLdhrF/d5sb+EYofXCO3HS
milcTBF5/h0GhrOPfwkRXHWAVeVQlUPHK2E7ERcVWn1YbeRhUuSZTsFXrVa5bNtV
EHVZI2zIaOikB2p1ebNiZ7wEjEjSYa+l2Who1gxXhjg5RA3iJi9HlTMP+Xlq0Dj4
rKTiXsls86e0Yx/MmwV69/gn5Zxza/aXfEu0aX6563XBzPKMBbmzAMwRM2mu1zYh
eIlscPdQtiZ6FuhJcZvqEfLqW8meO3ZyHXNkoYQoh7/P9F4iuPa21ri7WAk1tGkA
CIcUOEQF3drbWESOCvnw99B/RBBzi5y1QruPQrgWu+DcMbuGQxt7SqzPvmMPQKAF
E35Zmsp9c41ng8vU4+1DL57FcAkRO5W2srDqOU3itQ0h5SoJkVzQsQduk6sfA0VQ
4vW7kDnaY3F7Hpcb7uZUOU6VSGwo3OEli0AgNt5S8KdY/imMDn+De6zsLqDMqtEg
3jUKSzzock7Y2FIT2scgaeacyIpH4dIfQf7lIEYcyImNaQv9rTWcCBiqKae5L4p4
UHRA/ckyZH2g9hX09BEsjIcZ7b6SderJq+S60AUWOEsC9eJD+SsglIKhG68FAwSZ
XS7SFqEbDlU72OrkZa4cCtqZsHXnn1tw1TwL9KxWw13PAXukaUfvXLIv4aXBCJw+
n/hOnKvi9mCuxEKVcHTZIz4G1NeGbn0ViX6bumYSUkAg9Bqk7eZ/yjdTPppsDbBz
9LKGv3GJ9tVEMgRjiNMMYKvsa6/WoGY1d7mXCVXWjTDhiheLfkWPDRMbkg6pnylM
HR5ohI6YoYomZMm7rLKG6PgA3u/xpb40L4cM8LTSUJA69bvtKOKKk2lqn2xgBHGW
6Wl18Qnt4mmXyA4ga2HQTGpjPI4BdEjEpVQH5Trjd5ncbKsrouUFZLA3mXCxKYI7
gCBExX7bmXwNgNgE2tuENA/DSdSQWdxbXmPm1T8/Rt4XqxY66Xovp0z/T4Dafqfs
Drtl0HLaWBzT18Yxk9dGwdwGJeBaYqdCkahwL9DrWgsbGSswmra2tuUB/Rywf+yk
a+U4GRzzkRsoz6T4PZBYtkyO53sKSY2aY38TlCOTz6GGSlgIMj9+Js4Kg/G6IVVt
/mpRT+kqTfgc1FYc+jnIb93cspSkqwOmrUl9vI3rBO3376a8rE0TPqfgMyCYWvjZ
UlQ0BSUz4ucJ8eETW6GKEvaoOuDma8ld3OmqAZxGJqoKObVxz3RUa+GJSdmu+O5q
t70It2ey/g8Lm6f8h4ts5NR42yNwZKTvoX4t8dw6O+Mh/fhqJ3/xOjX/6aumYxk5
W+7FC+8nhp+cKdHG6Iyb4kiZib23sz/0uL7H4BFKRF6gnVwww2QDquiOH6/pfX2e
iw7IbtTud2u1vtmDbjVackgTE6X4dA3Ov1BBCsuq+cZi3gTX9CUo6ch7mTC9Xq8m
M1EKIZGLImoCZPD1MjvprVd87p4laiiy9dNSt33UqIuQG1lsRhulPGVRJR8+PuJo
OI8ELe5NdravpSF2vNR1Nmq9Or1rcDo58SufVFZ3cK66TgcXROJ+xgt+IcaFDYwU
mKq5eRvPiuAyWTJfoYp46f/N0TBmx+AuzkuXpMJ8CxuWsywvzqeWN9cZZn5p66jX
GywN3JpcUm3LTQ3Iy0bPipyFkhqdi8hJDwzfVF4EafpqZWn7QCbQ5SaWI77RHtXu
Q3XDfkvkYgdq4jtkqTTIlQSDiipEgbcCyQCEenIz9GyS+3meSyQN+fflVxP6VeNw
o8gAKjPHIW9A0n3PBPX8b3aByHtfkSh4MTzv9tjNvgYI97ZqqbtH8YFzi+Yp/ghs
+ToyuwwvcNYVBQ4nmlJgL7WOe8whFpW4d6LZSabPodAnxsP+m0cV+UxCuegh9Zs0
AjN3k/pC/BqWNEM5wRK7A9fceix9jCATKITQxd5G//38tAHqICyBJz0Xn8qeNW/f
uuzPk6zONYaBqzWqs+r5fc9ii08x7eNxwOWVR9WPjzU=
`protect END_PROTECTED
