`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5d9csHUb8kBz0X9Hq1vSSrdO0q1wd+/JsGq5rDfqrWIXeTs98lr62r9raVjh13k8
fwO7sVPD8C+0wqa+kv/ZrrdxvyhCOkag920oqQ/neIEZZoAsW0lHb5LoScsrIguC
DuXjsvm2j955DN2oOdZmbUjvYpUyNTmxRwOoLAbkl/4X0z+GPxOhdiQjT4vlaw4n
yxcfDBMviI3s49NrvXVQ10jCqjgyMnKpJVnf0t9KcHmaOR3VfbcfamJ6ONwm+PKk
1bTd4R+6OjY9CoiA18y7ZU4oWnxdmm1gWEMUKGFuomylHNs8KSkjFewljAvtNe5T
NfMowrgRURDWQpBFggZ71A4+xRsugf2xYW+7qdGZtBOUMEMh0az3Bs4pcdhsKH9i
E9E0PCJN/LdTRNEuAoEuAUCaXfT6YoSh3dLSlLLO153Wp/xH33kdYozSt2YmadIT
nPEsqSzzTM6Ast2FrRD9R3Dc32tt6rVVuUw89wfSKYLrU0MBNSRQoYrbpWccQXkz
utjutkRq4gGR6fVH3EbR8TR5CZSdDVZD91pM6VJA5dE5oS8UpX3xIfo+eCSodT0A
/5kztHw9JqZuHj6w0QGPD/AFSblrcLbaG4u9Mlbcb7p04DTcLZv3LSNpUL+yXe4i
TvI+WkYnCTyHGCf3rIa8/GZlC4jb+eVBdydwzLPB70QWLKQEoskau0ygKeBcCtlA
8dg+gFu8cUIyszA8t1XEnqYp8X2zZPVPgT8NzlIgCKe+JGTgglpO8JFMSWnI7T/t
vGbCzBco63TmjlzLs+rGzx2zGt3NR/SE5+nh4KfGdSQkXoPX+wYNrJbOQQ4fwyfg
r4GolMrjuAWkMmXEZPds2w==
`protect END_PROTECTED
