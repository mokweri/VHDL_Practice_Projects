`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9GE2fsxcNlMN4Yxjt9b6xpiaLfJHcNqNjxSTbR/nJnqMYZCxdtCNIsji2uy+5F33
ynYIynOA6c2K6XE5Kz49QVuIXeR8swqr072Vy8bQsTsYzPmwIgMcEVgzSrDAhYfN
RWEBuxUCZWHSUBa+XUz7x6X3MiSnex2JnRcQQqWdwc/ZK0+fko6zYU/olmxMj6Ap
KIRwD5KoPJmwv3krvo/nR7T7ErtsUgaApB3+XEF5yQqg8q/1Ic9euqdbOYXpTFXC
nUB4j8rpGCFZiKEIv1A2xk0KWhoMI67YZ3y/ilNVV9WGuxNO2iCJeQBnhK0SpUsJ
YIj2FYaSvGt7xWVtAr1FwW/971T/adugFuxA7T7+1EobOZM9PmTXVYHWwoO1vpmD
dguu4/EvB3Ny5y0foSvYHX/k3z2JGN9YGI221wNC96Voksghp/Vu72Xl23bg9isB
ZzZ7dyFJ7Mf+lH7WMHaoy6mBjiHyk++Pm/sBtlQs12YfZ2YZCW28OKaI6LoHJWvr
2QyD0fKYAI8jaupU1m94XFnwnRFsxKcCn/0EenD8muxFtyOGqgw9SnQXY8WcdqQ8
cZYdQform/ZQbldWvStEXEOwpazEcGdb8PoyqDy4pY/Id0jiZyiVbDxOCMk4U7Zo
beln0mTwSmnge0HnE5VwIL887p5Kei9MzbebXeVcgA9u9HOKloLBZ/z3dJ4jocxs
VnOJt3TUD6JRzVdDgp9wEW/6zEH55UYEqhsHfT6PwStDqpiirGCYzjcUG9ISRKF/
OYinN9h2k0dCkW4CJFjFzR2mmBRq2fWsOi01FclXybVdDBvn2Tkn/vp7a3wZ7CzY
kgTTaQJfUVG3YEYA7iIf5QwmcJm3hexRThn4zKpPS0jfH0AtrnumRDTAiYPdv61S
p5efOvoJuBAFZtuBxhHDKabPhi3GAYH9q8RXMiqMN44=
`protect END_PROTECTED
