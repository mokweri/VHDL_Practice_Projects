`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HaR6kRh9RuymfsKpHWOheSaT6coJDOiRg+cjfHaMzQ3ExLi4wx4oOc/5ULm3bftj
CKka0acRWCAlqPcQP3nBNp5UjnR5AlSJnHkDTb88X7nbxFdPCToT2vANei18czXw
B8z+qHcX7wi7Fk4DUR9CjnKAPFSCQzJohLbSvLIeIhRwgd/86jLvC7WKYlBn/2Ac
eUEMO4g9zcHgOTTgFG/sweDon5ReX7aU+rWG5TNBCpPi8WAeec9jH5M5GIMLuF5U
qL/q3J+6bXkf/fKG438XZ+n7nC2DPm//7QW99haF7bmglSCoBU1Zg5SoCtbizX4W
g9Z3PUHSdKW10azbrXg+nCrxAKn4zJrLaRb8qIYg8D5WdzrTWpXd1rlWXM5ZC6T+
S2q77gAyZIsXwsF4dUzVEmnLJneewm8JbrdLZgh1Sxbx2jE4oDTtha6CMjeqU6ue
W6hig6k97X7S1hQCVLSkbbr+KnqARvgc5uu844DTyyrqCAf6uVwpMvPe2GOjm9lp
JGaDCXcrguq7SUs3GCLR23prm2Wr8kRWhkstRoDr92ZU1AEwnusrmBZWjxdLOgrd
5xblPiA3cu6q7P6MLvgbVAo/YaQFl6xdIoD35BTJ9wWkS15kYLsJjlqIJr8b6QNX
+QPJFSLBPxodFrZjQq9fggptIRhslDX2xkqF1+Al98Lm/J7W6zTiha571UAgKj13
fhKK7+sj5IulBDDsKuGbeleJ1m3LmmxuKHfdpUDEGZ7bV46ZiWJXM/FMI45amDwI
0NiftbuodCMFbDX2vrhFiBc3O/vUpoNtI8C0Ce2nVcq/6iXBOEh4Y1TG/ubXLFzI
oVzICYAveqYD0BTM93iX6aIgtxTvOz8lOUjEVdvCxWVNMmTpWNLRkTCESXyQZwYW
epD4YXgnXvRUx+h9bzLartJA17fLKP12/NnWACUUmizeE7GK+w5uFggTvPO9uQWX
5araLbcL09NDPyz0omCICEFlgHkUhu90GTQIndVfRL2b9KpQJXX8Kv2wSj5Ho7FR
VzIlKaXU3NnCy63fuU4kHKT2Zrhv4NaVI2zi3zaSxvkBlmCeI464fFXP1hGDE0/2
WQ1Bu0zNRkwZj+WWM64+gBkbBK1MGHOqZS692qEGPsqUPfIr1RhewZNK+UXtrd75
guUH7BkgcIHo8CnISImXgIJ2GHZSMNZu0dUiDfgD+wjREOCSJdglfBWRYo6Lg61z
hFMaILmpdmNRiNMXMUjJWxEBxV84DJ/EPCprvUq+4bDhAaY8F2igZwcaNnsmR+JK
crpx8t0O9+C1BGWCu7YkNr0v0TxthApPkLxl3z5SdlbGGckGCJAPsUimDJo5Q6Ie
UQ+I5Yv6BlpZOVupCL59r+vblgj/KobeyDW+KCy1UhylIJOIOdtn//HXZvWRsjch
F4E2GqTUvLVmA8bqFFWnLQT81K+QvOeS5mFqemFvPMCnNom7Mr+kcnC4XSzfYuba
9cDapk8g7zZCUyjstCdrY+J6Je3fCo95WxFN0cveXhWXouRwhbNtJ5zh07WTPOdl
wSJKTfu+bQsNJjiJbeT9VfT8aupSsTQE9Lpx0L9nWT48CwaDqKmDywDCZnPQR/YO
JO1WzsYopv+fyRddSsx4Hw==
`protect END_PROTECTED
