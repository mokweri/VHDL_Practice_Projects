`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FhP4rUOi6JiAgx1LV9RyDtRm6Kn/6ksr6nr13VU+p2DpOwhk40AXq6tDGhe0QEx/
ZsB2p5G8tCu/1EOvruhZKuQaCtloW1rUag/5iGieO7MX0VoBtvdUGM8wQFStcAui
j0beLdo/Hbbh/Fju4eddfu/lmyNVn5MKrKKnb2u1PgoCyB7mWT2SY7fPSckLWa45
fLswJ1f2MBooMQNX5pyN5ShNBNyqaF+cNk7WO25fYml4vRbXSbS6IOcEjg1B6ri+
4by7E4xrlCKRtR/OObzVxOSP/qRrvUViSSj4gCVUhiCNB+ETDkMd5aJyTR07Ygwf
rBNXLcda8xnUSkOPz6OKLeW6ssT8k9sLwnkMZPCaDXYXFAKecr7MUsog/5heoMhH
7iAIzceWrSVSE5r9qhiKrc2rQ6xo/yhT1kqli/IUgmaaFPKR0FPr4XUbHPwjMf6A
`protect END_PROTECTED
