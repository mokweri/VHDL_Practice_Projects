`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQkUBoLu72pHiPcoloZg8ugz7ry0sceT7Xmof35oIwaR83Wo3X7PQtNIy3A+/ycN
/LTSjZRWsE81imBXRCDiStQ68U4RjoVkU8L+oH7rDFkpPzD+Dzu4ppVTelEmP5is
tE16V+M5syQuK/EOGiEWY6Cfpez51pM25VD2xUxt1x75L78CCK1oUKp19MjlCFKy
hbe0FMem8OJn5qQz1ZQMXDdbxmtmaxoMoXy2U45LeJ0fKSvrz3BgI9hDP4kD0ky8
RIfTu/CMwaRyUdRZJC/1FnBKw9h+aSxiJPB47fagZjnfOfpCJ/4K/rM0j+p1wzir
8yvmambZDYwwA48+zjxOA5JdqwP74ZHCkuXj9QKzHqnik7WBtkxoj/VURyzaoNf0
xZH7GDdnlwYaOkzz0IDS0w1TiIVsbES42N2W8evJeU04/sZfL2+k/WHww0RMCX8e
wwerAH0j8+BCxE+IUUeKMvwB1KbyWdM/6T3tNzcH+zAvdPEn2WNoBXIBKc4gdvYB
6ablOIFx60U9Gd9VVHKeFUDxKZy6MoonCHhQ08cm/wJHkeQKHSl1p9m54EWIbSHK
idXkEl8VWFrx9w4EuY6YCqBIXmiIS62TvOgHSLFZOum7ujsDWDWoUUdm9sd4nivd
YUUHjyvva2yApJ4OXZ6X5y+W62vBvRr0sBJ6dhvxtVpal7R3R2cpx60qc47b24ma
36Mnvk1tbCNaTQfPUQmg4yZ7m6+1326+YtH2jvRGsFmCVapbnf9Jc8BNv+T3Yzf3
7qIK967SlrIZ/QK4v0mE/uiZyN5aNewXCCiMy5WNGhHPWwYd7579eIfLGWglqA3p
YQ9d4JUT4elpVRpdr2bUTUnbeVRrstaLlhVsTkr45scI9ph95JFPOTObqntJ8EZp
bcfUiEkLbNl8mYX0rBAuj6g99QKCl7s35wxlts50sBiuq3t7+femH3sYyokC0jzN
w/snyDe8Frcu6AZ+nxR14WfVppHQ1m4nHIALWAIVyOE4IIbDATW0yspMOe1wFDzV
7oViEMz6YULiYIAq4asZVAzQo435g9riLmJJ/tXNIHn29ykgCKf4IhQ0bkX2+8Pg
AMPGpIPBSEMxZFxRvz7xKWH95R/QtNxuWefBjlXzgqkI3JEWj2Q1f2L4TyUpVHwj
JEuJiVhc/KBt+opMUR/C60E1z4a0tuO2HYZh0DrEcxsL0kZrorX02DvCRsb6bipI
IV9YjfmNx6com0VDN5cOmxwggT6ep8RUzKwewIKBDBaGG0rA8lONtzNGbNu9KUmM
yeal3rRoV3+Q/t1jJYW6C3vX2OnT8K5bhAudR8UaTOxX0uVdUWKCLjmkE/4GdlYU
0jUmLGGNMVmX4YfcSW/c6Hum/Bm52ixgjsqRO55RuIol2MhY9JRxDW7eXkoEguJk
+/TJtFo07qkgY/Vk7fftlyz7gM9obrBt44pwBKzuC+8qBwRw7MR3i8AKyWGh5ykp
+WOjsvyk/DWRW6+1Ww6d2C7vaGzt5OkO/q1WrkO0lgcK0u31MZTIDRXXRm/gghs/
H3feSAWyNT5XDHXV3gPVH6P5Clx14kpAfhRSfiCJz85y6pFLh8cFVPWnwJpeaYw0
ehW5DJmTaajl+McSE1TvocCg200kchvKwdTQPfoFHz3Y9cS8LAdVTSvee7v1Atk+
bib9PUrus0Us1oJuwARrpkhnIWXJpAtXwR4TbE4ZtmT5LcAYJAbEhfHx1Tf4RkAJ
f5dUaH8qFyrLMl6hYoe5Dw1xM822S8/y+PRqQvkH+oio0TXz5ZfXN7gjNZUXSLtW
hfkmKsNneCOQRXeC1SgWHjfcgi8Fv1J6b7MHxAYWX1IBwOVllehglzhgDEQEN3qS
/DCTSt36Do3Xa7/4U+luab2ljFE9wyqxTxLd6MCoR5J8LGrHkiJDX+7gUuiT+Ge5
UmQwU0Rj+LlPqfo4yy+TCENh7P4EP5lVVMLTbeXPQ2Zz0Vwql8DKjXnqK81ZidH5
bwVypfD1MuIr4Ue6BfWngN+SlybEBwEL3T8FlQUBGn1iGmE9J+Ir7gtyzbaQMp7H
dxXm3inHuIB/zrV2jYmClA7O7c1i01kFUKCo8EoQjx7HBSQZjga6Ih5YZeD1mGdD
RNf+KT4lUpPkRRSigRI20P0BQymEjoNwjJ1U+6NiB8auRHwx2lRCyyDnZewZN/Jp
Sskpd+Ob95MZLp7yttMIvGdvIvGD0YabqIE7HKpnbG3e2vSmRLSmSsP8FwsZFhyM
BEHq6emKd/0+HbRdhWD6IxVWk9gDGY4oFhV8USPrAdN3RV/mGYjXXn6zkotrdjWz
ipaCD6q0SjlmmnarrFpKhR0OihLoXgwRcm27lC/4GIID2SZV6OYNVd7wCIslWYT4
VzDk+YSODJo8kYhTQVp8MXe2yTPwSUZoHM6AbOyXiVaTuIc9130YEWITdpvSVcGH
3J7GkvfJnyVLvu38t/jSe7yl/5QmuO3Yu3Ktc/vUqg+Lpm1hQMgBQ5WzbWo5kHln
ex/osGa8q0xjDazRaoJ+dyAQTAIuUtylXgrX2Aax+3dE2Mhhy7TUDUe88PMsbiue
MMeqsQYNFdrjaASMvZXxJWnT1zTM07SioHKA7mt7DSFMfnwl5VdTyo+pNzpupmMl
Y2mjQEPEyEUoHHHddKGPpxwB3RRuvuSCXKz7YcFzIloJZup3kooiFuVUyGjIxkDZ
MhOvSr0yvBxbjKCyhs8xBmhrhBLRayc0IVevI+bW0xM4Z0BFBam+MD179b8wNnrW
5yehL24BT4c+bcINynhJHXPbPm72hOWXD98DZibdl5TZ9FgPwONJHCzBp8jrAiBk
EaVFWCurUyySDftZQNEWaHv+qEC4P763/WcosCIu3DLeu3iI0VQPx+zFP6LfjsIr
8dwezbSjROMgq6/cD8mUbGEOts5fA94Q0eMSxCReu/CKitB18ANjydVkKyPhO++8
z1lpvznqiOst8Ao7+U+mJTpbMBObgAdFADaMdIngZLfFIg/u7BDjuJYLgaIKYXKk
0PdDKCF7Z/uxs/DgrYC27zr+3KNlyVvZVLLddH+kU8UnXcT4WVx3jnOfjxvhu4WR
rPRKtHG3iHBxFPh+FFbhnRbaG7AHin3gidDa+mXn3ar4WbkTLv1R2m3Iqep94bd1
YXxCEk6z9HtZwyWhSPTV83pt1ePaDZIAb2hlN+pk6kdyTqOO3KwnGwrqL19Okzj+
TPrELLebPbaQoTLAzoCmGb3ihGFzM2oPLJtRaEajOQHFaWv8Ixu7n3L9INxTywFa
YXc0Lzj8BaChwFzwGuEJFrfUyu4DswxnyuF20/vJNJs9KMzhg8X02Gqoh12YamnC
gI7U0HjrHEEaE/P/aRAtfrH5Ph8dfADNLrW3dtqGW0VQ54ihNxNzyOhgJ1Tva4CD
9Z2YzIgJrn2TaJLonLWbVYW6tMSDvB7p4BDxveh0eVmxH60v3o49cpzAciD5Uj4N
LxFEif0hlw4VC+yZY3bMsIAlUXAWwrckmdSBix369rI87syjRCbwlMxOP9W1TMW1
QMvwKT9B9rv8hItst0e/Wf2LmIFSFXtOiJCBPB3+Bc4Xl9R/MP1SAArDRElIiQHt
vUh+nMSZ7ZxNUmZCZsxNXAKCzpBgJ+PNagSPeOlibZuiwJvwj6Ks+F+Inhb3858p
Q+I4yUkIJT52CRspHs9qDKdNp++Cnj8MH6Gjnu3u7UaNZPwnS1zWEWJYSfXNtaYm
eUDCNxGcANWpn5s+qCeTsOXtOe3yW+2etlcbSZsxL76A6v6defJqxpm/TRFKFUkB
9ZMVIALWWT+0tqKhPI7R19P5TSscjQjnEO8/G8V5MmO+Xj9SBf5siSKb2UUCSVul
taVTUZ5s/KHL511xJ/YJR6DwmoY+/URBgM6MxX2j4UhX0w0vMYm9/PyggTi8HIPP
VdnF4RHhWDp8JhSZxdTK2kBiBngelDzPd0J+8jo2FQbgIa963XjBwaDE91lj4ZZt
iYLpmqjTNmSAEDv4mWjJyzOQOC4D+1hcYorBkNttb9wAlPVG61X5fkxMgNpidBt8
lmLVaHVhrUMFeyYkvGUvOK1SA/K1uemfCdJEoXa5TbuAgagheOORqIOJlCOlvBJi
KjSys5PjlSBIic+xzIYGnFegtUp5463f/M12sbUUlgnNOhY9P0+JlOhMTY/57I8A
+sDB4GnPRx7zWqz65vpzpjbxkQyZK8peVkooego/i+d9iXY2wZFgLoYjuJ40DqzM
1EeO/qd4yR2jHr0onA/fAO6LxgcSStXLJTxSR7l9onmtG6DiP7nEsoxaJUSg1WjB
vkUfCV1nVKidTwMq+crjxyafDSUsHxfYaY2/f7mwWGuL2A7agqScGsU/2mzbTQtg
YFV90uYX4ljHyFPSGc/U9doYlCaspe4gO1sbX65Vnvzv8KKTcwsPE/g+3AKdDgcA
Ms+3x1Y6scTv65AjSfva8ijwMOW+nJ8mCdwOrIYHioJ9l2o6n1VRx75FcHopZFVL
JRHRQf0STop2fXm/iLsOa8rRHXUskmxRvI8oz1q8Ug0NUIrAoVg+PSOlKBGbxSDx
KmZhi2WzwHClWC0ZHL5NpiZOeIfQKdGL5cMffBxeGKS73bDOiWztFTSAvMOnRj00
nwVG/QRBz93FFU/Vxst2s2USn+BeNWBJsw01ROsH8l8O9BnRLSlsK5kkqbKboaIH
Rn/Tzqx9WfkMQ7KlZH1A1fBLYrGmLwD7KZ3C6HwzHc/9dQQDXM8j4PXWA33+iP76
6GYrDK90T1HDqwqlBmexR2NWE+lPrQIgBe1WUOxvyKLzhC9ED+qcAEp+3mGtVJ7/
OHtf1h5L4CNa0EjbUKjMVO5mOIXt2U7EgMxMnH3/QR1FEpoTWCeT8e3Ea9Z4Vbs/
oA9K3f3SdblP3qVX8+i89ZRg5v+xt32FuEpd2OGLtIBHnIJAH+U4fUmuMyKmJ15p
f4zfB+aLqQRTECDv/XE8OiPfDwTs73brmGb5NL6p4yQhbWX7ekmViiJOu/t62xkS
b7KMF5wqWIH+mnhYNPWubjhpkuXWVw51WkWrIEsVF++wyuV/Rg2qGO8R8ySxT7Cc
MYnayU0So67gxH5XKU7wXM1uYAUqeVdlIphpjCdrCZHvMj3dWfTcG7bDoWtT8gdT
ugEyYWr/42OLOUuJmZtQoZabsWPPzwRhNOM4s4HRVpPn28W2PjOJxuP21F7uVBps
M7ou+XuCK9SXX3CvNGdMvKifGNkYrbLy+vfZWf0eh6B/jsmz9stNFOD93N9TnN1c
13uphqWAr/ZHzRvbs9q2MzkLwEADnD7yeGUFzCX0KrEqdDe+BJck3Uc+dNmQ4Usv
8XSGWaaui+6HvqeDw1mhg1MQzS7wZZAKKcsZPcV4J8vXe/5uR+UzmYqSevSEEOjV
DHqpwAte2Ku3D5KONv8ZFhIlc0PnZhoSUkf7XRkqBjze8cSjVzdE6Nje9HxNom8n
T7JRvy7HLWDRPu1ROaGX1pH4QPamgRCVAypu1ZaMHfJkQZRHvTZX6PM6p+L3n+qB
36txfTMjHuvKsAhHnMeUxX6iDDU5IeHgOobQWZuWfBJtq++aT4z07vcEy/vn78Wr
pwISbCtgjGvQvHfaZTEsbS4EuSR19uliuDzbV+dPVsGWxr/I/8wFv35qM9AG6kAL
2VmJv8KZGVVtjajBQawYriWwoqfJ1qb15s3UdiwmIIlyoTQ/T968mbIQZo1090w2
a/npJxtqrQvt6bkQPIKIPUByjvxBiuZqiIUE4MaVBxbrlfYVtQ5ydmcSfxMhbPA6
y7nZPT5aRQgWVOp/rnRjEirlkAp4E0hftfD6bkgcgaFQiJpa6FliMEKebbToAz7c
yOHGb1+W1r6p1zj1pNTL/vtllnQSuN11FH2L10Pq+JCoEopEuoEHVHywKi8Z3iq8
EM+KjtyjI0bzO2I+yb4mbtS8cvQWnL9St/sNZjzOGpRBnMh5t049+UjSZ6xONP9o
Vtm4IhlikFrKZemkRnO83pgHiA3pu0t+Sn3GbVc1srJ9rOvXosMxJz3/TEgp7Vgs
T3XCVMCxCKY4NGkXOGhg/MLkyKyC5SvRc3XTOgwwrU7uQgTzLcLKXgmHnWIVS3Jh
uS5L1zecfZ8nyh80ro310wW0TeIX7mQN1DRCFrA5ECD+fphGi5y1fNTCTTsoh0uB
fLq1wOmCJpkDcy6HAu1zOJOYk8+Xe0lue3eGPRT4askZPsBkNAURFj2WLM69+xs2
3dTeSmiAOz8H73AYi6UHAZfo7TKBCGbIAHlZ3pifCG9MhhTM+O5Uua0gkHnoIaUm
cQ0dfTwLNVdDMKCWYNO8pPUPK/yoUj2C78wwZtKdnAsnnrbtfYKA7haObAH6T+PN
rei5N9G27yJepj8LW0t5khj5OxuKGTBXjmaHskEsTeb5lFEfGhzj2wKjDNY5bBp8
mAK2a1gtAwndgrt3uVxDJ2mzWqSpxd02jn6tY6PVIyIJ1ORiE1ts7wiWnroldev5
PGseXB4tImQuKmXjNeyFtgAR6S9rT3OcPpgsTMDWiFFl21beDJEEn10Z84R7mt1z
+exw3Hg/w7VEV33UACBlrpdIVxxMaY7+r04Gf/iA7Q4nVNwgvuJZ+7IHx8CWtbES
EkjlucbBkBba8MGIAhtW25ExxbzCpWTqF6QfW29d7bHI2LKl/rrvQZX1arSmk+fv
PXQKWwTAO+5wNlSWJb+oQNz6zhkNW7vV9qOfpBQJcrALMl5M5gIUz/hNvhub7p4U
oWziPMbkl4WcYbwtWx5mRNUpkQNV8xJZ3Pf+aJOAye4=
`protect END_PROTECTED
