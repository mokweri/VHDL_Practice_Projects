`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E6t/Yq9tcbO9wOMrVDR1c1lxhMQTRA3Wqa1MbXB5dgzpKYy+nf6af6Fy+iq1QtA3
8z28r/9ZqOXRN13F3KPbcBYghUOPEsrL0Fe+TfJwSF7C5c2vRM+/xR/JcWGoDgi0
N4OecsfKWpqONwRJFHGr5ARTK3ka9C6eWlWsVESHlpI5vTriH9/ZFMV5/+4Y1XfZ
sqRaroBK1Wtv25P00Y0adCYfYAdqnXNC0xqlBFYTJVRClr4kF3IU2jfDunUzdVct
qbV7m9djFtf5dOC/kjeIXg==
`protect END_PROTECTED
