`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXkfAze/PfDniNdSONFJf/XsQzoQBGPw36N5gsDf4lxfI8v7SV4utPVdXhxrAB7S
d1RuMqlswedGFTvpV4qBXiuxNeL5e6Hat+ySg/csTdYOUvbWLQ9g+t1oP+TcFbD2
WxehL6CXt81lsH13D71lZtMREI7mFxeTKtshi6WyJICojKoIZSDVu+QDvIg/zM+s
q+ViJUnf7NAE6ICRdv6j6BvHQgWTBW3KU0Cu8T/Gr3hD6S8ioRRQ+HEVHYsw4FCe
w4SJgf/V25NqJrNZUrbgflEviyZjzXnNG99jZofd2GM39auLbCuATvxq4CG1t6EL
k0/sYW361ukOTT2mQpKCDSwe93CUpHwLGQx0J72V6dRF08gQGNyLeNi8kK9xmTBr
iV3vFWdBy5HyQS+4bh/qi94sJhmFwvx1KrMDiBXsUhgCi2o4Mcs5mgRM36qsQtQa
pzHg45ouPGc7pfIecwjZJC7FF+zNCbuvnFWoRB+oi47yl12tHjJ8bzOyPHVA2siK
fz/eWQZMmPiGyVeIBkxr8EG1ChsCl/U1Mu+7CfxMzw1th6igNIL1EO2lhPawYusP
TjMUZijjsVRwQBoy06DrlOntYnXs6wVBmSuRcmwXEH+y0EcXam+cy7Wl2jFcfs7/
P88gy8lTlq1Yhw9BNOHRyj/sp1Kg1hxj0g67q/AlrQ+Eo966PlKnFU+mJ2mZ2Nnh
`protect END_PROTECTED
