`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCluNcMBoi8A/ZHD7n86HXxzNqbeZeqW0aNTQ97D81pbhqUdletm5mbhi6uW+yNY
4CX6DMxAJ3wCEXWxVyTvihYqF1yhEJb9/ha+GVsQR9ig+5dp2R4RrerzIqJpzsFG
QjZhNDL2SFSYhufV592DolTCJCO/r4Ap74OPocA6DeuZ67ojyLqQ93Bm6wTmxQsu
c+PV8A+B0qaWP0pa9Wff/n3KQmKeQB62qS/oc9R0dzWzo+s7fdFFvIcxN1yjdphS
EeWDXgDKnodPfmXS6S2GsGw7R6h2vaPoDU+hunoJlRPZR7DgaxUjLQlCPa9HYu1R
UcsA+5sEXJHi6TQjAsM+qpHs+uYEnGArWUf7d5LeqfELdl9+hiYNJfpU0537Pt4r
1Fn9hsuNAN2MKK37VKvAZf2Rq30MuM8gGtC1fATe0yMt9eq8IwJsLzC286DDpKOY
Vn+HFKZsQ1NlqZBwfUOq7PXdEG7kHGe4SO3dOVDffguqIr4n/74rVFp6wf/kbvvC
q4p5MSe8G9CFGuzJFwh8Axj2YO/DDS3nUNyOlIapPnZCKwIqRheXPW2koXiw2X55
vH0lL5YZoR+L2ptewbHlCA2gQkVTvVT5ehnay5ry1mgglKPecIJz+hIdr3esyt/f
3NznQdxNcoXbnku8ZmbPK9p2KjK9o5bg7aiyVpxS8ZUk/vetP9R749JoWGswO7ij
`protect END_PROTECTED
