`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dj2htjYrDye6ubsgPG3ekPGReUfGROwlBB/hIg9KJDAfIWHEzwiBofkcVH/Eqj46
ZqzTy5DSwhb3nJLUCWEiz/m1XSSAEVZ7xAPD2orIWqrlyoP6BvaUu1tOOoKSUNx0
TK3gURyT+WwMz7ESkfExzCArpwpQKn7tyn4mDAKGqtr/ddC1qf0Rzvjo/uOFmznR
NqmhsO5a6n4sJNgqo8lNngTpGzt42MvWaN6l7Nm9R86cHJTh+Q11NoUcJAOdjK1C
+gsUU+O3GKnBReGtCF4d62dIG2Mt3ExmBchGp9KjAvu/r3sz1aMhIg4061bcFUM5
g/0sfCant3MxD+Phrq/+atG30oVYxRW6w8GynbsRk4uRE71pO/mr1zhIHfVRIH2l
1Y43ieSCANSbMkzR5i0JDPUEe2q8rRF0eV4M2R/m0jBJYl+TXPuKyza57qWk0hFY
a2wLvDf10G2t2TOnXJE9znfwGnaDOiQrMhZ6Icl5F7wtLUJDHfbnh34KH2pftQmr
E1RdoYNot2hHWIGPU46sUlrSDUlRaupvvCZoCs/V6t5t4/IydhV9oJ6xBLTXptt3
yJ2jTVuQwgJVfprUFhbU20FimJMkZX0VFaXpMrW190q4qXXVoaljRnK8IIMLNoCc
aTBum1V4WQzXGrJwra1YQnCdR19SQzWb6/1l996wQJtzG0mpWxY2mTTkwk4qiMXV
nkViUa/bzknFakMFBQsJx9Gs/nWl8tIDHavOxOpyLNPyoMCJYVXgazmr1yN7Ki0J
k+KMNnNbYNbrjHtYMIKG48VOSHdylJptu0Yh/4T09tYUqRFZHHBWZtqcZQ0Ivkr3
4OJF7VxJSTmeWwxixXcULH+Ws4JrNPPHxtmUmlv1sMYFmjTMaoNCUkLiiWMBUbN3
jm/42TGT2zglbEE+S4qY0lWW9hVNBY0kCyfucGFnkGBZQaWk64txI/93Iq6z5Qcn
g+3KF9z9knBME3a2zpjYm+Ip+iJEbZZi0WveCuzjnxjvoa35BiZplwt7xhPDUyzF
8fbzC4R+2jPYks5peXrzVkwY0u7qxbJdjLa8JzMj7boBrJS/BsBimhri+0A6Dd4n
+sl0qmXAXKzPpXqSUnMnq3MoOfokgmewXn+6qPeBq7azd2rnBOKE4ovsiWT24S+4
7fBxM0JMJl8V0AH9Ix4plxvFqrV5YCCzfP5wy+YcEENDFeOwch9cBlFweUSWZS6w
07bNqi7mIscxf1T+jrFbHOx/fpptxlQKmVkkf9Vz65ZKgZqSITbDb0uDeed3kbQG
9UvYXgcWDBXMlU2d46pMDae601rPjZJrRo0CVwNWZ8YmFe2CWjQ3+OV86r0LU/bl
mLCYcidFpNve7t/bvrE5yhbSA0n7LDO/y/q27M4qOqsv6+Beqde7Rm0Dhpee3Ooa
AtGxlsZUjZVUw8IFYEtlGGFc0VqH8HUEc9+/UEFze4qtdoh7pQPbbx7i2A6hwVgP
/vHkdw/3mpocAdRIN6qi95r3CPvGdbFCKACr+ei+Zf3wox2dqbSN3fLhjFIaUx7V
Wy2BiwQaOr+okkMkBGOM1m586RKfNFibY8Hs5SSEbEbCQZCMf6neVfpbaNbf3Y1m
gMVHzG7GZ7qRNuekO44c5QOzspV3SO62Gf1JvhoErClW0oaVG6pupzHwsEj1T/KL
rBH032+Cy83S+VSoPjOj6M0pwUeQoNuDCQ8rbj7jIxfIT5kwmt0hlbJFikJT+j7V
cRu+NSq8EY0t+deMQygVQ1Cx0yigk7L0CV1xZOe6dVBg4U0n6yXClD6/yXgqkMHB
x0AGS6mkZ1ycyAerEaKpwd8AxfdZ8io/3ugOnigmamGkuxY27TaxK/aH53Pp/Lxz
Xru98bDHh4xGZ+qtysGwCBu32DKxR01hkMRqe5qbuht76+0+WYTXSKNTVopPL+H6
QidzaOcPxlOl6lum6qzmJYS4dI81j10JFZk9hyUq7xbAe9grHyaTFzO+0O+AYeyA
0TRnugRH/O9yV4ac/PLNeEgZOzERjtRHHWJILC4UWgzcA6a+uaG3xjWZ8+MRp6iv
YOoMKyhvBEEfwLk+bJuDpFFfcekiogmVtTJuHEUuOUfwvi+m520lA6vfoJjV6NWS
B1qRNg7kpMoY7ixT/3XtyqNcIxbHIYh3yrKXX50H7ZOWSdPYAKioqbJQPtGluwOM
PC0UVJITYyOkZeblKQ7mxnH3RDRpj6IQQvViAZ6iQ+ke34EXCiYdK2B7BPHdURvb
TxxPrDZXXR+PcIghXdJD8gdUOz4lSpdr7ZYh1G5sMucyAd8+ZM+bD7Ue1oH7kMXL
utsh4JlJQymKpNwdinjqjb481xMlqOWiy1jA8w17OPNQNtPgSq9LoNtI5z8FjgXz
uJ4V/3JbYXSdSYlMmpo/2V9tyQ0QnwYErOwSMI4OArUAVBsHocXCdp+p89FxUfN3
elLteghUoMXcp4gu1ZVJGgzorGtCAQQ/SHWuSFALXz4DV9SgsmZJcMlELpNJVNuU
R2dt9yMmTr9coDXk/Vx786yLfqsvFwo3xukadRzZKTBlCyjFhnDc7bmWgR8TcGN5
mqqPLyyHPG33AUgzkC/CJMGvsjaqKZdcZTqpraq9ay/ih2EaI8pFA6D742H69ayK
5p+xfZ33q+py/p8kqdCZDQKW8UGllU5wCmkA30Wej5xf2OJQwJtpWQsoBgEyApAT
Cfh7hq1O0lE6ckTXwTaBMXsrzcIrU38waxzdLHwe43egpymWef1bVBsGE9cZ5sCz
MR1htwBcJCNv99thiGIPjW2rquRCFiq/BvBvGHtn6be+jARoOism8FgTXc4yNWdm
jiVCrfVKBBHReKDpTJkFn/y9s0pR5G5q7b6l94E8DZeV6UDtk1FTcUQUaSZFl9Tr
GI9uAYWScN0T3NaQ4q7quwyqvyeU/7cLmrx4FXkObq8n3X7xWgYqFigNQhAJUrje
QKcluCExCMJZvT+Ka0dfrA==
`protect END_PROTECTED
