`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rjeY2RIiihEbwmPSQZs3J8hGfoMLDZJiKw1rklOl/ZI5S1222yb9DswGAbXwcSy7
jnyK07lSIf4lUkM3gMCG1wyRJ02cb/FPjyCTf23JaF4Aro57UgVGaUvppmJqqJ/l
OG9gjO6eH/MDSGDR5eIkOzzNoz1Th8iOBXB4FaYRqfZLjKVhh7bB+Fcm7bgC00Sm
GYSl2apDD8xc9KiGuoqx/lwU+HnSSv/HQKRAEdv7k3au4L8ZpuXJnrZGgKFsK/0O
dpWgXIcxsNR0AsTfAZi5lzv2d3pos88irR+XyW/E7YwhNxrcQMren6vBpwbSc20k
aiUSa9tei5ATLpo46g7Qo8VwB0UyswvjetCsh+la7ZSDyfBeJuBSEw3/9oi4mLeP
lvLyaBQdiuduo5EVLgq8EM3/F08QDF1c079e481Brn+veLHjBV3uUiDoHEesMqU1
zCbOFDDZYURYMzT0RgEISsM0+7Olg5DbLc8ffdF29ZaMwfw0GaUYnZYOKNLAoWKj
tzxNB6gMzfc6HfYlCf68fuhDpLoieCKLAWFYYBDLEMMPwkkHQ5dZctHS3LBmgQli
jzq1+CeKiRpwa01poOfpyAYTYtUFr2EtXikG9QdMs1CtmyKamHDkoHK55QB0+8MP
NLmzrRbqc0IkU3n9A4mebsbaMGGghlfHKWcUwjL2aASVZxYVUdIJ/Wrli77O0Hgm
x+Y2DIrHYmqjhQ33gXj6ekniEYwSS4cYb6tR74cLDSG4EWaIRbQ4kaE7VHJNKSfa
oHVaGt/YQcvSHQ+HGHxRXl87hg1AkPZ/40dqt+fvAjZJ5x8SeGlTrNM6qMaVu0h2
YmTHP49T7Q7CATjw7E84WWPJkPszBdznEJ3vUvzW5FmeLKPbvifWwiWTSbuS/Hix
qQoeaYmtRaEeGz1vXoC2ge/thHuOyFQUM3Udvnn8r7YXmbPAk/VTx3VP7E9gmotp
5Itz2ZgzNU2jJCwslXdKiXZgjCK63JV6ARmecDQcpxnEk2abBlg1VuZCWOuASoP3
iAQaVpc4MvfLPW5si1FQapjIqeCpL2m1CR121/4xwxBw1HFmaLVAJF4qxWq7Nm1y
/uIajJ7r9CrvwVr2C0sfTGwzqKKAMY8W6YnrJI2gLj2IQMXaXXTdpTna+Q5C4x81
APeSRhT6ULCyt4fSFyKZC23OObPulatbxDwcvbWAurb9SKhkUfjq4M4BO0dJpBG1
0mZj9qE+XPxVyNK6aKeseMqtEl5IZKq8Y2c73xOlYP4FNgugo0+aQqrDcFejXzqK
qN4B4YWs+GlnP8PyXYnLaqSXwDxrlHTq59a3d/Zbh3JWM0VievH5ouJePbscAtct
BB1PMNiOY63xGzRxz+GbXZDkwpBbmBZFZNOxknQ1tXI2DT5dRzYOBUYcOQgyVdAT
4+egB3/wjNu0ZnMJJ5brC7yzAefCIApd5H1u67fV1fo7Cc3u7ASY4OWo3R5OfWb4
1j7zM2c0SPGWpLcxJjyq2BA5xsf4l6KfNhkknvHv1a2IFnZXmuPUFpArtDvTd+/d
qtER5eDCACVIOp/sLwTchMBnyOoP2wekDT8gkQzwZI40kQ7HmtEmjUcs4FntfQZv
otU6LbckjvcYpbxG9JwR36Y/GxnkBi7H1wumkqiaqJF+Xz59mQPW6dzpbuAVO9PM
2dQea1eIhUZ4/PqOo+1pUAy71zk6Du7u5S5cfTySH1tWFlqSBIl772G4wt1/g7DD
uPorkL0vCmMYfOTl2hZZbZkz6n2Tvv+wc8Ob3eyOcFS22I4Wd20+E074RswpOzjq
+vQlmqciMr9g2uJMRB7zPfonoEGa9erz+lYlZt3D3YCyXPXHcnUaE1Exp1o0ZnEW
zIGCCVSWZnCTzyr5C9Q7MA4V4nhaTh3akGFQ1sjvClzUfqbL7mUiJnkjf5RWSbrq
m5iEYTUtGW4orl7QBRf+TOSO5Z1rV/exvZ/plwQoung11cZtOYHcMgXZuAHooy5F
tFql3Cqj6rANQo6WCtBJjx/7NjHCg0riSYwt+iJ87q9EIa1icg9obQiZvSQZ8AmX
41DoNvruxrFq9nc1XFTfd5UkmbHZhcNh9YkxcMJy2BUgSEKLXVcF1uuVB2upf/wV
938zioG536DdVyAvBQWqkGc11XWaa6uqbnAM1uDxki48VJzTknbhWgssdb863ag5
3qq+hZyMyEVLuuw40K5eUdjFoo/E4FKz6kp0XtobHaFuRfDDkiEaPE24NCT5hKDg
j+fPpCSFxOOmPvg5/f/Yuk1dfpyxVm/p2ztzdkHb8bLMu6anMzPsFT5AOYjBCJ5I
BAgxwMLEU6KEJdYn8mmSkRsxNl1dnsdaidiPRgP/vNnUKbFaX0DHADlR7lFvbrCC
qFgqcffEtOJqqcfSy+fi0IbLdTeOjF5hmLAMS5SaspH8OP2jgDaRBKa0IgUBlIk6
lcgcD/3PWihUgOfCuP9VYvF+8ha0liwBkWxk5mUtD0mKdTlvXqzI00Y6YSILv/79
gu9amZLfvnO9US3xXR9wzY4ypXimzQELsZ+bjhaUEoIrF9aVy8KFEuDIOjE5wRmn
FEuaTUAlnj90KX/CnPTmdo9KV3MbcB7n+9s9irUztCWO3fuPSiSmW+Svn5U8Jp5f
aRipF16hv4L5Rolla8h24bQ/bxHXIBIlIN1XLEjttcJNo/Kj1sx4HT+y9Envb5bE
0b3TKmbJbnX6MkeuYYl29ocLfhH1331MidPGB6g/1klWRewOggbtXOGtq8tyoIEL
Di5oQneukKJbeGJOQZrIfsgJeUEMZewilxwi8lFzyoX9ozNQZSppg1FZhTDSDNCa
Jo6pq8bxYeDKzs6oUpAZM+Cv+looOU/JgxjCOi/PU7BdzFE9ayz3ZWESDt9spZo+
R465je8d1SAC/aADrTYewfeAC8TjnxLNqLAy6RRvROf06iwLTS5ZCxiaXkF2uicN
KbDfJPTW0F2td5zeYVGpB+wF+sIBBYbjXim2+TTeQfi+NHZxIVHLeG9nMz3S7KQI
e9b5lVMFCPjBM6ciK4aS4Y8iySldDZ78RTAPo2mMPrJ8uh4T9meftNdCSM/IcJoQ
9E8b2c9qZjIlpOKFXRtJ3HdugsvGIgeFdNsMnZqyiuHsH0VXbabVF7EEJENrO7+u
hNwO0xRWd1GiKWXyWikzWkrOLjj+SQQ3/WyeLKfc0h8bv3jupgBY2me7ZcWDEHv8
kyefHxy7OBPW2OVB4rdex/7dkoECm/1nW50hcS6G6zekg935o1BQnduT3ulvgwfl
rVJ2lf4U3DTBeoIiSYaleRcgO7taP6rS6gMJfZHrHbUcR4/eODxC4SPOhCHGQ4m9
0GjO6+euMcHx4Uh7PbJZe1MQSNmkkKP0W/TZGpuMqTwNumkb9qy9SeBYYVPuGVnX
VzuPKeVU84Nxo2D6u9YGIGF4Iq51MmygXz3ULYs4PMDZKPTB8rdSAHunNAagk0A+
cssApIaSO8799joyXUC8SqVg3R9MwsufqmVLLbw6ireKWyYgXWTYQoWQRaYyTR6G
hqX9tuR3oaVUGBc3g7OyCfbWdqn+jdDETRAfcpFEqCAb5pjz6G3xUBZYT9V3ZW+u
9XtpELzEwDs06KpufIm2dZvLwlECONPceRQIdW8nLee81Gmf2aylAQ9xbVw2nzF1
nCyTSAbyA19xXzfeOcJEsXpb+9KUl8gyOGpphN8U5M95DGzuciW/x8SzCp6AvOQN
ug5SNTZDPLsle2+pzj8Yw579kvjMXXmVDzxjdJR27uLVjX9CXZXpemAVtMjrl2M9
Lk1O0SA506pcpZfKehwB7PMe9mGV1Mib972jy+FUbzdiOdEq3HW2JIi6JC4Uo520
L1uMZDzZWkUCuZsfekqpl0RxCLqcBS6X/EQcJUVK3qJ1DyUkJQXwD8vxRtOMSIJu
XvUl2u5qNj6+bdlA95rr3bHCN1vMOOUfr1u9PplVFnhQhh0W//+9y+as6nNmtk+H
4gl8sJe5BKfJDAI9U0cMyrUGnt1ugbsyed1k38l6K7r/uIrPel7XsHZ/OV7cLPFZ
iEWIIXOvLt8LBfxZ3mWbl0LmWXbCt4bC3uVn1xIawMGRYeJYzbmIiDqRNRtxzRlN
Ahf1WHROG7ls6UNAsXrUc/elAsybXcQDaj0i4ODdg2FRkRkriV+aBecE5WwJFW0G
pLM/v2YKLcg52N+DEITVlFss9n87MwCGmz10RwiyEutolyioQ19R8IBWxaECexRs
zw7WdhPvNauOSXZ0S1W8KVpW5HDxl9FprvLR8GIsFkSfidl+pgCAS+Y1tYZO55t3
1FyfcbNLNDDoIp7HuPH9BlKsASXPIJFWp3OECiBFPKR5CDMEmptou4LjKHU4O1cJ
dcYyXsLgfMBqxg0D+nzAIxrfOt/aPeQ3G467msnb+wVlN1tWBXre9IF5FGcBRLlu
BX5gI4OCFqhsrIb+vmhNpn42i2KScha648s+AwShz3+885oWWL248qNXsqIeKWC+
WfPx+Ae0BFpoavkjRQQ7ukDQjjlr/3Z0xHi6tYO8F32WPuAsjKVWs3Dt9c18EOqZ
7oR5fHR2mhfvB/4fO/snWLm7XVTtCqWmkYx6n06a+lYtJkPUXtc7QE4cCTrqLV4y
VfxUxv04d7Hl/YC3DjIPMNMA6S+inmLxW9y9M8TW1CPsVZNGMYA+qfmGJ6usgh/P
/fqNdgIzLDMtLQQTo1wCJjb2AFypBJzqSuF+DAhh94nRscKOrCa5ppgrUn0K9vjp
+B7x+w8gO1OUfZgfezvhrDSjA2TWU4MaPWSTWESThs8CBP+CU5jNeYuPKs4O0jo2
Xutt1TZccdCs7zwizQJEzU+sVbCPrv6Hsy7ZyD5eeWR5g5TzPMqB1uXXut3mT0wm
Ux1tyww428vO5KXJPSUu3RzN6YzIpOomSVlbY8q7i7TuBrmp+pnE0xM0nlV2ymHW
ltpOyZI2b8VLU2/EV704i0dmRaOfiReZSHv2bo+q0vUUyA2J4YgpXKvrZzjIDRo8
R7IiNKpLwoYNJiZ/v+WaBXKbTpwPvH5LHFPq02h7PJscaYJtbXNwx4gpyxAlwiT+
c8TlloBDdgd9aIGbySyTYFGalxDkKPewOIpEfcfUrx3RwvhfgQY8mpjjDharAlvo
jypnAMUuEAUgdcN3NY/pgzuuuTVVaj97ClQ7Gg28eySkYBcyX3AYJxPaxFyOwKUO
2Ue6QDvXkoCSKdSTk44ANYF/URUcTCG2E0TRM5vHMIeXTSHROVh82hCo16TkamLM
KX6DOo2K/vTeb1pWLzg8xaYlrFDWvrJySFnI7OR+VnINVfk5yUr7BUAVQ6bK3R3j
lh9KW4bxvKAYBqLoRjxMg/x0K1/ALWh4YXT4NXy7amvmUr60cRVBBFJXako6mnOM
y5DCeNaUO3q/yt1h42FVOwbefPKmC0fMC0D934H5P8YpiOen2h//yxxqujpncxp/
NLEHEB6Dxk0R9wlL06WH25cLz18NLUhbdqbjXN/Wjm9J8eDMw8HY3TTPsl+bTMA0
oewH1QSej78eJ2K5lwtAlOyh28fANL8Uk1R0qIANPXEter37fMab3ai1LhJEwBDx
Goj+RfwCdZpA/KaFrtaYmRsSNVYN28BEZItGElJAB30TMzzyDBimF/zj7GPHGrLt
HO3FlmRs1UUog4yz+99gn/8M/EZ+Hvg/w74zd8KLhw1aHs7LtXNYVratT81YP+Y6
E5ZlpGIfgs37DvqzNIPZ8ShdNtCDUcwk34Hr7mozRThK5EuPzabEudaABlTX9F3v
xbM8ylvE/eVzLDk4h7SFE5dA+fxtvEeAwQPFJb86mCE0UVOT80ClECVkDmGvBybd
mWcIdSkVmEXrX/7VON2chS46LM2oglKCuQvgC1eh4cXWj9kz/9MHHroaP8WFVRye
wjUwBf8sNs5MyQiZ73aI++RzJLMMEhsTAdUrQP7JHSdNnVPOTIdGNyAQU2eEJgLE
msEnA2yCwwNKP9zjWVpB6PSQ148nH51Dp7dAfD9d4PZEBI9hFskUNAFvbVHL1iU8
pJFpB6h6DZfLgIGWyLXjDTWhFCetiVp4J3MwjDD/tGPsQEYEpHj/kgNk1T03NCHy
Hmyd/ClHRkvOier1iZqYVTMaUIgIOv7cSmexDl6Ui9lGd/no1hrtHi7tIVja3qDs
8RHxUtxyvGNLAp1BKa3Atag+GU+0A4oDR33D/CJeBLOIrd2p+1BUQ+2FZ7vBKrrz
H5hpnnO128iRN3G1+x+3cxXke31gILpsgcBhrTg/QODi1EyzdX+HVXKpTBEcmL68
2hVn5HrCtSd7Au9zNXZYtTZpQg1gD6d0vV994tzcJYaRD7Men152I/OgzK03Zsv4
KfQqTlKqI4DjmRB5vMs383A+azwddvBEhiV253Lo0ltKk7kOryx5Tc6oAzgIatmN
Q1fFv2Cllo6QF1dffgMdEYXJ73Q+KCWSCpfiBsTZENEqufn3NsVCDOLCF/m+myKJ
FHIYdGpeu32fu44+x5b5PdULhqidk8kV7DcJTfn0Ic2D0copO1MjjfWmJZXay/Zx
MA50tLkchNsa4LLaKIUzPM056dj8fpFcmx6LjWpZZohBmeaQtcp9DXgwI1mSfRoc
N1OZVLOlgqeJZBQtNrP3ZBp69zCGME+lGVIDTvDul1/nqpW9HKlqqAN+98UBet2t
L3CCEkMrkCyAqTc/8DF7OrO7vdeA6GA0GsBli5ZV+dHMbEJuOvlpyn62Pb8qEgz5
gAyUPcwbHTJhLFyN/t6gRMWOvP/5qHeCQb8y33ENBMTfDclEDHg7o1/1GD3DsSUr
ONzroFjrbYSHfMEAEWRbyh9ztt5TP0bzK0eKNboJ416c//eCnTSiTTbrDB50f2UY
r5eq6XtIcW2WsMZpU3WXBzRfgIfVA3fOtQjhMlkSeyEgjB1Y46pSKbMd9mViJgiF
6KL+v2n9p10uC7+Os6PDy+sjKoioZc+OnNXT1FMAGrlnmj0OBL8SI/ijNQ6dZNjH
/0nZJaW13gNJsMe0hI1Cqgk06Tn553TOPz37ufUgV1icUB882TBwPvi3UGPbnkpv
TvQEfbUbw5ZCgc22LjlSHGG2P3mscmXM8ESztF9rc3FkfnB8fKVS3uWx+v6HwdJJ
2fu1lxcX8ui1NLiuFNMZKO7jYkLFW4aQtSnyxGoEHeYLWKk+iJMbNM+GMM8xKYwL
uR93ywNYaN/i3Y4xgUEymq8eYZ39w7mcUn2IaK4ZfhPAlzWIzv7p0dWF8d6hTgX8
84eJ8ImHm2Mpdi8IauobO59QzydQMmqL/IEBjKn3ywehsZOtZxF27fmxdhvhjYdl
qJnbmlJOYX3cC5noPHLhqS2EI7zY2qdSPwfSkYPcTLbvUbEDohVU/kXMeNqqTRUt
YgyL8gKf/U4R8BPNLUESciLqnrLiHRuDHgM5HjIbabDSvIyThEIrJfnt+7sGwOjF
A/DoKcw7xhYr1xMiVCT/JUL0N5etGt6AAupS0a9b4KGp/57cgie4ZqOYYzAbLcXS
tQpK5cIhEmwnIkZjiuUzCmbcCvZ1tM5a+zHWm2D9JLnQLYSTVxuG3zogXLoTcyMW
xrnt0amnRdlNBBIFvIarqkR0FXKf+hIcD+h2yOi/kzorqTwYdq+RBVxKri748QaG
gnqVjN9R8NXZgwm/5IjdGjZnDPRCNjvOL/8moY3oe8ztFKXcIJt+4r0ZVcJfC7Ax
s7R66tccRclJVXBeGnS+KsEWB6r0SjvyPXVmGoPrhuk7Eg/iWHPVsEGrnrenokHm
u6IAtvbd7RdF3XApzZbcD40zRyLID4Gnv6ncRRB4wpyq2sKLKPKGMg56DnuJ86yg
GXLeXoYqtBAv+W6d6Dhuk+o+fgFO367csLqn3W7OXeyV/xkJLc1GK4TP32EeJo9B
t5FNG4C6rqPnIzOfU1m+XIM86A8FpZlZ+bF+fWtaoUwbGyorI/mvnKa4JpJZ+COa
Q0JEA6cnyCaC1YgPF/YpJiQ9QJrUIOxz/Y8hCnLSQm80AUwBUqm7/ompF+hHQwI5
2I/Ux4PTyNcTBfqrHw8iBpR33Efi4zQOzZXQPnNUHq+wr+WC83bjQI+0nXDlp7PK
CDEOSAIdeDRIUJtZx0F39c4aj+TvyQpS8zo6Zq9GSWs8h98WTwvHvPTO5ZcM7XUX
k0kmwZoPphGDxtHJCdM9SXiSihlwwXICaxJWCH98ZgIffjP/jBoa+JzJkrNqc2Wp
Fld3TCKwsz222OGdCvr2H5MW8uXF+FM89kgTGnNWek/RGOmQA6ZJSU/vWBJVKoEc
d5dSF08lvTc1tBvkKW9VNBLzaoHz9KweCCA1ksfUYSOu2ry80mRjjjgrUsJJpy+8
FPeo0vlsMd0URxCa9reTc60peKtmKOhaasLnvM3tGeqhLSGQ18Chgy4Ddefs5Itp
EIbpGzzRzKM1jB+H/hPJimHJb8CJHI9233giVAfDppUE9Js/fhi20e06w5BCH5Lv
R4cfO03CSYpmaq56Tg4KYQ2o9Dk0ZIEidSu7Ni3ILDe9W2Qt/GAvLzip27mClDgD
zzxK7i44vHvDMuq7q/aX2sKBuIjI84ZBe89iAM2o3xEibZbvhM7Ql5DTqQvwnjPI
OdTPr/83wcDfGnL+7nY23IpmgsYlqMCGuJ2Mvt8Lqc95qd/jCINPM+WD8heToHBI
T9ubolZF93nSHed5f8JCGvd+juGtJxulZ66+HmeRN9gzL1+JWPerYG5Nhzk9AaSq
yvvXUpMT0VGlLmc9UQZ9OLpY1LjfElLOezkUHNosdwaPY4nK/YNIgLWZe4rJ2Xof
Zl1UDLcpZ1FJe5drVQGfEUvHigWvItYIZS5YpJSWKjRovlT/DPsZ0zytHOzzBGxB
ZrjaIYK5aFd5hbmPwb9r7SdoszgFpv1qmK1OvShbdwyoLWHojpQaypFbKoQ03XIj
gytjQiLIPA7uzU43jeHQf6VMHT0zaCIPR1/zammXW5+jtR92wUZn/HsUI3GeshlT
AaHzlwY+FvHqts6v5Aon3G1trkWWrMKUVWI82UAgOIfO5IOBbeNmzu8CZg1zscaK
5CeqFAj0nFL5da1lPrzkmRcuaM7kC7uuFuY8zxQnZVFOT3i02TbBdudHSOhtyfqO
6/vR0zsMsFANufbyZXg4qXg4pYLUxfOUYjipDhBNQcenI1h9NMgIYMLdvNZ51Gz8
3OE16di7lHZkgggkKw9PnMJFoW2t4FyN0lpp1tVJSwu3QJYLudtN3U1sS0TivcOC
lMkdpj3e612BawWHcmallIb2SiDKSccmrarRHDGkRuR2531+uMmkqCVYvU1nVo/n
k2qIu/9lOKdTlvqx+E89aZAxY/giVaSm7LTmc2C4hiNQSkdIeYWZhxDcCj/rQ3Pp
9p2yk7o4392BSjrc/E06NuENHXa21troxJKMjOOBzXSeu9L3Nid6ABz+OywEga35
i5/b7zPWew3kZWyb1mLVHBeOtDchtcUREf5ySveAZl6O8kgq4vD6kuJ8SioR85x1
mmXh+mdNvCb+ca4Xn/w0kN70T1N6oHAPIUvX982k8+IeMWLlh1ellksxoPi35vNm
Z5Gg5uBHgEoji/frCL/oJmQukR7CIsXo+64IqIopEobRoFAR4tHzCAPTuS+M3y9u
FSoFoW/dHN9KuLVkSIDbnEwv25uRoxNFdvnjtfICnPT4PKytTlHjKWC9eZcogSI1
2CEWtUynJeDUOtUcbQ4IN3uk8V/mqTGvRf63HDXUawiW82O7yiMdttFiKrYX3Pjn
m1CN5EIt2uQJwFcIUq5xVkG22YZ7AuD6focVMkNCOSybuM+21e7gPy3+4I0Ni7/o
0Tvwh5CivfwPyrebdH0o7yenaWjsHFr55r2Dc5zgu5ZYZYhpAX8Fd2poanr5hJ+5
rhXP6ZnYVRQRxRCw+sPaV/SMTvjRI+tu7DKggWz3AlwqG5d4xe85oNinEZ6Z0D6C
9ZT38RFdX+AoEBB+pRMXU+PWT0sSmPhElVcO+HjQmym1dCj49wJO+P27DmwhT7zz
x50Q/a39oMjuFYCapT7pkC+5Xw20Clv+JEYn4Ibk1DVDjZ8VrNHaIzi4PLOs5GA2
qHaPeE3kYkKpjYn8pwEHqRgxpD1MntShPUQfeyxWqlihN5G/5yeMC2sCiCJXLJXr
VLQ7HA30xt9fqDqvKgCOKUac1F/PlC0rClD5+dDhXLlL32zaiMz0+UkB/LCIBocW
Bqthyo4sD8BUr/lv36dpOEGSdzR/7JgVAPDOurO7AefGN+QjnDzyczgVED17Vxb5
Rd9CVct8zKVtoS66bogIUa7PQVYwwEp1JEeOcOql/vA5RfDfR7Q11doBx3PNEW3h
D5nWD6iqCq1nFdIXEeAtbpZ3sGr6YsqpfQOk094iTZW41qt/Jrxd8W2fW/CSB4GU
bRMGeNLfMy1MSY3YWpVd20GoBSJcQdD4BKyidiwg7twd375gt0nkB2SnvvwAGmid
wV4JjlemffzEruvJPJhabRCjySV5AGKRSQuQX4nmdBkMTpXf1hYc+FpyuFKG4dmG
f7q8WO67GlBgX2Mx8HYlsUDgveCaKm2XbbmC9jAkjhL5K8ejJt8jPPufaxVdjEse
FGhGQ1aJxBISui5kntXF6m2yimbS7/fvevGuBpOehjVZT8hQeHU2dZIK2JFwEAp8
3Mnpnpc67sgDvk/fcoZSW86STr1t6sVVOW5w1Lv+FbAf1e4EYiw+ph9q5Wk7rfPl
V/XgJWBdH88OOsBsYe7vzNQOXPqbk70LLyLZCRe3f40CHzjiANQKriDgS7EEbhHH
GWyXOOZUVNNPe6AREU6fNPp2mzDm4HNX0fu+89J+imou57ZlpB8U5+xskSilF1+3
jUT0ZOnB+vFsEJ+a65NPMaI/0Qh7Yxd6aXNOAdQzucAg4sX+/v1zbnLteXkhijT3
p1Z10yb/cwMHUxV3FdkkoXCvj/snPAXNqAdmEAnDjo+7VdH+KTJ4zeK+sKoljbfp
xdntgqoxpVVU7uEUJqCsgu4PS+34KRd+Qnbo0SljdQK46/v+rwIkzdvf8tLMTBrS
hkrJiZT29BWTim7wknVwzf1eOunKuiINpBzO426c4/SCQdZOxkm0EKq8m0danppf
TpDsGT9gulEqEW4rx9+dv1mrAIni0BBa1tlg2oMBLH3HnwTdt/MJ8frCJKrSvjGT
LUOS3lEDMY8DvNMw/bm6+XLZK4MWwdXW7V7T40t5QsGn7ktk54lKymEe86GC/eMi
dKRq98dwa9gn6QjIlmuq1l6CYYAvZYsazQfl+2FUWueUlvd5EnbuCQYlhlBj9i0b
zQ39HrzS7PkmVIhE0DdbzcSyDJw5Y4Giv7o0HhWZgquy8inELNO5fJTqJecsBOkb
tFRJcNd+IX1xvLN3UOoQJuNq88ku7R8aHDXrxpiUIUcT4EZlXV6NQguUiEIogiQQ
D1/V8ugD1tBMwCg5NvlUPxDCp6W+71aONkVcmZt9JHJxb3LBdMwUx5dT1H5j+Khd
0vrFw7p+2jh2JNl/BaT5sW7wUDx62ybDumBxfjyP3mT5uifcmfv+dvc32/fqgpaF
Ki7dnpMmbebwM0oFXSqTsbfrDXmH/aLizpBtRFjVdxnbfmMwmR+r//I9dtlQsWLp
afc2XOisGDhluOqFjaEmhBANCEBmzdVUMkil49kIE6JL0mRQ0r2/YFBZdYT8Pg/j
Q2iaGx4WDoiL4xJ1lJnarKC1KU3yYf+fKJ9X+2HquDH9Gl2fUGkI4kw1V0Zk5ula
35MpiLYML3wpS20svZF4+qzjShV45TPTZYstwap4wtZLsYnp00xtUN1S9YuSeSxo
gAczvYbfAhRkUIk/eNYdOm+Bo+EJ4f4Ex1R2CSQLKyzOiBGntZqEw6wjOhZ59pBe
NW5szlKOQZrS6Dp9qDSMLiz2S464TstSeolbg/dCkgsYN+bcdKw/wX4IXy/VU6fA
jZUJTKClouAweU7ybDVWlCSIoljMCCTBSGFrpL1hLA2nNV2H6i52wTio80yy6RNf
wjmpyRWzSWU0s+JDWhoDpFA7DcvepFBGMX9C4aASeGj4swuXKcT+a0PYHej+wpau
T0R1Up8lAdQ+ifI3aAbFg78ukkhmf6FqOpopkoQQsiSo9p5TmvMMgBuqUZiazMZk
LyIZwA0XkrJocrR/wB5mzPETYzlvQabgbKfQjRnxZ9TyOsiAMhnAq3Zp9g3N66Gc
F+LEDxfypof5trcY5bGK+83yXY5upmlZQoIXYMNCUMsRzxwmcNjqf+sr/oKQYJPF
/cVpwrsbE3ZxrjFOhXrmEu8/O9SUw4+HiZLSAxZsfeCEEfmhPxkvEJsGsyTezwad
6wAzGNNJRMdaoGlues/TFK9eJvPSj4s11Upbrm/se2QMux9OGXcTqZdIZFXZI92d
eUTcngr+OGKXhB0D1hDgHDnaPOk2pP+//xsbouKoVdF3G8cCCPNJxeM0KHY1hi5I
uv3kZ2Q3C3Y3+WTDP8jBgigxQNZcOdmRYjP+Soyf/b3CEYxEdpDqID1GUfOcd5Sa
G7usHJ90vn513p9OSMtDiNuplYvWW8bc4SyzjyOdP1PUZLtNOpZk1fMdyFjWNlDH
Py63m/k4guuQIavB+Mxst5Fpeo9YqzLO2sMCwSfbJSBi7Ts5tyt5KojgicbPqy6m
TDJGQq/6ETVhEMF4AtU3cAjDRk1CTdGIrSfeE1O8MjUwvFoFddYOq/5DbQWhRPKM
yf5Tpaw3I6WH3VOaFFc7Pm+b9ybyzYRJ0dPyV/hVod6wIiStwonj+u66OCQaMkTR
3fQunF4otjfXGVajjOikefBj7u/nFg6TQldslcHCsDv+4WmCFUZBQY988Xqx6woY
nNddzd/vVhs5ZIu1/pknO4RR2C/vZU6DSA+7nTnqKPhAlXTRNLbgr5ARnAUh6gqU
ak9crHa+JVJZQ7nS9vf/C2Q6WLp6ZnU0MCRtrRkK9Mdc0pZ5f3SlkCely6F+/6zV
EkZgHvenLyrbR+YDrxA7fWjzMpL9IOGBeCiiuWpinoKHT7b+z7H0ZYdhLAtlWWpO
zUEr6a/fNTfY8A2ERCLSTNcxHnaPheFZb4oLMChWopsmyu+dbY0SBKvLllIA3158
NMiKHD/cHVsGj2HmCoAKmcv4oPfEtPOqduhOeZx5AcllKf+ZIC2g0/pRTdm9nnIJ
hJM/0/wlwgrXtebkwo2/KE87uWg/fi/F7R9NBgd5T1IjtRHwx6ji2lSiLCibn98b
hduTyc2zi0ZQSszVO/rIsH2QJnDCWSP1p4wC9IAJxd63805FcBePYyYifFzOGLB4
9ZVELju9xuYcI5Ve5rqaGr8mMrQMcBrtf5CFEk5PpzyE1sMfr9olptBGeEAxbjPE
rih8uZAzr0mH0pHGuTuSk/OjzRBKBsfkfXSAxQ6P8IsCGITuvyDd1ldv0C9MI2E2
1Sy5hXFQpfGfaNj8obCpJrjeHA9dyRJchYq9NLKUkUGvGeXwXpcMY1AoVOBdwvos
t9Wytvo/uLo5uGoXgINHEgUzQAOFOQsPE/Mh9NqjUQCILNVVKowGtcXXf2aysXYf
e2CimoCGEjb9JU1P2dYkUthFAZFKlEHuodovRhNlkQBV0xiyKNmJThORAic0JWJZ
UsGNnLbohs0NBnVQpoBReih1Oj1NzLG1zf0p3Vti7OWkVR1z/Bj4BR6qtTmrevjS
8/DuaHXKIy3bxFBAHPpNhLKx8bi5nB6gf8WB6mXd1V+NuA3d7Jq8tCLr1iXru6Nd
hwNX2vx/Ia70r0g0ErOky938eCZBP8EtKq0S17AX0Ei+PO803mpfKazFzx7JDLOm
pOokuZOcIeaLupmcCRyJ0TWQXcRaYSAjScdWRsWXmuiXpLxzBGKmd0j/sHfq7E+g
s3yyHApEii9riHM56bKWNQRMGwhVY4PIMSBSt1dE7+v2xmppkqCIgJpS8iYbE9lF
P6aheBeRyp7WR4tg4fLMUtTXKvonqHaKPHSODwy/+UAhYUY4UuJgWM0GS3oLyfKw
FaXYlaI/O7++HFEDjQarYmx0Z1S2xRwMkOpZvM/0GjWkj5ZCUa+2+u8RKGkTlX0I
4j1fOXgNhNGv1YK/NLfUV0oHl/o1MfFA7IcaA0i0/RVhene7bKr7S8/n6Ofq4K6f
/hnLi6NIyRqQVNHCAnrbUrgfdFmXTEt1hCGDTXEPkplksOIfoc4Cl5011iZxmrpL
GTLwc6aIbpAUn5Cl2VfF23YLrZSHWnjWa2rf0xfZeA1H730HFWNTTFAvgNyJElsQ
EGL/9iV1OidTSYy5EPbbL0gd/bmNDQGLj6xlXgocZuPso4XXoTBysltheVxFpnY5
/CXpvIaxEpxSLV8CQ5lq4wJxB52Hz1+1LTSXfwf6fizOAnvCgetj5KNnr689lwXi
VWSCM1bCSDQcojtsnE5IV1xHcYEZq1S+mSu+rv3FD21W3Uauihx8SH5P0dMg3lT3
XgQ6Kal+/tRUVrbvSCfY4hU8NH21uvnAg1BA8J3/QBFVgmLO4w9dyi6rk1aoQTOE
ios2BTT9JOTvSk/h7QPmxiZY13yysdI1NWJ5YyXZQ9MB21sR6T+X9Wb+kab2xTe/
m48TmJA+iW4mX42/VfwEi3SKvO5qzjAaswcI8rmy2XiJCAl+ukp2XT3IeLqu+Jva
loivbVbZP2QSKFYsk+ysG7pKIaU0GOCnPwPbiwT2+BC4rWl521d3Ylo+Ew3TmcZo
EkPuma8Tiij99HG4GJhqSCI0edBTyrYYs5dfLsDjLANUJfbURfwkl7GBaOv73901
Jo8fNq5lHIMwQ+Scx9ag0rFqeciavrA88qaoagp5fTAoCtUSsgM4s5oVzpA9dsHJ
UgkzaMo1qYnJI2YhXQwlnPlIc0wOvLRr2g0vovGtcuHriIPBdaAJLpOqebcXyNCb
s6QEDTviHww2OAOHs2SPfx87GNBpxaeHBd9V6eUYFGUcCxuQ1Mcjwalnx2wOQS8f
KYGci4n7Ug2b8UoD8mBht7WWFuoj9i04QXEUjSfB5TC25+lhFaZT21F4qUpxid4Z
YuRi7ra3DGtIonx3GQHypeU0I24/XC0AYC3tnIz/nP1adRIbZ6Rys/Iyv0LOoEhB
K9WMrDujppkd9oZ4UieNz33pM0gsYqXXdbvgX1ypQ0X/qDIRacHFNjq6k1Szmmxu
FJfcANvts2sJSspE3xNNLcFl9mIapiB+6iiACcSq5QP/WALFabfRWNhbBB9vKU6P
7y6gaqvmZeZqNsxJGW6ecJ2Y8gPLPK88/0tBuvfUgr97phqDYyzVs3MupGK2CVS/
KDGJswXdOqAGtoeNpWD/1/Gi3/G3rCx6g4E5IZN+lZEYH108QYbq94cXzwlrdqUX
J7n3KbjhcHTUNveeFjAX84LyYSt72Bj2Ec+iwYqzTCaVcaUk3/vIrg8OIrOH+Zc8
B2HIGYBoh5fyOoyizCfO3h069oDBPk99OIIM50v5FwFonJH+X+vnBk0iobBPmeA7
jaO6H2RfZXMz5R4UnGH1RVbxdMmI0ho7mtR7rKr9WfrHP/H5rLCBsLyRPnHJwNnk
47GueokljUMy+qzx6jCtCVooRuX1Er180kjK0w1+Ewy+zlUG665fPUJnscerkQzI
d3EUAk+75KmNy9xegusHc4360Xefzp0D3AXcco5PsYhN+dwcQGbvJ1ENoPnK8G8x
qofIWTy3k+STdFvmXxhEt89PZOT3w5qRvnYKSsj1A4V5RzMgLenTtSy3yg9o7J+D
PyaT0iF7I306wopiwy3kUsamwjUDc1/i11CDH8erXpK5SvdRMQR3qK+IXTavZWTF
N/ja7BefItEudGFBRNpVnkldG5JtKd9Qx0DNJsEiJeQyr3DlwPAZ7X42z2kHiNVk
D9Gg9krXr+re2mt4ZjNEsxd2cc9tdFcheT88txdZCIaA8amy3GyjEaiJrHg/UFuJ
oddBDFoZy/n03NJeORnGKXnmWhckJ2vJJC6kKqUUNeF6X/wBmH60mh0I25h///0q
dOxEaWCD2rDNZTqAWSjP0zLFIUv0ys84iiPtm1UAOoBegcmp84qwFHz6t/ycawrl
7p5qbLVzBbrIxImEex8UO4kTrLPpdc2X4V4lvLncBhF9Ey2lNFrmfuhTqK8yQ0X0
hg1c/kNHrRq4YA2KL9M3vH7ctK6dI9TV+/xReM65bXYSgZGUomcUXFb7+mrcW1bu
x2ySzxV+vTnG23Fl7bPSUkxxWEb2IoQaUkpWlitjjqQ1eYRnsqMsB1DFJ8pK7H/3
klwybJ0EBejhyoNeFr3qG5pMuihAJlSwXXgkiWXv8GnJiaOmj93h8yMfyXDXteiN
+1IB/o0WmS43JZxgA6gGvbVibWyZcpWoSmHpPiFfCGiLk19b3YYOpYhF9S2JMg+f
RVT9+zR5GnfFfPEHfFpjI0SxpGhQfMR/7J/agLtaB6l0XWBIzYl6wAcsB/5RcBBK
P2yOP2Y3VlTi1OieDDwuVRZNcDjINdrCghMyCvTHrcJvO3aCzaGXKYqyVLqWE3Xl
WabJV8D+IB26AQiBlkPPXnYshTDqhRtSqsJswj02CCaPJAHV8BnqpqJJKvt/OoLn
Tb7lPs7Hw7mU0C5dYARrnLjUOKE9c2AmIcCsb15ubOjbi4uZ/CCwUhAfY8g9F1Uh
wcSWIeGVMdYq6UPucInEVqcGf44IANxnO8pz75Py2MN6ThJhBKrT+lU5PEqPqosh
/tjoamSnU0J4w7kw5qhihs5A1EtGKp4fFRHBjmII0uSUONJiie2Vi3vINe7xM8Hp
Gnd0sKPA9k0JpqrHeiIqmRldLRJXZdQ1eoxYSWN6P/jbC3FeMOsqSMepkASRGKO5
i9oymVgjSbhkwToa9oLkT8dAwqwW7vQhaHRUF/tTMmVnNmUO5/93osjAnlbjkx5q
OFTCd9Wl5UhbbGCy18dggKcEtMwjIYXhxRfge5oMx0e+WLwADIquVQLLyw/tBR8S
EBJCU0TVHSW2w00dhXwz+hUjeQ+Qrf0wMIgdBSFaaKW1d153xsM35lPaDOQKQXB0
nxRuOZnP0+18w++XQBnT5l0B+9+GZejjJ+a7MpbriJ9H6qRJdGq/QuhWYE7ERyBv
blvchAYZp+8SKVpquVgtqdqSo0dkSEpWEwRYml8xD68CmuYl0fUCHpBX9tPkZGVH
Ir/twAg5i7gJseJqpASjDNTz+Iyuqfo/+FKpp9aU1BEM8ttwKSF+/Nm7O2U6sKka
5HelpboPnRPKmA/7IF30HYs+aZnMCS1xpjhkP94Hw42pwZbgLYbdH+HraeTAlwc5
BFmBOPCbUQizkaYkGyeVBamMZZr/dtWk8vWh1M7dMPtbQqhsAE1y3+mty4eQNifd
6hvNzPD3y9gMWx3AWSOOmXnQ11l1znfmzZvsyTTmejyhZJugT8PjxBGFUA8z02Tt
En6RLMNCLcsNW4a5ikh5ytsmaT4cX/S/cPE2AQL/4vIjz6jVNZq+v+e13ODXp+Vg
dHKoVf1JxA2TH3LW/BwZEyTSBhwRjdBVhk9hhEC4Vg5w3NXGG9L4UxIBwqko/amV
ryif9gq+QC7KCuJ2CehCk84N2DMxQrmZLfojBwVgOGc6SO/6gROlh+VxJBR9CFi0
Ks2VkrwNJIXdHtwBe4D2P8g+OrTcmNE+eKEO46N/x0/b+AEPc1CBDgB3QMyVPsIU
x0zU1iCq5SdVMfJIpbIoB1ItnWMbIZ7Jahq60QHFOkNMoBQ7TUzBGZbbTlsp2WG6
6YSIRZkOq5snGM34sTZg9HZnqYYkvz7qPUYlAi/WNUHDpKduhVsQ9HRqH4nY/Z5j
VaeNdBce12FSxJlB/WjeY/l0XX0/PXpq82QeS3Z356bE4diPVmW/fbVuFWiMv3SU
7Gv6p7U0Ok56e+YOHbxfNkr7di0woebIv81xZk2bsukACWkSJL1mFICOJ8hGHRvx
qgoXdak/H43lVDZAKiitjGHXIscCCRDrtXt4w73Mxd3EVqQYbkwHWnbh8OEwnM81
3P6D1f8Hs5N6teMB+ptLK34t25yAVdLLveFkYl4IGa6h9cpqLJFqF94/0g3QhWqZ
q75e2ixJOlWq0/cQvtFBDl7mRyoQ+9tSI2FfG+m7g74nGcvXhC7GE9/Z9XmElyby
M2XQOf8agcbupRcod8BrtFg3vUBLFj4836pfGiUQIpSegBQQnvJMy869besLIkgb
3Fgq+hYtYC3JN4tZP2Kv0PcIl5mEToJLr0kQSlVCFF7INaiYN7vfhHUrqnjNIvuD
kXX8Fdcr4CuS7mzysGkq3jSbsED9dsjrCk9JajwKkM2oW6PsvvkBFjHIN7pQ3ash
BgKDkkF1tM4LY2j7/1ft9p2YD4ij5aAbLe9q6E6GIAulcdpgij+TAsuidHBtCcLb
71qBV5ASX2edVIRU5Fpivm+aKNKmP++XV95ep1ZwcQGlxbvWfjuQZtWYAUWBSIKm
iVW5YNNqp4USwlp2yf+9KJWEbjX84IMmw61UPN5NDxCKO15+yUYhqf++pnIb14LL
c4qifehWuYnHi90q2XjPMosEdZnBzPH5dC32j+BS+f3qG+IXeHkhxyccu+hxd33r
xVx23GuaWIMe3uKTuOaaz5i61UCVNqfZX/NzVOp9nfEWa1Yjgp/fYaeEK1BiQDeh
UyUyE863kfLC2Hq66Pt/UaINpw9B+PGu+/SNnh5ZwwbHPUNPVKK0IZIAqoMcemPH
g9NH2bSmee5TNT9jm5HlW+lucfsqY6sZujqTg/NgPs7DRxEul5JUP2CN+w3rjVeO
huN1igILgTxe5dnr5pnYO7rVvNLRDdmeFsv5GlS5uia5mDvz53U2rCqHFIoCi/0A
91+znKA5/cVXKh2RO9uQ1geVkEoNUCA1ZvquEoZskSjrEPWucXkFxAFYEhTc13rU
o67K2Gpu4Fwe3Oh1rpeIYa2wGVYKMSQw/Z51RDruxYurJSi41FTxpoe36Gsci3CC
TR4m7ISI4WNfTVDTK6kH4fszuqekk2H4YSqlv5iropN1YnTZqFeWNX9eA4EHbH3e
yg6yWAHYMxAKhk1tTrR6HxkychNMO3oNz01rAH2YiLu0H82yARHFmLyqK9UFT7/o
5CYMnFZAArXA7wPpb9Qxzu/gHkNJwnJf9C81256+JXZSrHyoUqNZluB2abxXjtPL
yhYqxDyjNgbcdT/Y0K+2igIE12kSj3fw05Wc8mXrEZQM4wqa7ywAKEEtNGIPNJ77
oa63f5Q6JqYg4bvEwY9RyB4CZ7RECwNVr+oigi/NXar9z24q+4jDpVqJ9FLZuDG0
+gUFrC6xjr0k0PXaRhWjz45BzaIM1+ubKYMKrVUobC+OgUM+P7glUvp2l9bBCzRw
T7fGFhTwVWPi75jwyrvg0AMz4ERhxqZumHVsFofY+p5zKQuhp6v5FqmUcoZEEXGZ
v3kmIIAYwRmCptkWkadMw1Df0gxuu0qJd9LmBcUjXRSGr0t7sBedVce46dvAG3PT
bNVogD4R0WTA+HqTg29ILJOs9C3272wwLfg5z9X2BZ/4Yss9B1lpItl4yEjUoqv8
Zq/8ajHag9D7bfVJxyhzazjeUP/pYdztRKb3fiBXL1amiidLmbryr+W37kLwxZGW
SiTtWo/wHsTkaG2qA7VFJn6o584HNfq+x/7LHfsSPcPpD0oLvQtzVcBBfgFNJgIx
yov15C+5CqmoYCtRwEhFzHmvKzo7QAQ2Ne6OceuhnDLudJa/asSb/iRgcUxrwD+z
eQ2AGObORzh+incPOIfTDP5/csZscn/aCKOckwSuufSAjol5O/+79svjBzPGOKj2
88c0VKbrNpVENjhRMIEZeQhSdN/s21sp7mlG5IeAzt35KIfrh7u53Fp9eyz4DNDT
Ck4nngCT6QZDNJFrG6OZ8z1LWv6D2z05xuMd8bG0DKJRnVZdiICKsOAaKm4+ZbBQ
YiWrWgWDzteV0vqN1qadAAWLWT3Lg/ZQLexeXNGcgIhuz++tLX5lljMSvP42kp1X
tn0pI3S4+dd0mdJmSgu1uHhANGm5mbwCQn/6eis8zsHE1IAfImtracWuENPRvcOd
DoMvuGflydRYWNkMUMSI/UApZ8qXG+5ijjATDs5YFkisfPqNAjOcrfSnNWI801+w
QpJ4GtVXCvyhRzFiKUiHQIeUFgj+Wav8OldfMApoUiH5dtTpEM46CwiNooLADF2y
E5plqDatW0UNyKRBu9wd20eT5yiE2OXaz1rcwBomTCAsRYQLSpDB+YFLYNlr9WLf
MMXKkhGrfJ6ydK7FjExm3T6gGTUu2j8tLvhe3Fgj2mbJb0842cZexxxiqlvVwU8C
qBbHCeBZUTRp3Q8dKM7CwWXBVJsSkrfxUlx4piWCqjppxg0RQpLnp2WzsBkdCbgV
FsWEVtK8J/rrfWjqI/chBSldMRKggIpLmqdIOJvITDI4/xeR3ITXg5ui52OzIf7X
29innbyColI5JJGCDc1SDtttGnHBCIuTx/fVZWySiSbXqGbp1V3V0PvFQ98wW23U
Uy+SVePmLis2PqP0alRy5+/Ay0fLp6qcd5gKDIqp98fn0pAYDOKL0B/P8wACQcf9
0CHScTkj96KhnxnBQyCaVLqGkGn29xXJzwzeOYUfsS2V9qEeuG/n2Ts1oGnBWirw
Iqw3lu9vIoR/gkB3Rzsscf678ZQxGWnp7qF+S3nyFRvqIU7QDw4pQDMeoGtt/zH/
K1HbExGNkYmgDW0lzu3HQHXdFfc2X+KoIi+oglyVB0CTpDZWEKeNIJyq5NodHepz
TeccRsDSw8yjRHYJT9ZNDXu+AQ7pf5yY5I2YjX7pgspmcA62LPDwss4lp5WH2ywk
lE27mXTOy1pQpPLXkaWlsM5zVUGp5BrfV/BdxHpVvVexCxVojBQAT1lRsbHXWVo5
fS2cdSNJDrHrkArA8KM/2ygpLRWlAPhu5bHPNaJ/F3CmEzgkX+DzZ2gxKUYuGGXa
Gwx1O/ht2YNocuyOvqMazOXw0xeuR9QP6gq2YUDL9PRpzJapnBUVQSjUV//G0oLd
ddTGs/noB4elC+saFwhyJTW47mnGzrZN0JF/m6cnYbAZE3KMFoZcDWu9F++NHkU1
mqRM4gV+Zatpv0kefRGDp47+zEzkLe5b7bRrehXyo+iWc2Bns7OnjrVsfiVsKCHR
wfMjGRDe0UnxhwHZh3E/zdjr3cPljxs4pEcHbpzPrxs3JzF95qABJxhV2D8lbPQ0
//4j3G+AQ4mZJECNSRDuAk08JDwbs3mxlwcwwNbyaRav6dGr9E8RMgPfVOpUd/HI
3KA1/AFYmJ2C1L3urml5c9cdmenqyPPV8DUrdzuziHr1MwvrePY1q6q8bfNzK69y
/IhJk0w/7FDo2lDQHrZLaxAvWcH8DAQKveMTs12RhSNH5PUUertGcFJ6/kdiFbBd
HGHTVDeAR7FHgAtiAGEDCe8nFmiyXmqX8h8VvtccgBherIx8POA6yqfaSUMu27Jn
rGpu2Db1gGuTKK5/rH7zUo46zvM26OISZkq1t4ZScC3k4qAQNp7g8jc7zOYOYk3Q
GkoCtPjZNGPnUh6lTBJSg76Gtlm2bFlXtOi3V21frBIthyp1+H2XdHS8WnSiHqlh
BZuc+9ImpjMAnCLZN7I69ep+c9ZRRpTaD7pax3J+GjU3Sqrdr7Kawd4idK+Vq9cC
p2JSruioHoIOqmvAlfXg/KBFtldg8G2/uSLajcDkJd1/XYBIewav9Cmqs0/khNFG
c+TzJZLM9XZ6/JXpJabfL9RMnj/JOr/biiQcALJ1RFoCPyOyYqaq7cIMAYrhEEbV
IWrA4iHOZ1bbJ1M/hs/RT92tZ7vt0kVkRC/08jX6rkBiLBkduPxAowZpFSyyNaZZ
Ih8oa2phKIxklieE2UzjQfTmeHb/hvrBawtbCj/0z6CLJu1ArCxmEKFk558dR8zg
0YTpJ8SYa5yvbd1TqrfRZJe0WXmOeI9kiXLMTNbxed28XZIelOGZ3lpBEjBDkh0+
jzZ9PFXzsuLslvckXEK0enrwd1tm/p0k+C0M7/29RIjl4X6bsto1DJz+qTla3yLD
+2et03sT+7h6clz5PsjCyx75cVe1sZvRgkoCMvrLfy+VUj+mbpaEn9sFOJy+BphT
yIrf757j3uYDWbNaG9YRdpgkksXpCR8tSXDjgD+9zCn9efLbh7zwqm4QRnANuHTT
2iETDRoeu0f+6snkpOpvl9enZ9WIdn5Guubj7KYeL0acs7kWjD1jrBfQM1Qg2jbl
zIExPhx9siCAYA0eWUlv3y+XOCWbnyZ+O808pFgRWIBM5uPlNOEkMYXnyJhyiHOB
Abo2vKLL8j8e26G9vm9+BYupTNIXdgkd88qNadTkMvg7KR+ihUo4tauAUPpyYt8/
TZykjPbEqqLdE0EvPihBqkHANkrfPtZRk2tW3ymfmQAZFGAfsqVV3Lyoqfs0nqzn
SuZdbBQfwBJFyK59NyILEdZWX5drLQqvRrEBVsAx6HLJmo3XZVLN1s5JTFrOjNVL
cMgu7wAWzfM7E+eZQ3LZ82QGxF6yTGNOROxozFPTXeq0lkz9DMZXf2Hhf3VBg5PU
TDIE/0YPG0fj5Wkkvg5NT7NA17KZuhQjcw6X5An4vF3ulwj2GHj499WcWbgYCjI+
DRL5Tgc1RKO1DrSp7/5usivWPt0Yc/uyuYUcQh8orPT/g8wOecnJ5vKgroZe1HNC
Utl1g2vOdj+Ia9nzEHfh5PMj/xmYBiE7Qv6969cHBr+gTBYZJTEvAgOOH+KIiHqj
QKjdE8vV4aV71PA4lLHbsH9BpXIjHWI/yXjFxJa64V8iRPXzpMxAYrKJv/wCVHvE
QQedNVGfwINaeO2IXbJL+vORofLtTm8++kXEvQKDnLBMwI3K4+hvWHYJW1AF8XoU
7XdUvv0IInXeTn49zrRzdIe66O/ihysQOJ4rCDnfT6ZAqqbeQIBf6sHdM/al9UA0
PF1+U/RQ5TKQ0oG+fAK9HmbfPJ3kKnD7aRgOz9zkOiHAryX2/vEehKXziuCR1BOn
v0YLJyjJvFrvITUwZRXN+fjnPc9D9UAR7bA+5l1T8RBtkctdE1ck/Xg2paplKn53
XDOHwGD+XgzT+MOGbERu4yaod9rRX3AIbZXP10TDfR9G8QPnHoy7MDT3p55yHzRD
BXldSYT0ikikr0BbuzVix0si4oMkNH/bNCKKWm5YYVSnPp/rmI2SCwWZBLdmGeSi
lrVNBsePnKrHDzFw+zgm1dw8SFcfW1YA5uKq9oETCDWn5XOIBa2LtIpWUgNAlXa7
4m9iDfntAt8dYOy/Dn0pkSlhjHuOOWs0eGrMWXXyREeP2tZdVQVWHj7vpzZ4DpBe
1oTN1Z1Ptle4+bvWqaLMtGq/ac5OadcDhCECNMDY0RLnwL47jlM+sw5+lcmHALgv
vGGv5WabaEqmmDr4gPQmwFmvD3YMqHEWVzBDWN+s66xSPVNKq8vpwMcrrzDK4QIw
LdzFvp3qW+MMfdDJAxgOqhopjl2i7OwJVLZT12l0G9v8rSf17erfvWCyZlpywdnv
7CyW5774wh5RRZ+8f4WZJkXbZBaIJQNF9cxVyLVIJ3yYHit5T3ejl7uV2ZkHDrxm
JtqnotbdFFFwRxSgK0jEtuHfFlDS+4V+zWvxjJHI+yuHrV1y+9M7OcQlC7ItsDki
j212Sfz849xVwbQbWayKra7CBrJXnG2G+08StvU0iTDuQ2NHHlN+ZbWaf1jfvDz8
XIoaZumXwWi7GZJmgl1ASg2F/PaoQIN5Jx4RD4P4/aJ3kE0fCk49BKlUw0+RsRbx
MHGNvPwE0cC6Hn1j/PIWEmQIuZG9m7HhYiQfC8qzBOObIwSvOkV0wiLYFxKp1IWo
hsF/3h0x/5tN8kcGyQbvvuukl/0mc55I3UcnCKLpj1aptYMBCEZfKu+vfcRM+azn
x2eLrAetjkE6E61CDLFrP02zNoThXmaEqAQEoH2rpVoKWNP0RzV8V2c2o6HFut0L
QquZVaCH9Y4vWocOktLww/X4lohoAXp+8DepVTk/7g+iM51+jzAJibQFBtIDUvAB
i7YBm8hpZASYPLtFt0CeBn0mR/NRglqy7v+KJQ8z8IwDCFepy4/8tbKRNhuD1eyR
+58jgXjTTEHg+l5auzsurRjv6IkCSP9MeK4CQ9NVFi0=
`protect END_PROTECTED
