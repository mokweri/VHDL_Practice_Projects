`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
838hoaYdukTXbvY5Uo8dQuKvYx1VNmS90OFGnOM2filhLk2XNzpI8Np7AUS2kCM6
Cqg6/RLuNcA2rRNJ4ADfBdW/hZgWGmm5RHcIkb5sOM2DjFNdMTNWtIXDzYzqI+XE
Bit5OR4YM9/ZHUHVexDAPud99kLeZDKG82+d5h8fhyzB4fpAKe1OIw4GA/C7tWDn
A1RbYbE/9caTMNcbFd5KUHXHuJUW7w7FkB/A6eqnEGRY/9YFFvax/GaD1EC5XXrY
ayTHpCGgw6HdqOZGkysVelbdy4u1zWfQ088/TyAfB/lTB/Vn1JIMYExrCvo/kqax
5VrGXDaaU6VPFIekgGI2CK7S3Fv2n/a4jtphh4LoBIH034kwYGydkiDc8ciAqb09
sHrLTmu+5xPfSn0/a6SZwoodDFmOY8XRjRQBcIHHcdQOhOxokYEAiYSYxkBwo+UC
KDenbwdLW1y/JfuyI1gxoASpHqJXp6WQJoAKFiO2Fzh0AlOYDg4YxJly7AEbYmNM
09d1Qti1my2rr9tKEaRDMo/+3DxJVpEoy1CJA4/WdPAcVi4JUGAgvdVcagk81Ou5
BhIG809Fxcc3y3HIzDDmLFpLdYN8b0JWuUcJkhKmpkCTM2/q+UEfjhfCAJ3csFA+
cFGLT1xUp5b5skiYM95D3H6RJ2W14R8A8RF/k0y/5KD1A+jJaYZS/WKnBje7Lv9e
NPnTK1dO76d/XTkTjF2fh6dv8a6Cej5svwBbIwz+h4cii1kTkzvrNEDYP1Dd+dTR
qRt3/GWrW2dXghvPQU2xBo0JxMgSiW8G3PCbwGSpZUu73QszdYY8wVsbBI4NpZoL
/NxyMIrIRwEwIsKL0abQ+E5UJSKi/NALEH2OJX9Q264S0S3nDSFTQ7mM7NHkXbVu
PrwdlhN27BqZenPyUvlCVdsaQkp4mVWWq5BdtSYwD2Kxq5Qv56SjAUYdN1krruZf
nWBjnQn3qAQfzGZjZ4bARQRpnLuLFq5fbhJ/4Fa0K9bUp8rtOyfjK4z/u+7rRyzY
fuF6e0MZV/tFlAdD7k/N7+5GQ/tRZzSJdaEF2AxF9MURRO1nI/8MIGpCwiRzq7ZT
7MG7HgCf6ns2mVCMau3yeuMCKUHFcoKwJPLfpA8iCdUObTP+RGwKGu4oswQi3Yfy
qr+X3bbhygURCx3yk823gI95Gz4SACD2oxx469KXC/5FNXOhUh7Mv7iHtYGfk+gk
s5/gohqGAMQdPRuNOLF+SyZp19f35L1NN+aV04HZKNA824AJppvZVATz4fCMtJyb
OPEob93cu9ff0NyeTKb9iaPcTq7IWVkIOC+cL5lIwEzMMpfzGY/V5edx58mVc7mW
1htrxw+ODiinno5EXSWQ9DhBZZx+72XukxOGvtzxDlkrqkYZ9i5npCowe3eOZxuu
+cWIH0Qr2cuW3BQUUHh5Jx/J5pN9yFdFsxweUt9QhS7dIKBdLIgsW8bDyreOwat2
AZ63AdeWMJrwBciPm9ZvHi1glfOb2DAGAile0/66kvDh5zieG6JgnFrG6EEIlWp0
QT/du0ykn8INXGwPmGjgUpknOXx5z+/TfdPMFTrkShexJzXWuTTJfp42ygRveoBv
vV4aJ+IrxxZeb1VSNt7KuRpQXZ8gS99o9OnApT0CLqcDukvjGL6xUvlPsIK2suGg
CcVqYZYT/ti1nd3+zIKrXdMo4p/lTb72AAHhhnmqiG55Sxv5Y/Y/h8mQnZhsfj8t
M7Dw+4Y4zMUITgnHR3wqyaPnCduZu2t+K5w9M1NZTGXpWURpPy9QIw2+QWezLxYB
DPzUUfe0VJKTXc8pW9YgZmk9xQ+ObEY8kXCvc71/0BzLhUNgZD67MNZxTN454t2G
4IqoBmSBplDqmIXnesqkYhBb9nagp5BzT0JE7y/aSAcvDtXVma3Xu2ke6R0MRFv+
N+8ilyfo3FrhcZelvFdD385hwXc/ptvzolHxTZ5mvqphbNJPTwOrUSXiWxTTkJBJ
yjhqeGQG7oAEnwIuQNAUAAu949y95WEbGt9Antd4kNCTArqNFMCuQPbb6POiG1jN
jyAzXtvpHPiAzsLBnX2+Z1PGEiZuzlfDkdEVQ3W3Qn//iZMEO//00uRdGaUQBxsB
i9YK29nxV7/sZ1iQ2J4JDOxs44dThZU2g2wN/l42MO2KIiwKioKhe9/jFwsmkF+Y
L1+iCZEKmL2JMuKul9dbI1xpMz+QKehYq/W/GUrL2WgSB30B5PKdLdaqCMzyBXhw
AvUDcrmVocTKmn+wlDfYgA0vjf9tTmaZP+90i0/tiFRv0Wu9PFyoqz8hy+HBWxJp
cpau1bYzNY4bU1XvpIqQAdvzy308D7pFkh2J5q9NIDXUMnCyrQfBpfG4GOAz0dsk
tNXn8kIPhiuVMR/zk/EHwG8r4YyQDKlQdMkPoGBH+YZ014iTCH23nTPPMQ5/DFnx
E87FJtfjo+PnkCkJ0r6OXulrwQmndGQJnuEwFRyGNDtN8VlquqR973JvpZp2V2Pj
umsn8+QGy8H9IHw4F2KjbK7DXoqvqcoG6H7XhtH793sOoPZ+J1xwgMyeN74IB74I
mICErSlyChb9ihy//tSHVf8OqseI/JayzWYEGQEQf9KsYQcWECY/5zrFG6Zg9XrK
0W37cp+1WkIaMz1JFcN5iiPkjdxkI0nLpW6uYXtue/Yv/lT3nmUG1wpk+DPX0Jwr
DWw/k4KRrhm78xjlhAq5aVbt/88UnswYjDlYTJ6C9UMsfI4ReKYxWN20I5pVPg7c
1Qsy5Cw2gQ1v0bIu5kpfT7Xw5mKJczZKiKbFLFbsmeWOvAQ2ne/KKlk1inw73mSt
WAZsqhTU9MqR6QxNuvEPZAGoQJjHZs8hGexbva7gWAoBUmMWHW1Vfe8ckKTYUmsY
oBcppmH2brkNeRqSIrnEFP8V+xK41IguzTpGmccgSM1ZNRBIv4lZK38WZ+fisgxl
/Ny8pOkvoUxfvmtSdw4o8V5sElYnGiKRV7X+ELaCJ3fwauGXB04E9Fzrag12X9r6
Jrgu51rjHeYlpQMzMeNPJVnDbie9doS7tY4OTHhQZBKVfZeaeuNN5n8wSaBNtBX8
Ff9oqpcp+sNy2jzA7WHvhR8KFtqDUOKgMNmOOKlwoneDg6Cseb+r4/kJyGAMq7zs
bIZom6ayT8Nm5KZS3fFp/pZoQaQXTpaQCmrDZqOYER88d1/68Hu+/3VNVIfNyxde
EwL3I9W9GTVDGb/f5G3DkFTd7Y72E8TMLSIM6r16l6QO9v6dmTKNOILzcCq9urkW
0Vn455bXEtF2K/hUMJzkd58jAULgvg2IvsROkV6uMq107ERL/bYTgr7tnkhgrsOH
M78C0qz5Jhce1pzxvoAaWQCwzDK4e08AgCxpz7RB2iWfJix07dmRaA7AYycQfdaL
bF70kU03LaQa+BI8a+tW/G+R8ov3BWkwG7LVlzkt04RHNFLBbKW82z/tdiMplxD8
YH1lalNFObHCarFsB+9CzcLoqJFw6dViy8MchO01XjXB58WIGYXy62/+/awZ6IxB
JqaLWOR7VKLwgY+bVIevkN61MSB22CQUxMFpdfuuBEvhw7chLRyDSCru9wW362gK
gnhFEi0SZnDymtBvmbD2AFCbubdXYse0VnyK5gCh8PyT8O5QMwLu04LGU/t/nOq+
ABFmGhXvS1vBySLUjjrYrlVR+Vz6SrxSxVHFv06sXZZjaCCx395GLr6ARUmZpRPz
CwMZTZRGIDc6NXSCTm3cjm8+SxBJf0KtrUOx/oIbmjp2rs7/417tklOCxgU7kGoP
FqS+vGR7g7Cf9GFUU+wVnh/oeOu0FAQY3dy23ZBXz1m6IRn5nwsf1/BSVQKfZ5Ka
OOgsaz1eIHMxr8nznGWiTNntYmjSsjkoX8WkoZgSbFg9Qp17+FQktdRTnNeKGEqC
BzGoSFgHkbWG/F5tSefnhoMmtEoh8PFKXlxWZgDPtaby7VdbC2AbF2fI3kam40Up
fr1oSwDoNfntqXD+WvADzGPZR926611R47ylZXgf1Z5q+Z/APivCjp1N4qrNqplm
SP1n/O1Wm1aFadHozyDy9ZV3KrUh5PwclyIcn1PzXu6a5LNJyHgJwovuLURo1Apr
v01Yv2sp+r71XzjVvwrWPYIJHrYDrt9UdyrQVdypCBffUfyYDw9YRcF/GG6UcSpU
xAQWQ7mMgTRg7MKtjgJl8ruPiDizw7iU3g6lgxu4714ME3Y0Kk/H9P1HFVPeqpEo
qm7TNw3N+Rr3LrXaqrAxGPNEgMgmi6ZCp1IQO1TH3FgzSEerIwgYeUeejmnjUxpq
5jS6OUUpHYf2z5/YazApMTeNbS1E/LcEl9WIElrAiycgueUEaPTMl7WS/o7bx1dt
3ls0Cp+8arULYEfy/flm06Fcbuu1ZmL9LjcsP8BNFcMnqpKlBZvfbxrdqQhggwtD
gv3x0tfpiVohviRcqTr875Ps8pa4Ei32ORyip3g9ruDdARCKf0/c4kR6ExNy+/5g
DFHQaXtsSPIWkQDZvShp+Im6NDg6/H6yB0D3jVldvyGKlL4r1EFkppRDSpgP4JvJ
24Nd3uTNn7KB7IBdm08XLMT84FAk+9pUwYL6dNpZpuaDmYUwSMT6vuywXdtqQLjE
rDjYnbCMYZyS5ymFryONpBtRaEkFPI6A46Y1iL1xT1AVM+EWCBKWzFyounz0Y2WD
5cXMd38loPF2SOQBEtiruriTn8Y4SOEBE042udFvQbByZNAyV1IxWIbjN0tVDJkJ
eidpJpO1Ir516gGXncdekI7Y1tku4qwyaudkOVjIdvoHShCBFx++ltP6HGsrhi3+
5dmQLTmYRWih0N3wiguNoYm0IcVFVpi+pSwNGbxXUz5IGWz5VBlklmPG7EOi4Bvg
W1nwbF6LF8fakisSZGXYU7nq1iGtaJDTjbtG7ziYji369VkI1UVxz3EySd0CLjvP
eJy2hENCmlohy36l7pxg5o80WUmR7dizkbuaHrqnAJGiokZ/Cb4NMIOVCdZrh7sb
DUcqFuL+3pJb97qJn0pLErsPZXY+YI/B4WTQcPqxb9PxtE8pnwLS+W7wcIrxiWWk
b4C0Clek1Q2GKhgAsU/hR+AtKx/X0mBDiGgwdmhX6F0P3vYp3vahfeFj05xLTcqt
P2BJgTCXdf+ZHUTLib6v6eCYG8xSA5KOeXCwdzVWWyw1EWllq/jstSMsUGAfHzA/
sldiEDuSmaWuJzy9fxO5c7m5tv101lTZTPJIyK9g4IgUH+HXD+mtc+1tr4jIcVGU
oBO5AW0jXTijfSG45HGd9hc6//twoP18YzI3XKqJ6kpQNNivju07R3AtPY4hyM/4
1WPU/0HATHjuzV3C2q/rYPv6uw3vdmd0WQC9Ses+xHFx4WuGd1R490bSdw93Qoo8
FFhfe1IF/1GnGtDI2hge5p0jkFDDcOF8IuGkfc0WnYD/gN5Mch630Q89zuqejZ54
RScWIaImKbd9DXCmoS3IF4bw0Qi2HRdcYF1GdCEyxBerGRZUcueLyXFQTggHDMyW
2vBEcZaKrf4TucZzE3fZkJIiiLo2ECNxpCz88kBatlnh6jM9XmchLcDTMRSCxzKz
mL53aUNBwJ0oXFrUrhW+1ypi2uAfcPyG+PRRNpx+JASVaNlIKXxgVC4beJQs5mWE
6lL1WK/mfiS9X0+rUuEyzLklhXiDFVzlhk4+W69gLzEX+xt1ovb1wBRjJmqpz0nN
Z/Y9P240sIbV+1dF/NPXbEj2RbT+wEZNCtZjEgOgGLMLJl5sMnuFHlBw9ntx8eKa
XsXmhrBpn9iHJrsJhlKUgJZfvyheWxFVBK7rc4lNh6Tc7ZmCN64RvbSZZQI1ogus
VxEVshRo36j2BPUPOQzlB0STD4Jq3QfO4/fxL7X9WFkBqsOyiw7FBdvgo1MFfbaM
yRitww+0rEqe3DFHqP8ASpRBssS9R0xDrDoIuWXbwahfbga723x0UtPtgW7mrLqc
thfEwcgqxTVLApV0VkZWuTVP08asobtVeqxrdIy40oryMgMc8w/8AUPgPoZOm+gM
+TIQNtSVxXmgUT7BcsWrSSeUbCd5p65IV+PdRMrzZbz9T727WftNoNp7kRtUFy+q
yPqFw5hsPoOdO2OQBcZLHWCpgqoR5e1y2IzuMzW+DlOEj02DPf6GoJS7BE9BDfVw
Lv3F0lNBPVRGlEitbRPMtAAcI579Uj+xPGkQW/Phw1SNdtSbs5DFOmOyW8kYumw1
AkSeR6/u/4ohdlg/8j8qyrUapt533hoPyb4tP9uW1BSfc+xbr1GLzPrm4PQWchda
K5uE1VysXV+OtPa/ajAJsYhAO4e7+pMqAfeZJjpFzzcwPLXSvrR4IIipT6oPmdE7
ND8GGtFt2RmetZs4c4OHJXSx+Ryj3aiMCHur94TBzinZ6KtjvlxOt7L+jGOwg20O
cuVBJzDqRu4H5mEkEV4FPkV35zXsCSsdA3EPsZX+6tdBoMrWlHeU0jqtQln/yJFH
MBIzw6c8y23aipkojyvPgXhrRzYQKgMd1C8H9sNsNuJPAPBdZFL33Q7Eynoi1Hf+
b2v1iw1xZiRbmX2iQkTTM2La8rkarlTNqsfdJhi8jiOZ7+dkq6LxKoF5mgwNAAns
umK+O7FBtKupLVLw1PAQSUK0rvs2l2gHUT5YReMnS7b5ANWh951anYbusndkoTFI
oNLRDmnddSPJpKChaI0VfYkztRShQXTaZdDSWH8G8RBIgNWsaEd5l0W7d3Kstk7D
snTp+2lxQjbIsIljsOS4hFYr0uDIyPeoe8xZo34DF9dkj3w/fDzHy/VcWt3n9u/1
BSyP+Fp6xAtanDlho83/eZgtYnVRyelaI5A7ndH+no/YaikisNVo7lP4b/wsBEou
mNoGdyR3YV0O/3jlmWBgt+eUjqPS+zznhwH/Nr3k/TIw3wxKhp8o8R1RbAHzJ/v9
03lJxUUa+sGTqTcgyWK4AO/SHa/S/jzrLfGZ7uwdVC6c7fS4asevIFhNWBRFcjxG
SMy7ALbdHcX+WsDqbrqztjOlxwuJbYKdztgZuO+0gS/saRntIclB6KG2HJtYx4NJ
w/3ZzYbMGk9HRllOBTKQR0DW2KEW/+GpifHjC2zZznhCEkeL4NWVmvXsozlOv4nn
cz9c7r+i7D9JSB+4KwWrLBJky5WxroVmInLnL5o4eTU9863l2FHwLrFmGYp+NJU7
npdXKODHGS4EcyRxWs8k2BmyWPztlDsuw1aSVeJa0VzQbsCmZwM49uf4DRrEMt6y
6EITi0aZ8KOObShoPeCr0dEE/eipUKhcdbl0FBuD/KY1PRC3jQqzK3lAx1MM8x8n
URbdqrtt1COivIZ6wfVS3+qZFQSjMX3ik6pOtfq572Vc0AzCDD88j8NmNR6zRQUX
TcrI6OGpXRdWIDw5GLu+aECwtBwZg8WqxkL3AVgm4l85qPvfRIRsfehFirNG8G77
bj7nS3B9RSzDSpZqUHFFe2m/Vf69wtbAKioktF7Jnb0NQo5DvlmVEAfE4SOQvKpi
Atnr6uYg5DbadaTLv8BR62yYH+5ixYGwza5KtwesSFBiDPtaICs6tITKFYN7fiph
1ZFU48Aza5uIFZ0J1PNO7KqlCG9g31NexIZ/i7X/WigAN9bcIUClt7k4uIqaRDOj
BFMQIAMP1OW/qtWmLrocLM6HPlIjmX98BtAp5hyeTyi3L7YEM0nhukq3EqjD7gCp
/2GN5W3tth/F12sNrR4Bp4oW0E7h3BOddmLzQrntEquK8/nLfIcK93Is8nDO3HUq
/SdATw38ODjzPU+aLH9FUVA28ZBKIPLvFnLeRLZNf4pH1n8i/7cleG9vAcyXcqoA
pFyRA5YJ9/Iz6wr3HcjeEKuVEZULo84aLKFnIWzc2ctFP3mBvbkhou4owVjpW2zs
6WJqeprRRZC207axyg2FQ63gINsqz8Plk0loMwCpf+o16bR4EOJS/YN54SXgnLl5
RtFENUjL5nrSod2PySVFfj9BSmtzMTYUywVhgtOPFiYNMBaCKVEn4svCr0D+GJpj
j48ei1Gnr8liSIMAiDqNCTUk3geDoE0GkoRBH9UkRxbJpuruMmAmp3J0iWIOyY5t
Gax31Y/yaK++OTTBsz32YOpQKxEl+hhp1mcAo3+jCqbbVP1sIq03ObH4DXZQ8WTI
8rTxP+DYAmCygJQvI/i1Cb4ZGWM9vVOkWhbulNKi6SNwpQeTzLv7Hn2uxzW1F4oM
giaie/buPpQ4QVEWOdaVi2GN7hJEuOPplvWSfbnxO4+yrEGeMh1Ek55XlkDEisyr
hdkRLtXndRPR1x1WWrySQE8Jegt0UYLOUoIEJ8DdImmm4sC5KDZxnmnyacN4s95H
+HozSNbFqfXglQx4xgwDsHXJMh/Ug667BxMQyxdAjR76cIK00qS0P2qLEDXwhKnF
1RCfzzlFxo3sb04aJvZj7y51DdMuyqD/ud0l0DVkQwre74CP8XbEn4JlC9Z9u1+Q
XGDNJm8CxMOQw+JxKegLWUdOFopjoHKpY6T2pvDzLaHPnjS9KI0WGq4rYQ4FfQ6a
gig7syWdc2WSyYIUG8UBVWObZavYNEFCiQL6Y9TOTfZfBttROK9SXfhYoaI209OT
P+68CY8ONwHPv3d0ft0ezfEihaF948Y1a2SesM5Hk1UjVxjGHJ5r2CKkbtIM6s7i
Vzo88F/GAYkhE0sYuDq9yWJqt1gFzw+gkQGuOo08cdOWTStkEd4SGI3mx+OWwp3F
W93aeig/tBU2j2vTOnPLCLb0DhBb9i5/MWdJ+VS/DAx39gdYE8ND8Sb6jXq/YwpA
9a5iHsKVFSwYvXBwHBS5LKgun5aNkkgQqE+XpQbMuM2+cGM3+4nNIW1dvtdlw20P
QjAh3R+nQ7PriFMZ/RVY8fJ0eUbxi7dr+q3w1p8PKK5G9FgTSldrtrhknJv8sY42
HLLrGxfgN80D2mmrNGRlOgtFJhoAbcq9bX1BschUY+ocWsWqiTw8aEQkrLv2orV/
BcTI6vH3iNzYZ4zbACHwgTd2/0f4PMRV8K33GNWIlVBRaCx4Cw3KRA++DTkETUJX
wM5QAdOYItUSxdSqhGLmnaFrpR/jmvxoYsAnYBfT1UO6GT3Wt4lSTF/fYCkBwfIK
ZJOwEdQlexmx7teFWXGbbOUeZTCPXguw7D6/yKBcM85EmiogET4+7TcJ0vzvlovs
g0SOVQatv1PW5DhDscrycxgnc5vOGN+0Qk6cwf5PhBp7HJZzcegi2s4zU01PiqCa
yqcU68x6SsJIzWA5hGOc3IjunfVe8JL0p5WVPFzUa12EMOAJcUDAsRIAMTPPY+SJ
CsX3rjRV10e1DOHx8vMS+4YYzC7g4VSMGPoJIqHcaOkW/005FoCbY40xS1zSyoCy
nEfdyfw49R25X8PmcJET2ZbgMVv72oNQ6xLoq9MpegM4eP5999OBti7UwBxMRZXA
aTpP6e80jMTTjmdT1FypzMIVVQ8Z9BU/zt4fFWlrqcwxnM6pKW0CLt8u+zEhn5yO
2gyT94iZXKFkPpeYlpaCGRiaWcneHFbk578fOCSWfMqAls9G8lSxXNZK/J9Y+DnH
Ohqzx0D5y/iHOFYmSHaYhuB5GpV7XeF9KgT1TeSjv+T10Owu4EI2+PmOu0u6iUxh
GwyTwXo1fXZo9YxnrppuOI2/YRqm4iB1qWhMtLX6Xu506IFrvQpJO89MXF3X/bMZ
zyyCGSlli+OSM7XZr60v3kXBtQfpOAlb9ldD6Gje5z8U7ZQKRs1wXLuy2GiaxtBv
wUNQgFgccXA4wOEgiQVUKzxf1jWqzOb/qVHlJ06Tg3ftx2MeQmtObae3IeqqYooI
20ySyKOsTq6gvTXGtFesCP/jrGh87tJGbNgVnoqZmV9okSfLebXYvIIsyMQHkDmV
VoHp1xh3gS8ej7i3THG2Mtra6BqktoFyrDPwN2sbQIK2yf6Wjz8Vzai1WuBTdSC9
gFTBjHS+HNRh1cQWHe92V+yAv6r2bn/non2RfEZaEPwO6Ep/bvdYwEFO3cLLALid
iI9Lqf6NIsTWFV4n/lwYrkJWOixt0ZA4oc/q2e4msqGKoyUtpZQAYvlRFYaK+6nZ
aaCGighh6pQeuWYhIb3Ws5WrpVbCidI68oILBQZOR9vM4cPIrihhBMYrNaEzVfEb
RBzMDZM8qZDXu+5ENbOmoy8KfDzZ5q0zvBxyTeUVD35a6bs+msjO6wAyR8Xf01Vi
q7kYquH79bH7KXvwdj7u4AaGeyKRcrVOg5Qvxv5fR6Qkr6xNIB7NVDUSAbsCvjWa
YWfJrL79fP5z+13C/1dW1FoXwBiOiDoDfQJ4Akf/wbr/oagvc3at6A6gQiuJpDM9
Y6zHpr/1jmPzkKaYvPhYsLOmnQRlOuemF6LrVPNDdPakdY5Qr+NjuXu85G5GC4Gi
TWmbTLNnaILaiWBVbiZ2y8FWGpdXNyjbFtje/5L1J/9EHLXBbloqoy7j8wjFRhXR
OIkNhBEWtiJ+IylXk6iGSvPWSNAon7oM8baZoBIL5EHaQ4veBy0ZawrUR2E/6/BD
sGn9VJuUqNwxf3hROdeG2elHBnum1DcU2RHQU1GpYGsbIgsDfjTPDGGIjo/lWUAY
1VP0jYmAS4I7fiI5AY69ItQdUbqJGLcSzu+j/zDjiQCuVRK6U1kOFtwkC1+T7wAg
XyW0nfdEXxH7GPDkJLv+dlNA3YewQ8EVHxOzebp9DP3XQgz8USDRtWcqgOEOTqkt
ogSV9Cmz1B8M1on7Rpaepqv7Q2zyadJ436Dzs5UCcsLnI+YGEMFajK9ldi2jvvin
6C3Z87ZN+JurjxEtQZ2jS2L7+Z03J4Q6cgzErAGhO67NBcPrPS7TIaN0C1LOM2Gv
GfwyEF1pTATTUoEATTgHwGSmiGRgySb0Ma0L9s9Mdle4oj41ckwfwKXG7AeRaXFj
ePaCfufZIoxjxkDA+cbKsK/o+VjW0MLn/7oduCswZUpZR89inKUBKLpOOG/lTnCa
seOAX1FBoH6qyIpgShKP4Qob6gi3Nygkfgdny7RTuwgPM9OhJhwI86GWMGSdSH+W
UQgL5Zwh1TJrTz4Zm5tNTVvqJrH84EMutaW3SP2ZpMKam0McKb/kkGSoFSWdQ+w2
/lYGgmM/3/o+rQwwjUhlsq98j3tZ2nDM8P+9Kpfcr/cG0MjEdJDdfZu1gtX3edL+
0f/xQ/PxPmwsPi4sg9L20YORmUxJ6jjMqqnc6/mP6QReHNsp9hObaDIim65rKK+R
D7OHUc1o7zr8mKOsnFHdTNvu+dZt31V8D+C+nUJtyQTZuzPWOBgXz/+GHF+OxyrH
IkRsDEZKPuKPcyhD+mBi47lkMwtMY2zwaTIKfS3J/q71I0/EwrMbgMbSjqiPiFAp
MDMMSQLjq5swPWWWxgXhP9FbLcHhQMBgfZk4obYpiaPD3I4MhJQuYumjyPBkhN3L
XIYhcZO8+D4UD25NzRtkUL7lUry9F38q8w4iQwaZ/dWApiz5T6GHsfFjJrGqcEeg
75xMAIpANz1pKSHbI53vvVRayMvpPWZGgZiv6Tp0RSUac7LrvX+sNCckVtWBsRdU
9S0HDILE5FuRX5ktvbJr+jBts6EVG03OCAmCclYUHhWq9wP9DiutpEA6EuR18SUT
SKUBL+aDAC/6PPGdDTFiFedrxAF7I7gW8DfM24QENRDVTxngr9WBjiJ8Xdw9kS6S
TZq/OgG3Z5MZGjLLSmGmb+gYcRTkiR8iA5+IdhxiHn+8QMFXaLNmxkwMt8f0DrfF
m9Mkp5WPumEOemgHU+n6k9ECcjeTGJvGwmUsp5bMRhuZpblSl/hLQJe76y1utjDl
KAGZYErtLTYyWMkM47nnE0zcrWoHOCPLiDaOLc7H11F7OichCLxaBYXf9Wfmy1Bk
Rq1M9JyrdEZpmu/xFKTXj9He2c3852JaXH5y3NVLTCz0IeYqVDxxztO4A0/FUncK
D9h7F5VE2gc37QbbSXCHrdnG2Pf2EtdEeO44I2sSq17xKSF3BXXH23O9fmsPmNh/
NmVYzdYyJ2VtqkEcBV4PNCltKoTettKsog6t4Ek0TL6XmB/Re2n84zjqPJqH2d+G
8nYHCzt7pZRF/VEXOwZ0dAlluOX9h/T8m5mjLbwNmYnM6utMYo9g5YkKHfjoIu2Z
QDOC+Andl+lYMnXRaQqgH6UicC6GKfDYaGlPL4Kczky6jnfTvozNOLy/RBCEOeZ0
vOs+cDcWITAQJHrhTjbYDS4u9utM1HzgsUlY+JhR8N2dEYUSd6RMxSiEK+VhrRNr
JU/Wgpc2rOVVnbWM3pP+4danjTHKYwY1DY/QTrhgFIU2SC3whPrmGjGSw2fCpw9h
/8ZepFHNk1BgS21BRxcdQZIJJOyXnSaDdnaQUmN4PA8J07hzSc7Gp0vdjkxSQiVf
W3cZpJbaSp28inFOtgTXTdh/5+tTHjjVYu8Uv1FymM2eqAns8gO9sAW7gKVXYtmD
2fXXXsBqsctvZNWkBTvUV4ZEHejk/XAFtnl0FEafnVH9+A8padm1TdH5LOWjF7gY
EVY4Nn1Tt/aVrnpGNh5cVGRR8GuMUru4HxIXCZ+em/OypxY+VEBMrnW665yoXDzY
4kUEafp6YQRCbeMWI1up9neB2886cE6NO2gY/qIvnqIlknv00xspehzYgd2If2WA
bF/d9jVdVmiycZhRe8XEG1bVDTzGdAIQTvHleqUi2vUKM+di8Vzlvv9ySZaiU2LB
9G0mB4JGzpnDaExcHdiW8nZY2vyowTrQwc/wABAH/96tPVFpmsmB26yVNsN+UCqT
oNN1VxDJU7nBg3m/Ir425F+gwQ+q6JXQwVzZzvhUGoQzjAXnsPeYZUlUxwd1GF4g
kLufBkh8XvihAGgfKV7Vqe98LAbYcV4WyX66g3/hZkJ/pw2CvE1pe7Rmp+UVFQxP
vbrUS2RoYuQW8JEYHuy3Zuf/fEvTy1uVWXn30H+p2ZW+HpVW+fkP+boLGMixVy4z
856af6BwH4JH6pnqQvyi4V1kwz/y6t4OtNZ2r2MY8QI6OVGYIPi4ZwaDQ4eJPXjq
8HB1Wsg8OmB2dnyheaxFZB4GzoGaG8WaBKW9e1TQ1ArsfiwpoOTIXy7R5H4YoGle
bkpWwKlUChCdPZhUuCKRamkbWb8FJh/9Fm4Lr0qRFLumV+5A8exuzuJcq6XJIPsd
+MiL6ptW8D3LM6JfsNEUSn3p2cGP3JlJWxLZ2flajZyc/SQQswUUYkidvfgweOTt
gNlG8JQmq/1vdOoyJOW+LI3olU4/ZbA4aPyfiBbcJuE2jFa70cfzxh0V8JbwMFlB
GhDx8XFJjc7McfyXepa5XTS1lu1U1EuNuxzsY2WVB20qUY3xlIKQ9ivqewRHLhGF
ncViJDltCKGMLpUKigaXew==
`protect END_PROTECTED
