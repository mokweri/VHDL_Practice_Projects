`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
26uTRlvpZAAhtkfk/KgGAq8jWqMNj0OawQQ+naSBSV/qXdZg58PXa2RMJfq+dCIS
mRFm1unez5Jvxqy8ChRDNTtNobbyvCaY8Zhdc5mJPeiSAYvd32bOiPNrwjJdOyuS
eP4hl2INur3gNlSrfbi8vPMiCUObc8qUBc9Y8i0VGkFeGy56bUXlPAAv/1SxQNdd
EWEQK6Kg1k1Zw1knqqgZbjosUh9V7krpg837rJ19CZIdEUrwAtTSEVbk5OXCHI9g
8Bj4Ys/tLp9AF7CNfNTW3qj5H9tmOZIzYrvreLHBksydoOrmvtat4M6sgSD26enF
F3Z/2HmIZ2ZM8PcNDh0kQdqecWBZOH0wc6pY7xFUGw7P6wyFfyBOB9jo0r4GfuqK
QW7npiQZPXmXxPBMux7m43SMyit3duXSHFqgYPPIffxN0hiAQs3YKUOE98NVwN3o
R/i6XqxjCPkaLPY1Lx+FNAsSYsKbqAXE6lZocjAPR90RqrJHHNWbokxhOgz/jade
P+dHx7u1kHOqBL5rb+EtqIREuy3+OxUV4RZG2FrH4gIL4mEJ9SVbQYXfx7nJ5j7J
V8TbajlIRZlH2944fxQLHv5CAgjp7+TCKYavsJVCNnuriJThKroHCyMhOe2xDr91
bjb4lHksZibsBV9MJOxNE42jK9anxnexb/nyYbYPyvJ77iaLwBbTGB/vcHhKe7qy
dAs6xOQ0xJECXT3T8UYrq2y3BEEgF5KiltkwFkRxE5OLBAaV7cZUsdIb5KPdmz3+
7JVWVjxEKkteJ8JZNOlo65po+7Bhst0vmyUGLnzFiVIX9SOlUMgsnC2mt1JwVe6Y
dF6JeQJArfVNEWjxGFZUIQ7bkCNWN1YVFi2H7oeYakBEfIVM0eK3PG7Pic0CG4Ni
2Tiw6VM0Ju93BokCW5uj32asYUekOjndOkJeFiIUYWJonSv7Gpoil8xfZNEPP9+o
YE5IMipAFXA3i9SywhANmO83NihEa1/ANx7gAJJ9eKXbHX5dGkWCKIwejEbaDJwB
LtzlJHzNi7ObK237F57wf6fNsa7HAfiGQ/2EkF4+BXDawkxcIrmYYHcoWUWgAvf0
ERlqVNiAXAanzakmGkmpWpdjpZ/AVEaEmmWjhA6TaFI5/X5IU/aynOP+LPbURi85
axaZg4Hmjec0hSCH4bHEXOQZpj4VMaS13NFa8QfZY9DiCC8D0usQrj1vSmq3vkGu
4NLw0Se3FKOzIhEJOSi4ng/yyK8jrB0ISQveRcUy4FvuGgyZhgJ2Zz0xbUijqoK7
NbXPnaX/iE8n/rfsysBTExnT1pePyd/oeCo+CgtCduxmD2qmf6+pSh0ex/g5XU55
gcFZeQ4GNf8urzKCR1wXmCDnDPyCbRFrOjaQCNX/RUSrapXbdsteljLAic2fRdh4
5FGuXCZZcB1EJcBMXNnXPCToAVpbrZmdCgLEZ7JYcDQOqQqGZ73rx8wZw86aFJvu
E+WT/8MAn1z4x7sX/Lt7v38V+vcZ+QgP1Rbg1/Al9fHwDmu2Ul7iStMORRgxSslR
rfSFC/gSgXmZkKqFwdTHx+klqogyg2B5oOp9Bl3zF6ZB3i4J2lXFhPvqDcP/vmlg
uqndn2Ltgw6CEMNjbManI4O6em4sZzPuCSbAAajnsVn/AIitqw4ObDk1U9wUwDVB
oReDliz3QKL+W4twmcfD9l/9sypRWH8Vn8mWT6ioIUsfJkvrQ3tDioxmNjnru6ww
VyqmBfjOwqY7asOMTraw7B/d0QxqLsqRD49W/EvUioll6CRaahGJ2hyg4bdMoo15
UzHGzWan8a6F10051G516lpmulDxXT6o6HRfu1SCI/rhzq0oA1Q502H933mkJZ1f
VlaDshOMtcnsu1DsDiCFjHA00RJIPWgQ0UogOidyx7yVw/uFLndAb12RTw21gd0b
am1aMoJ9xsv0ixRLGx9M9brldNu2g2Zwv35xa0B/xlLv3nRScYweMlOkIevfvmvf
hM0lsEBtEfa/X6jjsDyQlYxwZNsmF6LjbCWLMJWNeFGDnhKBd6JNZnta9epXw49g
o9a6plvNUtSKFqcmCJxKKW8NByNQpLKGPmKgnHFBuRqedHf+eDL0a2KtozdcIz4q
VBWjw5j6qwPxUKk4GlB+EEL+YN6KqdFswbtUkaKRVOBD62ELZJoOxDieyJczF8Wt
9vA7fjh/T6qwZxqXH4OwrBHSTs25K3dTb0NWKnzR08R6WJWmBQjsi+iUvOyzu3G/
arFz6hbWxtwQ77YcU3AnqLfyh6gb7nsfAzj/5Xj4KQo9c0HVtyBcUQbQbzbYjFBv
CoGdF8O4/nAvwCQe/z6kL/YGM2PF0MG68DEEWIwvRBaVCRJ1/Bfb313vYh/OMBz1
CfVbbrtbfAJdmDrOBnqP/o0AUYYbLc1AP4A7VSOptgIYSR/y9GVFByhIuZ7fHK6C
tJR0MNSpI27x9eKutDi3JcT6mIi4PrZN4sUrtaQj6MEtyFpf2WhIwoWR6iMskJ5G
GMxyAJr8Xybg+wfZyde7BJSI7+R8nYiLefUNdu7OHQFCUAizSU85nbXDBqKXM3Oj
GCGEp6Xmc4foEhRvq82NSHbFYk6q5zmGoqN//f5xd3CDlQ4FLs1vWKHInJWmDzku
kMXmgF8B3jWHt1gcSlk4wUif6SxD+SsgAkCcK5Aw/wRP6fZ2465/9LObQzDNjiY4
dL8UmBRZmZqWRswJkphaiTjnWYNL8fWhUJYKQjD6nZUlh1wj/DJ8Ljx8Ga3/5nn7
s0Z3deq5nlM/YCaQ6JrvCHZhe7o3hgMCn6P5lgze80UWNHtkIHcX1Jx7pAfk6OvB
q5+6e07M0xCBRbeoLMJepMx814z8rUxt6d97uwXMVyF1qZxY2j6txRMqRCDkCP7L
soEScB/J8z/qAP032B/KEWCFEYyfPMawsLTq8UGOCOX0pqEfdGxJ/HNf74r+Nxe0
pzINqUPvPkp3kWqMuvUOZdbThNAfhYvsWkYoduWOmY0bYjJdG5qs8VjT2ui8Q7uz
dCuWalKJy8y4IcSmbu2AUVHXQR4feo7how9HTA8XNyjrxc0yz0Pna46IGUeG8BKO
lQB/qWi75505tRFZtZ7gqv5dL3oW60KutF9iBFM9axJDnAzfDX72wCklZj/KJP1L
v/8UGai3BLcbUZdj117F6o/rigdQMCCyMt0gb3Ed1QjSDabZ2nf1LUaf91kLGsfQ
p8U3ekdJTEMGrkt5dSOD0E1YksjvIpA+zle1PaxWa/atqDd2j2571GHFUBAy9efq
kuusuvZy6EJ/gn0gX70BnXrLg0ZfNdufRQHAenmAv6cAeHl0zn45wtuknXXDFK3W
Vmpwsx9ksN4Z/YOhZ/L0JV7Dfj+9PXOpOwoyVqiSIizi47NNFE+/N3Z8wi+9Xbj7
Obt4zGIi7gw2hTX0b/bhhOpn99JgX/J0Nem9Imj0fDfz84/nnQn71wJoCVtan3aB
907rPBbmj4Iz8SZ1pNQaKQcTR0ewuhIuiHzho3qHlAuUERUvLEqknnbl9DczTiz7
Flato/z4dlv9QXkXxX3QB/04dCBf8De9Y0Xcqy7uw3Vkl3VWjnECLVdTJklkoQ45
SG54/a9YyEMS4zkSbN7sXUU9NDtTWVG0Xu04J2SUq9wgMgobHtRGl99Xg7TqSMxo
5AH8MO4dHxwC5JPKpEn5bMBHnLK2yVnCw2Vj1jX1iQIp+o0F0PfVDp017EGw50Cb
JhW7fykuqgg25mhr+E4dfEHTK6FVSy2poGfAmYyaK7DBF4TDs3OG/G/vHWpEz78N
ZRlZWlHTwRnvg+w6Mwa+vkjA7nPPcuIqaHz1OOs48giIt0mxQ/lguCCyfjSod6x+
06+jGZxx+0c2JtmYSwfqdloagFtHaAv6BPOHoSUfefs4950cGdByfgUpSdixXTT0
Z2Lk9CMrVMFboJ0TvoJvcux+qP4VMnq1aqa6yKXsT57CQdYzgupNO+lFbN3tRu9n
UJNLsybN8TNNFLkXQNaxUOAPVXRXM1BeIX8jmwyYfVjddcfobbyyDVUKFqNB2oyQ
LzRqufF0obREXmguGcPtQYxDNELo/MDOsxdkyY+OOj0oBlgJOjphXYSDp45r4Qy6
Br7+g6JyhNx1qxIV2VIZCifR0OIv4fsXmqIxhu4XVGz7qmayrOJmEAzd8LA4KjDv
4eRSDwTeQoQ8KrF407fizZSFISvsh1ttJaTLjbREqHePhCrQPovH6JKemPfxv6j8
T5asmNItzto2rkXkjHfzspbBP6oIcB8N6FVi01BMeemaDWS/2+z7RUW67V2xGYu7
cuXimHbgAJGmHT0HY0mIOhs4wM1gS14VmzqVd3xmVcwu6ktTSCYV2h9KP4lyhqIG
kwxxUzoUhav1u8fy6UjcU6NcMRB7g2gT/1AVxeJLV5TPB1Y84Xn3yRBbCclkr6IT
dYDSXSoy1RxGT6baayplpR5AznwAAr1MoKIzwBuWe5nmE27I2i3DXQ/yId93QcQE
DB9Yx4JHHMgN4M5EXgAcEChzgizPCedwPiSmdWSKzxysAq8nI3kL9w/oYX8+TYx5
WHerDFQHOAPQ2OAMF4WXWOsu66tqbXBWaygvRnL9AFNLge2lWJByAvmQ5nX0KRj3
4RyMsqyPHzaqTFgYL5KLLABTjI6iEkD3xCPSms3pTeSEhaXR7s9D0VOjPrWLn1Pf
IwdpUPnWZOAw+fOkflIuXFpFB+wu7sazLeawXoM3lnySs76SiypW+NG0QIiuizNB
0sr3UxGxAaZ1rPe3Qgqt4yZhwJobQRYB9S8YS21juuKdTYYjrrToyWNZHJSm8zcU
IF7488Q96Sh22C9ic57LbNOAFROyI2t/aaZIxL2QNEVYAiIytmjp4Tg3M99UeI69
DlU5QBRcvq3onj3W8HGZlbsuDoWIqGcM8SAh2wpUevrK1XKODag7WszTbOW0dOkj
4yebgNBXYAGSXB3ozo1tkafHZY/PxyiP/sy7hBMToIq881AEtj90KBCNzUft9lXl
5yzievoFnJqLr0udGPM+ccos6W1rj1v0wtusPzhfg3sLRsTTSsGyp8dcXlCK2Ikc
5s0BQe6/dnMw721czHmBSH6jIzAUV/5cheReEXdCLuXq20xcnL2P7cKq5B0kfV2W
Q7ziMT52AlANQ+AKig4yAqHpphnikf4q96ueybSyGjNOb6HH2hgR+9MHq0v6jwuj
E9dvOct+5ldwSCzzUouV6ZrqKghBASArEDLtke/ZsQYkiAuH2sdKzOLuiQFQQ/Rr
pcNMApoxCHmSiIBB6DT5m24VkPd2bWmI5Bx5oi71kiMDHriBAzqJpbOWUCzqIRP0
FEzJRf9tsvK4UcRhT5ZAQf4FtC/0YmALjAFpQQ2qUjwm7ji41SL14EbMaUYLIN8r
lU8lt8P887OIUF9Hs4ZhrWF/hpBzpnam2/EbcrGriR9zDCKoTzAtJVRZb4SwEBla
FCpl3ni0dyQoYAU50lTkc6F5Sb3PKahs3G3hyH0jzDOJFgoauQZSdhYldopnVGq3
nD5/SR/r73gtZ5gBYMG625pJLkPucZ6esm6jy0jJ0yiJtEYC0AOq040POf7qvYxP
MsWxoBoMEL7Ib64pOeVXfvRrexpa7oMElLf/bHYz/M5Tocl9XFJeanG+JkdkemPL
dZYbyEPLsN6eWWAfXXbfp3WpEeaM2GnCJTUSPosaAl+JYBi18s7mwnl5sVd8is9t
LHaURr4xpOTIBbqG/0AUB2W4kyQj2Pp1t3N+5iprdsTsFnwsFH/EftU9Y9aebu2m
oTuJJABWtJ02RzGN5Hr/X/RdnYUGxcvBHu1TCaCcTDeE6TWssBSEFGAFF2fH4Ivd
Np8AsY9meymDPZppiMCIJ5fOGIiBp9DTzDVZmsq3wb9ACBBxu7tjqdq5jT31foEy
VqKjF71qTgHunjCIoNmHJCMk7/F97OGNcxvOHAfSQQdzGXelYJUnBxUvHUfOMXJL
dn9Fsqf+DmqivBJxTsgSw7plHa4gRZ+YNrVTweGz82AK2E/HlPvZG+Ujg9kGXHWm
bAjI502azEIU6TKIhULnDtuQtOjZVbZeZRlu31dPMALUlArUkp089sddovDaWpU/
Zbi/vL6S+srLwJGHCw9zcXrwlu2j3bDHI9iUaK1NH1zMLxhf2jdKNp6Q9X3jwDnL
/As6Z8Jkwut01a3YB9ELo+kHVYXPS58nv+1Rk9M5SyP3oYJmhaYiWuQG552/bnlX
HwTXYNz5PQPna6IkdlJCRTLfM0svVvr9qnIANWFnqAjx1YlLfNa26MsgwGlAgfGR
V+ldru9+7JNhACtsbMuTja+LksqtR0kbfDWf0G1T5dIX6CQyf20BTImySvDX1GPb
iZMVdLwCCuOKh1ROA76fUvDgNSXh/vCsX2pzqqSSiEvq2pGYVRB9sQT+GKObV55C
Hwmo51Rsk0SAlrft+tv1z6wOy7YCoOFrsoxeYwLlCnkzY+y8AEdE446YcWwyHsYR
rSEbwcSlrLaU7NUiwiRRIOXBF505Af95EML4JwFlD10JQ1WH/AsAHulaFb/xHLbI
Iv1hnPx+XzjhaMvgGwN0L7VI9mfR2NC18WNYA3dZi1hG5WW58npMUZ+9QW8r4pkC
deJleQWVytsI8AiTAieHM773BKG467is8aAYJwSQgwKWN7qvBuWZAebdyW7DZaoG
YUDipcUErNsTuzdkifBySfs6WK8NzL9oboeK/B6fIA55jWbRJnKQPxvTC6as4kOT
whaQ4rIS56lyVvfYQ9NRj1kz3vwFx5vO4huaSwRs6Fk0Q+WxVioh2nNnOmC0AjJ0
57HvrDhy0SxjMFHIcOpAF0SxRyci+4mhdmo+QEB1+1LbhwpANvBd5eG/+hhmQbmD
s6Jqr5Kqv6urZ9+dMSK/MPblefbisF0umhaOAb1iEd8CwkzIU9KbBDNE+vjExqYs
r3Pj0y4qF1V4jM9vkFGzO3a1zG4bgktmbqUGLrEsYUXO6kOtfVuhFzIEM8nAFJXm
s+N2sOz7vMZWt377EGNCAiii7YGUqn1u9IibDMWCcJY/qU2v+4pkZq7H/o2Pe98L
h8qH9hSZf4R9zaktE6/YE+wODMuJRqsH2tjl5awvJcPDSZ+srvDki0a9uspz3Hqa
eHaPKTUtGiKbFVjjjzttGL+CAAImekTR5yyqNLySI7gQcNeKAaKWSPncZs0cnwvE
svgEI8Xd8sGBWcx/kBzaPsLxOptV82CSIreNX3YFZMYG+DkhDb6YLs5dRdc1eP8T
JsKVStyMGS1IuQoSeXL9wu18MsOJ+6nyZApSHSjR5GHwuF6XQDAo40PfJLy4c9Qc
GM3F+kowUboh+7E6QeYeio63Oq/Ib7/j/WZKJxNmyiW5hqdqGto7nWDaQVwI2U+s
mblkXED2gZeeHEeHjYcGfkmDayysiSQUsoQWzURQVUGca/uJqSyeaHfpXJgq+aoM
HgOKxJROENeK2My8hi3Eq6aLMTe9dX/9YOvSgh+OlKv+WCrkW/MehMTCHg5/97fG
joa2d1ISWaeUN3asrxLpQChb3mvWEBiLOTGsiRaylHLQOoYMRhG66FNeXvrTobrk
aar+FEETK1FQ12SziCt1k/4C6SIlXspKN22ENPoN5T9hej84WOfFsX5GRQ7hqrCe
YwbkL/aHw9x51O7F9EQIOaGxUHr1MPCLF+qX56rOsbhiqtEtSVggLP/9iPKwWKTu
OulYqP1TUgg0p+CIt1iol3VxWX3XG6+8QVUN+N4Rjj8UvuW5PtJDBXgFXRSNTOJt
cpn7rfXHj/6Fy/cQS2zmV2ES7Rg+6Kjq7TsIjSZUl+8LGMvixG8Qrjsa0XBviKLc
kcjewyQTJqu7bs1ZY7YgWPeaQqICaWVgtxbpWmHWiRPJ9+J0JwH5HlyUFbJ/Z8Zp
j+gIIgfah7MNKhYNsmFH9B8OD21UPnD3RnO/ikuG0/FuhRnVRZwB9a7BrqVuTg3G
CagxeH79xyORWXR4XiIqBlPU91ktUyYgK1U+tHEdPLrbu3DGYVeE+mhsNFyVu6My
LtU1uCRxYulGabNObcAa/yuy9MCG7PATynQmBc/WCsfq5ZxurMoIkbRrXi2cYhJH
LjEmSXAuH7GwkXLbMAkh/wVUIzLli6C8Pgy5jRiga3w9xJg/3s/LEbE0v1RgaAGX
3IOZEsajEOb46bZaM0j6WlkhjcvM1bdbs6/RrI5iVfCFSQsH2ikLcjcPh7R6tJMj
AZ0klwdZ08Q6ZFhPtFPTM9nRNk3fn/eKMzHK4ziLlmTbTrugOVHh0iFXsuqKbC4u
C+9wEO9a49M+2pSNKsSEd6vsasLuKIr/YYVr2vsJlvpxKB6WSJcfWdjteYExPrqO
t6uoBriHDIPI8dy946DVmRwoH7p9mK/+nTYub1RT13Z++72M4sYCHMmkD07zpnx/
Zeo0iX7CM6elZZFZuRlJRSWFz9FlcjknBiSqemvu3Ho8BvZ5G56+CZz7V3aUZXug
cOEN6xvVFTwiFC9WADoq0a5E18dK0QZiANikoh2mQtrMuZz6GIvRup845KKPVnLN
VewD69njjPXP7MyuqTr1xrqT5QTF7bYVOzbDw+VWnzMfIyZ/JTJtM6NdUdaehq/g
APuHavmKjKsRWP26K8kJZrXCQqqflD9tWcxM3hBgbHdIGP2ZBkARoI8sOZ7GZIq3
AoRBH6Gdj4YUmtthEHngsKOlWsDDac7FZtKueQiI3qohFbYi1EsTNBB85OKsRxoy
cEjVy1HT4sOBQ2eFTpcPUDw8YJ0GUZ9riwBiObTXTw26EPngEBylW93Ga/I/Swwc
mIukpu9NPhIKxhvO/Q1zasrQYDouB4n01RgrTdHUJVIy1YfV+LD0BfeqluIEklp+
grddxAQ1ddwKn0JjqYvvdQEuY28Ux3aainHlfkt9qGDkmCQTewSox7DER6qKctc1
n8A0V/RJEb7BMc96z5uM0eHN0cZ/BfdfJzQ3w2qvOWNv6wJsphmAmZD1myfPjRZc
LSBgVSUqW23GitYl/iNh5lbcUNXfdiPpXLMX2R85aonF7GvT6ozkZgNmZtb52s1U
Dm1TMkTz1D9NQF71065wckgthoaOlpjbKEvNk6kiJL4w5Tnamk3DiSYkhaYB97jA
WhLSd0Mrz/ILPHcXACQk86EtQl0fexhW8UkTUfGh6MfLsPe2/vPaR05rUspe77Mo
YbosMZr1V8IqOyRxn8+5NRKTyYEdUZy9jh8m65Rg9SY3xavArmNTAlemWSAjGIst
XzUu8EgD7MrcFRQFC2qdnR368STJv+5XfkDXeBBYEWWWqpy67eBFqsrjwVAGQWUz
XX1SuLLdVSGUgDzxLgIbL0AWyOTjOv44OQrq538NxZ6Egh4vQ46dJPI3ZliVMj1b
bleuqH6rb9egjx2GxIivbbaui8deQcuKpzIE11GAfSReFPoNI3HiwR3g1vA/bwiB
p2DbO7NlEI1Eqm3joAC7jxj1oND9+LY5ydxHBZDkFoEcVilvjwIyTWxXWUhMDRJf
m/nh/BZ9YRUTZCIaUcgPw1BfqjcX9Ixmemnml/67BaEzxePCCLdXYBgUSj9DIaAv
NSnm5PPxQggoYSe7ea3jNN8Pv6pEYIH4imPGW8NckAXr29Cw/XAn9IgnQ++t6ZCp
MXo7NX6zzumbyFSbEVXH6jWsClAnIT76tPksUVh4sF7TqajOuLT0qB6egGn0UFhj
PTvd242VLFLekEie3xEnAsgScRBgK77UAZiXsKihk7RwduYwXX4qEBtKz2Zp2pY/
kBkql+Y/Srbzz3yGt8oFWt6qn1AGSLxpL/xT11F3SOQ5H1oZXd7AV/FWk9XUZ64N
v4vPpwazI7MicRGB2ppts4qyy1GFOecaMhBvcP+EAqGf//wg4aQRF18/hymgaQVo
ALx8PXCe740FjeO7hopQUaPXIZqAkEr/GhlSsUe013N69HDyTEho4VaCP22Srd2d
ohSH4yzfPEIiV65MTLR2W26GqOjEojrygMq28HSFZErp6wEQssOf3sj4IF2U+ofl
WKvz1h3SMZjpY37fVOj5WlPS2ix1ie9Mg3POIP91KHDe15rCR4wdd0CoKURYLiyg
kE5cm8iVW17xSqHkzZDE+B4qyzUmVLuBuZa35B+JOzWBXOwLVyLtaze/z1LluMOe
U8z2KdiUS6gRyD9QtBCm58a/eSvpvah689N7PPGgv/mukrhnl5buWDAQNJ2TINDM
NAmOXJpG9Y8udDEVtY8VY0zCFsw+RsiKDHx3OWLNOel4KjVLkvBUicqMyLf7sXhf
iaoQyZ2o5VAirZBXugoPe/TbsbMCOfQiE7vwIsuDmq0cGdtmYLzozfRFu33JS30r
c9RMVSK7XeMbg9sQ7IDVFwLlMmmkzM0LD5CLPN/0pG82Zqb3iMn6wmp3QXSZLps4
9YPOcJUuHuf+xXuS95fvkn6RvFCFg83o+fGafumg/c9R7V0JqkXAVnDM3a9QydsB
rcZsAVCEXdNXDox7WXhxXQoDC+EJUAosQNguFCATbwGyZw5xpNRQNjEo98NFcwHb
vUsCVDJbAMj0cCYyM+YxMBb53/M1HjecAfaEaKYTEcB5PBadjfE5C66ch6OHeNdj
0KstjrWcsls1oRBijX0NpoVVBVrLeEEAcBYKcjiv6TMciHjBsJ4Ht0mjLYi84QTd
WgniH/y69uGtSyP0W9iI6EA94sSqjDqROHl1Ck0uRSbg8WVwoDe98NiqNnZFJ4NJ
AplnlBVcnnuw5oxvg+zIOpC0NTzyfnhXGM//z3LgSZv7NNKrjo0t210Fbqd2KkHO
dN6+lqa7k2IcZVnWAdCNbr2l7f6bNAUozdVVCJzyW813OQknMQojsj7uXlxbE6Ey
ADnvPvovMr8qQKaHcTM36aT3A5tV3VCO6qS7lnMzr39S4dv4YtBvx03iB6kjKyYD
V4nFPzwL0SyVy9PtyE6TwAf2zRxSnT/i0h8n29WSJt2/Y55kLPQPi5JoG+90dRw9
vzfPX6SRkVOQKMyY/xaPtSQNcHC7r5bWFPO6gDcgpTFpdc0Wfj8+nt2SapF5wk/V
6O/HT5WF69svt0iHeUTu4uS4gdiLrfSqxZouMTLXYzYtvqy8aVGlzIaDSiDpsBfj
63hVjtHJfKTZGM6SvyY5Y1XzGuzGlIPazl5q8zyA3+ZAdG6V7MmBAZF7ipoClbhu
64ELyDX3mkd+pBdCB/r65iLPbhlu1C9rhp4w3loheDOSHNy/Tz5DOWXwtDEBmmRZ
0Nbz00aa3MGtfkOXXjEtHGcdzBcEKrxtD9ZOE7mI5Bk+rHR38MVA6Nu3MP4VBVhc
vMlNOSHIU6HBMJoSMHEVB/pN/i/8xX+colfvdODIyb1coMXqFnLQOGxQuWEcPf8u
12FzIoiuBW28eXcHqhVNbDC+VCKf5yarUY0XSjRm8S8MhrEGGj2KN46JFVdFFfru
42yUgjiR/9PBc+h8lb99zEzqgiurUbH8fVjB4jcoGv59w69tvFE5QrXvADHkSnX3
8lA+D4cOB7V/R89bFj0PMHKUWj8gXkskeR3bcos6374AJo7u4wyUpSn/yjLVb33S
eYt2y3sFH7MFGVR1CsQB3GV21jnPIhKopcoMfZ9nG8hj8D4NCo0xWdx7cnduZ35a
DgZYP6uQp/IrIcr7vcq/988LauVwy+xyyMC2GdGCLVnSjjavO91RQQ6QEH/SjnRV
6qonjfS3beyIi/89NekJqjr5clm4Ea6VZjK8j4MvWVwYqJNCsh2Tsoy5ZfBamJNO
NClLMBcv1byF3t9y6cq1QEGw4kY+vi+Of2QqA0JeB3EWO2L5r2EHF/16UcnZSZTa
tCviY6SKEbE/DNBAE6wceVuCYJlVfM+dcGgVAHn968gfwosnZNHRjQpPs5MTmduY
fnw9flIl2ATG66jltTMwAvxqseUGAyrLkZV8allJsaUp8/gc40cWEYIbDr14b+O5
oz7OKckDtYcMa8knlNOv/ncMuSiJOaERcgCeL/wvSwX9l0iswNJXV5hs7cagzWwj
DJcUZMH4wu1hlcY0hIibVquuuqTiP7MJkzH2P7No1U8/liz3KalkTj1+TA199UsS
xt60O06uF4p4ONXR3Bgt97gUX8u8dJgR35cZxL5K8AlR6VUTdWh04KKBtgcivLNd
viHzJ/aAonGET/eQZcnAIoblSFV9YXe4gpSvmHLnRY8twpn4ngdFNzD8c3LsS0MF
XnN2pJYm8ABcPmLxha9aSQoXGlPVXJqEW8AQ3Bx+rGKEjG3j6yG8YvIGaM64D+Zq
GqYBA0sF6ODrRFQNyulxI8DRv4MSInlB2npaWIl22EkFEYQ1JwGtCLj0Jmkk2UYF
tYk8mp3Aa2CF2F7tsL9VJNBhEvOjZFnXjncA7cVPOIALbjRUoZ+slXCpl77LYhVD
ZDJgZIviYb/DW+EAQy3V5dQfVfxMzpsbRTcq6ojtz8MHQDBiWQPEwnTaTbCKPIyh
RiNiEDO8Y9ayL/12i1P1WjLpJwka6Lrq5+DGtAP2bYHsHuV4vwbpi3qJmlbTG8AZ
dtOu43hS4nVTzJCuFMOxHfEkh2bDHnX4s7Vk5j+WzPolNHWtApost7bsv8E7JA2f
Jp+2pwTaBnctTx90CS9ZRNWOzHrvHuOVw4rr/sP1deByVSDzk0+sXAAVq++dFiCY
t3lzszsIppN/EOVHkToHkJEtYclSLuaEcOtit1A3fyRvLRPoMcmv7X0Yp20kFTzb
xAXjlWS8Cy8q/nq9hLfoGwDPkxyV/xCLeMq/9vZs0ygFael+kyJQh9MpI8DrLP2T
7iIjak9aQYOW7ZBv7T27S6IGJvoGdV7CZCXqqQDg1+CuVXdFdjnCSAsPmuEO1MoY
iMq96bU47TPcOhNFp9lMaiPArjZJjCKCs8nR/XTslpA9NO15I2csT3EQ+201s3gY
ai9VhnvUzrtd2kkO2hnYFDqJgw7OHlpkZ22APmUgJa6cugaFeJ8lDd09YMwyZ9t8
Ri3e+qFEmrR0Kjev0gpPONL6FRy+Hv8cbIskPGttekcZG+fWklbvzZtcEcqiC8er
NeobAaUdsusiJQMgG3sldSLt0elWDg9pFdyaAIeR2O2YnldAuga5jzgc6L6SJ9X9
0MXTb003FdX75ghnkzLp3viTT/fZYqXCQ1PjP9TPKuIaxOf68vpOyJ3TG7EQNJt9
CfEC6k4WgunN8SLQD6OGIsH4frSn5pcazprqoBmX92a58uvCcvv/cRlhks6ief+Z
+SbZpAe+8YZJqD5PVIJLF7tNRxYZRX3b5gM+jWdhft2Kr+9X11UDj7/y2/R08wc3
OeqQ8i8ZrsApFE87GYzF8aDfmh9ITKrhIL04l437UAKrpGZl1izq++Hu09K3c3BU
cAWDsCyKRK/bwOmnrhW5So2arFGpyJNwQJxfS53+IS9CAuCKCDkoPO1Jb7CnVXQK
3n1/VdAl2+dQeDXC30ANZReAtyEjxPPZa4rsGOjSUS3OzLgvHrFnD/hAxa3XjYsc
icYibMkYDHb6Kv0odwHUET6JD1LcLYVGrGD8OarKiW0EncQ1t/A85C65ULlOw//o
secOORHbiP/tcK+BdUZhlO737WmWpcm7bTYAwF+VrNOnGCkvTgmlXGMEWhZGgVPz
DuXw4GcuLK9i244gFEcpotwl0pEhL5iYhcriKGdtZyaJZt86RxJM8qGaUbG8pG21
vYQymW3uzN0QCKsAFcNLxcKeBx7rApP5BSuJsvBPo0YpFfnnYk+FQll/j9SFym/l
98i5aoBBqHVcVZFUUKQomovV0Ph4mHXIyki7KBS/HxsnaXCVN+wuib9mhOCq8fS8
bnsX13arkKeKBpFLPMKKq/aGKmAdHJE9EtosNNUeNqtHqkq9SHAAp2y3Pqj4J8wV
BNLxaafn1ATDrDjqO8ZCY53LKXuC9d4K4XTVy+oP1Ri3TNIeTrdokbD8hEuVsT4y
oFpNx6hc0w5M2tu+QiYRNTOKIQqL/P6nJVoHVxpKVS65vjaAh5izNGM3gKLeH/Jj
wuN3Y33vDvNNTSiNvC/ysrdTQ78CWB8OGmT7hrZ98PMDbY2cHtTcDytzADMwYUhN
yceGXcWXPNhTjqd/4Z+LOip6Djm49o3LdHkGTEqgINFZ9kT7APD4eM2KHdICcYl5
A0PB54fiqGktDFRlc7MOaex+ILlrIrrE4rUAUGHp7rurJCxejYwJZJO07nFVr74o
IWo328b48fAXbE3wa/jvUafUJ2jLj0o0ReY5P7z5H3AGFmRXBCETPmFgiTPcul6c
CsGv0QRs/YZdhEGQjmxcicnqFOs81ekL30+29rI35KgpqhEHmwlgWnKDRzN1xxz/
qCYIAWbKdK4FgXlEe/Yt9VkznhUTPYV+5aZh7V+3JYL+Dh/q3ZZokKl1iRTkxlax
GQ0TPTQsVSXMMBlTZe2PHJjvaKDlKPbsf0LM7xNuRYcTdqEMukciB9l0ZtFoNG8T
zNVb2u0GLUV1+j3556AhupBbnw1YacBMxB6h9duxwFdVQ1/1SOq38GEVcx2/+tr7
SSW3SealWPXS75H8RpnA6go3yZQ8u1jUvvmzbhkVGRhymzA2euEOV3uQ32eaD3Jc
x2BcJw1e7cG7+mU+okx0lDmzlniC7Yw2un/iLFCJNZ7XJBgtb06lLWqwzSDhGuZR
bWZFWxpdPsMsI4peS+CZ6euaKURftpL4JJSXfZf6wH3gahVcKb+9bYX4wCm77Z5E
VwTAoLEVfUjXZwVCqJQpwszXaIHjXZoO7XUJGPwgLEWkrLy9aX4e9KRO2txPVVZB
EQA8/OdIxj6tpFfJptCoGGm7VZAKnVFJsnCeU0edU5IGONyva3Wpf15w4sg4cHt5
zmEMFr3G1HL7Kcmuy8T0VvrAH0nSZa4ldgPhZVuEUkZwjCQS8WdpJcHcRRifI3TT
wpbzPO6vHBB/cb9mJfMwXTCWvUGkB+oEO5hciPF7bgpXL5XR9Fi2ULrmn4YUH2mq
3HdbUAwQ7A1EyhEFuPuiTyfKI8VEbI7jRiQ2H67td6o1mJD7ngEiFEVMhhq/hUnG
lwdEFvonksGsXmukiS80qboz5MdMjra/Gw0DC99w+9OwD3aSDuO8iNwg4BxsMmyY
SrRK7Uhbovjl1rMyAXn1JM11u3KKfBIP1OkKEi7e2DKYzxCaRUSXiRIfhHAB5C5H
iHxsyo/K3koP1ZmMGtNrDWebItXI9yO1YeHb9e0dqDWv5/ps1scJeNAqi2y2a8oz
Jngd1lLrUha/o6JnnsodcZPtnFe3ArEqxdGrniQzD0eJdMnu3NFwNEkVPgkSGawi
tvifzzkTLJY/B4ePeOdUqI09ww6NxxSwJA4NLL77IFIiubrX7u3DH7TJweZbCTtq
05pYpDNTyChCxJPR3/lJXHm1A7OqVtCsOy2BL5TUN2SgF28ugqAiOleXMWG1UYRU
Wwe5dmF3HfTsV+k1KHa+rDtXbxPxLSXlKAbmXgwhcfPpqfCcxMxRUo10YWLxPKmy
bzzSDUMT2vd5om0XPSqdMkYA84wBCMyzQwZlC1Zz6/+P5z1Cuj5GQYh18omJESMH
ruRzqIQmp8iklSizxcAAB6G3OUggBbQprFE8hFKklSPQOXbxfPPfR+OdNsOKYC+j
kc5lP4WXty83xk3Gr3Uq1Zh1OSlg6j/PRNUtzhPSanWhWojx+dSVjVAHvMhn+/oM
dsttkexBczHtFHuKgJG+vCbELwHNJEUN8vlIZKkkI4yGhg1iAJgFkXkSMnUGZa5B
96fp3eT/9T/kNPtrjEb1rT0halfL7HmAlLE/dUHN7SdO21D15usFwkEJALnz4b1t
qtAic21/6PJxP78lfXi7E1tlLTBZ9kkRQPBkp41xKau/JRYsPyspOKcWaHoBtLY6
pGK0JRQEhGzf1K/jJ+zqyT01RhwctCJ21SZoCQlc2Z+0eYbMph59KyukbrGLxxji
DtxcKydZAK9VV66rm5AFsUclmHOQgw8oohbeh2Tp8UF87HFf8OntnBRrUik653n9
lEZgHColyPWIYWQDKKucdAFh7TxUyy7GIkJvhw1g3Pu5AbAIB2xUNl2OdKdMMBGk
6stoqPMR3EX0pu/9hVD6/WQT1QsqMLJi5cDHt9DYB6WiEWr4P7iOQBExrMvWZFmX
eSSne5GNHRHvt5iMSGuHF4TR93tltFK7cytbwH52AP7kwxy/lFff26PZVjLr6/D0
zdCCF/Ze+Reb6OFbAEMGxo+oiqnxgQa+IzJwlx7ke2+Z2I5IM5YNahc9yuP1qlK7
gV+Z7oeP/dsETPAovnkVROMv8FtcqpY0ux3d7sxPW0zhc2rnbU5W10ZBDRjxCP7r
l9JV2tVlxI06C34JlQ9Ah2FdnLdMDpLWT3KdxAKZgOaYDwSeTKM2jwkMjdzTa9C2
DHMA0xYPM2zBUO9jirSmg/lqYsQ8i5kmakgcktE8Of+/EwJbtgiiuB3IMFfCVhOx
jW0toi1dUFaDBMPbhsYT2+wCEQgI29qJ32yJFZAh5mkNezI3fIRK6muN7L6WGUbo
pzNnpMH/uze7Pw9H2UhU+ZF3i+wbiRUh1NqcTs+GQJteJcKv9uuBWkZr7bolwFsD
mhVIXdvcIy3Lga+kIZS0wStABdVQDTTo9oLlj+vDKQbt3ZaB/EdCKft8vfGFrjQ5
aqDoi16TvCDwCtRXmLdAj9EX7Lwcs/erqnANHKg8cOdsgFnwrX3gtq6JzcDx+e1V
Z9CtDYpMWcNY3rbBjo4AXlf8tzB3ZSuM2Eps+k7lv/R+OrrqSXxs8rJKw6YPLE55
KYyQiflXc6xXgc44xhS2neuLGjalsPEG4fV/nY0ZMHjvQM/iU+J6DX9GWuq+7Xtc
uErEONSGI8W5YJ1dTEU+10kpw3aK4J0zfgiZWX9X8LoTtwIEjWunTd354Q6iRcn9
iaidwsGxcXIqa240wK7gPyuDdlzQBvCbhfD+7/nJ5zvVibLoV/msZGG/OdochAuk
eIV/AN1w8LHodLJEFm5p8LzC28hC+qLGLLoZv6vbJsqnXPOZ/llwfX8TYGBMwhNg
F42BnWUvwfOMPfov1N9bLzdF5yU6NcZ34LfehX/29C/xT+RHb5/soRNfZObyc8yu
LKq2aqiS5vWRK/CiUsCGoPY//xXXwcxEkhGFXcC7EZPEq+KsJtcEXT2nEt/hZ81z
vjNA0nFOCbdhGR9JXtpNxJgEKG9qbUOARmJN73ITNp8FumGfJ8Ury9dgX5tfrdIK
dhmlg/gYrBhaLMQIURpWKxVWvu9UGNVjeHGi2GeigosCPaNjmerL/0nuk8qYH7FK
TzX5hp6iKbaQf11P0K+TqldT/XlS5yPuX7sQT5CDy/VBAEamg3ke8pCuskggvPKO
BP908hiyFHOjLi0m8ICmbTVxpADk6HAwNdCd9yolr/4O/IBG4BuIDGmMULTKGWqn
WGLcBWTZgMNZC3cD4crJC3goV7K/bkeIh8bxDPOv+VvDnDH0WDHU/3WcwKQa9mGu
QVgYYIjXUdjDA3SB/qnx+F9nkGF1lHgIX13DNfEQJpX9E0TeivGXi7BcOWpVNhma
eeea4ey3UusIpujHPpwI/Aady3gcoCM3i7y8CXBrMBYHBPsx4PDnSrtdjdW5zS9/
YPSmUXWh2KGjQBY39tnY+M9NiU7qdoFXwUYKh949LmuzDB02fSLKLdvT+7RKIMEE
JJ09DwHhJcTDV9ACxR9xujGfucFWlTyJ/pyW2ckogBcTEPx5oeejxUFmLKV8OuUF
rfGZbO0lUPWQr+K00Ovs2kP4YMo6TeB7zI2GJ2wBX5htDVUeK5yK0aJjhMBeou67
aVKXqSikWFMBhneQZI0mOnStIp1/V57SvfftbKCgU6y8yuRPRnfHlhJ9iL73Imrr
f4TR6or45JsRWnoW06Vp+kgrKObstJGBQMCTdAVloXM0GcfaUFObVgVYP8Zt6mLY
1syCMCztipvzXSk63jPc1/5YMaFQ6gXoPhkjmpc31XEeIPnutU4ZIvgWLMS2Cyqs
F8SiROzkT/i8FRuuUjyG0ODuSplnNwsZoigAVY8ZGERrMrzPIhHXjF0TFGWrlYCy
q9RRat/v0fjE2uBXBAITDLwa48oyaYL9BJxgmkzpcMeznaHl4N6Z0rE9fE1ndtaU
Vg4FrzYgSdKZK7fKZFDjgG6vt2nonMgzA7tMS96dYk1mAzxG3x4nRbOesGV/juFG
+mDPIgdFCHXBJKZi2DSbmX9ayKtsKpUwmsePweqJedVlzhN61zXC5TzxRl+ixqHm
TY6b57b6VU/juOQ6a9D9kgsrhUHANpd1P4lVQIU6cuV3WBoAd9R7se3VDaaqOczC
xyFDc0S/iyOTLb7XXtG3EmP+xLmWjQbZNEqZaCSS18MKyMdZwhUrQw/McprwAYRn
twCiwO7AgCyFVi7Q3GJN9VxEnm/6Gm9iHNyfnh3sCXLWdpL957c/gBUNqN7fb+La
xeA90ZrzKlRfsKLhRCtYpWd+sHV2XjMcf24bz08pkb2KdbSILTmgmb0s8ebwt36w
YdmKEUggFRm9t4PPJWcP2cx73ZqV9sNqyWY/gLWPp+0gAzvGdBFVsdaMLHhdwfxs
R0JYnvrXf28OGxNK7Ayh3UFveHy6L1qaVGwKIAYibu7aQUt8JcNZD8pCjApjcR4x
xAT6gKM3ciejAe2053qaKSSbHCzCmwSXwo9B6o2zykFK7zDhjRTkPAPNTGa9VwBg
gUZkHv9j/DOjWDyY3kzyIC+IIx+UtiyTCJiD9gxyQRuWdAzhoMxpBykAxyxhKJrp
A/I2VPJLjZnuD05RZRDJA8+D7OahkzQSQcfgA4Z/ywzngvGJe6IBxQ8ZCiBTTFn8
fzQJGFLRWhqLCFkR0awfdTRq58HupSNEnhA+nyotNJ4exhHODmTHskP5Vdc07jlW
sjAcjM+QdA7DKR8xb/v81OV2otvnnGOAL5VO7rPUcAgi5e+CyHVntA8pfzT4cnRX
dOx3I52dZsVbSquif6Wg9k86lvd61CslTZUg1hVnnqKzPOKpYuL4oq/fay5INuXW
uKIWNhW6N4LF84PW4cCiYR1r81PZXBuBgO1wRPzIr86kvtVxYbMUyDTorqki1lR2
3LDp2ncQSA6+U1auJ7PG9KIxqCbqt2RhRu582g7+Cq6oq2Qms6HeEBxp3c9DYheU
kmLt5bCS0vLeeCajfcmc0k9WKb6czXj79vno7PU5YRnReQ1VDgKIyvvjUCzYU2s1
DZqIrTsdrYNH850DormbdvI/qKuuwzmdoVxlma7ynM5Dd7pj/vhlSFNtt4mKiJZI
MldzusSSWAx3yl0kuvg9iDryt34Ekd8+QXuIa7FVC48GZK1mL00Ls+ATwg6NsWhr
LkAuQiTzC3x3EagMaLbeOeukhCpQ3QniG7t2YEY+jZSheRwVr5TSe+3avf5cQ7bt
U+wnCnh3MVdkgp79iri6Y2lBQWOlJh93XOxKUvFbnKw7qPNvAnLrsarcv3tQPsZZ
h16ehtwgjgJ+RRhyy8ZAaBi0NxIFVjaQfFXRjmvbgXaBytBpqixHXIczafF+jepn
1EOXVcjyCPF+YHH1llbg6QQos6AiMWyEFmbeuqYfDkIqKsHDA8VAw1RGSkqiKMlU
ZsJpKtjefz41r+YxrgPs8jzYTsFD9VBR01XdVOxtLDJwOq8qixto1fwCtyc5QDK3
E4nMRZmt7EwAw9swQhwrHkRmyK7Iixn8eYCbigVMVZBrU4yQF9fxYg9nSm90+GkP
tXedWHLJu2vNKKUZcUoIPkl66suvlHjU+dtCsn2lY8U4FHJaNRFeqWyRGmKnJ3RV
nMxaxz1OjJPZ0k54Vc4uu/nf7+faJbytsLaMRJfZpo0cxRdJETgKVGOTM75IsjNH
dinFoGFNV1weUVsHeyE0q8nFnWg9lx6V8N8R4f55xpFIwMql2Y7XKey136Z9yAqG
3WiBBSfuhaN+ypQvkolyAgYcRTZX52JcldyQN+138rQcdddljtjA/M1/RqSqlF20
x3RCKjIROFua1fmnsErRM1LyKDZ0TfO2aL9NuOci0dLfSu2q6HIotuub09aUyYzx
j182cycOSG4c07THA7TMjCmoKVY7NMWuj60Ad7epOBo9RcQ1GdTkqpYNJ8TIfnvH
APlkphgg4eTSHxVynrPY69FHitqhKM0yNYr96P1RJ3M0Y+fQ7U2srUkATyw2iR6Q
BPRVkdwTTHxcveE7blwXPzQ0Itdhcr5wRdR+SLO1bvnyE21bsOoqmvfvmZ33kEiz
5i68rKWIeYFju9Q33CLr9d47GNlkXH/X4rKtXMeNCIptLaHD2UiPZ0Gz3thwX78v
OIhwKXzQGeGMZ/85R8YgWfIpym2NU2QWdLsU5GX6R+y7cJv7yrkG2XkNOJod0inh
5gX93shu+a/JyTSrLb0bD1el6HBTSkxTl/KnENHRPGrCPe0cr5EmC7axjGp+eINc
VG9NZgowtfnpuupSeFmNZ/aJb1yY5gseZ9Ct1Hh1WZphXb/BKOHhiMdrq11fnxqT
XsWvWMF0QurZDGUcY1gwIXM8g3Kw1WLHZQZzHPv/SQ1iZ75wVT5ts4/jM8fRObaJ
smolUM4z088APCU2pXZqSrP+58M5607B1wl4jIeKwXMqInduyYJ8wHZEUt0GXrZ+
CIVD3J2ZLhGplumCo+J2m9Em2/xnvHvbWT3leeuqMTi5bRGqHXxz0Vwp5qZ5FuLS
U8xh8XfChum6vaw/2sb7JWmLytX5cNCoHO4uqOoCxc4Psx6fpAt5Ox22dw2NEuP5
m06PCeFGohtzx18Unan53/IdDLkFMg3LyUp++/k6DrJNPjmNNt61862MaI4uPD6D
3rWmj6w3T4JugRarZh9auyygNXS/6SKtOkxhGMQ9k/s9t1UhCjC7j4pivuSBUp+K
yLsGeYe6KT/EVoYkrVWuLMRE4QaSTxtrtD6Jwi1bL5pzCTYlVhkraBTeXUjwD9LK
G5R+SUOrSoktGWvXdLzjw2fJLCSXg4UY7FqzOfcIXRXHZsLrCAL2YJdhINmcuv1g
JK/D6eNkzQjm8IfRIBIUCuIA41GPLbyRjqPP6iNWgkcBB0mIH3BlSwmKV+EprLg6
S1BN9zd98zMlH8+LmwB7K35OlUr5AyJUSgH8Sku+QDVojnSTaWpK2JMBUWfHp3zB
+ntxUzoHH6hPr7Wrovu+6sM4BeEVK2ZYMASoIyA+AcTXm1pTkFA1Qk1erHtLHyIZ
djskw9tuwsBvHb6L/95+5FuWus+vnuU1KuGVcQO3jyiUu+FpvBEiZHjhL7W2tmS8
VnXoPkFgNVWamv+HDW7CQO9plZhXP703JyD4g92er+ndBzaFgVEcnDVSShLkIVyu
K1ssnrNY2JBCjCuwh5+4twHM8+3i2ccQ1FnzNrnTaH9YckFdh/jstFp4YvK4juZ0
P/XU4GP5ljT0R1ilH2gTjMqYffdtrom76uUDOPXtKhM4BwgfD7CkpkUP4OCnEspc
9EDXCOADbMZo4i0LstaJHbx988uOwMu/o4okJ69w0YqqoGIWyPdPGmucIfXL1fa3
mQrjCHM0FAmQM0gn0i+ZlJ8OAJ0XYIF2lT/t4GaQSr1sxA+KTCqdHxhJMKPV24An
LhAcgC+OAES//+Td1iI9UOvRK4iAg8EB/sbtLitVKRVgiUX221hamRxPK1JffHTT
nptAh8LJej/8z5FBsjxFM9wnuOUfLSOju9iISi1tr4y+9oFAWuWZfr1/AShdyNOn
YNqb/GxR10tE9Z4tArj8MC/ocOYw0OkK21WI/AYWXEeVUZEeWnYfm4WDAYsX5v/q
OlQLhNpl4+ywY+pSJcaFBhKN35qoRRTv6FqdGtgtc3Vhy7dOApnmBO9w6uwmFYHX
ZRjEMT/M/7IjylCdXFLpqPONpGurlInScmrp5vYpPU18pd5VFgX71qIWw+PKLZAn
gT2/CiYn1uUu5mqVZ33vCW+M86EKk1fgj1zsgRRbERKzDErRWdzaF6eiKSgKNypO
6yJV1GQ33VqRmioMDr86zqJwHBI2XgR1yMUD0zFbafTvnPmk8Lvm/7tPHQ4laOEa
gLQgU+1quz5LXJ8efvrLKRhQvl30B7+08OJQvOv4/JqvzMXXV2u+gZsy8gN5gBaH
PMtS9dyKRKlKiMRaixA7kgn4KBjlcfnBjDICBpGCTs6YIH0hQDCHNhuGQbIE5Xk7
D8N8/a3zBRu4RpPQFXM2R+2V1InQ+yLhKv1wgolg1oMVRENBBKIqtRrAGpTiBoiY
9dRXq+u+d+MFjK2ZH3Dwlm1SsgcdcWZcZaHk/+kt3LMeZrQStjJ7pzvDdPSAZMGL
OcqYqOW+sMSC2juvJhn7IBQREV8/b39hpN43NBGqkK//4VozEiX82b821MgVt4Du
fLPuzJoYmfc10xZ0GXbtK7eGdTpNBImHpmkc6sET6+7g/O9H3BoKyXxau5I1xl8r
FrPKnaH7bMEmMq4k1tjWBuG6WinU9IMn1PqZ8XDhwRxqKOY7k7RUdywonBsrkBNN
JMhbdxPZihx6gId7d/UKpXFkBHazpYuh+hginhFx5npSrzLaA3UIpTSrdbFuEmS/
Zgd5Cpo2DzMoTCbDah9jqsaXpsIQ5f1xr0uBAmUVQ4RzolRuvzZ1hdrSC6cYVCpU
O4X+LbsDXdtXsxzx9aNvX9XQehE9bD9puX5opwqQqXNkT9kewm+1XTYtgYXqJdJa
Mqa6vyzkgwSft+CAVnYzorVyY8DDqhLbNXeRPqBPFowjXZyP75qFkERz+QbJjxfy
EAC0oLkzhrwR/iOUZhG7lNMaRDjsFxBpx/k2LtUIT4IeTCVPsTYn0oLFeEBidbs8
JtyB0XmAT+mZFpD1EpSqU8M6dg1mW+rSVNBoJ4xvwaHdM7B512ycrI2u5gPiSG5+
gCKRrw9+ZLNpFrdUUOZ7SgBbNSNBxQ6NZnZe+EZ+aVhGWMYwt4txuQ3weOp1P9Le
VhJV4VUsPgu1UHjTYpHCPa2fh0LZpv5I9hKrUZU5ml3wS+4DE2WuGoIrclfmoKzl
n7bnUmc5Ohycimg7eZEyXRygRCAnkVGUWAmvgximu4h51y2b+vfxoQdAS9vYpBrw
Ba9BNe1K+LOkcz34JofWpVbapYhokxccPHra3QbQfBvCOEmnlhhc7JV4DNkynSPZ
VyDKWOjR/Abf7A0QY4+56ljMqCQV+IM6WRGCLD3CE6kU5FbMh46BBjm5PMJuzvmD
8NEXx+u601Cgf/fnO2VBs8HDrj233LwQQMNroE8ib7b5/5ecA0Oqv0mZbmFk0c7Q
hi/kHQm3McqOj8Qb+3IUOKrh2xyc7LvZcn3bKOV++dETT2mLpq5CfxRk76O8zDiu
Kqz9+GTE1YPwEtlt0+pMCrTHW3g67h/RVq8IRW/TMRVVpmc7CcD9lYBGJcngbMN2
9Fug5arj0uYk360kN05N18m0AF+YbPppdAvolrnqWQzyXUKOHP+/7UaFXTqQyl+2
0EnJo6U1yJfhsyswrZrGfcg2IC/kQJkYw8V7UQ1biDmWj2ubwGEBNrzhcQGjIozv
TD1YMYttzCgGwKxl6l9CoBv4/V2e0QHakG4DsAV4fJ+nb/Jv3PsWSemyzyIChKtr
60/zcq6ZsAby6zFqYmgcIvPTRxjfSpwqCLMpasxCH8hDbSzPmV4rHBwSqx+i1jg8
3W1zoZGhCcEmwqAKBILRBb/JQa2KRkYkjIZCv5WQAWMVIVC2Q/K/L41qKNI7Ka+b
09ZPEAWMI/CTgioUuxPhkSwk8tQQWcJqjwdfBgLMOiXZSXiIhWv2uIZqYVaQii9D
128BbTnIBxPJNBHcSS3AoYD2y48RtrTEZEoE4/aX/M1t6gZi4pCxvVWtiWovUz73
b3/ZI/xdEjuBApRkMMrcpIPypEYg8sqIbBqRZnYH038gueHgf+gKvz9Gf6vn9rHH
15fqu/Wt3qKN3yr/+4WYUL/3E28ku3wyae/Wmaxr3FXzo2+oii6FfI+9saex1nuc
PtrSncrkUxxZUXfEvlSr2q3MxzgZhc6tlWu+87bP86GjAsVD0OlpUxMCmpEQO2qy
ORzV82wj7FoMD7RfL4RdpWMBenLsBWbhFmTNVTMCsLRwnRDRAwi63swWzvC3tOgc
vxhUsHdHTfrqa9GjBjhihiiWWdfCByfg0ykdR0z67KHgy9b34eG9jUj9JRGvQbSy
zZj0FLTZZ1gs7fasRVf6nvDnh5j7n8gLdkWoDkIi55hinPaAKAZEUXpoddKE5LeP
W13JjfgNwaKNvlEu3kgBy4kSfa22VdK3zG1aHwcPI3i8bb9JC6BUin5TfakMWyQo
Wz7+5JU1kXhRukotpB3hAnNhKa8IxEah82GkF8pduYlGWp3nMFVsicClKuC0dPuv
JqW7zpUBUASE/CgOb6qtoKNTvvsiKrVFYFJfjoLFx/AJnYDhHEB//xzaQuJjjYDh
Sn0jZe6Fyx3+q+PIdZw4cym9ZmffkmshsStZrVUpbSkewW6edN66+Dk0m97/B6jf
Y3ou9bbnJzW1mZqCe50XWK/beTNgRnOTHpw/QHGVIbgXoFLECLhL6X2pTyPWhLTW
U8VvggWU/n1NN9pLzo8kr7i2J7kMzVNvhbJc5GkW5dUco1hs+iquM6Z/TgNF5lCF
5s8MJb3NyaInwarqpusv0TkGy8PuqJDT2WjE2gxNCNNaUUYHrlRAS9fnqvDLbSK6
PPpeOCFWBHVDzEHuG6Zz83WdX2SoXOqkwIhAxGh1Uwyq6QVuLFhb99eta6YMhl4/
YmiM/eYClXhFMomuM9aUFbSvbx7Sc2FrMMrsScn0urJpabqq7fLBOYEInxuGb3DI
l9ua09YjTx6krlmPUquXv8ztO1e0KInoDwCMJBhOXLthd+qnRFPs2enRrDrK3sox
tI8cef+UYC+FiQgW/kwE6D3obqdSFrsDPik725+gk+f1QElv/8RueM2yVezSO8Q8
tO2NaBNTHF6B6tr2B8Qe4mzqroSGjy1UOe1QyTjm63x8d4QIf8jojrKEC+xFpO1R
GHPb0dm4Tz3ifyIvKeLyhXYs03Efzrk3xvVpdqyphjMSq2yLWY42oBrrKS+Ok+Gv
pFkmzkxJZ79+fTG+2j/BvHcAdwG7dmHkLJ6wUUqHP/Hlj390hryYykzZmqn2AM2K
p+4yBUwZZ+oXksz1hJZx04CtjvieO4zL7oAxIPrjuEVhjulAe6vfkj01xTvFylgc
rcTPbjSNYM88dlT1CwsfDmi9pWjdVyOdty2+BEkBRuVS8Nl51y5qlbC3w4TeohDC
J9rro6diKfPt+y0aeF5nnh5VAWwaQWSJvgJb0t1w7FxeNIbulr4UrnZw85Tjc55O
wfBxqmjTK7lq4EPe/lH7bMoo1KW2Iuh5Gy2SNJt+iWIb99kZASLtNTLfSsLcUcIg
XDz4xyFVMBnMc2Sz+1SZOruaFathX8zhelA9vjKQRKE66PWIyhzf+LBNblNbXakV
01QHfR04WsqXFAMRq6iEYIA8aIoSbpwajQQEGL8GDpw7lDrl9kuIx9V8IJmZuI4p
xktPMJtV+gA9GT91yJn1QOQCavFRuAJrhDO5aChjsXEfhtW3faSf8IsAi4nZUgPc
a8as7I7sAYcvlX8bbZ0eKT6af7gpHkF4BTUolBlI6iLxix8lp7hB5koE2kGUIzdt
T8l5DhedabPm7voUBtG3/5zzEiQhmHIiBi5nk+m+ttAsQIVHHmN/IdLr9WVHEcck
RRpZjrhV43dPGNmwn5UhkcnZUTrqnVZa+tZGKHHthaXyarCOzI/NAD/FsS6lkSGq
M0L5x07BdC/xOgvqQ6UZuIuYSILW1jVX6hCrbjaFRW+I/RRRjdeOnNsoMSybu/UX
8wbDtV6FROmqYSCuWI7H+4nbC1zr5iXclPO2207Alv7hoi59lxiN6oZAIxKAZl6V
6WBegRWvScl8zz99BN+3+q8w86oAbn93M79i2YZeD5BXUQxznnPrLa4cmBX2harn
lWmW7gChZA/htUddWeAiy/G25AW/HNW1Sb7jzEeYzNKIW5XKLQRIL+R63CQwuMNz
uZrumRXqf67P3OvOfQ+O6xxsNb8uBbGEs4PwDM3XtWCc2hh0p5jky7aFPxTZV5mW
rhqdo8QmQIV/ZGoraj0MvfZDTiH0nGAUn1j8MjDBIZKOXvvGoQFOvnUAr8jZp5kM
vnuRL+B9L6B7zhRKT09vRvwXNT1PdiCVtSDgMltwP2x/rLUPQ3okWLNT9m7PoOHp
eHNX1oK/UCRGBFYeONKv1xYONx+DDC6zNI25L5OA8YxkPSR+Qu1zerW1BfKz41e/
leLmfPc68m7qyZWv4ndIlJogkX8K+ob249ENqqemN7/PLfHgXWnpIzS3cOHZsefQ
75r6caIUjCK3Q5N7PFbDCRXcrpymie9h4aBkYXY3fPDtj2wjqAVycnwriIoM492k
S+EY4goI2FAfTQSuyTqpbqj3AYqqkcGBZBmFPhj+DTQHKYEFYg1RdH5yx0ba67n8
mB0pQHeZe5HqnBOi5PlfyGrL15bFIqRMuANW4EonszA/FJB7pckQ2mtDm30VqXpQ
X1/Zb2UQ8O1r1H6HTb2/nE9JbSHtG546YWotiHxxLaXYt22spmkpFE1rN0PVuStc
B86Za49E2OYjbCuKMQVqVMs37FhI69v7fPHhlRZizYyFItsUSIbDmDRIztfGQlrH
UcuXeE3ehzXRXl3PRl+HM0NV/yIGr6HyNkMX4x1LqFBYzf0qkqXKY8sR+GCslFD6
ozA9kovQ5asmXRrtt4I0Kg6whBGsjnmLNBIFqcknut/4W6E9ABhlO3/99CQ+uQjZ
Ym4wpSAxe2YozM0ZEF443+7WDmNWm0HN76NErvxQUWITj5QIXutJnDFCs2DX0ape
mgd3KFn6sws7RyoL0sA3+HogPSGrZxlNNq7poRY9Ytr5AQwVBrxG+idCPARynfdR
CbU5SM5RIu7nf6Sh6ozPmHR3G0JSOAU8+S97/YeVh1KcTwgoBYpNFIOSedxqwKvU
pPPm/Y7FS05JI8/Z6VWl4KXDMnWARK4YgXMUJB0WIgWdfCvY0nqhZiutGii4NPEd
0oPT8nbYy8WLQNIvVaVYtLhWQ9MnGzfpo9cInUrBX+u2mq/WA2YxYEEZnTFEpNLi
dSIb8Dzxutj4AtPuxTWTJGPCjrRTqX2VFiLUXGivK131tOXBgicjQYsCl1n3XDwW
Z0+JY3ZXB97HraCi7nT/LAQsuq5B05clQKWvpWuOfOPBt2mGcQtBnsjLOoAu7bH+
12uxS5i5S5g0yRyMlEapISdakJKi6IiRqTG5DZ1Lov9gDDr7NVrXa916rkWARH9e
THsum4jzYO9ln3n2j2AMye1AFSErvgFNVvJXNb+QaQhnM3G3vZXhkfJl6rI8uy1j
nyM2S9p+U6+nsVmyn2fv4jCx1QRheJa8gmat41GGz2ztpiZeDfSesbqvrcOFJwZK
B5/39ipuQ14Hbt0VMc4DGhvJiZmpJAziiPdbm9GivH/I2wocFj4buMoSc6cPVTYs
5mEj3jgoAYlZIaMjKLK7jCojzsWWtuiIVBxfHken4JlTXXIJ5Hki8d+N3sztqZo9
DZeyBt+yEe+aJQ7zgsdzARlSrJKXsTCKkPlGvHDN4kyi6LwOgJ5U3hXHtPF7Kxlu
ChwBV64nT4Q0NYSgezLa5Yrb3iSSMfBgIBL2gzi5hasN+Ulagnjgth8B9P2vao3F
qBWQKRYVoHLkvdwKS6qC055bLQmFT+0D0vIpYN3q08GxJFecs7CcgsX4XhcUmGFz
91AJGBVbPwQWeMxjErJXqQDLEO3KinKrZ9VtrWG0LKskyKaYViI/QbmWu6YzV9nB
XM1T0zhHMw4bcsUDUR35XvJaV6+eagPHXoNnn12mq4VvycFbjS2YEl0lQ8bbRChZ
c3s85UQE5E1ZT3SMBdcQEjdE4coLwHUk9eSuvvLCy7VQxZeM/XB/dQb4IrUlVrYw
QYWeaCu2K7cbn8Ardm98RsafuKmHiVieI74skVMwUfUZ0XdUhpqmSBcfHO+OKw8s
+uvNv9mKoAyRckUD/qaM74Vc/qtyRQoSR/eooOO0Ay3F82jzJ30FtZ41u7d3cOXk
ujzWh6AUqxdF52kR/so7ukyKyad2v2P0latwRfh16Q7EHER6L/ozrxy4RT+c4yoX
3uSzVojfw2kYGn71JSa1O3Y/HxMSSiTGhoQMOXLjY9qJ02ghIcV3zmcczuZOeHvr
JiGYhwLeeDo7EaEtai0RQALm/HUxAOI0Sq2uvc8M6bdhGWmsBQYb5VX0CSbNboBz
l2jhKYPevAwluYzS4hrkg18YTOKp9k5rczMIGD5TWQfGi7w1AioVtuVzSFMr3t9R
NPnxEmiu7KORwg4Ra+bhSynCOXQvu0BD+0fc08R1C7BHVRhaupcueIdtyEPl5SM0
bRUOD+ZjTEdWqGEQuDsH3GfSN0dDpg8B38V+XrHyGN+2XMvEzGjtOX29hK2WwZKu
7SyUoiiPq5/Y0XCp+KtRBbU+OuN40b+YtOhvlWpf/DNsDzVEGeK9B6scaTAb7FLw
HBIyXCr/4tOMBaOTUFEn/eBnxG5hZaaEAk3klJNlpb2zyMQme/HoYKhuPxPq/6aw
OKZvvn5+gA+6rmPs7E3WkO91mYh5yptp+ewDwdA5uzWIOs0H0k5xjjQD8RYzmkZJ
7IMqcm7AbgH/vutBM2IvLm8Aq6JUIwIIRnH+h4MYYcqexHogPjVcenEQ1jwavME3
mDUv8V1HYiNb6/4pJqGnLtJj+6F1mUhy1JKaWc4a28BSZPTx6eg4lWAMzbxutsWy
Xld6yGyyWl0sr2xAaxLBmirlnioBVNIvb/xzIZlzxtMu/RYd4XC7g7oiiiSSLyGC
78WBYcO0XVhtEcVT7zP021WLtFRwLPbOkKZ6JeX02khCdPAjEninyu3bIzaRe+Ie
90q1uUIPBzJZox+QF169k2sMGeJsnu6f2ru3v2ogVNopiPvjjjwaEJY7RT2EL498
WPgt0Bb01Hwm0PF8ugWhVjlwVYwTk+wDIK6OqZSToZrPp2R4bDE45/vEpJHXB5iC
CK9IxKNzx7Z1Orxg6LoZF/ViTGDlDPdwii5yvKk9ctI6+DlVySeJpW8th0JNRmYZ
zWbPeX7pkzUxMNcso5FnhtIrHh0F7RXXUjmjS8fpBHttFkl83IDKxpSO+kuiU34p
lQZcxfzjGhcbWCBsFjZJIHsSssYz9JAHqG+T3xlNNn0lX3a577FpQlGsNwkGIFVI
UaCEWLz8Wid4I3/5sTUCSneVyN8IBx0+EZyg2YvtBxxnBo8LeWCyKfLOyvFWtqty
JTUs+bNqNtIW/YNne7hqqJtRMNtPgm2jdmrZayElMBk5FLXeEKvbs/+KPQMIhUZj
xatswwCLb/cyveEGMoFy4OMwbICgi+Rz8odQoNPK2gsvDy3qjCLc8RSCJRLZrggu
GkTnFv74/MPBRGY/gx3r7sNDImCrF+w7b4jpZ4FlTEIzLv+FxTRxXY0+QMjwIEbf
RD6gE7ka14dysfTig3Qyfdf0fGZVbLfgGkcodjojYtwQ20G9IckyDOxSihx38MCa
Pu5Z52shvph7mhV21mT63D8Oy1iXC8EQW0tvbbXpCnUr03NPHdQ4xTZ4gnaMHyr+
bPmImlOWO/uIL2Yw1mtvap6vEuhEwXBhNNM1Vm4kWTVaeRjRPGhFuL1mMED3PINH
6ymPk0vEOGguh95p8uc4z6JiVG4I8mHLQ84oGkmRNE1IUSZqZhTVHhkOvCsmYLEA
rOFItr8cRiV6CNiSO6KKGVQJj4ECJAsZC9HRCP1xysQdgqZ+Ts0Mt7cfnx4L+crB
aNEANc6UPcAVBiVuEvPc2x0at095p3Mb96GXsL2qyqAgKfQSPtngRbunrK0dOJri
k0SSdZMDPLhp2sYUXDStbR5tbLD/XKZHmhoL+nKGFqfXlc4EkLcUQfGzNoXzYUDm
QkXZCnilmsSjzddF+Yo70/n9fNEOdJuqMpZmKdO+pw9L3tiHlEWLciIesE6Wu/dO
4RsQxn8WIPVQzVnPQk5wr40NxQT94LixXTVaMahq0acNOt8EOhGI3GyLamsv8Kyk
/Yg15ug3/M82INk8ishzH/GB/Yh6jSGDe1nrcN5IK7oq+YLORsfSEubhU9BZSDEq
UrZ/lnrSy6PzEQWBfw1x8lHPX2BW/e82qR6pelifycwGr+oYVM469wjDahAehAdx
8D1Z0CHpGpC/eErn2uUdfCb5AyeOlIXt0VAIY6aKNFXO04vQLWElS4u6kuiBiWUE
c+s3wnIrC/dKBkvjqzTzeF54d5metNOKBkEIJ1VP+BpNyvrroD60v17OmNxCoXv6
8/jEHlnJNO2rimOfx2jx2q8G8UHsKx6DcElIq5u5GE8Vdx7qYatGIpc72kYKuka1
xQOZOvuHDq+vZtF2LFn9EQ3/tdBJ+axMgHH1jACfCUJmY/B4P2RT4pZ+DSC0f4JS
n/YMgHM7FsYfM3pvccY91ZC6b9UN3587grIJrf9iQMiKrOdKS3MqVpMACQO41SV6
YnEd0k9E1+UIZC3cUSZoeo2Edxw97KHBucVNgTes6hrI+Lpuei9Y8AXJXRZvqHhm
aS1o23X36FLrkXnJ82ZbO72AUkUndrxX2D/T2caso+LvpbqAdJus/Lz1Y7kqiegg
F6YaszXQSMKa6WJrhWuPHMxddEHDvHqbEVLn0/5WhDuc7/KHfFPEokqBie0UUfGC
WOqPoPuYTS4EKN6FjWnkO5jVFodaz+75EpLShmX0Lv1MDg44psGisiRU2KJUVLLN
ZHihXGc3Y2+ack84pAcoJ2uRsi0u45tKBhddb+WeiXhM6ES3LkKz5ON+Ooz8/2xN
pr8G6KUqDDvRbQGqH7hLJ6T/ZNcnL8lbeGxkeVSyxflSqqa8PqJAjIK9+NUz7mFZ
0m01u2nWmjuJ0AOTDBw1oNX077UCZogtg6YmtQgkMIVq0zbweFjfZH06EULyLYK+
wf9/EQ1pquwJtyy+P8MlsbTeQJttnfaBsZBF+zS6U3TdOoOQUT19R/Ypq8eF4VkP
RFpY1bT+9ziXHurR2FfyUk43UIplc/cgBcKafyqYGA6sORPj9W7SrGzG7uEr8eTZ
/+9h6udPZZPwP3/SEcvYa7ImfprzcM+uN8rEbxw2y/WYDsZtE/rgtP//edxHfF5j
k1JT2P2x0YPBG0fr8TLnJWyEMXAaXB74XfBWdkByMk6dj99CYeYHe/YERFLenOpt
6j4J0A5SZcFF5ddiqwYG4JDBnkj64GRl2BdqINH9KO/Vw8tS9IDZJYqnF6y2FG+s
M+6lDSFQRCRV4tp99J2Lnrf7mHXt52J7KxXLKdZiq/4GajrobC/E85Ioon4Rj+ye
yxrqRE+0mzOwT1X4tZ0KMi68M5ryv/ExJBO7cLiMMSvuMHhNNEFUJuDXrDABpg0v
wFJCS4CNeD39N67fRFxIV7mFAGww3WU7d4U6CClxtR7UGgrYgB2IliJ3OJr/Hx+k
DYKmmParku71aIcLll5EUS7hst03By4gYnY1li61H2yX2m9Q4fpv3gniqfFjQQGg
yZSz3XASAmqXykWENHU0FUaSX12+pUyQnuXDp+dq9qnrHnNFwTlFI7zd+UDeNFGo
qUKV3XGU7CBTS0pNpydQ2BnRZxMwqSb8+Rc4Mlic9wE1HbW7vez2G1WdSuUW1EfS
Z4dCcNKnfJwS7TeJuW1qFgoEtCCv5MsK1YezMKr1iarM8PRf4IW5lMF5FBdCm9C7
t958gDdVXPw+tI/wIoZ0dA/nkXF37oV7PYFkrWB5E6LRr6xe4rW0ffRryGIGHDxu
lilVhwXukhu+a2A2A7oCJd+4IjTWSvbYP8vlbvM92pfHuwqQAU6xEjPBBEx4E2gV
bireiHtWm8UbIrvdWDI/xd5dLv7fQ4AwOKq2Y+c+O5hPwKSRLtdyT7mDWZpcfy7N
qfy13xnzpxwpxC4+9SHGQ8nHTvxXT10mOA014bGlwAU2I3aMadqVuZducmdrDDqj
qODxRuGi5ZpE1W7r7VyeLNyQYIAehkwMrnLIAkjiS8cUvVVxloF3JdIKWUlaDyi0
viRpVYV3oOmpO6BDWGgJzxlt7I2uUsVuiQ2eDqm3soAkvy51cReBB5JJoCu+gp8z
rbbuX8+nftHEbM/oXZVWpY078oDgPA1hsn6qHTqZvVvRuKhAP8XXqQyJS/ksFsqF
Adjps5X6bQBrA9zm/jrfUxSnFXkOihLyK8qtOwyQ+AYo3p4muVLrs62XtTYfaMax
SR3d0yOAsN8pv/6Z6lTM56dFW9HeVWEXGG9o4J5nKb/Yf6etvRCpHLQtJurg7Z5e
SkoV6ghsIwE8/9C4S9E5+3a9HAITbskVIR66yUMbTTGswjGsePsuA1I+sXIi8byc
OyucGpHwOXIWeS9n+qF8AV4NFgK+s45uBKMoZiwGEniOthakLvF3lN1zFR9Dedab
g1lQLqzx8zg+iNhA6+iQUPyVo8KfkzvZBmDjs755Z1uH/YMLoh8tDkYRe/T1WvX+
h3WolnGcltafMoHE8Vbs688Tnxi5D1SGHMbzVU0xRZT5uJWGLXkw/0Q+hMVyotkw
Da69En6gUGm60rq3R7zjouD6LqShzrbSik9iaDIM+sC1oEf/0J4U5TAjO3oAuojQ
9kuH00JBWHRoJHTIL/hkTH9oVRaK1r5NeGGnKYg1uSMiip2+fOn8D/Z63tJhw2Ns
HcdztUAyiqrfT5uGemrJ3lXCbANW0hQwLr+32qrm1xMsVOGY2ZFWUOEoG9xbmAKG
B6FBstg/67ImfjW+zTl2TOFUaUczUsOnJmkiIQMDLNyNArXXDHyqvi7kkpISOnau
sFEP4P0NyrQH3tUm/AL4dfdkjIFhVNyG8lEWGncj1ejaZeshxqrEKTJJ0O60oQVs
G/C9hAiVyHLMupUgQmj7gSrgt+vvq0C4PLb32wvqmZGQmoDdoa9o9gUfYQtxzmj8
E9TClJUHZB/gPBuwlKWwAUyhiv38AfYa9GYzQLXzWzmkr22mDl3u0xEMxaKlP17/
hdH4NGEZwGKjlLfEzowHyyKBheRVkM1sS8DTV+VFAMYXVbVE/dn4h6FFIgPEyqOG
5uTfzNFaELfrf0V1B5mszJFgzWFvCYLKuBrUs5yRbeo9c7LS8a7fIA56gRWpX9pa
PXlOtc4jVBMM1CCHkcGQrXj7mgQVvjnlmXlCEYV8HJRxu/5mWg0SfTQYSnaRbknT
ov9Gl5WbtWI/gMXbM58HphtE+yf6nKhCf3K+tbiJrB13QjTx0pALOEhpExESFSMc
tKdEnPkF5fIm/GwtyhN/ohivYbbXpMlJi4ZUdeNAlEkY6doZVU3AJBVWAz0I1+jd
i/IjGHYAL8cpiOfRb7lHdQxHPSfp1OBROZxOAjDR+vq2PBf2sJAo7m7vcu2Asdaa
jgqTU80Z5TFXCiGQ/uXl4+0/r62Ws/sm7dkgMQIKt9vYlraTXEHDNpGoBLiGf3yI
qweQdqv/3trv/D0/ztRrxKtkrbp047dmM6gXneOXMsJfsYZgsveJze4kTFv7qj19
4GjfpLGZvy06idj5YmH5bo7vCLElqeaUR0Gk64D6RTyzixl4JKrkKs3XDSi20yRb
CnZqSSv6UO1SsBQVX9fcsQpZ5FpxauSfNviqDF9tsHMqTcpSbF2RdTndoMx8w5D4
bEX/dZPvKxEb4oDynCBj9jkm5HN5lDIw9t7MwxdC8uD39YIz8QcCkd7use/y4sBe
/mOHfwTGe8rpQAwb018THv6+Bc7fX5XCCInEkpIU9nxB/as8KpZYudoiuU6hjYae
IQYvRJIv4et1hb1//SPa05Kp3Sr1teSPKiRqnwoPaSCiHUQ8ba+iqBWA6OHs6CP8
mFSYcq9Znd+B74T1wulMvMArO+Ya0TzCS3EHyqu3e8BIeKlCEIV7i8ofR0CjSSTp
qeEaAzImPhPbiHtD875HjApE1mPH/jYSR0nmXu3jz7iGJRma84EWM7oYjJJdiyFw
+FrSu+rtwAiVSAhFC6GJqn32FZuWt4A/iBaZXQkbGTkdJF94j29mWlJ59m8c0PEx
VVEl9tV9uQGhZOZG3QllkSTO1ey4fQmqrYgQMbfuZbpWGz/p+k44ocRhVticiqoL
nNJ0p7VQspSO34ESxy9E780F6648NUHgppQxXwM+O6EsIYJisY989ypRfT7ePjfx
gCJ13mYA4r5GCgrfdxpFwLtkO+13afcKMWsALYWdjLPDhdFYndG3xMAVpX8bc5tw
sh6XHrcSBJ5SlOAGPZaDbpApdcRzUiMJyjDKz5z9IZHy5kyWT01ao98csHX9//Jn
tI7AauTai540zfxRBLg5rwgsEAkzRFvv84X5Ljq6W/amDyY2AjheGOI+VEmIwxSF
z2Orr2bSdBDgLpAfK+WhFIYtoi8AyX7kN9G9MX5Ks+thnLz44IBlPY0pKHzrRlGc
3cXJmtowO+62GdXCFb0yx+IYPL79wQbeR41bpeSzALawf82UuQVV+Ez3s3cMjcrG
KViW536bF/MJKxiRphrEsBEOe4ni9YGBWOd3NhPHgLFLNRAHEzO7YLbKpEHlU2Hc
81IwWieZKB6ZFuRHAtoC41Gh4Kng36cpKZfpPS3/B6LZsTI3XPQYgc5HRU3yNyF4
BYWqSjgUF01tpISMxd77824+Si3z3MG+PBSssCHP2ilGk0WPo7glLVZspJsuVjcS
onGUwKx25AfuoZK2Rs172OFE/4bh8fb8MN+uYoS2Mi0PFqnG2c3A6QE/Ch8O+z5x
6xvgTU/BAiLW1A/+ygzt8WTph3HOTnz+psoot46ML6e7PKXGRGYY/gOJBa4xiCx2
CNJGEY8rTcXzI+qXVKlFjfkBSwajmZgqPvfiW81Q5uxtRzi/EkUuZ1I+LEieAFEm
4Q6I2EHZTjP4Xk4WBbb5DvEvd9niENq9W0AyQchHR6WGTNbBf1QtBxufY5pOE7RK
Vqgz73jflGFtLoX+OxysSXuTsBUy3vTOd0GRwlXe2hoxFHNKxA4RtiTh7BfHY3P5
j62bgHn+zvgd6dHx5/13hGLu47q+Y/A5PMSGA4qoE/W+nCJeuPHyKZkYU62Ee6DE
eWU+gVGqnTu73BjnNCKN0BfPyCck0DjWw+tHXQ1XKSYMYtroucdy/oNlgDWkoqQA
xpe2Pgkq5Xe57KC4ZbYxb1GDH7Xtz1XVk3TlA8+sOpqsBblQ6zfQ3XclVtV4cpbA
Vb+AJ+hAdu0JGTmwtE9qaPzRIJpOKLGuzAActbHpFdyrjMm13LCyzrz7tIOkd+2E
WbWBZnZTsMbuio1njwLw3cLRE90arUIt9Wzqc6Rb/+q3tdMtNuct9aAgG8TS5YoB
+v3ZFeUdfGxhd6PsxTCVc1dggnyKkdc0IeEJJ6ssYiCLtCopPa2r82y4Pg8l817q
Fs+haFW+gAbxDbxuSwmZmTWBZIzjEnQyPn1YCd6Op1xiGr1jbVpqhoVBDi5D3R1Y
DeJrwFnEddXQUgbisL4ajdlPxsUdu5fcy3pikmtTMbQMrRavayJJjCbUZgUHV5HW
NuTLbAZdJBUeGGzmzAGoVlrOcr69mA3Vu6Dh7hEpxXcqwBhI/um//NSDM6mPl4NQ
42VOUw3zByNT4Kk3IyjIdzu/Bw2SEuM0Yix5cvq5ugdrrwphru5fGl82k6YvLEDH
IKFf7hkt/J1YrT72p8hv0pra4sIcgbvs3q6G+USj3TW/LboMv9x3W0YpKTgE/OWH
vVcnysful3Lme2xQYagizmlP+ktVCfOa9eH5PBfQtV053qogUnrQBjlQui9Be4Le
VCt2RBicvvQJksUKIutkZppSD/wmUtrgmyDy+CfQ7r7Eov/P9OnUsfKiy4lzZUVE
l3aZ7ZphchwCLNALcIx+50QIivpX/Sw2GasJux1OkA0pp3+ilaGOYmZhLfWITIJr
UonR1tCo6UFBUdOUllyTTA+nkLiVm9PLHWVpRiPDmd2/nQ0zSXZa42CKHv95fChH
UGF1Mlox7ZMn1haf9fF8R0h5cvE22toInNxKvarcj4YbahFmVlQEHcqtvF9WraMC
jW1+OXAF+atBJ4EOLH4esZD40V+0xjHQPx6CccWg0F8JSyhA/IszI+qk+B3J4pmT
ZTw03r0nywGqoRnkWIoSac4uBFMi9heruUu4wO3S66hAmF3OE+w7cafWNoVeFtht
2Smfti+N1Wu5ipigJOHyKEG4m49lBEeSPTjeNTSokkxcSfYk/rXfQJuQ5EdUp6B+
F3PQNoMhvk4et3EFb1+vXiccbrzy1Ub/wq9JX523mMGGdO4rtIMzYLruYrticPkw
AO0vGpBETqgy7LOADNIGYg1TzNffDSqQu4Gz35xhAn4XlSVK4nhYMwb9ymjReJe4
+NCnEw24pUbLfJtdYBB0ibvqTh5ZaqNsZ8TyL6dDboWtikIsLHQRtyIdVGtfeKTU
S+cVbR7BeOr7KJRpQkqSlcp04eoUPJoqjaaKeaJxpo5CjYiaH5wmv4rG+4umciqN
5Ue9YIcB3/APkw5kQJbzz7PFNknj/mpJuDqWiYlaZEOdKgALYcvQBKhOFATkpa/W
SWSt9uCTKNRX7Q2NUE+SswNhOJbnPp93I/uePd1W8wfN6+Xw8DX5wFNWyUWo+7qy
NbSzAoy7LYbqvOr4qA5JNwJBA9BSXMSEWtt5iXNrM5WwhpuZr0UAWwgnOCaW1OWF
cCL/btb0lxukPG/iBdDSUIJXv5+SJtbHZXfWzQ3C/Dzi06H9B3B+piwkiRnt7we7
xjmGqBI7OQrkKpE9RUryWB/TNteChZuK7x0HYH+Azc9XL+TV0YLZggATwoWwAqLm
JrEVeOmWNiq2phIJrEpVGiLewR7iGUUS5yl+BKQ5oTx8fVRJQ417+5YHyqPiSyO7
K10ET5eXoOHg5qlYeY1aU85EFdnle095Yv4Dbb1YKiIl2iPdh0Dd9AaNhUFjGJ+D
WNCZ1sz2Y0wiUWkUHp+OCx2u8qe6BCk78yj0wu/mvZH2Y1+vMJHF+BVN23dlMrRi
IKhZaNxjrS/NSomDVjvmUBJW/arkzAIrmYn4B7q2GSdKmhTZF0tiHsS+em2xgo+4
FsWCISFR/a4gC1+smlQS8jEiNJ6aYp+ZiixOcOMNLfxMzNg7tnWm1Kgg1jPzTnqR
XbLlZrWrB7qqh3UbKAQF1vIclkFQEWaLeie0WHY1RziAdsagXoESAunkS0LAJOHI
m28Ajw7rcibxg6ufsg5IqxM2hS42LG62B3E0IklReglPoS2Dto6OeFjvWHe2BMQb
8dpgPsAIhFIb1jIaKVPra8DcSa1JEosOWzvUA4kiX3Iy1XwM8FkvyP4KgmQITSLh
yqVGOpDxLBSzI88I5wvu0qXJ0KIBP4ysGJqipkwFT5B97AijymKACgscZrAnOGm0
ZohhOjwNo2XU8bjz7y2Iu4lNahPtt85ruoHItL4npbrkNV/acI/97qMj7kHpjtJe
Pwv6Psaha7t+++N9Z86t1+oAX1hFvDJCn49C9L0TMsowQX8WwR+oBkfkhlkG1r3s
nlS4iyvWhOwFws+vdtIDhEEuIcq17smA04zPUVkMEL/+NgJ6HNbQp969n3qUEkYW
T6S8hNm/whML/KsF2J+smA/0CY4mnAp6VHQzC/+LHrFbTZjsVnaZP5/HCWK+TVhb
S62y2uSuxi8yxQRnl9NuN1JhmdC9QcWgC1S5ukJG/dduNRO3U/yO0FtNaGsnvWBs
vFCN8xDpuXvE5igwXKxjGedJ249TwUFQJerBuzXhtbxAUU34u4Df2kKUX9acbE/u
R4rkafQQWoG6RjxwKRbdNm73/idWDng2Ferk30z7ci3QajK03GRfvF1zEwQKoxqG
jaG6kpr08Fk1GP1Nl34fTYtglHM70c2uvJsEe4FRERelEZD/2/8icVZwgrcWM//V
rGQEObKHwZPo2GOa2E7nSswFgmxS4LfjY32BY6GEwWT7c1Z8H7hHnFQMrxXNlmBr
2QmEZfL7buLHvewjKHMZHWl9I/GJw97ve2EwDX5Qf5Yt+LsGuXXxqPHpafjD61At
yVu8RnuoC2BiV3YKWILvMu9XFGr8YNzl6SqSvGx8Krnlh+dUyLhKJl+HrfmopOxI
yWUcLY+EXYqZ+NZeG/XaIv+i/Z5spP6m4dhYRaeez4tiARrxGjPZqYHtBZm0puOG
tg1Bw6lwqQb9r83WE4xDjZCM1xS3+hFU8oWnEJkMDsyO8/Y3sG6ZJi5ZSpY6dIGk
e7uF1a/OkOrptp4pTjENyDBvB9qqAZUdnO0/8d95dMMBu7ttXm3SmYu+qojn5Oud
xK+J5BLVgl4zIqqE1jjhxx290eEp0zeXUI9W2nw5WK7Pn55zQr9DIcLjINuOtwpY
e8L6pB7mJeKBesBMOgx3fLmPtbs+ZagTom3RzVYVbeCBJB4gCWiwg2saXakRcpPb
SfcMwFG9MvpSIG09gY+WdYrha6hNBeVBe8xXG6FEanpRuBmRx/cCoaO3MfDAq9FN
juuPPxeIcgCO6aEb0AHiIinaojlTZGHaje4O6senvNZdKg/LgcpoAlOiD7+937in
YKmNKnyX+z3ctPyClbB2qlwaYkLP8NFJuQAyqLruXEwEqvt1LhUQ2eNJCW2+hFEh
TJSwlQu/7LTWgMp5VoA8bJYQlV30UJQ20BsufNvu1uwrzmk2oooJsNFBIGdgilF8
B9c7mGVld09jwUU2frkRO7lXyO6jfwV3gtyhiIQ8mnLRFRQFph83R/gHLzRnzw1e
LBp7jU+f8tfGNHIZP7Qp8ipgQFgMYsF+23Yzx2N03bkLGB/9PfazxTCnOBAsJzcg
Vwr0nUU1SyaGsj3C/6Bi3DT0pu9HYpROF1s2lBI9L+lUw3kBDCP+zL1xpUfgelx5
eHv/VbTPEm7tANTrFrdj+D48y/tEnF9sJ1+9JbC1SETgQ+gMmOUQ+FbugC1n2Uu+
8zUK6MoIzYTcJiba+m5A3No2nFP697kVwjCrIe/+0/Tb7SAOoGapaMX9K0d8dMp+
N+Ax5eZGXzkf4ynKERLWsWQ8kk8btRPdQerMYYPOzXPnrpqPCl/EZV9ZV73/Shpl
Xa/zKVKcZy2NqV+jU/eb1lDN82deODSnZQybHKNHRKzPtkgquU9N9l8HBySfn5aw
aR9+vyeofE41n18p5Mm9BwVkxQknlqY/gYYmIRFGmGj+6LGmXyj4u69ZAGZ4vxI0
Go+NDChWJqlEicTQ2BK75nG7UvafblVAu7hHlOOl1zzKaw4+NPdhg3bL6TwnWlzB
WltWxmtDRUVIKhO3f6iAezn3DTmuNZDm2zJCunMcynV1qSVw2L7Sl04PbaYjsacl
KwihDFT8/+MxhmAvFzFb8ymVgHIXeqIROutPiRGDHttNyxqORPgAxeyUGUvsMszl
ELkFrW3K2TbzPhl5EqgBrDtW9YlaHoCKpWnA2U+ur0FqDHKohdu+sM/FDeB0eHuF
L5HMVYdIRkL9jcRUKwTrdLVVNRgFPMRQd7N49ijqcDEIMTBeK6vCpUPSMeiF6H5w
PEV14Z2/IaR0A/xFtI58HsJ0rJcpNii9iN8NYiXz/F8bKV1aP1x+LNn2X+EUHJY1
nwb34fBwl8zHn5Hys60I3KgqudmoolaQoh3Fv+enA2HrIID9JLRmfpwQp5MSQsab
YlLnVGg2LkYZQQDurhcZdgK5D33E37UJ78+0OA3spLDnk7KEQHsLwdHQmyrECPmq
udoiNrH5cMMwqhFyLux7XXenZzL3LjXrSp1QOOElPwkpbYTDkvGtPvAH4gwL1GhL
x7Y0qwQJMm27VXaPtuc10ENx3HM+f4+WOxNEl0mCgEFGBCZ6cE+3Su9+h+10WM4B
qDJ/I4y6HztM/fAtoLeQ8gosCNJcMbr9AgzJwQCLUVBfsD+9Ss/8ynBgN8z5QJKN
n8Ei/YX70T4Lf5eFAz7yFRr1OBgyd7pkAmEoK0wKwPby7vQ0yIeJCZDoGkJAWvdS
NgDn2M801zHP5+htnhXmqvPk/DApM9j+s2QON1bmGLHBy6f6msJ+UozOKRfjrGr4
pBusZSrbbD1rTenWXLk4CA+npeuMkmGNbVoTcncvCJ/nD41E//vav0afRu9jCEQB
QWhN/XP073ZAw5j36PqpAi4ATTHCRoHuVbEN/HnHmz3i2zKlZrkRRgpw+j1YNcRT
kXsF8ONlUf8IQEmvmhjOLDkREPd9z5xzzXosmpP76BVnnXXlWcXdnLj6DK2AT1Rx
W9h00sG+T2N6iNUx/w00qBoZ4O8flUWWUEe/DIE2P97ozERjdei21ruhxKiy3pNP
RxS3t2BNz2H59m83gwPewDyYVLMJTzAkaE9v5/Ej8r9XA1mlwN8UGe2wC3OlKN1s
UJSEnr26ZCXHT6E5ITltRkHV8i/gLqKRMCukeTgTIOV2faQQKIoid1QVr6QnqgNm
JvAi3jF5iceWX/vMKv9vRakBBaGkhOZC2Cz31a8cFaXlW+k7+oqq8EmGPZNHtDI/
UgOi+W+1rsgZbLjge98AtGXVkrKf08ICFuBimOQZWL9iU9nyOMjNYdZY9nSv1c8p
R6/FOXuws/xGwXaVotbcj/9ibacAqrVBRpHjF5EsPBX4SHB+zhMrujl/1Q+LxKJa
D0VxEmzNROzzZZQYCPeV1JVo51uE3933e6d3bZBCr+EycnwWqIc+wflFej5+lAkm
KM1kg1ezhnUCx8ld8Rk3qLDfTpuCoG2fAixFY8LUAhyIZ4/uxMTv4LhFGFlXzu/F
YPqcw9oWOi9OvXvi+IwfcJDd9IVmd3Ev9BHWxNGvtEtKDGQppP4rrn6rxdmhFZsF
rO+Cc44xQIIC8sQc1tZPHAIDxeoWycSf1PzWNeD3+NHhEN0qOWckumBavJmmS6HD
qmOCaPMjB8XuyaPh1H4jIhRdCj+SCui7HowWemMLdIHPIvRxUqS6AhO/Z12L0jnM
pw2zwkstmOf5JwZixMJnBOH0lxxG8TtbFKoDyXnRgtTKy7e01S0dG5ruXpwMcKGG
AXXayXsWyjNKh34VssUkV/3eyiswFD5ql0c5/a1YWmTBy8gDvqAIFMFiPv5ynzNl
N4UQSYQxL/i0xmVpcZYLLbd/EZeF2+vWbY0piS09eSl/v6zFMn3zPqfw9fAJ4wyd
b/JcHde8KWwxNunCqPXAH8Yfd9k33ErGr2bHKJKygkkjrIkSHLigLSUjlH6HepWA
Tu3YpW0rp9KdfBJzAL0cvuSYCeQ6p1bwJT7vSPbh8RZQ6JuRVVwMKFc1EafV/Yho
ZJiBDDa4Thg5qDGIslyl+xG9Pe8hnJryYH+8wNWE8zOb06b3R+XRja8Igsx49E7c
EgK+lKul7E2sM1KVXVSb6ZE+nyjCtv3bupey5tqKj6Hfwp78xPGZOlHFnNRepUAB
qEheOlMlA8+vgJXjv+WhDyxkrK13iSz678QXFrlU1g9hB+dQcGlS8IOyueMsaClE
spRfxF9HnvLU3gpKCnst/nFvEw67pnqVCAkaso7Lm+ThAkmWzIB0MONx+qT/uC7a
Qit5pFnWRnQl/Grk3Q7BEw8lSELAByqS3j9kaqyL0ERIjw4cPA6BgjSZRtjysUCw
R5eMYzZCEU29ocCgSUz18VtiHxFBrztdd4xvZDFnjhKpmq2GOgadIWAesmkAJeeX
8WRKQoTgqvqxuBU3AuiQAgIYv2+2GiG9ae5Qc3PnQdLXvUzvKWLUGoiBDCpvV/8b
4F38Vx7G8UhLmpsa05FVU+OQB7IBlH7a5fWFcr/IVpIrnqamVpA7HCSqRWvg3/Yq
ULB8VMq6hVIQ5I9ReLfOmbaOdgkuYrPAPb6MFlh1KuOGwNrIfoB2mqA/YL1MNVi5
xx8lNpvMAgHtIZ77RKbytpHhz71jII8919u47W7dhS7Mtq7mVrJdJrveJolcOINM
1TU/KfK78Y6/dsclGI7kCc0cG10wOX/iPAfLkNLbO5ONEW7T5o9VkuMB+QySQ5Vt
6iGnPrwTG/CoQLU5nF9/29EpahZl2DMsOus5gY+wZzyNHNHD4VNHflg4WUTdaYar
KHxGaPImqSc25TqfE0xnjEOqLLJbBwOovlAfurIAgmq3OrhEMhnw3q5esBxDPUwy
IfleDzACoLQTvJLfEBcrwEBMTQaElUDx+00TknagQlDK8Oii9ZpeK4JoMySBElT+
nJ6a1/QayZE8U7fJf/MUIKa3PNhaEcvA+5A757fkUG+oIyGKPBEIaxiTWZDx1zZx
N7svKyKHUg0vz5eIHRjrz6FWA26BuH3OFl1E/3wEmnHFdWgw4zvi9H6vbUcKQwJd
ZWIC3hZInbDQzUc8faZ94BeyKCXax7N9bOPUPbzz3nmR492fEeOTPLYcITpSjjYN
2jb0fBJ3fKAlZkN89PlNjx3H4Ca7VRRGRg4Dov1Lo+XNiJqMrA6QUDL7lBafBWjk
H1RJbFIaKYyAFJHPtLyUhQMi6BMMVdEUUagxaSbAbyoyk4Qd3XHH9Zn278pK6ZWc
YLaXBGruCqaAA0shsu7MZ/ogqM60fdUDn2gTQvpSmi+r9GvX8rwRXnaDahgkYlKt
yHmk+T9oMhpTDv1wNIlUVxJFO91oeCuV6J0I1M/Losl9edfdLJTB1L2kBE5yZiDv
ZE5ZqetrFJy2zIL20q5mqWP5LRYVXZc5y4uzaC9RqmIN1ljfG2UuNPNxKgoKplpW
QIOruApazqeJhKDsmre02UF1domu7z0+bBPXgBaVUHTL0cq66aoT/pTNtRS/vnaS
aO8tEsKum+wcV4iWC0uVWlwDNmj9wulnGcifi4AGKqIE0tyhK5yzP1nDlPgLH+wx
NaxAn8QImnpYXHEm8ppS6PavGJXvQC2pB/pLa6ysbgdsIX4sMetCwpzGqp0fHehg
1SYecMLkvZXyYbWB+X8aoiYxeGYp7GXP/yEt82tiTtRF5fks69QSmIFiHr/YkcX5
0Jn02Ms04r2pkCeI5Li5al5IrbEMy0Mc+29OL7dVS8BC4ZGymGjpUKPqYdraw/rI
RbqQS7bVTs1Oz7VQ5skq7jslaDojokfmymbY0TI5KYu3jnmhVVyoHRKW3O171CxJ
QJi3pYKNzHX69falKT4J4QJsMswMOvr0YZ03KmHs9ksHWN51fZBReB2l/MF9rmzS
0fX6JV2jS/EXn8wvSx8jO3RfGOj03YtXTlfpHP//PbVCzeL325H9xHg78m/LOl3A
6AdIE2ykorZTucI9QYgPS2uuvmn278sEJ5bW4oRHHCkMdgvcQa3a+bi3hyofO6Wy
Vsf6bjKeWiJCm2AvCiAcKFC9DlpR9ZAElKaicBQMr6ZXFfV9W+kmEI2wxS5lRAAr
IqdRCTORk+A7/M6/aDNXmf6K6IBqfUJD94B3oy7JTIV/hVPrZQ444wZWqRAMCGho
rGEuxUSEjJuUJHnRKkq+PpAeIabtTmFxHUqlB/SLexlj7Ozgd/1YKj71JnihlVPl
274V/IzQGxOvSvZwfHsizuNhAUAfNZ+wj/sku6JCeqOatTdeJrWDXzvUtuPPRVOt
fMGs5ipK9Poy510pp/uuCctqFyfx1YLywU9D6XxbCKhWL4i2fOUBTshLcwID/u55
Lrg4fKTKe0xIEn7I+IQxYeJfzxoBi7syFmgACIbioGqDNShU+9gjkAzsjF9UL0k1
q04KivWoDBsbaNnHQHeycwe4rz1MjjFPks5f7P0FeVajxOGTaaDLmog/PNPkvIt1
pnXY032B+zARpFklKw3vmigeu8DEy3GQ2msdHcPtoh37jVpMGOyGTirqpHPUm9K5
6E8Fg0Mplg+HDXuNf8UOKOPN6jpSJnCfmSnV5/x/kOhENJgESnmw8gSQ6lUnHx3u
O8zsB0KifhYHB+G80V77rDDJplJB2ZYqB+TTDztTAsalp3tw/nNofGN6kGg92BPu
9cFm/G2cUZo91MlrwE9F3l5Bp3xhVsz53e4iKbcICUCgAZtQpHrlXQeSkfGw97Nc
VoEB2mPvDeEonQ5t9TTjpsJ0ALC/rgmO4slxbihzDLQrfI2V59m86AiUTS76gUM7
/hmGQNJ2X0cp6o8e2mwLCsZ4RJItG6TEpHazmC74vVbTiBDtPby3GucBMwd48tC0
s2m2TNb0tJ45YoKNky+X4pB8EJid8o4y9i4B0WgB2Llcw9FM5ZRwVrMqWXloVYke
XggdWy14tGmC8ufzH7WYCRoxXPnIRiN6ig0WZbB026HKy+XlH6m6z/cDiTDZl2QU
2XDtdrgfUZBr1rxciJlA1AIAB7udIe6M6kVcS5MLd5V6Eu8ydaqZFM9O4OBMnIMX
twZt5j6BMO5kBgSeK3RLMngzJ/JuoonsyxbY9pCs+dmu6izIRZp3U49fHORAXuXA
Y75Bo8XOqAfkLITiDkoe1PqzGYZtspHRjmvzvY7r/bdcM5lcWn97r0Yv7d+HzHKx
FHe9nwQ+XnNh9FK82DPwMhlC3yvi45zEgXgGyIwBS8Mwemx+3KCnhb+FlDypcA//
n+5JWJHE2dL7HMHe9xZX/Rn43l/Uzlh7CocSiCGqbowihqgTI9whPPsS7PErz+aq
lj/5Yk67QpHE5B0aav/Qe/Pzr6Gq/x14ZI4yTZDWvVZJZI27GQKsIz2y9WdmruUE
k4OPx4oA2t3+H3FkhOCTEYEPBFnuuEidL0ht7ggMeBwzWsprI3tZ+EwNfGe0ZHqo
wVUtl4RSFwhgImTwMhNvSFyJVOoNCjdJp30kbu19nQuhHfxSH/SmrkFWRp2Nwvx0
gSYbUn3MJUXm8tLCwX/LfCdndpR1gpURkeHJIu89NMvss0A3jd82o6Eld7iMj1Y5
1uktrzTA0UBkIpw/EUJ5iR45Q/2ixcG2lBSUY9/bnCZ4E+R/tSt2WsM/aXFPTFLS
nPLWp8xqNa6ZKnMaWcCO+6NrKv9iKveWunfOwMFMtg5wV7zjVDmQxSDtHjP2VOqM
7lwhbnPnKsvqzveXXjSXfVzT3rwrYqEDAWC2V/MQ2ajpDx9V4muCyH7S3AeF8dij
sg1wnp0/Hv1RQdvKHIExB+8UQm0MJay1CglzNbKLbjg7sccB6elRbotCzfqjA229
ARZjvbd87FUWVF8PP/6n9JruEn1FZ6WXvs563Z6ID0fymF2fFdGSEJA8upfSkovj
Y50nIhsT8BpdaT8bDs4cxRXypzEXR7DykAZxgFXTgx5L8E5U4Ir6Om1to+duDr5a
BrUGriOvDAONbsKqdsRBz6bwtB1dN8RKncDQnnszQqYVs95vJMWUY46y7B2H3iD4
Jq2MpelZTeSOLaDLDo9b+1ae/d9n0mfV2xKxYOAOfTFpTQXxWqjtbwshmveIzNpE
Gtdg4ICwWXuTM8xAG1bE1XD5IHVMwdBAo/HWr730Rq1g2OCaZJDYaf0dLG6iM6yp
zT1S4S2EjXGzvyM8iArrWJagMdVywbYQm+KnCxRz5mH3LGgQD6uBjNBAb3DHjNBx
Axqqv4/RtxgALQtzZc3r679quIESXzQ0JqWVU4zinXkdutfZ45o3c3WC1cRldjzw
LcEQ/0UcxwbAbnErYqN59VzczILuPBraFnydH8bAXckxaB5z+4vo4eM8DJzYPto+
sDwD9dl+y8xVJbn+Ter62fL5th0qN7Lc9iGAoz/FKvkPs4YB9JIUWO/Q2yo2yBgz
E/NBYU1WBjcvvp3t7mUHhau52B0TC+C4RzmUJJtf/hiWLxZWn7ezJXmeOM2OgyYJ
+ZrdwzgcfAFAHLiLFwiq1Gfgbxhn+oTflaKvxAWev74a13oU7YI/cU4SOoTf8uzw
Z68/eLIxonCbpB3JAuPyXYkU0ExCJuYeuuHlCfQ70KVVI62avkyedEnbD/4amrCB
RPxkUc4ZzgTIhfifQrisuabYPAWOzJyydBGQS1cI5Ocfmfif6sIjEG3KiMUzpvVh
sG7ZhMhhRDn8U5CKhwgFEU8prgAPg8RylWRMFjotc8MDf6WgNAdn398RoWBgyeU9
wr9HNSHn6vNyGHo8L/aoXpVo2yrM1+U9MnnyNqjmmh62YMgUtFlJo0by/xPp3gS9
WOaaisFHdSvDK74b0ada4SZ1ui7EY98eXTr9YgnWz31uOmliHptC6Wxz78df4Mmh
bmnMNjoffP0yZdRktkUZtegLQnMWpaceQfRZDwIHLS5967jrMmzNzZgclqN3UZi3
fkl1QUqNZrdmJJHcfjrdOhsKddEKy8s7YpX/ieYRwIwHkkOcKdE0y/mJCYxMPCzo
7jAl/rij3weKTSlK2tSBSDNgVwIqvYzotA6NtFqPHWJt97YDH1FfaCbRVUU+7MJP
sTXOCH7lsu062sQw5RtRrdcftdFiYDh4WgrTlxrrVlWW4Og+jQkzSaG667K02pJ8
8tB0hgpNNMfx+sYNFWsSmyfacvpxWY7ZGOox9l6Ue781CLweUNtsN2/2gTRXBOJO
CserYzP//wbw7aoC/PpwNsnFRns9HM/pygBM5R1YUHIbceBTSuUoeyi9NW6Ql5VL
nmpF/xqdFV8rKX5OiX8SoPnptwju/whA+OfusOKiCpRcM5/24hcPUjYijjnORQcE
rxurf3Tg7/uEok3HGXPYmBg8ugdLJ75/UPoECUz42MUPYMCpEXbX/RspUx1MwpPR
FJMsFCTQzCmeJ2fpVBHX19SYhwMUl2JMDlJK+k6fGxkkaGy4ote66lwdmfQTUHTU
KyKToRvNwiSc9yXbRQnurU+jz8czCFW15Hw0b5LjmNLUR1/4QnrPkd430N/cdkWw
mOP6MDnUUmSpdnkjyxvGG1qlwhog3RVGbCU3G0RovErDk6tQyJo+mvE8QOGrtCoQ
wO/Z46RWGIK3nNH56SQ3LUXgMILILthhVh08qP7pZ3pEZepODSh5jgfPjXUO73pW
1aSPMR8uQtyGcomkk2N6OdmzSGtCdn2oXbZgXEH9FrrZMIGlb0J4uBecztt+0HAg
Y5vUM4EYHc1F8urpZ+4IeO9562qzfK63DzrpkayMTelssaVztFJoiECWxcq3bnIM
mYGLCPiW2pQM85yL0qwDXIl9a5B84nNl+P3bKMagN/UYHUpASgTYiomkJDWM3KSX
JZSkK2XwgbbBxpqAcWmQE3VwbzstAtnVb14mDzQEbfk1bdIbTHixzkPvZg/S9NJD
jOgEusXCAyzf1GE6POU9cUQJXCJjagY+sVfr8tCjIGAz0f7UR8Br9ptxIikL4WR5
dSDH8ut9Qg/5qDpCq1UJJ7P1L/tKz+Z49kYZMrj+tZ8Xi4elwCkjtJlXe37wFpa3
bX8E/Dtzk5lO1Aewyph/wYFTTV0AXWzjMkHGhrvSLmslcAFwhdvkxsuwY7zSM141
1V2p8jjKspCbubc2QnvGhhJ2ZZvhVxBHmdXFypWsRxopVMzSLWOlfuBX9VYW3Km5
OL4twRTWq0KpjTvnHZbzVeC2+wZwoPV+QWtJTV/p06y4vDbgdxLBfs6kxgHwpdzw
OZwf0SFyFBEZvGEJl7VCYnWKExsSFPuX+tMkQJ5uU2buvIB58Y/QPFS2aZLN1TxR
QuBMtw3EVaBT8peoAJYGLUsqxBq+dl6M91hU4SDl+QtVb/w9hjFZpQoszKPPUoI+
63ak6cuMmOHuIaWceyGlFgqOrqXt8ReDWETx10Zvbk4dgpmph9FcWi5PjVMXHtbv
i1KwToj79dbiXzOUd8gr7HrTPBH6YDXZ4btz4BFUN3eRv1wJOpL6a6dY8ed1O9+S
miO1eY6VplLwuv2taWWXByhBXPtbtx4x6uuXDNAAVYHsThUjY7Vd8G94DSsHDC9T
QU9kK4uwODvit4+UBhKJSV9lRlKX/O/1RdxAkzsaHy6/C2M1pbSCEHq+0V4MsyEC
/F93I8MGSucT+jzSFqdQWjI+WBv75yHrHTLzQQWHwAwJ+/pRGO4rfJGmohYvXTQm
tRomVm1RI9jJsuW+jz/RjP6f2scoFa9TWC+d0Uz6U/jeq0lG4WvysNfiAH5PEmPn
22hcSM3j46oHZAJut71VVW9j+qD089KCLEVqjUhC1kYYRZHT2H8nIYDRJ09acwP6
yDnxel9Z0QmOQk78uzga7afqiTSuPMf2lYQkahEcvIaKQwtvlR1Qt0gnHjlBge2N
uTrJJ2dkJ4AMgWW/IcXL4iRQF8psaMxupZu7Y0otCzQFbp9Khn8O5ZSPsxhWYifV
vOI/kPueWIkHnVTyYtROOnp//YF3/MF2FWDEqQjBFH5SVkrkmFDH25yM+zoiLswJ
czOoS+3LOVbrnKB1DZreG2iUQjNKhLKSBNBq+UI5Y+OuHEW1ov4WnKvHEvfGHsf+
O1VDe4/yguEf9/Lpa9DY3Wgl11DzseaTcmIgc1PuX+AYdjXA43sZrq7vWcytnfHF
QJa/sm7u+DHNVtW+B423wVXbOo5mp/oGT0tLK+J4HkdWlTKjKz/p2NznVc7K48Gg
M6ZHbpo2jKPYUqtWnc+/5FWyZqVz50sZk19Mcli+fWl7kCLx32baNU9zK4G3dkOD
aXkeMV91nUH4pdwNn+E6jBma/YlfP57lt6cE8RJsNNPe2+iqm2DRkvNAQ2Q0Hq8y
ppg3dWiaD1bxi6WCNf352b7njKzlZo0l1GRSwqq5TRNouCCD7Wuy69faf1PhW07K
M/mSx+YplyShVkCkiJ+F/ClBRKl2KfyiMTbWCplrzkv7JUlGGFnOGxDzGBudPqhW
nvLqan5NLV0Ux4JujEY+H6PibX4IG1trde5OjPLDVJBG+18X0AvaRsQ1hYiObsXE
RlZ33GC3cf6kmAgpSmEEv2UWYA4z7woIUoJnPxYhcI+/3rVyq1YBvctrg+bPYDAM
AkEGE/Jen+UVg86uFwDOIvFl6dZIjDVgFAPo5dmrbmis3o26vdYXzG2eoVRCL7tG
mYP7oTOsiP6PANdWyg7kDhvKDxh8w4POL9wy386QeYDEKWCOKgsMuJj3hqfd+5kt
131JUr5PJpZkbXuNV4SUxd4kHzy1hzYuzhc0nJjf4ZQYbHj7PZmioEIiaOVl5pua
HwG7cJafo4B2AID5euKnWkVKbP90dqwjSWKDfXH/XQuTx2qLs0eG6s9D7J9cSxs9
8l5mhhLWTph/B8hAZfhwwvtZhTVMfsAte7y1otUjN4lJc8TV4D/hHz9ZTEfD3l61
fuo7+G0Mmq0kWqvw8ySQZvj3iVoiy+jDxNtYPWi6xuvam+/q8busUbwA8FtUaWAy
7TgdqaqvSBKOxTWFKECakhs56l5xLljdgqEacfNuiIvvQKWaX5i4tY8UiPj5aXs0
mfE4iLDvnDNIsYfmVxfBo43EFae2+EO7Pcyu2ugmTuNpK7Z/N/rne0yqjGAQlbGj
+aXhQ5FAqo4pl0myZdGAnN4U9WKv8NHprGA6eEOZZW8/mxHCOOCMpHoyQXbXs5YO
Elu/fbvieD2LBXPXJeBVAYFwDkKPGsI8cC3VNliP8WRN8LgmAkn/jMRMI3bEcdZg
iMddYS2M0//RfOjXj9Oicj14iYIZcYO0ArBcrvS3scJLco/cA+ezlT2KiStmcrUN
yZeBNM0E5bYDhUMWkUbQXZYuyBBCur911rNu1kkb23LXyanJddbhGcBXTIK5fR/N
Zqkd6TDWHespWy8G8Bt3xj/5o1nqzZgwC7dNTMUdpZZzchIiP3xxT+QnfOYe6a6h
uOeEA6K1z267hxttiowiSOej9QvqjyG6K96uIKEFrAIYiDfiLoQ6b01DrNPwLBJh
v/KJjjoYzy5dX36QlGAxHevguju76gTnv2T8UFecPBZOIfY3dl781qAh2Ais2UId
Vc8oV/2gclduigRAV0LjGVF6BFePAUYsJdJ/H+FDo2yJSyFZBepghwDQGp40y6KN
CSM3EvZauIaZJCd5DhuXBM8qKfHJvEX5MjabCt8XBuyTkDVWa28nQqcHbD7KEDuJ
jFTltC0mrpl6hUpZ5I7kq9rSCUV/QhtyZCphZH/dF6dSf9SlDF0GucNauMF5wAAg
Jyi9V0QvR5TfIpRQPwnMHjmslKFTRL+PCRR49x9l7WZ0vxbtIqrfThdk1iayPFKe
hNd/xsy+Gz6sWA2YuPM9ngiYgS0w9AJmOdCrzxd6o1nMTwuN44aROjwQXRdEpp+m
EUPk7NCJy23pTTyc4glFyz9XFyhzLLFrhn7nt8sSrdZh1XhrhA76jmxzUjRUpYNP
QdgFLin86oivrFTGJlDwG2yrGznZxfmXjWX2x/WgUEk+NRK84P2ZVtaDAnn16P+v
bGYlFGmK96dH6U9YjTUiQpI3KtnOH5nMFDcg8Gh47bnM/OCJ6gX6PrITUXocYzS8
0GH+uWpZK22l34Fy5HKp8OwheII4LgSdHyGvSOFPKRgZVqyrrCkylLDMGEfvo4xS
4ikdbhd/8Xt+SlPGqs8zjS/TrtBV7uHxSQud9uV2OCudZy758uNf2oydpfQgXC8S
A8pw/YyXyxj+AMZ5xGx/4qH2ZeWCwqqzQq2jAJpJS1wi1tbCM7oDwRQspI/amPCw
2QKyCZqUaGb0ibrEYEtcHqkBQ0KuEyKVgv/Zy3Nylv6YtglpR/JS3rDrLJheUWE1
dAsK9qQ++vq1BazcdENIteEy3ipw/M2orhIVQtVNMZGuRN7dyK7NrA08OL8vnKMM
DVGWw4yv+6rojhV+DRxV8xshp0ePb1ReCsMZXvmGzJUY/ysOM8HoZQTOCsXvaIYq
Uel7fTYY6QldWipotBdAXiVKVzpYXj7fpBZv54pftNEfE733c4ve7FeUxqyeoXxv
XagaP+1udgSK4bQG+JOp2F3oNcsfobP2vJEufSTm99M0WnlN2AHvch6gJqVeU75R
LC+j9QXEDRiRinibayz4rjSU3rqQLNLzpqIF2yYdG3c3pm/zwdYrz/+Iq4KD+TWY
r9KNiP6EI+IucKdEDzVoli0DnRguauzQtMiWnYbl1VCBy1M0IqFohI/05uqkOfdA
kT3g7qt4jy4kGnoja0LKb1JUeNa0Yar66MBwKRzc/D4plC9eR4rxrv+T3XsNNTc/
r8BivhBrhO1PXMu8jaf89qp1b1ESsY4T/AllTQCTXHqDxctbGLRoLIWEb8TaM38A
KnRgrrAYP2EMYEvWYqaAmYl7PmbvrncePeZHOxVg7nK3ht1La9Q/8lH0GfgxHXlO
KgBI1/dAcuAq5k3m+IaNkjE81IwQSnNCakXBMtXsGSr8UuT0LsGU1Swk3lnzDK2N
Vxl9whGhsc/CotB13BsnA/ipfg9q05lljRggXjY5VDVJj9qHVWfH2LZpjsWui9rN
i7d0cUg5aB2cXnvJdSI9uGLLo30XQoO/VU78W9mhQ4/slDJpNx19f9fVR72JtDqK
cNHgFzJ8T+8925pink37d5AALbDUwh4bqHt4Bc9XJaoLqZfYIb1UKf0dFjOiO5sr
7zgcDXFbCIw87h7JXYTJAoJlJTXo5j2xfpcS8qV3+3SaGLQaYfAjXvVtQdfAqZGv
NyEoVJp2aJ/Kbld0qXtY/4lR2k4f9uPOGQNMcUo0uj8rg/rN809SLctFf0PRBPZh
PHonknAAcC16R3p1OMiTtE3lYJpohir0VoAi3RJXZxjh/x+CX2dzzar4YbwPEh4o
nWI2s/v6wlzrsmdeRQOUt2zhWat/0WUFbIR50OGvnhYqVJRcAWaw8iEIgzHlcq8R
vKnGZYBFUXLZqamAR4XrdpBjcZzhGZM3DAxEpp0SG2r0XXKcECiS0SjSDmFesYXh
eE5Iwhjz0/fWikKidAwrTlmDGWC6SR4T3BRS3/r47Nj+fpH86getsonOcvPh8yB3
zB9u/9SlJARUsEe38MNxVQrZ8gbBTNfoXdTAmVP7wchMvQs8hlefJ3A16fKYX/cK
i9CmeTvfiWkJyfFaQAQfc3d+f/Jd60nkheuHpHGCjU6cEIjYA1nKWoTsba+I4LS6
RdOXza32UAoIrn9AJ9yoKHCIxSpyl6qHG/VzqLTlH4ekXE6LW0zXnaYXhcASo04R
ZhaegoWyMqw3Am/OBdbpeCkcTSOz4WrdqPICjNOBrHxGKA0qhg/3ko0cetauSwi5
g3WzWFKT95WWp81qQ8bI+ODmMyhLmE2V5pJeWzqFq4hKqXlEHcXM5wywlhy1+V0I
8OpTJB4XoZZLu6XIgevzQFzgJ5Gw9wnsIbeQKUnmHtq6D/hhwwf0uZqVKZSV0GIc
CPLMY3e33KWDYx+LSk2L8znzjj5kCASHgbG8NcwENv0q+M1+0OYRGj6teGeCT8Pl
Fxiy9UptGIuroPlvPlRdyCDNJOm2zKYFCJkL1KL3N0A+1SkWjRYcL8DRiEg8E5c2
P3Y8EPrvaC6q9L2n+b76kT+I1oSoB8tQ5LkaKFixe2c/uLXhWyesTl4wyieQeRjy
pOFEltkpRwIBBy9RgEPG0gnSrpxRr0QT6mjY+uqHn1nyxplz5wXBdwJK5nRBwNXV
QZIxUZzzxlz6P9T0v1lOIepxj4aAwhsj6NtIFp3kpZU6G7NRzXKWG2B2A1CzcEWI
BXMB81I4A+aFGQHmADFR4V5vmYGU0mNMbVE9ILLKctzH86uSWd0VGkZzr923Zz0n
0DTQUA3d69DijUUIFKgKxwSFtwdbMHby5PxQ8xJvy97rQykon0FQpQdz0xuIhHBK
tTDpQEBS6TfSMiieeOjaaJ8JRatb3X2oXDjHOas+8F1LZW1BJmHxV+h2tbhUP4Wj
B0GZLF4vrYUi6/ptGTa/rehGXRBxfydcXuj1aUbLddFu0eja4F+ymD5yqAIE9vWS
OjQbqM6a977J742stTf/05OoZuGpz0x95L+BBvUUe5qZ5r/qsn7Vokb4tika5fR9
Es+9fFcPqsxqUBciUDrnvhpCZGJI0KhIwjZTdbo/IcwCYKdp5r4puwpbXjM14UIA
f7W2j5PJA6ZuouHXo0FOpTMpX1oIGBCtwUqbcEp2ryUzVz7F60rpQveQSDcc1Wvd
I7rv4O3AwJ/mXaf7LJk7EuW6PRCsF5QxVrsUfuUc2oax9t+7qh85gXsCDQbc7bT7
REdQGgVun+/I3+wNJeGQ7Usn6/YgJg+2NT4yaqvPIZT5tvg5lsYB5IO98J9KaKqs
1day/kGn2Xxw8noApcrdGzeuAQ5lMt4K/YDz4pAOOfQWzdNHRpaOrycBN8mzE2kn
aQ9zzaICgMLDkxuHGUfzRdRIuWS1JgOst1QzRUrAHH0/4eaCiMXR6cKMtrLAPRC6
oplfmaYt+iVsXyLF1oa6O/7ctwgYCKFaRZ2v96ez0jKzZ84EmucjHBhQZADmuCOC
faGpzS4WcObkd/0qmk2BslD/EPiQlmbCgFEmXrs3D/5d6sRYG6SCcpE05/7DSfiv
1CXqhdzn7IZ6TuPulfhUzVdr+aw+Elya1mVtnubUq7MY2joWKdu7GSuZo6BxWbF5
HWDHuk0kgPE/QoYYstK7Zu7EgEnztUh4VzAFGufMKtYm1xDN9EAv/FDu90C2YO5g
Z7m2i97sBBBohP4VdZBwZId5jQcX47gx3uTlS7bbFphUC1su8NJEggKVu0C0yGr6
G+DYjApi5hwCuGmjDTgdEczr+/ZKMgFeoaAOGtVTLtOqrHd5uLURMons/x8ZZsHU
QnCQzYV+eruXq+8eGw7p1kl2sPl5j47NLxdFNtGV7CE+TZK470i8K6ATyCY8vZFX
vbVZ470OgX3LugbR0d7fvX74Gz5AKfl64p5XK4FmdIA2mPlSTQk4tmA41oeYJtVs
jJRCXH+HKa0rgJujcXJafma0AMwX4qkjMxJRO0/ou4sWJCOKXLzoW2Chmmq3jHxk
KfTxI5wktL3w5NA5oS2Q3ABvyaWiJmvusL5NOIuTZKUFBaLLHchwqelhlWHRiDJX
MvR9ZywlEzX8Klv95Ea3fMhRs1gq7ONu4jqq/GhctOa9/ToLMT5AMOIHNw+sBWos
prng4ye5x63x15L/ZHD8+pxmyeJ0Q+0dB6XZBsfUYW7ZL7zVyx7eK21x+svRP6KF
sShaYlWcaTWf2OfQT/ewJMRn3GacNpUxpCC7pJ7/63l8BD9XkAoCgG58JuBdal8c
Wqq0AUx/LKpa5/kCLN0JDSjinhm9fsS+i2LnqzVY1Xys4+VDkzxyafFn3MLwy1qC
m+0b5MWysUqC11txZb4knXhC0zTTii8eBde9+wcAKwZuMIZa2DebQDOpX+EY8gBv
SOYA7D2zq/P1zAg+FXo2Uk8A0d/f+vCFpvUx/Godm/nJbBrkro93NlTIqqHySitq
Oll2NkXHAOiGnCSn+8JDVxu4TmKUCDXJ099V4YAISepFJr3QlGniv+y1S8dDQi1B
O/hbnGissnqd7J9XZKIe3YTFl6VTel0pMvrOh5qLWs6xvnG2EVMnVbYoD4m2b9xr
uJXmPVYkvSURv3IFEd5nkV50wGHRUWL6O2Oe5PCbqdG1i7uQEkuQ1GWYCstCOWKP
WrJg0FGoCUfieOFKLvHSr/zmObC4lI8orjk+c96P7ItQ1UVucUKcurucBK23AuTL
wFY3z8CVJQHCA38aAKr9SFV7zSru/LKk3el/Id2TV6xpxxFgsBkxxLl1JgE1SWWY
FhmtMa6yf/5wXrK8VqfUPdEpr44r4DdJVPDQ6l7VGTZtYohSPYWLQTMgqeGGdFIj
xXtJTz4O0O2+vykXn4dxuGK+Mk9NLMBGoKTYVV85kR3n9DLpp7BO4nTxv0r+cLdJ
CG6k7yfIqMwpXcVXzjMN+Bj/fpYi42l9NQKfbYAcwuXh4DPCbPVUYgxiXkjhHke1
3gMoRslwyTAkWTtKS+9vASohm2iurb8Hlpav2OON91ZHJej0mTaicW/Z1KCdcFkf
5AKJWAaUSrQ1l4ib5xOgOVMgaFr18rKpDn8ON0cbGQs0vU5o9TR56BygsjVsOccd
sA1jGwEDh9JcTzmbGgA5CuqXT7bZ3IhAF8maQVJYdWxS85NhtCHReMQ+y/ATiZ5w
ET0eeSd0MCiYb0A7VtyHZyvM0hMCtv/TDfpzHqUO2kcr73/Bg+B/Q4u2xSyQfEAv
FQouVGR3rsqH0AwYHrILBhFPMaRVRh4RrfS9xiuZBAF7EXCGu2OjaTff5zXZcqK1
q8bNxf4W1+4av3zTzsk/nm6mPTjbhTql0ggU2TrMO7WNlCV63QaMr9R+88t74E4K
Va7rLLt9i0zR9jjOL01/00kaXicya+XlzqAM8oG23ezqjkOr4UOaZEd8tndHYWKh
5BNKExK6lAYPbpuzluLyOjbrjKUB5V33ABX8lghzvsFOtCcKxWVDPJIXwlCMYuOQ
71pgZvde50WYwtqRmJVYDuptd61Bi51cdu+UyX9o+c7Cq7gUh1/1F6uhnd518mdc
Q8E2Py7ZyRP5CbD7krrbRzHvIkxO/YVWDld+hc/OUYDN5jcsuacND4Tr0EcXYLBC
lfQzxLnB2MVrZZfBteAdykwpchce2Cub+UisUirbLWbDYm6mn8MRi78lAn9E4MDZ
VT4ideb6P8uX/L7MTVpeY8K9tv3XuOFMuYM+6EVbuPMC5aWwB3rKiQAMweuwCgoO
OmbEWxUrySe4zBGgxtqx7dwghuOHvxNbOw2a32328DRggQau5hhg309VbzI/g76o
cmpXLuIAkL+zLYKj2OB+ggGTcZ+zo8qaF5TI14uu+kGgXMaTUQYHniyRMfLCjyBI
A2hhQPl7gwVzElM7hFrEJ4DgDIzCKJMVBd7cHEDBvVNzHCK/MzW1KQZtuxjruKqA
dkW2GxfTSMkmdLBu1ow6Y0GUdMWYdVLMWUegPxyL/VvrLkgSR0miF/KiI/ma1YIK
lYcvqWUaYqJpE0mr6Y7XcJ1O8htzjX0JL46StnGZQEPmD9CjxuajINZ1vSavMnit
zVFfIF54WKAvZgumMXuVpzukao31hXBipDACdkRHiSKExxJ64rzuC3DwqCpV54qS
0hgIZIBiNo3zCwFbYTH7s5kPPGg4JnpYxxwgyGsKYzMT1M3MS056a3wGnZt5C/kW
rgDvrDiz6IBmMtXPLj642iTDYRsauLxiffLNCQTcng2RnXda531UgBLJwm4aPtQB
c+osnKj+Xec5StxUTKYSZBLVddodcPXZeTD7ZfNnGJXDo031rZGvZccXTeaajyzF
bLEk/dMWltEptHU1D7jbLteUu5xXp+yDN/IyPSrbCdUBFm9xGqGrMLX1ll4JMViA
Bn5b42VsVYWWgP2a5mehCYMNJyUBPvnVBAilxIxs3vNM82lIDNEI6gagfMxX1kxv
tEfLt87bJYYEQvRffEk30A8E3r37n6hJH6ARj5cjM7+h2+5t43hNrcUCTN0dt2Fj
mm+1n4wuuYKuSJKk8VQ72ua5ux5H8iQEKmEZg2fvfgQFxScMsG4/eYNg7LnZ3wvI
eNYB68EPvFmPPFbQJ+288iuvVLq5RZIW8Z20swRuBqHykoBh+Kj7qMzgE+zdzxmA
lhKpmfqYhwDEqoyx/XMx1PYS2yXlwRDZXNtgrlzqGXUJgVgjP7ftipQ4bFX6EqtL
ba1iWbKWBVUDruag/NfLqg1jhBkrz9Dn6PjeUmTKyrt3jKyIGFW1yuwVDIREzyCM
s3qI3ttheL1Qv1Cv7WMd3fYfe+Q6WBvcbQVmQ7ebKjKlj9ay05VXria7CRTTDHgX
Kr5H/QqKTnyZqUjPoVTrVv8A3Y51t6sc8zbkK15YjsGAO2ZyRQXqcUrz3Nyfn1jR
+Z8y36+23VcXiwYnA9+EnJjbHobG7DJVcTrMy28pI3V/PWpq1iGGA7LkiJ20U76Q
6bvbBxYvrupQdaXFL1U8xwvcEq8oA/R5Tz/186LO7hjEG7u3rs0Dly1gK8avfRKh
aU1JOdWB7hw5Mp3DK3TKTI0KWDvCz7pe7X6dG/Ibd3sheSfuyM/CMDU8voNbH2DA
kmP/Po/lDCLhkdyUxOm7Fhgz1nlnmOGRzujPKcXOa//cGFm0px3s8BAwnd7l1RbL
8CXLV417b/EVHTBI9UnVRlwChJu7w/MWds5kwvkjrhH6cunQhOrDcEWFo5wqfYzx
XmFvnHLsz4lo2/o5s9mTBJpu9a9nCXU9WKJj2eedOlfOcCXSCNkWsjgEzPzYH2yx
vEVQmNFYwSfBai1Lc1hadqKrWP+gLJvxMw5UHT8bNdc/UJmVdr0TBY+JSA3KAvc+
vjK56yT/Y/Yl+N11SnTvwDrDXTHwT7XMLLWfT65eBQQbYF0V9QEwJpeYAsS0cGrD
iGGADDXX19SSBqcBppHOC4VVKo/uc5lD0h90tYXH2oqsZcXiDFuLU4NzTfL/VBM6
yNAtFCXMmG7ukSqAo1iU0MDAbn8xKLHByVQ1HJSmIYAfjaoarH6LzZnXcpIYwgJJ
Nn2YIqQUJ2D80kIKP+GBnEVVF68zeQPS4fsusrF+XpPPvwDiGuhbC6FffR0NQ067
rAm39SLHhWQYWhz0lYtiOPTAeV6iUj/LA0vToAaGbJaqlglyNJeSUJkrrgfPzJLE
pyLkNyhHARqpnzFEScWwfPROOQqIJn6Gr/ox8UzpRrgb+hn45ET0ac7Xcb4JqfmD
qfWKfyR/4hqqnXC+qOxAymarLdryzOovumcwJHhMpcXaSB9OET/Gabe4Hc45TcUx
eW6TcyjCYKdycveLnZjLWActXSWNDmRmk1MjGgUcaH+hbjwvZGFeryLCUJSlUbQH
HF+bNDYJbAAuglHerq886W/zRRxAPVV1sUgSRd2Ip3/4Tv9yxUPGPp5WA5X33dw6
z+zwR7CGvnXt1n0Q0MLmjBQvs6fjnGZJ3BWRrT7+g/+ikwbF56L5T8kYxoRdd3mb
Lwrt53jPAJqzJY6VqTqbcFqcqXsH9ifqlSXTI0/tjcXq1jTK0DeJng3rr0JhGKPr
T7UhfOnzggdYKeamUBnti9xnOzAzsXDpP4nJRSHBA1aDourGIBT+73kPs1mUMhIC
syMCMvFNQ5wDf7M9tsJ+E2yXQynPfAuJMpuZ6jUcdABuYNmucyg9UrrfsAD0XlvS
8hwwuEY+VIPhYDU8dJWk0DIu/ZTKFWhQtwBKY8088G6BJpPR/1zQJLoAWfOxhgDr
bMYb8ewE89sWVKgGFTQimvxz0n+pDlxR4LjyKuGeso/a8a5ECbgF0tN+eIiGirSE
YbFm4N9IDgEloBSFgkp/GhnwuxX+GlyK2+Gg5M//lrCVMbMsPaykY4Ldvrw5+X3D
YbAXgMeIP063bJsAUz+DFmLXKQUcyq9sUTGFpgW/cQKM/FWh+ARyZDJdya5DtExj
i2Z48CrovlkTYQIk1k2qNA60HIHNYr/WOQHL1GOFZcRnPEp8hCSaSmxBHkc7XblN
hKAEbWHZ4N0Kzbz3e9rY/3XLP4QqCBEB5fQIytEg1JPUj7icuRKuhuvEPIWJssPU
nSeLeMZPT2WD/3AdW/dDiwwRj4XpDRhYx7h+Jh58c+MsFXnSis5nzhvI7WJTQUvv
nKC9AMAEt67fzr9yixRNM/Y9oLskc9VqgbALis4lTGfDulZVvHE5bABEijkw9G7k
Aq7rdjmIQteiLfYJU8H9V20GFgxBZONSsTL2Rwou/QnRedzFgrGqJZ01bxDP4vjf
QRKqx98eo14cra7NFtOfHOvg6mAZkYj5xEbXCctwzb1YN4y85CY/FtxA1JUcgKkQ
ORv344pFaYbRtGUve4yWwaaj1Gui+zDO9PVR+8D/cM9PcgTAoMV6gpflwPIgETHS
ROK8ejd0oWMwdBIr8dPR2EPu6uD8pm9V0TUAl0p0CLdlfV/3+Vh+qb0rsG7Q5FOd
ZUS1ar6fILX0L0TtzSXjGmm0/zmBtwUtYEKx6jUMMrPUfHk+o3J50NtpykJ48HEx
dZzFm69hRk9qUWuogPEMJOFN1vTjRj7vAUfpX3YO8Emlsa9v+j235OkiAGPTW/Wm
xAG+G4f4WyO+hqh4+65kn7k0nJZs0o2dVouH/dF9di+pF1ubG7HDqEyUBnd5jPMP
DQdoZJwKH5W73r61AzzMCQrCnYAIo5ci1IxZ4vrI8rUPNPjusECLhr8i76vda89c
ybNwKq35mC3CQzg6h9asGx5NM69jM4RVSvymk2G+GZOTzWXDqLHXGE7aoG7wqnuf
PwJL9EXZns0TM0yDc60Y5T0S96Ex4cwFRWVL9icVgkvbBLClOp6UL5lD2njL48Es
j9H5V57IFzC/75ad6tWP+QBMWA1YrzQVpP5ZC/t8aGS6ZL/nS6Njda6R2g4BYXst
hlTLlSigbWWhBJkivcEr5avmNj6XIZptmx71dbC00P8gHONF0XEMJj1WGrJTcA+G
wBk+dkW02TkJqll6yh4vx/PGEFestQVG+cXXJ5ewKRlrFFxjJ6vFqQh11izJTDN3
YPQtPYm0nVOeFuBmQWFp7GO7IG1cd+ec/1FUDN1VMjUfm/Sw1N4mUZhoK4i8VHrJ
tefOucJY/cmCS0GBp8rOprGz7n7qqpN/ML56y7znZylxejopXY2v+izTxod2NEJ1
wFThHCk+E+qbweGcrllRENBCmo1zVwOWNHdPAWTnHwP1G2tnh84bv92P2uooM3zA
F7C8og09+ar+LgYSSQoJnbenYWIic4aLKZIhKy598fFYQ4VTyA+KUzip1RK5m1ur
RuIOtugFbhguBeOfVTgj/0jxv2eP9u5FbtFWz+ay2yS6XCSfl6giLpNWSgSkpArq
IrJ7/jH5kQwSyOT3JTcKiqtBbhU4nQ9M3IA1kVLt5UO6yOIrh5h6QBXY0Y2Y39Cs
FfqO81CMeyF6ltN3uvaolGzzEDk5TAnnHKaoq1qzVPS8/OzMISm3E5adpZZnpFe+
2b6741M/gJjBNC9isxBNh5yjRMZOL0uDSJfjw7sEzJOKHNtrKAWTDtJI70tDtg5Y
oaCThbpzVmS+K2pqzI2zS23AW0cJxdoslNqwfeAf3rldNlxa2enEL/9DOXaAE/p2
LLo1LiY4hjKYfEzd/3nJZ3yMJ4ZYN8W9Z/Ay8e2gaE7vmc1lG5Gg2Ky92/SEYANi
vky4rJLrC1XFQ/rWgZcoKPC5IF8b9+m8v4iXDAe7XV3dwuPqqs5xBMJdsRQwQPyj
rg5RcD6OP+J062IEiWiypbZfatWcNYaANIHEVqD7bg6vzLZ7frYBH4Vk0OuYiXta
aJW89D+dCPnAU7aG3RRF64jNjrz/BkTsz0QxSUoMH+RSXcvCXWST3HJcRQHOVOaj
177YiWJFSRQyXAZvmftilcaifX1AP6Rs4Ggj9HfR74iAk46bKLO1GwLAjW+lBWD8
WpNBeEJ8SkkIvP2PtvwTsCyLykp4QnTEY/BJwlD9EakCBjYgHLT/2h5dTYpslJRQ
yGqPbqUJodmm++jU7Kt2b3h+NQiJwO2snrKUqiYSmQvDNE8kQnNRwm6G1d3WWF4d
0EJdcIZC1aHL2fEdX5RksRG20j42ZyQ4mE38I7hmIwiS07+gfShoEQrlhtJqTzoH
Des9C21oMBViU6+2AvCS6s2f642p3oFoLWMUA0KyMrL2wyn6YrD+BKS/TUOixpvv
KWk7bdoRAdXkpOjS0Q7fchCZhkaNTsV554jedjZTkXC3y42nNVbthcpUbM5MvEw/
5qZ6JWNhlswYL8NpeJo3ZzaiGdqi5d9XI1//klACxzfZhFltbdxCr9H9xZJ/h3lN
lZ+cjbn4BxMu6r+eQkeHKymhSeezv9AJoPEGeHnzOIpUc5TBrtYnhB9PjQd4e8Ca
ZJtJuAL2ftYe7BHgSyL7GPya0gqmwZhaUP1rLjRNNie6SgBn/AZrsBCQ+FQ8c0NQ
VI7DrkoT1N5wpAiEMLl1LAPC7F6dFIl6FNx1gDuj2pLCSMyArLFJz8+e9hdlOBQ5
CmSXBXIlJbTWTVoecVzXZBCoZfCmQYS4+PNB9FXwx0sfL5Z/eKBg5Yw5KrgGxIVa
xRLd7BAqhNtAZFUB3jv1KlDNvkEgxmi6TOfvlxC1De/e3aempxqWFp7kl+zDRKl3
4A4lzw78+ZGgnqIufElvVh3tZEtW2e3I+PMhJmdfJInfXgQoeBzyH0hCwb3o6Vff
fPUqLOThRV1YFAn1ST1Q9kTntGjwH+DiLXuAwupwV3+YKYyG/cUHBQNkUuJiONcQ
FKJWQ/iFJWoUIkKwbDuaw+rhAi0wuQOZYEhbeqf1eTr7VK2bU+Txdj9qa16zSLJn
CRFDWI313Wy+oimcnPomGhdyUF+mZsYpUzb++ChWIb+zdmj7jVS0ejhTwgX1EtIu
9faI0WhUMWM/wqO8CeLGw7pFR87sFbsibkPxjKuYAiEavLygnRFIJ/3Y94AiVS21
SAwL4hjDnrPUpdi5WRlr6ep3Av8i2dTD6HAPxNxrg1EaZ3RRLW3LMOXn5ZFPH8Yt
nPqAQmsfS6qkEluuycnBVAOI3XoiKjLKmpmSfouXNhMrcvq0qKF7Nb8ZhFAMHNgR
auvp0g4r/5Xv93huf3y4rk2dMrjWbrS8i1qHGUqTJZOJAmvl+h49NyeGG7fBZoN4
iEMPv2CVzys/YGiKKML5MCX6mklUDvA0ScVSzuJ2XutVgtjxe+xhBqra6isNUZLm
5ygdg1kexOnagCJwskc6rb/SupCZPIZuTmXvm3L1dkVWfwDCPUg/noqOH48v/Uqb
QQAKvSotcd2Pb1uRiCwffVzEVWGOgdKHzJxWyBb7+4cF37fk1RQcG6fsYiZqCZoM
4/8lRvhJIr2e0QPpNx5ATo1BTvKm9uRRo3ORez3H91M1JWHHt8MFaLHvieoz6whS
kU010YI68y/HmCJbYktERJkfWLH0mwPspW17SF54uyBnhZPsOmQ5ITdUCy2skd/x
ynro0uxx8lU/FYLyZFYyYQ0WK5UavXvYo2Yhrn71sUywCRYUvQ+iJaihWGIpHGZ7
QLF77KOOTizT40WQxWwVbcXtqwCI7hoSv5rg7IqKujmiPLyc63FHBtZeZZJMyqMO
H+IrPE218uxnJIGdaRWrlvzse7jfUmSDN7JnKFmBpTjXfOnW/tLGFz90T0ZZHNkn
JEy5BAWoMMtPmIsbpdt8bdBXHIq1Rn31nlRstIlodFKHrkYpSQQXPo1LZ7oP65gu
kr/ZwWrY0ND0seZdMTZ+PfGN3nuEAzODFSrWd66LbfHYgKZ6bNvrx4zaP5hMlFLi
AHQlAiWvHJPrhOA57REHcViEG5LToElukLcuKuiL16yTjIAzjTQZtItHL/W1cOrD
9rgTZ6q9QTmaYnhZQximzs5qiEU0ZyyDSkB7Ec/WFDQEyeUn1mdfH/cFkmE5Vh7I
J0QFS0pIrWrTN5Uk7NpbL0Un5VBgrMl0/Q01jdbBOGvZ7mzSFhXu3qY0kjGS6jaR
SN4ro3s+vkR5Zp6Vkylg6aKTlfVoK4NuqVwFlDJhTZJcRYmDX20jn0K+ZB+GIyVT
vsATRz9P/Aq8kOCNLlWCQe8rL5DgV7KVJI5KNaYd2wONj6fC91oXW9jx+Qncbak/
q4fVC5Zprv47juBbdD33ycSFU/e/QuGB0hDgUqORFife1wpHrNjl9XNNNiDfmA/v
YRRZuSf1mwRNC4Px6LBDEjhofczgdzuYUs+PFCdIEk39uJyPsnsnssk274ujQ094
pA6c0Sne2c/SuIOYcSCnCijnlUyJjmtcFZa1lH0LHcpoiFnG4zuC1vSf396ma1E/
kyaQLIntMktc9wK9pK9+8VtK0mxhPMCzuRSo8k3mclxQFm25CPF0f+jzr0nZsfpa
bMrnKyJ0iYzIWDtVoBKn0D5awfIq11nymuCKx6VdB8wUFtX/hwbe2JLK2rjIR5Rx
VQeBZqo9BUIbn+U1/Qep3uct8h9/1DSz5qJMZOuXjNEnG8GlJI5+IewzsIQqQRAT
mbwqQ2Mk+T2Nck/P/0gJw/aCC76lbtonerWLhdHONvXcgcdV2m0XlM2M9za3hi6q
61mvKQMoSAc2O4NEBIn+6fQmMM/pchfZ/V1kOIySqmm+E+6FwCO3tbQGFrdRPgff
1TTT0lX+J72Ti1K1htOXBaEgtzlQuw6Z7gRAxsxzlmZ/Vnthy7L+YCbKjBINWBdQ
OXqkh03hUQe7kRdIrw7FTd2gImZoOFwhD8jtUOWuUNUzT59yv4sUTRrUiKmdZT5v
95SM1s3eIHdBtEdm3TvfLfF1qWL9qsR+f0cIPD2l4iGpEHfRgH5xvy/bpPZIZq2i
hSQp2hLfcFVKCD6szayUo0dadiWOcGj1EsgYgfxYJySSKWblPyNEHCCGdy4EF81r
jxxO7/29vugiIcJucuGsoTEMrYdPpmFyMN2YquqS+fUv7a6B2GhP/hTK8JuRCce5
fQyUwMK3pZc1c/hmEnV0Zgyyo0SULcEAkhldh5jjJOhNSRtC30I06gxJL2vsF6zs
SFykRdRGJoZqo8B9tgFDYYmzr8h0RMwV5VmGheh1X0ItKDt/PppTqQHAh7c3NJVJ
QMjItscnCvEv+OM665rP6LAOlSakA6Gq6COkIRcEOLSirwavpWJmxLDPp8MgAD8F
eFNF301WZfQHTsBgFdD09xAZRehG2zZjG50wynkMAUaBNLXVTqNWneSQr4rVJub6
mPxnnBb96nTClNN7LCZkojJoQVw/87wTBA9vF0TWGqw4L3BJ5eyn9sMOOOzEbm+7
AAVc2Vp4lpSADsgVtAdteEzwbPyYNvYByZDjrUQv4hwwnaZGQ8O1jJcqo7oSKcQS
M3SE0r/qtev+xdhCgTbsLCeoyTpoA1jzbi4cyVIasWDHu20mAmMysWO4PAa9PLFu
hL2N52/BWzmksGvr3/6uuGDL5tjuFhQPL7WKGdabGIyPO/MUGFKOjhyCZhIFH0IO
MU4KTRXLOG3v1c+5XsXc0bVEAdOV+Jz4ddL7ptswTbaw5kvszUbHD9yPSlKKxsGz
cD2IrscU7wxJ1/8H9S8Twea7h0gUoYyZrsrgP2onaitSxR37JiHHfgeok6hJx7Lp
onkwICFuf6MD6LXhDfP6QS9IbDjOW0DFo1OUD7vQvDZ2Yj1YxICIdt6eTDrOSzXS
vqlvgipxINa+aL6XticIdJmJOhtPlSoemaUbk0gk3WZJng5fAWHdIap4OWzQ7hUN
JOYUrTLwRhpaDfaWOCQmE8euOnh9GT1asFxUYUes5TMI9sah9mxv4wOrxqH8fgtP
eqdZ/cDYbTUcxHxexgadcoUM3URd1ZVRSo5Jn8bg8Msd7O93n1DwUk/d+ZsrQZJ9
9eJnfGV82H+37SMaQtY5V94xiGbrjDLVR3Vsa8/p2jKdCp/31dI9dRAHt02wi33h
yyBWjLLblUxxg+sq/w7KvLdklXctASe0mST1xi+5Hs36qFCllaljMSHQY5MdGAHO
Wiw3ihm6I3cZ1tlyxIbp3d9AAlnLAmD3iDG03s3+85oCdo4DGavDJZp5W3PkaJZh
tIJL8ukujDn3glnqReMUcOfF9BUYhsyCllmds5UDzFgXJoOBe6ieVFz0MxbM0kDp
evMX2ZxJU7WMGo7dEozFfEQnB4PbtxLVYm5TrNccTe6mjgE6HoUg99/PpOkpSgli
620kPCtT6BFvvlAKjECegxubVvTe1/a/OQy540MLW49/Asu2d6gqfwuu6e1YCOfL
mMkppb3Iiwso84rJMUT8I+qa60nGTe5bLeq2IIIj6eswjc8lH61Gi7qBKOboumx0
whdXEz/tRGXa4NlJq+1Rts2uXCq04zRPpgJcMY2UmUrkXdeDxqFRAD7oRlt5NBHs
4KuFg4zovygGL5sfELPGZ/jy5a8sACsFLDiB8z4OoVSBzAM4ZbItjFIPbRUf4myn
crHQOpN5VjrfFM0SGUOhQjleAkEaNepiT3mwBT+FmDL3bW2dUBOQ4pxxTg10ZWSS
YwhhrMBcjQfJWt31ozSDsSu9FKzfZ27VXOuyS1z6s0utNnN6jFbEcErmjDGZEBjd
EedgZvxFBBuHEf9/Wplp4sQ3nw1nE5b3cng74URNupJh0pAyS0DM7T+HPYlG1sgA
Mbl14tfr1TIqIjaika3vz0kkJ+6XUXz+WorJGdyHGicLS3YiJItK++BjR2QYPnXj
6PIVnptBuv1RPPiFgeLeDkLladbEYRA1ts/h1rtVckVvvmlPIfjqvAa28hW6dFKY
jUJCqPqIWlauoF81wMcc9tlO0ufbvsWTmVkA7Rp+fg2pW3REFfP5u8oRyYMoia5Q
Sg8gWA7S8QiTfnoUHJxoy/pTHZE/7ir0OH/I6yK3W96tOCC1sPN5v8wvwH3NXkmk
28SxrDjO87OFxCb3D4YAX2plBWy0QL7Pes1BVMlmdSKmEKo5v8G4ztLk54vcb4rH
BATuDui4BD2na7/uaoW4waw26TfsmIX4zfmaRXdxpnQadfSkejRcdXIdyUxREwtI
ohHjAcAHcnoOVJm/GdzV6Ceb1EnGAv1o5yxfotaBiqDb/ujCgU6ft2hLvp9yqCiH
/xP/rnlwZuRIQJq45TWoc1WWk74RB1a2L87gkubWOBL9U7xevGPPX/uJLsHoDJnT
wlwwVRwAYRcX7bxXcYwB0hJQUM6Gtdpg4RoogQ8LoM9pcwd5cWMCqO9MG27Q0dks
cQpChE2xdaF3cYeQs1U7KRUtt+Y9eKO1AgSXd5kIspCf8nnF8qY8Q9ExtaFQbydC
XcY/hta/y6pqo/w/D33r6+zzF+auCXfz5u4ndVZ2pQ9H9C+IJBeUM5nDIXM3omrC
tDTCv6Cpum3MvDd5RhjIeaoIc7NAB59qf6jmcL9pvNxBiWDRgeHqpiTCrSS8zB/C
riLgESssT+uXHEXjPaHLa/KANV4BeWmh7lO1IZw5sq5ERCrTUUFoQcCbTMYcUzOb
I18Pc0mFTjX4j43aXe7hiT56J2KT5Tbz5QikGbHiiJAQ/tsFS9MTmmPQChSGd6Z8
1v0bvQZy5ANDtq/TLrBP92fp37IjQsB2R6H53wgWnEujDzOwucHmxT9kk3KMznKG
Rx5KHmjWE2q6gtooOZhEQZZg2NM+uIsgQk5urDejji2Zd32YtFs6kS6rHYsiDrz3
+SJQPRrNyCiqbAj+qDtCJJNJK73QNTKwAB05qc8RNxhXwjKm4rEsOyxq69nx49qY
aWlxsdNZHDh3sXpO+1cdXdshgLn8lIHXiyOcuq2UYS6CQSuBHapiVnS59Z1+XV2H
mtc35QHy12fVSKfno4A0sIafBtlL971rFC6EG3Mr3rGL76QUEZIWLzKoOMr4Xjv8
DPcFO0bzZgQTaYtgvtaoHhrxIpd4M2KNs59mf18IdhPKi6HfqQQk+9P01Nr8pcKV
MniZxZOi+g0/s9RD9EJi1GscBonAcKmEz+/50qyhpUdrftrCP8GfVzU4lIc9se0n
lmnAm7Q6GyVchNoUe0Tak6kh12lkXXFYHOljV7zfYosjxyEfu9Ri+2BjYtVBOqno
rAI9RL38M2QCl5bpOgi3tyjxxh5u6Tvsh0tB4WnUzgr9V7D1R8LFG0ff4sfXVncS
yeOKWL9msAROf2X1t3T0BZdanWB8ML1pLXqNCLuno09n6SVAksMQcbELqPuaOHP2
Cvf932IzLHhiMz6LB5IE95xD9QwPyZKMg5sZWPuhMFrTAS705FLqBbY9RE047q78
ZU24cpgrf886CkzzdTkUCqt7NTEB6qW3f5uPSvikWe9HgNeohb4JtnwwBXQR48WF
lKLjbKnTDtOAO/jWyg0n69AtBrAq90DSzBPG0eF6l21zOAgrPB13X1uP+lCFgFqw
EjNkX8qON+bj3mvDPeUq2WOR3oUB8ZkG27PNRDMWmKcb6O58KGR4I9Uxz3ZPJ+XU
TQgkY4aLw1qmUqerp6VlpAgY7bMUqK4HT8K132fXXCcFSnqKAehfy1yl5IM6ih/K
Gw1Xfzula8OVoOxRRgDCEi7soI9WBS/ND4RQ+iQO2opiWjYg9fA05aETAb4yMiXb
fSmnEzmtpxnIvUPgA+b4g0zViqBtB/YVm8266hYl1Vnlr1jptFQJ/qRf1zSQKKdr
dfByJDYg9B0Jt2+NEdE4nw//+RDV5haUMnegs1HoTTItn6LuAgr5mbciXApkdtbT
Xrvy/EXB218nax1By8EJGNkxXj4JvB3iWEiqz9QBk/sGWj0IrmwyMAN7AHyXPThO
q+zosdIWk1ztDX5K+MwZdZpiBPGwiGV97PiOrV79ulYJF9yZz0aNlbtDCLHxJ+nN
vOJug3VCsFnrBRPiNApwrvx5qHemzVFrA/7s93oR4sk3vFxqmn2qIusuu5egL2y0
Gfw0Kcm5WyGlhX3urXRo5k9nTKK2jGFTTgwClYlylTZFcT7IfwaIqrOAQW+YFgQP
PIOp1avKeTn0y5/y77XWT9+u5fg4CP/vYoCSFrLvJWwYLPj32KkbHdUdqxmfLDoc
eZ/TaeE81tL6/hM2RWzxC1UUabXkO38jntHXZIbL37t/fxdjZmDTZ1d3zP7HdQUG
5u04bD49F+evpyIAneeXpeKvZnOPoMCubZMlU3Zz58l7K2eI5pvCTj1iiX6bGfwA
1tzB+wHIf5riNf0hJ5jaquMFpv0CZHK3bupfIJyKKlsVI1xqbzYbOMzMLFltuqkx
XJ7U4V53FH2oBrJVila7+i+xwTd52UZCgcpCohFlVfNrJ1/qJyzOTuKQxweUp/PT
cx3Gc5a/4dsr7NZfZ5yuoHu8wfECGpSqRlsxZ3DOqCr+ibrBjYHjzdqoGl0rDjDt
y6Wo5lI9Kc3dLmwthVb0ZVU2uNm2KDTYWsjwq+nLMvrT2e/wwydx4KB43nytIATs
4xPtBLXiPTPfmPjqEROJvygkyO3JnnVaPfEddHK2VAZ9bvILdztFNgPjmCyGTDtw
FYzUJ8Iuy5rfmAs51hXWMEIw+lvmKVMfLwJYLdSZ6Yd8qWfgnrjOeJpECTo+Cte/
+5b4rPsf8vqSsqqpQcYL7KoxPBi075SC0HB9pER2b3DPDEUpZkSh8MaXsNx9erXY
l6GgDlj7nCtoAt+Q/rSZLO34K+P8LiOtowXm+mB7vZGALCpq4pUtpPDxSl4SG/EB
RhEAFJvBaxYCEk/4MzzIC5eMSH6DcvBweKcBdijHqFC95JUKHovAQdVE2o62fV9K
uM70mvIilMLE4A0QWWIrt6re2/rAk6Q/6ZFW8oW6eTNoO7f56FoO60UEfDNVuKUH
La1V80SNvSeSplk6DAKAzZFCyoZr2slsALeIWCLOuhuqCB0VwLPTFkOVPt9tdZgj
mr/OoAAMH3BLsjWPuVSDZMXoSwtuXBCG3KQNDgy+ozgNWc2pgZHPntL8D/nL5G6/
VmwVwmtY5A4cJUEdUm5Wv47J508TpRKD1SyLn3ws2i6iQMr3fRSyL/kcKV1kNCYA
oMoOcMBSBhBxRkchxKxSfOBGYp9i7VBCBUDu4YmyiQCSYarCZsSFsFzE0IPbc1dT
YeHLO+EMhISIeoD51J/oETbD2eicsr/sgLTMJlKABItcr8N7Xt3YfjdZBxSLs5Cq
KzeVrFGpGLQMY4LSanr62RnVIpx9ORzKLStVJsYi9xB73ShkAJlP8qX+5BpkKPRc
bsvW+NKGjMeof/evMQ8T4aVxCxhf23RPEAlRjsg0NsRxWOu+47juBuu5Acv+6oTh
5TPjw2prpxKA5fIUP7owvMI0PXkE01H8Df3y5ebBxlMuqqR76mnEdLSEa/e7c6Iz
F3CYYC+BeFoTK3RoJdey7G8q7d8U8TFWuiHuZ6ODJI4sPVnrlC8Ag0sJPRHYxCcG
i1HpRnzboa+jpjuC2D9aYWze7X5iZYwPoz6m8mxGiE15KwsSAm2M6hVoAw7VFxat
FZd0tsAOlBactEos5XYlee8I18SFwS1ZurhlYoXjnA1HHf9cFhaoQRC6+XvgKeSi
Afqi5OHCpljUp5T38yEM01S6QdC8wM/3ASuUh843MtlGdzvc2I3Z7lVixHYaXiyz
JoGrso5AwxXKsqXxdf9bUjvUjxgwr0poOO5+GZQmtlj4Y1TsmZjw69RZwqW2Yzss
gPpjoKvYJ9edSaYrIHVVFTJraK7ntICU1wO1DjNtzsSW1hnQkpairPd6skk5Scep
eLBsZsYg6AMKG6cu79F2npptiG85YIrfj1Qv+kJ1CT21cOwkqMITKd+Qb1+q5pwD
9RBwWxtfa+j4PlNBnWpVdE0QrS+C3Wm8ulnYfs9bVss1ObwV9+NIrnYutJo0d15n
R7e4YkwfircKBJllbJcTmTvdhgEMs/YdzlWCGOcSC6Wb0Pca3E9i1xr1rWJG8rmV
UqsdQd+gp34qZcS5KKN20aXwZKqUn+Bpx3aFsX4eQ5kZ//oxjNMgaQh4I31baJZf
P3WpVO6ryEyU7432RdDXwNBsYkOYAN6JxZ7UpK11KT8ugaybL/HOmCSZV5zmOPZJ
Mnxcige0CFsNTPR7U9YlK7FrVaEjs2TFSQPxxYw85hX1S3QgKx4/1DY9u/EtnU8W
5el+kVHum4C3ax9yoKZ4+hDr2b7rTCN4M800x1POveS9pqvAhpcrzfXUTRDggSJz
+T011GnS853iCsv2U2u/+0X5RXAkWaDtN+TdMnBgKfER2kFa8q/PUMrmWI26IxE5
kHwVKWHD9Jimr2rsYk5HP6B5zCq4au8vk1xBTbuY29ZeFunhzRdL7UbaugHjydLJ
VUemeczGr1fqDUS5tZizp4UDq2Sl/UDswlNp2KjRRje+IxKJaK3i8qacitKj73kn
yVlcWYrygaKZ1Fg05F7Wh6nDKcm3e2u6XHPdNQAavZWOXgdyL3pAzj0K7o4g5+yj
6BewS9sB7Hb2c+fx7gCxHsLDJz5na7HkohWQvPNdQS8a30+9B0fc3RuVAwiCakpH
NA+sVWOr6EDgSI4nH4lcWacnM5pK5JOaNWxc8DDFtCiYBTiRpCKkbRtXfQ72TB1A
Gk7+i7JtKAEyne1W4unXL89Aqki8ZN+KDDgpghf50TpcTUDse/IZkDj/9xv9Mcw4
m+wEBX2t58NCSf3UuwknJlkJXtszcYbvIHUHL02XFdnkFtaRD9I7T7PEr3SD1fEs
y8Hyegvospm1yxWfB0paekAFJAtKQgvVJ1Auhy3Cs0FFzcYBVbB/HxrqP3l2rLKI
Z4Jl8is7fYQHXMOH97V6czDL/yPUF/TR3+w8IZRGx1Rnry4jjBV0vBCuS+qwjqQj
J3kEs/OaZPjp/Dir1MAQ9hiaCmdIO+oqOuhzrYdAkpLwlvrlElAo6pw7Fk864lL+
we+aTBoExgGINqK1aKlEWNM+nHdhiXPmH0HIhWNtIdA30BPYM9/G2I/zdppf+pgA
2HfihUIfDJxTaLQhwCB+55wUXSCcz+Gi0lS3zXN/AB2RIHI656YznxK4PQOfgx6F
v1D3mvaucA+oHQDoGsWLMHoY+5y8HmeS1nX7vu/Rf4wT0EPKwmVk5WoDWzYc0/Lc
d37AatsmgfxrNKl1aLWMCpbSlz3FUG0PKnMvGGwsARy+YmVdRq8BQTLoHxtGCVQW
fzaQb8zYOrSjnW7Zx37tePY/LctXO1kQf4QslGOv5FhGpnMptxEKBmlPoG08zXPA
Y7MTMzi3RwDKHlqeVu4jorbe8gcLWdleRpaxO6AWRnrXhtiyO1Bhh4jZLqR43s2Q
v/y/8G1oKl0/pYGi53DylKKMOIgc4eWRoG8A/tOUx6T4jK2rki9oC5Mzcl5LTxlN
TuBZwNVwNagGriQmdQgf16h+Erib+SCSJfhbfUcdv3hC+4F9nx9j4/T1gWQAbWR/
3i65npTXVjXSBSLUzTFWfYwE/Qq4LtrhyZ28o22mnv02nD/Y0L2SlSuqWHbwm6YL
/xVNzqn1tx3TOzUVvZLPypEUrCNWn+kFpV/GXNfV2jJ8L4YhQopM6i2uzKjFYfg2
iA4D9g9G0xpKBiA4X1AErISaSRQ36RB9Nlc/lrHfq/IeyeiQgFWILH0yimR27776
MCWa1YfSFcE0HF8YIXKRLD3TQ+DnOjjjbM8suxySWfT3h+MoZBvXnRuDwgoP9UwB
5NXyUltNnwNtDNu/VaD3Mf+/g/X98g8kHS9aG2td8a40ODTNCliKHSCBOVeaCrE4
6EGJ5PLAJiovSO3gFDMhshcHTib3xGXqASeDkRx9GMOmSgrVgNk60cx8BpikTMbi
fBgqL5qz9FnulVBpblRU3cb5eQnrrBq8mdwshgE92w4ICoG3M4eVTWh5MchM+SJs
ZQlQfVQMvAEhsGz+WpOZ/4c+uoIYhSYdxoEdaQZL2GGqSstwsdecQt8BJv0YwD6c
AP7LtbqlhBvSpLezgE+eq9QIXTx+m/VwrUBFbblVOX4nJGvQ6Zkr8iEGGlb4ISaX
HprAHwRIqyTdTSnqpG51KYDBanpFLESUKEbP6ma/NNlOOu+K97kz8rLbgTVLf2iW
Lz7BOxQ9A7H9ncTykEoFMzkTYnNnHWEk8XN333uS51/DVLJfUeg64nNc8avJpHFP
2KCpxi8bjWHVO9j70Dw26FYKu15ma5j4KYxI6KO76c2OESyz3mU3POXVhY6rQWU4
E7BjwHrGelsAreR4VR1N2fpIlX4ZVP6G3bnJhTVOSQTDfiITwN8KzsIrEeJY5VZz
WiBtcaIg50aNjaIPb06FaiZNIgRjjo7HB3LFSORUyOGPUQzswmiTiJzF4yORHBwH
qKTxbW/fhPbJh1XL+unqXYVnt4MP+3axe9xC/rTs8Qn5ay3EVoB3p+cHAPzJ4+Vz
/SguJXyu5ndVkQvUEwCo/C33epwgRo0RwBQwdbrxPxScZ0hKdTDx3cs7dbwGg8a5
iddoZJjzQBKiE67do4/YcIQvqdU0W3yB8Z2SfuVVmMoIcibsLkW93ZYMyoVOTiWm
+yRHfUMJwbLDSwbqn07+YmbkOtO6lqms0OzL/q6cFgv0DMiMOQpRxTyyHRMEjlPn
OlnhKfWCPtZpsCBF/Af7qz4z5ax6E5ApFqNaJqsntBJcQdcXWZnoL6v2wTbiCUZp
QlTaCprlzVtd1+VuWyJNKEAF848dnZ4nTGEA28FfYqkAfjFyIp6e8+pKYDqNcdAi
Mxfp8dUG/PXmPEYKMUIsNsiF13JKbWPXqXYGqd6z1nUfNHRDIvchkMB/RSTKm6V+
ulJCspfE/edef4PPSlrA2mY8n4mC3c3mcOHdGqAAMlL5NcQxDYavQaRRDZb20uAo
RTom4Oa6UOaBxauHpyadEtlm+Gw5ozj+8K5AdBaH6QuTWDNN+ugdcxf4Ls9WICbK
SvjJS9yfnCvxK67REvk8sPdzzDDyakddOjV/sJGUuP5hXmsfDSvlnCjS3oBYX4CR
eZAXxuVlcMS0ETvac94gAWFAHV9JoyyPPN2YQ3NJpxd9GHrAmxH6UBLV/EmFI4A4
U5WB5r3Q4vOvKjxeUZfuTpXafyE5zEXYAGAqnbO11pHjoY4vnNuE0MtbWuFgsZp9
meQC5wUJS9OSgNEAR/VpeseRPde6P9Tn/EywNHoAD69g8ycxdd02XUMb1LSiyfTc
2UN/dQn8v8Pzs74qAzVbR+6YAuNwIDFqqsu/jdaHVovbcRukZdDj4reBsffRdAOD
0oEClWnK+SToPRE4RzLplnJLiVjp1KvDgdeMrY78OdlxGvGIWNqq5f97VyoLWA4h
TzH8XbtbO1fROSVLIsTiKvjvjf/GsghIOT7QnZCPCjVCoaWjuqyWKhjVkas9xXcG
iv8w0+GqQF9Kk4uXqoW59/LiUuvjdnSXx87klXlH7MuMSawnZQsKO0I/rvNwemFd
uenb3v9NXaaLB0/JL8+sDXtC/DPGM13mlpiDXnnJP9CzjFVg4rk2TKaC3NH66SxV
+309lW4PCrDmryXReTF+on09M9byPAxJVzBpqwrQtM38qPO16DY5hQSxHCWFuOcT
mxTtdju0ux3U9O4YE834tfl7WJi85Z4liYiMqqJA/9fZqtgOfgZOoZ/X9WDPWx5T
XfU/3FiJZrTGK1YMvVJnKA1EQD9oNUqTVRLcqFqsBZVf5pdprsjXr++GJQfK+mp2
e+pBRpvpDWjcq8fU+AsEkbQSyomOQX10fQ9WAWkOJD0iexQzoRsYKhGS4lOYem4n
6dkSbqA1etzmeVh1SJ+RxlUnRABgzZuyFDl/y/yhJTf76NL9wH+nqdEJKx8YWbwS
6tD5UJ+RdwRk+d1fup/nIt76PkhdY2AuWfbfDdNLp1Mqe7fBVvU9DQiRrwVroU79
Uf9dxinO2cE9hjhhUCRQuI5uohCWQ3zlCYOPSFO4CqZLeZ6IW0jZKb7isQdHD1I8
fNWVE3o0kZVHRTF/mhfViEtxhjdKw989LF2ye0xs+RZwdGW5r5eg0cd7Rl9XLHLj
yEp08KrOnO4rc0uFYBMfMdh/E7mlrIx5B23js9iFHDjJau+khlJYJ2mBSjqWGe/I
cbKaB7Im1Bh5M22x0AM5bNpZStY0EAwm6WEFXgEcX9zBl9eN6iighGlaqAXqR0HR
S7DMlBFyGze8TAozsuzzLjEEVA3leCfs1QaEFbB+HYCXiXxLD1dG3ANi8cvvZr7Q
YNPr1LsrHSQ2vIWtFa3zxzjhOzCQHp3Ty+7lOkDvPw2gKlcZv203DKIuwvJlzz7z
5f1PkTPw6qRTLLxujemGeED0GBIR1+UgCrVw+34BZeb3psStc3+h+mLnosqJgfdx
27ex83om4vPWReMNeXfY/3eyEE+bnmZ2SG3SxBANavtmPwjObFSdopub8D2eV/5N
oUCkERMsjc9exUDQYVZOCQX8o1Zaz+eDxSSR7gKqmPfvzhv5Yg8vNw18R3HRyzYo
9tErkehSw7GjJt8XzBjJIEa9L5h34CUUtJFzcIi8Vh7tfikPUxgw8GKzlccLkUqG
5ow+3Jdptyhtg3mwcLk8GmIzjrtnCGiXoOHXKZVqkbbAlBTCW+gdhMCH7q2RNoV1
zHgzH7+BlfIpVAZbrjl8VxsunrqquO7QclKpY5H2PxIL6uyXV+VL8bJydVKFVrHy
1Z2ecRTI8QcdAacu4YtIZURCs8ofpbgg22r5Uxz3K1e5aZHkWYDaby7w1TpT1IqC
xr8g3I1G+8ucVMCfGXCyDHuwHWn+g78CQ2nd4YWRE8GZMnhs2BwrAR8potuELTs8
22ucKZ3KjI8rFSY3H+iCikzjaDrPB16KWeqZM+6FSi/IsL09qy+/wCkcAweP6N76
/5e3pK5SIBSA8DeHXF1mFukZzk2RF4vIHvJvquprHRPf4nziORf/4sLS8p/KLo/I
PMjTLkRdmmA1eG82tVSXpmKLejakVKY1mnFcpS3+yEPTy4p0JhxKtlKXjuVngZI3
XQoBIctdW9ePEX+Rhp+Et8UViXcXOBqhSGVeJ2A0hXxI7Sw5+7cV9Vgnbiw5MqTk
N81ww7jxn/9JOC+ApJwZKdJUZ2WriBI0EQ0jSkm0Ulqh+gkDXcJf6UeHP2+fIU0u
GAOFEz6eFMHUNsr2SywUzpL8YjnEfRrYg1I43D1CABB7AayKk7gH2Aiehk6cv6wL
ytuQFHFLZcpA2gZQqe4YorixDkeqoZTRG1y0g6MXIWxllIk6Y784h5FR8rRQeNVD
77/4Oqr1MzNNs5wAW3ub29wHajvmMjxwy0W6Kozru5rvvR/XlISnWiLN8U2ndolI
K4hY2GZM4PF58j7PqBC1zEsNbywJIE6cpu1M3fMkmCrlB2nTsN1B5vbJwScsGQZ4
fc9Xq9Ro6/6eQXhyfyjvOgaixTrCqAwMDALiu/QKSZJrgb5eFuRXT7VmDI9hhONs
RCpFtSR3P93OyLy/v/NasW7b8DaJpdFMSPVzJv+Rt4w6v5eKvn7Y+5IEeXyl1vMG
0pTWzug4xb5AMt9VV+X7a2FUl4XiFNIB12VGHJ41YAx/Fh/3H1IyL9rrlQGyWjuI
AwPdhx8DLMuVJaKV+Zc128COR4mi7GWeHzLsfCCzCPkICuSX/iH4lXwot03RoITQ
Ck4fxID5sJS6AhwFhh7m/TklSV11MAzc7bpjnkE0t334xpqoO8IEM7dYxwXUK2Xl
DQTmow12107KJAG82AFtOZR01zvHDOa1q/mfJRQOgLvxSt3RmtFmtUuhtaFjuM8j
QgMNrbxC3U0MM3G4uZjtnKY2CLgEBhb+cORouLAQDTpFBmkUBEUCZuRGbe8vfbPV
vygcwIHexTuCE7krQzZtQjqfiwteLgHbb7lWN7tHeXstqK6hevhQdqggGvB1MWi5
hY1gUScWzV1ZxKVtYWqhsmy1X+ZqtKlScr3hnsLFSWGCGtigh3mL2gAvS2extiGC
gR4h/p1V7vGeC6cPJbErR6N1f3c1anEZ3zqqZ/V6SCD+9F61eDSo5gL1fz2kNF2T
7A/Ik371wKBoROAY7t2FVzzl8vQ5QILTg0pyG3A7BG1OJ3x83C5sCAXvBJ+s9r35
YeAY++1uwArKoU2AvA37enBSq31KFU5adZT2CjlrO/SzX/9xnXfmzzl5p5SskrCB
92UVZQyPMprDjvc6Kg+MsHuJ/K41FIpaclp4mL2yl6h+QaH45tvlDc4aK6Kdyf13
PJ/JjGo0GTi0w8+sdrAlN27oewZ9ug5KkaEMpZqKEG0F6MS+CHDQ4lDQQlgKYLYw
LNbSrhhdGm6brqEd6rHBIz6vRFJwK4BWxDEenmvYw+Uta5rD0Rq2eCAXemh36Vty
A3Act5InvgPTjnXlvomRyMBkxMu4YQRDCu6CDUlsrpz3fkCpQMg5NaMgJL+V/Tds
do/CPCEXk7vQDZiAVBN38a0eHEN8cdUEbPh3Dyix3xvUy8G6BrnwRgNiHbIlS1J6
hsOkzAvyxF6LLTspZ1yESlCCXQDeupxOOBipA9CtcCb017UeT1zlH3jIvifGIvid
CBRr6P8AWVUGqscHKv5kA+OfiR9LSl0ejbZE/GcZuFIpzIm1UazSf/g+H5fjFg8M
7kAeqJ6tj/BAyxy03u8Rix/bNYluD1GKVTkvIIdOf9FI9r4XCkmdjj1vmu0/61cp
7mewIXXjVrwneEKurXXu4au34ueFZqi/541ryB/gYoM4K/AQttx55TZBIE/QVo17
gDLlaKBtNLJWXB9E2SQCoU8r3XYwDm2vpJttAHFXZ+xqrn2FXGwf1mj4fGNSGaGo
tF/iiA8MUehbrAxyQkjGlpLDySDlBM3MTz8ok4JLfTsZwD9yUkHmkVZ+ro7l6gUC
ZTfRuR/DYg4FtK0svIrwLVtcnm+Ema4RVutD+hDm/S5FhFjsrCx9UVVATs4dAmFd
ZtfZ0RlxcENSwtuYHZQG0MJyTd7GaxWIUp2vaNd4i7YzPnPK0mzY5iuLTCbyvURV
kKhex+pu2IIbs3R/i7MoCtrIPtIv0eTmwJSnyyD7chP8l99J5cgK7DFjXoRhswX/
xPmILMtc3kUVxxN/1l2MZaPC3uO+52Zin74r9+ozoWio6XG592FVnbNy3M7OSLqk
BPp+CWdMMpOKWpSnl1pFJWh0IbW+lxXvfuM2TfBoNiBlSDa/zYs43w1aJIATF+jU
7UFac+sZGDSi6458r7urdCPZrORVh+os9RCTimciyUpOwAaphe6zFXaFHN78qItw
AzvwokS2F24kBvA1bygikTJ4P7r3neLs150Zc6EJmYtZez0MwDIwYM82y5B1wADE
a3sQgtNCkEvKEXZ38vGNkZh8ch6VKDUKlumIFwRwD1fG0SW/jTAsS9qNa3V8uIRl
rRUTKMb/AQgoVYBjs1bWaLCwGfBBnBYrqb7pAtt3OM2aB6A0ud7VIS7NDirze9F0
HR1iDvzdV++Dg4STVQn4/F7ofGPQWWamG9duJQ7QHG9bKo/k0U9/EzlqInnzVuji
FGwzu85NglaOf02f7+j/ecKIecM0iOqQu46wif9BuYSCdoJTaHxFRPYpAAugAsmN
T4BOLrOltW1bjXNe4DRg8/I+SERXnGW/HH7NYlJzFM8YRYeq0KwzLNXfj+BaHXot
57KfNwMxCEVfChdPEpl2Kbxipo/arsgx/gBPnF5hM4GCrru5bH6EQFeo8OG+INdo
8EfAPvqCzkU2ji3n/PMzi5srH8NhN9lQhmKFKXQ7FMvV6FcNMhwcArF3p9Xx1Dbh
+K8S+T9TM2nHebrqUqaxJNVH/7JR25GrynGfmtPeoPKDTZoHoWE2/YOM3e+dhFjj
BYQ2OVn4I5czXwrq4RB3+jV5w6Seepb96rt4QXMW/aatFz9pDLW7gMAIPKXUDp0U
4FHx8gbkbIlTp1KCgKkgw4MU2z5w/TGr85i44X7CzhXrbcfOWODQT127jENYCAD9
AdXli/ZCWmAtsAF8nOaOO+vtyScVqBH2L6bkYjpvZ3L/YJQiBU31aO8/xtNwIMIV
39tfKaqDfmDhFcYyeNt7Zn8Ud1voi/hkofS3yGGa54tb9glDMUXgMo1o/dxrX2mI
G+LEiNSlie8Ap0xurMuzf1ul6GzB2pLUdfvu7i4kZAOaQeHKwtOuGWGXNt9hv1Lx
LEPwQf3aQoYAyORTFu7YkPpasDocZgT7awdqqHLUIU9U03vhEp4UBMfIvgTbub8F
SFUEh4U00Fm3JJdFY3OY9ZuPZt0mjw7aKJBNxsy4ET+z7aLjclvx+ieZ7x9PWTwW
wzyHPx/FQKxR1yRpPt0Nf/5r7U4qMBop9lrw8RpRkBRTrE/4/akeQGdBo4T9Vvtk
RDgMaTErt13xGv8yIYrv1ys44IQYzGo6uM8Qkf2dGG6jFqIMYWfb7BZbpWxCY1oF
XhNwkGKRu5tK8Avcrh65NHrZXpVHIMrhZRlR3fbpwfsUPB2yXEMSjzBhM6NUYuAG
hOcUAWRqpfLhX5EMOYWM+4Lr5HeoWQ1OA0wC/0drsRXasJ4AvXtxLAtxxLYDqRpu
miK6rbmzHJFuixlqgEY6zdldd3sbDoz5kPdmvLgXXnRUUegurHgxuGvw+55IqG5c
lrZ5d6+lrxXmGNKX5ZGiUy6RP+gmNJi3n6oASOly3jD+Qx07/3CNkk1aBttgNN9R
BVZpv7j4NlMJOmoKfKMtNqnyyExj2JpSCfahTwn2goqoGYoDMBAutXAk/jbcnFDV
02fHMR+zl1KhWQNyczsskXnhP9DKzDvwSBdyunBtY2wmtfQcn7ibtzZPEzd75wAK
kTtCLEeNTjdJiT8OdrHYKyTCyOdDOb6Wj1R160oGXCYE20SuEr7haHNPvLR/+NGd
lQzStWaYKcTyzhjs/YnG5ed0rxmWh1hDKDvIId2OzRbzGFqiBYabkUwf9iT2Mdt4
+JM+NHCmNFbM337k8lW8MXMM/wSz1xJt4hITNSYDJa6zkQy5vuIleh8j8aW+NYUq
wzTU19ieNKGHFL9Gma0hBgi7pODFMCaLdOh1M79rAqOQwDcd7w+fBRXzugCMSPdz
jkuijmqApFFMZnC7kU8hktFq9H5ivRo6js05mEsTcf6NWniZojnFsLQkYHZ1ZApe
xh/RU5HmuIaiL5xVSk+WwnBz/+gWVeV8eWv5C1M8ekmp7z7q9KCJGz6ux9buAmpP
tUkJuNdnPlT20WMt1/U6RG3WBxgJuM337kcO2Su1ZghXsbgd/1OZk43Le0GGqhO3
54LxvLgoXvalLgzeOxSTW3fenh7GCWtLG86yPJCPxEi+W/AWEwwagNd5PSPMB5Sh
Yh/KDScIIX1BZR5JqrN8ybu1Y+PSa4YYgHvSBQkvDTiSUOKpZqgzxaCIyQl3vIow
nbbxy2Y21OhhLUCawfuEUG7sKiWTcxJubQ4b4dPZ3uo5DHkQi74IbEB3I4b4S9Pv
LLTGp4DIngKCWcGjlz/0L92iwv0WWHs4GTlP+XuDa7ENtllozHlozSNGJ3fljrCJ
cWy4DIVWPri60vtt67VnMErCAk9p+W3ZFTLzqf2bsIbE3AWDczz8oVjTqIem0FtF
Itdw3NMrXXa4EnAlELCUkbOyTsRNKj0ftSrs1CfGS6LDiZj9lFClczajis+29Mw6
DATy44LhWzdrsdt4ky0EoOz6M6qO7QnYrmFT5wVCtQLnLF4v4dBTgUrdncCps0Y/
VdmgTb0T2PW0EEfjDm6okpSqteuHs29oNgy6BOzrvR3PgOl/+X+Pyyirs0foLWO3
/auzHYttt32bYY9OQ6kJHCkYqPSIfWWXebkT0E/6pGmrIHQSch+9jjd92ftWatC4
20u9pXEqUvcLM3xYNlXSCGt68exhvjG/l+qpjFxTnLuF/7/SCgc5MeoXDsE6nxeN
7utc1T5MLk3dfrwBfPWTDqqPvQqxNgWPR8snKRudT4fqOql5rE/KwhEYK9XLXeme
V7q59zfRczHmoMLTL7S095HiPWv1OtdhucVr6QgJnB9fSTtDq1t3vVlVVgTqWu8B
QZwSY1hbLTjnX8ux22LHWyISL9cUfJtEr29nSk+CEZUtW3nTabOGm13bfJZxmnAq
zsro3cwGPADHblMTIKIgoQNZFu+1QEMFU62HxN9nRs6mIvYyIyFX4uDCAScAnH2D
K2cMX0jaWMhAJp/w13NKjO0KtpT3dRbGcnFAFEeS8KUAieG+NNpE2puggA9m5ZnJ
FId7jekLF0oZ6e2KFXuO25oFgTHihZs9XacxpAYTbs6WKyiwIA7X48LHCQ7YS58V
uL0xraapcSW5BOyO8e/fF67Hn90K5rXaicSIir0RtYZ0I870RlC+daotgSWHF6Ys
nBqbaDvBIRSOHENU0tvaCoLc3EsoQQ8DaBQDoP43zDjqlWBZq5nNQQ0NIbu9iMvl
yq9PWS/ox8/OTXTeQx0P2tvgydw/bKcRfCYUUhVtzfOLglnXiAAp8ptA7htmm4aW
CZ7FR7E5dyW2dns+NAtVoyKT++0W8mY7AjnsxMCR6u7vaN8EmndNgUJdWJviErFH
UZ/EAbSJpdXKPnJ20VTWRvVpkCMYG4w/p0WMjuxlsFDLuqBk3bngtLGV71sjg5Rw
UW32r/hhf3+JI603GFMRBEt4/ui7rsnnkZlnlGLwUw0/DKW+81z0cPuAxCkWTfXE
l5sBx1LKLu9qAwgjGHo3kPydD4NbR1AcqxpNU3dfEwoY6Jv9gWBxZuQVkGSA3j10
WiJiztDZEx5a+QnKF/xxsdM9nP7Yd0qOQH8ZLY/6b5xZUzOS6g/BShRElCOaM0aS
1p9h6pjQHeENmIJ5YzLG0h+2MbOpDS2KWuJzF9IFAJfCIq9iAG/JfaMdQVpL2vtX
8wO4Zb0ZNA0+ar2pbayYXM677wjGGrVE16r3N5AaPIpQbIW89lVM1a9QIv4ByraU
Kv9J+oerH6bTaKqlkGvcb/4dQCsskqIRRxRKY19tj7Iv0FvKcTqRHunQ1nJYIVVt
KN7fd5T9v5SEFRrrW884ZV5P0PicyBh1q9lzVt98Dy8HGX87tzbbgakhEZx+9PmS
0pSXZJ5mHG9u6t8rxVQ/gr1Th9+4v6y5IMOGRt/6+44vVKP6ngWSyXqN2nRYVKOL
5wfNlKpG/Zd3/gOQGFd0lW327anzFIQxTIcJ52iEG/ebsP/S+hTvRy8QvrlVegHY
Hxd/pIONNDdEtXkkzWLcnvcPPAwF7oY60YZkFw7hvhjzN1NrI2+FIZtaEcZjcrJm
N6FI+N4OOqNPu+TnDXoXLakt4XjPG/jXkLHNGEEs8OUL/hHBefLLa8iarxaHk9QC
R8PyWxaRUEc/nKJwuB0Ans885VXNUEeOIsZP4Anvoo8PjPaNnCl+hr67hLf85jeW
UH8uUzH9vYHM61FXLwo36oWRbkXs5a0DKnmtgLihMv9mgIEfss5bKGfPJTC4ullh
QN9sDof5D2ddSZU4xRAwvnf1HqPDI01x8SJj8scm1O+/ISio8L9dXanI1Yq6il/1
HqaZoazDzmKczvVBVy6UL+4Cl90x8WIUZ9hYOyqQf6VY5FAZE8OhdJk27RJiqQDO
DXWRlHD4BnwAk+uXjibYLuc6lRe0Lugub7CLqBGSzWGpHDgTXunKuBuPN4OD3Q/p
QplNqdwf83A6AytzOcdoZ9VAdEhmXVMGD6CFo9YLaact3OotPrjduOg/mGZCyuWk
KJ6mTkspNHBP28ugjFInU71DBLEZEE4Y1DDNDt7dKtu58dXrKSddnKNzDoBbA1wO
r+o5JUmzkb6dhKHci+C9A28DrgDjw1jyrWnRQ20RsmkB+klNaJz9uLOUghGHEShy
CPuzgtyUM3VNPyP1YPDxbeX5ueHutq7MbmqHlIFkJ/M2JB6k1P/43nBT6HLimWFa
EqvGHylUO1kfDvRUFKLi7TMXp6aAW8kTPYw+UyjWfAyAl8k1d33RrAoaQ65KBxj0
JFfJ6Om404YpEDtJVre98oaQvKLY+qedYV4K0bW+jrgjYGAPQv4v1+knMBZdhcJW
YUC9k7weK5eYyaQUxTozr0BZhUe/xX/DBNMC99DO5h8GfYLxmm1adkSp4zFCZYsu
I37MKbs7Qprf6+3vvkMySy13y+crEuO5MA3dFji4OUdsg6Xo812tcw2OoPEN5ycx
7navvoH4Mr6cX4mUJ/g0d4wMBDgGOXN6UEMViA7+ix4FOrTI+Jlu2JcK9M2KmdXP
4qUCFCbc6D9lf/wlVwys35aEbic2VsWz1Vf0GI0O8p6EwPEcyrmjELLeExgpLk2A
GronuwA4FTrbQ6zSYtPmts+U6ZFHugi4UfQvKVU9kMQreAilYDnyoUPlk26f5vpa
TtuX6FLG+rixHVR2M0YOTzQMFYmYk87S63TPnzbxZGyH++wiSEvxnyTO01u9wWgl
EpoWpwH8IzKa5Z02YSgao2+wXaqytTl1rtmEdG4RBZ7UUGIruNYaZDk0bgGugQoj
ezUveXd1sg9X9WQJEq8skedthe0WLt0dzI6lYWju6IoUWWmzVc125Icgx8DUjHxr
a473rnBoPrQ2MrvXO+Xibu4RFXofBFgd/rwuFIWIuiT4RL4K7ZTb5uO7xLtP8IDw
Hs4xIgWrLv2eC8IEXywjyZ1Xgtmy1ALGnDAOoI5ETPw5pHsXPLwJHT1UJA+sHSCm
DaWX91z8hAMHcHzrlFsYQ08dCHPKrvUtzOuYqoGVqwK8259eJpNmVaQzm0P2dA9F
47mhbJ3cXdTsdWB+x4Ck1uPEGKabLHSP103TVl1xg79v+UaCSQPuhaard6myf0na
fnWMEa25FnXk9GUGg9M+fBrOtOg2mWMlqSbadVcFC1RApVhwtAPB37H526NW11Wb
aqg3JOa068+OP29lHGSPh7xoeuSNWIjbWAuLOdGYOIekOPXXyBeWeIB3sEapA7r3
ZUrWMKqEQIFhdlXNsgg/ZOeNQiEdWP82ysg70sDW1tgrON44vGnfV6gSC2ayy//o
Rd7Zg+O8zK+yeousxr6KX94N1zN7lTMnmwSri1a0b1J/pCHiACPKnaDOKNC22MKY
/D5okXimKg026l55PfkQ40xUYFMm+xm5gBAtQnKL6xjKIt4yTcJ5TCpgpqOAnttq
90i5WAuTGsNMqNM0+APn1NHEZ1GNpBpzuoIK+gjIsAB6Q474m+1LpTO26w+3IlIF
qeb7pf8ySNgUSbUGk98bFxcXSviCKYbBuKaVpmmFOHtd4csB+VnwhyhWsKNHgnvj
LwRvQ2xfx48z6SKr5c6j54iMohRA1Y+c5yRRJeUnXrJWRiqWSuqKHctwPd1tDciS
edfb3flRlFY3i4SAyiZ/ZelBRjrcjNQYjXl9SFDPPswcoNtuWaqU1ZKtBXPS08t3
UN06y4Va/JXJPIXSEicEH3WtwUYyky+17779vvHvIxzrRs5rc6CRHH7z41ju2GJd
A4x6cj0VuQGMb4yI/Xd2yRhEfNFnTWcOGvbw/18Hznm7T5le83GhEKk07TIHnn8P
MJEZxJxiWoDCB7kRx8zJM4EZAbaIGJodrMFdsJ/0ggATiAAm3f0gueVcvKeiRFHn
Z0QgBi4mwIyicTsRj5m3qZ4BXn6AaJ5GBJIZziZKD5wKE+E+DDp70nzbkjvK8+P9
4FuU2zk3xWqIZNnD1s0VdgHyKeaF8YWZQx361K4cNgRZGxVtR7eOCWP9z01jR8ED
Kd80d8EIW1HeuavA9iz/WHbJfFryBp3Bq7Ebi1bwFWxuYhycais1k1iP6Yh9Tt6z
liVeXogjgYv8EBzBXblrubkiYBi7cuB5flMq/OzKbTkZwmrPaVT9cMHiwqYxsEWI
rquRO/7Y3Nm0Cc2DBZV4dNqnJ5L/jqEOc+WLWbSFZskGShFf7M9yZM96FUzu9neP
BimeNS8BpbfE7cHV7yDdBUnvTrAW+35xTEyfFRU3WtuhL7cT4BUBOl/anv2wgweH
Uo7BdiU6BXsIGEsSSjTLUJTIIE1Qz4lxFXy195dDYMtUS2gvxwXivr3aMpfplTpa
tsSID2pIUyJy7hx77elbldjs/DguXT+vd2W67ZOjPd/kosbh5b1RS0odfHzZWb2d
YnpBxSW/qrepPoMR0RW/3LsyRtDrn2MGyq2X7cAnCINn207DRCnzvLknk8z3Y/gF
qsVJQLti41lN+aUAbQRqGBhkC08YziNTjfg4nPTzgNZA1Hd6wOSY+aYRuEhsnOvX
wX0H2Sjg0sEeB13otBb7GC0/dAxkcbyhcOTDcJPtm6HOTiBYb+VKR+yuVMB4bGL5
BjkGm6a4KCLeiYyQHpkI2MEkaR9nTlgAJoxuz1NFOiT0ogmBQpnVkJvCl5alx4aX
jmyflYwoRM34CUSYw+uZB0LLSCQXakcUhtIUw9I05M0CnMShChYukytgtV4G7GZZ
L8flaK9JSIsrT3jx/DFhVOf9X/JyQ6Y0L9bwI80A1wiGv0hTZgLfSAbt+qPcI2XC
a2bkSklIY4JrgjFYqo5QuBFDegn2jxVsbkGcmJji1VSk/U5Ycj2m21VqAeV47VuI
0rXSWCaMNvJJEXE75jNn695Xm7rYgXvnlqVIrBk7dkpojJaZFUf8uwSHs7y4pK+v
jaICfGfRdAtDAsNvMiwt8YpzTMH3mXyQ1GzfhU+TcHhI7w9J0N/KP5A5MFYY0SvT
7Ys8JJQDwaPBHD74Yh4QedHMGVb+LdThTutm/LOpETBQqUYpzh5XQ6Z9pPphZMF4
235wA3mp/Z4LJP5OvcRHAkzbP79uffsWYe4Klm4T0S+c3UMUwImco+ZvLQQcWmb8
hs3wZImfyy0MTUVvC/J4LepTN8Esa3XsS964K1ryXR4T8HX6Drc1ghRIxT0j931q
lMQJDQJ8xpU45BE5wmrFIw6eRb4XQ+rJIWH4oxKtvUhRn9KuamJAVeCqcvEKvivt
I9dRkYIYIfkv5ShHrhOcYx6b+N8qb/msn34dj8ixfVHnsLqSZJeWElhTEnsq6J/g
XeQNS94m+og04dMMq2u602R7Y17AnQJD0wJ5MsBwBHAOes1lT7KvSJAbvCPpb1l8
RVQrBzJlEEDTFpgD0NN6HDhaiR1rEo2P5jhMdN6Eh7PhU+wIyH5fMnHzSbVJF4Tx
R6xplZHQVqUvH3pPoh3RhdxU500zo+b/R88Y94Jg+rX6d/t5HDourXR5ZhY9fLSE
nEsX5GmNPN3DD2e7bomgd3DE5dfJP/9gHQ6NbHOeN+Tx5U1hLtuoGHd91zI7mNXe
d/9vIzwFPDLcDe2kSvrKKP1rQafU6T9m7OsqGTAlbMS4DtQFu4oVoSz2FkVbsjKV
VFVR6a3icGnl5+unxDDdpuJPOIv8iM34ifVGFKASlzUVOFmsdbqA5GfzyWm1rH+6
nXxc4rDTe3h5WGLmpmKNWPOeV19XzxXrEzi4vv4/9TC9wWficxbKCucAlLDDdI0s
Tvde0FMQBEHh8kM3J63h0NqoTpf5Dnpb5DCgmg3MFA8FFmXOd1DXCQs+8IGdbGN3
vlKzeEZcyP7P1rSZxKeBdh5FvHuVtc//JkLR5zi7cuMK5/psXhdyoLQ1PGgI9x/x
3Qgi5N5NC3e8EtfF9AFyaI/NuMMwXZMpGYFbSecdtVXZg7W7mIx3XgwV3bW7fHs9
jP0jZNX11ySZBfQzGHzGpEB8tSQP7Kd45zUgn1TlTaK4tC4zj7T5+/DjgyH05A51
3FLi+AuhiXfTmpnV4c7mxnFwxRAqIeXXPCVKGs3p0htFp3J0Qy0fEJXGtEQEjWW3
F0KFD5yL/NcA+OSocY8j5OWfxWfzOM4G/SN9p5yZjjfk2cJdSAUV7p3sUkFhnn34
NW8HO54lqro2Fi3yT/nieHOcP+Rgb8AaFdH3RcO2CJSj6UD0YbdwVPB4wk1XB0Jh
R1gfv0y0m9lV3Qgm7Ucm0oXPYovRhnbjxbzQeFrz3Yn5g6Fje8mOKSfz+JIAY2uR
J8i9p/xoZhkjx01AR3D8Q+6zHrMsxVcTILG9cFbXmeYuakM3tXGK/d2GROMpQkig
DSpxZVMyCAZwF4qUFM2VlWh9seEfG6GXFbLXRAEoetrZQFxqUZEuta8BCEUOhvWA
PhI2xNSayscaYAxC4Di80vVl9K4izTtAEYJDiJk7++78v7ArY3kdM9SCwKEmmUai
A7q1GlgSZtIZB2dAKnDEZtD6gdb2nWSmwvL6MZHX378FcqdGtbvUoX2pfJeJWvwn
8ra3ADwpltPohK+cZfs9r15HMkHqjgVj5SCM5QLUdFdl9wOIbSf1pLe1MiScTKlK
vR9AAqIPWCNY3ZL8Lvx5Ic7bqlLOsWCIZCmaj9HHSwWWYszmeekoz3s5Eb9GuZcq
d6GO+fzmSpXH9XkaVxtCVDbzT/SgRYWu2tkCSsgn0KAQY7PkSb0OLWDpcagZxNX4
ubtfkkofM7U0nHDA1+r3uBJj8YoWKDQ97GmyWRi+6WJq2bv0KFik+pr9LrWRsK4E
L0pxsXiuVvQ1Wv+U86LWbhWMO6zAoV1DYEess6eMT0S0gIqv36q7PzkwDsoN6j7w
JlEDOFysJyPpiZI79QRf/id8sNLXf+/on9KZFX0vvrinf/BYbqKuvLjdvWI0Z/Rq
xC3s49Q0bHPIcEr8Fl4BLIp7cS05lYro9Lk0BLj0U+etAOkgPgT+INnUHhNdjjBE
+O44yZTkoE4vqaUZyFpb6VaLB4MEe1dJG52vpTS/aI8BmbvOK+qo8wPzduvJMRyB
NYkseu2ISlWWznD+7OofH8DvVve+d8bmp88zFeW8/7Be79GKUHvJPU9AWiPQBMkM
2SwWyQMPHzqHvqMI32v1XHnmTdIwRd/mRFMg1P/liH8TJ1AQD59p5dpo3UwZ/+1i
bIs8/z2HyG1No1nSxDEQh03fukwfvCDjmvrI9nYbfIT3HLkseUP3baSdsKG6tmNS
dlzclR4YMDXXY08Eho+drpfOlZiReSvjTD/ODP5saT5S6aD69kFmgTCyO2Xw8v5+
LkHLuktLR47lwoE6hdzcwN6LqeN9qgntNDc99VLzlEtRjb2NVRMOh4nTD1DbBsDK
QYR8poCs+i0ONNVD6CeDtdm/SftcG4yOC+/Bs1haRxbxjHuBV3W1ezD2GOQwG6hA
iz60uuNOBbZHusrXMXkgTwHTqnEnVHJQxom/hF7NPBNJHiBfh11ap6qJ9Zu5gjhh
vV5cZHnGU942DBCVzDHwoeyb83kbQg5X4XURfedE29ROV0CoFPz7Rmjpcj4x733y
NxWxloyAHUWHnlwc7LRoJE8X6AfbBeloqEoBYc8HQZaYkHNPx+QJ0cEcEbjgFBBl
WwLrrl79oXDR0Naiigy1Vz06+fcJyzfU0nQedE6hEjcg2Nb7KWqlwQlHWSBYHyGl
Yjcd1Xerp4aFs9ubMY0+/0/LFb/JY3ViUy1KRUc3/qzTtP8l3SODP4Q9i4hjbU4s
w+WnjTOhlEz476ggGrqPZ/Nl/G9PveuHO1O0ACHa2clTTRwI1+bPH4AYqn+0X8q3
E7T6vICO61vqXCDu3mciz7L1idM4FJ/JLwjdhGye+ppDqLj1UnzOcuiivIlcmlfP
vVSiMpoEkvfLEUXqMI+J1tb+ZymjvCTVxY7qSdWM/u3jC5AEJPBxNQeiZ6ImBmJH
6rotmKz8n/2fdKKQINWdLwGfaGP0VWdKDI2QAB6Uv06BEpYHGLz4V4UUZ54chmS4
4EAVDsn2n70i2CsWhGZb4YsMT82qB8UvLxd7qp42zDQDjq0J4Hzm7cXbHCNkpzIi
PH7iY75/02Nyb0RSmPunJ8O/ZVasx6rgES85btrFkyi3R2WWN3sE8S1cWgC2Kh2f
4ZbckGWKnDJisT5hSERPD9Vzlj/ycVmALhef3kDen/IwOAo0EgKUo027YrsdxbW0
3o1Plr5+4eFlseaBoqfSsnurOSeV/8C2pTL9zvsGJixFGYvr5JziPLC4kUAw6lbY
r1luIFjb/s44tG5KaOiOH54IdQdKg5/KJH6NyDA9KSMRCvHkIRMcJndu+vhtTXPY
j3g4Jp63BUV9UbWlTdM55Lu03anI+twomNbfb3oZyvTcZ9Jxt+XXS/lezTgDvhbJ
XwtkNKwzHHqq2GpdDBKkQ0vMIWlH3Hk8dlfeeLPEBLFqaGTKlT2N9Zg8A+1W6GBx
bbimmzxS8ganFka0zMBK51KOEg2DJO4u//t+lPHYMBiQ24jQp1kEt4t+Czg7o9zQ
MsuPDHYx7THGGrC6033UKp55srRHHbE52EP1V+3DvplLkzupFfSLb6C5NGhVQVZv
CcmUfqkgRWTQhOpGhCUpDXWfPZP4QeEs8s0/UFglTi6GMbWpGWUqXIiQBSj6zBnf
AAzQhRtJWElvfkwI1CIYPj4HJnnkCKJX5tCkDNdwdrrGXbV6YCF8ggPpD8CO6Xno
CDDNKVAXkF17dUNqEZVtXtz9N+755VG5cqrncX4fjzvfCtnqrJ7WPAjwHN6wSIj1
NsX0wpfHTrLi8OkEZzf6dzq9wgpW89sy1sG2CTilEfklVIDT++jNn78+cnbC3fHk
PxV/LZG7sNe2YC4dJYjA0bW5y55+eKx5Ud86xxisJDDmamRBxEIHceuOAbgDfFkw
oaGoh6shzH/W8laVDnLcPYDypuhE/1Ss4w80aouSO2Zgl8/EeEaWHj9GcoNhjp8a
X1g0F07eMtvEgIOC07ekfMkbrSdYc+Cr1Rx1tkolA8EYpMQ9SSt+K7UL/NaSxYmf
iijsf0otsrxY+++hYRzIGp05Gpis+KWG+49JSC8gGQCqTveZPTOQgkQDwCqZ6srF
R0mnic44ya2mnL2YRRrECYIC/I/aVepTvtI33g2/eAX6yQxbzthOgX334elo3iYH
K1EUMv9Ffxm3f0VGkwDf+Fp/RcnQcWbW9+uIa2Pvcm2Xa5Pm2hdKvdXf52OFN+cm
R9TIHhNA4GhdfBS2P1SOO16v9JbXuTF1XqjIHRkxwYmplRqYU1iUszPH0zV13GQz
rm8A0Qn1MN4RDb56kj3JV9orc8NKUnTPuYLzYh3gC+mFyat/ZvIbB11PjP/BGAA/
LglswP96j4zZqQtEtSS6ygXN58Rr5PLbK/hk6uF/t0OAQigk1+Mjd+zYDrIsIOAC
pfLtxDpIq+rYv0xO/TvazM8r5RA/EVUDWb9M8G+BFeIh38XjPj7zo+nut0cvI9Tx
Uc/E8BZlXCpREOIwbT7vcKJAnEmTAXpuHIQplL/HlHKhXegA2T30fwFxXtNyilbU
0UAtMIdAdKx9KwDqru5EpXMfTCacDlzWdvk2KXu957X8vNhBK8l8+uJA0njun1hE
hfDIezAv7LcHFoHxjzHZfVNuhUjgmq5D2vF2S/Okh9CGcK9HoT/sPnoOB9FZBblL
U8+ltO0uFa4zxpbTJC6lNA6x+PGvRd3aWNiZBBxvPBFc98gIoPbNaEB57wtXk2Pu
WXWHcmfCxeo7+oxPdb4MmXP72UDwvnZ/eafWil72301ItIbAOcSlDu/7O7Z68Y9h
QJ56XAxh3LYP4oJ2Q2GxawodCMXlH4ondJIzpcbFtVj0shpPebl25WIbXZqcqTVx
rTDuk9IE4nCBPtFwOOQ8Jo05C5zj+kZjcf7xDzYSy46+pLWq6IVeIebAM8GREmnO
wh2dgb0EPsv+lG4OtS2F7M7Jkt+aHnG7UKsUV0AcBZh09SlZNEenEZ7ZsXuIiYlL
cOpnzyQJFVuA0wAR0mxC2dJQjxQy/hgfz/U0y0rqNJiAozyF0PG6qHASZe6xvuYJ
+8Drg+o3yQBLcRIRcCIqAeufjyVTxslRVgfs0tBuIx1rS3uQXdUh2jrSbb8kSHeu
hXXTJdZ19Zg8MigL9UH7ulihUtw4KEayFeTuh5rKZDplTk9YZ1zEOhwEjZb8hZDO
XMX0gMkJr6CzsW+ybQjJYwolO0lw+oui6yTSj2avOvDKdZiuep0wlm97nRAqN6at
uoA76exwhOW0stxdLnE9+BxxrT7A7yISoyM/F3QT7jfwF0mg/A6/lkRwdntfL16z
CmVyrKBjWhuQmZ3WxJz8YMyAAlk/wWBwyp2sX0B4MCPti7K9rWQG2fZs770Y8vym
n0NigieuGZ7/0XGyOcCILjVvSPr+R02iMSdm1mRkfSU9meZV62Pwex+sxWr2QyJw
4jzRag5viFawUMacJXp+4o1tVIAnrPXU7nBm8Ih/8TdJ5NvjrR5yQQT9Q8VFD83u
/ipP+7cG+LJUKqh822fjBaf23wn2piYBDtU5N4qrVJ+bPzw5suHvg/FGLjeUqh58
rs6Hua3LpeqzDILgtGxPNN/vSRLjOsVZOJV+/2/xoOVnscv8Uhz4P6EwkMDE3RJ/
YIlTZePszO9uEMgqWbtilf2a0tWkEWfD7ecFGwv8bC0Lm7mpfJOIxHtf/nT9IHFN
JHkVKzs7Ru3zo273VV4CEI7UvfhEmWbljADoYHsQzJRneo4oh/W0fdx4e+NWC+Sm
7FCagGpC5XorWgStp01oNDZHE0cKvmbcf5oJL4146dI3G7/LBXDsTO/q6sH2IDma
PaSbW/uV+IZWs9rADFuAR9JT+zpa6LZvVQneN+DkQuY5/fwvR0cOtKejqYr5t44A
qCdOLc5Xzyp6oSZudkYjmhGtDiWnUsSFQtBrZBCi1KmQ8op+1gYBu3bi2zSbu+QJ
B9r27xuMcdc71cBDKUr/DgVpQSHyIKCV61ZkJtq0SpVrvYlTg1/hefvGr7xHW7HS
I8w0Z9rOFtCX9JrBheDFH6cd7knihhecu7Pd1vNP3TFJkkFvLE/o5oXesLGq7+dF
4eoKSNmOOST/oIj/E00gRzoHC2Rfflx0qhI0iwe3bbo2ZS5ARl5ft9qa5Kw0cNLk
PJOg13qNG/IGDgAT5yra7zRCet9WGtbK+g3FLUdRSZgTOtupcYghgDakb67aHhd0
F6bxIqKkwsiHtsqpLaR43KrDCH3zueUZHGmS/5Wxpn2PADa/FtJKLt+jYh0dtoRH
DTmCzws2zcYABMsB6Qbgb2/VYNPbJ0F7ONn31nFUNosg8pVLD6df+BHaTgJqoO30
4WeUGCr+IfW3rt/54n0nCXxiVDHyoXEraHlj0HHr5L6lvZoiZKMecV6wCrbKSyGZ
b/O90TDuhntgvdEZADG/vnhTSfLs3CqsqkBJG3MTnT0imAcAcO28PUFezRvPoiyL
Qn1KHhFLg2V0az6M7CC9MGpX2IQWCecMV5Bv0/f9RGY/e9QK3hBCav019H0Sj5ty
J2v7Z4IFMoaMWmcr2Xm3h0+rLf1mmSCu8GvWMHl6pqIk1FbeuwVgABuMtGcT9GTA
Q7Jn3ulVvpDUA0v8vDnFObIc/WqKY9nhqNp/QrqbeXV/k02U4KE/4SaKNUhwa5UX
ZoKXbMZvc6wZ6tXgZ46d91GWAQm83vBqC4GlpVmE2bGWa4exPIapAnT+cVudQLA0
8QmGFIoMag/QMFBY2u91/KjzsN26hWXSjHEmufH1ipQq5zawh2Miz3K2JoC+IBgp
ymRDnBiMxZpg5+vSMUmLqxQs3VM7NThEiygcIgZk2ZiKTc7vNQSUzPMf2Bx0t1tF
tuzLwUHJToffLPh3OycCj8uFT/1PSMVs47EpDR2r/u3bMxccDyG4jM5npfDyyQIO
tm7QqQ/kWvmz4BDA7Y2bRTq/L5np7+FKSHdWbBq7BTosZXuggdMigGJzWeh81+6l
QgSMgTGVu/iImCLHwYcfpM0wVcHs3QVybJ/w9u13LPIOKVRFckKPLNnp+kFfZN4H
+JmI1N6s4eV+f13sPk02xa/0pt3EBIa6FusyEjUSkqrdsI9ecDoF8a7Jj7wMqBGa
Ftc5kUcTfCs/dKXPFzrAUzznofJ9mSxxDBqIRY2Nh99Yd7uK6+GsvfP7CiAhl1i+
heKOghiuwl/DS5YNxfLWc/DLkj4rp/66PlLCwEoQViFSXQijTmXV7Ay8Ij25DwFf
7nt8oFudjcfUSV6bNWFIkm6BIIG8wJsnyJlJWb87bDRqXngy2BF6AGU6fPgwABD8
gDK3LsGKn6p26hZpKAV+GO5VoBnrJ3RjfxlbOMFCLjMy+EUTK8Q12GD8vtCgCT9u
/GPQN2NVMw4Ipmh7XKSAHLyGFtBzxCsolUvsknhwj2AM0yw5a79Yv+3gPHEr8DiL
X2QMyQfWp86ye/I6ErP2RIqgL+o1MXmUY2oB/zte98IoknFYoYdMcLBQA2GvWaT7
z6JQMgcdN/86zrTp1Kbjeq1ISf8zEnZ4QPpHv9+zjuayWiqszKhDLgX6ZCKHRBjr
8/bYmOPBaWr9DWg15fYlAeYiURftsCoXyjVjVVux3iwPfjH9WafA+KGIiRBYtMnR
Mnyqq/9gVUrWbIcUMdKmhDZbNyoGQ+KvzAvVTPhgNYn6OZxoxkLqc4+TDU41SkrW
GfT8qSp8QI3l0oJiYoA1iZRFOU/gICF77J6cRxAD6NS/hRUW2J5T/cGd3bHXKlka
huIK9OfUmVCQ7F3xSFYxnYn6BMJmLOUeSnUeTrDg1DhVf08z5WRL5KeZFyc4KGXp
M/eOwEVlqx6mZQXUg/vIHSWvLGthhGqXi3dBS6NFslVkK20yBNtY1dRIfOeU/H1H
2RKXoS/49vXT7ticllyyQ9Dfph6stdKsVtvaFIM1u3UqPYu3Vq4rIrczLJiyjyAv
ya0WM305MQe928379pJYwUGfihsXRN4xL5elTe+EmpQBK+Zb/nth8OGN6t3H0RFL
5v1xQZwiZYtK8bV/OYZm7KSq8Xv4ypkHMjP5S3rg6WnNQvJtJiOLlK3KC8rEDoX1
CYb94KnmTcjSiEApdduzx6n0SWmjLGXtow4CNBbX0k223CyJeWGz65vZ80QvF8LL
vhaVezQtnR53Vt8o0Etw552Q5CFT0CXVSOd+pSqEGmjddBpQBTfEdNek4VBqnARr
xZLjN2DG25f1L7kCbs208Q0wtghsHuToLVtyCcnK6YXF40TouzONoFNwIVW9P++6
yk4Ttef5o0O4bKeZVSU9W3Hca+7hsmPTAhnyc/0R9PYCbmosLkeDfwAPi2rql9tv
1i5cVu4o6/JdD9S4P3OkCNwR32aLCMgn2QsPRXT3T/jY8gm/lavxoAp3BrnuB0Y3
Vfwy9x8waKWgBW96fHoWTRZ/V14KlyGIPR8x2ljreOvUm7t3Tn6EFMAvEuGYnMKK
UzEQCuh81oxzjYk2aJ8fFABx0c1gOsamHrJ3qncX+Vxro2ggQtjkBt0Q5ZDdQJL/
OCI8j/W6yqca9BNoeyH/nmg7WF3X2YvzxkAxK6n9RRKcfaRQHsM4MSIjtGarJZ2a
tErySkm7+0XTX9eGvVOjyHGZLMOpfLZyfq2+Vm/2b1zS2i/vJCasVvB7ssby8dFS
NkyEbO8clkfHKIBaWZnhXpoluhWY8PrKfoW89noyLbDxU+dUqJTzRWQaEHHyTplP
/Q5laxXy8dmPGPm402hxfUv/wnE1C/bP3pDVkLoN5aoMrC+9AtC5ugtUUCUJQCfp
r7+K7bkq5+rVXj1RtbaXxdKEmesFOt8sXkwjksV4KhQWLGmeP+m+KW22Xcp72yfX
KeEK8KE1C4gto/zqNxHJYufP/yY5rf977X/YM5F2mXiWgQinTNDY/BsIf39z3VGo
cMaKrQn2UM4v8Hh/3nF0z2gUy+7BVVOt3XLBJUe5CFIozoE7sEj6IX1VRPADrAfp
qYiRVVzzqZ82WVeKjU4TsKdabjDrneUVc0/MMu8EBnAhEfwZBbK0HsHtsD3GlspJ
PG57Fac30Z/TXcBydNbMPlSLVFIRqvsC39Qu2UDBW+NBqhoQ7hl5kYRvXJE8dpff
F60tkdLO62ikSlim+GBajKBcAYcPKJu1Ixm4yJlSYUuMOOUhBorrwSn3fr5VEA6y
g5WvAjGJj0m4iK8YnzAqZlM8RuiFyMOZ+PjkfhYsJI+55DqRBpO+jpU9zrCLLY1t
scrKYOtXej92bN5j7qGIZSP5DQu+k/DojfVY421hWNYKSyndOpcexRx/cqrRvj7B
tEriZ4pbdtWc+7DQlhH/do5+4TM2TQgmA71OdsRIDvzbPX+IXw3SMgEaD71pKCE+
InPtLqKi4s0J0icuEfg8oOcO71+xNck155I6lXSGnfxUoiJY9v6VTj4Br/sAP8SL
Gi4yXlCykqUOXj+/ovFQvcQODS77tLzXDn/zqz1EEwlCy3LqI0gwJD0+wZvAKO/8
zBIhwn0U0do7E54r1acovsy9XHdAPJw8yLpA1LO+hq21Jg02l3ECLaHKfW/X/QnX
oh5b9jSpjPRCn9aCiaAfPy7SF4kZLOUQOpgPRjobdBOLvT/IhF/TcdFfc5j4lU6U
EaYoJYtSfuHFnLvGDJM0/iwnQGj5LkrsgBOa8i415GmoGOOo1vAiiaveGup3Zd4l
rCg4DrAhClBDOBJ2bP+FBGafPBS9Lg2tfc2hiPUY9wYKKZd0UbmXE0v+sg4+DAey
FwCgSm1GPoDF1YRgmOM1ioyDyo73QDKbDlHwD96OLy4erXj9+sUAT8Hz+0ZOwKjN
2cUkUmoZmZhE7Dzdd2yu6nUFQnQqa38pBCBSHr/fBPjdncfSl53ayetz4ljYPo/+
4h8XXjZ+eO9mvvU/4+KpOH9DgcTE/vlBcpBbHkp+D4b4omdEb3fKk4fO9uQtCXPF
tn0sszlH5i0gcs9GEFWhat63dRcqfYv55qwF0YXM44aZ4Eabn6J/o00Lw8h/HKHU
ctCrwdNwJixV3xlVkCyBECI8mVnMeHM6hr5XfBYJimRPnWSZd6Jb1qAl/aLOY4WS
3EswE0zTEg7Zdk+GdH2NBBosoAJt39XY/P+ZLf7lPVn5bI04LQbxpsGzAdPv4xqO
Jb8vApHBaaxqEOHQppGZw/7Ke7D4+cvs6WXIksztCxxTX3MldyrkzCRH7ssW5lro
eGkZIqmb9lzHWt/Yij0EN9aq3LMVRIP74IMpQtN4Y3PRwqquVf332ZkfaX7DIebq
W139OnrtQJMmEtXBSQ9qDEMwkp5TaTRipAmPSORA1veBEJEbnLdYS9uFQkPNp/ND
Jc726XnaHKbqhQHfN9vn/L4JLWqHbJOuz/oqnzNtByAniI5dWEZnNbQYTLJqFw5P
JRl26bgzYCFDZJca9Hee5OufWKwtxfENI/gWRA7V/QiwpHXBzZUrI4KorOP0VAg5
vk24nEugsPrtiY+boGRdDLSQwAtO9WDaRgfGRsX/6dclQe08Q2eBqpsYqGGbxDZz
5pnApnJgOafeLgr/EnuvWkdtMAK6myxVUTL6fxL3pZRJNkDBOm1b+mrjJDmc623j
kHtFun0CJ5KL9S6CMGGtJmDldMkJQ1SBskLT84g/k/8njS9mtdKyZiLb0vkD7Dhs
rKrSLUXbFlf+uXPhYuMRwZgzgJrHzLhkYq6KOqjls8l6Na7eqpIBrHCrmXiMSOBa
40kPBbLf9UwL/gfmrFNdU1DQVMGnPuNY0Nm5bshEqZw19fd4YRkcIsqTFksi64y6
/+byqz5vHHA4oq1ttHAfzLpZo7dCOJ4Og4JsXxSW/+tcHMKBruqtb18faJQRt5pX
YKMbuXJTdXA4j54dNGK7pmLLFIKjxxgo83zYZuo+S/snAaEn+1y6KA3cM3FtB8wi
Gw9b2sGo1cJ3looJnSt+HXVcg2byYHWkk3lzzUHfKLYpsnaIj+KCdrgC8rKmLxoU
erAt+UFt/ztQchzgNL1tPyw2qGE5Vd9F1UDKxJopvNYLyaDwDhDbG2BfXiWGizuk
X6UhyhIl4grmHg5Va6KIj5XQCPQuDxIrI8ESw2EMWp2DTDycVE5D7hYKI9lbAbOf
yqqYMmGQamia6GIiwbzDVwa9Vbgao2QINvPOTyynT3cTKXGgth4x8zHPt4dJjFcz
0+XRV5gDyK+tySY+0dePG7qAM96fQ0/HBTTxrKXlfQZsbsCe1dEdqWrL7KqD9nZd
ZXc1/kO9t8NblOL/JuAnbKp4DIhFc8Uny2QOh0dfOkbzvD2+uvLd+Pb68yEuI31e
xu84RYSrubmsyBonTYepshuu6xgVzR1Wso7thutm3fuXqSAyAxb457befuMFgnJZ
IJkdyO6LV/A7CqZjZM9RbwvrEdRLcD1BZlHqmJTAfIG3T1v/xD0xmGaFdeKup0Xg
LvgjxgO+EfwWDFX9xMg3feSK70guu25RLhb8Uc57y/BiuXDkIGHUpTr3+6KK2wf+
cU8ujVF/F5yEb0OZcSkBONrmA5tYTFDCix+g6WwZffjNvHCXh4hSEpmU5rCPK/0A
0Ak+zqU5F7ptHRp+Jozqb+3QbxmmR4zO1ziZMd85F5E9sZri2pZdCmLUKBXmcdO0
Tqo70RTlC6GoMh8zEZd7BizEASPWZ18znUV+CiJj4pN/BqA8fgL/yt2Q7RGbjnsj
qMvFbsVr+M9vsALGLk6HMjEDbCAAbLJXk9sY1nKIXsUO25+n9nF76Xz2khMLiU27
pllZjKYfpFV4j/73xJ1b3iQmtPuZ4kNvooVJS73S4kptSmhX/V+CpTIzOf/pMwP5
rdQdE9RDiJYRnFVtmIiaTGrVv6bFR3Bv97kLjnoTD6hfdVcnNnkIhHK++qZfadtE
Lz6DNMWShtCLJmCRZBVLv/4jh2/UoGp+NaegQaocWQQ4mffJf3naInAd+hc1o9m4
JBYWwwOunxfHHoZi1hxvrcF/hjxiYHE/U4Mn391gHL4iawZyG7IQVj+lqUq++Dt+
Q0Vqp9T8Gh1z22UFcvS4gTD2XUGRyJ8pfcyk+t/M+vFH4QjeszQaVjP66PPri8ap
ykfClQTrVn3rgfjIwX2kUf1Yh5JOitG/FzyJ1GIMs6vlrLmyfmjkRJ+Yc3NIAaZ8
KGhwu6lP4lKaFRplKtExynTKYFrzAFnlljQziwC/5tm/rYtgUuO0fHKWYJPRtbDe
BjWpTKusIweEkcLixVr2Zj1CIdvPIGo303D4HEFJxE/IuH9jYhpWFOgiBxw0EdUT
PxyE7OYStQsGOX3PEOBaXKI/j+tBA9cdBwsEyRRPMdcpKGqAEWoPBo3nFG4nBiaf
3dvHa6jgbvQwbXeXA8kSPtmwT6/9nYDF0BhNUPgoKBK4XvTioiSt3skbJEbb0g4u
SNIfvNJH8C6tgRWrHHOXSvDf9pTHECaHbWsMmd8NJf5WRZj4GJPi3cxbEBttcrTw
ZgvPU3GYx5ehX7jH9pbUibyrozb2nOdPMj8Sh+wND3QjeDXR3v1S5asDRK6gf5C+
bG/4+myOv9gxm6yHevavuqShZ8/3rFHfdOXpgMRO1l3vT+X3rNyfiKdSlTtuF13h
PtCkX7kHdTq5AMIIHicpBj4J79vKHCobIC1ojvrqY/GYNZSO2jNh7rnVIfjYWX+I
PWjlNVl4jtONppYi5hXMP7XI/BmY1Z+qZaFxhagK9SQXBMttvjkNoPxYsR2Nhu4a
faFjbUYx0tx50tWIq0lMS8yhytHxHGWtN8n7buv8fHPO5AT+i1EEZf1FgvnlXazA
ClUEg2wsB8W80GfmLbe3uvv6D32OnJlMQBiPAA1tr5okG5U6LeqAsc5HCPVU9Ymw
kc8wyl5461LxqMepD4FMmK2AA5031bDSDm+mKZhVUpPPE5whZ02N1dVtuWDkqvaz
pKsble8BdtKmEFc+5S57FlGQln5wtkapLPrGvJs0x30tr5D+fkfvQmb+0kQxjtRG
U1Fw/Z8nPJ1xebfiB7xsJYBGg02MZFqJNftPeRCNj01qCtKOBP8VzdjRI1WlZtl4
NSImI5JhacRGm4aXUkSzX6zHHvAxHBFqXWtWYNymVlow6Hp5G3vsnGQgogqcHTpD
RmTNMSsmh1oZC6RjAyeS/fnt6s64wHk13LP1uKw/2ZsF6nPznATSY1urYk/8iD5z
KYp4DpCXqSEGN+x3H/HvW0/MOyUBehzJh5sD9Yx2KjlJ6o9GlxNF37+7mEKAe0kq
qcEWb1y7U1BMswkqE2y3mcBzPFOs/+OOc1A0sP/UhT3cOLqsW/mYMLJMVMd2rM/A
iWIsdxLRiUckomIoZ9JZoMJifFYjqqx3XIy4rKXoP4J8KFITMC3IVcbHp/JZC/3v
ZLu2O7YOGFHfV2gFuK93XnnOkS887FvdhltC+V1N7UiVLU1FuvlK7dBBhrcR927d
J1eOUQkik7xP9waOKzl1Y5o2JaNCjFAjCu/+ViHTPfofXJjrn9w/vx66EgSf7omV
P5aQjv9i+sJkVQhtP/WZpBV2lMq/7jZ7E/Olldw9Obphtv7/UaV58JQm6EVGpgr4
Y1FCSt5aMawpSXEnFsCiNMW4H0Io9ONNQ7BvxDx0nS3+XHRMNEl8jzQGuigRBJrt
U3a5L9GvwLTrTR8ZGf1YYyqoupsOCNVjhr9eu7VBE39YPBoJ2zCxkw+DVLBbwSWF
nJRd3bVYnD0dp8lbqrfxWO0MOMeD6Th3XS1sObSj7mPsj0/dLUprSb0zXVGQc9Wl
3wddfULvP7IiP06gBd/on73+K+zbaa3EEZQHgGh3kSZXhyNGRvVOObqy27+mI5/I
JzKFOViHOoZnlfyB/Cjqr67s1dg3GKqbZ12sU20Zc+mNHeCGeqguZBd8igaT/ODL
ZvuF3ID4OEiqmJF1n9tokXtx4HVmbD8nXRUhzoi9zY4a2N38UA6Njvp/8JHcsEqn
kD6rbM9cIIcvvntIVLgXogiL8Q2ZoGB+vgOCaxfLUkAv4AJWqynOszbth0Xi8RpP
jFO3wfFlNHhlGmBpjxsh82KtTJmHCsf2+/+SUBeHaCPAM8+QIClUAsPxBYwyBDWS
ogIWpE0N0BTsdvA7h5ABO0b7Av/VL9FNZJcbaQHzbBMHasLlRnTSm2NBUAQ2BAf8
IKIG1T2tdvtSnU0pXHPxRpFV+LHpq9ryQXcw4iqmSvmv1QtURLIuFAfI5QOy8iYB
rRST1rhZK98wF6zeIcreFVlAiM8Ng+nK7HmtpIJ44UDnE8Yt0BLOiLkgmFEw6Mq6
mmYto+rUkU9VbCBSkkmV0jCkbKWFCYoKRpp7p62vto7gC1s9OnvT5EuWhP3xsL5X
q3wsZIGRWBaT94CwiwJShX5KCIwCWCnehVb56oK8n1Q31ipYpSoNLUZW/GQTTrU/
2nqLFk2uaOaZJboBYH4ftDslS293KDLVbhXvLcEFkLy4a1Wet7z9U2c1Ipr5kLRG
OVguei9tChlvE8kx2KueG39J0XMTU+yehloIHtkSiZuhtF/RGGfsEWj6H0+lL2mC
X8gUUeEPXJgixFTaVXJK5GYYijwMt/E4l1wJJsvcub748kZcwnuMGLvsy7wj0Vo5
iOjU2a68Zjxz939z/Nwd88q5/AQqf3vW4Gyloy2DpMVZe4TJ3yRJtolBGr2lBkOp
9d4wbSjz5P5gJ1b9Z46/wkvf3duVu/Iacd9LdXZxD/7HB2SJEcRAIgJVFiqlGlwV
BxbGlMYtAE+afn0+X/IZvLTDq/fjucIFyNl1BFwP1TQGlF1HA968MWkhyAqBFs0/
m/ljq6wkrz3nbvAlJ5WjSQBofYz6FHX8cZFcMOcS/UrBWW0swvHtvfW3KSxZhCtd
CbDDwFv9o8qDNLKkVYkD6c8O2BNUzy6HEJCUMukLvwDPX3MuEdb7KKHJsmfh096y
//diCb5BGBbIt0QSlqlsdNC9zNn9wjZqryOfY0kqynYOLJyPSNU8IU+eh+aQ7fLI
zlrl7oDfeNCOSTb8Qw3PCITzGqF8L7aHHE9nQ8cWAwEuhsimbF0NLYOejmjFTUVM
Y0a6LDrXbO34UgMoTG//57KrwaGMosQiNzPJxQXjykJjW3ld1r04MtYpVCzbKBLO
Q5DstWIyWeoo6G7hbn6y6jgtIWtCGL/I8FdmzUAqJ5ex9jHxTl1HxA7zoFt54xiR
YbxoygZNgWV5EhxBiIZ3AItmpj4m3bHYp1pzLdi/ET/55DjZ/riMy49wDhJxTihg
uyfQzowlNXJxYLADuNXiICy2MLZgyn+hfEW64K2V/G1C+bYjpwKB9Jmjal7RCneU
+yrMRYlqDa4Ib2NWbxn7VJKp23w7caGsa7IZlbIY8G+JiXZajkspph3SReKhhwRF
FrI5eLTmsV0R7qcbyP1oqlt/+9Cars9Qt7YaEvv+jnLHaVUxTbAL8PzhoIg0Sg3H
Sma1IeP2Qy4Eh2kp022F0eRL2NRWNmPb8Cl1uc/v7SNtBg2dDzSnAfYaboXc5+Hh
m5ggC7GMWWa11k2VXsBqgwiLYBFTz71oKcf8FQwcwxpNK8/5jktiMX9X5o2n1Vqt
YN7UzcNHGSzoB72QnEhjCtGINECC3+tNubtW/ywEWlLC5/kuEY6N6xwOTju3txqr
hNn8iEMJBX8iI2528lN6WZ6TrFJNKQYfZoehv/ctdR7qLwOrzKdu0IV3naKaaIMS
GEFGHFRiJkKEopNFMP8BUZJ/oVRC7/zipDFJNuqqrtPaAH3T+EgC+67xjQEpnug+
chng6NQvvtcBFHULW5fINIVC8y87BDlo1XKDEr+fhw1OWrwDN0jy5t3Q8s1Bxxo2
fMGGDBnNnW+r08szJosbtSrN7a/4m5TdOGBG/+7r9pvUp72ZbsNdj5ipt9Kw1NTQ
iy4Yi0OSiF4fanq+D8bXWCDaPq6aUjKm+VZfQrIyX7bwuF/YoGY3aLlzpp2bdltu
m1FSYoTB5R2W1bRAjEiiizjVKPA6h5K7PbpHZ0B/0dNCZisX1GyqhOF/RZHSvmM7
P0+kpqKHUQ3v3wHW5s8Y7+TweqMMJ7pkyeC7exnqLUx18eYsgDEC8mk3OS5wU20H
Qmy+CYZrGOzU5uFLzzVCG69l6Y9jullzD8fE+7nGVE9FYvLf7hJzXofqy16ycgrB
CP5zGflFGMXkHAdA0gwVTfH8S8BhjlPaXNc0mH6hXxGE2ZYKUZtTeytbF07XRE1v
0HU97JdlI3T7Gc/DMViY6F5M74JqUN2Gp5otqdtwhndF6xPQaAQ4NeZuSRVE4gpC
TklojJKUMsf0hP5WpcnBvY7fkr90jLjHFlJKOWrbQ+dxNpqsFuSAuJTXCLTVrf6K
9ZIOBigpVB0J/kGQjs1DYwNMu72BVwUN/lskp40L0nheicrEqYb9BmfzSpR+i+d4
YAd2hI0fBNRmIfscGMehRO1+pHpUH2zjLFrbwbe72Rdx1uCpbaOKQYq40GGdoDZG
yFxorY8CpCWzmcvd3PM/+Zcv983CqZKwsbsZgiMUnR7yxX02SxVDSvA8X05Vj4bf
lOIlLmwWD+aWl1L1vFW0G+E8BXedE/vzeCFpsgWnL1dXerFmRCI/JbVZN1h3TXal
xWHv7J92eVWS2xpdFysQoVOJdg+paF2oJ9BpZfeQMtezGW1iU+At24QRsfv9xfYW
hYawF9AfNecpJ5c8DxXlT+cUw/8Xr5wMTTbm2UiMKG5B1FpOjA6kX0dvw/cHMZJl
8jEottmE3jqlh7EWVb55viyP01GC4Vaf+rE+/0nOHK9Ga4KMap2jzHR3YBfwqrKV
WnxmxEuJvAXuIhKdo4iBUhcdrz1zxtUh2EFaKoM3OrPIjrxuLNn6wV6rg+IOlYeC
a3vRH8SMv/y/FHe4+DhLGcZdfoDyNiTpQcGYL3g9p/kc/ebo548mogRrdZ7qr21P
yEI0FSeS1BvLIdG+4pQuYVpB3iGbU6LjYYb7gS6i5HsFiZNvRL/ZNTYDnCvlkitt
ZVnkpQSGVWWdq13MoeM6AeEl5AO/HYHkOkFCyPGAmrML17wPVaVhVGeesJ7SnPAS
YTn964BUd4vbAfyxvdaKMvD+AzhWbB3fASogKXnZ3vugkICszfc754TpRV2fvenY
M3nao43ph+qDB2Mv82WlNVrrpjsTrMuaiTzayhXus9PHUGNSOb7gV9tNl5oNJgk3
W6cxVH5c3exccIDQ3X+8ajGFBbxAqctD9A3w8qgA3dqwuBtpENdl7qR86DA8X9Fc
d1DV2iZLroQorSjKCmSfmGXtJ183vHaTdihAtOJE1h+kbEFb/eo2YGE04q451Ex3
sYD5pSEfkKVAp6+2UJ8UthjczRlEeukA/EwohbY76U2P4MwauaSQA/zXw5HmdeZ5
dIy0rM5AgiACJYpgcEMkYcMZkmanjV++o0Zrt7ngSII6HM8cE/T/koPwusvRBqO/
6Z7xkZdO4p1FwMOvm8O23wFvCfJDetk2zUMgWLoH7HFDEGMng/pQKNSNeKp3eSfo
vi62N+62seJ3aXrGhylpN6MH2ioclTPUfIC2V7CvD/PgPjZ0s+lcZneEkur3BzPg
8pUaXrWR65iNy7cSuwEQr5ZvI3vyyzuPsuAG4fE6IFjOMIlvt5wAHSKyhLuLIg2m
1SOzx9KPau7M/yDlC7Pl/aOfiA1AWsGu/wjmGAwSetTeNSnBXprwHgsAT3XnhKuz
BEEnCG0t1Hma0tuphbW2hqN+cMyNbStcP/XhjlKfFpMWdTx63bamYIsNVaZrrzsh
pfJMvHk2jLbSqgEdUzGLBIpX/4RybbLbe8TUCqxvjusiT0Affglk7N8kXrbC3u2b
5as8wRo2kbsrKaLnzD5e5T3CdxnkpfBwiuam/kRFkBEO6FmhwNYXDsGwY279MON/
dW5gEDqp2n2kRvZ0ROstcBkNInN+f6weuLEmGHmTgpKWgYY+K5HdBJy0agtzICbh
k9OP6w55pfYDKiZSX8RoJEQ1nHjvThtV/TpQYHNydsl4ZoCHS7jWPrweqA4tvn1e
JRXASnJ3Aoa7uwkxMk53OtF6pMyAAot08DdHPKcGNTXe64WGqs3Gtg5E+a/c3a/V
LIqoCXYLG5ZC6tReivoAXHGGuQ25JMmPRY17qeea3lSpZzoMkf22fuJo2iVjs61m
rxa5mJlwZ7CBT1lK6OLYYw6esCy9tyOfN/XE0vqs8QgmFfWQrkdMI2YhKr9fo8vu
YYRYg8qx8lNtzHRt+iCFCED0lQqHFH4M06e6XQptJZ2n5t2lxEW2ZA9fnqOcmaUW
9MBSZ+H8NMe/680E2sfMb8CO7EMeqR3DW1rwb4WKUP6P61fX/0xVZ2EOIrq6P/t1
34rNAs/UxbZBkDWvhFcH3uksxPieMu+OdQbbpk07rB41WJ7vzvkjXpqYZ/efRFQs
spr+/e+lSHWVrylTWCoUICfIH01qJQcbZb7Jf3OfxdvJ+ynUoD2vh9qDkaX8iy2C
2Og921Ri1fQN6Az5evpXcJ7WVKX9R7cRp7kLSCprkzgQvGCG56pxN22o4FsWb9VM
gFvdpGDvabsJsc7mjLCi+auH10Hj3e7XRXUJb7/V0jxdTfdMUdIQbPcv2Wfq+0Ed
Mmdy80RJ3bIhgG7u8zAFLF047fMxho2XAA/gBcTz6rPNzETFBbTyVNAzjleYqHvO
3Swk/8/FBYSbb4oxXIrvxWwUvmmMFRaHRNBysjhIPMPhr42mttTKAPBGgj8Pktmp
+f6+sLPS82pMD/z3h25FSarPeQ0HZDElrDwkiXJfEGkmkd2FuoNuGJNIg6LJ9oyZ
N6edyguLTIhQFISWGre83SElFrBiW+DbdyZkI3J6Cm6vcXygoHAflmwGAOazH86z
ehmlGcULmttExZzduPfdP/JX92d/ebwYwjBceUan1RUJ9RBnk283PSszmg/FgzuD
Xj0xUvQQhyWQZzv2pyFOCsswDscKWvbRfe9VAclK2B1+g++opBiylDlnlUy+qugc
AVfcEazkaC48NzO90LxapAOPtvGhX7gO1yWoSSuVFn14VW3q+7M6Ss5ETvmmv4VX
M9oyYcTZccx/F27WIWgtvA6WiRlVYsvx1YQWm8HDHFs/vm8Cox58MPTDH4xRrgzG
FXA2T7c6KzjlXW6f2eoEMXP9XnVAaJzvSg/P+a2hDeKMZy/2mxweFWISxMB7gwIY
IeO3Facz0Ex/2F4TmAXamlkaPG832A3MBECGjNI3weI6gfgQzSqgpPOzmTkbmBpP
Ix+lsUYEztBK3Wp2DFJBJUlepHdbc10c/Bx5wic6DLc0h5xUdQV3Hp/0nEZUilJk
oQhjr0zQgrruIVetuqYAhHHgrZDxkYZRVCBD0VHM7gd8gUd7izJayv0OFe/Sur1r
rBW7Z9alqGwaT2wWTNUXb6HB8d6X7n9HGdAFRiGjMQWHSKaz0RZr3CvZyeFxJDpe
ScjNpK7BhcSqybvucfBu3pibWhvCqyxwro8K7gh//nR+ae989S3rxH6kRV2S2IY/
ZgAIkAe66rs10UJm5G5l/9eoWJX22McTVT6z7tMZGolkP1X3EztV40ENvciFW7eg
muYlZp3mehVGxPfu9ebQxPHJn6w78QsvUXRiYVTuMF+LW9OopfGf1PlLheBdjfQq
kcEvDvCUz1Up3f9csjiGUbSa/1+Hz4T2j4wejDowRc3SPicqGM3zrUXYf8yIjpgC
FaFJjwTt2rfQk9shKtooLcoVQT8NgeyMcD8VXYikq/vj5hU5fuHT0YLOgdjUhunu
kInUfraf9DgVXX4Zg5khPnLgcQivLiOD/EsqL/P/zMhGcdObJ0KK+tJKojo66NWU
zpmHyb3p5NPI4yUxL4ieI+8WJIMIOHMqsZLgSJ8AR222+BPWd+8JiuPW18bXeVrG
09W3OJ/NW56i2JIVt3j1gKaKFVc5xmMVJAIy70FS6C6vHMQouRqFDF2Age4srAl5
5mVMFjGPovUzZT6V3K8M3C/RvTdvVuoh2Np3xrtbmNlzj6d1Rd5FYmuBgsaMYz+b
RGwbVkqHdMNYnBVbof/HO4kvAROZR0FgM4eNgPV38tL8tK/m/ckI9gbVI7s2q10L
+R9YDdLH9c0+H2dHD5v6T9XAsIvQL35a+vKYfpLxQjP+y5arFSCmPKzgTR9gup92
YQARSJXbdpgnMXpRvHEqCEQys1FVs6OXUKLDxPT0pmT6Xxk4EHu9m+Qqc+wahKbw
1vP01FZi26/mNeSJ/EUKYOx87Yetb0YV49MvZAQGsiLSS3Uq+zucaEy2LA135p3M
gpc3g/mjyFAn9WI3xHdPK70HDlvtzsjxzFZ1gnU3sC/D/fC2zhAXspWHHN2xrAiA
PyAtFvhPxrzdKEQ/l7VRdBqVS2nhP2fsn5Uqav4LHAjoRerQoZhcRzm/SBrs9U98
5mffrVbxQxjwqaHJUo6RsOUJhZTSM3M97pki9RQa4WQ4ff/uUMwUkVp8Q5I5rAUv
LZ1pWzvOTgwSWvpT2jvfFUpBE7Zpa0G+9SJIXAuq2wxl6SZ4f2N8DVcFwFdYndfx
5hzkPlClRjsI/VWBc24jTcoBjmotAVoKVvVBLngS67qpnphaOGRkeoq09DN+sbAP
dguHjII4twXQwNI1nMEk0oQEBM04ngk/jZD7A3xdJvdpwCoVD1NSzSpT42jhNaCg
au+Vw21qbaYh7EkqOaUJ9RMf3TZbd0RFrS3QPEXze/tBVuYfnw0YrXA15cxd38Dz
PuhBYDiTqpb8Y11AumSn6ZFWSgXaK4d6xV+3Qo62aHmsDpNVXDAI0muO1xr1fE+i
18v+Wqt0rl/OtkidgLSrmggC+8UInhAtPAuWPvAsEb85uJt0ZJbeCxW2f6AtEB7G
0+jq8/dYKLRQ6FKGY81UoaHdQdPGtIhocoSH0FwbytTjlsC/U/bcBrHhwO6SzyQW
v80hcVrshM2xdtaK3JvcH2YTxikeqR5K3FAhlBKXgqII2lqqHnjvK5d1Upcgf4+e
PpeFRbOLpdJJirujx48THL2WPFErBsCftjZSI/6cqIPwYsMxA8O4W1qeJXc01iKr
aRLDcJgvljObIUjlzv2QUKZbCSV/hOGTbrIKnN7lj2wEFnvZlixo3b8r+FZoci4h
zclv9Cix4dU5ghcwkjCvArBFRgueWEoOiygRjmIWn9Ql9u3rduBiKVzpzJT9wQP/
SsGpiof0Ks9V/jH471QXEGX2mb7qKmF9TlzzWIprLT6df3PsF9I/Fk0WTAPKUviJ
5F5BdGcqT+unUpM2POaDUl43fW9TAPG+TInn/hrGVMTeLMSKKeGSUqo0XegCvSwW
fL38sjjTjhNmgtZFmZ9CuvhXN88L7mngrN5t+/u43BrfDQnHFA2zTeM6I9Q8GJxs
euzckdn/eL5b2jmNZkwqRXsHn/uAeFMWxI8Z6Q85NcQiRl9aKg0fmqBLtIp+yghl
3WacCCT3xgM6TnMCMcpVu1mFbdTE5BIvdJTlE7xjR5Vq5YRAikEVOQ3XAq24twXg
7W24rgp1GdVLb8WLoUBGqN3UL9Ya5RlK0cL0MzadpPOallnc7YsJr5x7pCFeSlUs
nRSTx4FXFT8b8b0b/5VYcXP8pf18mYFbab2t+cWxreA2657e+WCyMW7zUa3q0LbH
ff0vRKaaOZSUFLjnGWISSTnzg0B0Xutf0nsjIa48SEmEceQM2X6uPDgL/MEwQjxV
/VEP5cR1+ZnOn1cDOFByyIaWwXDJzjMrrhKPL5fn9zGleNVdNmvx61jMjswdlwMn
i3yb/kjf+tKHW7hCfIoVv2KUZvuKUciB6QRJlkRuo8T0UvUOAlPEeMxUslDDrefw
VivTpV3SLVDAhJLWBYpCfg0EEAY7UTQIrBmwRXlg0rGfkaTdeOVj+8GSL8RDeMto
zWdjNoyYDciitvwad3p+y/CzfmmHxvz9LiqUwkgB/hRgrrNen7U3fRXqezlTEqdw
tiigiqGyTDR6rEbOSHcjDVgfZi64mY8f4NLD+cjtsQc7l1aN4XqJhAUEwJaKCDFB
oao87QojOUWn7pWYPgr9rQ3+l3zowIpLY+NguNIdp5CMv/HNybFJniQOHusjlFms
L+HfAkU+82rll5off294dGkzdfbylLbBwhF498PPfC68USK2hjhkQBtDWcSjx3G2
LCnGkZA2A7zMcwyOS60DnxZtOF98mGunAQ31EyJZoh4lX0V2n3OhCi/cjZhL+FHf
2ocGKN3dDxOwBYcguPqpXx4Q7nrmSvRRm7QQh7lxYPbB2NlFxiCMqyPh3szsNOec
y41hYS+SL6nH0uKjCXrAm2grNV7hmk0olTzszjrBgRppXRZpXKo+Bdo35XOTaRO9
scbXTVNdiCk9GUd5bXvXk2p264Qzl1j0RxwAGpf7jwYB2YVONUwRNP+atX9YagxR
Bxkr2nh8BuRbMmK5koTH0o7yPhvP96kZ4o3HIi9l7IOrszZXiqmdPKoP1s9yZv+k
uptrzbzxOSfJKBhb3v8UnKKTVVhNZuqX/x+lb9CGVzkkgJCKK8I5m4OZzesWPvPk
Yyh/mv2R3naKj2uFGiHTO8JPVt3BFm0BMIPU+M6gETbwErIAyXCu/mPuLHQOJDpt
A3huehA8fR111598DoW0nG/o787tcxBZ0SONq+6KkojxDX/eYkKAlBXdiBBWRkyF
IvdeluYVLMxvmHBO2tcLXXT814Gjw4jE8oLHmefXrx/ZNOoCfV/ou+v0wglII0eI
rwiai18DrVNEaGnOREMdHlV8kiGnZDsDv+ODVRcbTWEm5/XSLjsT9EfkmmfIFatt
dRI8T3e5/+kmdONSrOJwb5rj0Z7whSuO01yjHA/oeoOeyS9+hRX5nIx+JK4e/niG
fImYAhStDXarhvo3/HxJpcNoZjEu8EUsI1shQO5vm9FAbhAZ+5X5rGHJhwrzqnuQ
vWLLwdcG3GZo78QUOEwMYb0ggdHK2DS64zt+YBk9uvNEU3QlzxljIHQzWApe6sod
urKZi3hshXTH6blxpRb+kI6K2IeGrJf0rSoTyH/saHEqcCWSlAcRmO09aqyFQmT8
pe25nx4yjGCKzdH72gtFiVCjb2cKE/L05vI9YWRTGjTV83d3BWMJVqhb2FiypE/A
GeF0D80JVBIyXwZKfC03njyeAhkODpuxC4IMD+N7/FTMm8ENS4XzsoVplvPEqmtD
kYPwgQQ7NVl7Lgjh1ApZwB0zeXn0M/qa5uXeoh343MLeIapHp8MaN9R5IxnbabrC
g4Qa7zJ+o6D9qkvq/d8VNlHdWNmdRMBCS6WSjUKB9BDpZbkcbBbG5Uk4Cz1l5K7F
aQ2Dt2e4J5kGCasguPI1Ic5U5wpnIKuUob9SgIvro0qTTDHpokmouv14sRNEM8fD
ZhKgU8JCwMmlSpPGYEcKtdBWDjDpmOOPvIg5xMiWHbIlZhqX2dfgzxuxuiICHEQ9
vxY8WYLuu1BaR0Imh7awhh5yWjA5S9CiK/qDSF9lwQXNC4irc2sZgaXP+Nj4u5Nj
BTjOJRtfov0AMgzVeXvcsmgz7+8TkHe4sZqubnha82pmDR7adBgKWpkZuh+2L2RQ
qN2fDWbR4L8bUYVmipvUGPiDgKT7wHq8f6JcPfTlKxCZ8VRfH0jRbfu9R5ggBEgx
0cmhmgUUaqD69awBM+yrjmEyS3rFGxUo64pE599aJnO79BEshsrXhehBOPWjpAgu
HUfB4AIt2YqaJx7FNn4QVXhzJiFADVAJZyz923dKnAgOh53Jl70E1bpRfm2tx5oI
eOdCb0kGVozeBF2Cli5+dS6xC1wmDGWk+jLSXzCYiBlUwg27eKOj+wWVu/w4MSDM
crZsQQ+6pQxVN4pGknb2VDISXz2t9BM3//d21wCjwRITqczo+z8p5x+o5IAm76eg
r/U6biYHi0HGz5MLmCylXzT5MjKsTajWUTN4bP4yMbIcGUM60fhBDuxhqt57Tbhd
r6SgewVl9ZGPYJSUdt4SfTEjlxQIeYTRfkXrSvXuLlhL55aXk70wX2tMry383zJE
bPOgwSzVRJFIpmdB+QucL5w2CqQVxIi+HMKLVyrFUcm7S6+/7RoT78jT1gPYDxj2
ZnVc5ouXQtwzvhhIJlxeI+Fs3cLaZHQbCzefRaptkXhoWRsqwssUUO/E/grlLSHh
vm9M3jCE5L+CCFk49U49ChwqZDoC40vXCOezWY2De+PiPIO0yveR3zpMcMRvIQD9
W8ffvAKHtQHpzLEVVZRL990MA9QtHOVFzhcAjWBM4KNKpr9S/RsLRnVI8ljrhkRs
ov0+cAnqNIT13Q157dY+CJ37JTXsIip1Ja2lgi3A38DMqcvLRjwG+fzjeC8cLLh3
GIKrakD+apU5jkEi6s5TfzRbhhq8FQRqrKkEiKceAhO/vAoENUq7OFxDZiEbUCpK
STEeUKQmBCdQWB37mYbRE3RfrzXwPI52r+VgR/DXLxjtpDsNrpqANhpEB6O93C2X
cfsoFcC591EeqF5yDZaikzsTlegWNBvQhRcETfgL581jA0RP+/wBPwl2wURWn93N
lhN+YB+sRVWzACx7P75phd88BHIMJxctMbrCJ6L7jEVYOI3CTorkAM5xHU00qINA
MfEINFQUPeXwNJLopqJY5n44OTz889uE/Spxh32vQE2i8AOSNTPEByIG7FCRGTze
WNmacNWXo4LI/wfS1xKFVgUg2iuMZG+aJzSChuIODkC/5vPuwoJho/ZgjO0mSwm5
k8Kj6fOM7L1QSgfuCx1DELNyEapkL0I1KBPG4/G+P0UhcxLSpa7Z69oObifUveZk
YZE1yxRCzGdfoL3dkdWifxuW5uNJHZChHCrjQEfrM4KGz2VfmxbeGaOMblF/3RxF
GspzLQTitTHc01M7wMAXlC/63x6dazgi3fGI1/eaPHXSU/R0p6qkt5OnEnytZhnm
qOejsfq+Ytk5xetslVdDjUZofedTaLW0xyLtGN96r5J1xmvD33pwMhk/awIeF/eD
j+hsDdHBqqnnkfoRnbhY87lQkzyg/KGj9Kl6HGG8K/lu//5bWW3yHo0fObpm1aWl
yXtA4G8cr4UM7Nk+6MajppEKxiFL30srg1mBbAF8nfQUICMw6oTa7AsDsoBk7z+d
2vmcUu2nPvmmKUQRfQ644HPk/SmMbYXCKsX1Od41cltLvE5mQcw/m9RYVLRg1GNN
26GhLT8PxDh0tqLd+TN317fvwUpitap6gMsGOMkb6l414cV2VpNBcEuv/xar+grx
d85JL21Co2FBbHoLYNzZ4b8yyxW7C2pSp8kDknu/NGovlTCcTIDhnZ/A0NBAJhOO
02tMY64PW2tbyGX+AsJFNxR7VnfALbQsuM9ZKkr7cR2uccGz7cUR/4EwTbWCJLu6
AIEZ3kitjb+//FBcRVRHbtd91mi0VGrVp6ShvO2getFL6k9IwYImmueams1gjzm0
ajTJh8qk1D5rSQDTlAJTbhcXIBqHZ0wVJ6sQ4XlMSzemdnh2ca0JkOwouC054kZN
r+J6QrIuTJdfHdjCmKTOybnRzIKT7K/bo1p+Hqbwj0Yw4QAJH0YIQWYbX8tvCb3O
TcE8vmfDW1YxfGoCBK8mCcriwLXEFtg+8ykT+Rdv/evrdF5TWFV+NLtz36IVvHnv
vtSVf/hnvGPOzQ27SDkzOHnuGDNl4etNnZTI1qMOBUmUhHJj/rY3zHQ2B7zEIk5/
rycOq8Na8HtUQ98ja4xif92dahXq7x9IYjBz7SS6dT8ECMdrt4wA4sL6yH8dmorh
kd7WpPOZ5Cn8pNPYkGmYA3JII3YwKro9Mz/LRav6qTHzTpq9DDf/h0nD3Z7IJTnU
xQC7LQG/NIXl4uio6czFKNLIxx9QjNWjh2eMll6XQsZl+cVHAKDzqb/ZtoxGe6T9
zAPD2box08vt0hMdGlVuYb/PJKOH3keVct34sr+N4Ti4S6XNSdbPOutclLVOUfsj
pzijeyIjzL2BWVCth2FM4/v5kX+Fy08FXuBIqhbNSWjBhjI4joTiOf3x9ROYm1p0
YMvpsb6VyUox0rydzbxahVIUXDiYlDrNFZJO7B3p990G+iiJPV9m3xL95MT+8QLV
UciAtVaVBc3vQvgovcE2CJ9AgDdQXvwsjj7ln95SemYMMlWQRpp1K3K0Cny4zOwV
Ta0X5u+8UFYMoodQpmp1Am1ztyzP2x0aLwD/bUNEpa9b4hBhdoXI0regdUZi2Th5
uDUS01WfVwnpADe6VEpdM9ztPfBOizGCUm1bj1CQBLVeR0Lca6Avsxxhji3jul4h
P5gICPQVZu/aAEaNx54aFT3X5ltOYJXvFzn+iDjcpikYrar4W1pWk+HcLoxQ4+RB
vPUksxc/2FYAt3R+ROIWc5l6EuW43poxiH6lOuvucbYcyBzJgwwYKldY5co58oTn
J7+DiQXWSTRMge008134BwfqL3QWkjMzJeNJFPIjOqwSdivLHvdFTsmdJuMA15Ik
z05ygTrt1Z5NQ8umqEC4AsfncDaq2DrLMU+cA2l5W1SsiDZuWZzJ1grsW6vT4O2z
mS04Pn70nb+9O7GAnAEu297WfI2Te9XEyAaOZg/YRH21MCQ4WuMkwaY6sNKdEVG8
vREBf4h4bRaYxKaYU19UyNiffxWR5jo7hMh9hVptaGzRob6twbbXT+2VRxdyuvYV
LblQ4yaYMRbnKSBtaIXryx7CFAvo4A7BRZnC/FZ6a5hA3VdgaHLWbCyEzGrgflLM
wYckp4dw3HbrA9Qr4VOmr2nqepyTdjTU9NnEhw0d2tgK9FT0BzvrD2gPrNKHduI7
HNFJlcGMiinO24jO3GgRWGyUQbEh9K3wpBhpuLFiT+2sj4PTql4p4DqiQyAJSAql
spr6x5cxVR0fcrMKhwPvYal1ZrMHyNlw0mJ3wXpFojZn3WEUJhIWvzh3EJBFjIWl
Qdpu4RWB//N2Dmeo0RLamA7m50043Dvzosm1vPRnYmoA4w2+1WvvK459xcGdDM/c
/U/1+KduOYse8/QzxPaH46Xrv58/EvuA342gBH6BAQlR5az+LQWUYN3MH6bty53s
Lf3xoxAMe1AZlU1PDsueh/2qY/3B1xvdC5VF8XY3loDQbkIS9rTtjkAcCDPUDINE
nlMiC/fcpkXv1H0ee6AlqbzLijPwMsRiHQGGEXRWWmNWh6tyJS73jSYCoRztjk26
pnmlyaXFqvLJ7VZ50l2iTYdJ0dYMD8L7hd/7UM5bhH8tKMZgCAr7PAVvHmMukQds
578QaTCGhW0SDo4w/kkHnUi7OWa4nN1Fr4MHsz0exhiptZTd2sCxRdnYleoHRJVe
ioeQDzbXR0wpS6LDsZYrF2YHQKn7fDQ6teiDAcoqRZ/733jSBpCbZTjIsY/xgrrc
aqvL8AE0Lf35ti1ZbIXcNR5DjsIbRcU5GPp67yiMG13q2k9QZh2DxEC8rLf2QOi8
vKoZihke1SyTo/hcAyG2leaE2n+LrOGa7v8nnAsrZ9FMb2mm59o8A3Jlnhq4h4Cs
pgqWz/bmVeaCWTxIzjOw8Bl3R3fa1vAHIDvdqN27Vw8mm/XVLUDonbBJz+5pKrNN
H0n7ITjx5qZfhqKnLqbtx9c4dIxixgp8yige73P2X1KsMEvLPELvEqkTQKzVW8A+
8kC0lPIWw5OVlE90VdDom6x62YaLLWPUgP+yuTQjTzJAOV8EbQQw7wAcWCHy3BhM
hyJUW91cTkEj4sAXv5usgd9DJI5n5SkdN/4ir63lbl+LqYvqi16E02DJurAHPVtJ
2yoDKBYsEockJrJ4NfdEm3CG7FKy2WhNS/x1xrsF+IJiH0VgcS6mApwN5V4yiXgD
OHsBc4vyv3jnGErCfoyCWuI8uHKG50oP+u8tdk0dVA9K0GXaV8ox+THmYqmmLNCH
oM6yNu2LuDcSxEzEmCAwV2ODAHewW+vakrkIFawqtKlBsv+Dl3zKUHhsoOZwMui2
mLB6PEeugSIRyVaoDhDq5a4SMItMsQWrCrOTPRtgHDAXYSt1fPosidY3S7tJ/b6G
NUu50fB/irOza01XIk/RXCTjZjTSIWFVGOf11LVdE28ETTzJeT70yd0eQvaV0xtn
yFbNwmviNh9eswCRsN1DbSegVgetDcPdQ3LJAFb2TzW3bJGC8nsh7bbrTwc3Yia6
4AYy3o56xFa+SQUkiW+JBvh8Fx5rTSVgikh/f01EqnlAFEQhQJJj/L6xSl4eXMDV
NZDfmfb+1lk4flbTmbYbRhxJ7aNvPa+haYGU9pjfFzSIs2qWrzAGHTDV95QdnTuO
m1MIi1jv770Dyr5fO7Q8NMQbZLxRrfloimkbsRjuiOjPUOEwFAuokJG/r2+ukR3+
Mu14YArf3wUFgmVgz6lXYvtLYla/GjF2l1jCLSXVnOgI4ZrzSMCCj1qFWci99Mno
ZlpcSvxsFb2DEZ1o98NqU4hQPNrbG87BwRPpBCb+9xr6AS0rSUrDMbPBm1yd+SNP
cvhtvMQizOvc687yuV9xXLXZIjlExwSg3Qu658sYUCg+tcUnEyVmlFDXm5gviEg3
fRMMgSPqUwKUjTSB6tf9TiLSD6UxSL9YiGozCENmXZUfOG8IRaq2o8DP/jtdCyT1
fv9L9Zp53is3uu4gSS6E2BYwiEbkBodYgbCjjOREXtjmr4YaGQPXvG7A9GdnjIm+
NCltI1CpSJplyZEcAn9Mbs2coCWwqpptnBe+OatzDEVwQ2qK5kMwWfcjfEYS6oDU
IC+Ppip9QLBdS2CZJCq5WyAuTuJGH4uRxkLPNV7jnhbVLsw+fNanVYDFu/UDG28e
rMuI5icEk6seA8dLXkhBpdBTvwDLlNNUs/Z9p3egPcvFBfl1GpFAjhkEJYEeq0a/
eIJzaWDVmpX6XrKa+UpnKNUbU4qwbQ6lxDYvyxUfY5VZ3oiCUxRK4LroqQ60wWWk
LF2jsNQOklUUP+2YgpvbDI9jt1Z4NSXaw9X3+v0HoG/Wa9QzcXtsKJuDGAKl/EUR
UKAovb9jd1uLBwwVMSP7dZe0YJV43+cChEQ6qMHsipwUdiq3rHL5RSDsyHDLRs3W
4Jfknt7rUirQ73ggqdT4fsUPbiUWLEvwoLJft7NZ0CQW9FR0PRrB/zL5/BR+mhML
HVAK/fWp5NFxJo3AIdAeH4/b/7eBqc7GmSck9KmV8beP8seBvhYAr9vlwvPRiSrL
/RIBYKmmF5h4+gkV7/jGaMrtQ84T1I4WyTv9RizS0sjgo6N3o7R5tjLQuKegZAhl
82Qgj2i+Qkx6p3fQHKLsENJ9pscptbCJgSRPYR2We8ARbWeThEgHasFm9LRjY3Bu
3xUa8byIDXQCId7dtmZ+gb4LeL+shICfhQXLHctHiKYSp3ck0dMYNgWQFgTrrGYh
4pTqr0+yB18qKBuCXvE6Ph0tK4mjuVjfpEuIVOxiksBo2Y4E1gXAh+Q+uJ55M9TB
vZ8wgWvfX/Vf8vhfs4qNKd8pAQXw7UlSQ5P4wCzfWOJujPUm+UGEdVj3HjQwbY0A
RpubvdnsYNZi3u6ExWZY/jBJBOjMivniX5rxWJsiNmnY5WSQCKRGglHzp6InSjiG
mQbeKLAQJe4zt9kXfy/Y7AlIy3LTfG0zJSBOMZdroEBrIIjEELdvfE29zT2mEdU8
7F1irFgf+hEo2ZHgEw3GWUwCn+0eaa6RYEQh+VhdUgdmDMuSEKALZeLmXGdf9k1y
tL/4RDzWtVthalbcAMV0+QR3PXWPgugw0hROh0u0fgI8Ihc635eXevNq/bbrvnl+
nQKUDHh/uowBxpPukCSAkGJXIdjHDGqJaZwDJ3C2bnJO8o5o9QmoEhgZv3ZMrODn
1jrKn9ivi0zdGTUtrXHO+/F1mzF4OOnKef/nKypNObDHBjKiZ1xSgayNwJtXBDd+
FyAL0Th7ATP0zThb+opNnyeWoF7WSPWT0eAybBRkjdJ7T2TZE3ThuN4Cj7pOltuZ
AmdhiNuxfEQ1m0RMl9ewLLvML3/CyZXPxfWfkhvQ+m8QjiEVyvxO2t+Cnor2Vmhf
K75vCwUNEh4PQvSo90aglHnYR9yLwbKyDpl7og6TjTQsu69ScisMlr/5nMPEw2YF
mIobQkAGdlWe3qJ4HkGL4ZMNKfl3bDbIlxDJjs2d1K3DiiDX6o0XkDnQiPCmQgWS
5+3wKb6RsFtGifAFqCnMMpdN7BlQ3KR12jXi/trUlojgnmpnFAROK8dzZmuhmfyx
hi8croLwkuyQlJjMBiinxLsMgkn3++CMBOhBkt3iv6uG9QLEWxUI7r+z0weiL5Yw
/ct9tujv0wS/tzI/yh72AnLLncDGRreJn/Ct65q8yAwzRe584ORSUDbGzUqI+QWn
qjteITjmQbyXCPYwSKF4reZ7dA9GXFiNCX9CLo8Nj/jM3ubwpqSSayU/9FW+NKpv
bmfK2sr5KIataw0TMvQLoldGv4t8/ZIchjq9fdPauOv13TtujLpdzcT9l7tSVHjd
Mu1WfY0Q9LU9a7gppcg0VemSYNUkqo2q1jzjWF3SduuBfWxCs79933/OXwd8quuZ
JI+swcwOw9QdSzliflO6ZxX/pCEYVvSTxG7xbgaJRL/Gs3I5woUVIzko/UM/JR9b
ifmmOtpFdmWopdmJXDr5G7PtsrMqwmD/lUKcRa+YPz7gVAwP/nqBcnQ95H/gk7C7
dyhhEpZFNmBwM233Oms953s3EN/yq69l6SZnfWh7sxp6rcTK58JG+wv8neBoYnR9
4hKX/EmResULapmP9FIUcuzkg3mMLSDJgdv6Elue4YR+ZcDWpqbVO9LjkW10TzgU
W5KhPXoq1X+0DfypwVTzv9aCvoXoWi+ZQ896u8rQD7Og6lBDs0XKvQdiwLapiPDR
DdXFBmSPpu+qONNh89L0ME3pRA+1BFNFC72qcGRkOKdEsHnkHJjk+a/DHmu2jzbE
RfJRmViMtF98O1+U8ks2Qa2zZec+oCEJKDsDeMtwffKsImHLpF7D4zfB4QegVCYi
QffduiUfQmHgldAwjP2ZkC26HdW0sZ5UbJIcetzbQ4FQFmu3hCB0VnEmJ4XWHMvt
PlMHvfquqPdjw0eoVPcOyUwnBageKkwTF5oh7reHBGTeMMK6eCVvsHV6DNO1M0cx
DBJY8u6rQ0e/GOSYaQOhp86uC2/C1PA69YJgNgHU3ZozjD4/PUCSX5JbbQK0H1ge
yCuWoLOdkt51NAdjaV+IwzYNCRMw2bwv+8HOKOfNZYpnhZVWnDv2Cao3Caww00Gg
zP20hEKGnKCjokZlVRwHSutGXp9VEa2oRRmuozPVA5E4bAOpYjxcJWykpQ0bHefZ
qE7GQZnYkdmrl+sgaK22jQS1bD9TTs97Bcym3EdDeeIdeIN30TIDfh0k7ghYXmd8
F+RMfjRN46Jmr2PXmXniI5ci3szaS5FipaapwenY/b3t42jL8WdzMf3c5UlfCbNF
uJq59fNTpFztM3d1c413n9I6V37VxSer82oSTmU5P33SkHIwAZiKtTE5pH6hvNCw
QKQEr8kcSV3jnIVY4B97zWrJZ5pK013OhLMFRFDG0PyIeQz+UrOXxe7tGXSC41n1
SQWVOMh481oh2TbCOmLi+NgftjrQ7lSH60u7oDhGOlec9GG7IJ5i5hZmxdVw2RC4
FX/LdzcD9W0FAcP7s5jFQMmB84GDwZs3XN6mr5RkAY852FoTM/Vcdidb0nMlXcQ/
Q7kFKwo1KBQAysAbr2HN19IQUysMv2UO7MYeyvNTbUX8HU4c0vtG2V8M6uFWXybS
nFS9m6g/u9UsKOu+bApsUTkosmHrV7SfoDla3e0XJwbKJyUoZyDeju1BJZgzdKgY
T+DHwaDloM0i2NTbNCXOA1SFCy0RTt0QqrJQYwJs0UQLrymK29w7X2TVrRPzlTKQ
wbBXfoAyZ9Sma1ntuEsWVRnJnqh8jk6oebQQ8MxbpSzSLhkglENXMl8Jtu07kCLc
KCGNSM9tPbIlIvogh0+XUt0+MhbLu9hVXi2uWel9SL+moKaNrWV5SGhfTPFQ4vMY
A6UaKzbdZ27UTnlhjj3KWlhT/zLYk/40GWRGMMm+a7IaHrLQxjCDaX+2ZSUPVCJn
03Jw3Dr0zQu0E91cIUXhrfOmb2jrFS4ueBjhGlFFwNQNsB3gS4yOpxNiT63Fr6Z1
MqsJtGaUM9HyEhXvRbg83iTgDZVFNmGvCBROU2jEMkwaGlBRzG4CElTKvm1veKOc
/xtpsZqvnAR36MQmqja5qM2XuP0vGESrfWMpB/n7LIXiK+63/KbqyqO/vEGscmze
PzmWRLMvptvgYAmQTrJj532sWsPZEVdDUv5FZTxdaVTrRSxB8SpEietAYM7BUHpn
PwxjAKIDbvetEfpu7MzZJJknGIBRDV+2dbwaqWr81YucuZaLUX3+rPL5mFr+iZ90
wxBRJ3wH5TgOflmDwmnpe2+QMQTBvrEDi6LPdWLI7n0dvv2mRdaOZkFUu8F1IAA1
PVExUJ1E1cDab/UwrI0GTf4+E++enJ1/CAMNrJo6juNzgWeOnji9gO6axmlKZepV
VJ4WoQqFVAb8DG1ckf7cJ40C/AzT+BzwmL5UoowpBIDcyJX0vgSgvg2rUaXHRa4J
Ih8w+ZR2QcuCx+T3Q/jY1b5fkYh8LdoeWrVSNHIwIW76AycHsbP5gg17gq4c+RbO
cjOQYYjLVL+4AWs5SVaOM+TkdQ4vLpEDIQ1cDdHsRBO5+zot/NBa92QO86wRg5Rr
E2ggf2Y1lP58iLoKPErjyGHPslHHhnf9L3/q2RvVBEbHvmEqHK/mMFGUWx2AiuJR
H9WOPxVq/imghD5aB4D3pqPNK7F19ywmdFhnL0tttK0mpAnNub7XZBRjR9V+lnso
aCkVJjHO1sSjPY37InaI0C3QdAHDScnOVDRLbJUUZAibuP1fKwsNuOgUsczcbVs1
5T277bi1pgGHEd7UCbaGDA+FhTbP4O6hcBHpq/rSF91wcVe6kif2o7iYwdfE2Chf
tTpDKcPpnHztCW6Pn28FcBwRhESz7FVB5IFJqdCXw7vHVulzFDiO2OHIBPTNP0nF
D6iU3gQQMOfRqHdSpfvEJI7ogTa+welliQfFyDJymbnxHzwQBQh6lVunNtlhbuq/
e06Gm3Cos3AV8yhnkwf4UPeHw8Ix4lfMUAHe5J7FOIs8lDHCFUcoDlSmZj4KseaJ
65are0Ho8JMal2qelq71w0gftQ3wctxIU7MXN1zuZsSfRiqmBplmNAAssUK2LNqV
x+G7G7vv5jpjxt2YJkclIeEr1JEBpGriXUddfGAG2A85PeFMk+lZBF8vJGk06h3c
XHZAQzbuHaCFDtLv8TqdgBOvXowlcn+LRFnDajvL9L1P7iG7WNQUbW6EE2edJimf
8ePfEfPuIf5Mw5dGuSr0aHo2Vk5ttGkOOLFTqLbMnZOZm/HeZTcN/flvL1/U9WMD
T1AVyI3rP0mYHniVZmLyFiXoW0Q6P7Dj7aoDAAm+3BxePvOjn96DmsUpJFhRxgTP
yVcxRsiAHDB/INYuJf5cs+hQ/3tUFdCQnykjS8FIqRPDHzQN/IJcwU5hLriFS4I7
U1Vvmhlrcm15OmVKwBg1AQYiSj9lEwRBihbXDRaWs8c8SvuJWNrXxkNcJvrriZ50
ESe3PbLTq1n4GbDdKyOJJaR8Sx+NKH5+QNi4Mq0J9rkxH7Uta2bmtbuxlu4rB91Q
qLDoaYbXOK4uJ35PIoeeBIKq8RG2+HKMkm/ycplro3xUve93O3GiNKcVMpyzB3GR
NMFGNZknsjUKSET+SIbRUHIgJHoWWYG6bZua9ru402ECmmk0pioSjA3YFhdQ47ib
SV4EGa8bLM3dUxb98kEUuwRSyHo34UBA6s+JDTM+lO4ANLEgZMy+e796q3u+MTEE
EbV5q+9QWIq2DK1+8cWkXcRn7jdzTVjL0Nke7wOQiYcSWnlZdLXg7up4QXqd3Ueo
QVqf1xvTA/SowH151gRoOTyK2GSkhdhaetCo4c5uA+BbDqVM6dvXmbmzhl7Kf0GQ
mrryFHcElJ150SY91E376l1RYdnoU/CTiMDdJHASKhbSz362Dwu2VX3wmwOyHUOn
k2+hgB+kKmpUWwFYAnpIWLXBpQCBhD86ZMcsiV9sjSGN26qYX8qNFAWnnv0OqcF/
fxzldcYQaTM2RDRl3d1MgzsmrCUcATJbrbwDX4jLwnmnAJBnusR1jEP3dZvHoeP/
zYxS3WXy7RAp/Fnb+jfAk8CKOexH5bj9YxIKLCAPaR8meAd1t2hdPhk6ybQ6Tneo
xNPL3SNuBO/+wmty/1rO4RTxufncx52iQqSBgkSOCpVgwwfI4pHiNWwj1NV5Ej3W
McELLH2thKuztX8o9UFow3zNlm8CIoKqsTW/yy42rzpNL6EzhFd47YScDULpuGtu
zmIoCxTvGRD30B0kgeeeo488zb07YsfjyO7mi4YIVo8QF3w6Y83U3+/WXT1khm1B
9IZA3zNnxSJKHdkv6IR8LIMh5Stf0Xxh45dNvFrND3pb/BZjmUOJUWPO79k0fSxx
Hdn9W3CoACjCH9HA3UQoWR1qBKyMIiErOQI/VGRuYI/tyZLKE02EOFhYvl9LldSx
vIIecyvwXKcM8g6urAcDzf8C8p0/7ud7tLZZdnR/y/rKrcFRVJcmtyesiTpY32Bc
am5B79xwVGVVslpaaopLGaF6BQDOJXi7tSpR6iCwLvFI72Gu79tiVtE2RVoXzK7X
+Pp+lW/W3lcoXQAGe+V7Lyog7zIYeFRzNN491dOQlbu5v49G0ooSZCCZjZGJ9p0H
F3NJ6cVJuI1m7Vy0EyoxH/knaOYsyi9sS2PNBNNkDigLzKYzVbe8PN6J4mO65gI9
XVOd2Qe4Y6R0giquEa36jMIEso0T5Ikol4z9mRSUaNXi93vPf+T4YUjW1A7rLfUB
tJyxtvyCUgtfwWNkYubkvo/ZH+8h0iwa2kTQGKjJ9I2wMHsw2uWFQ+sA22E2qu4Z
p/7tmkucNtLdHs6HzDj/t+296bq4n8hzONgutQD+FnlZZBNG8Kyq/EBWgYo15oxH
fxUizENDEnDqvMnaZG9fFbsgDngE3OnpckDk4OXr2PJvCctRepjTnfplBoTitpDB
eDV9bNECMBP5yOAS6K2Uy3tBKgb75IoZWLoWHTbCExLjcBp72fLZ03QJnIUsudpK
1QKPoH2HdCPbWPWL7QNwGSF13WrH6PX5swl+DETiwwoLIYQp67ESBnhVnc8kbu+U
9OK2Ogctq8tJLIgaPPTlgkCNUos81iWLKC3XU5XEdb7AyaD9BUJpM5mdAtqOVCNH
cg81+Low5K7ITSaUrcOPxIqH6GWE8kjUj58AMIyl1p5dC4q82NmFD78alfF+4q/K
pGpbJYHwrvk9YquVChhuAcwWIEMfSCeoV9vMmcs6TauqXhAMP3AwfnyqdW9h0da5
Ww3Ckt/8ZYxyMcAbeJE04kfmwi3A/x4MHnIZZ9uCGza5rS0gfcLlwavm9n6fK36v
l6aTGbrHClABxxX5AgglG2JEv3qX9TqyEENFKd8mqBgDFK9NMvtLuBNI1ElRXbLW
uPuquUHDI6umBsZsvAvKMNoNHyeIIbsMrxexHgoYoRXJfesE2wwJV1BtV3HG98lw
xiKHnNT60TUxicI/EsqJf+vdX8Nd7CC+xYw6IsTDbHbtXoLSH5iqY469qpB02bhE
ToIYsyaeCkYxbH/WAjeZYq4dHopcHCZDnRyoiOgkuDrHF7KCk2h/of9lDaRjqoTN
QZAvSuIUFUvk/Fg5AV1B5d8E642R+RtxKFTBc9kJo+9GhY5a435oWaHZCEm4KokS
/9roCNLafAeriF4En8l8WaTYNhZjvWiGbEhgqAWRePPXfuRSRm72w/aO0SXysbz/
Yz9RAzmYvqwaNTstFkgJqax0giZX2Q3ugxtzp36QVcQVdteo6qkhdMtHmExycYLy
/9eKT4uyRlHqs4iohZV5v1ZdSwVKUKhG40bFqbNiawQ0ZLKjRMFUR2jd0H9V2IlE
HJcz/ZzD7EKH0Y6rR/LaczbT1+harxfPeOoORokEerzzAPPlkwDAH36NdVqRf+2Z
tUe9CWSOUiZOmTp9+X43dSh//FYn6habKk2h52m+TfgbqSRNRunzxKsJse26VqnT
IyKFZjLgo5FgYB0HBgNRt26UJSTp9Jm5jda4/cJWvmsEp1Gu4uwfstsdR7T6nH1h
CflPYVib7xzbN98/RJDRHj9w4mloiNeStQAXg1o2eanimHlwQmwPRt1XxuOG5lNJ
blLSeako5NGTWIUSkCT4RWj3fdSQtCmHUi6YqbqLB3ljCqtEwmZ4YkGtWTYtwUTm
MO2naqbalFB0GNFNdjOPr/cuPNLuZad1raqt4YbhILLk6dY0ribwg6qqdCg1JqVF
PaD4nkZzFcNNZplJqlruQPZ+YlE6knKUdL6HSPY/1mfkGWrRu916cmroB38gHnEQ
YZgamFrf39RwheTt1nsBXI5Pa3NyZCM8Q4MXLFhHNqsiiBTTLCLaMbAlIVv4/+2n
rQmV8bnlTgkaIAcC5qS6Fkzy7CH8p1vklMu0/pyOpIevDZ/OxOPJLLov8JZ8nA5L
AA9wD2XjMr0QLpCNW0N4FsEuf/So/dYVf5hgXEPYTosCmtOZw52fOVu9QfjuhTA+
wGVyk/f/6sb3WYC4ztGqPmB6dlBpJUygUMHO1JnXIkjyS7OiM5EQB3KLxAveEPun
k2ASDtUSyVraeg7TDw2GcACJXnOYkI9yh8KPfnmOUM6meCrR9TQ8i00ur1VKkBjO
iu+ySmTPGGw/RFYw5+VjajWDnTIahF7nZhPf7O33ZWnazaRKu4gZaJOegbMBG3im
+XVBpiPl356vpMsc4YLd6REqA1A+i5q9/c1WTzzQrh2TZEazhxCwTTJ6wxnZTrwG
XzjC1shyEcgYFK99oTiDPdIfV5vW/2yjNnx5hy1HC2MoNwGYl7vyQX2mGtAqdiRz
40boqQ7HcsB9szIVy+oVmoLGf2IdpWZ/+MQubaAl5uBFK5mhTrpyVtKl28gAGzPX
u04Eevpqr2wLGCDmUVfUkbGKrFKn4ouvrwupHuK4ALDmqRcYs3/ijTw2p54kQazN
TObLcdqIqmTrFLmtv3Se83/roNIlCLe4ePi6UGRpbEOClVdR9ngtRa9tiZZC4kcy
pZcNYuFQoSu69fyYFIaCwCOKZFjOEmIVfTm4Wd9EyW54efSrV4GEMLCUbVdfo8U1
N5haqsHX0+l2dJ8bviV2foJKte/UYHWsBIKvvFS2AUki/k22H6PSCJshww45IVf3
8NBUk/bN2+L+oW2TstLl6arY2xae7mTnDu6pCdDYu4K9HgAiBKTKENyTiDdHdzGO
VQBQrjWlZesav5uCwhKVEXOGtyfHI6kbT1b3z4Nlif13fUdzorg7bvMPdIy1IPSO
MQLr6rndbJyacx0shNrkevU6+RDgsZt6inCTbiW23AQ+yM1WCq+sF5dX0PjIkppZ
FTU/Rld7iI9OuvuwInvbPGAemoTWtM0E0RBJCVxButM2IOzh8EM7XM3jxJAXl4K+
GdFMHg8JIwq4E8kF8kzVz81mDeB7KuFAjuunPOU1e/M3qk7Azp5WAsY+f7K/EdWS
n1qOPhSD9pmSXP5UC580wB8iQmnOTXIQM876jtNjcBRzA5L8oLM2xcr/Zlw8rLKh
6VpBr+l45y/SgRDiy11HpHArXGaWXc389vtZ+RFjgDNd14Skd5G6BQKS9rdAv/j3
MYuE7pbNDVsab7T27jK2JKgbAn2ZmzL7H4b+YqynVo74aL74ywRSL4NRnuu6LZTD
6Cs3rJXyYeE/18VKM6Qw8cdwL9xC8w18Rb3IOfki4cw6Gnf2/TgBs9OtytX9RACi
3hzUoqGaslqxAJWg6Y8hQzKBIoR/mCFJ9T3mJ+Skoz+OBImnLf3GP7Z3hHqQW2el
X2LNIEudWPVKFoXEBMfjYZhZy7y4mWUakUGj77XGRtd0hWoqGG+qLq+2qV3K8zOi
gXtVVFJz+MYcUPL5C46toocD8wXW9IgGMKTdtocJlqkB7ZSss64jRSUlYvwN8YT2
FapPsK/uqZW9lzzntHdogJJ7LvpQhGkTvU9lDReOjaMvmAQ7otOEp0rkgVgzalrt
B4mTFBGwME2LGspYFfkHDdA8gwVBXiWSRHmpGk4BUUx90uLWmf7eCiAyxtGlG95F
MwAvc1W3Er83Tyxjfd5Mvza/goJSWx7Yif3GtP48ntYtYMh5JHWyL1oe6rk/9gEH
57Nx9BR1yfTR/4FDPIXl38qzi17DH9uZ1rlEQxfrW0bym3/qSLmivTogH97Cit3h
SeUdM2uNRP+3kWPZzahA9ZLp4Wn97WioUCYOwEXALFWQU48NxHbfx6Bnop079Pyw
jEZq4cpcSptc1Q0K388IKYmqHAsdLcdVQZsN4YY7QVDA9pvqtZVhSNGonfomC27I
GWDv1UJOIkwMEmeRm5MlkWQsbY9lNzVKOjLiU1eTag/p1vcQN84J01YBLeZcJIDy
AX7zDwJfpd88eO6f8QRuXjqNMvUm3pjJdWS8LK6fXIapr2Lc2pJexVs+oflibVo1
Ji2x0MDEzLRQS6eytJqOI1Nqn6WbTM/rtA8FRHOuGQdVCPAswRMa5+1MhOpq952B
jw8j16SQcL0oRU4VQq6qeKdib6qWOpagpIgbHW0VF3udXqAfGHZK5xGtQtM3ZuEq
ny9Mr+FWvTUrOHVUHHKUR9uPzbXsPV8fCXQQnrM8Zh5ceM4yvfCzf2FOVH57qNjg
cSLu+luDbEBOezrHEAHl211phtsZW3+/4ULjEaOcbZtXNnZ3O2stCN5hAA7c9wGP
iMr3ItMHG/ONvlQaG+UqgOoNSnMeyiNjUIzgxhQkMQfacNYD1mwocMOPkzvnSR7a
mABkQ0Pd7YzXdh7o6wj9ay510kv+LFCvjsjKkyBu+Hkrm6JmGOpXKaLr/dN3kfIo
CybEa2aw8u8xhg9zvIPgdNIZSE/9lOUQz6JryJ4J3yFLMO0bDz0fu7x0TuZ8hNpD
dTg6W81grtxuxMFASvgeCjQbTeiyURkdWZF9Uq0oqGyG+XPrFUU30u+BpW3iRBjh
2BiCHF5dIa3V+XWj1xqZwPHHqAGjS04yI3obdLuavcXuRsDrjGnPTaVsZr2RGD8O
2iL10NX+b2LhqV+JWCkR5kaR2YgvhaqqE568BZFObtNg6yR+l1XlKdUkcQ/cGXhg
k6U1NsHi3MSQAV2+nKfZwh3pvyiedGYucinmNC8aKl5baUWMy+NrnPxAjH83CcQk
YrOm3+CDi7uR2sOa3yXGeTQZenyX7TM8kYzdqJsLmkn+DLP9UWQh+81/uyuxL7L6
YccStAauddRq4BX3vKoeG11UYIMS7feu80kwlwbPBgHSYZglfzDmk8l4IxwhvTz5
eqTckvyZSnPyAl9SGcl3mJ9vLeZdoslas8/4P4kBcRdL8rOQOa3aNxS5TN1XtNH6
qSVt0Gpt5E9Nbsi2SlUX/8PnT6ucYdPceD1mkeW3QmMLkSOHE5hE24Bn2W5O2H+k
+qx3DFG2GTkCMIN9IZZakkFHsuJVRbqfQUq4/xgH6ZxDDdAA0CoRnB+Aiic3dL6o
eKf/G1XdOkbyjrikQIfUw1+LBXVac0SOBwf6lzHxNILx0VLKKWhHmzCFJXZICDzv
q12oLP0eCS0ACigoqWogsu6zahLUEExxRvpXHXEmSA7vxKeIBLkLvNYG47/qb6T4
fcJtgK56pnrNsKBT62lhKuKNHnZLMQY7Sq8b3GSzvIMtXcPpCng3GBSLF61w7Pul
WVUjdcOxnD3fiDP/amDiurUQEsZ8cZupBDMYSBHwqhGSUAC/9FCT3iXoAx4HWQcy
g8Hnp5HkUYBAbCAbEIEs94MLBDr4fCeqwmQRSsE9KIBYSi2thI+3CqRXGYf5noh8
pA1dFGmT2fjeVHIn93Zkta8MqlmqpGThXaozHujSIde9gzu6chYdyxVKEhkXzEhO
Ym6vtxJNNWiA9YagJ6PcKuSrL1Zfv/y6Ug8xc//U3T9+hXsy7gWZC+S/hBIkupFX
UA4FAAT5IfyepZqj4dfzTJL9CrRyix/z3Q+Sb7VZmxVAIkjid3BlUYKAoB5RcS+p
rCVEXsjdoffvSXsCsrGnbQ0r/Cs7KA9yANW3SHLVN3GrZzP1CLGO4Wek3x2KYDcy
LUO2hChSmJTS6tw4MaVqbBPflR5yrCG7fIk7wYFFkCSbbjsr9rNohomb4s56StHJ
w14+yHIE+wLZCQwEgZEMAAVhjavebxZB4aMoZeVC5MqRTJ7sdRJ/l8NHuPVu5Y/s
EgEIOp0QzlMsZfu5mAxpWXbx1rif6+mltFF5tjU6rVxrGTGpsTsmk2PuRbordDPl
0KwClot6utlsGNATckDv85m6UIkSkpd+RWJsbjaE97cQdv0uyxfoKbNIzBS4QC29
Cm7pB5TcQZmi6xrJTyl+o90o4UTid03kVfJiS1H9BMBsMPg+Mrf0jhYy9qLZ7Knz
8o/fikV9k+Nt7Cyrxlaxr1f6tNgJ2qdkFok+2klbkgtcrG6h11ouhWCf8HvVdvoc
uo942wVakoSE8UmaPHuVDQ/0APY6hA+o1ymxAtgo2q4c6LJSekaCNSe1HoLVnXEh
dpuJ4mc/IpgVWOL3xZYHrVweNfKI47BJJNtyOCFGIIXG39NzYLeINZw4biB836IO
SWGsPuMvO7aUI8DAFVdQqlKjOUsKYH3sYhEw1E3s5Eb7QELqX55/IZNSbUw9XCP2
UWZ0lrq62ELZxi4RCCGSQVkcHYlqOFcv40jj+sRnvLMjqtDsbgY4j0zD2lgHVKM4
ujpEZM3Hd9xGT/zjomhWPPJDRKbBXz4HbUk0RXkLITIxcVW5EaG9s64+ssyNjv9k
5wimTJxvlrOY0DLAC+J6VRAYNICpo5R21Nb9pk4Ortn+igR1pss6ztU2kDIfSoTd
kky895qEilChp52/pSxnqMtqo2+mZJGiPGOo3WPeUdnTE/ajBrb111ScdQ3Vr0CD
NlxfYAtECQNmCCFCdncbF4p8mXKpEnD+IwnCpd3JrDnEZcXtwgGYkq7O0UfL6Ra0
cLr8cnlucurTxIOQ2Go1OjXAl+Qw+UW/qDbRkR8cBpNVA9aW2cpY8d7zW9jwFWAy
ctlfkr7tVa0sjuM7GTd5YKBu3DrgfkzjWPZyBiXX36zUBe+WvQVMDD0FgiXb4aBK
YKpNaxMJDZb/Gi7MKBKrGf/VBVMHjYNWjIWayrGNEUR6c4ljfcvGw/3mLTKIZJTJ
REnsn+rLIwIWdQegi3sd982y0iVxtSpYwp9i0Sh+kjb+f9Rj1RJnRbjtbFkU3nIC
fi/3KEPdUhS7A4aStD/DY/ly+1dL/dGDCWVKhYHd2ks8Nk0JgBb6glTP5cEbGIOn
fnNDqW5/Ouxm0sqhzITCwhXAxSOV28Orw67r/uWbikKvB6YMZy1pOnipfq82VKf3
DkuDj28HG8MO6Y0uY8L+TxY0fLc5yyG0RmfehjYNwo+huZCkA8iVmUnUjqUs7GMY
ETT1Wi+HBB7LiJLhar5GgjilE2P/vw2va1N+JgUwg0h5pmIXTOKe6bsxICNaslTh
u2jvcDA0MYCO5Lg6CZC1m9dqLNde55/mFPFLoeh8F/SEetOG1TEK2bqoDd1JS2Ub
UFuVcJYZJkXrSTBqwsNfuj51w6Q1RdKoi/zzs5xWxEHuS3c6dS070qNccWV1W/Fc
grbqhZAy115x4E1S9fLEjrAb2uVn7Qv3i8jJhttWn/GutpwL4RG9dxA5oNO/YpOu
L1eYIJtOmh1FaTb/Rb6WhDV/qjzA0Q0pylVOkkZdOetRmL+Vp5Wjx/FeoNBxG3JY
TugkESnTA1tinZY/zoT3DeeyiDAlnQnsjlq6Z3/gdtY1OmnTXjYnrySlfhaCqBmw
0XCZeiHLj+9d4xIdPlJ6B/9ToWex4XsEGH5Oq7XFfvyqQZVgWoRNECzkKMGGWUoy
PlXGVIoDDDLYJHKd5FMHH2QZZfS2tC9x0tjKnjQqqvOpbQg0/KZeibc4NrGAGndB
elRMR+h8risA8p0/JVd6O0LmXWRy6Gr6XwQ73Vcy0BNEYLiwPcncrxeP5loEMl09
j9wLEX4TM4MF/6gyeZxN5nv6Bef+U5dDh+XLT7SmAS0Oqg2gjCaoNMWnF3GY+N1k
kaO9RSjMCDWpLE4eJbtx/u3OJQCS0sRigMIZt7Q5VEK/xq+pZR//rAuhAYtRfE64
dLzaCkQ80TX+zNWmWRja+nBj/vleO1SfUOu2pJyLew04eJ4+Awuotb72zvdaG2dg
v4neIlfYah1YeBurNxqnNFBTqh1+33/9SHXkiKw2PtoX0KUw79sQk/bqxNgIzHVX
XvcpjsrvQPYB2tJD6CyD1kj3nNYdov+m44XmbNY1GCJ94L89r6dBPrxmv39BaYSe
vfQaV9VQRXGeRwpQqZ3gUo5VOlYJR7FYpYiDb9juXyyxhj8lY9KsH2ngD9+o4gyS
zllQbLgLXF9dAecR2GPWzVHeJpYJoRKs3hGySZuU5SrShYmg9wmCcqmQGVmwE7hJ
aWNCs6qM3RZ1yKz+yz+f21VA62hEG9zmSdypNZ9ib+NsEBlunYviJyCeM6wTTafS
3pFpEvYWFvG4CBd6M5kfDRrC2Dt0TDwkSk0TuyiEHwvo6TuMpSLxsNKTke4Xdboe
6+cWI46OKuFhAGRau23iggtuSTzTL4Iy2LL6EOuBcoQvXnw4TE9s86NF5j/t6hfU
FCaMMCPpT8szDoM/1g6JjlMsGy53ePcBP2gAPdh6Ryug7Jj/kUBSQQ6PpmKwZIPP
TNiDeET/WVnHJ9NGs6zw6ThwDxr5xDtEvXKQ2Wane2WRrqaJ6AeFTSMyDBzAXVSY
Ca+ToSC8vMfhWI52R28DykTbgfdrPCiBdBE29jUFYQkE4vGEiaDtYqNonuFkzmZf
TnUl44vJLx57I9Xzv+ho4pZmr5U78bppCEI7DlpwdqNKXlxeEaX/fMOgIoHCXFlS
ihLE25tBpHFxK5GeW6AL/SXoh4WhhO1PtIzWFXdAQO5DZbRJrDIIXhpGDU4Ux5jT
RzG4RTm7zvz7UcpPnpQJvR4LE5IzYcQQnoeEHcAROcXg4VU8O8e25/rCSjwrxDhK
9vP/0FZRsYxy4C3Q5U3v9gvwS/fq0+7i5sdpyGovZlEdquCN8HsQpK1rGExirOYq
Rpnt+WVF59I4Fk+a5rhqhWTEciPXOHF3eyReddznZdA7+nI3KQ3J9awefqaq+pU4
RlD4s3WOkKYWKv6ywERsJHJlRglCmFl8azzHr463RKlfed2SK1IxQ0LVLT4YzaUj
l3sp1hgsDreJo8VmD+iV8jccyHZ9qpuzLgkGOyEhJ4BRU/ZQmLsajgCszNb2EMjH
Z0ydfNJ4NMUc4aNaUVnDkaaEU5uAoFhJE2vYMEY2jXvNmT38gCkRX3k1TmyDUbMc
Zy4TWads1h8dm3rAtrXsUUglTMWz9MAM+3R0lOKTxOjmbzPKKBRJ8WGtT1J9RUz5
qw0vIpX/pk/1E/vmiDpiIdpcTOO/TcQQ6Ih5bl/exSHITYjQ2hPZzy58/WDEKQZ0
wujkdXADi2/buUkX3bEtcVV7k+l8qPeCe+vAmPZvuzH7v2a8KnGhLTwuvf51jvIY
Lkh7u5KokZD7Z5sL95UF6vKqwpxYO0Wy4iN+RkDA+jkjCOO8O8xwOupRuMq/sY1j
odiFlM5mS6fsU+ak9uue7m6kbMZ3gLiV5AgHSbyRo9/DlxPoMSHgpARMyU0vx2MZ
T4kPEwuW4lmIc9+CF81Cv/N6jgIfT8ZSrIYpvA6rRIIj6G2H1jkJBWdSv4GoipHN
vxlkb9FBCVhgOxfwo+2+qyxoAjqhdjA1cgluwjvITPqreeoQ8Fjj4qpgjfgIAj7f
Msko3zikHNfZ2QvLWEehFrRqWn6LYIpcwiFeUwNfmQaN2a/6qaWlDpLG2gDO/u7q
fmbANkzfI4uBitNkHDVJ70iFgIgL1ZTR2K4gnQHA1BWK+PAdHxjbt6F4Bef71+66
xx1W5an3IKzU8TGhcpJFx8WwqADjik0RJGmE/8eY6hKmG0cqMEmgCZYCckqoqlXc
LrtljQzV9Cres0pt5cvi+WTmJDSGQDkn+N1OsxYu+jR9l+dFnbm44axIxE5Mi/e+
ee0v5RtEj5yPqqyji2YGJcanQXeJgS6pqQYYzNKNcvmQRBv9QMqjb6E9pb5GoVWk
Lx/XIGb+o6QR3JTmYv9/QuOfZL1zeg8k/4fxbq1J+X12UGxo2Tb3UDKKNV0cw1CJ
/WDrNGp45LG1c2b75AwxZkBGElp1bnSK+q0A5FU8lHchXuKnH9ANF/3pb847r7co
PdKuxzmkttOUzZB0lwvi1m6bcmmlAfaHnm4HVT+xbffCXnDdzioHBUIZlnYo2dk4
HgCP094twLQ61ghSdyoN7oYmMoobGwK3RolHfY0aPcgDjeF3Lmw0FBOCFPAkpGnZ
+viyVEYHvYUxAjmAV2V2MZlPUtyY9PJKMAYnTWiC1hSmeVdAtVoIspvNCsByKvUV
trLhqEhjuSJ3D+JLGSWAAPkK4olh3xTda335va6qYWaRto5WgpNJgfBBVEtRBtvJ
J982mG7jrnwj1CTANUDS2Ij5LBUGuil95H+Qq7SgowvUDsR0zV2HHNxJpTmYozjB
4Zwo/yQ9z/GkBik1EoP0TCf0RogfrXFfjsQ7J5LHzwLfQwJ9EAbNBPHX0fHi6KpJ
kvbiVLvAGzMj088KwH/E+MrW4cXh23GD64TU9VWqU7jG294oOkCcxd2shuhlWSIs
nWcbroaEMC0BTS/6fWYKU8Cm0lCzqDA+LPtjqD9WHYGhs7SCiyWuqSe/JxmsbW0B
Q60nnldT2a1XBz230PcIBiZOgQ+ldedJAJ8Qx2GyA/3KSGRbQKUXk77mnSFfMXqJ
atMammBS2zoxFw26SgX4HA8pWRZS6Zh/3PaiUfybPo/jIeFaStRfypQ5FyT40E67
OXnfL/AxRWJl3XUIz7nAbYNa1lhsX6rfkY1wnuP71q26eoGvYSIP14qADyJMzeMM
Uk4Grx49IzUdWscYhwKik0iyy6KHuxpEuOd0u4WEWCM9rNmwbeZn7f8uEm4WeS5W
8mWNwgua+6fusmKVuy5vE4M/hZeRVth8z5ZxiGjuvq8VepMqe+eoKgle5rgeFcDH
VhUrBv2mETj3gROUQYzquy47lp3jS5pT5en2CSm/8PNll6HxS6vO3mg37D1FtRjy
FkootUkbDwD1dLgQPZEvOUrLnAr1E3MUzTJEnPK2pJDiuSuQKo2/yzSasz1jR64Y
8wdSZ3INL0b+GJ6riEXDasxlQpRgccpyWFud7fLya8eTtM8Zepbm11Cx91fG7Oni
AdEF4ml80X0QJ68+wu4vlzsKvFMiLtP+52GYd9VEex6V3atrPgWe9ODCgIUYusuo
PnDPoHd2u96m7icILiiAHLAeK6vWvIgIWwGcefYwx4j4fi6X3TmJsf0cahl98egg
p9exJZZ5pxhJBJ6EmogPHl2EvDfr4qSxfg1npKHT6/3zG+Wa93pZKG+kb/S1bDd+
wfXOFrhugWefksiC9238/BMS22lPfuTWFdEpkpSWCq9Esv0J/jEtI9UujgWqOoP/
Aqea0Q6PdD9R7j4z1WeKk5zH6fnf0kBnbpqnixZvyDCCaqSYyRQWKQEXT2FDJqld
0FKGcLxXoFBwm/15dvG1c892uaLoFICbZmtRBGDH+m2o1PHE8EMH43/dwN2BFTEb
JTJzqGTBF3kHTQxEuztV9KpjE7LOsnuO8GTdBdFkhqN6VuewvXX4CQ3Pw4xYqhb3
xXVnzcw3W+CfQEKjXKU8XYuG2DCAJyA18JHIA6dmcQTr1RrbugJRvaw90hMviINg
NEmKcdk/E26lD3zgtnz+WvhOQip+nzdBA0Th/u1NCsswDSZjmYoZcCB7FX6qE9cl
aex9DCK4mB972FQO9wHtdYzOz9KVtYfDksZNSzW04mqTBLccUQmuQ2SeeKxt6vPd
ymd8dktlbZP8YpI6HWNBc7J5mJEFgiIykiXjhGtJkp3kC38YbT+54ZBIXdvzc4ok
vpyB4cPGxRoDYBjQnHcriOEZ6XFY4NpOZx8REXGV6Xa/vDRtKHDihKHW/ur6NiG6
KY1Wzc5viO6DxsBJ9IqXoAna+420EpAC3KQ5XeQ1vQaFNLHjfPTEpfYQf/gy9ymJ
I18LRNgm+RgnJV06BhSGiNWM2am2SR3jmg5ieeT+Fng+ST5OhGHqUyhXbe13W9q+
RrutJuMrLnqpsQpeOtjMFKlJSMAdhdbXtyB6KVNDWkAua5xcQRKyzG1WglEFMZ3p
T0CtTZfYfc+1z2UG8RpPPQZlrpCN3eBSAYQ3FWVXrpCeRJW2B0O6PMwwrdz37SXP
olS5hdHi1ut8OGfm2bakrGGb6iegXaPPV7cA6VMw+ChoR7pY4Z2eWxoNNenrZeOf
2Bwrw5UVFsYj0a0LTWdW2JCJxGG6lgvAThFTWnLE5Gp8Tn1xS572IxWZXslLPdt5
uw7a6DYLs8kR27zfHaV+YUM9wzZWScMs7LJGlpecjTyVE1CxnyVEQFPBC4dVHnGU
TxXHp/20Uwxj/sewfc5EFM/YmbpUzLKb2nufTwu7PeUYGn1KjflX07PaFVL1ZUZl
tlEmSYVjvl4Vv2IPrpDZzXza/l8Twjtxr3/gVzq2Cbq3Dzbwm9k1FSIJBA3071uy
XzJN59BmEATFh0NIJElRnWqAxgeGjCmVoBDxuyt9ePxVrwJQBRmzdGbz3E37i+O+
v6Z//LhlHszJZG/ES9ylRejTjqLVVmaOTL5BFlyDpVmDV7jYM+Mcuokju4hRBKTh
iNjzuDP4bsCddJ7dO7hs0+kG3fQhPTLJlEEuWsi7Ym91LZyi+q0nXlncAd7gB0Lw
UksGDO8K0hOqqUw/60qFzSP0+jzfdAPmFwujKaeEyWcbojWZH/iVIgOc3uV12fCD
Ug9xBxcXIJurIPns2WQjYtkIw2+i94yEnSZOT0LYtml4nehrm+g/RCts0G4pZbW7
h5cbm+tnRZ97956cRKZz4CfRg+FmkLFiKZeW0JSSaD+m3HSWxA4KHApFqbRJvV9l
Bpd5AAVI0Vfm8wLQBKRCLXlHhN7uj8O1g227oils1JDbxjk6RDIh/BoKkbDuNs8D
k+JUvdRDVL3I9fSSHiTS1QSkqUiYj475HKwyPhW6fIZXIxifVkqIblLhufwmwfEZ
VCGQTswDIiOmyJc49HmDdaUWpWRbUWHDJ8FQEBQkRQGXu6vaCLI5BJ+X/ARSpyry
WjbXyMThZZYE/ZRynQ98D6ZH+kwjeSZPfziGAxs63ZjfetO96AilqY638nvRabcH
7SuuLBWpzEb7q3gix7n6b7JsnaB8oHgrTTHNSKtdLiFEv6JMwRYLeS0jCbx+688o
JMnaZV5mPaSbYCiYO1uYV6CQ7is9krMBteJpN5yQMg0qw8NUzq9l8GcDjoTJjX29
bdojVJrvdlStPNnAb+kTzNEdudNEAXqbony7FDklt4+XdreiU98UDwbVQZuQmOeE
q70Jp3ASIaHOSclbZe8n+XnTLBsIl6la4RWzbIOSOvWuTeVsxiFk+KsVit5jdGkN
ppR3M0ksrzz4M/BDh9+zouS7NBqeDO+G3ip0QJL4skpFbAMQxsyQenzkwyK3pkTx
1naPl404b6EUTsPkUWTRY0hkwXUzDSDP8+7nsbxm9gkWQL1Ck0tIUpLIbzHSjh8a
imLR08jUpxJu9s510QICRVUaDvo2upVEIflD6CqJz3XpSBmpoSYnV/Yv7lN7/8rl
yO5dT3i8HLRkYvPqnmswLWkO8999YC/QdCcbhOQvWjNAXjGvFH04L2XIUbndhza4
VQclS8rxYGkD054p6h+mfAdN/6YOyF/y3lDaSzsFyVp/OQzenegRJLOkRnOmCjns
z3QXTl8xPeKWTGWPIqtu9zO+VnIqkq/BeHTW6L18uC7K17BYcjTZi58fZ9Q65qMu
XSktiyUN1qf3HRXm2MDlr8E85j1nmGP/xICUANNjJ0J9e6di4X8BG07HSvINcy1V
MB/drjGsdHzCoCyC7RdgHpR9HVktosu6j6KnQl72hVq2YG9FMnxhXfazd8r4ZpkQ
09McWr7oQfjDLnHBqCp2Mnv0UNw3VwjXpeqmSoJguFIAx5BAIGHWVm3EcE7TI32u
kJtNR2dOJb5W4xwHP5puAIu5Znb+R2lFF9R/Rz1PEj7fkj96Gpilj0l446nH07pg
kqFzoKMpCDe4KIlGRG26MVoVKSqXQ7poX6EtwRjYQ9yqe5b5MS2Ii8Ompslil1FD
Jr/aj/4MLPirILXva6NffuxN3UiD878WPOyM5M5PKXXJ6yA3ch67FtceWMaNd6tB
Gz20ncs9D+pUpair2LNKDf4y+6iux5jodBBVTIrLXKo0h7HG3P53j81bKWGlvX7T
WbekNwjgMqE9nWHgrYs/PAzpVnjhQov6GkNQrMLvF2rbKNMXXQH3o22BWqfbk3HE
TPE9UqLZ42zYTDfuDKFZH2OYP1zNp/AgFVAXmInt07CzLM1ghLV/5OGA+yjDB10m
8iookOpICVlPqA2gdPwXzLRQ2UoQe19myBYqeGK9TRM9dDJ14VyI2yLKXuhJkFMW
Jk26on5D2WzhI/2q7M+jGi7fGe1+SgIuFT9UNTzYo5xjqF1f9qrmpyoEPOq1OEDw
H+mTILg/6TkQCFXLI42UYBcCNs++cs2iJEZSTlr9byeN1ZoNkF8+h0pN3w6BBUKi
xOUOcuXQ2GXMG7waaN7a8aadr5VAfHqaviIOnSkK6L7yYkpXyDvXoW3UVtD5uPMA
eSFC60MWu7HFSXornR0eieYCOPar4jsWsz/5Mmb/RQ9ZmBf60tVOLbrK4uYNQo3j
9d4oii4/2UU5+kz3msmiDUhxAWToGldTVZIigp6dn+OpUcWIuA4PasD1SPpYBdD2
7eHWSt1YIzpRLv8QbfrTQYQeszRDqAsiESkQtJ3wLNlPrqZAXeCy5H1Xgm2DMe9P
Xc/BWjhmUO18a+RLIthNCjA8XPrvwTEmxiKw+gygQfu/3BJSNa08brYrLrbgrRO7
kxTXXZy0QAcksTHUYp4x4NnO1g83fX/RMEo6ZUC+puttM1+xWd7KjOsx0lZXRMbz
t1R8+KC7mpTYY4VMp/l8YsZV5mkL+ZuLY4h2HpZg6g0Jnt4BQnnELr5UI2w9QD+/
V1+eNinbXFdk+HspyaqQofzOmya1blS9EhsKyFFApMy2a3ZGgQKcqHuPJ43nivZL
OOWj87aVZiL1xKiE6FSWFeTNwins7DOlNIQ8QeKxNn00zy+VexXK3JJ9Y7VoOpko
BuZgQ80H7lYiX73/MQbb8n09gQTKBUNdoQOjDujkyJDU+5qs+zj27OUeL/6TjLo0
Nz4PdKs4Dbedv5Dm9IkymfItH+kOqslmN4mIONLwHWDjqrwx200B1/yiLG9JudFG
Tgiv59P/Imja1yhqSooYcx4vSjjG1hk6S6IwEqu5PplhbpxwhpwvpBnRrImbAGf5
BiZyLnSTDE2QjlKc6ms3XM5Mim7hGrWLEx+6vD1cOT7+BRwrzhWC3ugqy4n9/RHC
JBxr5cXdZ5/R9lIcaWKVndl0T85tg+uWfReCdScpVdBjDbi5ja22uifarIML9vNw
U/WX93+Z1HBupnGpm/aUB71/20maBbYjWXMPd12m6+T1hpX+1h3ozPjJwwyAWzc7
S26ICP/1YJ1ur9HrfgZYCTvP6lWtVwi+qDACeivpPBFZIoWWcuYEImem0A6ICKf8
SUUE2l385MJj7BZh+YoSgnVgVfdxugbTBb4ueREFA5OlBmdVcDGOLLHARYPgljku
Rzlct6X2gNra1jGVsauIRrgabNab1PNXf7UN9LiYBGF816L7RjFo9ShiyHLYLeQi
3tuB6r2JVxFUSCCEwKW9gIyr1B5GEDAh/bdyG1lGDBrOMVVXqudQBa1P6u81WLs7
5L3+6LFp9EekqnDw1bGDzMu9j8bS1bjsLCPQmZgqQUGV+8T0W1EPqYLk7H+dDt/i
nG31oGtCMhLD53XobKnD4w+heDbOZGA21EcFReISfs7JALWEYayOpWQfit8yfwOx
wlFfgIjPB4s3bPBdYT5Chiuspw11SgBaP2cTnncGLWhtdgpc47k3lSJL9LdRPD6n
fuC7lVhougRn7E3SyYRWbtYGid6YEiTfcOMIMMPNFLqpRUUwTv0vXnFXZkg5He0x
A9o1VEG6JI4zwpZwtJmGhIMLMfSvnxNy9DNyUNjA1FQNu26fJYyWaETYATeDuYgd
xpcSv+x7Gj+rPJKGFE+224qr7+2Lrw7abusYakA48h6Xn1A0HuMkZuBaAiatibMQ
YaFeS4jH7E/tI/FdAoTW3b0ExISoiadAWAZGvBlP0m21dT//7YGCrj7C+4saYt2t
uxXZybEUA08WXNZP7BSQkykoSrC85n6TPne7DiBvnAiEUlOFGH5IRgwZZ6vaIvgn
uvtGm0/2e20OFEq7xJ0R4rDdCjiTBzH9QP8L922orbSBIU6t5Fpxulq0OL12oHMJ
iDXjBcrsleWCR+Zb2I/P01njNgDNbk786qFQzEKqYFtBAwjKOx+HMfqbypN/YUYo
4x6c+y4ncXcybGoPSv+qGXBl4rq+yKgpCJ7brGkqBCDC56DEanPZpFYhKLErjffE
ZcCriYTDJQuOtV19H+zvexLr41JRoNELBl0kC0mq36vZUoWYW8PeGqwYOAHzBwHV
de8T3H4KNfshufLHU2pWo1eOz8GU8Q2axLcKsJritWx35Uz41yqH0FNA6AlKa3vp
OzxlKwxgO8jgQVdLDKFqEXUCdEfC9/pw5eaDDkA9okavwPH+dnRerYoLzOLxu/fU
GnbPzO8sGoazDBC5sZ+AdSM7FIxiAAfwrd7I5BPOYzXbPX8fFNF2lxAyiI1kyIml
2V6bFU73FQNewoyrITvxKDzyQh3nhofWFVscExXt0chuLRGNZGlr+0293RDoZoiM
4ZjT3A8Br/HbEZoTpgcGMJAjV7r/sv1sMzFmW+3XxyYlcGlmRFVYwMiByfkF/aDi
t8hk/O1T6L91B+zDU7MxSxHrhITaGjvOF5W0ue/pV6YtkMWT/231VmRQBFon3PeR
sM5mxhfWbZ4NC/awK7hgn2GDIxN9o2O810JxXxk4cMzAXT+cy7KlIm8rOJVOAIA+
nC3mr0ngzBEPoJl0ZVlBcotCNpYvZjfqXZs4lKBOQ0SVd/vPKqTZD0hh3dBmPLse
lWeY6a9/YxV9PufakowRJR+24BLWM+lOrAtysCU8lOicZ6sVmDQIy5pW6854VDRd
ugST1pOAvXjeapJq+pif1FaO/QjZK8DeA+2uUQdgynwuXnjQ5a7+iDdHbEazavRD
+EFVY1vGpgIfMGIsmkbV8eOP3bxB5TMnIJRbandK+UuPYtQNsjzpS2quEqgjnK6W
JiM4thIus0P9bJ+xCsCu07HvbObvvQNfbnYRHh2OIJvSAwLmc1oNzhdqQu/iKsll
FqvuQG7Sdn6ojHPCb8ETi9qJFzZ6iQD9IgNdKsTQlKJiLsO+XP7q6uRAm0DI2qAa
Fr0LZFLeSNNSHcZah7sqpgXam3sqGMw3gUZkS2d+CLBAzT3aFDeSjgoiqkHVCyjD
4CQgTLqur53/pgxDYhmz2QYyNEVMHML59/ollXE+rJ8CTVqzHLxw0SDB4wyiPCBJ
tHhFtzr1D5E4I372kRR7Y1WcV/+brjFEEgN0/0YW66Vu+gKf6unDfOPrIj6bdb3U
B+wsviR/6O6z9+T6ziuKUM1d1XrtumUv8CLJySlpOfmJ5ZaFnJQN3iQgJbJrkbe0
TnixLRl5cSN6FTKVv8WXH3ooEs6V3SGpuv+9f8/e0GT9z8Z+uu2aQrGBiOG3kPCg
1r9IjoL4/SnpPQw720vETQEWbSjGt+rjm6EV3Z0wh9PiolFMabCDbw8m+tz4W8qN
k0Ehy3VJs6p9zDmCkta/pPiGEIouTZKSih0JbF46bP7FG0uzLh6iR0Vm/IfKUpuu
LS1Wj9CInGnzzg/8lw6ZMeSu8g11ee+zc06AHsUNw0pNLleKJyTS/NQ6k8OX+3xv
1aM9xErKzDhbaAZQsDfYK1rXRwcYceTEZqDE/A99XRLnu2z3j9guCLnlWvuxxlNb
j7ZlFKEROnlrktsF3xdOOTY2nQQJezsWuNH3U0iGd11Ull5CEs5YZDuDpcRno7Xh
lcjzf47kggagtmKQCmRLTaWxrG4IZek3xv1qUWYU/bXlkLjTEjtHH13LogfKk27U
O8ebV7TH5814QEItKumP7Khyr84HaRzcnWVws5pCqUilYkgiHFSa8mQvjA6aSznh
2gSjWSwiGuNmTGACj0AiEVgWw2JHH/JJvrI9MXunNAI25xv++ko2Uze4jxmPfch6
k5tbPTSCLjX0aZq3djw/BSzyK5gwXtlCMkNhPrRZT+w+RZNl4nleRssXbTlealWW
G9BE1zjAqD7U5lrksAs08Omu+KmcMGFLMi2ZvFYNQYn+21B5Lkr3w6dmSKzvc8FM
9rXFajzMgTl6ew38RU6bRlxpGXkURnOtbVSSExGwJf5VgtbhkWW5n3A4mYYygEVT
2VWyEPl2TWWgfkJo0dD2spaRKA4QrQd9Nfk0B1s7jwQuF4eriRJUmI08v802LA8r
+5bcR0v1fHBNLIVsGczL7JH1sjidhpg2q6tpM8yOCbLPb2bS9618XRwr3r32xNT5
dhfyG2v8KzLcBzcKIWM5nyLaBtiKBzvfeZNTlyojJdP28BE1dOdJMIFxOvukhS7b
pn2VqEv5HriemzePmfp39gKQijmInnb/rOC3RE8uTFFDjTPz9W96J8JBd3+RCWFm
FJuu8cC69X2mAiyQQYvQWHR1DSblcchnFPptFuJfLLDcwRthgAqEMxoT7x1KtmcE
7mt8XNiOtWzoHHfnqxqXmst1RE1ZW/01mo3kCzt7P5WAPfIPhJA0oAHPYt2sh+Vy
o75JNMBmwC+gKOsKadsZXJZCxG8Euv1N7fKdk611QainrESrNYId5dOLHXuwytRn
3Nx6umlm8VUemXvSe6zNgt6M2jpF6DFRa9FQhfgbsXgKkflKkX0+ohGdvyHYBPPg
1qP5p/rj5CV6UAlInKA/h0u6IQLMSU1FRpC1OiOv7YvV5lyvidA5MMjdHYOB59Ij
JhhwNimv/23A2gZM7jheTnZ//eEznLmN0+u7cVxb3n2KhhHVBZ0zlCRs4c9IpItx
I1j0q2MlJFZ56FrQNjfVreF8kRbburLtUa+ReUvW0vRDW1mB+gHF5tMrkoZTl80a
t2COoZY6LwRrsgAbdl+tOoRfp3OBRQeJsC944+gML+bYBmOQjVGv6AnNXEYOwS9m
PeG1LXxnO/zqTZiV+ap3+EFeZER40WI6ALAAS4/xghdnZGE1MSs8i4gbs5PSP1Ug
ssgn/Z3I3fKca/2CSG7ezYGO/cETkWRKdy/0UMYjSLro2VNZh+8h/fCaT6sdVa1G
ouYrMi35IYnYQHLKmIk7o0YTihhSa2q4YZFJnJRtWMISb+vHmF+Yfpxx35JomMWu
BRFNg1T/3lS4GZz4jffJi1qBA7XxWSrMODr3RDeWKM+ysDgxjaqr9dRbLK/W4hfK
7KD+0Zvw6R0yIKSkFGu1gZK0BVQmMZ6P0mF5pNkvVM150A21fxl4Enmllkmj27ST
g85Tn1RlDAU5rT128NuRfU4N7v+gVVUJvOXWYLlkgm+le35vzY3j9oVfSeLVY2/g
FijXT7iK0LwWFoBDhu8MMhkBtPiPmg3tfChAHhihMyZC2BEwcw60oX+zgpUOh5j9
OodS7P3lKa8PYozrm+XIEl5gcf+SiBpMDNvdhV+uXdUqOkpbGkq4YyhO3fbAHU04
VK0924zDAEvBYE0PjHcXMUMulp4Nvi1Vb7dGJm43Xtn10qW9MOnkinF0Vhe6hLTE
2zfnrubYP9w8bCqcMOUFyk/Ra/kwXOB0xNjti3vlBg5ozCNyMDPcdY6Om2m4uQDS
qbjwDbj0SuTxzBUSCiSrTG45OmmFhGvjwYEiP6B+wYEEbqbysUVcTsBWcVKtD5mY
kRuSVoZony3FkcSfnRPLpfem/PRtuVQUwp0SaEytyx2jCdUwxxZrhuKNKauqEe5Y
+Ry1linKRdqYWHDb+w8c19pkkUw1zsIWaaFeTvDF7aN5qpztmvJt7Bnx7q5FI1T7
RHI6jPWD3LKCJFy0pQJSneWNsEajc1GdOHcBFjWp9T3J7H3ZvSJcKe0NEx1Iz7gR
MEWe9Pok8UHonK+1GfQE9CNfItxYUHJxixgrMLtAsZCQ1H75Hs5KYlB7uCthmVuJ
qJZhnhUj6DbjyOVhPV79K49iGCDXA931MH/s8QBr0EgAcq98a9rhdGIObSEEHJIY
F3aqauwKNa3joggi7He1IJQdl1wofe6c+Hdu7VMrCQ0gVToLqEBaWYwBMav1GCAa
eKMbpAmS3WdBTmMslmWIJgTnYXdJ1m8duTi8zY467NEiV+y9Np7fV/JGmudx1uGw
HQ3qa43djDxkuw/8cKPMEXOPI4RHTNXS7EkElZXbjc1kwD5oFnTIk+4K7dsYtn1R
lXe9Pyl+NXRKQdlV7VkaXH1wquUaZmeIr++c1XtxCuBHUF2sL7ve/TtQrT/oY+1A
5ds+glXw9/okBYZYz+R5Lgia4TiWj4ygsjUKn7Upm/i/foIk8P7p19z6Kwwdlyi6
OU83UWbS01KpuqYHj8vm6JUS5A9KW8Y3f55QCu1e28CxHc+6eJB6It8KznvGiTBV
XAd8Xw4raDlEUCU27ZNggEX1BfSs5Q557RCeqfbySkV6ML4c0jk7ohQj9V/+XObK
2FQWlymC0exYOEHPIH5PsdGj8CY+55uEqAIP1iZ9KYPHcYjUQqSOe8Qvvoq0NNpk
3/gJfePSX9iZhqwXEHbjoYUa87ClfyaDteXwzf8SwJlCCU8Qspl5vFN7tOzgVN62
y5ZSRMUarbLc7mB1rHTCSGzKv0a7XKEgPf3nvn4BIvOmb+0ms8x6vEkBxhSpGPk6
5RZb3LIp5b8a8kbtv3RkGOJJpbRE8q+bgcWeCvGm0I9Hs0TXOa17mZid1HJdB4vp
WlFOTcsHeXJCo3JdEQmrgUNNtQ+l+4c4ofHbfU4/sJwjoFVJP5N7YFqiGqgfSgsx
NX3wytFxq1zcjgzP7hGAV772BOuWkxHq5nGhUWkN+79vUzDAjazERUqStpft2+ad
ye0DAC4el5JyuOZK6mCLkelOrmGAga8WhNRfOKx5z3OMQJQgxSsAlsR5doilr7in
V9BkuEJ60O86WqsBgt1d0VazHL9wQa6QYI2+vQXCT5TVLpCFds/GHCldD1PjiHMh
E4Ub0USxOBpWRV9I+tx8f2VjZUCHq4fWgtuahUD5YE7GOrhFOXtrv1TALclIVG3o
rqxLsRMe21A8SBJg4Vugv9RLzpk4OWSGLdBPMvSsy+v6its0csgP/fLZJfdQ40Xz
qAXbV8ftwUKRyShZI/EycRorS9YBFF+Ttg3WXlkLy7dFx4vAWjjP+Mdq0Xq4WsYW
2CC+ubPhNRqWbKK63Nph60pm9C0H203VSTcon8ZHeNQYpEl1Yit0vZG+c8v3sgOd
AZwHAR+hZkDb92PPUgCQCchofj6hBMbsZ35vSWbsFnw7EpkjbWROhqEPpWWXNTTr
rrWZ5R0VQd+9cl5/pCt3+8n2eb1rYJhpBwXZ+NT3wm9n0ifvK+JXZMVzj9O/loEi
Avv4wz8OSQdKOcwq0hNrH42VNTIUaqfoO6MFV6MIZR0FCAtBe05v/CvsFOSD2nJk
zduTTsRwkCJH0/AU0z0bDFo30A1iK6LJsYH6A2lQ4w55OOq+mqEIxH+5UAtJVcpj
V7m18swUn3gBHqeM2YYDBE9A7YU7IX+K+tJkG5Gw12s+SnLF0XyZqyMEg6ymJ5bA
/gcVVm04UNKzZE2a/ynxjID1supRsjwMNbS4StAnEwIl2hFxYaIgqRoVGFSble0/
o56Gv6gHWEo9cufLwo/wFTGb0wEROcX7fZIbUjJqMAA3Gv91r/Fh9XZr0+/sUCEU
NLbblmybvWUk1ylEPgETAsB3hSDWFHlrJgLg4lep7+NNOLdJnReGuiCi/BrngsiP
5oemr5vJIes4+90wWxxHXGSQefuPk+YjJSFWzSRCnJpfizNEdMSAr8rjwNS3Raoy
+AqjLJatifWQQVPjwP+0Hu6VBheAVOI8IxotJevBBqLWUZCVGZLflhR2VGyMQ/Bw
N+SwsNzKu7lwpC8/M//o/UoK8HjhP0xGDtsFX7utshvItBiaFdzaJpDNkuoSGlpx
yK/1H2Wn81NF5DwHMkpmMvx8SDEfGLGwA5xDXIWG3bVuOz+AB89UfptxGFPLfhyX
ytWy7a3yE6VRTDzt9c7Om1Ihcj0ca2T6jsZ9P8GR080P/ydY7VixrwRHyGABavz3
r3m67G+Z8gpn2PO/DzJDPm33T4jRFTnqoHqLqJtze05KZ5vN0dwVlj6m0T+At36k
bYIzQACCwvFExy6xS3B0+6450am5/SUAj17+jSmh6hLKSwildZQp3hx0WcAXolMi
F0ohppKiDaDtiv/rdIpjwGcbvVAapML3Hu1VScsdsFJKnhIfk23pbOVGluxBT/yO
C229p6VgvBiM0Zdz9bXUdt+Jf6j1+HzUvhdAdAsAd1h8dad1gNLkcVhHsuMLp/8C
5kSJm1nju9upgkoPoSc3SQt48/feEdzrSU+nWujM+8QEYp/uIUfQW33I/cKf+Rv6
KP49KAsz52bMCycCQC+gLO6d8vrGYUuOP/dYYfFGxFirxk9MNsPXn7RXQ/dyMadA
3o/iTCIRGR4rY/QX5I1OuqQuz+YqQY2yrnM5nWgMm+JyX69kha/1HhcoQayP/+Nt
XGNBLA6YGYj6uftDv5UWaNNgdXAEzYEFRguM7mKVyH1auvlToLx8JISNHkHUrQg7
F8skNxvrQJdK3CGFDKUjpvaatOVquEm/IRazIgCI0RuVFTteG9WRrWvJW0VQgYT0
I+cR92HbgRXHO37VmQTGZM/os+UXKIZZbIq8UR50bBvcWzcy9L8fWFdyIdXf0Dce
1Zc9PaGPcVVm9e+k72dt+BurYYLwjY4zA/+SemHBg8OMxFKpfRytjUPvongALl7D
SmJpfYoBzFEJoZGqQiZlkYh5m/deJJg6vpwQJ4V4BSin9MpaMuUN6S61vYc428/t
mVfYII6676do5a+Dd81YonBeySxTXDu0VsJmRUfoNwvicEIYp+NlnhpP1ev1aTAC
Lum/o9RPMTpbJrGXdhYl87faGHV3d7FGr7txlzPxFsLGy3VXdNdbWyPXIJIv/IfX
DR1Qt4Ffy1LLXmCuOYnG0sN/5U9KjdDItBXdRsLKCoHvVHPC7lCW+Dhx/WoDhz4V
sgdpRRhiRJCcSqaN/1cHa/rB/rXQLFx7TbPwa2mfE+MEG0/5JURbRgHV2WiII34Y
NS/1rVW7lflnbnuHTQbVgiu8+H6s942GO+JsZoGw+xpOw3EbaD4jJ2Z1XOU0AhG1
NVzJDh9+xCWxwcRhBXjVsbR+tHm1gKYfGl+snRrPJCh1gJb6O/ZR0KkWKQVer/mm
dFQavss8qM9l8X+LIDa/TBIetT7itoDxttcsoXyyJPUDNyK+kjn3PTtcja3v50c1
q0Ufa6JfawH7iGTeB+BqgNs9L8p6lerREqbMCz2RNNSly58E9kyRrhaHEG3nLQDa
gRPSmDzuh8/IQvNeWFDmzBwWuhxei3Bz8iPY4TRjZkqNwP267ii+/LemWBDpS9bb
yul2hQXLHLM+wAE3e2pcTPf1HH6rwoZelR3fovVkCma3UejKHwvpzu8nUwRb5WKK
zVpMCUTOBAAA2NjDCrwAzV6f9kUpaYctQtx1YL6tulQX25VrCG+dnlYlGmtE7QWi
LKKgj3ICLdXv/mJImEbUN/CeKCuIARl2uFwHQMNvQaGcSHBzJRHpouEDbqrH7akR
61xn78DRsPlJrNdAbC4MeUw7OXoRA2ZqaAvu90JIpa3/GTP04yZUcu3kGxskmUdf
cwjERlO+PoaGBijeAAEx3lSuHsa1IYBimdX9S4xLAr4YpceHmiVmSlMCAI8zayKW
7w9LF38IJrj8yfJonbRfqnbX47KKX/eMHqczFe/lGb20Bw4RzJ+R5RL1VNnd0vgg
TZuDfuz0FSb88T7D0kXaw7LH14VN0taSUoOPjYzKBoyFr9ERWNmRYo35xUVLZ7EP
uHnAblL8QD0XXWrrSMIFhKO3vn8QaA3+SfPFeYipxcq5Yriom6wg739ss4pmzVf0
Pnbhr+ZA8ebi2k20rehAVeIknRHHnDyezweyqkR/RjoCrVTxKZy3esWyFMRSJeVj
Ipdoh79Yqbv+FpoOk03PBKYqMkhqgZNZmYPTBC6GPGDqq/WZ+L3xqZ6F141URJBU
iLdbJUFyzE0JRS7tkl3p5UqZ0xtHg2w+/7e06iYp2uZh0wUonbFCVTI0EUwWx+up
oqqU9KJgu4Zg2r80uQMwKBj+u2bxY5a3FvNsxoqcaWZRvJdsc1cjiDRaoKMA5ts1
L7Ywk28VLBVWF3ZPXzgwHWkiWtsgMSmJAM396Ox47fKomhkrIYVh5PaqBIDLHFES
IX8/ZWkxdjz7oBOtVoJZrFYYvOKuQ93lZ9fa7xxzdGZnIlSVluSl0KYRrHCc9LKt
d/oL/SxlnDj3sKIJhPgqzsYtVMoBgrQe6Srrdux9Pa4D272mY2Vot9EewIKjwbWh
a3yZ+itFYIbr9h/owiTW7Qo+HCQXZjvWiZftuZvGOu+NtPu4D7CODoMlmNmkmI+2
z+i5wDsHt0uRkePKZP8xUTscEVOVDUNDh4toANfJ7NSOxw0g4sqnBeb7yaT4GE+b
f+pN5lv0btXU6yveDgjL007FD/bYOhjdPdx7ClqFMf8G3k2nmb/402pnF2hXNVdU
bjLvVwnGc11FOuv6gOXIVo3D2DKRjbJWd3lnovNL7bf5GxZIO3xDlfV7zo4Awy9O
7ujZOKp2fzfORcxxRbjtGMnv1sfowzACRgxZyPYcBEleeETRfWYz/YNNCGtk93mv
v/dS7+IM+A8ZUFt5vuZfseUBT2elElDBVUx+rt6d0XLsi7FktaDztK38SLxkINin
18cPH1QovjkiDs29ZabcwZhj1BjpO7pPUKnrm9yMc1GmMICbbmVirZGR1JKjqXFV
G4g1lnu7jA8OXSTCgdpfXMKoEsvDVOzuu1cNHmHT5WeRdWCQVVJrLjvGO7c+pVYm
nGG5hjnM75sTpio+cqZWx3+vuwxmdEGkJ2XV89Fv0/Wub4xgDFb3OkumbjJwUeiT
xIwpBpTGlYTBL2x6tEMJ5B6N4luQKPeRF1uCCB/WHexCjTExIeZlvvOkzgrt9DKN
vrJJGb7CFXMbmbQgax4bdg2tvlCTBZC9YHffz7CWbV3fW3YYGl4T9NSl0n+qTQ1G
ZJ9kK+8296X8JM/xIhn9yOcdLzGgsiSBferC/H60nqtX2aGVzPaNaUI9yjRPzgem
ppHB6c6a8+YRZXuhflP0MvfDTgwxglH7wkPURDg/9OYpmMdXcaXrNhUUaZfmxzUM
RlVGGmRoLTx6Sy/rnruee6t/UZQ8J3il9JT3jgT1hMdyyRacRjeG4/dKfv4/nrC4
Si0Lamqv4d5HOXDToFL4Kd/DmgvQf6udkpljsxzpOUw5Tl0m8Jv0exKNVGK5ptah
eTPm4xhMDVsqwmWeK+K4I+u7wm1aLPTeexwCqiSF7l4jLQN/0ha8ESHi8h0ETZoC
m0mM9aJlWKZyz0zt77L+2Arz5L5b+YYp+GWYvOa6nK86PA1KRFsmbAI5syAnggdZ
BN6FJFDw1zkl5j/YcJyMaxc72G4ZnyyXtgff2JWa/vI8JfkCr+tXyf6zHRFOvIxz
cHd/4OWFOJj/lhAxwpJyH7bDYTqhjs9qKOIrGMwkJWAwwCw4+2TYjM/vMu38rro3
S2gy3wovAVpysJI9F95zjVegSME11ARsEFtf3+yiP56MLyPApQ0RSm+s1mjl/RPT
Sfh+/mY1RVu9uRPOcByQgsX+3Y5gejDInHc7Ds/AwHe0dnXh525nmsgbxeKvgKd+
w+X2J1WawR8jH2u7TOWiUZcUKmEwPTBlwRA+jKn3t/pIsglp3zE7wOYva4jQM28b
X6jWM7cMh3/7v4NMhQjr+FP205ahnZc0NYxq3jmvvEkcwfBw0TF2zXXpDO3lczHQ
wvA35b12+93tPuYcxawqUFyk/yE/njKhV9C0dI5rQH7ev79FAszZmW0gfz79bN8f
xZLGM2fxEKnXMKAaoWA14qCdZZ/vgPuFwbxAQBoHBClF3mJbcGsiSruaYrWC214F
CfAMMcNCmFQQSO+6wa/ZDzAaEaEf8Zb7W0phhjkyu3qGvzVc0pv9CMztGsMwyJBl
LCoudV15D0BjNWFCv7XrhU1J7Bj8QA822/wUQ3W1z6Ahd+WFrD4JJcH5+Fwdi3nr
WvJVMDLIk3OEos/Ipr5Cq2+Myq+qeyfqKoU18x36m8ImS2RgJy+PE/g9ofomFn09
YO3Dgl8idAFhCrANa7IXUbGYCx6h4xyjji1dtLxwjKlfru4Cn68Godm5uSKCif+9
W15qly4YQPfnnmnTtAGc7lkNyK0R1107dy2CpysSI7LfgeOXqMt6kTTGnoedjas+
Dm2yMYAU1jhFb6g36Z5UMpyi5cBgieB1DPfy2LMELBTWkavQzzwl3kb88HAvO4dX
YrK7lKOwBbcKecQRmUrAf1wmuUpqoyluCPk4ByGpaQnbvSC97pLWG4fYXJnawFyS
WotwNRRTJvjmCCAkBFNiaZLircCUDHZBqGyIEA4fbx2/foi3fXmNdHi4HCOMHshv
diy3JkXLSmK9g8vND4AwskHbFKn91H+Pb1V7b5LQLRoom2icysEB0376Ab/rrcjC
1cXvtzfbvt8lpL/AkqEf/z3Hp0Ltjjs9GyygvlVM/Qz8q6qAre10/AX4nAKpVnyA
nrrSgpc8BcVwQI0WE39U0f2JdK2t8pyRVjQI3/A/TzSmibf3LSSgKrdd7JGSl2+r
H6kiw4ZtufxWFHLmor9DEEeCNPq5od+2q8LTUToxph3E/oHqJ2zMVlknAEx+tcaK
wudxUnv4AUnbltk+BZ8uUBBE1MwB2JMwokr57vTuszkSBRhmjbT07DHLmDMwPij0
o8Ib3nCSn40MwMjdia7YJDpsdCDmDMcGfhr16auHLD5RSR9Ia8r+HQ+mXX4qAs+s
vH8sHs3zx+6pbK/2jLMLxgs2k+IrRmKMeVhHJASfw9kW8igGWUWWSFw2UrtllDya
Dt4zj1NgwRTirSdcaD+6Qlrsrr4kCZzu06H+MFBChB69TE30pxamOVKoutlxBlX9
/l7XomS9O1QwDaSvbl2ohC8mkpgevQfFpHW03WOacsU6s6QccnGkf2zWjx5XzMIX
llz/26szYKIokCVlcitLAhdgEipjy8sbbMz6E2W6ZcolRCr0AGbPR/jNEU1xzTzl
qNsl6LKSs2LFWJrJw06a+Xdm0eIQWC3ZN6FICKVVSCAzkVEfPA9b1DIHJffAI+WJ
ScNbfuMIs6BZEEYAVtfL/LM2QZYTNwrUDhAR60wkPM+PpskDXFN/7x9Tmcr52FA2
5CakBYSLpSjA5FuLqp7c0nOFwpF0FLcyr7nwb8Qi+jJdbUjhUMUQJQOkDdHCKY5z
hWpMaIqluwqfzGjjdge/mRehZoOLoaVaQ4flm6m4CIslmmaPCAsIkxw7mHUtAJi8
a4j51FBmcRsUrTblvI2wi7LtABAgR+6GhA/4o+jxpteFhbKQjBjLI3k0T5iFr3ZV
zsTyHFRFEZNMmGf/95cDBYvhhZxxecIWemfFpp4dMhLyRTjqV5xj3OMA+mTny4L4
2CuKjG3tn4tG3oa7dBXk83U0WMLDF3c+of1Ou8taZZxbJpZtMPrKwQQUMfXLRP+U
DA6ySf9q+5BaycAOlHhR4MTehHJ53ZyMvO6ptXM6UtpH478OQxjwl1temvTGaBjw
WOQf25UrQFV7U7nVjDWDW7mrVhU0Ib/r/ivUXwXW3whsQSPxoC3qbPeeKPFCzsAd
HB7zsakVxJr8zPZg1Dc/7EVhDDQ12T0ueav8c7V+f2lYEP+lZDcIUs/rFeDJYm4z
DWxXrcDP9dORkEu2EUB21nUFbRo5dIweAK2H4HBiX5VeNtS+vT75VMYmiOfQKmfQ
wgeeOE6vVv6onLf6nOxGD9SOXfvi7uxBqNK5rj0AqYDvGLX7y32RdJPzJDISBzdB
Dx6AO+fey0+DY2gnm1kHyLd91V+jquVhAIsMIWWqK866t5TQrqK3knJ/nzTowtyN
FaONu2I/1wkAo5lU72pFpvIcWdEOkYzxdPJrtxumdB2eXNSdl+TKRmKLiS3rAWIY
exWEZxz1/7qL/Mxp7HW0cyf+An0mLCYnuQVYAFsErtLW2N0qY2eadvwQ1Un8hL14
4y3Re7dBx89kzsOdoZsnfQNJrPz90pnJNPzHAutP3kXdX791D7wUIy6IOLB5izJX
uTr8AnSRfJPjKheejcPjSRAhu0eL02DxjINtfT7AtdNsUkfbU5Bw+6lwGCiRNUaW
GcxvvDNEeZVhgac8G/3ZsMNJNTW65cpD2GSHODHhNfdd67B7sOgwQNtVpOnRp++M
eBnnncfIo+DzJ5L81RQAzThSyc63tvaWhD1AMGdhAoizT3M1U0uS93iSnPW6fYtI
1CXfdbTE9MfKLtijIq5sF5LC4kW0dxxl6o0G2Hre1yvil4Tq719VaK9iZ9s2yvzi
cL5mXWkjpI0Ermpbnce/vLIlETYKQDZ6Fo2K2wa9MYG056jhgIwKrt9avNAUVeQO
99u0E9QH1+Ge7a2R9beiIPdPYC20ZPLwBPimVlEofs6Runttn3xap414C3G/pegA
f78i++deGOnQ4nBPB3OpE9zgFYOj0H5EyDXUWBluB/mGhv0hf34+Vtw+NMHSQ8Oe
zm5tVQSjo5c8lphJ6RHNYjJ4NsI+kkR+flbZIoJZVJtKq/4oNoEarWA5C7QNZ0b/
nncOHC/4aJIW5RxH3YuVlgS4RrGJqXmLRvCX2BflD37/8WQXFwEdPocr7GRgCqyr
1BpHRg89GpJcDJRYSTE31K5N0pJ5uKKVN7rLm8cz6QdOGVCmXMIs9pKHDTcLMsqa
lGvl14YKGoFxGrc8zdt+D7n9heFSqcye7HFjpBXzuXr0vZ6U5kVdYDkzXBPgUlxA
ugUd742ibnh7pc/GFsnyZ/Q1oB68shv+G7TnFe1tUeXaMPZinOBs9k3NAW98djes
RlRSK8KteqJFiU5VDz6ehw6AmCJZBc3+SqdsPpPXsEAoTyoOPohPr6Zez+/PkCEA
8Hh9pSURFG3mU1X2Vbrp7R068IDjWr+CPOjbN69Nuz85KV6wvVRvMblp+1uvI90Q
jWcemM6hcY3HELGBPPOU8pvMZFREqMb3j6JMXeiDV/AGgI5fZFigdxwnbMc4q6fd
Lx3gNRxXyOhOLmWwnpi7L8p/OkP7tK4q3S4XZrGJCxfWUR9XichLm1FGmkRgjdU7
eEvfrHi+8RRzCw9up8vlgGsL8a4f0t+mfP2tyIVEPQG/2kyl7bajPVYsUgAPJswr
KR/7kcgKTG8Rs4eZnCo4A3E1Yq2mY5NFT/yxXWgcg22Z8cyJEp5C6/Twkp9L0jgE
yGtLmfeNF7tfmANQY0cJId3YDN2XXtspxWQLHzurqeZyPv47d1ZZdar5SQx1Tsvt
Ou65ZMC421mQjc+a4PyfKJdaxUl19b/7J/cbcVvgxcQ2WJgxKW56yB3oF2nDVn4Q
Per1o7TnlAaiX9QUT20gxjpWXaDfeyIBsUCkM8HvRPTndFtmoNZHVS4a1c2ezIIb
gfjsuL+ZFchVKgl/dzMMMGTfkuqSYoJeIol17lRpCCAOkHaxxx67lvf3GHdxot6y
P3kBxTcARd6XfT/XLQbs+CVlIS73EShTzyvTXSM+DemHFN3JA2bbY/dKiKSrpcN0
sR6jhT4aYi6AS+a7rxVPLX4S7WF1kKjCYfzdKt9KLxP5uYXm9JLdEQL5+YWN2qDc
XyLNEQYg+i4i6ELJ6hacSpTRmd0hXzI+11SwlTDXMra/IbCNH2g2mV/eujPbg+DJ
WfcCxv3uXLAh3dzWcjU5YTyTdzL4IJGWJVNsTj1CFXb8gffm7hKXKHi8W3SY+qac
uhJdzsLHSGoBufvxyY8PBL5UAVEWb88o8XlH6f931wPC8UOZ2oFso1BsarA1eDdp
mBn0XKKLej0BaOgti02YiQoxa/vxgF2H7ac37UMIGnHGBTDbnQXsDyUqttuQH0+n
K0FboQ0DDs2IRCt7+Q8n1+7HLvcPkp1mQj7VSNqfH+B2IFde0eTIGaTR3GW2Qnc8
9akpILGsTzxSfbdVrN+KMY1WfXYgrpWl/8aS+MdI2Zm7Rzu7lKw/NJTk0225xbhQ
BFNjlC43CfhKDKgSCR/1yhY4GXu/iVpc7SeMj8XLZ/aSaovm0gAF8ifr1jwwP89D
WpawunPURipdaQ3vkE0mhXWB6Ngg2r3/tJb1+0p3OFIh6in9dKGH2IEjHluVCgE1
0ctJTovLVbFiP8noxJBiwxm4O+gcwARC9AcDJGH0BtHnnxrqQbgqMLSSo8LKSwuF
RauN3GmH/5nzaMItQb5jUg+g3ACK/slT7iVtHjU0FBQI5Vj6s0eVDw61nfvco2j9
mvhmrBDDWtdjzEc4fX6UckYAybymditc4DHoMaKxoaelbtH/2dzh1qnnHMvVFNt0
oNcueatbJCxN+BvEGw/UMw5v0NtpkCAsXbEwQtji8MJu080G3DWQFz5pDhfe53l5
xTWGtvpxgaibR1otVPrh3ryP3M/DGB4HdwZAeF8s/WYmfcOsF+ViJJp1QIFj5d9L
jVFa0GWP0M3RE5AbJspqdmZ1Qe1GgOqVrblWBNq941JCNvU1C1wpgaYpQUn75/0t
5F2luPtYtYfucsWu0vsL5MfiX2+qb39tlMkGD6cT6p9QEffqXPOFaX8w2CmdKS0r
zsRwsp3PurQ+Tqpz8iZlMZzzeARm/BnyBMyHTqDew9RYNe6i7C47NTqZIQeijIG7
Z+YeOO5Ext/o+fnEFDreNtcqzYw4/PvxdYzuSXEVQ/3ZxSp30UOoFY8xOB8pq1sc
c8Wop/D9cMSNmJYldQXK0uRSno2O26w4QtopuBtnJB3yIJjekNjjyMxLaRWRiJg2
bCssfW7Tq+ey1T/GgL18sDC91OK/bixpnPthgIJR7WTG+M5QOuwBsbebhsnW86uw
srsLzB7RijmRv//3r3jTF4u8XYc2YoCDB6VkMWVxpx8J8nFyIHTqnLt8m6JQzod4
VodKnnQDDvQjJr/hJMMZ0BJblHIJh5HDNvvK7g1ijeBcBOrGD5Gq1uzCPIXbMUiH
bapqKXy242F9lYGuOE6S9KUO+99/op6i13b7EEkOSr2LQqME3WZlVdlejvAJOVZ8
id/W2sHfhLcsxK40ZB0AT9t2TRhhqDHO8Pd1Nmhs3ePouJipCORFH/hbPHgdIl/Z
kAdgI/70U55N/clbg2dUx09a3m8cdM7bVP8eq9Hv+A6JQib7IKH2QFtMVe52GCMh
dIoaHdKBYarw7N2nOxLDY9Lc+7zR2HemE2rXsUhx+Oya2bnilfGVUWqnziwLzYUA
2iI4UN0eLc3Ni8Hv1xBn9y+P8XxEH1OkiAgyHCIO/m5T1hM/qYTJfrG68dEkCyAS
GkFwNxUh6VkugWnA1GI7QvxGlFSqaiy6oe4F/sif0SoyA1mbdAw+wX1aKU+1cdam
X43CmA4HyEk+dm9Iz295xR6KRuUHa95A3OnG/6PcUuPinoorMRm3Y/wiQH6h5xNP
yxti5yLdz4Fgsa45AmlrTIay1AezoORnewM/Rff0cj5AaSrATucdX2+tpvXs50Iw
xkrogMW7Ub/vV4w23UbRkm8WTMRDwYGo+5f61lRlrPiWhry6pIlvCynheKN7xAa1
Q6OITRrlGEXKk8pXg2+rZogJDQI4FvaWX5+eaJe+F/2kmN6Hyf0SDPwKvDGkc9Cx
sBRSZtRa0sMaPuqpkyVEchMTddERd1FX/wZ7iHaYGwI6G+fX6YOZlYh2Zd9P8Hgq
kHAA1xtuebeyITqmw7se8m9RINJxWkBgPjqt180AP+V5JneXdl+ebMOJMB78tDDG
iI5rKjpfFW5wqb+wKeyoitG0wwyKu72IX6coAxUaVMUV+7OzRErpqlfN7wglDpEY
v7oG5n1I2tDNrdhs1Gzc4fQP8jT/9lO3X3rqc9ZrrGcU4bEPTxJQO8Ov3LaBTQSP
mIYFfIgJY5hnrEb5F8zgji/A20jIeBLhG/4ytW1v1PMnPnlc8aORvSK0r8Mu2tQK
8LVC+EoW3ZjTnVkfYH6LayMS9O+ogDjH3CZB++7sTZ4Y+pjYGMNCskt6UdkDr9Kp
fatAIBvRdjfbh74cQCxZApElG71YIJGsvCkY0vNAbsfgtPX3O/PQGZ3DlKSdJhQ+
nB53yLlMMqeRsXD+jiuhDNbftw4lbY85GFxXF23Z+9UwAbCW31ymhEdqAfBujZgJ
ZBznkSS0UcFrcngKHWZBDyuZ9rzswSHqyoBGY8Rd63OQBbFyu55edBCXEDSkRWzw
dgoKhBwphNEKj+GYxuDzyhPti8hUcepzu2JSBqRGAcOaWYOUfdOXZHUp5JajaZcg
Qo8CRufT2bHLfRSKMy/Xn23Q6fqBrPzY63JSt3T/Gl088ol9w+dCtXtgghc6ukD9
aXDt9jvgUpejh0x9Qt8IGvUGNDl1RrJ2fcPrfl+s6JfVsTpz3+uNp9o0q2GWNFDw
6OP4gRKzS7L6amAHgbIuc3BBU3dfwX9Hqg9sd7FsgrFrCpnYFftdPbZCd0tlZO8A
F7nvhfN3Y3iG3lTqJ3RKrUg4MUKRVNpORpp8rEqQk0ztYTQjJTPXfIb2yd5gUUCP
qSrXCR4tnOwHzjCShbTa+uS3teAckWaacR+fUBtg07Tubkv6RZre3ziTvZxO8Fj/
ntl6FLZtPK9KdF0eifNBcUwZqiLF5jVkWjqncY5KThtrHC1fFDtMwR3Tt7rUaQ07
RJpMZhR31G/Z5+/vDooBm+XpA+QbWF4hi0QEOn4/zp07M4ywTIm8JpvhgwzIRf80
15VaLqFn7qw7Lm6WRpoj+OkvE/QvpARi/cncXoGtgYUa/5A/G1pjdCty0i2q6qqY
UHeFktPbR45/AOjkNV5GyvFcKHbuzgxHG/x61CR3WbLdc9GqufaYG+6+Ir7l/I1V
5uMPVt71yzO2xBMe70jXY/lAebF/QHWWsq865Dm+snizYVE//6YyFbS9lQV52nlG
rewKT7atEH3dTDSGsNLeB5+dWhRAfuJUJq+z7aeCiPnhRIvSTLSEU6Ao6HbC9Kab
xk85AAvbhe0S36sE7aK6tY2J/9lURZiOtDqrKHZ8oOtA+WDcpZsWdkgT5mYOekm/
RIF2jMairq7lO9x8HHsxPSrFys/iqqNr1qh+cDDy3dCh0YSzO6x6Xu5hriNcTpm2
8GFhmJTo++fqZbR5cIp1SPlZs/m/OaoS7lQtIaIALUixGBj7v6p2opMOp0k68BJT
otkCky0YNta+z8Ks5burfDrKNt95lt5zIWoved8+gJmbX3JdWVATDxzmjkw6SsOu
q+OaQWnjGDXAp1xgUbljH3NFh5Zl5aq46jbeXw+l6/qGVy95XBsswJCPIZMvmnKh
2e9E2s6kjWTYw1pk4/2Bwk/OIg/DutaxrQfWuOJA11PCqyuqoxA4LAdXu3GsXMUz
tryOiOadCejes3A9pBTf1gS7cmGoXrqAHG5DMdU10loeRmZouFDf7KHaz14pmkyM
fHHRajTABc/CLm7KWkhcgx/Fy6XZijfgywEGMrj1vmqX7gjC8BvHqEWJhoPkMVfG
VyAu0QI7kqCmaT2D19EawGhcpXLTDQP3ZTqWJjPpTFE8EvTbGgGWrRjbXMmZVQQY
lZVzMX1nC4TjzdZGfOlb7BNYgMPiXgMAO3BYnPGjle2j/mcTEF79YymgPem3IZsW
KMFZAgZZT9law9nw9VmBACK7udEP3tQTDw5OknG4p+qlFanxzU+AJJzPAVif8Hm+
o0P4QNjk2vq+2hWMdm78paZowb++9HHcVUf5j8CDFHJeAk8wndSJ8JYNOHvkw01N
CuvXEa2hlUtaTiVBbr+46j+p1wSdVjEzf1MFWdXEP44SWKPYXYoejM+Ci9OYeoBC
Utb+6kXE5drqz+J5rw/q5AItv6zGbGYnr8uCRhrLuckFajewZAjMUX0doZrqeNP8
U5QOdsCouVe9pNyRfHuxVcL+5yhgJKRGHOGHBd6FO8snvSbz4PJMBIHpqJNx9wnv
/m2M2jCsfWKTMtGI9iligVAY9rJYS+VwPzuUo6NtrP5DqoqJ8m2mMmO7N3rhXDV2
FULsBp8mkcS74vUqF8r8jHbEUyDWTivUYdSHTXlenfHxAdnFe7hgeKOohopfL3+C
FwOhcvDDj6jmKZvjJf0py+6AyqXucS39YPvNpP37B1FLhN9xWjXhh8xluyEHRD0S
QHHb/PuRY2lBczTxWg4P3t//Fg23+1c4C0e4XQORfZtc+VdzDmE6b29wZ38ADatC
ARHIMeGMGhm1Ag9Otd2bO66CuDPd2HEXcTDPVbYvjO6C45rnxTO272QZOKCShazd
3babPGAIFwBCIh/EWHU8Qh+LZW/BXErWzVBzneuokYWthqwmwyP/pNIO/PgQqslx
8ciBtJw0eVRI3v0fvXDWWiI1qqZp6EX3dqAOq0arOKqTzEWC7VRDjNqq83dMba+q
WNChnhH1dRPATihfrXZE7Gj2liXFAhBG1Zw/GV34jdKuhrAPxaefyueWJtm4bLOp
fTo68vlY6aRvfJwwbpjaiopBaT+cBglTZs8qJYbYYbrdkHJ2LHF6K/UEAt5JBDCY
wtArz6C7dHkc3cLxSPbg0lT9ARienqrcxponuWdLkvLE5Ei+kTzxaSD8v4ulanEM
NVMVSLHn9UexJCPgvcPDSFpGqr+Oz/mX+4M/0PoGd+o1jc0/R2FBYA+nHYYiqBK7
lN2V1KCZ3CGj1zj1YDbqII+/NI9iGTs9KXk+EreK6jiEqF5HjCq3DYp1nv4bDqG2
F2BZAAfgoN6b9RhXbQvOvvyduzL7n3Zjc7nztBO59NaQ0qUG8Kb/Oi05i8EZcf3D
7VYMvXLnhi8cJJaR231FopjWBJCNIjsla/WI++qE5ZkUN3EztPvSoX42dVXUAH2Q
tVoZH3kZ9wDJkqahJtdoDyaPk09Q4hMOjlM+RLGnMc1Cez/OXll0gKmL1CH3I6IA
yfn8MvSDVTiwywgbRlL3GueWeeKqFjf20h2QC2k/PyTAgjQGf8YsAaX/TR1FzeVf
rQHWhvO5G03+4H+EcV6X37gCAWW7FVIaIZNbZXow3GfQDL9MFWWeZ6miKPc7PYZs
ZVNgd+XFX/e/ye2A7qaO2vzfcgVVtZyZ8j+9j9fFAUK9A2Og6jXTR5YdNstsw0zX
RGeBOwAQE4FVuNyCRMYQTq9a+Ymzitrdgd924eLfU7ZFZpewEhaiMhsq+TQcgq0X
XuPt0pa7IyNhaQpOQccx5/95ABYtcdGs1KyPRVHmd4qseFQUQdsmJC3bNzfWSlSL
q9JoxZjplzCCrZLbrvtxtX4knQjWSuhyF1ANMhLy0VYsCh4mgPO/UrCCEoy6QBM1
B46kmDSlkg4fUpJY/c62CQFTv65eAUYgv/cpbmTkDv8/3EcT0oPFNtQsOPVu8/io
bjsBC4sOHL1ekDrJ7faOJMDnAjeoCfrXZQo+RMs6qny4a1SokjVpyGcrfipfsaEB
CubnlMEnI9uboCWJslZhFrDGq3gGX45cnQ5me6yXoNI1lhLo6aPsjcXN6vzN5XxQ
xYmq5am7KJQSbHNcs+5iTh45tflc+vRg/Xhyl92CTnRFwQnNyKe3iRy5EXiXRsnv
tPGSeT3roobvqohqQNhql6NR8kj6MYPJk6OEgJuqquWe4GcqacR1Lo62d2sWYBuG
CUVkFUqRrLI2JyswrSGZuicR3pjjFBkIg0Ejb7ARR2J4FN8zPFVd7zgGN0XceKL5
Zhi8dmb3HktL4++AKQLNXoM/auGy/hE6NNrnrxtAL0/EdzrxRbN9tcxSLt0z2jf4
HepNj0NeTCs904Qh0BNUvrN4EchVo4Larns575uMlqn7Nd3ae/IdeTjiRIsQIy5l
n9U/ooG7Ym/fWPYCodFzzYqRaQAwgsvDeyjT+PljtnwmGh/jd/toOjKn+W+cDlYy
pZjaNII0U2vvz146QvvSNa3M2H+OGQuwy9UfOwjZ1ehH7RRSzYluo59iqfG/AGZn
IarjV5yLe0jgCP6x7duban8byJugJiEDH4c8V/tWks19w39fQsRpRVP/JyCPevbr
5qo494BUsrHhfKUgrA8sajS9FzBMRj+qRCXBETxeCODlugAKkVVnkVMwRNXPsFUz
HlnfzJHnUIAFWHjUHXlrnBKzf7b+IW9wJ219+OUTYhBDZGRCfqvZbYKGUWOq3WLN
5WJQ31qZaLX7AWu+KUQPkcJVoHkB5qGAVUNlGswphHjM6YzTvXp6fg0lu8LeqHEX
tSMKp/8USQ728UsV7oljiC6g5XiHGI1kLOJIUWiy8HHG8v5XBXbpu6vO8K/8Flaa
aS7JYS+W/hdmwHYFW8oFKlhNusw6X4Q/wmUCZslY1hXyXsBQnw7PZb4RyXBM2z8R
L5GwV6M1284FoqoJkMSzQkpdeUGXf0fJSo2/HmLm/moMDFWgek7lB+9H155VF9gD
LahDG7fNj0p4uQz3oa0PHibqWpBDT+JBmCKpRJFwoHb0pyEiMVbI9pqvfwf1wMmO
drMwdftmErZzOtSLrel0XHbDGgN5uB/pMQmN3F3LyzSbSqm+ULT4fW7po1mE2Zqn
uyseaUW1RGDIjwIwfcdnGWzqeRSPqSa5KmsuOL+KdFX0KQBA+Kx+8KstaNJ3NCUE
CWP9jOMtKB72aimHFvaFzrbRZTD+Xvw8FkodskKstEMKyMXAOS27nPnb2QhI0kzr
7C1xM83LJWCDDEU4yWsNpYh9eV15yUUhpncuOy1rHio+BqAdcfvavHNHujvyvD9H
PBkL8sp3D76/4nIm7/XWMe2IVTWyNu3XB0h5nGH7mZe53wBemHO4YYEMV99nf74k
IdLqtNpiqWQJXhCt/K6C++Tz9LS0Y6LmOfodKLpq51rNKp5QtiIEByFQmdeo/Obl
Pzq/fEm/TyFnJ+ZIhNgP76Oqssu/VYHv6ylHqaNah0QPRKPI9j7V6z4efq8WUD9R
ERow9fcia8vMiOrmv3UPHAlq1ugSegVL+S8OkaZqQDZF8XBZn+sKcfo4/p33XTlk
b9EMsg2j+kAJcO0sTc4zNPt4uq1zs1wU+cz+C6LkjnkGft2MALIbi+kmjcZNRYSV
IYo0tQgW7NklLenSpo0aPaID/yZBngEJNiXgvq/Y9QafSUo7fYERhQuNIYEswsvq
LbPVlkVU6u/4CVGC1+wm4ygxnOAWy7BbreunuIlvvEddhdnaPcyZ+CX89q6Dv1EU
Ki5wpXvwWN8fHcALMhX8TtkXgGQ+/728bUe7c8X9z3XUoKj4FXG+W8ESQzdhifs0
j0GhxV1rWgu3NWo7/wwX+lgUEem9bzf+m1TDFtTEQ+a1KLcFXGY9JrTTCT24Dfon
BSomXf0hyWGLiqn4R8rXfGW5dradvjUdGV+FZSkwZED43q9A65lh8WBWY6u8R9aJ
S0gqkPGofq76Gz7LYg6LKWNntsiPTGAePltI7xqNyM81ho+8ZRzHM/coLwpEiL8S
CI9pWFT0Fg0SJ2T1xWsC6Sr11DhNLlk3VUs32Pp3Ri/5sk9bpbL3IXdsgeCtLTfz
45DoLnRodNe/mkkl0ZJXhcnX48r4wHWlepcQei8mkPa8ymD2J4etkmqvanT7Ehn2
0qcwG0eECWyvKNC32fQYfzddy11goma3tYr2Ts4U1D18XRJaVAiziJwvwlAe35pS
7Hhk+5hC0ePeP6x6OYDp9GNkNPZe0LiBbfLkXiAyjDLs/+r07xunZzFBuMmvEIO4
8hQcscUxFJXBFhfb1CVdrTttdI5o2k9kbgB+AQgVXK269YzUO+VuR+JjGEhZKIb6
dlPpaTTxeko6FVqTgIf00XY6EzpZ3wZYPu2v7syvjVyHfZQhrXEfB5EWyh3oZ40O
oj03w86k5trkiF4ZCS8z6CFvPhfWiiwjj1J1edQzQCk/Ef0C2Tq4x8JO1+4cWQ5t
XBZ3o+iVdCD+uE9gUJ4QsnrZIbEdY3FvbpAu7o9AWHmQt9aSkbeBYOqaHK6Oh75g
oya04EQFGwVpWA46jZrytMYQEnwwSdT4p78OcpZZiO08//o9AKfv+U2Ej1b4aR/b
dNJkyHdMQjG9yJ2J7oOMCWbnRB4H8WHun5PIoI510dZio7ZGb5ZYOtDVFG9fdVUf
eh+6xmb+kZ5pbpZoHOULBFVrC228pjCVV7uGl56EvuBHRf9BrGf37QtSqzCUj1Gp
8ICrsIrjnvwhzBJ7B40eLoEvBfrMTN3BC67UonAdB4EgcL5OvXYAgUPdSiE1dGnS
PaLN2AU/9IA32l4DWzBFQ/IYWDkc2h/ouFLj0Kt7axuNEe8M6HTTJQH8Y+V8j5E3
ooQc/SCntX6V+Lff71s+bjyg/LPqSs/3jgNhRmFKVPKwNjOSPMiNHpFS8T9/l73I
DMbUxCVRtCL5iPUB8T7tXO1ju+hDt2CA1/RTwCUSB7PxZld4FO7O8J9x2CDPrwZI
VORrmc88QtXLQ8qneGOzxgZLURtpGCcI0EkGWP1a+5ciFTsShHCzf4zFXa7lFCmP
59t6T7gsx0olu6aYZh7drp7vk5yL1WyTe18ufe6APSgs2yP1GCSRNL6DLNFSFUMY
NqwVup4inrCJCAVvEyT7HeD2cS8ltvGMXh95aSpZKdR27W2igeiKxzbpgMz2lP+H
bKXrztfSSD3wrhbnxr24Hzui51W5bSMNeponh0IwnuWfrBN+t4oDYBEfa53FYSeA
37nJVxcHDetSLulI3OGBhj+1jgEo0ZqaD0grhfxLKoSA9g0Ur8USO93QDWwZFTRu
NRFyWcEpR7LLxPeb4Xv+c+z2TpXt5u7Cysp8c0CC0Ql++gNwyn3BiG/FZp2LtjOD
qxhyDpulTtii10Iu5WTaud59CWvzBhN/NzEx4EUzJyXk+LVtVZVfasJwTL0y+qJt
sC1kSnShh/x6YTiaKEQff12oU4bmULYQXqgoc6r8xOp3cA8bB+bhK6bYfBiWbKMI
CTIwsKxXA4+JRgFvTMUOEhxw7qJhfGWKsAlCIGYPN2pxtJ2fop0xvf6y30NU5vGT
kq2HVSLuIXbHUrWshFhdVFXytqRPFfBhtbq5Qu4xyZDBS4qyjMGHrdfDGe/GaUat
XP8TM7RghWh/362P21YcYlfAJAakwbFVNxJWUWD+jTyGR8KGHpOphqI+sg2Zru/d
7RrpwnMp8arNSeGUrJWKqDG8H7mdbThQJn0KQ85CdI2WX3aGrK5KrtFXgXZ3hTrA
vH18fwLwQlYg8mJUjMj4NTGFAskEqpDfoF40yhevjViVZ2IUdOhK7TuGsP4qyQXX
kRu+I8YsFH9E1pCfmmRZ2PNENjGpPWF399JMIfgfgv9rCTLzK2h+0CTGv83hZdHl
1JXzJci4Um1Z09GmZO9JEAUArp4ee4WpZj+aWohF/F+0uU7pqI/PPBGRvb4Jke4v
BlrfEETiqnUe5OFOWe76ErHMC17TyxJ4zLMihdbU5PzRlMgKutJKdfzxvC+fmRzs
rLiz08WW7453aq+vR0W28Tvm9cdqBDbAg6bgAJ5G6Ohd32QZDcjOzOMyrmA0N0Q+
sbVOwl0bnb67y/ecpk+zqq7GxCVqkIF94X31o/6H1Bt74Oz35FYfZk9B6xuDBsEO
GkTrmj20DYc9Y2kBTiP6UsHbJNA29k3ILXCkvldxogkkNUv/tJHvWFe1rUz+NwfB
cg+rZHKzwO/ZFUf4H6yy3vPrjmMABUFSqSo9g4wBCbDv7z/hEfC90jW/37ID0TNK
fzFKIH42qQPDv5WulQ17orjn5Fjd8+z9Mx1YQZFnMqVrZSKxqrYLK8r/2Ys1zzA+
07Z7cSKgsBWks9ofanHTvzw0jNtGaLNklLWm3h1OVF4freLEuHO52EsOxYyQ1+lJ
9CFLQfXmHfo8DS8dvzBVHUScg3p2RfW17QIEyT/Ia+NYGlw4o+EbM3j08oPno8bH
pCQTigIV3rDpWLjncqH06hNEAFERe34YRyGH61ofeQ3B3Yke8IrCKX2Kltnshme8
04PCJX0Dse0Lp0oGpcUio7g6rtHe7K8K/g69oWDNkpbBTRHZUvHp9yfqDMHgwOLC
xl5vvjMYZCb/Az5LWQbZFHRBPRtySf0yR5A4B5enYU6l7HHQqaKDPdpRFl60zteQ
hhoCUq5PhM8GJy4MOJE16ThKT8+mBuOUr/lCztYB253chlvd81XTAuVz5cdcsZEp
Gqp191relOzpPyOXxYjJCLkWl1BKAT1p6Ta8fwlmSGwl3hMx0xptJbSAS5n6TLVn
pYFHsM97kf6e7bR1SRKnXFpe1l0PKwtomh1rBdMgAoaF9JHg5TBi9N5B3+Gl4rD8
vrRJ/tyHAsc9AJaWv8I87zXRDxXHkpzerLw3fMPdd9rtSpmpZqu+vfiE1vloLzP9
BfEUGm+fsJgWpmg91YXBkFK7ECWoDZTJJr76jcTaqC2JGR7wpcmVVxrv0h/mVzbO
RT6eB4JDywnjNHg8IV9auwX3d6qVreLQ8Oosl83KWSS8fKnnW8zAWkzE2P9+R+uN
/bFnLPaUhe1de5SKVKtNYbQI/CcsR5C0gLut0MnJOc1IW98eSnlgVpiXznHp2m9U
WXulppLp/JJISuYBAVXJXF9r0CFAiHaCxE0LQfUWJfOc5TIliM5D1bNCxj4iJMIV
6naeNmk0NRD5YXLQynqCsX11Ul/NudbuOnQMhO/yzHfVcC7l1SMksBqwyTO0gyD1
RSilRQylYmpxT3ckNPvHU0Q4Fn5mHNrAUHvX2LWZSZk/vXJWDEbGtl+RZN46crqh
vARDBZt0qKOAncGThCQj43Z62EsYkDvhzT5373+KgUgFlQvXL2FwAClZuukmHPFX
YoJ41BrkuzBpPCvyB2doO/lVU+6vJBOOQCFCpH29iYM6heR+pHX4xppQOBcuQJGc
qLWtqSEBoPpAxS3NOWMbAAos9OwsruuEP1QzRcBLAx0s9JT9+BFLkIQ9JXBkq9rC
RwgZ9npjY8g4BUymj7oQMBrI7cDZ7/yxRtStQxM9Jta6+OabGpWCy6DOA4tzpXXe
jCttECond9t2amaFeM0cKBB0x9Xfe/uGPdMog35ByOd/Wi4QUhF2+bbsVNF0dvwH
iUr7hu/A3f6oli+x2FsvJW/BrK9EluEX4LFtQgroHdnD7U3gGiXZEmsK09SRCyJh
ruIw9VVcbVbzs2O4TcB7vJILZEWLELsa5u5W4ZcpJHZ0y/VMTyYe5pFgq9uQ5QnV
XH3Bmmq46QNRRCiJglUoFsrP4HxDRpwcIFzVMYJu8HIxSGI59qBVENGyE0GUQNb5
TU47s8DacI5H3Y3rMv49jCTrcWceqPAop+hzskzyXSZcsUE5QeZokdjD+TqgBC1x
xCrropfy0aBdoOLaks6zYsgIOC9jRJPObB2iYGoqeFcG3tai6376ittzVd93Vqll
XN1rJI397eYkGOSgVEMpCBbD7U2GeF4OTd0o0x09hLzAu5v7SSmtPSn2+iOU2ZoY
+XZMce9UmGdbXylOLNAhbvn37P7rrCFn4M4L6IP4bGylMgzxP98yGMHA+Q6WltmN
5i+lys6CGbeL/UVLl4vTs7Riia2A7ErZQ4FmxQ0H0Zt0ofT93FITkWP4Myijgf67
LzN1YshCgQ1w5ZcP9UOvgNgztLVh9TRfjo+dVk1+qT4g9IVst3GufLSsED9QqOxm
MxYmbw21i66tjoigEnG4Nect4QtT68XCmva+3Wcb+Ock5OH5lIU31gpa56C17iYA
5G8yRSHSvEiRWwRY18Q9f2xCW5GkqF6QnUQLc1cOFx1YqN/Aph7TK9oiYSMT4zTZ
7rXoREr3LuuikeC18GuKsQzzGcyzX3AhO265lt3roNJaPh5/d/vhcsXNgOACqbiH
FJuBsPI8Ef/Ft9p1AvgEtrYSnjgRGdVzh2ueUSDjqEh5aRTM+WQtRHGJPjoJebpj
XWE5ckuApR0vs3vpdowZHfyD9WC/ovs0qacbNN17Od2xv02BrUkHF5Dm37tQXh+f
M4rYD7n+spUXmpsVwhe+xgO1ShwURtbnI5ETPSku2wsLUWlmt9ZeLo2BEyeTizgl
iWe3ZuqNDa9Xuzyar115S18LOpXRMuHvQiUL9k+CHHsZmaXkZRh+J7dOiEZ/zRPN
+iKsIGGF2kfUSkc+ctR8YHdiURsHKfKCNVFsF26fwjnBoM7Hx/p0ypac0oLv3i2J
+/Efj42lQcr6286/isWivdxkZXATDmdtrBqbDcz67Wu0u1ddJZRAK5oDxF+mQ7oj
TJDhZZXp5xmfS3cYjiARiorIQGwdd1OmVgvXEkJPM/adb4SRnAPqhW5nNl3bKMOE
MY4SYZcuToYGRW7SUOo8gbyL+TlW32iYH77BGy2sk1ZjA39CYXDOttBJ87ApizRm
B3tJYWhY2A1cUKPz07DvW7aVOnZS1MGvmHqq3rfuTZSvpee/4WGvahT5RMkzqPMC
qOV5gEZZ4TY4BnNL1fj4+kF85QGRT04XxN70QTxqbjtoDKgzNIyxqMgJTWx5pO6b
Ppgs+6tXFKCPCqBkWWDq5szOWjbZN07TdIcqk8j+7Wi2a+n/BbqqSd3BHTstiWKe
wmz1opsNZmjc+xN8JJjtdK696iDC7wNk0ypInkaTJD4MmsJ9KsGoUq8wef9Q0blr
t6mKmVQvWPyIIODw3CqbcDNjKi2acq1NeZBAPWeGPeL3jJm4Ct/dxYvko9KJc/+3
JBI8rcrA/n9+FqO4hiLGD1TCwYH1o9u5WgPgRDIIZNjieSw9HYq+GTGAN0vP9aWF
iEvDqt/kfH3yESVLQF+43OYKuGB+Op4XPs2bcn5ygysGyWMBZsPIdkT2xOLCYj98
8WcZVjGN4riRlRvhYU+nccs62zLdANSJGn93OSiiu3iTLnzmmW3a7IbKFgTySXJk
vamVM386oQz4B1j1JZfhvpikHzMaUVsACghXgFRqza/H4yZgYT128/9mWwsOpoIn
z9mFTmiAFxarIcNTIZgnvNitgFovr1NOSPSqui9vZmkyJh1s6nm6ZDhHFEyKvPLq
LkVlNVtmI7gQuq7weCkpIBWI5kjpN+jRMFoh+LyzVlfypp5rdM6gRkG07UTYGEy8
SBPf/DcYB6BYwp8BOONOYwGQU4LkcJUsAvsUF3nP5B8IxBSXaMA9MpccvpUMyCdh
MsapddJAftF0pbeu64hvnpbIKbN3UWtaztTSsEXbh5mFClV5YJOkZSOdSkymO5Oo
vYh0+zh+qyQwMVQu6dhjSvPxe3nDu3Qc5q34ZUPWwKsEvs601rq3G+5HxisH7d4v
ocIp/KSYfD2+37WeVxb7RoJF460guZ5MhPCEgfK8iftkBD15kkbIGnaGTfH29xVV
JPhaKD8HjRx7TcVUz5NNnZRn8vLVjUUWufq0bMNmzD/zGVigNSgrf44q+XRpNQDE
Jr3iLZxkRw/5tLDQ4HemzvxMf9jmc57iptbguppm2y9tUQ6Ceszbp3mTOVa3eqjW
sz6Rk+B7LFIdDagnBM5Rnk2ZqVY7Wbk4qpZcmowQ01UtdUxdXl/osndMhlE2hiQs
1YDxWjJOffffKDSLZEMCMCNOEhZbeo/CDR5OkxIcGVisjLUWjS6AGOEhwDCMYsPG
cnMRlspOgwLhEPXPXQw9J1IlzwCpDK2c3ZZllC35Xmg1vwcdD67bjERClMLC1yBU
/0eu3SPOvn6tNH0ERjPyatCXNt6It/2ps5HjJGfk5RKumnoVhNCDPbJaO0lmrftv
sUvO1YI/wozFf8xwTsp6YAbpH2xnrrt9zz9x1yuzor2FTO+7XArmqhet671mect7
XLL22k8Ds/z2eJv/Jh2Euw+Z70d3mkAZVOusepvLy8un/qi35/8VvaX8pod5oKr4
4NSsEH6yvk4mvE4dbpmNYVov0ybB1djjRHcypxI5yL+EVYYcACfUaxcJmyzACVs3
Z/W9iOlm7H/ZJgI/TRBPn03qrMc16nXAV+9AY6FR4Xs3MYNTN509W1aMP/oegwYX
jDKDOLOWIeImUxz3bX9Zo0Om52JOFQZQWZlMdSt/EZBrGhT3LcS0euh1A6UE6Hi1
e7Mv7PTA2KbcyQLw35dNcxZJxKnckWZfclvOqu/9WV4NuV5wEv754EzOuEq3KhmC
RCMSi0USC984sGMHn1yqJ+jCkSUWJSJkhFV0aJF+0dMekaR33QIDa/eemNASq9z1
lEizUluIAVgweWMfM0KSOEFLYN2lt8lBfZGUufWvQDx3UphtEn5SAsQH91/ql2O4
OyaxmTWJCE350yz5TbI5WjoZnlX10TTbLCgHZ4zJsWEutS7eC1w/scChIl7EghYr
smABKBW/JyEGzzzv4WnOdvPG5AxWKGxs/G8/OL4CZEPCTAo4Q3k5T/DU5buTpMxs
0VR//3PQb6xKKtaSa+mQXZbGED9HBR4xy7FoRQP3gtpNje08WHL8jkoGRZT4CJXE
LW12cJaoG+weujABztN8H1pIvE1ujFT2br88as85vTGbLK7wj+NaQxsVdJ/v5UK2
i6SfzkZPPY3Mc1B+eFh3T3Uh9icJRE1O0WpFtGLuRDlBCi0lIK57EdA72i5EwoZy
0xMkDR5KgC3pk2ipsxaTu1h0ns2fKAHqhtM+vHPGkVqaPrfOfvtqj147nWoRt54Y
dLCI9wuTAvXHBIJa9679d5PiNQtA1XTM20p7QonLrQZjqulVUPAUL7iNs9qNi1Qs
plGdadmJAL+vChVm7TDC6X1K9I4POhrIPfebJycpT5975Wt4JiKah4BaYLShJgBg
x9+tiMe/DL0a7reMwgFIBkJUbeLmv2mPUrU5AwJyzy4WPgwIAlVC5Ohhicx3DEBc
SjLCwce+aCD1yCCxui1s0zs/HZBrOwkLb0yBEU5MpOzrvstNbklI0ckWcVR/GuWP
O0VHW45ldavssHMykLp0CFFfMfzma+jhAyoncvCL5fD7/GSXTo+7g3z88tcs3/CC
zWmukDgDhG7yZGIav6rASzr03jsfB8naf88/bkHD+ksyKxCTgwFgtRbCQXf48y0S
8TtrYrJ22gkzxflQBI1t3FjFIGuAvuOWpcrKWYcAjmrJxStwHCyhbvXqbngw/bht
pfK24B428MMg+T9weBrcDOCMt6vgUa/JxkvFaWc22Dxso/AibtZL4lH8md2mdXUg
BT8gPK7pRpvKu+bhbhy5uudOHDAAfKUrSFGCaqoonNuLhn1bVUA6pQQcao0srs0G
az0U9AtjXg0InmNTzniSZ0HUMpRIZIBncdmu/LYy++tpHmZPRa3UEmg2Y0Ikaclp
ScX/EWQSWTZusdnH/luJFd28aLZn8LLbo1fJs2ejvH2zb2gTW+E4dHOdiK60Id0f
xH57UlmGoCYuD6B7rol0zWFyZtuKXQCUnLsItR/NuNfnJAiKb5EkjkzyLiPJvBE4
7a0BaHiZaNy/626FVUmx5Cr9eQhdsKtRtH6pln76YoCGYcL5xnfRweM8PBtkhaq5
QYA8J2/6UKtrx2QOxzvSRsUQ8Eq1Fk2NZUKMFhAyTGfiGRhy09u4sChyerTS6YZR
9rybD5dgUYV3OqnsUfKmUCwk/2cjpWIbSdJAGPVdQpSH4T8tcrkbLmZ/3vhMnSHO
qmMLGBzhKgcg6CrpVWp2igiIuT9gnulxq1MQY5iYujvFjTnEilqTwPI+MpkA9xNF
Z3FRJgqwNvvI63/RmrfLsF6eBODRsvuPp286tP5awiLv8y0hHBbwHHo+4kHnsZgh
jj9j67IYN4ovFnImLOAGfBeilIaEb9xcYG054n2Qgu6ZlhX8NcQYOt7HGPmtDM0a
b9ybKOALVHK8cpwZ1X78pwdYsmeZD9ZELewiIwaGQqV9Wp9ZP7xeGmLFWA3wo+yW
hBk55FYneCUoMh09LUy0LnpcrZP6b35eAV/w5o8dUdIfvWnTCf96uoaaCcGkzu49
D7VD2IN1fSOuvsjyJQuFowj54knuk7UV0tTWkrLXZmGGZ90CcufrkF0PCn/QNQoC
MG2lQWOIYmK8jIWvG69HDpyqb/pnFQd8y/vvq9hcdIe+WcgJkYFslICQSY7UeKN5
lT6dZtbsPLR1YgIYNtv9yRTCnBh9AUhQedH3AuTCFeTaYdX9R/tyUNQu/nR0M/0A
6IDTdwVGdyWlH5FGER+3GSoU7IFKCk8EU7yhQuLpgV0aPQR4EutozaoPi1oR8gy/
80F2mb8Of0BTxNr0l4tVS0pLfqJCCH2hrd+R1aoWP1aQxjWD7j7GVFD6jT8nBMyp
Esb4syar8+hZCca8vJ8usmPc3ztUWoTEBJMis4SzY30GqmD/Nz+/ipQ7ag6uYJ3Z
Rq/+dxtbAMmA7K8J8aJzciqtDKadwkVNmMPWoIH1yizO+dvcVdZIGyKlpofkPmio
xUjNfDdV25B7oUtvgHDqDBAIb3P9xSqDzmngHqi1HucUTlvoBZjQl00LVKffFftK
mXw5+7XNMm2SgvmDAa1QLkkERt77+3qUZ5SrNOsqhB+Pu8kiHthINUFARf32RFS2
9IDTUn5/k1rRQSi49f43Gi2/SPkNCUyoDt/Q4bQjiu2dNHHKkIk9L4nZI02Xx/FA
46cWE+8YiDx5XX3WbfnaQwcxuqz+QEmIeA4/uSZwVJoX+LeM99fxXVSoZlA8JkiB
J29Zrb/8hiZfEahQ/7mLM5sDxFwkztyyJWj2s1SDxQpvUR9LMbq6oeTIVmCbkORu
ZAIgLl0qUJXveblXDVGzzPZuMaE/nsUfrJLDFCu12hkWpJjmKQ4D0KyA1lM4dU2d
drhsv8gToRnb8oEHfuBWuK6Hc73qK7yW7N+IACokfx26wK/kFMAScNb9GTXralr/
fnHj74FvTjRA18Y5UfF+7rZNKgBIMPXygKdpOJiCFuTg2aHbuTHYa/YJgQ8IYjKB
t4Mi0t/Xd5FWiHshA1XFhCRavsWI9aEFLDFZHoLxqf7MFzfJ4djkpvW6i2N1JyKq
d7ok3JokSlVfNR/1sqUpeGCCt4LARM1wcUvpA6gjIdPiwujQXx7KCaWT8tMwn4Xz
UUzo76W/hYkfbcS9dLExfoaL6UWEQK1qpp4/4IgUs3Y682VCtTW4OGPsfWtt5yzd
IdSJ/H1rvX0EvF2krJF8WiRIvn5cqhm9zYbzECZ3vZTbN/OVN2pH2AXcLahDhTP1
O+foyWbJIcgmJJZYgjivTZG8Ec2EgkGHDfN7uifOWRq6h+EL9Do6VSPmMZjGZeLJ
coaZRw6iks96BKxREsu1HCDULeAjNqTyV7c1dvc4RTmHrRgRgk02h92mlVf1fPda
/nQR5OVS+fiNmbaixErf8Rj3U8KcoEZX+K7VXPuxmZ1bYWcQGh8BBnGvgFY6xkme
i4xMja76bY6nB27SoyOEdMlPcYBG2Z8pgo9FiEMtZGuKAtGNyRbf9nzJtzYSKtGE
EqyvtFqQB3ghXmMthGoWelKMvlqkhM+LmZJZNB0bHTlhaROM/M0lvWxbgc6ykfPM
AOBQhxMNvaX/7d7LNadTqF5CGVmRjtGlN8UtlCaMjJUzDXQkmc3Xz2qHhkHZ5JkX
vieLXY83eQNaCNq8uN1L9V9Zuci99w/rtzfiG7TTGAyyVnv0MifkSUUatCJ542Eu
p5sgOhIjfhlhB3lM1pInYTyUcp3+QTtIFsFO7YNFzCMe2VNLJ5/j17ji/MwqihRu
U5LWzlF2ZQ9BEiOuX5hepMiqtELQlfYKD+zizkOxYtMUgY0SudVBkOb/I0HaA52X
IZUZX0dGn0b8ogGUtTe5ZYf9g/fw0f3AfgHBzfYngiW081nk2ZoMugGyB9AET291
BmzjbdRaJ86kohRWWMeGR/s2APNQMMY2v9F1NhZdCkeerQI2mFcK/McffL1HErI9
wGZ9tk9bdp5iufNhxCIay/PIZZq6rvJFUC4v8jeMQ3nBrlqhLGBPrLDK/q3iO3dx
0vJqT5IvhVTevP7Eqi/SkzJGO4He4nHPbfLPbBz5caWhkfcds2VQb6FE8k8/RgH+
sD5falHit05AdsoNIn7ueSgHw+XtKodVZxs0y3g8kkDe8AvIWvMSV5MzXg6SEyRw
E9pILSmCcrYtY68Es06lm5nUF/Asq0QcABqTx1U6lSiATM+tT2DmLjzhqoIHccHW
3L0spKSEKOf9bGa5bK7ZdqJr/V2Sq4Q5IPDbJRWjLoqPZMjUyqUMBEpjdf6Rx2ed
OrM9/Oi0XTpsnoF6AXoOdf/mWuZvwQ9Jlw/pE7bB/QFwyqDQB0FNOZMDi6Ez74iz
01EdcWBiUXu4oXLOd8a5441z0uiWPzWAPZbYORk9AXEuXdMXHCQ5+kvKBQuujJPE
AwtI08FwsfxfN73/b1p/L5cIzR1Me4Dx7f/7cyn2doE33b8LFZhtQ9QeL/8NI6Or
qa4V02nQdwsojFoV/Ij9rruFu9uPrbAuwg/Z6BJ4epJdPfqIJKkwsU2j/gHP4LVM
4I9z5BdNPcdk9z1mgosT+DuM4tiHkTN39ZaN+sd3govzJxcBoOIIXt2MpBCG51/L
yWEo6DZJIKRKcGv0XHFIgfyk/Fu4iVgzCACka6ufy9cieGm3RODVroZuY+Y1YT/h
/U2HKA8L0uZUZKHIPknUVIPEtomokg0qnZa3WUxIju+ga/lVNcozfXCAxT9zW53y
tJmVtrWE2dqCVGZMx6UiNuWEvHnCoHc+nuoxxo66Li31Z1GwP61i/8ePq/a+4X4J
GqfAC+6dq3MrjBeHC0xCm6H+IgsUlsGyKIne31OXy/gwva19iERitlGlUhXNPRGe
sXFUU1NaYugXtsz7KoF2M1aZNLgW9Bp6K++1zIWh2GbBX7IDi8BNUBq3RnZgbK/q
AA37+5ZrennJ2BeNkQojTDcmLoEJIQ4GIpgJyG+1aRXJ8rcS7DgecliqJo0JUBwz
cJYyqoistmKBO7/bSvDAD/iKe++U1LieyFQZrs1uWZVbfcGlXY9JB2atYobOA3zU
k/d6f4g3OXVqMss3bsxhqdAN8tqlgKKv3H8L/pG6CDRzL/nx4QCr3TH928ID4H/8
Z+BBX5XUUNxC0ZG34lbAMK2IDfWeY/oCBSfcM2VZ+DA20OLI9o2Em7kMgPeK8OT8
rkTRC+ecRdpxqw/BdYy29sTEXaX0DKL0Ucdy/+Pxl6uAzrUZFoB8xKqSseZmnOHi
dxbv9zliU9dBPIamnqr01vYc42vs/HUqfIYXp0p5NCRONRkUtOneMVKUIq5MxDZV
KqIRlM6Id/J+1nq4tI3IE40DIVaP/VDnxlPxYALOkMMNGZUgPV+h/Ur/KK4b7aIn
MoL2jB5KGKdnqIdKn+M+IAOAepJpe8F2Lv3E29WmQF71JXYuYXJ7gnXLsVOeEZpv
D8viuUg5wLO+vh7cn+argif3U6wjfmRCoQT8u4wJSosMq/hCCmxzQ2QryIPX0mPL
tHnedOp4sepcx6Y02L6KQ7PORSpE4kWm19zhoilseRnEY1PzuLEpqBrfudwtHqTD
ih63LBYlNO78s4DPaCUWKUrOSixrgOGFwET9pCw1kWBPkmO9eJ2I8ELSXcY8PB4P
5EHDOq8wejiKy4SdBRVYAzhkxK/+/2h3PHL4HYa2wEhZS66qG5K2FdQA2v5mkJqp
t/qjyKQXhV8EtKZ6ort9qb967tx4n5W5Mag2jZcILxsNyvFyi8AN9U9UoXKp6btk
K0IZwIc1aTt28ioLYW/iEM9RLJcTyahSo0olBovQezXIJ1MRqNQuftKjQypjo1cc
rc86yb3dcMavfqwci11UUwt9mkm4JAQEaCy4ZFR4Bywj8i1jfbauikLWBYGSMySf
wH/PD8815ikb+3TDPOEdllJ7ZJKh/nMDzDVsFILpAlrhm7NSS5qoNDrJg3mg8sUy
CUaJKrqPA9y/FD2MaofpXZFkoPsRS13+ConssKWujDNpTxKXs2BZGlTcMgJTN6Eb
43khVxkiCBNhUbq50bjC0gUQ971WNIpnY4HmyHwMStnJ8wtQoC+ZTvZU0E9++LGM
7uZ/3TEc0YZYIpETZbsLNi+mpRI1NCsNpnn06JwV0B3054W/KYOWmLX7baO0vxsb
foMKZp73vZDq9mZ1ITrMap2EhykrB53Ik+ooyGkyrYBpbjcYRWQBhsmXE7B+YguW
r/hSUE0DhBVHqISfjPl6WHAEUrwOy/0wBUM/dIFCP6NEATNUKD4+rCHSnwSMvel4
X9n7QCiDH9O8YQCO+d01fD0ul8FioAgkj+DO/eftNoeJYvGwI05uYzQC7EDy4YEp
Pfg0gjoOwwJSyzO8K58eLTHZveVXQQg1KiMvusauH75OLoXPtgHz+xKt3Or8FVly
9L/VFxUNwJKcLAlFZY2d8inGHmZqdFAonM8h5kD1lmBPVzlBZ+LG+w9WshfHIwV+
soTr8DoHleLnMkX3wqgkAifAgdouvs/XKXyrHr0ct13su/ttX3ZbbB/aOcYiYFGI
72w0wGsn6HKMSJyQoQT9qcCgdfR1yFq1tLoe0iGj/vhnF1TK4XyB1QbmjchgdWAJ
jqhen5pe2VKbyeWtbySt3Lg7909U3hVc5CB1ZgrAEq8Ik51OTNudhjrNdnFqMAcx
CObIqnqtDpRc0k9y83+Wjq6qUsX1Me+vQqPW7GJJdbGZvfLjJt06VDT/11ofj6GG
k74oHZ4cAEYFiS1M4NXmia1HmKiIDCwuvC93LqBuET9/myihZ8zZb6f/SjlkJ69O
TwSENMmpnYGBEav+CR+75YND2ksQe2lwn1b6J2r3trHYtJ9X6nEhZPezxVugRl5Q
+BmLcSt4krFaKEsbS4KVv37jrgg/9ePgXkIN/jSQOzlGNgfrb9tLYd/FMMBsUDvi
X/fqugZfSdGTASiyur0zdal1czqfCZLzSBcbmtIow8uuVSbmB8N0Svy1j94TUcuh
eAoq6cg7g6uNW/ou0RheHdowNy/yhIXkSAxuB9FUwV424H8j6AgVemxNP/7xFEeG
zZWyHhYIakeQAJ5YFoIiBGpc5hgMch1fgKg8HWIC13mtLE9mOaoT7SrwfOIJPfye
DAHnHrKa3mjXKOMjeFdmgDxpfwupr9l+iNVWE6abskojpKXRLdPAlI5lXc8JhaPf
0s87IjhpC/pUI3tXpbnAP2jcQJSyc1VdPT7mjB4zCULYuvsKLEvEp87d6p/k5xq1
mZWR1g1Rmpugl4wAVOgqkKFxxel9gTx6lpWh1Ui12MTS2uGdWZH1nfREc660pgAS
PYR7j8r+iRo1kK9HDgBeY0PEsCqnKy0Y8KsTW0xa/4jGqg1pnNVU5D5Svw3/mnTz
9aUdyomdgStWuJdtKE8EcvIj+yAhSfEiK97GA1wPRlaJeNdH72pQSbuCHfzBv8GD
xTB7QaGjPepBpSw///J6QSt91CaRObHfQPsUrOIQuUqDQcr8xZXUhVUSK+yNs7x/
U0H6+B6C/3JFmwYVMaZi0NODXvlhsT8wRdj9F1Bdi0r3oK5gcPR7fa7oIQxIjx7i
sJa+cKO0jkQfGdMNbON18FYQtqWQyspr68ZdYlFXovBBVk0umCQorw/gH5kd5SyQ
QkfrhXoVAVeyGntXSUPoIaETN2ynxhzIR7tQo1fkJNacs2n8Zy1AF5Ys0YPN6dWY
YwcCjiqLhfARAtV/BEHJv1mh2B0DivjILNFP530vNwu+o6C7wrtL6zO9gs8vUG/m
geCOK7jrgiAn1zGqYfwxnuTaQISJK4rbwNDGgB6IRn6pV/EuohPt9S+LlazSK3W6
Nyb8p1ITuH423m2QkKATCXD61y7SqEAk0D1LwqrV0vYuuhc3l9+CXakNRLTjJalr
0O6ZmpF9O5KzyZLxyNzccGbEFwwfm48aW8E+Vc8sHUIjZTsMv2msIdGS5N60Msh4
ZWwHWtWmzY00RESr93INDplBNdIuxJCztJzvt+zLrr9N7BOsreQ1iFdX6KQGl3lP
esehZuBYcXJAYL9uuO+A6JnmJg9XrTKBQ2+u8eUMRs/0hJ2dApm35s887GqOx1Am
5xx4pNw6IJ4Dmjd+SeTTGSS4l1+Uwqieui8xzrE4lACGqq/o025IlmNEHUNU56W8
tTQzzL2LZZgD6ZiAXDlNFV6bV/WPFRwKKRFu+XgrKBpPNhKRdFBNhj4SDa2vlyEq
dhSpXnQ8Y5Q0SmOMI5GcjIJGjgJm1/TqJngNkjzqaPrcT4nGEGHNvY7LFS4TqpGV
k5jDEBC10a6aBGHUr4AlX2A/Y8J5Kvd4YakxFoCmuDi4hhzGw85C/h7YnEmIzVKX
semB6pY4cZmpOhpCN/3OCtvnCQizWy+H+xur/z3ySBRLshNmFQ66JCzHZsDP/REA
rkU7Z1vwdF1cbgGMp6e8NFvzZyYu+hIZt5BTft4FsKQYUqVaNactWd60HHC0UaCw
PbfjtDZgGDHPRTr/v6GsPXuk4pA6DDaRs2+IaIfhl6nW5H/JZxro+1tt7SXUtsml
rafkcZtgonA1yl6VXAFJdYkMKrd1EwMwhs+XcabwVls9q908dpZM3wsPX76U7kwd
F6RG7XVUohnToSgP0Ig58oC2W2Dz/J+9tHxQmtnD+plCA0gWCmccsj6+3DoHhBqa
TukJbLwOGS3qezAuAvDQkD1a/t2rQPsbq3x6LASPsUrfPg22oH2DvAwClga3+3k8
/brcljgZfvfDs1DYj7Flg+GKuDi4aKThNvI5kvJFKep14ZWyNf650E8WF3GcNg5p
/3gzUX5Luc/yQhauTX2xs1OTaiPLhLfqNgvL/oTx+V6UMOQWtuJITPogJUIr9iWs
xgrdX5FsDOZ8s9eUmEC+ntJLqW3hGg+pafNzqnZgZpjkhjEXxt3eWqfHX8fKJ8hj
s3FVBY/KlHmMqxGBMV2X9Bbf33IbBScxd4HgXLMXrHuIVO+8ItJiunfJlzcPBVqU
QVyE7A+l/BJi3ygAAgTYgejHV1MzDkYNZvp0PDbh7+SdhPmNfQ+O3QaQrtZfwZlR
Z+RQ92KKooUHI9WGzsx4v7/yJzubPSqsC3Vq+vvNzXjpVQ9Ihxkn1syQNCXyW4N7
w7iOop7HtpgbXZyXtTHgocEBeWpqpw9mUnNZruv15ectoWxYVQasTjpAw3kBlr8I
Pu9KvsJnPErbqWgrq6XoW45FV9d4ulhG+3g4JPd4hClp3VHuTlXNijAv7FD0DTLz
ZFv3GF+PyFeLQ9szcGTMSxAnt+GARyfomBxhiSLw3sBUULAArc7EN5ESCtdegjB6
eEuAMgOaGZhKCsX/QElQ30Zzf3zr9bKz29vTd2m0H+hJTUUYyKJ+WlRSyGqC4Dgx
1yjhKeck7P/SMnkea5HzTXsXVu11KAjp+AaimSuyY654ToXEBhOqHjYYn4uPtaoD
aGk2RFlszRW3j8XtjDdrftUFMxMPtePPaYoH2uNgDhkajFFLPFiPezW8fqABXral
/2EfASM38LLdDxv1gEY8vmL5D3E02UdRg41UUHmFmMT0aJ1oRFyYFiBz7SHePtqR
3/6HNU9QwX9FlThBwZlpIw5lwxwO5+v0AB7FC6euyBIVc1/L+5IK2eaYTLx+Ycxk
hcINZMxO+XNnHrMG63q+AJJNFc8jFxiZRUPtjYLkkoW1kk0OZaLZp21siYiuDBDQ
z7DSUWyNIp4Bk5blqcrOzUp/gtbV02XqufIVb6X5cXFrK1A8Azm6IXbrxmEcigaH
eDiCkSNYgsB3w/XoqSY7yIHqMpzJLknue6D2SQqYPc1vBY4v2wrPepzd3CdCkr+S
mlgEcs6sISe/ORFpchb6ZUWpGSOteu55PaEb8TzTB0tuC/q9R8GsMWNRPWANtFtM
EaX2o+LgadGTCroFLK+IXAM9obOYE0Y9rRVGaxpaUn05eIzpDqv2GDNMkqvCNRJ5
0KZXDRfEfyStEuuUrjStb7/x9VOxrKv9b3rFU3uspkDKbTeVNY3il8s3ovUplhTq
5Qe9RVcx0EwaVgKPACJDDhOb0Ca+e7DznWAxyhGfd6GjprzhDxZABO2e5WHt9evQ
eQrfmXRynWGnAKunI/lm0aZNiNr0bcj4kPaoSJe3cajdHAvCAw3Dgy8Bp9PKrJrR
iR9BaCEsJalfjt5ZwZ1rpDxQrcD/mjj1CZQwdfSfumeyzHEZ+wJiFzPikNRRJRy2
aCxiciXb+oZIuoAIg37Ac3iaJ4FlZVG6yJjOapRu8gdbSrcofDWK/sZchOuFleFE
uPywGjhgSbihGb7h18sDQVysYGaHzapv52MYn7SXWzqrmUSMaZ+3U2AHqb/vxvlL
h0l9/2WEFNs3LGo3uhkLJ1Sc3/3QCmpA04xFqdIaPNsYg388MOyw7eiuq7Y1W+SV
NCgfOp1zzeWjccAQ7I0IZ3fx6VO8er9R2dJe0YTBHczzsF4jpLlB41iulH44bXqR
uINNidKAApWg6LjyI6lsjTHRuY/Z6ztqYGEhdo8v2LFvRiEh2DCRFyn1APdyr+Df
AalsaU6bw5AtkPVEC05tj/6tSltSKQU61T8iN+5n76P7nKWee6a2FdCjq1tCZQ6N
0Devad3cAWHQTiZaKGR+Wl4dPwJPcuB2jRmBYvOFvTCnod1Vv2yKixBVAfdVPeSJ
PEegVkIOfPEfm+IVhpPj0KYOlnfVUL+pLoVS3C52FQd6yqNqWWZMQF52oNjFfzZy
IVeMtl+k4maNXEwlp49PgQhyVsUBDV5nrJmp0LNFpZWtoKcRUgZlIzg4D1p5R+I9
+e4ftkS6gW2Ww87LsaluNty2lQof0EfMT+6cnJdkDoucF9Vr5pS307ZFUYo4mG8A
N2JAaPDGehSyXL1hfFklKD6uwAjxmtpdj2oZ0TTSjEUQB+MEwKDYd5XDkTSB0qyW
7IN3IEQ7/MjGLJxgzxz+mV6flXYLogAIN7tAG3kM4YfSQB9cnlI8vjUaDLyCGLKl
CYGdHRqOzTIGlYk3hIGWiQaMqILt8gPfuV1+rhPq2DnUfHWaPJ0zyrJgoq8tP7fk
ECgczIa6RxEUeAuyETFYKn09EXh+5W+G/Z6D5umbCIHWThyPh/vyIMU+52W3RfEz
SPi41Y5BAXosPU+BJrvqJNzo+5aHMpADFOfZzLYfqMqLGNULPXbG5l5m9xsCopH1
6+ZKUofSwNCDn9N0KaV020sWBo43JOtS+rjSrAJ6VaiV6CoWyW5flbf+zRaEbuqJ
opNf7iKlfTYTIaOZg8OHPZQDGpwyWwKU4D7cuD2WnYga2fmNyVeQlpQYhqgEI4VG
tIHyQJf0XzAp8wl7j4I/IfNrMYDUS26OjdYltHj50gFRDsJMCI+fb1DBuz03i56/
WEM3jkNEdDzGthde3OORU3TbUdCtXSX5TWFxADAYQRrnfqHNuXKDOfnv0kG9q0sr
eiTwpmWPMVjO33T3LGrG1uXmOK+GCdJwsLRkYvJuEtj9ZzlKlpH+cFc2uN6KpZsY
7eqs9ja0gMUK0KL0cPMKCaWCV5inYdn3WtZJ1DsuxwU5D30V9Fb8XjDKcD90h5Kr
rSQwdsebkNW9H1Cm7rWLCfGBNpjX16NiwEfvvhXRvke+uee1bMpvTBQheFbRa0H2
WuN05gvMChoh/QpvJl1yy8t20F2LpHyOE4IjbkHZZ3WlevFRnDxgnK6wdWSIgQNb
LVZHrv+b8Fdq/Zu5P9O65paeU5ZNHClli78EFJyLlzuYcUK4Z3Ikdrtmz3fQjAu9
KUccLW8M52AcjeMNYRCJebxQQwJzILJrx8QdeBIfARw9inLFQGS9mBQfEk/nVjnl
auo1lmchvbcjYTAmW8r3pt/jm0nmZMocIiCI+Ut0UItzmKqosjBByEvvdGxZrosi
fBwkEnoYVf8FTXRr21JhTKgXxPMV4BcX8NyIJgfQJAG8n3EOzGxbIQs2OkLH+G7U
ZLoQ5NllZ2owJ3nGzlrxtKluEZpBRcvdh6Kv/oFPOJHJ14z7CXPHEBSbQb+P0FQu
miEYg7QMZYEWGrLZ2nwsyuFD2CNYfQ7d7lHH1ol63WpTmSSicNHemU5UpE8jdebi
a21OpFczesBoeEaGYH2L6NNj524uKJUfatsi2OesVUwx2Et1Y9Spmu8ROACgfV/6
DXmxWgOyk0dNEbZ+YN3itgr5IaAbng1TK4yiWqc2VRlQ90cy+ZVcViy9c/jI4eZv
Cy1Ye5mOaGyWXknov5/THLPR4n1YBJuk/m5SSc/Y3v/x3nlZkDCd4kubzRhh1dBd
vgbk5y4mMDZnFAY89/HdQzVBnZrN8PWCeD1TuqAsIO14bxQ9mAMyKXqhCMC/cp2s
IW1JRlE69h/XQVkKdqGwvhWTUwf3He0cTJ+bfmtDzLeRXrAKdtpNMS+aKr9wLaji
al4RY40SXJ3CQulH0k41f5FF8jUKX2JRnrEdAsukZqXMh76QEhwdwBCWZjt+Lyub
VVRELrRvnX3mtbpBpGLCH5o2XBFcLuT/4V2WznfCvS5l2b0T/f8C6g46PWfwg2zC
onL7GkPKdqgeB2AzzARkDw3chE7WeLMUYqkTqtTZliz3gbjGu9OC/wPSf6U7J+3F
P25GIDzuwdeEO/rxZAFdXz02hM4XggIBv8wV8Cm5ZrEKYZasCVRHm5dgFiBZaOVa
SCIiMBRRzAK4aW1dwWJ3hUjjsC3ZRZecffGWZAeS8B0McmeiHGyxyhO9G9fPuTc2
o05mdUUQQVCfu3TFO3XZv3DmloEkPHaTfhuUzs06DXHbwGkkk7Onfep6WCc8g6R3
mjFic/Fe2yJ1xc6/kF/vo70Klyvxpc7gUsdq4RQMUq9AyelJ5rAt110VIXxhEakp
xYppjjA0Sx0DZNmBnSoCKrCebO6LljxhvjxEueHu/WunIHfCm9gqkVx6DJBgd4py
zExu7tfqiTFNPxz01I9NGUQQ4VlIKZNFtgYIM8fUDcMpeVjhP3t93OTrUvZL6FYm
rNqlBxAT660Va9QtdixeOLdv6zVka+zJHjX+YiZqQCRm7lGrUDXKybn2W504iSZU
f/HOhLITSFO1BGRWKdaTbJ4lT3QtYf0FeMY2YxNzQGQ3V96uiM8ksxQ8RQC9ZriQ
v5axkCmyLYEbhPFM9BXmo8nCAop+8OoPgINiT55qBbbmFuK+uJYH5+4kvRbeLXYs
Yf5CVOMYWm0BwVYiZWJj6YegY+/HIjnSr9fQ59sRPmK6ryQxlRTfz0sUpcH6PUBz
OcEukZNXvweOzyHvAadmu6yy+T3hZFDdqbkoSvUPe6WG5xGL337fIiRN50z+n9Nl
/AfHXDr/rgB/hKl+T86IJuad5DGoK7ur885lOHNwMGYc5uJ6OjgEwnD+rgyDUhSz
m4vtuIC6e91fTN857Wja6zoGJq/HRRCMrRQ//pL2eG8my/Vg+E8E1qC3cYhCODsW
s/7wbG0+NHAZi258HWaSxsJOKkAtpdyjfEWaqCezIOLI/uwcb1JlNnd2+CiPs77H
cGzhZtxPjyqypc973kAfFhfjhLoazliOzOQfZI6jS/WPclZ6ccYwvOmi28SQuIl1
nQjkUQiuFJP/KeAVE6P1sgh15FI3Bdl38DZC/I7OMgVs1TMgcAgHWa5RrZWpyUUB
9mDLYohlzvQJwX0bEpzzGenE6qX+shbJXeOIjBGDdtbWZpojciYFK2RPP24NOKnp
PYEaBwyJa1QKB9VBxGsaZcRsyG6D2VhQiIgO+C384WcN34u049u5TjDbMwWPOa2J
M47ZQmjQyJ19+IDAKkksyhsrthV6XHWXwW8fAIaHvbQw7Bd0FUXsi8ui+ElZ5EBX
+CFRyb7iS+TEHQHTUiqnKKachx6X0MEG0Jxe64BT+IQYIt1pI6AIBiXbOYj3YNBI
ge4CS255QLw++Yh6umyHrEK4fqCxfCrPYeU1j+rgUhy+WpMaGcwgHChb+aYd7LMC
Sn81uigWPenh68pKPY+LiadwqM9WEPyWZhrSMgefBUTR9C0OIXy334XuZYfJ9GS6
4INS76IPjWCr0RMby/MVYcizpBC75qA16PISnoQKkvkFiDI7eVnfJ2IrZENznQal
IdC40WoiiJM2CtjAL0ubUPnF7dn5U/wSVkuoH5UUDfnxtEYsLAHVCYMaFpvUDfBE
1+9NvctSBpZZemGKig600MUa790LxplbJidpEaYE14t0SekBHHkksTJiPf46ClY4
u/fJyYCGToBNwiXt2qwSWoboDCre7NN+rO7ptwx5khTupiE7h3HgLbZANLSnoCUg
AXs48wb4m6gSBy0JgzXDflHAPlV/xTTwKtcrDzxGxpMRYkkjPUG9mljRaAr2zdHY
9QaHwHvOnDQ79Xu9nzRKi+PL5YSDXSdfg9GTiZWZBmrM1Y/2dEZ8HC9WBAjF+62R
YQZZnnsMH7+1DyUYzeWTMWk4NXAoVm69l4jxAjQIsdQSXPXF2lrfkJqgwg/BpUnc
cg4t+h46tNPBCpJV8DR+sffeakFlPAaSzSSpPnfQXae5mV+vfp6DMGWgBkEXz2fe
1xGJ9UDPYrWg1FFWPLx2/KI4gjspAdhiWr4McVKP8ea7AcaFcqtj+pyvGwk3pOhP
qgK4+LH0DHoBDCsn9de1FcWFeLt1ZsJmkxgGnMDW71VfG/BIyLfi05N+Yc36+eUl
MtaYLkq9Sfi+xmf1RuNnbccpa642MJTSuS2Rp52Z2eIX68DV411nJkRN/rns75yz
Vz4OsUEIe48hVtjvu8RYt8PNF/x/yDAwite8YaTU5kzFye1CztGZcpsqXWOnok9k
eTh/Rq0r+hNn4g/gjcHN9K/YnewqBKXbxAldO8Xft0CNBwdS+4oFUkR6t9krlstJ
tcLn5H9yQNdlg28JTT9YE9jae7QGOdweK2Iiskc2Gm5a5iaV748mbTIomASYgrDK
dO6POdiRMZu041bxiFwoqmrnDQrol7HnYcmg4fjfnBu2y7Tj7p76jzuAF2GJepYD
Gj16kkTICL+S7HohbhOERlwvsIV++e0E8J7d78Ekx7/7LARP9rQ0RQklbVmc4bPq
wpwCPZbOp9ArMd83I4JQ0qmuq46CB00hnFxXYK6nll6AN1KnNpog7qu2yFBAq6Hl
HPdWBRPivK3pRIkrFlt8/GFjmZ7v7uwjBulCjYF6KGYm6DXKrtvp9AeSENwfOeCw
2OWy8Ya9uYLVWgHSLotNO9hRrbppyieccTW1AV4eOxJPXNSeRbNG103I14vo/cga
aLoFaEV281IA/xDqoLp7lbLSfqeMh/LRGU90nOponlopK1aEzD2oKpFMUeXvNIEY
QRfTZ01VsTnGahXGsb4jALgb7eZJn5y8fOaWjQxedgrXEnCfaDtSVaWWKwo5TiX0
RLCZtFif0izbQLpFG/dET6naURo8knyli/gwKJX23+WC8ZCGQCLQDo2vNwdqSB55
MKRuAxsmF5oE9Fqyhdzj0+TvlmZIAwvNtJvIeWbyEm+46K9NL1yjUe1ABDhgzj8X
BY7NssHa/gEsaRPy6et+VeUMexWzTc34Cd4+zrcy/fNT4zK81DjtmaS19sgFDk/m
c1e9C1lTW5DGt8zWT/wBP2CUSvR58M5DLjHpR5SEwluJoKdFIYiYM01XOzdkT3kg
T6pvIfJ9PlimE+pZHZXFabdKZJ7Zk9ZUVnhU3iX7kfnW75/zyPgSewXWTzzIKFx2
F5WLwyYRjlYcWF4RW41AekVtk3b2+CQoN/Uvaoq1lSl0XQLCdbZcFG6BG8D61CMP
YWFg3s4E4IphzyajV6xWDBsf69xduggkWH2OOr6l+RWtEa6GWrWSJkZFEdpqY00C
uint3FB0aKfJiTxQR/4dz++vMA1hL/o0gio2MdM2mOFlZhc1TDhEliEWWx4i9ZJy
69UHH/xXjTeo02hHKLYQsfj6VIS9vGycHxV29XikRrUmjatUocY9cbrYUvw9G97v
SFMGTkU/8IMWAqm0XtxbD6YJUGI9dpOQGgH6Bk95bWd9iKeduRBZtfnSFVgWIyDo
dhctS6of/AZm+z3GgLLJwAMTvCO/NRo/Z860yvasVVaQlvGZUC7HIoidf/ei712N
KW9JQiGruYHtb+rVd7FZs3m5LNRjszqDUiOZd44mnkg1WH2pwCa+ca8D2ag9t6Sm
DPNJaBJZiv4Lv7rmYKkPGb1sHQXvF1kcu4GZr5mKpiQitWrsWvkxpmLbON5mwqYk
jEBNfhQvxJnL6QnpAXLKKGf72udrXQBrF7WXnS/54GDhBI9Usio2w23PTeL6TjM2
YScLDgXI4wWkPz0LFHsveS0aa6bSG7pNmRs+eDsLD2t/SDn/po713Ji5SxPRWbSs
Y0PH9NmKtkuZ/ijE593axQpNF2Tf07Nsjvo1lSG7HQxo8xGYrfTeo2/SiegoJbYq
pQ/3Vt90I+5ZXz+lWpq0WHxKccf9Egin0/QmwBr0eGEL6v14uewKeHZO08JwDta9
owrGDI5o+sW/tDDOlcLEAP5OXLGkFMERl5lJ0vzCcbLkOWQHKtEVcFedU4ua9Rep
nZHiXd9xMRHMmf5NNfGCp7GSv0qQ1AF4EjSccfWpyn83ijB4CRgchvL6sAK15poS
SpjBsiXZw2aGV+G8qZ1W0SYQtOKZcHlmdKjkm7OuXs8+LD10mPj96AGpc6aK5RjI
1IeDc8J6ZiJKBXCQa2YtOYtCc3QKNm2/HQ0b7sxDpjyZqg5MJnKhbNv7pGXSIEkr
1uH6UjvoC1qURIcSyrl12+iqxqhuIDsDuAfnRVEfhaEEF2yR9RJWVHiU0eh6Vjbp
H69Bl7fodSpRIqhAc6ll/C/nFKxDGlKGDZsbauUvCbDk7SMf+x9ZQSGoJxk44cFa
dPLj/K1kLBDf30HsWzfsSa5QJZzUJn/fwb0EFl1wdDyERTmPf4ytNo/25yJ8Iuf7
o1hUmDZW/Jvr/hrsAREHaWOmm5wYPH8eFQBh3++lr8EGGOGuA6otao5rXAICokkz
gmvg785+6tzhhx0PbDTkCgxQuTNYcQXdwpMPJT2foX/U7OOjnG3Bt16yX9y26DuE
rUYvDimHlf0pgHhYWLdSHcNtLWKGGuyXcY7HjLROgVkfVdJEiM3yL7aF4kTera0O
0yZyOFn91GJGHcMFErRmIC9Yxzkns3TcLGb+Qu7dPmh5Wc83Fro2tepzX9eXifas
bsjEVogiVX+SXodwK2LnQJMePHddHCOgBAvTm8kWjqDvlrb3VyMLd6/Wpr5VcsoS
94nEkYt1Bb/MEnR+3fVwJdXjpzVtus9PDQDsolfAAa45jAgV4883r7TtBFi+4InH
hwu03RQk5eSxbZ+aWYIgzmwtqCOGriRfGno16Mamqv48jOjqeI5GbHwdrKvJHB0X
D6EFEQm/YE0GMV/FFZNlynjOW/ofA44gf8K/1OnJHNzy43K1JJ921jg8x+/qQocJ
MVl5Po/Ey2IfFzzlh2JGCeCjNcJTUGU99sqLt0NN0cixo1Dc0xDGtTybhbvoGYE+
yZ9UYasp8Y5o2LXoM0WYVOfMzncytaw1bZZQ+6S+SxcQf1pJ2ZfTOnDyVWxolRVE
G/T7cOTqbDSz07vCcQShzQqeJo9Ihgz77VjHADOTn8p61Dt3092ZqLqN9Q6Ny5mx
HYf2/SxpN3/1+ladkxYI8OCJ0A/nfSzhgHmtWROFMcluVRl2xDuiMX8ag+ec0G3D
uTra+47dqOJudWQQ09OU91/WxhFBRe7qUJ7N0XHs/u1O7C9IXLwNYZ6bYBx08636
G5IsIbQ2/XD7sftYyPn2Yp6hpG9xEQTJh1bx8/QAz8ool/XlBT2B0RnoMjfjlnz2
oWhcZUSCEO1iKyNNLjF6PkznT+927sNXiri7XgGYZlWN1n+IEH3xtVFcTMhjqgeu
d8OtspY9tV8VIzm6Ysbr3lBjiqKjnVkx23Tx9Z6tzPbPLXDrp8WBaj2vegfbEchX
Wae3csEMHVRINJeU9lF/6297ZYnNgPB2e/4eepdkeQ7/uNUpGhfsbCbZlj3Nus0z
VLl3mBPa9Dyz6xNfFjF0eQ7PLmTuW/9h7nSI4EWb6OqmaFKdtLCNGPgtIg8Gtiqy
pNb0nhacIU5nHuwwifC0Sl5FwZH3Sg8N9I9s9iXdwHtMNJryj8hu0bhDavOe7Uaw
8QTjca03m31aSq8hX8R6laW8DrQJLYyqKZ98d5vYS5uKf0L8MsV9HYSzBx4DExQy
qujL8tb8PZ7H7VtEUkQUf47mEJDoT3wOCsX7AC1YTh5ZCkcg5CWNRSs/a/cTTzUv
95WzCu7MzCEXQ5GViAhMubjUo7QBh8klDsOLUhG6w/bzwHXkw0WtnTxlM1QAGTbS
lwY9X7IZGfM8XaCuaSf6Uh3GmB+g9W2YukrxejSBhLkHcNfj+ph6Iv8Kul+FVO67
GZAhrdy4gy847ZjEpr/T+QTPO6Bmy3YQ2eVs0jeAhxSVPLSpszS5Hvc86aWOvhsU
atGp3SLcLIVB5vf8jSdVOM6Lhe8wJxoHwPdX4RAAarOTK9NH7ouzd0B9CZ0Q1h7c
xQCPl9/B8NQ+ZzAGksDyYBYayy2c66q3w0MbfTWn1rXQ6I3xgocCzg0hGFIfzllY
nFYAh5L4cL+KoB7JNcmBVB+zNHbnH1+9XjA+4710eIw6Tp+SW6wLlaW/+3FMvFcA
0p4v6B4kGYE42wtlPKrGLBAtNzHSdhgnkk149ECWzgfGuYVfigfa7yhFhPEu49mC
YS4FC1EjhVakcL7Io6lX1AiuQiRRy41ABHDfH/6myzUK10ceCceQbRo3mJkOnTAX
zVDlRZDGfSAdbGmXZLR2odHGdiPvpzJkdtNFOcj3EYC2j12l5ZDDl9YrZEBH3dHY
ATSDeM2dWt/UKVzLQ+asJc43H7j0huZtaOkEsrlpNhfh0hr4SjK4pvrafpnysCGR
IXLVmegas9h6R2ZqH+JDz0a6ve1Qg5exK+RMUngxiYTgTtWbuknt/aIrcfODd/49
78y3Vk4upHdE4mZqsQOmFSSW2aJMUPXszEfnTtjOnwM6f8LlflnWRyGYJ6+FQGih
Ja1Dy0prCKcsnTOKGtsLhTwyvZ4b9FH/O1VLl20OiiylLnxr+BzYk/cC65gZDAH8
sxY0OYuBBOI9rDDQ8ZM73h5TfHcAmdDorf27zYN3Vpj/1+f7tSmk+V4EihCMRrQA
ynlKCkosN692zdgLzXbt81KqiHIJfcbJeKSPn5ClpvP896SSbApWBY9mvrXeq1jx
QYuSumacS0vzV6fRuhdepG/9UypGreRvfuC3836MheT/j4N196T0ZEBslgNLqG8o
eC34EtYotgSoLytdexyk+eUv+GNIzScQkDrpIylC4ox9vxs2LGYUa/vVJVRZUhjK
xJn9X/evvfl4kjD+y5OGpBmXp3JCsbYEnRYtM453Q4nvFjMtjZOIv1Nh2+aCw6CL
YnZC00ILgjjktqxkwdMGxyJQ0IQWNhh3O/y2NeaDTJsQgdtLXP7/rhupmg0dwsIa
Wv0v6zj3ytgZgRe/nfn5xZfKeXd9Yl4NIFv8uDgv6T4FvLSZp+qs4vIAhS0hszrP
GWw5nJ4pZJNn+JwiMM5TV9Psv94O1Kn3yDkY2TdPNZV84QMHTspUGdwfB+oUTovY
VgGNeaUnl8z1QksXLLWrE23QMY0vG0sqwk4ScDAxqoQQPe8zAZYpZxXq3Pifa3Wj
dQ53SpnZd7TQ9nAVfpxu2upWsVcOFnenJbsUSAqb3lT6toeGx8JWMQyVB6aqUQEt
ekBOHitnfddFZm6erSDKIG/YlgVwRxP74TIOkeLmsTZw86Y9OXdShPsD00MUGRVj
ajeZeJmY/mnrgdkw0YYCgbFq5Y2gCfxLpnEGRsfc13H5tjkilRQ57wOiJV+ud/qo
uzaczLBUPymzVkDYkRsV58SfNNFd0g5aSdfOZtkILrOHZmX33mgTBy/Cg/wdsBfk
AyKGC+k5L16HrP3/Oh6JTs2zGxr2Nfesp/o5lX7XgR6Mn/v8mY4AXM4GtEsYRIj6
cE98gza/bUxdPppEQ4ojFkJ2jyJZ1QH/8JwSn2uJDISDtuvg2OC0B+cNOB/fgPz7
xLkyEFzA8l5xbyXM1+AKujdo+5b9Zik8cndBwN3u0A7yFZqu0DetUvzltXyPD3Nj
LJYbyC3PciqhlHOEQvPqN1QpJ4BhVQTdC086/2DcvU6fHFmLJjq362hVrdRUDx/k
O23aZq5sX3eeam8JeDYVc+Qhu7ms2sLCtbCDsfqy6+AaBMn7wdLsbrZWrS0BL21J
sIAy4xkW5PiweLW8ZKpbFips5oDimwBRc2Wl51iichN3DGV08cYk5VFeASH9Lz3I
8yEX0whkzN5dNatDvxuA8mvF8eoAU5Uk0f8ArFGn8iZ3zT4abwZxPPrF1zylVIF7
kxlWW5JAn0xUHusWMMcZ19ZCDHLbGN7dv4Lxy6TB0NuZArkV2ex20jv42FLGhMQ9
eaTZZmqURT/0piwsWldqS2OWX19qIq2bVOjak8kYKNyjjnVhpf5Qkr2y0KLExq1z
doij3J6Zu9W9UKYTrCvdByudRN5B0W5ykfajl/ueZjy1aayOUSind07t3yRgEsnM
tX3GsLB2ag6DjYkPQq3NJIjeuPAsrgg4SPjDXFSi68yBgn0XdZpx7gzRV2rAJgEZ
1rI0Zb0JJ8SdddmWPy3sJr7UAvkiNkqklQ4lWjOa63tcujJzgdb1rBWrkMvWStB6
0Vxm7FK62Y8sw1fCoR7+CPFFSr+6IYDYn091skGgsjmWT6e7DHN46ENmiFnJd067
g41haJ1CaUWj1ehD/pngoeTNt02p1xiEttmpB3TZfICivIsLc0TJTqAcjWwQyG0y
DFQS8G4N7Ma8Ny8h0LH8xOGSkSPFjkgGLqlbduMwT0f+pNduGAkcmAhBWLubDu9S
CodbYrW+XnM65DuDklhMN4cGAoh0gPmnRK5LWNayWvGTsMsYv8oSzgAYFlUAqxIs
e/plxFWS4V96gDVBMzX41dtaf3zhZgGMtE3Hq7aRf2MPxO7zEn7fr8Eww/dqAgQb
gpfNfSfZakyFEYY/wvO7rEhculpMvGuyh/6GS6WyxBrJ2r8yknvl7v3Tb+F0zVuM
l/0ighvaYt3M21YJIM2dReTvonhANsPaaivVNJo8a0kwbIj2lW/QWI+EO6/lmOQQ
knGIxJl7bx5fGv3pa92A5xs0ctGAVaC/812uG0VOxdxHOg22dElhDUZG97gUthj/
VoOQQ1V451hyixlZtyTqNLCmsQ9M8AGCgo66OVzsQCSCMhuzkYfOc7Fg6UueLh/3
8ihewjNRZoXb8/SnmMMYz/zCECEb2FhDkzOamX41v5RIIVYekdoRnO06uRyKCL/Q
d4oDn35QTLJ8DKlddnWrEBTWO6Z2yDqh0l1hZOm7WpzeKBzu6Ej1F+9vbWjVmnwj
WxoKJz7ipIR6penWBbPOqcRfF6aMbJYOJR+WCS3UuTVToscotTP9T6BodmH3NC3z
qPM1EpMAhZEsAL6JH4QjPVaN9z+Q4HAi1cjXnxHxqWB/nK2lVeCOJdhlpG9VEKEe
1cAIIj9utnqdUPqD91pz9MCt8lgjzJEPwAzrYzXt5rKKEiOdCGVfnGjGFU1DzbxD
IWTd3CtMRVpf0j/8PN8/DVws5FajGXUAZPg47eRiBK6YxpuioVx/u+eVxkBwkNwk
xAcxbC1T/YFGcaXaDmWyWwNbBxe8aX1aTDx8iQR2MP2f5iS9vNjjVIh7Ryro8pF9
VnIT+Qj5sBZeCnaWX3HjMj4mqK7zqtVLur3gh6dnzpeeuHgaOaf6NLIaAlILiYIH
aV7/xinpaUXFVQSuux2LaJY//G9Tbh+J2CcaxjAIv0DUtcCkbwW13TU3pulvvXd3
rWCxqayEqfw8u7IbqiiXg5oxqzup8C26gN0CfurUJW4J2m83LrQYsWzxbmc15RvU
2HREGw0KttYt3Ie7RnzH0cIc4pk3UPKFxX8ZK9arwYKeR6VfXkZ7JD1uTk0eoSxq
PEXq+Z3ENdx/bR0X2sGhmARjIKOMnEpTMictUOnJRGlTLjsFvI28W9f4Ol8BuS5V
KzC8PDrF15OZBC9dNwR/QMvO3hlnr7ECcSvFBflwsym3rnnvZKaIbeuj3wwmWjxg
9wAiYceD35lgy96/Uh6SWbRuhLTiQFh6VagVePVjrxbozFm1G+fJAvoCwL02abws
rN2J/Vih5iVbHTmoQ6NPlIehu9OBPoDtsUCquPhHXgOC/35JfPoBIftT5ylHGPjR
yigEKBc2+RPKQnb4xB9+m/MXKRW7fuby7uddoouLnJuRosLimx3ti2iLzIFfxTi7
HlUW7BdjC1iFchH/PYARBV51IbaUyueJiI+Xsghx3OxKPIwzvudIqOf96ASGAg61
4oqv1ypMvjhxT+LKY+v7zYU3u0bFzUb3TDVIl8AGWrzq1dtYU4bepJtoIBRJnXrt
/KX6m6ExssDo+tO9mlUdrOPf1X9Y5ko0BbGs+rGmPrRY6EalsrB3ufnGSgwQkyUF
8/nfSjCF0l+riCVg64F/JiYHEEiQFUnjLRGOhcuMMq3z/fHfJrVffQUyAeJrXELu
mN44auWHRLS9BFLgOh3z02jjvXyKmSJcEwJUXrKvO7JTMazwY1+SMvLLKNKAjcvT
Y/WQLxTlzLTeK2tg0OX8G2LJKivDLRrrWpZp+efTKPQxXRN9D5r10JsBkv8B2Bcq
DtKjFNlHUIxt1ZJ4ypN89itZbVB1+qRu8zUBhzt1w5zSnridosLeJ6M8uc5WrJs5
/OrFVa6dXH4jY1oiJr63MprUhrBecMOcOcLKmsYR8M8J9YigKavGugAiNsO4+D6Y
/bWIgNv+E+ZzOHYCyTdajPLANzp9xOs8jfq1x+Ihl1IedzO+JcSQe9gVFa2NMyuP
PmdrRqAJ4jdmGP+F78SaqGs/8o1zV6lVW+tj54zwrTqGsdfz0R0zIHF7eLb8NpIc
RAVYsOur6KOqRxeh1G5YAzLpYjUN/6RfGRbMN3EcsfuxMEibyITv2FDJlM9z+LlU
yXwwH7MknAj9Zd7YEqdSmOEbeg2IU4KonVUk7OGdglBopj8H+apZ7gc7bnc7ghG4
qCrib9lrrtZm/cgT+OP5fg3dtFyYQ4orKpoI/L9itlaLswAP2r7KeAOg8NtMiFEX
FE5yof7RvS0HV2P+vttW6Sx354n8qbeEf7SyN6+A5s0ciM+OA99S0+zV7i32IKGV
47A00IVqIzx9qL1q5FxS7VEHYLBLonsFE9i3cjywHDxE3uvkU+uz02Ee6e7N0vun
Wh7QcGiY2oJ+5H9yDPEieI2eHo/V4o5kIX06D7s4dJYFWkchs+SErVMy3UjIIpGf
RqPDEh3kI+KCtm/HGNNucuCX84CcUDr/9gJOuDQgGRbLY0BQMkRE+1I74Yct+jp5
dQ7uEmpgwLAJsl+AJEAL2Zyj257TEfDj3QYPktofJZRwOdxuFjQMeAYFhWzyec2v
geb3GpB/krrPNkrkHGh0IKV3YVYKnvWoR35hFEBP1SQuwxpUV1jzCjiFCAbeOdGt
yIWGLdrCuVMgEzhd7K+tvLgM0fTMy+Aix6N911EBZX0M0Ls4hj0BUPBaSU7tYAs1
VHXzOOFta6rm0Jg232D41qrnpn4/bGDet9i4Kr4ZVaNcUijkCQCBAGQLle5R+bIQ
MyFazKagwblCdpI4IGE4tLkqjd3BZLaEahoRB5Kg4/w7tqx9dTla4VWhEaQ6zke9
ontseQnVgLLk/EmktdzlY8fMUctU/i6dUQ7V1MGdkt0uvLBeMtdLvTvaL2i3YRNU
furuNeSN3A/JNbpDdX9U1HLLmqDA/x/L3DclPwbLDWgq2Tn1nhoKAuYJxPbw3wMj
wjthix34FMfm8zQZDNGValJan/oIDr9iFtSKEpmE5ue5ZlRRlnilWe19Ajg4BzOd
fMGQJbuktBIrsKIagwgdrG3O5hWajMvnstVZSGJ+U3vO5blpP/okID57Cm89OO3O
GEqWZlCfNlfyjGzoeeGtgX/O0Ab38bPmYUOqBRUHf7N8QcAs1x0xbf6EpcY/zNpk
j9kLCl45qstZu14btlHcGI/eqgDMBzRAuoRozTn198wRzUG+xA4e8b/I2S6MpVP/
9RQPqExPPRRYJDOHPGc97AWPKh7tmGvRjsF+KqQLi4K6cZbaVzTJI5dy5OkkCFNM
Uea5NDLNS3wLGnfDtfjXnT59P4ZHmpCB+BUsGZktrN8BZPmUVTHKE15ORVW5tmQw
zgmVUDXNg4m0xiR0CIdbx3FT3ldyTM4E/dzjICyjbVSKO5kjOxJCvxjSL5ojLLZR
QaXgfUMNfGuoTyAMwQIRMlIPr2TuAK+8RPv3Q2B/ftfSsloce/cX0nzQB9l0wpe2
gAtVqXTkn+s05r8JuRZakjYT+r90lbKXDP8nciETJ4im0F/nUpSwhoBwRP9qKMeR
LetuHH4E81+i4LSFQVu1UPhEUQamNQxax+c3U9CyK+K0NSKgHVU3jBcCMlr66wuJ
wzihbDxXFHBor3FC6cIS+nDl5irYObfl35NCQOlN7BlDWpB7fWkGB9n1nOtWjpe3
LR4y+feSdsdi6k5K4dGwkXXOTMwhd7oditEiHPcPmJoX+TsmMQuAzJoiDTlLDK/W
RQ+GgO4q/kS2wraCdPO9EI9O05xgN36uLO/wExam/pnOUxRNOVvLsSYtWkOiV03a
m4k+Y11qG3+fx/DIynbVwGCVwlVf1nrQshLJfvr5E6LEaINhSkr8gbteL3pngxLC
8vkbxckY+anAqpXhTwLdZJCKkUndUHnZEHWiwWidqAvqCfFTOxkA/QERLe+pZs+Q
MrKNjucHQcYrM+AiPcroWbEt0vqJSeBuvglumvQS3gQuLJrEAxtu/cilM3WmjRXc
ZBwT3SPMk7zwX0JZOuMgLTEOLttgnkUiuEh+3ZMM/QYZ2ciz1MmbWVKylxjsFfkO
kx4GhzJ5+iISECwMkRXD9Bc4qT3n9uJqcTBKXUle0cfd77G+m96sSDELeNxSNbtx
9+a7jDvI7xht6PBwsKalfKsgBps7zuXrXCXcn3o0P7yxqoiP0DeP0gUKoAYqZQA5
tAHImn0PZFKSDdXAOq/lt57nuQz6UISCxUDPH/JcluNeMCTdMKE/bIJ2x5eAWHb8
IpS/8iRi7fwTn/4oi7a01KMpOMLBIiror/ef9VfFXGc=
`protect END_PROTECTED
