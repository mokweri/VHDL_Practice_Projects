`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coX3ATSOH2o3z7TbIHdrfZ+v6BJ6n0hKtICwkH033fm7sKb4J6toJrWIK4IbkHzu
cvlw9rcPYfwI/Rfvc0H+tsdVruRegGNImsskJTAy1szREnmr/ArYTvLyRu5UWFbR
kZpIoeUpaVOBddOLv63LOz076xChqf/kMpXuqjfhqibiTR8Dp0Hw4aQ73Cak6qY5
3GHyWUSx62z3GeBRTELv/uGDnSpBKCGiF3XC+uSxNUn1OCw1DFPMvV38Mwy49MNB
71vji/orXDAvSmeLrW9INcBgQyQbaCBPpXgTo5l8h1qKeBK+XNXCV76Glriju1QS
OwJJYKk1udyUuSzcNudAjhyxJ22t0CPFkrB792vTCMwMKnklBCwmceYnIubdf6aP
HkSOxocLgMCv9ki4TNi/6MdtMVoomfqR6FuIWW+GtWu39bG8v6C/EEFFhY6LlJmO
A5aeK8LbjO5I2DULt4QsCt0zymc1oR4DGe7qj0aIyjHULerU5D5kLWSr9byXPzBg
G/Q+o43cRJQIznet8AhOyKWgh8jr2txS41/C86V3qQp0VS62LzHWRubcdxo5pT5j
eMXWVA73YFGQn2Xs16/EF+39mjaUzz2jcUnlWFglTwmOot39YIU483nsJsWOEK7J
4dtaCWpNwnbvEBglH7naalsIkYDmYWCjLF7Jyqybi5ZTNJpcRoBxPiOzwbg0x9sl
1ZoRdvgJWo0qBnheVH4m8FshUFJ0SOQgRPBRZRjunP63iH4R07y6mBgzgDvOnGib
IRPZLdiyp5rqCcZ0yzk1UGvCJ73Ri/B4TLKjFd5/1GCqHXqICmp+JxMlLlVFEkS1
Fb4ng6KwgjK4jQC+Gl0g2fUAjLhV0Zm24qIxLvhlAA2WkRLLMjUhV6ny+CTqbhSw
aAM6TcOMa5CVII9l8RmegWg4sMo8/CwWVCfYY29cV08Y4d5z2iqvENzliSV+bF3G
AsZziBXuit8XTskfc/27DtMceDZAAz9XH6HvyVp+BpRPyJa+hWAiCcRJEKI38DAd
jhlAJ2wE/vjZKMhIK0fyUyXkZAzY8KI7vzOFdj+CmSnJCilQUMcGABcbHBNOgP7X
YEzKincVii5K5WK/LUUln/PaOEoIDRRVgbiialABQNkwGMZTgGNFwJP/xf9BH8KU
gHB2spDmP3HsSdA/WgNHnSVJza3rXJMFuXS+yd9Co8EYZDnCwgjZUz3tSH2wM2gS
cmWjFL8lw7LuKfqsrFcvzY8D4u6RnQy6ifTY36SORCr/flox5ssz5kDN96j9aCsO
dN+NCCmUyp+8QMoq0FyqLf65bzqUZYg10E3fVfZzri/6UDAfR0O+u4ZBvDR23Jxy
cMj4m0E9lUF19soxxZNexDZxXBhVR9hmgY31U1UEYIsFQ88Gk7uPBxstanE9NWkf
tSkRjWJUzmLYRRuBO5AllROjfp71FROQeWGXgPJQ+cUH+20GqmROnXvMN6KfQreS
drG/7YEYqik7XueGXAoACFtXc+0rerImHRsj7CYHkYKaKJHXbagl0mKEbt+WLmzo
NbX2E3Nybm4+isKv0d+dguEa3b+ZSSm5vIQwL3lOxCCH9Fi2b5PT33MtSPY+mXmC
amyGn58mcWXDAfqSwrIgIRQcs1sC7ZE/C0q2sl/L1pRFk0cAfFhiGOKgXxjtadIY
5Mb8G0fTqCG4zglI2v5Z8u/2qOCR+ZXAc4g1cNmgFXsLc1d47/xHdg0LhjcnyEt7
OJ7ERcLgaoVTBVo1EHHjD0Eia0AhIkZwTaPYxex57P+tOelrceeaLvRcmK4F8cv1
FeK9o70iqx7hcSxk2kfTk+7rHoJBqVugr/dA19wLby8YsXDyQMn9StCDpgMK5Z4/
ounUKyZ4z3JeL/WtRd+qPmmMFYopIKnUJWAW8hEbejFF8LuDXhd4/OIi3Z9gjyLM
QnK7IGSuJDDl4mXQjGpsmHRHr9dc1eLEVeRYLW2RuuIPKJUaIOuXHMctxGLsHTtT
piNlxRmk6XIrcqEfMC0bvxjS9YlPY2xCQtO3ulgNjVTGeHW5ZfJybrxpyhAGgGnk
qPNhrTo59nQLrSVBWHdPovv+Pfq+OLMqk8xgRqRg8Euz/ukxXZdzvEGQDvX6QCBg
wfVlze0dfOsXmdzcX4rwiEK4h2sO7WEJNPEBIrZYLDEU+15SwLLDW3KtH6ZeysJU
aby0fVf4lnuGBQcpgDC0HPH06f2K0QHM898fFUZYVuWW6AwSghqXkcyBJS5Cq/1p
saNkJ2MdjHSvYu7b3EZJzhAC6bTAL84x1wPqao7BCRCgZyzEYwh/l4P5Wqtbmqo1
3fPgYayf+j0M3UlyrbVWSw7DDX6cD1KQUCHCFb5hQ4hxtyXQfu+qzGNF1mibj767
O4+CVEduVR30bNm8+4FaHvzQzH94rlzTr+DjAc/iqDk8Q0YsZIBdTukbG9Cqr3NZ
PZqstQVA/jsAKbIPnsnNlt6E0VubgWFKmHwOwJzRds23IPRU/U6ZfSAG65NyZyYD
h7vxODwicxmp4GiJh2qfLAba1DqCVjgHuhzYMTGk5IGI8HVyxt5c0yZiHfc5OPC/
8tP1fixf9XurhYWrtxGSCRHkVlTipCg0UKNUZwk1ai4FrJzFNG0TEPFflNwCbOD4
zBVBkMaKWgJ2CkTMK0rUGtilQQwKrMx5Z7d/He3szdD6HiGrjKJZ+Sc4x5huEs5M
v3GJ9bQjbSL4xYzCqPHWGcs2ZtZENlGPWVwT5FRGWEGBE74/d2wwZpbEtKu4+UoM
yDEQRLA9aVT5HEmLqsWH2A==
`protect END_PROTECTED
