`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xcO/scSDxMbESiv4JQ/lJA3zlbEpxdMSdrSRtQ/rlXL0hLawlskHhuayPNKUYBkF
Yfk1jA2CaK+4ELdXhk7ug646Cc/y58eWp2rTaF+huqEEkAxawkekjv0+N+cxNowQ
LitxA+6O7UhclIaWw2whdQlUy8ityLx48ybnTRpGCFY5d3HtKfNlf/YyJLKH/tJl
YE+HtXhFqsWtZFshYBUlQrDyu0i9ZGSpk0m2e02kLYo9QveyZOB/GgOP6w7ee1Nd
+pi8MGUc8PHJXmLesOJBrw1vmCeWymXDiqkqxdxbUObdPEsOyWJ1zRa/9pAZnh3w
MGbzeDB6hVqj9ps9or4twJh6PgzG+7uG+xDTUTS/dZty0TdPxrBcwEj+KLuTbYNS
+GcDO4MAlHbxdwSWolx1F0zjTM1Yw1TB0obz3FiScnpN+KM00HXdjBuwPqSXAGfl
`protect END_PROTECTED
