`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vxWCd0Xy790iqSMk2hdiOXl+I0ybF8uly4Dgc5eoSDADvs+tOv0vxp/Z0cLPNYzA
ZytuJqlAi4KaAJHng02mjSAhTC2EOliTUFgW7bAWiGVqP2zG7numHxVmzVxEH5dB
HgyZoZdr/uRecydpSoTbkLlnJARngSRDoSoKt96FaMxacBjxe6OfXHO4BgDyLJVc
llxD9maSz/FEagTSw5MGMulyQBC/5ggqjyHeMyXRu3QFRTW3hcDwqe4tCoiDmOTB
gBPJiPJxjOD6sbfXzTOMYZUdXIXiyGeeeLGO+u/d+/Vvs7XRf2rb6M1K3JEb4apE
MSMjLZxfIavQqTK/JiTthUwaCSminVcK9I8rEgCv2RPRpUG9IoPA+mCbUycPYutJ
891bLF2xaRBnf0fPJLMbQj/0Zb6Lu3WXalfthP1Ac14wHOVxUE6IMzumEExBRxT8
hQysuxLh6BpzIAPy9vqP8wL2PaucqcZg/aOcb7LqgFKnwy3tDFhoqgsBl0w6/Jvz
oFLM/qwtEDhUOkKtM95lSJZc+0AcSb7PDlE2kbDv7UsBQZFXkMmxK990M0oAYlIq
Yp30KL9hV8Wa3QF+CKeEiTCjy/rcUNWTOo030Epnotwu6h3JhBi0jAXpdsBaZXq5
FUUXxbVdF6V4dnCmu+n3gAWzgeu1eweSFRJ3dD+w3QTigSpjUjdr/d6BFfXhZTSl
RDGl/63J7GG+attu92Q2ltzTq6ImszhFWjSJDKhVz6tT212ap6FY1rq/Ga3CTziK
Lxz/tYUDnvn29Eg4lTqm9XLDfFIk41PTBrxBLW3RHQs1/ECxDWA+pO8GFg4WnKRB
bS14VMVjupmG2yQ2HzEFz+rRXln98UuRhs53gaX3sUJcxCBI7qQ14QpTKXMTuqvb
YadLdApLufRqAD/cWacTLoRNfgbs44U25Wob1arUBFadwH2GyKEM0ItWh56qHcCJ
CZRLaAy+TxlhvgJjNzHNP6NvfNLrwZ9tHx5rq2kBBR+vmoAjfg81egFwtFjf6Vci
uHXP9EKXQR6iEDg7D7BaoiCVsL8WWUr7u5b37ReKCFVDDgZWo6kBdK6m8fzMnrQD
2I0tHwGQ4CX7Kwqe3Y509s1PV5p57qxPJm1FPlf4yjID3h+u6nz/MDZ4NAwf9NB5
0xWimAGjccTa3IPCahFGX3uCbUs71uuNskXd7YchOo0K/zReI0xzXO5CjyDQZHOY
o0rqG5GmKzOGLXIxiRT/o31HG3HnJQ0MPV+d4dxuvNIxF2O2vjl8jsFWvkHYZGIs
VmDfNfst8sq7fzbAt2FukzG0J22EEZzhtY90GFauFtP4bZ4eNajOfPGVu4UW4jb3
6d8mSlSQqLNDCiWc19AZtz6UxXAAEYerTTr3JB/bxaUPVHqRhtg7GNEIK+9Bpzke
EGrgwOveAE2/hWSy2EJdKv4CvaRvKIGDzfMrm+7zrzESkFGKn5SX7i8l32aWe52o
Vek+5jhp1jn7XtJizW8wQebFqoZzubEJo4q0q7JueLfp0Yb2qFpchzv35p4OTX+6
CFVq3vuVDfSGXG3NjywSS9PiLdLUgtrGEpwAcESUBe//UbjuZjBMesQx/MvJJkax
yFuH+M2QER2QYNxo3wuo83qzVyaPgjoyO1z3Mcw9slo=
`protect END_PROTECTED
