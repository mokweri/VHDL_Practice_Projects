`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlqA1U2taA6+7hHb7yLGUB3IeqisvYBHAu7INalkgiG9pfNnOTJtn5auTAkykZ+O
8/VGUjKqrzqohIrLogd0CcOpWRhV7Fa9WanRDYZDv8UAwdLy98nne8x3RKoEBUzp
xJuRiMGa6IA4sCs0Idbk2glUtidrUx6KVs2vpeX1iTydFAts3RBFopzH/A1KtkAR
2IuKnA4/Sq5UAjrkaJvtqIy43hB+AKjYaU6sVb04L+28kGHx8N/vLv/T7FlP24Yt
AjhLLSLNY6XJEIPh9M6ndOY7jZUMNs9PfzYac51TSwANRCHZAAq7NDaR4tBWkaUL
nUCJIleF7IkC2lEOQhL9Pg1JxzVbzOkVy5GG6yU28vOKz22P7GljCF9WAyb9gMqA
fSJ4e8RNnenYhR8f6IdPQ1sCM3nTrWO+V+cL6R0PA/DfqfeOq3OvBAnwYRDCkAJq
QCUmKgPjJ+mEEi+22q7rNTrnnqVJvH+0LIvyA/NaUJHnwHRGEy+10CRaiD9YCGmn
k0uKfpVUYwfrUoOpL7f5jrLSvviIbZufUwRp+Ng7gZV7Z1PmEBt6qcKbjNl2/BKM
naDnFeLl0uMfGRAW9NbDbYx/mOYgAVyd6Ny2InOrDn+lMokMyg4VAtlbWPAUREVw
Jjo3NiBYegi6BXxbcf5gh3p2WRl7iZ2L77qme+NaCRfGksjxRowPicobb25YxDmh
xnQddnOoerI+naAz+vdEBNSP2fULNeVxLkgkfHbgd8O672mfy7/zlAZRn/kxTL5B
1dP81uWngsHYg9KTUpvClT3qsfrRtVi7ryCtWTyT9CPyvOekvwfCXB0S2Ie9vT40
2s4Qwie03OzIcdvVLC1ewGPzmktFVdpqrflmhM4HQvUe09A5WSIKT7KQueHFoVcE
FFGxemQzWS6ybbduz54zluneuFlm0xMveHBrYfEH0Gyc6kzy+hTBCSYSpWInB3eK
aZp5UMSLMiw00DhcysZ0af3uw8YglRaHk2dy2tGRb2TIkh3MVma9HYQ+bL2g+4oh
BXTEKWmuLZVhVt/f6beZ6yUiJq9EE9rSGhslSN6jfvD3zv8vczEVYzEXGvGe4Jol
zv4PnujlG1Tx9wACgOEfTwyKKCOTiZ1MAGJ70sQ8evv9ZPD/+1FSESqAO5fxM5jK
0y+QFnKoNtl6iTEX8VjUYyr2pcFhbN/VjUe2/H70mmOmBkEKg3lLfKyQ+RKXdXz8
IH5bKw14yktp4pdOaCk9kw==
`protect END_PROTECTED
