`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jE0daMD5pJDhluw41oAB/uUvvdZmb4mqbVQX65uU+KIHjJIIDULKcGoTfv0sxiZP
L3KmIMqrVDMviQ8fUb95wo66jsZOUGbxvG22MIiqtN/CJjoLJYoIrPIw450mXC5h
EcJfWl7VMJYNcU3vUDqiUvofBbKpb+CqJI/idaIYDdWEcINB0KxZ2a3/SgCxbfny
hoj0QHKo4/2E58ds7J2gupWcKqnH5tgGJ5RyPVTafqNLnSbNageKwdwgBh+Vzv2h
OGW3VVjmiXErWlvkmLZC0yhqu9UXprYZzzAFwSNCNXMkY7lzlUoUlBUKnvrsGCxI
KIrHISt897Yev2yWKOWYpdWd+ITNf5xMwsHxYZIZFjhAgsLFp91q8YMDlClDX+B9
+SAqhQ6+lkKPxTlHtfxtsWsJFwD4tRUpaxjOGkaTmrV1j4A/IZdxfbdVRAvPJDg5
aIgrZO3eZEI7x4x3Iz9EaqpwQhXPMgR1YjOfUEYAs9WM3wZ71JvH9VEne0MFpA1V
V+AlXLtJBDXubh8ZBdgnfcG4au3yHFJEs8EXbtwAZ6qYdNqpa0w8CqLBRmdHo35G
HNRwAfmVNXc5LTtWm4SBBaFwFcsC9AXu7+oXBMMJtMmZCjRPFiIn/QElBVHAsw+R
zTboedSxAZtSxMYBz+dAJsQu8WwQnt/YSt9uYqp/huH4cY1yh7MMcoZh81jH8b5K
/+fii0K6Me4A63ZxM/+SyqFws/O5cKA+w4PLKiMZa+PQt+1uX3FGOM97aQDGdysw
91uweTUmiMeiG7cPZhiMRQkwrXUlQGQ7GNSvTj1Gn9ELOSz1Xqi9yYbPYXjr1geE
7tZaGy9PtH5AiMfTSJESpugiF3zQUfwDqP46eUhnvjcmub0iy9TH4Y85KF5D/thW
AmLlzfotg5h7eg9IqcYcStioCftup42q24hHRXHi09NhKKzFweunoTT1P/WTiNcA
TKYlhN/nFnsx6dBk2qCJ6beREfZ7qa0erKVjVuu5pQhGxFwJHdOAk58H7iMUrt8a
nDLH2oo6AJ3aP2WtMqxExDRmXYH0fvJgu1Fu5Kyl/wASD61NlOzygeViPcKG+SM4
tzuvr2mnflu9QvyxxxA0wG0RLe++GpWIO3LY2E8ur5yKRc54vVYc+4bTe7ZjuC+A
y2yyTYrycUOXnFeG+hWIVlGSZuyZVL9YACb5g0Ca/3U0YB3nOFsoBEBt4SAHU+X2
c+owbb+ibxLgaYzdBXMiX9wzN+tOUTIjdCIBnJ2XEm3lp9OWkHWZrENyqnWDJLt3
11hJvIFnCtxW0O10HBE9gXy115jqCaHA9fQVUQspNDc3R6DBvJjTGEDsWRuIW70T
VoGXS43HASWrhji60tcwHRHGQn34gfNCz5kRB7ivFSvcxouBkVb3okl6IjOajvmx
2J+tdKmv//ogQD6eaTqkvLiLkOOMH6LLRqdvo8awtYkdoa1miTe8xXVcz008C3L3
CkDl6bA1gcPnO39873cbZ5c+DDdg+2LvZi6CcKeg6VPcudxktIX6bNKrQHKXRomN
AC80rldfedgQF6otPO38VZp5ZbXaGkFbigs0rVd/BoUxVy3DH9RA72kzlRw1CNAE
85DGVfUUaqE7RqHLpmjs0ihJ/Ge1iQC2dXTt/RQl7n0KjZ5TmEvnvCYreVj+y2re
xrw1fR2+89xj74FzENtFBsysWFPt36s1nt29YAAdJm3lDWaEiG+zjFWy3t5wbr4B
HXqWUg2mP2bSJq+cNAjJ6pIyDScmJLAjlB+Uefi8XZ6uCRg1xXvUK9N+Qz7Latm0
lVnkWZyUtY0/1eDz55PAoqWxaWPbSig2lfpJFLcROuChJd0d3jEAx/RN+6hMBmlA
prKSju+C09qizPvX3MGUmwESedUefipKPY04S8f2Ckdp+rcfNJwrnGGCPQEDKe/L
RzGcIGOoMQweFV1fdZzJa9rY47mriY4mzr2hhveLM1vxylR01Za9F+AmW/wdnYMK
VzHVHZi8l4cUVXHZ64Q3rIGuqdeFSzeLGrokMTDxo1Jd3A6t9taF2HcxvJ0bqIB/
mhU4Fy7gQDOQeLous5wK5dmee9syooAqsl/oa+MQ8vEUoZ5HmG7pYMq2u6rhrjs6
pzXwSMf1i28SBJ9+LbLoRXJchonRT2pE6HbPFW5P+4kDRPVxwyg4lp3XodX2ztOZ
bAVPfY2fnIkHpvqO6d2dosUp3YxUtXWcTGVMdPXznQR4dCpMEDIrPk3Yt4CR7nYb
lKPGy8RHk8NSZVF8PbMwJsO5E0hEKlYLb1/iaDI0b0ps1tWhXatMdPhXDHcxY9Fx
NnaZAnE1lGSB2ZF3q0dSrWPcmlFub48oSHPUsvvp6hEk5pwUrQxSNUrlJKIeZo/v
nxuN9PrUxOZjxzKEtGmWTK3khUHDuwfo3ctsO/1UIFvNZak10g6WoGtzKFTbir7l
I/ywahN2KV7VnIwfva7eWi5wTwgYctbFopDzFkV5QSmiOKYv0L44YGGaufyUopDe
TKQj11Pt5s2+noMMpQ7Mt27IxJV0rtP4qEt7cmduW9qYofPeDFY8sJCrXH4tqodP
9anfIyFTvLUrHqUf9y4GPV4izXLX/xvefHRe9WqBkFdto8B9E+22xGM3YBLwV9rp
UBGvypg5RK63JDiJJQvdD3xFU5g4HQblXK4M0L0aDXQ3t7vm08X7XCqIR3Sdr+Nj
fcZOZjo4qUv/fXPVz9xEi3KzEka3BPvOLjy+WHW0IsQQf+zo0ir5R7e+s6ehVaZ+
A9C3qkHEROWMc8EGigrvvj03PtQYUif4FBLlWRsj9Qt/u9E7TH1jIWq/QrteGAxH
zN8IQpU0ZjtuUexSy+9iCWDFHIyaWgzILCLYg1lp2iLqM9NfWPa1zZYxz0MVKFM3
u47MX3mgQNRyHdM7BrvJ49fmoIIhn7leMyFljHKR7vm0lZOl7zZGP3yOwBGo9Qya
YrpqKCE45Ur08qogisv07Lg+zJSepzpXS7v2fuq1PW7B1c1sL2CN4sotgXGHZjuS
9r5I3QxcYfagCi9XPzpZRLSI/Ehhk44ZaDWYmqJjocnzyQx3goifFzxGEFR+bWda
KngLsXORAT+zxajGwOku9A9y7ZXPIdkU+UjB69mKQZmr9Y2PcpaaCHGskhOIQtXQ
eo9jY+GD2J8rQRvXcSJxqQCWPpYaIgp2Jx3pdGcssFI2F3DbkK19DkAL1XhFAD9Q
XHEWEJ7cteGQSmuYJDMXFw0dwOI4u9+OWZps9ZPZR4HnQR/rqRzE2sAbX5lemyXb
s1zzyZLbcSu9mEF52Oa+g/ClriZ3uwuWAY8h3B10ZZrVvVkd+S1NvuEXUd6Yi+tN
+sH3U6scvpeG+a7OB2Hs1gFoZ4O5R4Wzqg2TNMIN/YMzNVxJNCMTdwAgQoXE6LYd
lha/aZqjBaXToz8iRJJBEhI1OA4VG9phF/1MPRI0/ki5fMv8ypFqMZSJF8mg3TRc
bsEKoyqRW+lENvm2h6HMBY1t1P7zNprX/yjYjiib53ghrJHPlX5w8bH3YEFW/pf8
9u+8CJABXoDuiIS4JyyCA2iIXYWc9GI6L518MDzmsOxlqlM3d71ckbPsFfrub+ve
Z71SpOXAk2cevK2MvGZDza7zkx1EkSmnP6vL3lauMgbib+xummvFmgk9mIj14SqS
RYMl0MG48njMEtVMsc96UtfDwcG08bQ8COL5/P9jS11k9mx4yKqdxb87ZykyuwLl
XqOelIw7qDyE2WW6bbDEisKzadRaTcPpEj1vxSnyNIbAPX11EN3JYOZR9IVdod0N
xVFFA7vXQU34O4T19slEaMYel8Ls3TRCO+0S8is/RvfUfF35W/fa9NOMd8DJtQHR
F9P2JwHz06OCLSoqkeEWUnNyWKhDzJNvsQImr61/RBxyaeh2vQ4xOMwDOHg2Duvk
rpTs41fx/F/+s1ERzy/pG7pSSdGmg7nPeTtgVlV6NHb8LI8D1l48ltLoVFNwhfNI
m9hHSqALb4D7qXGqtfhTWMJOKlsOXOHUnEpm63P9M47rPy62mguO1VbPVtgLSMtm
NnEnWSFKx/p1HiqQeulOSwQIxRweg4Pp2whFR8BfWGLedhxJldFB2xA4IyBFgItE
0q/5ew7cA3yvJsFGOYvSnXrIIuMJzN5AhAVu1zMhTBHHk5kQQUVW6PKMOQuiEFh+
F4mwtdcsIuGfAzdSd2KDEVrEhEjNVm3ajj4KBer1zpRVJ9P9hMxeL6L/GoACdYCj
NqXSRKDI5Y12hF57i8h9PWrdJadlPNBESEQz6wc2vjGrTHeW4v18U1VKAcNMYDW9
6WElYOIylHH6GOPcfviBgutviCew+wVKRsCwKkl1Z7EYGbDyb2s5UEfu5FIRZ533
JCHkNIeAP1cgL5a+4WIKJjImwMKCK5X4LQ4ncEnplhcoZYXuGnrJ2+2Yf1qpg7Ge
IZxv6W8uz80GP9iTYfHZgUD1rapPPzfltTIQMvbl7sQ+mfwaq9PvSZsGpWOWwU3J
jo+Ae5n4VCuKw+GVpWCk/I+UCsHRJFZVQlKKiAZ0MHjd1ywsce15CCg1jYC777/W
5z5gIjMH4XmJPkTvJvU0Aw==
`protect END_PROTECTED
