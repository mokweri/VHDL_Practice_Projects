`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGleRIUc4iNlocOitEMAufZat5G2vmlSJAsb9Vz8eqQlaGj0zOSGoSKGOTbc9sP+
2HBQDBJSc5dR0LCN0qykGip9RanPZZgtYsKvo75LV8jRjzJYE5Jufi9rvL7GmmIA
gKhCa6NiqRh80OR0ABRyu04/S+0nlqTUBksUKAw40mdAjdulh/dYXsn9yK/GeaWE
WSdGk4lHLpWFAzcx/Ixp37JWkMdD1MpH+NVncGzaLOogrfXSRdJMziaTq5T9j0F0
KLmoiUuPx8poZ/K9mllGrpLk9d20SjNBQDe/7wsfqIR2/QtpP0xeAZejV66meREt
LqQs7CPvA5ERrEKpnK+mncWQeaU6baywr8Cc3sOTZHpfzg+N/328CX/eBw9ReXUS
+ezbmgTNQpUUsoXnwA2HlYOYU6Lh3ppr7L5kB5XKw9XqQ4wXpw1jr3piIJnuTWmd
jx+h3556PC0ImokOfh/jsbPZWQDsMAJlBTqI4RD+mbwZ8Pub67tSwrL2bB4CLU+i
n2x8DHucwDbc0NapioGYzzskG8BIaBVI5HZlKfAWHEk9NwnBrtGrDzLIwXJhEohS
sLAmxLND5ccyY9v9ltNfQhCRisftoajRPJ2ClzU9dz9wmMxJxG4gf5ToNSrMyyDO
CsaIIsQ4fPCYfRW4TgNgru0ylaBu06B4XqqpUwNaxoEukWjjIS+iZUs7Pw6T8vZV
UVxCcMOWrunb2lfqpg1s/zh2m2dQTNRzpFNdPyPUs727wvcq3CefTHLDAV7cbTo4
oFN/5LSRszDzimm3AKqvIalj/OAs4k9imy7trmGCSxHiixxDxohCZ8ubQDwSjmWZ
APXyxZi191JUW6joNaOMi0kdql9wJ+8NmqFqxBlMnYH1ya703evnUcmAYMpQTYxr
2QGxsEH0J3SEXlDyPj+dM4zI5OOfPEfly65v7+crhs9uDRcLsCdEVIidfHL6aNce
svb5hvNmT9dhf1yS93Sqf6KTkzva4kugHB51a+fzX1IMGzyJja/KybMa+Kug2cZz
cXDsG+A08illUWkT1MHzbdBzKXaAXsjgEKtB7taYBRFmSOUhqGZqCNu+d87qF774
nwAROZWO1NPjWa6bC8qUj81k6vD1Xl2jf4T+DLWuCvhLCF1peMri3IFAHYEazFsM
LtmeIh3muVEQj1SG7BK+MS8qLzwlrC/bI0G+0eg3od3tfn6YHC8e5pDhlRw+i8ke
xnSq9FWnSyEX4P0m34z/niCsk9o79oDJLgqqssN46SH9dayLbbnwbXyu7N0JygHQ
356qNPNdci077Ausn1yCGluatkmH5hTDSgYXAjA/naikY1yX9wGN5WDloRHx553W
1KRq5DFVlf/LZNprht6c6KpDwnUFLTYQ9UCHci6M5pZko7XmdCgTjBBoqFf1+X5V
ZA9fV4IhFRdg6DtJO2g+L7KuN6+tpZTLQbvpudzVbernpD86sCmCOmdnRkG+cHyN
pRwyR4JDBNRqhu5SiM2hTLSns4Ctyy2T79+oyIv0zxUwECuOnx29zGBbzJ/R64lo
Vzr+GoJcZCMBQ/6RRBo8g15CwV2OgaUsqfbP7DgQBVL3dHb5wLbbCO4HlJD+NF7P
fljs4RRdlq/f2DUQttJsFge0PeUw62DpXkJez0GH1ECf/6oZWfBnWTKgDj1vCTv7
0BEuqE9Fm4AVI7hpgDteYHQEP/KqZiR1610wIdNG7d7Eq0xI8rFKYIK2LpNkxP0y
WNI3TxN0ZTI226Er6rpere7r5vfsmNj+L14HVBj9JJhURrDvHTySYfsTviIkP2Kn
P3upX3fD2JFRiWN9N4q9AhtyxRyFNq+nnExqHRrmGvr2Xg1juEdvcrLOg1yDC+1u
6GZLmRfHCuWfFaWUjyVbewtEA1lxN+013cdoYDvYgagjwnG/+uE8v/5WtKx70eSL
ixkUxiJ8ElzJON8ySj8O2ewFY7huzSldvEarHg9u0jtIVrSW2bQx1h15eUwD7mSx
dy0JLJbVoTmPXfTqoN0zuur4yXR9qUILGHYlGSSbGrjdPEXQTggZOuzmrLOeWR9n
ZIg8QKS98dNz4Ii6Lpyj+E9QLcRYpnFVRo7GxvBufJjuDZFbwXG6ef65er2u97PS
JyQgaw+S8CvPH5zjmlFTBCnzD981Qeg+Uo/7WdGeX8HvvJkNGNA0S2+YicJDA64m
AlonkzvGnuQWtqfX9wUFahaRNWxjyJ7j1hhcFlaVVtO3qWcnZO15r780/WSrw/82
zjlZEg9OfRRKvURDq9vL/HB8b0eJDJkTjVQgkCslsSpVz5a1RUH1KH1QXaBWzxkc
/x2IP1j/tFiHCqGWWy/AeGkZoDzNFVwSK5J5qVdNExCUkr/CgGp5YWB3iC+qhIBH
0wZEFy7MazCsjk/ANR2kZH5ahie/wqPp8VM4DrpvNnPYkWMtGtprHFG3m8aLfvU7
N3yu8/4MwuUf3aKRY5J8WrL4lWp+f17jGGBbEfTpSDXgGJ+2UCC3AxKKRa2vwcOF
CjlCgzMYzDBSc1iRD5iG2+0c1to6C7QK2FEUu3fpC3t7cpMXRnb2snsG6D3Iw+Xy
xJgtm63Q1YlM8t8J+bmqX4j+fTtohdhjs+Tl5CE4ASGFwF72XYWzAzPm0QGY/iFS
Jc39NnkPKNdMzuayC8vNN0l1daUKzW0lE0GhwIeUYwCT5vByhBtIBbketwAoK67o
gtQcCDMW8km/4UX6uKcdDsSbCAxJsy2EXjiMl67NF1N6tRFfmwoMpbnRNU+/ATbH
+fRF8mrnVJlBGHvLeT6DmTDMSDW269fOnszp2U+e78/Vqp99OgUuXZHiUMVFWkEi
EqukK0tkd4jJ5b6NixWHmfVwwz/fJey53TRPpedJ+D7pRR2x+UTj/uo2COyIA3W5
g2De0HVaB6/O+Tkf296F+q3Des9RIadOoYaRo5R1d7k1q5wLFq2HIA9V1VAADPsm
MAsnhKWC3vCgEQAXFcBX+iFYyTqhlrOYOoAFh/ANYGvotb65eb4mcfiGyMq5/c3U
ktjPEfB7IMnnOBqbIdIo8mz0VmmsFfD9y7r52igkH8+iT2ww8E8hjr+GjQMxPuiv
W26gkGzFpj+aO5jddiQgMKYL/M/r0milspwFlj6qpbZf2giZ3W+z+dkcXIDy4R66
0t5OBiSLTUwvvKUz+ou425CEAkcAxrQF4Ov+D9vIqIGd2nhuQR6yjmbXsdCAplTa
3oGU4j0R+EbkgHnZXunzZVCoUVVeOXALqKW/oO0WbwZwZX+HnmKiTWo/79CGymEV
mKoDgUtKkjyhoAyk4xcNmqTYSb2Qtzy6BESPoFceDtwH65JjJk4dKxy4mfcQLW6q
n1Z5Gfris3AK++jO2NnoIBXdXWnFtymC4cTZayMqiwSs3wPNWJzCGOUP/isDsXBU
FkqchRCTYZlARyh+LSVGIyNbDBnJdHfalxlqG6UtBL4FVE/NxV1gfiBajB5qcd4l
9OHmHgqPqW3T0pRKZ8Tvr0fjzxmO6ipdzLk01Tsd4VJH/BZFQmtglm2lZjJzoMxP
+lWCLxk9CFZPhM7hZiLQCBDqb+ndP9049dgnu8Zcm0bHtS3FtZc1qPxKsyyqByk7
miQzNY38winuT3H56qP9IIbisyRpqGnpnqc1QHH1Xd0TgtxGEOPJcrEIXxb5IYsc
1ueHgRsDPb8wMI7MMj1+jwqscvDLKtI0k1a5ZdqfOlp2eyaVb7Q01+cXB8Y+Dqf3
Y0ypZCga3ecb8pxxa72Tod85/41zZ5bYz6kPl1rbkMsjbuAX1jcIl5jbHlIPtFFh
kIHQcnObrpWLCBamzXLswksFdi0sOJCpAMpcr0FY0viA9A1hDjCqWBm3RngvKc+Q
kr1zQmPaR/gaHYTrBVEaPfbaY8bGv6kt4vn38yYf/HSA09aF8jp1WLWV+CDTxIIn
58QNURBiAMjVvMw2/+REUKh/BKmUoFZCPV6tpSSWAwHdtgPBfPOJG5rwSgXxBphS
7P1NP/nuGtKyz5PrvDXDk6eDLrW5lfekJeHR9IBOece2xZjaPpVF4mhWjziHABhZ
FBpTqV1QbyjAEWFH7L5RWDb+3AFZu8bpTniqNSo5yI0kbyoj6D8kNr0rn2zxwvpJ
MiwMQ+4SFV8NGvxtRszAn9rVLw3qoafBNhGSK+iF+ct+T03kjengUEsGWeIaTdwQ
Iq1/ccUUXhZUx5Ch7Nhj9ufbRMPBoRkJyjGdl86sve7JICVZ717OFTWetoNNg4CX
WkV7NTef9iXYu/p/cSniGvmKwnD34keGsPMXd8hjWtGAeiffDFJb4+gDRcCi0K4P
Py+HTD2nq3pLx6TbUYWpsM3WS/jQVG0iW0fBfrNk1BR5ykRwCTCkLVY85Zaoeu1p
1wACO9vcbyiplyeLMMB2izN/ZC4K4dXxX0CvhJEb4kvp5SkgYR2sc1ESZaDNLcdW
fSie1QcV1siB+DZsgRGQcVyyEEV4KMBUBcZ5tpE+WgW03nsyyf4hDP3oBSugpmF1
OVuxfr9zt0V1O3QgLUSFMhTI/BQwHOSQXddw0YwYsxb/eBDbjneHmI4bkmkSgyCU
Qv0GCeUV6NQSip/C+oAhs/2O7WGQwfU2EafjD0O9eOht0/pZFoTc3s996PDOyL50
LAzaWxNHhLFpmmfZSic0BQ5ViZJmTGK6p/PeWThFaYRW1Z+TVH2dfpbC6uff2eDT
buv2yBJ9ZhRLmGa7qGjGCldMmYwhBdy/A9lVC7KPGcIpgOMtc9Pd3JNxlN/8lLmP
Rw0/c+AGK00PqWjWggNHmMlgPw5A+cwQ3dgbF3C5DaUOam+HswJkf5R/2uflhkNi
1biObNFAxstoNZOUgeGijL3n6rWGhUql+jTdNiYq8iiUFQgfYgr6YY9WLALHBtok
MNsghZVVUWSw4WZiXuLUH74C2fADgnNkdBIf+pCovgnz5CWgAP2Rj00+v4ndsWS7
tnWFupUNckb42YOG6gtCapQVByRdzEp3gYQZiw+sjA7LMvh8kMIDMXpzxt2be2CC
ZQMs7sNdAFs1bYHJ5wFAr1Esexgv3ZN4UzzLK4CRA5Bw+iUFpJtwcauEJGkhH/kW
mLG3xD33hdd/HjZjwz7mCQ==
`protect END_PROTECTED
