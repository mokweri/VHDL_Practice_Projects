`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O++T7o9GEP75HWo+2gxsiEA6wwnc7OAKA3I4dBpp62NPXuDrVi+85u0OwlyH/htL
6FyDBDR1pgIvrT+WkMvqz8wVZ92ixW+Zj4/uJ17oi1j5naA+9GJ9gb4RDIM+G5yS
88HY9AcravC3pCuv8wf4G2Bl2/m3xMY4AXSztvmauXfB1FP3Qmk5VOovKfEF93C1
5Yg+4SWKX2vdcFC+AWyETdr+Wxl8xI009IfjAr2QvZTzPXNQtdhDxf76U/4EyFXQ
WM7p5lk+15MFWNed/HCsU5iorneCV9nLfUgpFEhBuWZNNV41vaYewAWZZ3j/r+Fl
urNLIOG3lr43f8lZ70KwRzh9ny5Q/FKcde4B25Fwn0WyF4FIHR91yJ+AQ/z6RJZL
/iiMKPTV2tQBDZ4CqhmhSIrRV/KAo3MsNxh+il45excMbMZ4VFpudMCHk+lrVF+W
AwZMfcBgkWXXz44DUjsFVeOj2EomrvoAeC5D+MVHdwDqWujJZ/mkUdz+UPfWyFAM
WJEEd8HQy+iwgWL6Rk3GnOyO0/TGALw91NPi7q15IvEHd0U+ndPbNDcSxVd9Wu27
bxKQQ2wRySqqIkhml1if6k4srErGyJNZQuzVIDwaekxCus69j6jiWYKrtHs/6/Tm
PuZjwoLXNhcveXTzPssvJmuwLKuQfQ/tbIDFcr0g21omXjCBLqN/s617SFfLTW0g
l41m7ubzB3zHeI6v/3USNL8i8tSDU3LHk5VdqucXe1Xd9nQ4aXWB//DPdQu/QDtI
iqtgV2TV5aFTveFYY33Kh9N/c8xSgO6/vny64ePi7twPuSi0ZXucZoYtkzeyDhMv
fiZ0OmrcVO+l3rl8VSXArAXoeG+DLnQJA/DCIyYx7sP/UwSKSwpfm7esuNC9n8Js
M/j17uy0GasKIlnvWT6obMrqguylQ6CeinOLQrZghKp6pdkX0kOSgQlon9SP3UKp
`protect END_PROTECTED
