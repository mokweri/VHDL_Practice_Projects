`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqzWnOLCdYnfQeixDl/aAUdW8Ae1GYJNCGMOxqIzob6EEAhdN2QCI2T0m13JC7/G
gfJac04ZYush65ClnBxEASv+OHwlh2zYj9/gZgES74deMnKiFFvhw2fdHAHzVGTs
oNowgb4+KPsnU90anhhhlklrzHhFU2CMKXTZX46Z0ieb3mbucwxpMlw4dyBrBeMA
YtFkAe0UrXdLqWc0dli/Z5Sqitjwo4OoYsrUPDjuaKKixZNGjCw6yFWPOIu+/AYz
ZLeQtXXA2Dp9ORRsk6OJIa548cN4A6G4uQRxA3OqEF3rLLIqEUlJ/j9Jh7chU+o/
tq4SL65sBY0A4PBtjoT+yTcdsqQpWV8Qv4WcWHgr0+PTr0vfq6VIJIMz3fX9djf9
1q9pYBcuP5PW+FLEhKdsnl2KrrlLHx7LtW40asc8GhOfg4wlSA788TN1N7fjf3mq
gr+ZrRlRqflww0mJ6t2VmRDKVqS3CCgn0yrRXkBhqNp/v0q1hvLxDzfsM3VbPBeA
qlG4l1d5sX9WyE+05E6AqEMg3d3cZIx7N+8qWM0FCBzDWcZ+MAwebIgApa4Bbw4M
Z8GvNvQbz6mSBrDjrZuAr6U4KAUuGbjKd4zjJTE/VHAIeoFNyHzvo+6UvX18/uGj
TG0SLkcG4cLKlYfAYnbKa0/oJ3AQxn0InhSp8vMS96/lezin3rjIyy6FnkPp6BVG
/heAx6ZjE52Lu+WRVkY8ow==
`protect END_PROTECTED
