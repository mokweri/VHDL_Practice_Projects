`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VG8JuZiwd7X3Z6u05/r2tZ5+XXJJe6hOTTZatIRIscQdsQi8p1ulYc1SjstMM4vF
lianQuQr2re15g6DifOiq+n7x+a6xSDPKEoneTX4HLHf7KRt2J1u9wgPsjH66gz1
0wRjt1seRiHoVYj7wJrVRdXmx7D6+kUsVtdtbo4kM38FHCJV01zMm/gKY21kvzJD
3tJO6/Fa68RQBjRRzBdRKj5k2qyIh1tQtTVKXqPQubw30y3cFTJ2pChsyjlrOgbr
H0VA/1OW9SU5hAhVyY9BZp3QiC5WuAH5uO3zVXjhdAwtbLt2yqsKABm1mgSejmUX
SJd2bmEbkTh/QnYihs04kXii/V/p0CHByB7yXCSmmFguno/8B76SP4yUCMeKS7HR
VQIhaDTjnWIMlKh6ckRfouc+e63NL/R0frI3sjwR8j6nA8oRo8WeJXQMuz5OciRD
EUz/ONBiB9XhvyaXoxcolCUouMziS3lQkb1DjMqMP78VGdbJmF57uvqn4ZdorxF+
7hB93OMKI1TKoUDgzbGYT544uRUKcPOey6wcyMBMF13r2+kajOdAUycsSatkPp61
Oa+GXc5SOr9CgsruuKxu8kFr570oue0syU57QFgDKpHuGhNQuzmC4pfRLmLDPIBn
BUaoHWv0fmqQegqK2aC5P/+Su8P0RuIMXr9Q39yNlXIpDGw4dDGgzpsBVlMnJCdo
TBqdBOkid40o63Et4kd770QOakF8peNdkfPw3zGJSF7H08tPG3JKcbpDDZMuE6dk
mX3/N1QJPTTWj5OQoI+4gQhZcMe5ICfFSOeTh8BQsnmUW9pBgDksWpp4aZqTMEuj
Xnloul4H9MdTqH2gCEK4RHEE9Sa5lqgtbDovQRuCIqMQQ3NM/zWlXNlyuW076CQs
cOxFkoa1M4/l6Eyo58J2qHi7MTu19thUKcCnMgo/pyQv02MiS+TZVMg5Tn0vxR2k
wOrJstl/HV2IGNjhx+M3onfHYqp1tGOBEshL6PFoHzo4jAoeA3zJSFoqPYfQ2XE+
c4pdTRc6sL07Qw+poTLeq1NpT/rC5Jb/LIJL6pM0tZnCp8aTALq7o+L377q2nFdR
fZF1typqVAqGHNPcv9jz8OuPHpp11k/pbTbF3tzrDl8WPLaLmTYW/cv2W1VGjh2r
22wPCYA3QZGEhY4vJ8q1iHMnsOqzF2pdhYx3fams5yjaUxqwG9qSikng+mhURpLJ
2Yt64vQrPNMnRCNiYQd8qQzSoYS/2czalwuCLVyZWvqDr+XlBwWRonHHPWw7H+zF
lvRC/jux7DraM/RgpY1jZCkLyBAU6myXeWfm4FH65gGz634v/jrBpV3KXPqvWGcj
Y2Msu5c5ALPEhN35YvaV0O6Dfw+FjRwqwcNGdbxCeYLwzSC8IqvTlpSCMnSbUN41
Ya2G72RLUZR5g/ZwYXmgMXXzF/hSta6Szcj3fXASKPyv+XuhzFDVAR/2H4Zgnrnc
FgzWW75GNT8BREpF0zE8nDHAwcaew/tywIpZdDwaHoKXMJdupULZwQFCZRHXbbEN
EnAiWlUmnNnwLg29KyaFRUVCDy7JqkHiV7IIAUThUzq9r1O8rmtX0IEAtg1QlqY+
J9bQOb7kWLc7c8LCsrprQThQOM9gFJ94H4sxZ65wn9mUKPU2XMjjhh9r2hTZl71k
r97gQKLZI+E/2fL/COC24g9lQo6HX8c2BGSpqQg/1ObyDWz4Dt9I5Tr+CJpoEjPf
FLewZvQJKp0KiURZbbFkWJ+aFmnV5zWc/ypLCQG8SKSE6KIG7k79PkVB6MXX7J8K
AV8SCzYTQWtKRZ0iJSOdnECSZ/eBq4H7MZ3EJZngaYqg5y+gJ5tcSsmiaS3sF/If
X+lqaQy+Gxdl5Ho5woS+JaIp/S4SfFjONnMgGxYufzkGZTlh8XX4h0R3zWPCoHjW
058cZazIl4OFuRpRWHi99A==
`protect END_PROTECTED
