`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1dA7Ri8ykrJciyoFt1LoCogOKUjFKyzzuJt6g8QjshZPBoHrPnJFPPrPdubeTlzE
YkSBKjlk4IvU60Ed+6mdsjW/lWWRRuYTOqHEsVH/xeLe7HRXab73Et+VIArkpmYF
FcLVewrnh1Va1YgLbZDNF/B64kRkIAP1Z6ewfgzgtycXcW8JAT4u5uVPbOa5g9df
ZJceUW4qwhdB8fLeiY/8HeACOL5Zv2zKh3Edy1MI0NtLQ/8AE/9gOUMLKiSHNCv3
HeXBRqXz6f2F/npRnLBw5qt7tARXyJezd7SV0osRZKZbZL9ogE/8lyiqQQBwz5RW
0z0gZePOAZDf3wADr/J4NfCVvUYOmutMiflwp3JmAN2PU9zA6TtLL69j3pr6IbEf
a0Jl2F8NGVSJWOYyhvJPWP7NAXgD0Uelqm2FD2PiTDPQlhrMdki+1ks/UXX1/d6j
oJIGZCL7PRNtrQZnVJj15kTVDFjx1sdxoO+jZKMTWLOg6s4+tme5NabamuIDq0UW
NYyt6Ubp7dDvsL5bLfCmMJ5XCLmPd49Z2e6sqUk2MX/VzV/sHdOErtEGLQshFBA0
mxvOy53XrcNYwNh0y6cjKhAmpa1r58wN298wKUMMvK/Bj8347VJh0IBISjXFbhRt
9//E+aa+qFeJVm1TPxvWITU+w5Ct0QAbYrB0XKOat7t0542rJORunoXR3VbDQK7B
CQqo4hsoiry5X4P8HoCjvRdK3W790VEnuHB+FFsqiBOk/lDhpgcANpgwb1Sg2wih
Jen2IQUzmo/1PsSsY4g/d0vDvkZvzUBkFD8bX9XLNCG2Aj3fycbjzwNeLhMBOZzD
++N6wKIPQbp2pHjkJZ4yv8t7HgwF1/3+R4lxbHmnyWIfJHsnmng9t7J7AmB/VTGy
BxUUFhDmghfsnYSz3mpI04oLMLQMjk3jsP/wYtJUXeNN4n8B8d51dAQkySRFzCyR
oFJ1wQeun8JdUCdV+g+0tMlKVyhA2qeU40+LgtLSC/WKIaZYvpvG7160zdn4Krfl
g2N6lgjpKkwMnAY6s5xdMduVO5Upj2AIYwAVOoWYqXzzSumXwn2zBgVTjOTF9xt5
G8f2zTicAKKtDDfqZ+5ntqMYziYhwZMmYlFonmsT+NOtQyCq7upGujnqy+VKh6Wi
cO+Bpo4N8ywVFT6/IZEcMXPjr6muCb4YR5Ih2wcJEo/FcWzbNfRWELlNLZzNwGQk
x69V0Sg+NZkR3zz/pV0IDYqNJFcl8Uo0MLH0XfN/RPUH/pKgGGtNhI2pwGChHwQX
No62+8antsPqD/O7J1pAPWcUZO2YIRnCZtMs4dil6H+6WCtXz6f6uh6Wxm/508O1
+Qc4eshCS4eeQmczkx92atb7fD8E0zDaZ56m0PNQuNaLf3aUYv7z7Orye1eDka59
GDOLJ7kUuxY4x08YR+SjpMEWRqIfMhA5iD1Q2cBvE7C0FOFqpAx+uNx4gi8tOsqJ
JHCMPTVJTG0BsftQcraQKntZHzhwuAD9wwbbPyXB0m1ki5QIj+jhVWOhfy7l8sXK
JSPXUqXz1JFIsME9fFJnKWYEzgSjwbe7YroV88z/SOzPJJglFOwwzqXxfeYFFVYj
0mRI3A/uPplC5XVCZFFi4y5jPR2SWtRrSXWIRVFBqSqYIGqBmn7UWI0p5AkZnndg
BAT28+xLsERefiQqM3LPd6IyH1LUa+0OLDhxWXR9nu6LS8/2+8f+DWzA1fKB6MG3
eFCnfl6VxAuN4H4nJKDYJOVYFoTSbC5jckerw/1Ej7WSclyh32QeFjdqOpey/t1P
va5vpsbBV9PskG97zvBKj1Rr3JBT477kFudbjQJYA7x/3/AJe1jMQqrC8i5aqh0l
KRdIDXJhCDvKfg4MFNJN8XSjx1zyswcsM7HsviUzMdHWgXSnVXbVP7wCoth5iv0M
BOZWlnGmCWhPDQJl3gBTBIpYvr9AUdkOTX6Xejvr0jQw6GjrNpeX4CMheMuYR4Ug
U7RBzasmUGhWIrsNNuloyRljYpM56+LKtZkCagkh3fDqlICtl/DNY60nULvYJI5q
U2JBFj5+dxnDMFw0QAUjgcaOT8kGJpfCrgK952A9wrhn5k5RmHs0PEhdi1EPzPDo
To66MkBDgEjKDNyppTMdKeS4bFtOIe7VvOjYBGh3xhpsydULCXSu/B/fVUhEU9QX
BLJPJNKrOf8BoRqyZ7wlU4FBQ+JQpe15UgNexEY0HuywA+sj9h6sGDtgzCwIRIUY
fz4ggt+5RepSZwmoYiNQSOlPTSnMbKHAADphPUFMZyh0IhQ5Qv4MK6rZJi5o9f2v
lIlbwFq8FVYlRpJJYIRnjG64VyXxVJJ+QH1lTvA9iWnmiU1MDRSu/nwav82R7Ate
qLj6CHimHQfB4R1b+EXI1LaDat9h6JWS9S+rRsRAD4+masY/4xbmxNECAljJF57a
W05o94Rk9Fc37+ZygJWHhK9Xtzwxc2lbnqicxpzy7pP4h4MnuABahtBZ0HpXfVSa
5NUL+JSAjlCQXG1ixCzpLJWrtis06B5xGh3kb5AesGxivlnevhid1GfDmWvR6liv
UrC1NmvjEGN69MdTlZDFWFb6UMRtSYzErxOMloh6b38vVhq8XkThpU6UIy6R4A+r
5QqhVaTB2gNrBqhue4QsSPVD8iC4uOA3aj9aQ3f5xlLgyq5rJ1K77PUXjVovVHVs
U3UXi5KVn5wJMpxJAzLagiJofRVpL4gsFFTy9zdlL5O+GpCmgXaQObWT6eRCQME/
a4ac59BJos28egV/dLWInWHHKW0gXRDoOl8qfykdipqeTrfJFICzvPq7o84/CtQa
0kstaz0M1ZOdeOwALObTmMCwSTt75lo2NKYM04sCp+Y433oTlbREASrsZG8q8Bnj
16MYIZqY9WLJAAX6on8t/nDj1v1c+8uucEZ0F71WJfNDsu4diGAlY5OXtnuwvkMJ
7qlc7E0tH+AMzxl5jDxfJ7IHeOZpHkMNkgBWlB0Ga7L9Iku7TBjH7jLk3n8NzrVS
q5oNXSGeZwE0MaXqVyy2/RGSNKUPfIXnqABUpGLNIT+v0XgfjDImPqZG+H/dr5Yq
/4zjnKQXSRVVF2UI7SYqW+S+xP1w4A6BIoyx6nFTQd6ckVoCLqUh0KyMXE/ylsFM
LyJ4JKG/ZYU6x0QLPKslzRH3aYjjVpcbkSFSIufqVOxwOoBzsef0BFcBd508lNSA
siUdT8mFSSr/8Egoj8pYbJn0F9RYnZ0YdW28+clVkZmqAsihf5AjAuFpGVB8UhZC
eFzgVH0zGJK5XVMxjMgmAQBxgBKylrmNYag13mKRYU+z43506kspWoJH8P6uOxBi
v8YUoPagW8tyssCZC3/LkD1ODNhhyHrG0KJjU8n2ETN72U+UNbRoUDxtkZjKHdJZ
t/F+mpIu/nn8YluNTBTVPNbH6+FRptzZHXCi2kKNXuh6x27CjkLWLCrHVZeuLeu+
yjFQAe7qoyAVK3rlzZMKqbC++7lhCEbzfGEo24fnUIPlszFx63nMF5ZDEhUVapHI
7zWe7PoDOTtJbWczP5i+zywVizx/tp8HGospfYgtGA2FW6/qURZo1wZ8K/TisuXm
xMZbZjWW+h0wS6Df5hynvlBYjHlvNLDAQaWrhCjfaKXq7Tz9DjQAxjslQYOkpFBx
s51HdozjTwNFuqaiazRkle8MdpHXSzc5GyW/+jz9woa6JExLOV2XLQv6kSzrn0Mj
a78JuJq4mPS5egrssisgz6NaOpXPiObTQoLH9bRIpd8+ZCi7ZvkYc9ZFrDHD2o0l
VkWlizz2OvSQ5o7uIoB20ZTMU0W95epX4wrb0p4Odhjd0AyXddX4CM9NhJRlIqHd
JcFjy/KZSIpGqjTJCFMFR5DX2f9TbYJpqBBI63Z/Vtzmf5ArS2gO2KamBnTnkezo
49nFMIDnr5jLEE7HRsTAH+DEo1o4YEEyHkVYT97gKDZ9YPNF+AqpLG7sD3aKyewk
NdlGFOaD4UBbrJdCZfd7+BqpgNOeYsgUkgh3MeFcDPHxkx6HWrj5XIF1cYBpQWdU
aKVq4E6a6CpRRORM8yvDayG9IGxPP47drnQ50WSFMQPjTB0mvehaFFbD2vxsw6jq
vjS/V5RxN1XYwh/XII0qOoC64/L7mXZBaAIBIWUhQejyoxdNnD17nQ6fDci1RWV4
k42c5zdAtRLqxYze4JBGgxc2PblPaG+2uoIdvIaZKdyP1ZWT0PVASLOxmZHx1iSU
5jr/TLCLkHTbaujBa8sB7fjFmrpLLPpHJvqRiCmPyOaqwG5Ky1DTJteLZotZYpQc
2LMr+frqoVR4fvP6avwvRqNcF10v+TgRhqTK/SU6xyAPG/H5ZrwzYY5lxrlVwJqy
DGOvGTlzusnA5qPpdbY2uvIePkKEuER+T3aciEtzUqBiOGje6SCiGtaXTXus26z3
E34STo4joXTslJkXY5lH1pmK6zJDUPNtu2Gu7e/1CqmbML82vo8fKEdVk/4LYXJg
l7WXMxeqvJldt0kl4pgCtakDp+6J+YJyrOKjH1MjXSDJU2fSznhAzc31cPWLNcTD
4aXYfBAuPbL/W79xUc+BOcrGrjkaFSIq4PhwejFP+oleuqKOwrht5d9SnnJ8R7pg
C+3Du8NQT/j/KQljd0+YGrK7UvCjPaPqEPE/fyIpvGjd5qTsAjcqlAIeiPImB3Z0
lpI0HLNuyCpAYOO6Tsh4twW4ghAhYCU8Ox8CsNBxL5pQhcd12qKwAenCuUgsDvZA
k/bhiWNvEVncScAqSTdeTRdZijKaNqYFASsfYyFi8IksCCSmBpGunKu1yq2oAZHZ
t4SRXA9ZZhd2KbmJfHxUMWxEIpTfuuOohMBgzh2CAiTTjeNaDJshioJlYZYYEuO2
A+mgoRN1EZD6xVF2mIUfaWkZRpkZpBQSF91fOXmPxSZ4jrSrSAYWHXV5gkKdjjHv
KIld9OujIPw/Diuhz9tVVuft7f3+GmvJIF3Tt0MCBYBWoAmmAVLPJ4GYEOykXmup
9wS0NDCA2imCI0JuAtfjkeDE/9x+3puT2BCn6e9nQtZEYH+OUrPebCfyq1RYKNYP
t8FPlWmP9auEKkAQgonX/rArcipWiXi0BVs8p6QiXN9NQiwySRliKTWQci++sOrm
MVf3/v8Gc2HW0GcoYqRJ6Bt1NpH1UHj707m0+RyT2xP96yvAvdY8qk0obKtdo3Py
2zriBe567aXN4S2rr60snmFS/paI3WgRWoULzxamDRRCsLxpN8ArkAyzjs0jmugt
asHRIckVNoewNkmKfovW7DgAtzPaBKL0Dy4EPYfVzzlawY5b7RG+wSbcohIKRHtl
GE0Fzk1ygrtEzRajbL/bHE3L2QpxVZf1oVLUe4yuWrlTeGmw8bne5dt9gMMCjEup
6PazbzYOPKPs7ufrX4ktvofwKMRuo+c/T+sfVyah3nTvDc+93bUHvTmckd8bzBEc
ZH7JPRgZBIravWFnjgY7q2/N2qf8BpCAUm9FsNGKxHiho4VSQFfqRH+WNutmHTtx
JaC4oHtwraj8UET0S3xvQlWpbIIr6C5KGPb6ThwOKenp26Ekop/e3T6Cank8qbNH
fWZGgJ3ceY5ug1sKSGh/7tCWXJGNJYjB8E8FyWIi0pCoHiS5eb5ABnkUQ79s5kKS
k4YMct0sg1797Jd7g8KEbEelE0dWQkqSyBEeC6sBDcZvR1kjI3L38ohMw5V8ZrXv
UV6xDMOVTE6NBTDK6FT5aXTJFD3yWEzxvdaqALO444cz0boPcl9pZ3ukGt9WoIAG
hAdf5pTyFeGSWzhskxhlYp7/n3s3d9OwWs5TUs5mG0DmnVXXnR5FVv14jHo2+XYb
nDOhxj7Xdf+hc6utFuzsObXbjwbNg9/OCkKahlxeDoj/Hxsfz5dGxXoTs7OHontH
FB5suKDiWwaOu3jwgkeLHCwTTkTqfMX9QKG2S0Eq2SjdZwCUXHR7FxT1F94b+sX5
JK+sVwtQMfTYk/Ktd5fv/s4b9M13QWyLvYMFG77TBk5b6N3p21pzKWAcdYyY9vOS
6VzkV6mXgV63gnGQy2hajPD1/U/yJVI1zqBq/nYtVQ+dAt4+ML7uBrGgKmY9mnuI
tSjMwWrbaHSQtOTJOAYrcI/TflX1vWBclhyqsFqW8YngpyU/iSIGU2035L2k9ecb
lAsrSxYYME421FtuD+QN8/5HKbgTFN6x2fhQ9Zjrhzb8KLk91wpz9dVE9msyQy18
pfjW99TefaTKjAdQgOZaoo2ECu5h9K6xbYMcUZspOWbqHSkNSROyTcYEZntpIcvd
ljivZfTt0lQ8wFBNEO1McLPwksIa1pRm2n7h0YX2U/Vi32dDcNtw/yVsxe0h7nSF
ef4I/1u24kXkopw3rKmGzcIl39J3J/yA1ttz9kA83XznJaPqRvrDvt9yX4BUEbAQ
CcQYj6pFWaAZ0vtDcjgosgMG8RehQbZazD4xkKB9dKDCC5y47tfcATdSNRy367lf
w7EPADBQgFfU9RlU4ImNsK6YwIXnYa07H1aXX8qtNoxzIvHMzLBVIZVHXh97hFL6
k8mmKV0Fook5yjyKGzJD+8g0LEZSio+feuFQiDLlIlfWUqVAYzb7Yjpz45+TCTxZ
/CR1wMpl93/Azh2NGTZPT15+ASWg6fmWP0k6KP9kH7c3W/Z11UrypoT8rQe51d+8
u5RSokcxyuWDx4rs8Yde9QIOm2CijlQzb6RvysD3rua5MUHULcz1Kk+y8bs4fOSO
Ny66yNaq1FF+o/3pNmci9zewBSKsMAYgQ8dAvEIlHGQ=
`protect END_PROTECTED
