`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2uuRQE8cho11gi2Wd9qLy09mNP+6n8LtdQr/aFeI3kmb/Jv3l2RSB1f5lv1njcj
5VuSVVPB6LmMqH/tdv+gCeIeWnCmJlAWAk/iYtxCJwgoZ6HWNaZMGsb91rhnBc0y
zRuLHPiUFplEKjnkVMi/cSygjHBFKav2VFAHSFgWcMrz0nA83t5gikgQ1N/iX3Dl
Z7/7d8t/MjLE0Edzvt/5yJ7LxEAE063TtOzJMKNqGXie8R97fepsCsMHqvgo9DdV
Z6W8L20wneOEQbuQrCRFTrJt3Vd4994ojWKWPYf7E9sJQpyVOLOuZJgQtQhJFkAl
JgNLlSbDtompP5uZoHsasQ==
`protect END_PROTECTED
