`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WiL//a91rzwcdTc8QI9n94w+JAIpq38IsUoyIVhFMbXY3e5cyiIuGBLa85Kc00gU
NE1t5+x9hRPym+DUB8dsh2Um6jUnJ1m8mh8Qk+l7F9u+MEngMIf8DzfytbvFXM4A
NbXINSt1OiBY4cRCIlJSe3j3CDfSklrixTTzIoC3fCnkB44gTb/rMzgDo7oui+82
i74+9Q678sZLRo0ToE9erRzRkbV+H6U9ZL6Dvp6O1htVuTFbn3273gtjqW7bkDpz
y1+cMocF+Xn79Yk9fDWTN2DyDCgfh68i2hiqbxbZ7lZwGB+ScsEVVHII/5PtH+3s
GcCwLP2mzw3zDJlNM1mUqpaUc8MjwB+9u1X11CMEChQK7qpzghVQf0WXpnC/UJyF
KhtV0WPUzFJrItGTXEGB1wloRcjHNnoVknjkMc+h2iSXQFktRia30EIZP/z/r0+u
yZlH6IGuJYR44YhfTRmiTsJAbDW4lpvn/WlhEZWPLDru5tSQNrHwHo9q6kR2ylno
6ya6KcwQHW0PWsw11H7nG3Nm05/fH8ko8DeMgqpOs4xoGMxjQL4HkXZcIxOI+h+z
tR7+dWPU6bPuudrNyxm6z8OGWFG4Pm9+vwhciUSGl8dTxjSF7h9GWw+k2sjHxgPT
q91HFree5MDm87JyFv81RJVsnCM3HFxqTWCUWosgBEAvhoEJyMi9y/Eu2TTy+pmh
FRj64wNi3YVdbNscn73dXzpL8ldeeF74DleQDK6s38iVo8PF92r6S3OYYr62jO7y
VyPSa76BAGmt3MRqGyLQi9WorWee6x97kcPWvBaRDePAGKp0ygg4EQT5bnI8pO7n
mq5DTIsx4tN76sJxOQ2yAEjXXxaAVQAZMybgvKqYK8HdC56jbJKRku+2EsWbp6d6
rNE1orzXs/TaiqcF+zMCHFDLNd933oc4ncmil1g4JurpGXCgauuZMSU6AayZDU/U
gtJCaxyYcC44V5yPtP5Lw93SsMynDCaed6VkqCkkRBDT6q0nyzSrGzFKfG4PKCi0
XxFkIVvqIPkjYS9FSzV+AyKnSPzW/9hmJscC92FzUZ4YYk/PWnUXVZGr7wOlofC1
Rx/1xFIF1vqe8k5QsRTlgEZCbvPIuqQv8rRjQAkvgIxfDoJMEB1GRFw0dfnz8ZLm
vrMXH5Q5wQDaenVllsKiyrdGqyzR+AXsZwVCz+IZfE82FsXPet80pCO1n6Z/L7MP
2xkMwtcAVenQjxwTSBcawW92FDrJVNwQpPbCi/wi2W0mM84AyUHgCvGuSZJrMhz6
sJToqRZurr4svJfGIl43D9JBfREWqzDu5xoI8v5RIeBI7do6cItLoISwfFDvuQgN
ybY8RfxlENc4pb/b/Vy6weU51GDe4ci/IPiNVfW2ADW9+mNqw5tz3ofJWXKHZyhu
CFG7ADeoqLDtmZ7WX/CFLqd8aNvcNG91gjp0Z3rLQV6fGrtjHvloE7nDdOaWgZab
rdMDuTfOzmaUvBqsQ4KzGMkL0aElPbAQZYLLFRB+Am+rttwnsb7g3KcZ3IvvqUxY
GNrixgsCZKXmuPlig74ARYJvb6T30dBO1lT4Iz2C+hg4B5xSriYWhqtMNLz4OSIG
JK3OHCeJeV9ucUcXhtDTs4gNVeGYKKtskn9EoNtQ+lPSXPkSDHBhTiDtk9MRzjHz
QcutwN/Wa6zD8TVgm2a3msxotYmciFigT/o6fupFUZ5wq2HU3FJYUz1Q6mOjgBVS
kDDI4zjCChZ0m8ZW8aIWfd7XVSMhNTlIqAiklqlmN+2+c+vGSL6ShMAWATPUWemm
edO/XYPdm0NvPtX99t9GwG06Qn8Af73ESwdeG4jvvo/6Q9kYS5zBd4jkkLQpEhW6
xHO7GqXuJ48cz2Xv5geYL22hrcqF19q0GrT9obQZioYOB9QA8zMneY13bswMEJjT
y8X1WzXZ79zhVNCPWM/4U0qQcWMS5cpsrHXXJSWIfcYUorF0sozo5TO2+emLKbed
oJ8apg2v2E0BYoi1SBUmjWLUv1SXtX8OrwPkmnJ/ew/ksoTwzEmMHTPb9p/Qfa6y
D9lplrUFuzDPZObm5KOJzlHUFy1E1g4Nb+UvpuoBkwXYjSCOt/NMwkNPdXozch9Z
T9UhM7v+BYWslUEhCyPb6FYiWVp8CqTtVr49O/+iRGDq7WKRX2p3mM9n/okJt0Nn
GmmvDbtfEdftnIUsE7jZiHzCB2c05nqQlfRQ9IJ/lWmO2U4O0wS89hFhspVsmbT8
+qNb8yUs/rvFZas0OMBXqF9bsbz4u1JacCAr/wLse8Bh+Q/voKOOyC+Rji6H/e77
FWsqEAfc/6HHt2ZWSweY3GWIHG421QkhzrVyMi5hAFEDkq0baSe7Zb7Rmb6PneCA
VhrFX+kBOheWlKQTfSDvtRXyIAIIuoOzqt2iCN/b7CJUfREQQzgmtHs/F3pNyUmz
YJl4gvjcrRB8IwQzvheYJa2aqKWZoyK6EuE48shp1kY++5I6yIqXUUgsA+bq93QI
Gydn4ZN+M2Z9ZZaI/4+oopKDXN4458JRd3Oe4P3sgkl2rBY12vuXy+SprWla8GeU
NypQlGqih50MSYTL62OpFw05MLZ3qnBeAX7kTZWUn2gslJAjoDCBH1BaN7tCEEoM
UKJEhb2DKhKETVzDj6SyOPJXVtJlmheUMHXhxEolGitg2Le20cPsLK8NWMNfIxjL
ZUkyPWrIpu8er4Bmj0x8PcjFBYs4MF+/jMGQwAI9HiPzzU5N+V0hbPRlAhch8gjM
tWwh4KWrtIJ36PsZsdtYCo30xGgzuftSumEnNRy4y6uoVTXMti3Bjfy7twbP3+sJ
Cf0P6J8XoYNB60fYGB5gj1jnXSYtyTAfNq+sSMKJAaa+90rNA90mex46cZIfyTix
8Zda6RK/HaAJlBDZIrY4gGzPF2N0xSUgDu2PAJXyjP5D0WOodYbskHhno7YVkR9A
UwEmdHW3OYRjJ4hWHYio59z2bnJOGzVFcFitI6+NZRwI7HWEHcspgy/yU+Ri5Jvo
KKKUBBIZlp9Cg0dwi1gOtOCjs4yNO8VeTqIFypnnvMD2nw2MCjp8kFFLYw7FTnKE
hdM1Yz/TqsYvfw39LzLT7ZEzOMVoeW1ajYrDW1PctG75NPnCkFbc+LpQcG1OxGkl
/aOi0iidyaCHbt9uxhi11ZTjR+OXYOWHXe+bmpb29Kbpey4XdGTx02EAtYCYXmCd
H7cQIz3gtcnEe6/qn9tF5mECTJRkfKjclOaKxGx35MrngBgZkMCDk8w+xwvvV5Jl
76y3WUbsL578wdwpF6tQxl6LhT4MAfymauXaPOUCAKdMa4q8VNIemWQlSxPlBBRP
7MMp/q/LCV7jExBwwPUx027s1PSvwbm7k//U5roNAZ9drXJ4fkdxzXBtv+W8ws6k
h5fJc4+Ob/Dfz102zPMo/i8PrMSw7/kiXJt18sgtpRssnp4ytqLXvJICSPWLJqgF
E+hPcQ6nRIwBMsyY6G206CNA6/wUd2z+Ekq5vXvzEzx6v2d+KGZ5YMCqwZ/ZOnJ2
TxQbf/Dnvf3JtieeadbQ+l4hFuzdC1xGHJGwRcXmGVaNBNKd3MNt5mKGSbCB3XTo
RQ65nIHyiAyGQPwc2PZA0qbiOltvpVVWy1qhUdU8WQcyQDb8ZCugVubYo8H1yAEC
kkd4yY1AZQSPfsxLd/d1XF9GkH3z/yUVtDKLeEPpgAJtZ2IxZaiklq66Lbw4qVhp
8z9r+1YNNAgE10HR6IKuil9tD6vcmwOmoafmHK0Hb2bJfWOrSvrA71MzwexL7yxl
Z1vbqpD14vh1HXW7gluRvhk/Ud04z+WG4eVqr1KduAHQ3L4/6MJXFCGGgbxhyZXe
snJYj3uHvBXICiU61z++Ikg9yo4GsmTx6cDj3lqSy2fdK1ARYNlcj4ZSxpGkOeG8
po6vFzHsero+pYtXqvq4duxn1bpVTQ3N74Ybc/Rgjk13k5FKLfYMBgnWdb3bwsan
S0j7/RCZDbWVkM7Dp+T1EKl8qsQe5yw4zU5RvPj0I4RqEqAPCr/NYSq9+4nJbKQu
RuCacIukwsLdxOEymM5RFYawixIPv/K6s0ij+hDgsAB1t5vrVQn1ZXEGJuAL1rRo
fKpgwk9BIv6n+vpNsCHEzuSv8yArDpLsItdmekSCyZPbHHArq1NDz2zT81nx6Eta
eg5j4k5MVHrw7nqh5c/1zfpFZG2qHiZZTi81L5imGnAc4k4vY+N2qeTncwHKRUZz
8eetUxN3wT+Pp0C1sbXYu/MqE7et6G8nevY7n81e9v1Bev0mzyVHhxLb/ahDJh4I
/Tw4D/jNneQ1EB5NvskcVTRecxI+uYLlbQRj7u+30hpqGDSMPUc0zWVYSULLqH0y
JpWSKz7/uS2yjxr0vMhMGGSmHBFegNE6rg5xQnsINjnuKmWTiNhCXdsETYdYY7XY
1ynwWVl4Qz12ULgBrXC87NGPBgMjbGaua9wUK2XJEHCUCZnZoaoPudSN8TVBLIW5
Uv+hih4yjlDFoiPGwmOnIUdeL3Fqd+f/jxCkjabUL7WOmWgR6ab4jI8L5+07FFwu
SPTdPvbNcb6+cdj7TFJexoxgSB3Rd6DKe8khxdAVcLAgnxU2ckw0lJivuc6p3pj8
fTWG6ANX9cU/mOw9DnyD/DWI3sJ++ywIxMHgEKAm5MLzdWtivqym8bQ3qhrQbAFk
iqZXJARe2aCZroclA/8A1XnZly+hBDZwE4KrO3dv9qgIwKtQnYBRJm5y3Ld1Dz9o
t2DNCGaeWY2fOqaZS1/CyUDgM6TSdmU+aXGNuzUz1jaT4w+8XHI7323V9+ca0Ann
Ee9dwnLWigCHa4ne59e2oGWxWTM2s62quWyn40UBHhTHKXr5fmsVbxNUbDlwiZ7c
Gif4cZFOmGgO5RD671nGy83BVRIJxLjb+A1eV0M8/AXwtg3KxPhNRWxlbC1aVpxA
Ze0sulaX5LHVIHbcLnuvIlHqL3UzsLfUu6c0dr0lAC5L6JTQgERu+OkvWRe9GIMr
7knM54YQrEYJ6bLfUK1fnw8PPw3HQM6PqN5imzDHaIKrtUOhsgIyJR5cPD6X/n3t
s9gDpP7KAizH7L0xJR2YhPJv6/C6tZbceoFs4RACefBnnVotyXKHtHDU3PPjYVEJ
FAbS0aay0AvG5rCW81gDzQOpVan5kOnTA9utFJKTYkxwqMNO6jKyeCL6DRmwJ3Q0
e6lUMAyEHfflYu9yRvSalpjThhlcLd4bL5wPLjd+v5zjjcYWyJ4JQ+tdqYph4McB
S6s/fCgHRUBDn2f9PV34uGz/cboyEr+0woURp/lax5Ws8fbZJCVmBgl6Hg+VuNLn
94IT1ehkOB78DrqHPWolr61Se0zYMMqc8ypnJi2nWQVgdyqvWfoY9aJGuNYF2zrh
HZYsFNjUrH6xS6vUL6A4+h7CrFHxxEpAHciGcck186+HmLhWmuKhRTPoa2Vm6Abm
TygWL0mKw5p3fVuu3RXpe9srqLXKWr7m5ze9GDZHBWoymBcoePQRL08rTZa6+R5J
Xdk67NobJ4ftkCxqC3CxfGYb0izZiiPXdWfKyU985LHeK6sPvXgb98NHM2omQzhC
4TSYOo9mLtF4ieZJzWqdhdfsYCBwW4RqjQLX01sTo7lMMyzsM2/+MA6gUmoLQOXr
5DUaett5e+kuRsoBHGW8/1JCqBx5VERnBC/lbDQmHbZFJPg5eg+odC5ujNDax7vs
4rHss87vBwNpZHVv/uJz1IQ+2++RuLoQdCriIOkrCgCFUCdyolBBU0pS8QPs1Ovx
XQumJ9r83aDxP2w9sZpsDwzmzaF/qdTo1z0l/IRaWsHDx5PsTyoZJC7wPqgTDWH6
buKYwY2mg+hIfxoRi3MAuJ6zi9EKhvEiNzSX0x9rdSHi0uph7rrnYhb8RV42n8M0
wP1Cabzdxcall8WguNGq/qbpZ7xnwxQCvwiu4le0oRAeuoymvDRl/X2QTaHpCvUC
Vg3FhjTw4ZO27UhXoaeO6Y12H07k8/ExbqR3NlkZpVPhw8wIPelY6ULcOgI0Elc9
kfdkR6sFbfxJyPs0Uy3eitN5VGdET1vG9mujLmQmKCOve1Z3Q5qKvtdQ3V+49Dr/
ZMkkJh3CqoDVgNuoQzaRV5K8gvb+bZdfqctySk5JB18NfqPDavyUyFZMvl4eqn+1
MkBIuARqp+ZacvTdMsSFwrqXPndB2np+9IyhoDRpGjNE7NDGVM4g5HQU6FmoRlRt
xVO/RjzDLUlED7AyA5pchVcoorct9sSKJbOvCXJ8Z8oVL8gv+F2CZ4lb/hDhMbh+
81pHz2o981RRMmD/UorKd8NhrrKQr9EhlRub3OXAns05QDgYqXP5Ihz77gDltpFR
hwadDjElIFi8D7tTYKIILS763oJvqGjby9wswW8tXW0unPagVCRPCQ8hoQST6hIK
Fq+UbSo+3O47BMBKwulUi9gJKmDiCln6OFOUVC8uL1mNQZDGlmcMMe66lfEJHe27
2mFk8R91RI7QvgqGQPU1qgDf3Kq/rt3IUc1wP2MU18UWkD5kjdFXp2QerqcUHsqh
aKOBlljZ7xJc/scXRayykgl84W2LtBNUm2AZrBfGLreQX6Ff3pCc1tUu/FYTjXIU
mKZLXZHUFatkn4utKRu0l0ycTlPmEDEE18sjiIG9hScIQyBSV9jCE+tNNFkgLDFn
fimH8yhlQzFMvSdEqPT6nnfTW+pPDJLriTcMXWReOLsjH1Sp9aAFehI4jkpcM7c9
DjVGfhnp5Z1P7pQpAtKq+nOOaf39Vs2VDNA/bGBrBRclhxDGA2gqKSgor566Kki7
bF3TphkhKxvlKOqcUCpBU/tHT9GhKYM0a2N02pLrYNfzd1vdcQF525QpqlhApFPi
I2FNyM+aXNcJ9pWQHre6skTbGHUtpyv2yxdPDZtQ3EemfuBptcfqmKYDUpVj2VDb
c1aZJOcyK77u7rgV87j4ptN25cD81s5j+4dOdhw03e888dwYdn7H0FefqoWOQC3r
E03rB7LbT2jj9EUFMJesqPp10ynCyIOnNGzJ0c4hIFWrJ7GDqQ0tVo2ZRj/CJPTb
vZtZE57krQX9dSjbfej9qP/2vXt93aK627aRQqRtpgLowy+HHhhW5+8Zv6Bk3eKH
IykQMHfDIp9vx95jStoyVfIaEXBEmJw5uB06B8LinJycw5ftI0NB+aDzMRemdfFF
6FNYh9TJuv2oWDSRER9wPAtmQEkk9Veux2+tebRNIO5iq/0fGvYAUIAOuJk5AnbO
Uz8o/o3XGfw6i0di97qm8V4Pz9eumDQwI3i6cUR2P8ZXp/TSQnWqEWITGBGCizE9
3vuCCLXR1JJ9NGRIJUZa3NszK6ceBnhKym4x+Ufeq9G5b6ZNe0Baq87pTKyWl1pZ
NfXzZyYcW3drcxp3kJA4FKMwlZZx2eIGKfwItRJR3n7FHhHVjysb8PNudcaVZT5Y
eCARpg8uRz22d3wIWRzGXMKvBzRj7vZ+AipFFeof9OpeFNkk6xrCo5GMHHnfi9EG
J23n7NEEX7zoCWftPyT/sImGGikFnj0Up7lsahl9QxeXM2yomJn/owTea/3HGUV3
5N+boYV61rCpN456S6jVeuySCbnB0mEo+xAsIlVGXBEU60VbUyTt6YYLpCUoBMsO
3SxKFFiPEGmuQbu0xgDywFXOKb88lnDmUm1bChZC0z74Gq4AV9dUtbUX/tDyH+S/
GM2nC87ZY6QEmzJaCvfHqxu/efZVVEzlNMf0sMBlqJUumQiEcopp9CcPZO7ehXtz
EvwdIAI27VagLEYMNy+qHh01SauCiI8B+RAR4q569AnnUmFPGde+Euw2i/KGStio
+PHczbPcHieUFs0+2G3djncHsm7Z0N1mU594lbi2tv2w4k6cWLYy4utGXSmVC0Ee
sEqwbIqPPfQ3E0BKmb3zoskiaVk2N23f6QZgkVE34Q3OppofDWinrIbdTQ+FAKHL
to4MtHw+y3w36lfcQgCOGdD32GvWljsvS/EhGnv7RBS6y/b8JurbjaTdkZfD/VIb
ibD/rB4pm4cIw0zwefG9vaK/HTMX2J9N/+ynKsm919m5Q+RIIwGmEKbTPmkxivAe
xuzZByPjOUwCogGH57HdcN2/3skXjK5Ls+vKpMdI7ir8ZjWeE9SD92M85xAuPlr1
rdtCTf7CFeXicPE8/Ug4Tbh2NtOMcyJckwlncgMSBenoN3DZ4TXDmG1T9us25Ecy
8BO1kcNXypciyM0U6KnCbJcoKLaJKhRbdxzwzeqxdpl6h4Xs/JxRvBjUx/X3eyAV
viMYeMWfu8geHlnskCpkaw67fW4v6ZkmPhknep6vwUJ6LwFdWMYtH0DrITpHu8K2
ONbohbqQ7Jy7heSMyghYe0FIvGasPZtEyQXGd24AEPLw6JaJ1ePXFTlFC0XIpGGW
gOzzdLEN1osvPUc8f0S1x6DcRH9m9ej/NyLJ3tNSWqIFvwjHH4Oivsuso3JwW2wi
KlDN/Hc7StGLu5qZ7Mt/BX00JP46MuScxUE0LsFqfEANr9V3BIH0l0QR0EjT0vMa
AmiYC2NJmC23QALTH8sTzCmmcRlVWECSJEWAxn3A9B5WkGHV0vo1ginWg1v1idZR
7YiCyUZkhOe3wlvRWwrPUiP4trxWefegAa/gz9kVQ8omqtqpgjK9A4khqLILhKtz
HFJoJcIFfdvCYefxAVseqguXvSGnkNXueaO/vjBwhwuDxhnSnhl1e2b6TtHO3mDO
TRmu2wAHrs3/XPuCtFPAL559WRejTrVQyPpGsPF2b4Iml7XXR53uec/xw2Z73nBk
xl/CvlSHFFm1dQfPD7+7mUuDLgYubIvGEVGDJ1EbxFFaLwkG8CcvZoDjGW8lJv9T
6ptop+vDPE+6auMf3gFVBP6iovpU07IUcBF+hROzeKAZU4k2UuCIQ7RatZLU+kUf
OOJ7k3dEktW+ATai3pvLLzelI27ymRsr+gb+zpc+QfEqzW1K8Dx3NnZn4SV0CT/0
2rXNe0aqtNJtBovM7mhHhSwO8jC/+Z5poBj94CJfYHLto5yAV3fa2josSIb8fGsQ
uF3mKlgipbZjKZD2AkxS70+2Ex//gwEqMLcYzNc5jDbuAF/1i0DzcLgjnFQxUUCZ
7tmb4xbAwOlmcfWcurA8kt+JLp7iiA6hAcvxb71mu4w01Kx2HuHpags+H9T1WI+c
2QUVfNMdn4tlJPMwIiu43oXMerzh2vBGXfuh6o+k8qGxvMrJAJ8lCk+VQB7G1EgH
iMUtJP66PN90R9iscKroOt/87HX2IYpqAzzyXTQ4EUlIqJOl6RuTnvpgFgjcm/gh
5p7ozifGBwZTeBbwIGiWfbZHczJWPdXm1VigyTs2Uy6p2hjHdnQCas2YvCzwD8bz
VRZJrr3U4c/tfnaOxuYphJUzQN00vB+HiwRNKnlsUXzq711sGdr9PecCqSYUkgPy
OyTFrfN5+eltzurv3lIqP+g16lrcfuyk3NQzsHi0iIXn4swwrKt0ysx8y1/zG22z
BvIiFYXFEXnXKm5Hepg2bd4+ysIp7Jgv8UZlywttVEhIo7THCwkHgxFSESHJd56l
KAoDYV0Xj9iPKFXD5DTDzSjW84aHW8phKX1gVk7TPBqLIifhpCLnuC+Ry3S5wR3+
TyN0kx2gu0PeiCahdXS4huCP0hQJrO+dcbEtiJ9W3m28w+oMwexK8E0BQs3wNR94
jrsCzOfSBrYE4MEwT7+8lQW1auXfbbyhlwu0ECvd1NDevMamGk2KYezGUi8yQYZT
8eaNYg+u5xgYCOWMrfU5wtbFOTZxOSJCQIKmC2wVJkRuAnFVAk/qu9j0Xn9ukHe+
aPDkN4TnxBE+O+6fJc4l1He1Qw1IIMI5XJs1I96zooUokZKTFvoDWdM1JLIZgb6f
tK/XLPIKeWWs/mzh+7fzqu1kSjDwCs4xdq58V04vi8KYZl+RlwoUTaaguW6X9ZRK
xNpDxRAUEeH0Fw4Xnbqk5N/DTSjWu31RAyuA+t42lFzIB+YT50FM2kSRepsyjFrB
T/7tSp2PrDqkiF6m5qIjx2uXEjI++PssvLS6abxpNu6fkpT1btADbRc7CQFUNv96
N9NwToLSKf8/e4RGY6wMyltrYhVqrtBtTey5f9wZ+eLmV5d0BDJ5gzG6kTjiVw+4
2HEDDD2sQ6uSDW5zfXo8lRdNrAto0gyXgNMMfDPTt/wuEEzHR4cZvMb1ltK19Zuh
tn2zrN8pkknYVLn5DmJmjq/TPi1N/DLt5BmfPtxD8V0/1D9cvLZXb1sNwjMpM4aa
FFFB/KWugewx5KV71cqtM46tJqkPbTtE1Yw//gm3AtEixlemAE4b5Zavmzfy6eHM
D6Sm0Yx7V11R4MYuVwxv+kyMpg4xd7UicSiW7EteyIeu7J4dSRfFo/XouCcB53wP
BbAi0eju1EcPF5U/9fLUGg9+1EMeZB2Y/3RnE8WisYz0FTOW9Xr6zMnS3nky6RKN
MhylC5/wbOCWKcDXHn4ITXIAoBTN5wm5A+SQzi1oOknq6NWG04RBXoCK/jky5dHu
gakEmxjiDQazgXKlERPRCJ02my0ymeU+OQBnXyb/wT2+KmIAmO9MlwAxLlPeh7fw
gZ5QSznI7VJr6uyTqNhUqbVpdMAdBwbU2tCj4ptUYkt/65tvMMODH2WS4lwVXI5A
xz7lr9p5qL4Ms4qLqVxOKE0bhz3WByFP5NC18WlhGgsrCcPY9cZLlqaMVYrrdyh2
qz9HxZ+ju0Kiqwcf2SxqgRzZF7RDVhb/zuoqNmLASJBjiV9Fzt1bg3mu3HH8Lg7q
Z0f5KNmDvTfJgiTf/2sRx8//3kZvBdyb8jWgOCK0VgLlTKvHUskeW+vNqzHebuMl
no/8FiuiMWR+HnSdFSg7zQHK9pNVlJ+OZ8glWoEXtppLrSarSGfAWjndGb4QSsMo
oW5GB9oz2XvoOlVOadlrf9JfHCLkjX6mN6wciR3PwqAU1UhxcA8LaZ8YeN24F6t6
Wa0NQNrQhMDzxxd1v012n9gEPbjxGfvsdy6HrEXxdMZLGu55x2iIk5niqbLO/gKK
Vxd82FBJIqJ36O7Q86dPOCyuQqSAGBe6kcKrAg4ZQgZhIZt7zRXhEIdrZsk8nq5q
dcNkChMyR9V3A41vF8WCNEfvSOsviubCJwOPNRksVOp81/En3A9F7GN80bH56OUL
L6T2GseznxQD3EFuB2tSTllhAZZpddq8P6zCCwSB1vWMd6IwGDvjL6lVWe8lFdQl
83L/pQ36Rz2oar+YGGBkmPzY2zH4lek+ejJb+Wlhwf0x1SAuSuJ5AyfNvRDo+j1U
z5nrLLlN0i/QHZbIyaU45pHUAV1YuiAT8e0cnORrum0fj1sBdy+L3KFax72aUje4
uKbZQAovCoJZ3jPchuYlAxJTcf5WFmVy8hV6dT1FcKlkrolv0/YiuiwQ48tRpT5j
HqYGIiganmc8PR/la9K33Z+0UgJyZ6dQxOpGYr3FemRqwNsHFKLMWj9aybYkKH0H
WmeAs4AEx9KYiUzx1XeSzIVZuLxH+oJXkiFa9CTrXQnJB2+TWgmwDsfzBNBVxGbu
jTSY8s+TpFeeUoOyz5LQjKYrSWxYvJmEPZOTLSJY2O/l+KwnYoSYZfx8UI7P4Eyj
2DX9NBgI644v/eZleK3S1wqBBGJpFUqX3cdJMTtwGWu9nB7vxv04MMUe4jXBvLB1
nsVmZCqiZ2GS2G3AtC0IXiVUhNfdqx2nyIOyj4jVg51pzKtiAL4kGdoSKvJ+bLpN
mj5UarBb4bTlX8MFr1kf5h8H46exzIK26AwJfoKEvAS728Q5XGHiIP74SwmvuNd2
kd10qTdTduoW8g77RBrf8qmc9Utsbrc8iRvbcHaSo/fwN5EfHsecjhzpdCUgCDvV
n2PxLg9SeyYoqAb1XIVMOqZ2Cb2Q4OhIMw6zVUqEvQtQDES3I6iYX6uiLTC2LKcN
Ip6zwXaz3P530B7tNRI1VSiP/LUhNz3pNUMi9z/lyWODDvPN5DrPu9QAldXDicdP
AVaMh3lHbaM1TzKXgUeGV3qPAtYyFIJyzrEXvSH6/mjRi8xf9w4kAqkPr5nyHmuo
1HmamgoqnaCiynS9dXn+/Qu8Md3486jihxERSNdVtKUcVC/AopAbaaz0AZMVA9Eu
chTo6kHknOb9TvM3QDnRiTE42YY4B9MGtX/YtQtSgVdX4j/iyceR/3M03mWvqXIp
bXTFt0sjKFWtx0KODdTFBAlpTMAIhpusp3bIz5VXTO92qwKKUNIq5D5cdcsnnTdd
Lnzj5f/W7ng8LWKePgeOAstvz+5clKX60VeQ4K+D0EYReW0Wm/qYU1ck+mDRxSW3
2zGoj3zGmT4R0gMOZ96bPYazggEaV/9UPk6L2guFW0wdVUpg1yUXc1/q1Cviknl6
64NYhckUn3e2XuARTxsfIim2Z7d5/3DxYZRtZVmIweWQi/NhGoZFhhye5IShhez3
v8d46jqNAaAbIM2loPj/JDZisAlhekLvhCtmQRtHh1+PuY78TeoiXygeYUgUD3Um
vZb45Yiyj13vxduO9pdTzi0r1FOmJMNYTSGR1T+YD77aI21Zwl/Wc4jQ2+36MxVA
TrKqB+859U03POW7hCuu3IhjxTRp+VuXYbXwMvwhJF/11JTPj9zbg4Q17xw1zqS5
MGGeil7xEsKxWdePKEHMB6Nh5uT5pPGnFNnso57BwMOGw1bNuZ8diZRlKKYqkKq5
kHHLm/czE12u8E3J0w0pQkhSV2nYgAz2WdTrdM8nO2iVuYfR2bxr9Eh62teMHWNO
BPtRYouAKhAqbND2lHTLWWy8wHcnw5FryagCjO9uxPusleTNzL120NXsx0znVAAT
gyUhLuAMifImpQSuSpsDYtqp4XsheYHYr7zk7enWnYEnN5GkZTKSPXkrWe8vl1kd
1icGEmPKRnWM8uX//BoEtuzXXUyML7+SQgRRX2zWnJ6tKuh9e5GL3xK9xHGPYOgU
GbUhTNMDxPLjqw+GTD9xcBADCC6rWc9LAGw8UTCBuMWZCA4MnVKrWsO83cEms8wj
w5/geRTjn5JUeCHGiX6ItHUUPu2+PqAP64g5FiItlk0NVgnmF5DK3YACUsNljEWv
APDPO20Q+X1PRJYhNLKOnpWfnF+me9U2rlbSdHJZcfmw19iz6gLRFe+rLB925mmH
1x1/cWp8AWuaTodjq6UDg9+ghrC9bCQS3SAfOyp8A03X8mi51vzi/LQjHLilqEy1
XRVp3iYTiDqXxp7CZu/sB6yGduY5la1hOibf+UiwcVCx8mZs8GA2oQni+r864ARz
A0GuF9L/DrGgGpfrqHBUhO76k6dkNvBWBh7yY87pRpMSBF9WbPH4pwVKPJ/stgjq
BQUmYf4kIhUzU5Z5gImpZALg25Ow4LZNtu1vp8wwhSOv5evel2QFdyEK/A9fBlvX
PPBZO9sxGGPBtnx6Uq75xnIRmDsKLLfzyKry24LvkRVW+0xV9G0OpSPSX1EYkWle
WbvNL0mt6YP230Zv8KoTagdVX7i6bp8vdsKmmp2Mk0D3hSLehHLK7XLzZmRAuPKu
JeDppJ9w6IfUkm79oZif4pjLukgzWPtoVYyH7OJVb2U8Cr5PXlm6eeBXMnUB4BtE
Xb8fPBOnIT3j2ga0m7m3E6OYM5Cmr7YmmosMIhysw5U098qmU3owdJpb/rzNgaJU
Dvr8JTPQf7vM5RGWjgZLM89xFWnY4cUnstt+fA77DHpM1KNEZWuwpIyhBJC2paN0
yAmyh++JmtAgw4G0XonwyurepTRBjBfBBgSEC3xvh1XeX6fbBRewkiBNHtaEQflG
QeiUO7hP5Za3YTIymZkKnb+HmYftLs7gIHaX7R8TioVwbMDgYWh7fVWCZa+yYXMk
8Ser2JyYOFLLWs4FYYIynyStjPZz8P8ePXtuDMOfRkGTNS1kOkJcl3fBU8jqtY9G
VLOxJ3KtKS7r3l8CA7YL4B7l4f5hD8r0tglIe4E8TsklH8eBertf6VWk8xAUe1L+
cxo8HelUwoLij0LXtENuyOZvp0OGL82w1+FqSCw4E0h3xM19B0bHC8kFsSOdh3tZ
OWzeW6T0X11YY8htrCgCyNqf2TDIvBTERW+bXf3q3t9yaEuCCx9VSdz+o8vHCzMB
QvBu5DPI1UgleEPnni9B9d5J4DwwR7AaMFNxn6sx8jiYLuyTZGJplWoP5OCjhU9a
hleovrQEn3rplZlapVNSF2mxTDSYBhD8G81nvJSoqbiscVff6gaXBzXaaXOdrys8
prubOxHEQt5JO44njt3z/zUnb5p/8SxVZqJ02codD6yObFwLZsEc71/jvsYVRNji
3IROEwLbEY/fYa0HDHdrAUxiKcVWOxxwsvr2pgMf/iIpJL5oJUyomp6DdJ4TbOWL
hfY18IPeMeJJewZPUrxRLSs7Bc8lQFrrn25Hnq1rqnOJWimSXB6J2xhgaSg8fcJ5
nLpuNkjEWwQl0U9uxlv6/slRWkFeBfzyXYQRP1y+B2Vnt0Mcq0S8NtFYsh4uL7WJ
oTJNgmvkSA0oke4VyUE5ntQ5Vg7bvemL33w7LuzQ4XIJKQlmgV15kwtgQK7nAz6O
vsFffkOTEWCoTAz90ueT6/sZQuSJsc9AYQhVqve8QMaq+Wm1K4pIOJ74Iq5mXE4O
7S6H0u/iWojybpmqSbgb37qGJ5QkA8gLgD/ThXTzp9P3X4iiuqRkH4kyagRj5fRA
Spb+aivRt/FKPog8DrI9SqYfWPO2VTfOjy4NWteCeMgqyjGR79EFSyjS+wkR0ee7
okg5PKKtrzSQwxzU01KS3A9qC4bNI6x3T0I68C4TZqGS40C4CHAMXBRFFqpqB+Bu
DnEasXb1h1qvdXncxdKm0/XBKHHAl6JZ309dUUTlUisd96tIZLFRcBRXvbXItXlr
mjxdCoTNAvFs0+PMY+YgDdv2wG89ZBUltbnFtoUscQFx7vkSe90KappDwHqKRe06
yj3okv2YTBIV+QATQWC2AjwZvxdnQDfkr/vLBHpK8RMMIV9xx7UD8Q78HO+DGnzJ
I+yf2/T5Rb5VO0pwT4qdu0pKwt2h5AewlgPcpkF68bRQl+UY1PBEcR25zlI/6GSr
qPOB8+6QS1Ijpj8gJydzjn5d3OMGT81dbeyESZcdw3JJIIKCnbXeL/orPltP4yMs
7E7ab4Aer8zH75+KH7obJWOICo6KhLAdlLw8UazAnarWKnjGOVro4L2V7+U5Qqlq
hksLr8vrK2DoFS8zao8ooPKlz/U0GOQ1YGco2warkBbGfQ7Z8rz9NBCT34GlAuC+
tOZRNnDqhYZh/AMZsVIWOfB/4DOTxgrSofT0v3T59S4z45rUcyhiIIOYvRJHYfgs
4VWc+tr+0DJykWAO5VNHw/dvpoCrcRapzA4zFCh7+0Y52AcvhnawRN5IJpfNdhsy
7ZT+Bp+329Oy0DtDwyXxqY+xlg19TyVThSnT6+lFyv4c7R4/niypIfwk70FsrR8H
JW3NPub8EggIH5ruUMDOX3xXSXHIH5Qc6vBTTgjK/UIDF5b8Ozt3+K+I4IjPu5Fn
84AOS9azuMhjBn2yOpaGEB68gbw7p7VBZY/oBk3/f4QYjSujYyrxn1g6Kz9Uy3Bv
t+Nl3hyHliKKG7UcNdvlu8nzHXKGpJQ/YByBiKTBEJeXjXZ9hDQaNJomgDq1Wn1M
8+1AbI266fG/QGeCiyNXrIuR8lqSDcJyTV4pbnqqRslfslw6UnMGrJkUDq/k6U/7
qCCXVWSknoip1MwJFLWH45lHZSj7ZAApXfirh8YZMlDYOFTlhYfQ0I/6wguLQKez
joesIRe8I14L96aWx0wtiXt3Cd7l4tCrP9ym/lkfUeIKCD17u3PGzlb1GsQPsFp2
QoTU8eOWgdstM0KVggcyYpUCa9CLiYJxafRUbhbiEww02CIZ9ECJCgAIOF+Fxskl
CHaPDT0crWfsJ0dUHNJsR9q11cvB1DRMjcCbRl2ridBZ4B9hwlXd/HkU908WaBbK
K9H2W8/et315baoFqoGJbWjexskapEhfy+DrBuacAmI5ky5VNxKTj0TxiixVMWnX
LYlKhmwWifeDt/E6EJe5SdV+wNtEg4WxI2pRIIA6YSnMsHt+xyrNWT/sx2jO/ja7
xcFptV6IiUoLKhRqjZXilky/sUUOrhetuVMRVAGI2q7Dwp5qGBjybZVE+G6QohPF
T4dXxtRxfqo5j4w4WloVvmCCuQK0zuLpzAIEXXpYGOFAT+LdcWRcc26rpr2Bd8lw
l8ti7ZWdw+42TCTIL0KMzz8LZ3wjaCHOkOJVJ3ta9BIBBMDrNPpIv4Ghfjzb/13Z
g7gB7gO11SjCLBaPycZuittQZHpJyWBnfQUrqqc+d5+EKF0et8YUeHdMq5UGgvmN
aDgfITVXuZi9bDCFHFtQDGDi3pkRY29iDbZzrnkc9P+ehBZU3+A3F75GMX9tmbPJ
g1bLAvOHg/6EAGpbK8O+6+ump+kqKfMVrVOju25CIHhKoHxKKPzecxq0z5HLVgXh
04oM026Y2QKDOFHWyp5fF92Aze2FM2eW5LYhi2NotGRGj5N0rkqL8j6pURzSzJXN
0F67Zkpe980nA1/0/ff4Ek4P8z0NKVlbIAF0FO6tI8Wh9tEYAq4/pWncUzYjFbn7
BBfQeokLCUm6txsG4I/O4c1Y/e89LhLNsfo/c7xoYEJOfe7W3WPqgD61+doIfPhX
sudZu8VzDJicVlSVuZYZK72vGwAulzQ5Fe9Ely7ozXeXxH4A93R+He0RanbuZQlB
ix6CCT1sVtVHCe/HDxNF/JC4Vv7m6cffZpWiixQp0y+bqF5Lo/kYHexjN300H9a9
2yWUIIohMjLYvo7pmMk4BkvDMeZEmlIhij/Ez7M3/PF29kuofej69KpA1Y2JJURb
D90rj31A1lB/YIOYWi68YS2StFllA8h1cAGDXVWnPGet2IX5/7xyu047FeHSaj6I
Hw0BPHyzBqmxfFIOrht7B8K43Dl2WLWRJVKjP2lwkWx98pHrqx5pQ0elVXnetv2P
dnO7UWmhJRPRi7TbGymPsfUCOG6aE6ovstTvjMFHnCuestkgfimrGrmtYY+US80U
WtXSBzQQRQcEglTw0zaa8RkGPUIPOGKYy3/kT0WdBYQtnal+EDWidRBL4r6HD6b4
s7miTJz+ivC0/d8p85s6MBAZjYoQ4fp6FJGYbpnJEMNmvWNFCXDvSo77c/NXpawU
I/K80fOBpVKtFq23+CCNlGWYvD+naeurTeWmTGWVAz5EETr5ew97gfE8Ikgh5hJf
eKtGGV2IqhcH8AZy4M0o8LiBXypcyahcbt/q2YXSp4gQ1aLLCNgD3Sz1qhwJ8IXY
sZpbl+quU3abXZ20v6xrPVSHbkn8LjU3dNYKyRe2Oo0OjTm9d3e7Dc2b+PCxrb58
qTd38rYp/aiQT23yXapxINpHwnHv1GG1fGFIyfplys+klNDkciFSaHjx1eC3i1os
TOSkaCWvsyTd/i6VWQJ77QDM4qb1b+1wyRjM55FydcXCRpdSCm6erlCmkas6LALB
AuervfITgIqJMt0q3w6G7f5o1xLBFMif4ZpBBKpsR+XRP+DUgLd3Hbblu99x4ZPX
BULRlEZ9k5OwYRgKZsVg4WhdWYzlLhASOqEClppOPklC8dDyD1Dh31PBRsLcqrzK
wVkQgnrzqiahiNTo7pTkXYscDfnLwRT8PhyQYFmWSItu2KW5qYuyHnQeShrVRJnH
QM8+2R9GKYdzNG9y3E8tdoXkO7ia2Ee42Xrn+zasXNcjWa28JmlCDnPAXkCAyruP
iVlUouKLtaBC7ppb7emGgxphs17GI7RA7m562D6Gy4CZq5EnTaYnk8KcWnLBDoDt
HRkUWXNmMe8H4LcI2gDhr3AFWzts8SzUpdQ5EGjUincZomCracXz1Gdw/jWL3+l6
ipLQ2OrC7XfsWv+DBOV2APD3E4ZNoA+hL+Pbf6LYaPJKAMxtosYkOxz/KWh1lewZ
QaJsdd2guR6jsckXp7/ToCdA0bCheue5xwEzT2X2w6QsULfRnLir7I+yw5n94EF+
ZkeXjVnwW2ZCAoY27UpDbT5VdzMe3Rv7fvSgUxA6axJFOVEBfQxvj5VffNJeCed8
PVwfBiX5f6AheVw8zvWAKVB/P83oGiU/HZTqyWhjLDBft7Yg/H4uASlQDi+1C2Pt
vpvERBc0H7iukBzh+F4tQODjf/10dHxC9IFciD6e9xlg/8MbEm+NBQ6J2COQErhn
zbBX01Ktcar6BNnvRrBjoKofzPr1Qt9APCO7NUTGBu1UdCrWQjlW2VcDRkGvUk9C
PYUIWlcCiGHpxadYKhCDgRnXGA2mbEjN64xfgIoD0Jdt08yAvFsBPDIImLlCbXW+
2gkidY1XDHiV0gMj+C4G4ITvRTmggrK+ip7CrQgcGCVCMxAKQHVFwlfBRyenlDS8
hCj+QIWXuBNicG4Ru9iSORogqiXUPbvKnyXQFEvOUe0uBn3Qjc2tmJnSnB4Pkg29
8juzn6+FboT3R7ycCy3zC1jhWOg1qAJZvvxFKLE6A2QRlqXKvvfSUqdRwE+udSE2
bSE8iD0SBqe9J0IYipakP9ubHTJTQJjg4RCx4DQvN+5NF71lLqybtcF6jnwJBgpd
Bs216xJr3zggp5S90Rcjm7cT3wcL4MNj+uTf78qXDkfMyCumWvPF4zECmdByO/Ha
ZJEaFaiE6n+4Cz2UWsXt/mcJZGaaesWXAhOuqSzx1FEkzMEiEbkj+vie+lOc+4UY
xpNpkjofNKqdG7sXpUsSujxD+jGkd6Q76XeXbQ9+N0tYik05HzwULPTigl1fWmnu
s1WF1WkPJPJ/86Qz6GjwA1HBjiU/1Z49glAcfHhAdzAZ/CF+JOMO6nccvnD3gifV
eeJv6cjVtYm+fhX7rLB+yovSdu2J5PvsQ3M+LW+vyJmetrCmNrPnVOGtYdcYKr81
vaYBt0jxjZmIZ4XJygtvT+TDXFzCt/dd9YDArSgG79xEpZJqBOnhNiUS/9PfVm7d
//bawkHN76AZibRddQpdUJ1aR5R6LOg9AP94/yHzQwkLvZTQObRsRmWgtWFCH7dL
mGbCquLVVfBHLxGolmswRU1mcqjaioTQ66LgnyeOpVCESAq0mZkaLWL3aPBlKHzE
5DC0yK0iEGvwDNwCPzP1+7FvAg/lxlmEfzgJRk8IUDNuXHhJuTvwBq6qN0hT6+B3
xLb+Pl0lRg3fJPGKFM4YyNdVnPUzxnoTVvuU/HzfvAOmOrOy67UwD6kT4e5tMd+0
TrxE4rbcZ4zWnLFRam4KQPXzkeN7VVihUcA/N/a+oQ/87CM2nzDsOimM6xZwWlne
kDHLNaiyrPiEH0REEnM4TyPeN9C++T28EY6/GHjkZe+XtbwHxVRzvkSor0BhikOZ
UcLyfhzdA//NWwtzPXPZBwy4+FEAmRzorFGDbtp3o5RKny/tPgVbSK1sANEUUJK+
0RCSMBQkZE9Evrrmr1oHVPyV6GvkV4XJRXn/feyBad0TjsNZtglc1IILsuuiBt+H
TrAqP4bUUiuXzcCbckKINlAz7z7lMAR33nch+PRGR+DEBVqjVie/ob0J7U8Bw884
iSE1CREZcVznAkTPCEA9D8gAlwTxZrzxYqhY2dvBwhj8/1yIp9flraSIun/cjgO/
RMgORiSxQXr4woyGh3lYRbrndqCl2VhUMT8v4RxF/iW2vdJwC8ukzmaqgiXGoXD3
Bom5NF/asI3aUDbSBGkXrxwXfUgMycoyLwDk6IfkS4GdFf6WLT9A01Thc3XInV7t
dpkRFjqXr0hg3lvPylViYwhu8kBakVP1irAneSteJmIfPxpSnocZZWbWUgLZqrmP
ufDwY0VYwukQx6cQ+NwRMDilr8xklNzyYrhkGiYhURttKWA8TE/5UW9fLtB0MZrS
RU5Lk4U2jE30VwxMpFRaoSViRPvBhxOTzdFG/nSXTHSRbv3tGZu9GypXQTEhGTIG
gwDtpkjVp0T0+SSlQRlWoMfIY/sr+T3hPuo0aeRpaadJTP8jWtHd1Q/OoqO9kEmH
3MX3aGraC/ggosLdXsKEeiJDsQO0YMCD1u4qcG2JKTpskPCKCmpp4VvMAiTZ6kBf
5gyNpce8N0eQRvzM4ULsa70/Jp38zLl+FmBMiH8e0bvBF/7Mvjb6/PpSAZI98SZS
yv4jKPEwPVrf9L7B3CWiem/NvbNrjPP02LrXN9KK4LpIG6kjGmsV+zKLpbq0OA7b
eVPo8qElzlOLybkGM24OCT6FwfuroMfjdLce2JkxQIcuhs/Zwo/vJJk4h7vcm8sC
Ysbmynbx8UzywdatK4j8IGLMCubGzDWYPTu5K5/OIHpML9A2lpj1+nxx6NKk4fuL
V2ZwLV3Vcl1UgpWWEuB2hmP6nHK1+sz+EUAxuuyBI7S5Zdv/DWi1GDTAjThkhBE4
2dx8gpFXZedQoBv5sSacPnkA3sgasxhwJrmnQcL0OnucMC52GlnzqNs7eqgbhxPy
oaFJNyUaHI/n8NcHJZjuk1Tatz4WgfdQbUJ1Pq8tQDjKOq1dbjrTZAeyrDA0Q4ir
SdwC8ucSb8BBRYPGQblEgRLQi+Te/krn2FC709la/9Ui8SJZgqeEQVd8g4JO/PXR
KRp2eZyN0mM8M1KFB37vVFOBAmgwbShLcueGhPU/N9VQ8DAsS3nrKC1b1B1eZBSd
tJrvizRKxLRsbZZnr26paNK94MoezO7xY2ktK7L/NbCmBbYHKBZkdcrU6vXfe3Jw
KDEIkm2X/8Y+6DrbnSB2lQx7IXNN4U3bNObSOBHZ8QSkImqci7Gd1qUXQL/aHXVs
5KbZHTYYq98xqOLlJdu3Gx8o/6ByUe5CmDoIvSoEYY0uNg8gjLBAAiNLmWKfgw33
HMuVqQhuF3C+o/8784w5Dfwy4cISdepSUN/bTRQ+uHilUg2KxXl3JXxUyTlqJyLp
CwLhwa6mPM4Jy4alhLUTXSyaJhu8FYprfjhtjQcD/UV1JkxWpx8D2PwuYUGXDGkE
IrKD2kms+anVFdzl2lXT9ZCw6nqacQYjQfYJF7iuZwkaEXS235dGPLT/akkitWOX
PvAc/SmomZ77Qn86iglaGvSW9FSBbIZMTNcanqxaCvikM61IfnkBfSlPkrDShP+8
QYk8wYlBIc1+ACMbMX3qYN5SDmcQM2UB06Fxo78D8vsRDcFakWrH55tu8rbtnchY
NbbU9EikjN0wPqv1068C1NkyjNCCIuyLLtd0TgG4uRs=
`protect END_PROTECTED
