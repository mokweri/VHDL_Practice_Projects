`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rV93p9PBI66kulS6EmcUSyBDe+F7qMQa11NeRbcgH0h8C+cibFrx1PQ48+//A4x0
4UuvyhX0ERIQXKmzNvxYIyyO6EW6qrA/nUexkUkkHYXwoA0xvnP1AJqz3LtDk01l
VlurkDFVufC/Puvdne3QH1fyYOxkQpiX4GWgDbRm7u+Z72An8GcDWjHpR0XPIUCC
/Yat2V5UHx6p6cBdu+JLA6KGL8wiT9+6m1E7uLOg3ztAuye4XXZCFN9X3h6Ux0bS
zxf2UVl8wOu5t4BD8//djm0MwiYdCMIKM/xKYDImB/7WJ2NWQA92MtYDnHrMIjG2
4vp9xzPFm1+xo1rPLEFp77+Zx61iwHi94C6i58dgot2HmjK6uhEFHaS4i29UaeLU
JynMj7TJ1Uz/OckFtzNvyuW48kQUEIzqBR1ucJLFcqvF//527qY8o4WsDhxnISx+
lr0IwbWikD8sFz4i7Y7AoIDYjfowT+cSk4p5/mK8Fq1dSia0mMVbNxKtZlyCeu4D
AfSUylV16pwjn236g1p/U37a8MpyvV8DOEdV09sJJrgzaXGBNjLos2cRmkevXlvo
fqH61ysgH9EsxGYHi+ZeOFqHq8Ma2OCY7CalHV0eUx7zAbOADH8v9WA9FRbFDMV4
dpaGbBs7IgcbDsD7Qv6YDpebtUXuVv16DhNKWTl6nzMWC2ttExCTSBA0DehqwB+4
qKvnDztrk660gSLpDIY5c7mUbLGmC5uDEeNztGRnFQMJQExKcKkUn9y+selit+oW
RiKoq9JFJfNYo+bDEJZD7xHijt09I2PfKZL+LWgQqJAGIKymjwDrLjmKh7r11pjm
Fja+C+FOtGmdGojHZ4iPMlrVSO/Q6K8RNlvRHN+APY500k/240/26Qd2MNkQiusn
NXeJYs9PM9phOb4FQxBTTu1DPl2gZdehU9ugonpnTygPZ9cgq/JAPjg/ae7fbsrn
x4qsuYibtZJk1/t8kqqI9koREG0Em+p8Z7XfgoqiRRJLrTUschcRPRsnDpOqv0MC
aVt4NNe3c+TDxFxTUNLQKVntOWyAIvlgT/PJ80DTAfUPHUdm8czYDitpzohJdsBH
RO7wapOBoVMGJsdUa0vLw1gHj2OLnKPrcn0WuncBj6xRZZjqfb25tb8TVZr7lk7U
PbVmI6UzdH0HQsQCFDgJCB44w6Q+rjUBx6+VfBe+KTt/1Bwee+YpJi09b0MXF2Ro
cPFqIQwe6DCAjxhp75X59rHQw87RT5E8Hx7BcT9II1el74dSBOylmeNAHG56/N9S
feSJ/aPr8aPfaLQ3XQDf2qZJGxd6CpqhxIVr2hWxhVBKRKOfOM9+nnvntbrVvvq3
JkKai2VIiQGz4I/U6jIW/vyfL6GXxsW3ZwvgyFiIygXIotMIWJivimw1bFaCopr/
AEcmnq/KSZOBU+3E7kTzIJ2NSc67uUydxeu4yfAjgYRwkvl/xdGACRLV+KcPX14A
P2p+knv2HFhZDhJDEznzQSQp567m28iMT4JrwX4SpuO/rBswjV7CarYjDS8BmiYV
WfckhLbLZiVqCg+XEhPWAw==
`protect END_PROTECTED
