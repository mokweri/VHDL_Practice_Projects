`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l4ivKPNEUBgIMntQM/aeoPyF7ESTMlcwC6zItq6FO6pHI1m3DoUI1qR+NSw8votE
CAFETPSywyO+aLY+XgGSz3yl6F3wxfKdgvhzKwRecRk11DthK4Byoo2K43zEqAbB
Kp+/C78stxJUbrLfsyjnZgjRhbztP9FCBnlABj2gyONi5jCaZnrNSvv7Y7i7vZQP
a8G6FYm+I+RFjzf8OOuzKL+8yXgWroHbnwy3AoDzDQ/uKQ6N4W5hdZptriE60Mp5
4v8+T0Mua2EDLODMdeGNepV+XRqSiyELUpyqHp/4kwX/Rw9BinEmYfFP2m8V0HCW
f00QB4gCEgPDhaXakkYfYCYgmZkzexe28ZemAUfJvOa++bW7rrOHP6mqu1PKZ7ci
dhO52kCTKwWaUq6NDsM23/CQfQTT19xdb7d+jMBRqik4InS5vqAGwFkx7Po5cYdo
3FRCxmhOnd2a20Sw3cQkcnV4NPmBoNqS2qAXYId2QKnDj2ifyckLsJzO0snu9n9E
BpssjRKyufr6mcmYltn6APo4EbGfiOYs20SR5Y831HhvQ8h/Un5kA5kiodTXWgXk
+lSE+AmegWKFlgTbszWKnNqge32BXovEh3yV68h3/TRqmcNSqBYBBnadgUPqM0SR
WnfeLKvrmB3Xgcupvk7G5nHNFYHis1cjCVBIrH9GyTi1Pmf3HXUodUPs0ZA72Dxb
AAe06ppPPQOmBCBVPT8V6ZA4WqKAyeHqT6tu7DbRDu5d9MJTnF2go2xQBQwoKWCs
XUu1I5NGrIAxdPOTK829PJa+ldfbtNihPi14SzyXgrVS3Q5ELxIBPx8OD3SHfmMW
FPm7LXrqGTzTYVWRTXzTrs/J/k2z1AQXIAIM0h5ZsRgW4EGzGb9WowsQH4MmQdyG
kQSIgt9Bdrvw5rQawjfryETDgHdnhnzBSZWnriojFOQNn8lukOgvGSgRzIfwE+3D
0nVAlWBbjcWRDbfIatg4/UvCL9ST6wOviXZZykplPIws9au1E7IjcCFtNj3gWc1Q
Z4CrayPiKiEPSSk6UkbSGk5GhYdhbpMwyVX9slmqeiaPJdduq8pUqv7xqpD8tcKb
Wy028G8H33g7pQwL7c1swC2Q1msWKIinO4+WpVjaRZyAWtyGI84QX+W+OwDcHy3e
8GV4QeZAj02IGulR0tCqYRKQdqTpEky33wQGZSQedL0xV/TsVXpmUspGiRwRI2Iz
noSr7Wi5oqnANkpKPJbpPjXVq4wUW84i24/W5IjUJFH6uXv+9m6jQOtzl2REJJmw
KZg3QctVklBRasrx8tf23QVA1xszQZ3gU4MkT5qpdvv51ZDV3U5OqppxyKpbUWtk
TqWtAk2hb1oq4+6eqLLvH1KDwOGkxmNlenugSLRrFGUJfepg1ny2kXmOxadyFmbK
T6l3sndvjvjGTLuuPy9vdESBpblc/dTmnHnFZyJGIWUGFOg5WA5RRFMhKcTVb989
Pvp81Ir7FDpHBFlpbzsDnBq8Q+L2iq5po7aZY/zJpeYwjKeS7Rrhn1kfmBbIaLQN
4NeQXjlZmVG/fHqJY4GIUI3tJ22xz13N7vbzjfOnlpey2cMiFdlVWgy8WMfHoMdg
gTEZOHQ/Eza+Y++H209X0bXx0/d1b5ObCJv4ybYRdr43tcSAaHTZLiqgHasCtX++
C7YsgEHwNRONpzjUhZxl4+/K0+b7s+YHo1A10DDezQayGiUEC5Y5zejOo8S4DPsu
Y+eCoEoy/W9mly1ZbWoLVDCrWipK0yUxZNILk/fUT0D1n6F6met+kJJJnv/+tyR+
ydNahR/fgJfWvIvH3Gj2+oluvtbEtzQMqWe4Ilq/kXNIqzlkcxCKq2nnlWw46zaB
iKYojNKxmkDxeztOCJBZByyssWUEWmEkjiFGHeHTTvpvmLNE0jE45RBCRg+xrD5t
6W+IRjt5ZJk5KRK20v7A7XwphqV4vI1XtoMtaMb1i6ce93/tMCXAPjAzL+DWz2Wr
LziFIBHWarVGOzPPPFUsmQjiVgL8VxJCdMPpJ8uMxy3q5aeMTZzPIEFbm01FBnXz
WLgi+2zsLGZn6FtcyO4MvY/SgHf6o/1I1+qePOYZ2NKJCNY5HBBMXWU1WLPGJxSI
ajPVyYsfXob74FEwRf22vlwLp1QS0Ye4/hfLSmTLyQaWW5of/fNdtESm+0PgPVWd
82uraI7K4hd5E3cDKUqjbWSS0wgF9hoJb5duA7LyQY/5o6GkcGAsyQXIqBB3VxRf
2r63TwTfy3svFl3ldVQ6dGFLMKGe3iJhUlBnelColLIOE8h9lSsnVt3qyRzfEOWd
UKIt4NNEed9XHiLnCOAink6viiOfXpae+bHXY8+swH+gR5YEVD0vIYd74UIzongh
fu5yZC5XL66OnvpVCpz5BwVxrBmTfmGk0WIvdmqkkt1ffa04A29bmGDnVNxzNaPj
WJwgPxgHidHtum5SKA65hMJe0LYev6mJkgXB9DhvQSYJFXuqcz52b84jITr9hc0b
wz3JliBZEbiPChj4i4QgzM0ReyMreYJWxzPzhoNsJxBTeSLJWRhPJn8Cxrl9SKL4
CXneSRdjaoSJVFtxdxPkHN4kZhhWIThqzT6lyhAn8MFYaAw4oe5ZQeCh/9r4b4/U
BE64ynF9l+mKuZG1bz+eln7vuPMT47E+K/th94NEkVFGVVpZaovPaxclGTmKSgzZ
vZfns3qKzBs69TMP/FVoKJzVuZm3EcoO4tQ5wjoCKhN8uawuxFLdtaFC8NOrnFg9
OYRrSBdRYFp9iTc3G1P5G0sxy1ETmZVgWcD+ZPiZ2QvN9Wu/wevVmtqXcvj0QIg2
4EsgbmHLlHoKXN5zvoZl47nyNSkpbP9OKGtRrJj9uez5DPS2Kvqi91qeov5s2QwH
/vWhHtG8IJrggJpa3aZmkwgyjJFYBg9WJqqk89nGuOgLzQRbgM8cqhAmQMELBTz7
pQBjWiP0zwm1u6rZx6yN6N+ZBKv0+9KqKVmdBeymx0eHV9ntAPnphAxc3MceeE8R
yTYRrDYwUEg9jHrUIQj6gz/14Wu5B4ok9tq83lY8CJhfed6Qn6OnxzniBIOxPWOW
f05lwIZ5LXVYfxZQp/7WwSmYwL9jdmtwKfx1sh2cdd9lb906avPv59gqA388Yi1X
jaehjsRnx0qPro00+SoV31zSbF/pad3mzLHFH1ArUelJrE0/akZeBSL+yNX6KL09
Ev4TlcQqpKBr5mEVxzpPHUNoLRb9vIK1+f7UWGcYL3X97zjTsMVZ/mcTZobZ00cN
KkA+qqlPXuE7+DQAXTyLSsB5YkmGvRFiCiOcWpDJiw2gQfJXsQABzFfcew5zN4yv
hzrydrUlR7mL72h1P3oz+W0cZwqKH6tYFM8yCcpDYYdQ8+MJMFtV9rXT89MWn15S
DPWcCQ+is06VwHGrT7YjR/gJUxTgyFuJ395CtP0zeAR6uY2HdtVDfdTHkJzR9uGX
otSXtAs2C5uINerIMealmcbyrSGqMucnEsZ6JKD5rmjuO5IyAHk6h/JxL25gksPQ
fN/mhLxbQVXNGNHUoBII2LpLoVeRaaJR4y6RIllXG6SKO6JMntUL/i0gG5y00M8B
cSREOpQkF8ms26UT62tHDQRogWnrVid/x3dR3VLPyWF/VkrY6YTHYke3RPAd+/nW
Pf5wCmxOmHWsqwHYqJQv59MXWMIHsZpwmbC2zUiEZcf/27yzB995PxBTBNb0U/zt
15+dliPCYXl0wFza+sgLf8RQOZC+qqi4BGLKC9Rjn9HAUqYqt3TQ21yggdqUjEX9
6u1tSl+TYhjTNXjM/+JWGEwUIRDuAHtlTnHDNYMd438jccJEQGG6JFLaREwgcLYI
3/ylcbSO3f95CKJthgk/hxuQIsin5tD9pwX8W0/3YE7NqzGSOMAALh7wD7EGKmg+
huplEi769oCiewqR86Gxu8+voWOKHBN2pvz749uv7KApkYmMn2/J66BM0PNfM/DP
UhJ+nclJpRgTr/HIM6zvRwU4dli1v7TS1ks89/hmWbxhab6GUZeLg7IAKJhCPJRe
YKdiMIEzkpLxJLckTckEir/5y+EubIkzj7QyUPiNFEf9TUGLli4x7RsJIFRGltZr
Rw5MrHCfSNjSD+6u+9hi60W8oTFfGDfE1mLvv+3UCli5/E0zfJxWwK3vA4wH4KxG
HNDkLMz0ozChlfN5EUIFrNZ01c5PR1zAehTJJRxWY9p8HLdJk+KjJMymF8Kwj76P
67qqKGsEveyl9+E5bfEX5JHQ/HxBC6dF9DLdmfA0xJm25kjH6uMVsJ6ZNPRQFlC+
fS/VgRKq/QoUgWUe5IQs8KEHGPtmYEHFEm4mHa9+tPn30mdlf+24aLLWPU4vi1JF
t+GleH7z4UEyGAFW0L64EC8ASxbx21UiTzbOgfg/gKfJDBuVQ8/vBzA03GHz56Ql
3KL4OcQ9B2aRQwHFQSu8/lHRskXPJxJ5CCNHbVptbG5pLARm2O2iAwUznYt66of3
E2egJrlf8NwWE9deIQNwZIwjDtZhOaZjeHAVcfUPLMKEEX+7ht5tmNX6CByHN/zj
IM00giqgKJAN7DlQP89xUscx5A70wiT9XmS0iJqD6dc/N5vi8TovNOb+xlQJXL6R
z5shxMnj2aYgTBg356pADTdDJWxpIvFOPwdJRTkP087SH2JDaiNqgCNHUR7C8BoG
IqW2JlLiedyzljniaGSTTrhYj3CZr8t3RMRGixRlnGCGBY4kE8YLaL4qFoNycsc+
w99MTyeUT3ps0YkHdAyQSvv7IIc+ar8yUnZAYztWlGof85O3h/EkXeUJ9e2r5Qx9
PkPwWZIzbIer4ycZzVL/tigNM8UE/FND0DwPIhiqllBtMZT8hbU5zp+nyFPj30PQ
LHvfyyLN36mCgbZv1WPyzdqjapNSIWXTSQWfB819Sx/2W+XU3fTDXFD0D1FdGII8
1jgHzeAhu54uMyAXJD/gA/qylQcd0/CtGimFV+7sqmrySA7S6xKpLIZnyhIYnqB/
LkJ+dddwrBX8SXy1FjYxpDCYDF5yIqE99G2DDpfdxk0RtBmpKx8qguUVFz5Opfeh
0l/p5aqj9izcs368zv7sHfpJl7qWni+nLarZ5MIsS/LWEpxDMXbtNtEBnQfGoQNy
rR65wAvQkVi/+0CvmayWPUiwl4g6Y6BKx36CahKTHcohiAxEOZzsmhCchg7hH6hF
Dj4N59LJWXu2CpS4p+JPby3or+Ow6MZpnFmkmCL099KuPt8JBKmZsOl7nS4zc4OI
jY+1TPqDwqUu1iYdrKDxkMW37q0eWkRV3mwfvk7ZBpCp8Z7Q1jAfeAoiBShprCeg
+Ck1ldihInED7XCTpY1zrP+boD6FH2ZDtNNNwB73vg3cfQQeDxzMo5pNG13zH2vy
k9rHV3Psl8GVcQOCF4vo5kXoZ8Pbi95JMKxyJeOpGC5oyhKaK6BrkU5NO7FRk8As
6H0afHtZ6RrTXkns4gb1q/a6krC+sG+w7WnSrEmlxE9SuwrEcTZraYAHTeUinSGo
PU4aE/9mWRDInwzyn7AlumW686Sv0N+SOA4ax6dR0Ciw5G7nV4iUjYz/GehamyIw
YHYE4+8YGNsZtd7++7Udn4mGVKLpzw4LBvrfitqYIDZvTJe0j8qmjEj4e0r1NAOA
GtzVh8JNLUeItyfk4SxDgSwASRykKYi52I1a48FkslOTXRrsXIIr/vuEIOCubJuq
FtlaNJs3atdbI6n6Zv5r5+t7ked2QF4m72bcBWYe9qul46QV2lDRLA58aHc2/zz+
iFLu3NqPUfeSgwM7MXcsS55omhcpQS4VwbTnVGHZCCa2gme5BXHloznek4n86C52
cPqWUi+HGTaVBBQq5TLwCXI2LUfKKpfz2ITPgnNIgp04Y2wr9sb/E2GmnBy254qu
st7ixEcc1S1ydqQ3EStkpLARDaG4ylz2hmNoMJ2WeuPFY73pjLBtXcg03YSyX774
/g0VcECw1lIA/23xt/hEcujQD8Teiy0Ee5V6ZcrAcMOpzX3+bciRUERKbNJoA7C+
vlVrtK4r4Y1k/8T6YxKWLArCEDBtZIpKBm/g6KVIGT4=
`protect END_PROTECTED
