`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4PTyd8h5tDjgMNPg/lnXZN2Pp5ErpLxONOlSrObVbBx//g+Ms00eKH3SMb9RhHgN
GLkmx+AkrihNrV6kwfv0db0pDlXpuu0IoV6ckXDDIeOjfowsBO9fBHJ6DHfeidv5
si23LAmaCh7EOkgelos/aBBELuUuWLjCmZqYOxQtWRXz5ZxyUEeri2ZT+hbCtpVf
6JDWfxZ/cuHbrmWGEdInsBVduXGk/Q4Ovb45uZtAhqTqGEPyJXgiRd4xXe7L8Ndb
TdO8MCAuSw5DHVpe1WRfHi7AEiYMifdI59baVLXMSmSI2UdvXU25QmkSFT9BTJyO
JiX7dAA+yR6wQD00rpbn9SSOgt29iYkVlcakdbrGLsA67dyzSzVQGUIrNKkpN6vn
tPYogypwDP68ejpZXMmQh09FfoKk6yzwnC7HWesaTGyvX/fw8WSi9ZvauGj7QYt7
/k8Af/91LzjRFPzxeKyUW8ZFVoidvI/+3MztuuE7UepJ7qpG3ZBl+GGYOHPuYWJY
TU/LsgaYBbKIVf4wt1PRv5IZLkyHwBjbbEhwE0jprJwOVr6c2ET5+saONVRXcuO1
S66LhvwAmFyR28HVWj6FtggxlqWYThVuRMBc/ffINhxIl8dFDRe4S6g1vCvF6nSW
8ZCrFvn8pXy0WpP9zUlaW/LGNRy1yPjVIcICMrofVYS9ScjlwmZIPprJGxvHoh4M
ACqxnra+vS5YHbD+AxVVQrM/Ce2iYRmdbB0cfNhPwVPQyZpmCW8RPjHFX9ikbig7
sMB87PG55DZlg29dbhwcvfl7Y5MROWNjFDr1Vbu48gakARvcZlUZC0Rlid49dJ4Z
GZuYPcbjnlRFN2kA1rEvAONQGWlUHRbLukzRDOOQ7Yx42+HaHNQbui5x2sHDVe/b
`protect END_PROTECTED
