`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1N0OVcaYy6vw5JZAZ4YAxb5YLpPMcp0IZ1jAhIATFVoQf7uqdrjlzOqZUWqrFbTE
DCk84syVkWobMkgjB59DwCnNElGqp+6q4sYii/Trji34v1bagXfoXI2xpqxfyl1k
N7W3RMIJLh2quww3psCVQdgzcUgsTYsPwu2aoyC9cmA0YUy41gS9VrOq5aUrDJqP
6zUgx/oR/Y/rt58IT+pWbl2Atpo0CmbPnDRM3fmzGaiFBMVIUEqx1Nbx4NYJMH0f
SpIGWpghCQ7/Vb0e2iQPYxyeJwLXbZzsRHaV0YmOobzf30tK2l3y2XAVTuURThTC
g1/jCfhn4UeQ/ka6EikAmn2h+i5UwqRxI/X7pzGptkK7eT5dvQv5/vhtiG719WbG
JJow9YzLy/6D1UVXDPbHGzYAOFF6rXN87+sH9DaTWe5J8YsQnGXXu9zb/VpiA1mI
vTBSC0HfJuSRdbypwvJk6O76gGdK8PhotggdSaEEpImGq5JP0Y8DP62jwy74rgoQ
ue2NprrfLrYll0Gbx+N5In3AcuFlIIu0kxNSTGbFdDcg505k5opHkGZdIB8ybnXm
Ob6jvr9E1ftIqpkEddTipZ7f+E8fjHbWxrV57yQPJzOfRgqNzh4Q1ExFXSN8pYBj
Eq1yeiYyKHoO72x3cCtAaxtlnTIi29kLvgKyg3iQmiJlAWA46qsMX7noUGac/mTN
XfmNqDYnTOfp/mzfO5hJhW91LNRF+fkkvCyq/dHdGRmHLNuHZPMMZ4osI97cQ/sF
cI01+4NhcxkmyBDmqETF1C0bX5usjK/1BB65n7f29tsjOBHw6PocJyvVx2752sfr
4joEALgeyRNl7agSsSDtON+T149w9a94xIwcttsUqydRurXYpuLCvmaTBXDpl+lT
zk55XvPn67gC/Fn3Z9dabyJTSqMS+MiLIRhC9NsN+EfG7KCZHX1nuKiVRoE8+N3M
diaupsyI8M7LjnBcQqvt1l3DuA3cNDM4ZRZ/irdWaPh2FT9IeyJA2rNV1I6Dv5x3
I3Rn5WKmrSbjhmNO6wXmOsBTw3df4H0Z9Ap6mYYEOLGgPJnKI1jmg51yekPEgpFu
mZJs1eXFQWBOD4FE2/6Ux3GFBqopO5xrz06eRo0k+Es/eLjxw28uPq9fCc2H5TNF
`protect END_PROTECTED
