`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hWcYuNuUv2Lp8XdmfOiAKxWAnrcfJ/fWFogNnEOyr5pcqPegN4O8zwacJJ+rDnSJ
K/HqNgZ2jNdf/aYxvj75mnJZsYFjEvpOYWPxDmMmhLjJY5wLjGOhuw+UXPuprNiw
tfHJ8XPHp6OO0+52p+jfglAjbBMj/8embmttru3GMSlWBPNbx2OMfpi7x2MX98iH
sTSiNCIHgcbQiKjhyoksLLaBYRzLGRA9d7UyZWsdxaf69coqsCH2/OFTk3gNA/Hd
xLcdymbvBsbOgOnuGmiwAzxgvhLwvx7R3xfmhugXA0gNqbmjAzXxPqVMQZfLsQdH
B99ipsQoNj6Akb6mpldWa3kg3qYQvwyeITYll8juBtnBKiy0ujAZBdjwhgIYcoHW
eAIWt8VHUu8yyiys1KdWigQh8FA5f8WON5zrm9oR/mIKO8Y6sA5Vribgn1oea43N
ijNHNQXR6f4M/+XNOnD8jCc5TAQkLeC8HLmhEBLGX5y1LzOeLFiNkb2B0prYm3YQ
OtrUF5bjKUuchm3r00ZN7BU615mZDngMRyFVVqrwwmO6NdIS3NfUJg4TCKseFEQq
4qD+tLcG4h6Q4glsce6HPzQCMaaJoebBXpoNMuJ5jGMdQYvvIW5WzmS8m+VKi/FM
xGmYc3QBZsL77/loVySaZ2QQxTC3Q0qDqPAWbnrm2sqGsuWRN3Txi8G7ZYqjBqIJ
GaADAIFc0TMibAuStcGCK9TRbabX45dQJmLrUXjWb9lI3tadFbH1a6L0Y3YdWI5H
gAvWStUWLoWacAvXNOzzwz9czgzHyqMiZGTFZNZ54RsyzlqdNEkrLadbrd/ABIrb
k3NYagO6JZ7nJndF2GrEvNA97qtjc78dAzMUoIjv07n09s87wjR3zZiAeCrJ59Z6
H9RqFgjpLZyuW0GhiTMHstdNz1+lr9LyR855Q7v7LCnI4vbFQ/zdMz1tincB996u
IEb7UM5J4fHBt76nt+AVOMjw3CxcTaJe5fK6wGYK/S4KoWuQSSLUGoX0HMaNmPg8
rShYbpjYC2+u8R16LYkpYKRgC/FHrPaba4ychNASJDB4SJ/aeI0plRWERQFUhVY9
4GE91RNFmEcAUHKUtFpMjab7kz/dRFauVADp09dYuEjbAVdq4jvQXRL0gzBNpyfV
fW07CXhOs6ThuMBudAvWIZ2d199JeyPCxJboLS65WMri06DXYruqdZ/yaoQZE5tT
cN1KzeFIV4L+hJjWOpuzebwQMkhvv0KZO93kqcIFxfB7hOn/aax+G99MKkuVqCKs
KbxEWtwEqgsyP+mdl8R0de+Aooa3bR2nImvkwXMwYEySYl9eJ5TqWAL79/hWp/D0
VQAMGgb4e4vR4B0hI5cfTftTryPeNJ8JzCk3NIMNQmpEfOtKvHqmNMVo/HSFuRvJ
kWP4olXXvLGOHO2W3n7Jdx+7WxtpfNP/f4b+5XB2JT7KNnUod8TaQcUgjIY85c8E
qkg8xXnVJ0bvq5hVufENqaTLeXa564NBf5ur968UBcem75kVW8Og5SfidICGxbQn
tXA6Ym+qQjAdI5+JCpBacStCF/vGRrrNvMaaoOCuMDisw62ZOBkXvttU18BfYZI4
9edJw9XgbhH3GdEPYjFtB4o/ubeVCCiyac7zsCD+fuAPg+dP7MpNOgFNIe/6TI3C
x0MfKtK62ZszR7/c14ON7VHaKN/TfbXNF9Y5xWgPkfUB8CVEkheTbDjbhXRvb5qF
brWSOIitAXY9NGP9qc2/nuGpyjD0QOrqV3N23DGhQn8xVyteQNN9Jk9LwONLahdk
9SiYKJ5AcNqKB5vhW5wJqOR8KfsaATaEtus3Gc7fd4e6JsoaExlQy1vU0edyJ4YA
o430sgH+ZBqbF0tnIOK8SmESaUYSmDrlN7WEgPrIcls1erBTCKFYfYeRxXzCUHCX
JqhpxJ5dTp9qA+DJkeerLQ==
`protect END_PROTECTED
