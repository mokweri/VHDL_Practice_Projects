`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXOV6enEBQzy9KEOTDWMd1/DYR+2dAQGDQ08s4uhX7o+TaCJqRFLw0WvDkJ4oFKy
KjZQAdYsizTziALEo0oyVI/5pbKGcmbqNxDt7JJRdtPgdyHvUX3wtpjH167hCsyk
jX7+W9paUJ4fCFMT8kaeF75qECyt9TLvI/LVq2YpEk36UYVFaKfhZU2u58junUIv
kmsLti9AE0c4BvfZ5Nj+t3K5tmBu5yMA59f9hIsT7/EKBay8PqLodf0zd8rv2zRG
4Zq+I/Q2hvRDprWykqDXxalwrdYx43/fhaXYhYcwS2PxqjGJBwg7m2Cp8OQJyIly
GMA2mQxPPkLf4il7IG4LeKEb4m2P0eInfpLX8rV43YoYF+yLO1T5oCOizOAO1LAe
a/sDuw/j55jRNkvhBBJfpvcRMlD2+mcNIoWYj/i+L1LVVr0QkGqsrH9Si3wW+2wM
wXXXD9+mKfur4gRlap40pu5aimQi98oT4jyOoz30w9Yimg5aFlmVX7nIClSmPmpp
dyEFGgw//sVsmbP7NKrgHcQrelbMM4eWyq5/Vpq/0aMl/u/acUQ1wHsokmEPbdG6
L8yerwmMKrgMJ+mnwgfYYpMvwC7lncmRWWYDKrw1j2GbTsZWN/e9co2VN331lfws
a+/dlXEDseecdIIZbgHsCMT6J/rFyjRkyT8G60ijxIoFjXAiHhDaS3jnjtNrUbHc
ef6Y2Y9SpoLlPhxzDuqkZ1F/A3RPis3njfPQJs/kRjT5toWbuwO6Vy7MWbvKIXub
/sp7GF297IRU3zU9n3jpfjnCdaLhxxq5yNqaNN1ChffQ0gjduOzHoFf4eWY7V218
vtH5WakNT9BOkqosuf+ZVSQEI/HaGy5wT0SBBJNxcEeaeUYtTQ8ZhN/EMq+qu61Y
i/ZoGfwijOfEo6gftfE7utYdA7ieHfxsPermIp/T/7WSXlMfhFdr7EGDhzgvsBmb
vEmsKtbibmJWtFXnUMbFPPByB8+Jk8oWfstNsagbetD8FCcWKrZOAKjRuk1t24jx
6px0+4jYDhQMlynzzVsa5GovNfeSaZTE1WpaKAsE1y312pIxvOSqFzv6LiXO1VCF
qsmiHBJd6Z5MNl92F0+WSGf2xRYbesxLDUPmQA/Fgurr8fiGl4WoZ10/VaoJW5Td
/heovu9yB6C5W1znt6FpKeN9+ZPnD+kVayS0bmjRjnhIuf6qCOoSuero5iItNPUi
Z51fsQvEYLZBX//1Zug+J1rgW3AEhNFxuDM8h22JoDAsU8nkZYtl3bMuHRn68JS3
a/7BkvwrgCB4W5d1DQNXrMInsadpyUvZs+ULiFKlgaLowfxtARPSxXPh8EKHdgtK
V1/uoNzbMC/kOTlvUBX1zGPsf45iYoG4jchsieAxmDMeP08AWC9N7lwW1ifBQNdo
UilNfxVAIGDdldu5RSwd7SoQSWI2a8drqNnOzF1ziaNuPQlO/EgL5xKkm7XFGPnt
Y2FOJjZih2BZ/Ddf4IzVlpsm3jp2brQG+4pdM31vEw+lUVqK9tB31AmnaWdmqcoL
Qfjo8fAb7ENR0uHM8ssk6m0tN5tYalN5ZHdbPu6cUlmFQlSFFDxIAdnopA5CpsjO
uYLNdxXn3mVVJZfyCCOr60ED4ajeWS76mgsMSDlEKrL9syFnhxNDB/KjSnsAHHJ3
swrGisuwU093CSmn9devHABBcDOvNC63aCJdo8PyCWxdQMzjquKIPpAcE9NqY8Th
4mk9F2oFtuMSjMXPT36hz/umdoMvXB1UWJBjxUEjerL4rbfIE/s4RXwiRtJXYb/t
PGCnTN4/+zJYPB+RDa1Ft9fRdYq1zyzpUvqCazWHqE1XuFOzMeireXKF1KaVkgqP
tYsaD53/UH8kQZCKtnXC0g25OHlCCAIl2MbMGYIFORGpe/NJA6r7/QuljwTTTvum
gqEC+AIagHHJ6fEJ6HDNPbcXcK+rkepVOPW+f9EW51cWxcL0AGFvRsM8jaSY5GNV
TwGRBntAYRhob28EmxKn1Im6XqoV3MCUdvcdP2swYPq1NGplzDrV9cKZTGHnhm08
KdCC+hoANhM2gevPPZMfCx9wNiDql0jrg7FA4IOfTFvR3XS7TMDBivfr1cOMUyPW
FvgBGUbDvX5bEj8IUJ7dBv9UcGMxf0vz6YzxklCKpuoH4ls77y4NPHG5b+zNVOVz
kG9ZdiTLvsJV4SxW4+j3pRwLbvgln6WIxdqamnBSFcuY7CZsFb5+QZ9Re9tlkLMS
JC4OmM3jzScgwyL3VLyGbf5fzyS87DbW95ULzNM7lNtXx2cdhOPCQN6BSGa4tOtj
lOwsEhWjqRVbC5/YvTYIYhYr2T6ySXNW/MBKE7TbWm5fxH38VQ+eQPLXRZa7rIeR
2PwNB6mzNuCjxlCSfIjSoUH1tiojU25U5/nkX6F83mbWHRIG0nTg5lyNeXIzr2wd
UiL21twyr18w+RzXDulsD6M/Dn2CaHjmmZf6OgqtvGgOjcKiPU/HTTnCbn0JqGbj
mJVtkEwx95cierQAVaG6xEERLiAprIsemh/hpYjs74yuFPN8oLjdSZCcmrDlwHUb
NAgnW1ph3830tUgT5ArJnADD+WrCMEk9Bhr4jVItHVSZHa+2Qi89L2DcXY/MlZNP
NKaFbR/7A69GKKq8HYdaJwEPN+xhGhQU9dbvR5/uzE7qwAkTB+z+hRSSvzJYmQL/
A4ao3XqSUdZyVBWEISzN8T3xUj1I+TSUHxCaVht7ke1lcNDXFRIcUYMLy8rg0BVv
F9ezkJmk9QJR+1Jqzl6FYOzyhmjyaKnO1zY7efU4hkqpIUjCrcfNrXsnTu9fnarV
+9imfP4rmxI+j8wOM8s9QHWkzJGmzpxbk2/2ykvLrs7sOptQkeiig1//y57V9mkz
0E676gJEHaoQi8gNP0TTvcaI6Ik7NX+2oneWS43WFm//sjOWAUlsbX291DVZtPaE
mOXrLQbsldwcXtr/C3wBmQMqjzgfYQwl+3tuq+HvRCewD0mqB+9ACbzZWZNgpC4m
vUKIdtx/J84C1FTtpCYE7oLTB/X59AWS+wWc3np1RL263GBfFHOboDDbJ208L91P
lBNQxK1hhEHSyhq/vv2mgtkIfH0CdjPq8Ds56fm6mE6G+QhkQDhAiX5gLgv/hIkI
D42QeBw0J+vH/hmddCpvpT/h2L8MbvqrpL1fcjZ1uYgwZ6pA3L+21PjimwjcZbG1
8VrA9QXYCKtJ7+c7tu9z2CQaFGrqzw6ZYRVFb9xp6Eo8Ofovqm7+0/K0nBmH/PY2
ojr5AXxXwStG3CV54Zbvg1o5PGC3IexEAbTiaaaHQUU0rTmsYVeIU4Q0fUbrBPgN
f7bP2PD14PmTqE2gMAZqmQph4RcsTk/PQIsll9+F8zSCwj9NWIpb61WUPa4cz7ms
yynY8mpLeGJjb0ZtP73NPcRW2TlDMXmeSMsFhUiXOI3r0fHsxWUvn0aPH7UXVKy2
Yb/QZD6tuw2haQiulVJHdICc2/SuQ7dRlnjDLF7XWcWNWwp37HR8n92upNlFIsMn
y9jMOwsAQ3+o36UqxYm2s7lUTirGqJV/DwQUyZiUEGxg8frLZ0blLibdX/nrLmLN
v8y+Iqj+LLBEI3HZWUzmrMyme1lkOm8obs6FcvCty/Zpl0IfnVdniQ0JIfKvgXhB
SvneOGUIGZ+TA9bl2/iLc/rJA/asIh+tJ1ghRYAP1AiNcolDksvTXhztYWyp9L2v
6tq+q7nhBZrxA07/IhM1fWu7+DOiObzesbZdMUPRLnhIP/7R/WXHiTxWxVPUYMfr
/DU8dV29vGFvGOyJALu8RnruSxKHH4Gu/iYexqfFJ1Vgb4zt8PvDOjVRrthihLH6
Osi+OabUqIQztDr0WS65+CMO08R4uvNCwbkFYrHJ1rpk7qc7fl8z2aqvezO3cb1y
kjCIyNbzBOImqUsF42J4laXgncNR2Qv2QbmOASUJbr48L+FQyR7ByM2XXe9DMQ2v
wTlCG9I0g7PE/lJnScXFTEsfbURAxhaY7Oj6fVVZFuKPRh2/KIB02m+RDSZ8acIf
XUii1DFEP9C0GNDQolatGAu3mVzgOfFl2cJ8/m2Fh7rAjDxg1KLlr8xOzfxvTlE6
P+8i5oaOALzukxnpQGbPKQIMHF23zDQ3bBSMR3uuic3+uke7XfOQLGbEeHg7dGo7
ca0Nw+PUE5mRYwtij1K8Iw9BKquI4Sz36mij251bDAkLYPXTImNz+1GNUFnkeb3Q
OMiCeMFuZDHQL/MbEI9aD9Z5446eFTMsLkdcisyUVkhgH3MqeRXc36uUHzicPqId
rEKCb9NC4hCLQLSFz/jdwR7tPIL6oAV9zmw7TUthz1CUwtD7rQFkbHyE067eM7ur
ujXdL9HAdUwZ/0ejNhOiMCaqNk1llWexXCzInjLW2cvh+U6eOKOzhNmZNauJyNjr
G8pRJHQjrCSHMcUFj34zg8G9wvOn8r+7pvQ9eTn92+z0ilfUAJb1yu99GaMsVz2s
okH+QUepijT7U5j11xh+ZVDUbF7XmV6aTZhnz67yxEUgHF44uUNRXIK8kSi8H3Dh
uNTIc0fw3RiNo/jVYk9+IQpfCx7RBiQqqfFPmtaEKADdExBm7LPfcqw3iMkeJn0N
`protect END_PROTECTED
