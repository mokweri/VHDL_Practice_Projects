`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a0of+buI/LUPtXBr247Yx04CqLPnf0cp3u/cOqONVgD9PvAZNCjlXKcD7vtfZLhW
U8j7OfHBca/An+LTsDvZzDQSsQ1Sf7cPlqsCqJcaZ+TiOXhvbv/tLbbWKScJum2U
SfdMm/M9PkzMPBgYVNkzBkzXuMHuXolnWRJcTaQucP+l4eNcUPzGDGGcqOmu9UNR
hXADhJPbTZv4l136tgEIi2f08gT+jKzQKOPDDfguN5WaTna1Y/wYgMc/uhFYWBYL
Bes5/rlm0X+BuyVF5QmBYCgyTSMb3t+3UW0w6i+OZHtSCreokzUuwkR6Ofl3ajji
6NYj6aWkkXIr/29QwmP2K++ijcaMT5jux9e/CZst/oJMeaTS3yjSfyir9JQaBqYN
w8NCUCHIftm4nCV9xm2ZnXQQDrFPzBfDqv3Yrzkc/jPf4459GAc3yyAFZ63vdUCi
4YoA9sMLMlDRqij+9tSJcMjchIhio5hMuLcmkVF2XvKKJEkkPNIsD5Lrf/AM4xv5
dSEgAk31NttXcQDIl49CbxXuj+9EMGJ+4zDUcqbXLWVnC3GnMJ5wJEIVSl3P1E52
8MAHuLO2mpPc6nEwINO1XaRV4w5zAFU4g3pKF2WHP3EdHeYtrnXMVec6rmr1Wx98
79WLzjWfOj6TMYeLCYdA8iLgpDfmte+WPyPFZWu2HqPXj78qZwnBHn7EnKFhqMtR
`protect END_PROTECTED
