`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eE2QwWKHSoICr5OEYhImXd0neg/NuUtlCyKD4eFZtzkYHd6QKrX2YEnY6u9+pUnv
vA0sgZdcHc9DTVYcFcEUQ68e7DlAGJokzQNzc2ydHDtcoxol3lwIp8+wosFGG2Ry
SaYkvO9FkeW3cmbrSUw6chntCwtEahVkhzzybJqLRj6maLXbPd6Q0VXpx+zVDHIM
QuCLyfkmAh9CGVmaXJUL7vSWbC6QQMP7BtZF5U92oPb60dhCVBuSIXqbwQyTpMom
wR4JhOCwfxKMeurruwLibSTjg+W0ZVLSHWA+8VJBobjxnypZyWk6WzTaChCxt2Tt
kee/KoiKWed3acKJOQxRuR4lVssoyrwOSvUp3yDixza9Jy5ykSGCWPu90q7Yft4O
utD/L37TnqAS2zajcnHkLVSjXejD8T6GsSOQmhpobEZfs2QnTVq8P7Fvmi6gMQYY
oSo5Ozd7md17DglXwNQGB5jQwHQwWvL1tE1L3+/E/o/0ktTBEMRh6jVthlcEULWX
bIbP4N8qax4B5zwiXoxTTM4T+s9Iya2OfVX/AP/1pjHa3nfkmc83HyN+l699UHr9
cDTOPBcqYlXugeiMEJYdlpk89ZcWVCjCFvkw/BY2TJWe0Ty3gzqXcyztFLTLj8J6
ZayvsYMq+QN12xC2EenHqe6xGvb2ov1sFg5G2bD2MVIQR9FWLqm/BPRMsgEK/tUU
i9F4psgParhUcyLhZUo2vVqlC/AqfOkhXPXlWr5KA7Y+4AoQIpsEPhS8D417KW6y
JWPvFffGYat+IaWeVpo2/Eu4mtzMjYE8if/uYBukVaRvpMAkavajkNbeiUGKJNWk
bC+PbE2ch8EY+pFR3s6vXK9GPm/ixu2ozlozHkaKa91mLm30Gtso83bxYsHxrbD1
qQVT/7E8X2x2aRtoY9x750CYjFxMQpx6AOBC76vsFR4G9h7LbxMVYksAAh48Ghos
6pxBQhGLAjpt0SirfiNfqvyrdAdBbitukQrlDqBteif4OvfodmT8TFhybM5J31x1
rjpWE/MClGtHOS2lcdodMDraQzTMvl59a5SDsUVD2gnTPnpOfAOiOKdXRM/MwCW5
FMBkTylwpyitQ1Nh0GjRX5+tR6FVi3PPEB24x+E+YV39pPomQ8YuJEtpPHPdsMKO
TrIH6AWCP4Sl+vn0MFM/7hosSDMW0KHE2kqYrXO+nGD0aaXn/GlSCuEDyChr0td7
XznmIEF4CypE/JKa7YJA1w==
`protect END_PROTECTED
