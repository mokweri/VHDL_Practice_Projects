`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFhWbQF0GOEB/OhCFsxoPKvHwp3Y/HaZhARSqBERSFCMKZtu4pYwhiy7HFiZZgZP
Bb8eP8/fQVJgqQT+s14ClfhXSFgQC8NieccDoTv1VFXBkQo8plX7+fltQTCWiIAN
U9ISpTnkkB5BY6kFHsg7U7EPi7PfpcVxNtqn2biuPUMPOYS2OzA0USjqoZ8szGPA
aZ/NANagpwn8e4/YAGTaqkwSqVI+Zpmu5nblqvioueKO2DoD9E1j050oHyjHRwi6
lTKPUUjZIb92aeI8yfYwYcjtaoeB0Vxnby928G1tGLWRb1xdKfiBc9L4lfI91n+h
freeDSYcA/gnMmOXU8np4f4qQtpuVKNaz6p5XWduCOvqped5HNjbcd6frkqtKPac
fqi8e0qh4ReacDuIwsEDBHpj+JH+8eYg19C3iiSpITJo7pybUvR6n8juaxhMwK7z
xEboUoEiynshkryUCwN0QooX6eI+QS9ilTgf5Twcvg9yOHpLti3dvrxZuQwAsTBH
Ik+Oa1sR6IYcPre6Qi+c3ms4BkxVswsTlss9WnDQ/WMBj/iXqV3DaELe9FKI5xiD
ZNLAGzzpofRKKLLzSRs6Xonluaycr1gAMOsMXHR/CJN1nMNi6punBOYne1niHpbc
hvswDfFHSdABnCmdZxMJ60rFQYl1WjMEleWfOkweNKTwBKb74bNqmPsMg6FWusty
6K2RxiVvieETPqumsxzG+o9ErcYNn8FUHKzytox3taqtcufEmuhRxmuGqaI74PK9
dtuZL9JTNUfJmDa/z6D0WHCQKcvbvei+WYt5WvhHOf7jld/HUOJqxX+cQYMKdRZC
L41BGOHKf2IIz11Dko1nz8lg25ttGxfUNKj+h0xVaRww2vuH6yeHgL6Rr53Eawnn
G26QjzVTsLsExifBBJuaTzw4yx9dd7OSB1xyjiraMj7JOLs+8wrBNSjE/nzu5xNa
z9I24jROM6M6DQjfZzGP8AtsGRczUU64LApwfj4DLgnpo2E9dKDwiUZR1AarJVvu
11ioK1zchE9SCToDQ7lpPWXRcQdPf0iyDp5ak9ASgd5ZM7TdWz2ovaOUDq4/03Ah
zYf9xL/P4s7GXsmDzmZigx4ZNmlIUA6ediF5w9hF1kW954oL00hrc4smoeNkoHJS
+98x3Fc9pE64iE2snRyFg4uAIVlRcjdVOYyK54b3Azgx8B/MbOIzNDIC4osjPFxU
mvZv5rpz6XZIYLkNT+HtkPu6/dMhbsrRCCNzo3fPhYUn44XJFf3CSS8mIPZCgJho
qQf1NVxuk0UyheemN6hRuNNsE4QPSIj5OW3urn9rHIHyaIsQ4LO46zuBwgCbVuZ0
EanAqI+6Pcbc7+GrxGgd02a2qpvkjOspCfB8YUxCw1+tMmStgrwZGy/BDtgMgv+n
SpwHXqR9RbaG+GdXDiti8jFHabWqfRk2ji9Ero8qnT1zv2nxO/YLCDxPFkmvnxid
eurRU52P5lPz58E4c7Z4LXvmpYleatipsfp/cORV/ksX5jkxoCZNVgcxayZRjrh9
Dh905N21zuNx2NHnuweoa6XKjs/ZmDapY8+x3NP9j5OT4hfZSdhwSUgNYpUxeX2O
HFOX+h0tUtVOgfDzGszV861lXcfFMrd3q/JhxD44Inw36Kf+jwuUFpF04+ZRNIH0
iaMF2iQe4tsZutRblZAtVO06DEUKuoYXMKuaQG8jfFHXnYKT6zf3Bw0iJADZzk2k
ZmWfZEJ74R4BPK3L/tC3gsYomh964Kf824F2NzPE6d3PspwzZY3kX0cSoojfyMF0
`protect END_PROTECTED
