`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yYRcDrFq0AnzfFr42Ht5O/CFjh+pYg1fRCIaFm67oSJGnuvo+iq4f9HxFzMQJlPj
y80NRzCJ4W4VH8b81dF9aPnrdSGytsnPccsYrYVXKUy5loZVuGZ3ATiXJCEsXZdr
X22WFVMGsFFu0eksduihAPNiKzWWXGVLUYBr4zkudABmOBvUxEs8U3XZUiBbOrux
q0/ZQHpn4+ABMJ6JtVB8bM4iWikzWExk4JIWD/Z06o/c7DW3YRMyUaTDffdwU2l7
xt7W/kU+tcT9+xbyOhBxUd7/qfHINA5nfwvftr3P7dUL/qvQZTnb8ggYjE47GFGx
05jYzGaFZ1M4a0nPAnowiBARneIGaCldqMw8SoZ3vKy4oKEDFsD/c1aQsrF8460w
hA0T6pAo1QHv2RCwWi1BqGVbVVG4nyCbO/BU6mAjxcMyGg3C+fr31zEKRDaA98rH
XGCxwUivsofXBuR+5mh5hZcMepQHDQCOpKCwAqAgwt4LMwFdL8ZXsUEoTj5oRu04
KdqfSj6UOaMlq2mfBzrEFHV2ibuNgdS3Z2pzFFpv7f2jY/DxAozNrGz04jRzDNpE
O4tw7Jv4UC0sJLxitmUAxHnyuNI2i5rbH+N3mmHQeh5QSVuRNvFo9B/7scy/gTZC
knQZSZXHOa7GobsG1xtFchF0MYqBEupX0WxzNJvOdhLHlk7OdKlfyiwYt3Kj4OsY
GOuBKdFKjTTTuoUWh65OQm5TNSVeP7s7c9zb1CzcErw4pDwCBKWAG3qi/ShL9Q/5
jsXfOWgcf2a2n3exFk4s170nRN/p2Tq3k19nRpDDbvAS5mLWrukeOJm3wW5VkLtf
MmuCZqD2U+sHyVAXv9k4k6L/25vj1lKG82hYiQBeABo2Tcxh2HGrMz52pUpwHZyI
OS44M6plg704noBWsfLgIUWRmOtT+2OyzZIbLHKJuAL3dvo9Og0Z/L1Mb6FHHc0M
ofNz4bTv7x5Tp1k+25PACwNJAAQUxHsf2DLoz1WuFzD1dOrto4yzBHUY3BwccY1g
QdInZ81ax6/gczBXzqnqvtRZkDcdYPk7h5HurFQeFg/DAxKIeOTES166SI/Pm4l0
URDSY+oeW0wmi4iAH6ty75/XSoa8SelI2cR0Un+oqobbla4aZQU4PHFjrsOfLeeP
LzMnIlnIVwFS7tftI7QZQsY2RaPLoyA5r/WAP/ZXbozqRccyWYZIuR4Z+ywah2Sj
37qrfhIun5j4F11MFE8q8L3kQ/+mwoxDxMwlaYEAbYaMnDfxKHRLV2+cvTOetI2m
faGBjbz9SkA6NZYk7ZS09lxXMe7iPKFQePnZLoO1OrP+YyWo4R9VR3AbiKaFZRwy
SgCr2VaHW67kpfwNROjUKNQYrzW374eKpDaSbNfxSc85rBAOIHSJuVG0flevoR2e
nzMqAl3Gj+DXEoFMW3bMzflVfcijqa7sm9AvG048q5XEdU3BDoEWsrW/CFNGeaVe
K5oW8Es6dr+lAfvxeWPEpeQsSN1X8fvI/al2YJNHyrQdNnTAtN9GIfmVWTTeZHcJ
R5eV31kFqr+4sjzmWj46u7oz8fwwuHw89ZZqiXQJmTZdXBhT99eT/f/EI5Fof8pi
224FMRmldw3dV89W7EXundN2CPq0PjHU21VmwcOQZoFtwKHcaAu0I44a/qvswmMG
TDcYQZluTdyoaDtTQW5NLkC2hHz5C2oTCUTBc4TGO+1j6SvvxIi0LOWo2yS7xlbK
ZPCDpgkcQalZSi2TgPbsjp8bZsBrISUiWUUPlAj3x06oU9YyecYw55ABI2gyXa0k
YwFwgYqrTmrEMl++U4n05sRP0c6MdWN3jJQab8Oo9B1My9/NLiLX7BD+/KrY4R5I
6fVqwlL1Oe1GXnjQWT5uIK5cDc80+iUnJERQKNxHekO09N5Ed1I5hR/IBQ1rWX/P
st1G7HaZyFy1eEnGO/nBfvWN7Q9ZvH0JV2eWpJZbKoRrGzZjovAYpRDIbwvVxKtj
bbmmRq5qzAA65E/ZDS7BcPPzCRoPGkEZXP/fxxEFkyD8DJFkKW+lH/ebiHsEPOOh
oNz3BSeqzh6PtYqgQ6tkEU1E3OkOQPYN5XkSXxr/h0KhWQXe+PzLq3h3FnB+vOy1
05u1/9v8jkfhnhoZeWO/DyHhtG7yXgQ4CWBpELd7wGSu4wtgKREOXLYw5H2h4pdp
kR19ecaJq3EsguymA5bwYtQ8iTAXG3iYZuMW8Ot5lONJqrPdrcfNwyJlY8g6JOoa
kPjg472ps4kVI77OmFPGWMMoeaWnsFXBJ8VxGb1LxPSQQdp62QotmYxcaOf890RY
5QIsGmYfx7A/qEyre/kntAc+uNu84hDv3Op/tzqmHk3n+CIYxfGizsK6R+YbxKnL
bsmrj2tMn7YR7eyQEglmFboZAPBg/Lm2NGTaz2hviEESJK9rk8wrOW0NxQBEJEoK
`protect END_PROTECTED
