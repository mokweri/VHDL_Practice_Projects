`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnGkY0+bHMK39NUppkpvUBn7zIys0q1aFmqX2CW49F15LMZ/aoN6uq/YFXetjwr6
bhrU90sgBFfR3pFK1dlS6jtzTT/srsZOiS8AzFle2I2Q7hE2kp9cF1sbyy/RXFVc
ZMgY8oYacpKQgbhjD50GEFKgEgwvt5MKo6Mex0KKk0/crpn9dZ7BQvF3r8n1hhcE
beqLVP0kLfEDEYWi4Lekro0CPf+rjym7fHZKCMBvYqi5S0LmYf5Mv1eSGNOnh57y
vD6bv3vtEuaRqGzltVvp9w1fyi3L+JeoE6ZpEPq8psfid4MyfTx6mpkSk06egS6D
87h5NLT/rukPWocryp5Kw4jOCYGidKSGXo1BbMp/JPfAqnSTXgEMYM62Gx8LnxOu
Q5mTF2RgSLCLLYrpR3OnLWmHhSUm3bRsVjNQwaZru+YxnJh4QN0na3nTwOyuf9Zf
Yx4/vgckuUlqB66JmtlzISAW0W+eELCI+AeW5H77FxsdNCiNe5Olvbg5oUpEq+ij
myi+ChoZh2bWAWb0Gwui9hWKWcOeo59zooWqmSC4iKqOePPNekETuusk8ECwPvKI
A/rr3AnUizI9lyj5mv7ELKpvVhUGR67gOC4Flb/f16qcVfLm7VDUSeGhoaoq20M9
Cuhtnvy8qGcuOlT3Zr1cC62CYh+M/Hs3BZWvb993TZlcnn8hcjfyMho1f5FJFkHR
WEemmPwmSx70otWaOgH2SO14cnR95mO6R8HVUKlxjFGts4it120n9m+zzfCfbM0S
VEqBdOSc1ROWsQzpZq+uGo2Dr4hmpJIuAKo0e1HbXZI1l3u03d7L0fXa/eqssqJr
sMhfy/uQUeZ7dNCTsEcTt6e/wkXObE6I8goVfXkjVYY/ZhjupHlqJ86u+4CgaTY/
3WAJux2ZNRLehvz2rWty426q47jIJs3aM5wEM2iDz7EEPVz4XkRAnkeqmNeS1I9g
19yqqiTihnl7000UDsbvjcz7RE+VOMAEACUqI0pmAaZd9eaF4URrlphSd7o5BXQp
2EXb02wnUP7SSLT42of2SEhA9MRzk+QhB1NIGRAGOUX2waSKr6Grlh8tHWbM8Idm
ek5y9ncdLGhwdXcdSpJbzgsQUQzxvgF5RhWTL80tRjI4EN/tjXMlHVxPbLFj30WK
4FzEr4/dmcf0aHYCTzcovOLYY+qSOtu5b56ltXtACa02Kfidol+W0zf0wDN9bR7v
EAruYIvzy4Iwq50RgOTdBo980czSwiCyP9LaBWPF1HYyPH305z/ViYJFgtfUwL9C
RyYJOeVDS/wW4s6zI7gX4GSUdiGOyqyEMgq95zzA8B1F8JL7ctcIk2/a0/cc0/Xb
2M0jEFcLy1kaVxltKPCYbwvmZEs4L5rF8Q/YlAyRTo+iw+1OVAZq9MJoMn7H/dO0
WsSqJWXJoxH3Z0TPYLdRTUTWDFGbIaV3zujme9essuE9PXKlF39GrueP8j0PZWe/
gf5UdEgRFlV7GHc8YqJFStpaBKbeT4JW5JP70TNRy4dtnMBXNrjsDcUMIh0Svonb
rMjJ8h7nfRZQAzWCKCpeY6YEVnnzI5hIuwh48r8LtDdVGK4VDhfpfHcRUfqv43mP
dDQkF/qsw2OZuCSQpCPxAVLNA7TmJHN82Ldo6qy2NeuiXiTkvTNG9zJurjEDP1WP
t0IzmXx1rhXbf5FgshTQJGBVLbP4azu5IqQNF07L1h8lMZPDUs3n46gSfJ+V8ph7
W6vVCejhCz0WKGrqb7IEjI01ULqLfFhplH6WtxI9vPLmuu4jS9Gw3S9VDFUII6m0
XrdcKyuPYtr83dsmYcEWwND29zSWgCkM581CG1o4h/tc+h/NTHk25AHVXaFDnzT0
MMXrTqmexCSYHTLhQAI1VbeA7ERYwcitgPHBEz+JPYaabhHTl0TmQ+6vHiy9sejg
DgHGlQOHBnlnyHCXZu2s6XaxUiDuIZ/yqTbtxDzDDEqtxvGaIX5REhRIR3pVB8yx
Q3FYAUslemMB4VcJdbPY77roPQVsdC/Yt2D6j58ftc4TZU1cP7FZTsZ5p5AMJPMI
hG6mZC3wk41cuFdDm90SBY2kI4OznrbGl5HT25u35W86Z3MA8SPhI/DgsMEN5Vpk
2FXURrpbRjXReSaqvGUBL59m5IJ6Y3AzIotbAhelI6RcWwp87qpccpoVko0/CY1Q
dbHkaFgPTIk4bw/CUBoicvS+IJBuIgD75KmFU1RtWCrmLtmlgtXxV15N6r5dhqxn
NOK94NxwNqhmj9rUy4eCIKUpRju0WFNp8da4Izva8oU9T3OQAoKmrGzkKVzCqO3O
zp+jEvh5Mn+D9S/RVVnl/GAcwIDhJM95ed8HdsNlvEXdftSzkTvZrDxkVRUpJ+TA
gfkWWjWxyLgVuAzOcQXNB4B/vVoU/8REPdjOW+xXx5EZN0tCMpUjexsu5UZnwhjl
9b7fl1ZBmsAw3kZf3cT0k+uJ30uzIGoSCJ2YYYiu7gtEIz2AiaW6rvUMNj0lwzrs
bMTqKGyALx1u5D9Md3VnQj2P+bnQsCyOvdTnZSQKa1NbjAg8gQYipOqSTPQsd3Ry
QjUs+qAbCa/8I7RkzCbrHb3IMBmSnJX3fikeROmuoDApSsFk5EC8Y7wI97iTcCOH
Uu9pV7KpW1sZHh7x7kLEbuoPAEWyChwkAc084VvqpTqiIUBLq7a5me2qAy/j/qiW
E88AQpX2Af2qwd7niDKYiZXxOAejq3KmBuBxvZyOqgL5PtV4W6T8qLX4HGUUfrRo
XiQQIPXcYYrxfnUcHR3eulkqXhSsDw1wrABGiUlzcBSBjOaFm0s7z34qYEXyq58w
U3ct64CgxrNAAm5gam8qxcRqFnPi9zvrp7OEZ03rh5S1GdljFqcQoDpUKliFjnbf
c/Om4xuAGVVun3rhDTzv5lS6NaudI9AVOQiyubJpkAJj4XjhIlC5P+sKQnPjsC8a
N5XtXF8uw+uKTkEyPA+QlK97bky6eBPE5at4fb2pz0ku12DPPPVhGsQzI0K8CGaz
zK5RdzIMtwjqhBoMV0203ATuRi9/3DHpSsxGZvOtIrLCF/B9ckLNg7GU7s9h+Ukg
AVajEHPHPoenxzrBtQ5ZwUP3GOn2Uq+Cvkql3AxK3yraopBGh7hz1YYATgAk/je3
Q/4Yu4p8UCT9eIn6Ih46OvoSOQZntI/qL9710RTMpbXYJyxEKMOZoAiTt8Z6ADJW
UXDaZuI30474YM+mcv3lvpXq6fbn4Zn396jf+EJTGKgX6nZd+6Sf9ch1R49v0j0y
m7CkhI/1PrbupWkRDg4UXvH2sRaFXV744ELSdbLghoK6Q9odPNiTwTzRQBzjZ2oy
Rx0ythHslawTT072ZarjW81H3pc8i/yVcgVtfGUi8nAiIDjGfuppbvzwOEpeLV75
BN09G+kajlB7CfOpT+qr/ZztT0DyK94XdxbV0Jejn0evAUK/8IJudx8GmedHhFN6
VC9A8oqj7pfl88vlXQLYUGfJmObNGSaCiQ0lrqink5ZvjHZBoCe+kCEfY/mowaYY
3txw/uQaVo02kdvNsis1ETZ1axO4c4xRwX9Kh3pN1OVY25IPvQ/fyzZRi1HtgdrY
85rgp+O5bpZ3asWoEn5CmbsccNRkQ2ftyDCi2y0zPRHq9oHhLKqmOXc8jm0yGENj
ZNY8OQzmMtyX20flFHgE6Wpt+jRTPqI+63ykZ4wjHV0qpwC4kNRrvUm5rg1cOJog
JA8Nvoay/c4ycx8xyciK5igqo3t5Wkmcm7wKswhONcQrC6LB3hVM8cxumWjLEoGs
pf1E+2H4LZmKAnQQnLEXz2CzdGbQD72SIMtQCm4xyLq95rvASnoFWIOqE/Yu6UiB
SKgQ6XEGBGIJeQ5kfK43ydWyKQ1Unqy+scrdG1eW9If0YhnJlFZWBC4LCfjXC3WP
rSXUid+J4ZEzXjdNkM0KrsJwQl4kS6ZD4/HE+Az9QogmqnOkqZVbMnFMI0Jqj8jd
MoInpK8KKMqbh/+RYcMPpotIjjovPrmwPLLaYjvHOxVf+PG4bg3oPCiXidSrJxrL
VkFZWBJElS9Opw0LeE4FV3omdHalxzMzBGNIlu3b8MNmAdTPWWFrRQq4u7g4tzdB
TILDwxv/gApOb5mbeUFRZ0mFBJUu5SkJMuJhmjUnbKcs+nCTVqZpsXwGrc3x3YPw
a6X8lQ1UyPpzXRiS72QIk/qVmEYkNuBGOAM5PGvvf4Wj8lpPFNmIgkTv0BMIw8ev
XR/lzvQVHvgdyTPCDExcyJcN8qY4vka7DfJzbcBaVWaGWN8fGWyM2FA8HQpqsdRu
I8zE3Ug9rzXz0A/fLN2jfbXi5UgMeaDXeQQPBtqJDKAmv9U6NOKa6LT1YsGnzoC4
9n3/2AlMTbY9ebIVqmnyAxUH79HPG3sJ4y6spfiEctt+j+Xt2NeUJpA5eW6l/52z
+sVIOb7v8Dt5gyfTMunlOhizirQxMb6rHn1qQFnHBJtQhvsz4gHrbjMYkCKlmS18
`protect END_PROTECTED
