`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U6Rd7ubDdxIshkkQ0I43/zuMRDdUwknsyZYoqClErgGGsA6x/YBDdWwkiGaFclRz
oyhNqU9bUESlwZyKb5xut/k3R83XRYrYdeQbUuJgrL/kRnj5ErLt25hw5Eq/6pQy
uFLWOXawRopQ2bJK5FwFGEsNSciU5RtDJkbukO4ZFvphsNGX/Z9YXCaXELXHOG7g
R5St5F+ITIOnRxIK4WnD3uV60pKfPO0lXpzRCVxaLKKPBSLNBTPyghFNnQN3rTY2
lgOfz5PIdmqjW64lF3SVHML1w+DsiSCu2C+71ZUYsCB812cqxTvMnIUW8xkOkpss
ciJqLzDuGqQ9eHQMcAffHNVXu2KN4QGlC8K0gaQQXm3lnEB7JkGcpuTgnOushSH2
Hx9EYVmkVVYGzENhNpR+/O0S2eSXjNBXNVDlRQHkwlbqWqYtAqW/h53ulDw7XpHK
jm0zGR2MzmUqWbnB31Eb7AhNPot9k0bEeZYC61ccNz1h7rlegM+Xd9O10FA3fGnq
2VLLf5JHxkmsKb4mGI27bpalI5qF1LiUcmOxOsCd0q+cg4ZjVnYsKxF27daY9F4y
+aRDUd+FNiSU/Q9SqQ/8/3OqXmb7t0/cl092jJPgcC4WM0loBEDC5GRVnOjB7Ara
Dja6sjYw79ttKD59JClcBaLV00TL/Y4C95jaqBL182ETKcymLikN0Bssaj7iePGa
0xpT35g7nJ/OHRcafvee4KQg9k0f4o7OpnQWn20mkihv+7jB/8R7ExJ+eB+tf/vK
a2HWqTHYsVDFyzltZAHypTI8z5tyzFwhGdKL7iGui8vngZAfuT0EkcWoNeiRc5IB
uCzPHxlf872W7L41zxYTXFQrYO41mmJ3Jszx8i6OBJHfaoRBCGSIgzUbBexkeLNW
Pq0yAYY9VvwokMAfnZ1I9b2nmsbZQrWz2b8aHh/29x7u9rF69217V6dpvqAVL0cc
GZQWaJVtc3nEkirBl5djerxfVGQb1HntWHESYtmi7l+4CFPHmtES0EqNPE7qasL9
gPPN/XktmEHCA1sipcw/qiATGNB3pCLqPaGJa2f6GiPSOtNGVCj2PLcyyVywErBG
SlqVNiWzAdz2iIYCBbCev7OujEOayjlzneY5J/HNzT4YEmwPzJhaYym53V7hfSPb
3enzvU0SmCtOJJGm8IwArDmOw/BdxK9KoXCwG6HnlKcHD/iooLxLMrwB0QOeJzpy
I0sc4oKOo839gepBNQza1BsY5kbTFFxJUYoqyardUzoQQoOVClOd+2b4zAPOF+aZ
dNyzOmvu+Mw5hS3UPzZt9hOvFBGJg+rLskr1NhE0LUPp2pxO9XxjJkqh0iBIk9Pz
0+gzxPo/1dtBYhglPpO5jbojZEsmVkrayO4YbRFfv3nq2ZELVDlJ9ndfNgG7QxOI
rAk+mF4bsgT7fPmv29tEvduJypYmDwphQMZhIF/Z/XROBi7ey9c3zxoVPmpgeANT
G3+X0Lwx6IlFcipokpvFJ+XE5/QUlS761UT6x0imBg7lDcHRTFnBZnQOWl2F4nS6
cWSesSVutO4a//lhKbLcVCFP1L3Y9FQNdI7oyHzq6WOIZjeUBDWSlm3m5h9d+kPk
r5U3eM76gkfP1Jt5q2ZYTvAP0bgMBPeGce/Q5K2Sm8xtHD3yorl//SBJJlTIf74t
LIQ7kWvpqBPJMeW4XlqkuseEOWZf7cOKchNKziL4K4k=
`protect END_PROTECTED
