`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pq5cnAaEsIuRId+2Q8bfizTTmlJvB05XY4St0wTrSNArYs32NeJoGsgHi8XzF+j6
4lX6+w6jyRe6Hn9xsrN4A+0whDi3sM9BxOMVV610E1OCxoFdaeLKxpdDQ8Ud8yht
RqhH+ubHnR4qL2uq0qd7lVQO/bxsn667RtOhVETFPgWcprnlwvE5ahnxSHYWwsvN
eHqf/hEk1lochB54flWADnVTSpuN5dNczcbZjf0jpnfgnGyEKnKIyweoYozjDtWs
YYRrp07AZ8JKjASt33Wiplx8qn6aP5mvYByY8OWKwHXqWSOMiCC8QcSQcEtBD9C9
IijPChoAp7KPXzZGGVl/H2XK8rD4ycMoxKI3VMmcZ59gA1he/r7vRGpDZPtF0jev
/5/FK/QZ/+5unrhx32RR+YyFaGGmDvOronEAYH05d2zmGvTkFeRs7rVmpThRIM8J
pOctxOhnFuegiSul5gPGm+FO+v7YdTjWNpDMjv+32uRE8a/jDpfGqgOT607MKalg
6OE3W7+ZyLzh3PJAs0Hj263L8xWPQqXAXr0l6PrHsAaBSagMP3M6/6WFNzcKLUiD
+NjXmOZ5wVeADygneEuBZrrqRLdLZHD9w9qUWwu9Gk8TX1vXoavUDv292BTA+C0w
N3/doKElEg+Aik2x7c17updIgDRV/mXri8n7gI/I2BwL30iQDTPQJ+hd9SBSog3u
7INALZtQ/X7PoXz2N1kiE4NWU7+CyOUHHKPh04QmV+LoCYrd+0S3h0VvcW7bnMuC
DEDJ+i4m8O+aDNLK4Vsk+KEE2AS23/KudFyXL9e9zsVfZLxMyw4aStwWoSHHz7AC
hiI0euAQ2VTqVazfn6QL3DbYMHopx2GySI5qqff4Rh+JOPneOlwF0Cr+C1Nw7FrG
7e6R/wegpkzMHo6HSP+Fqa21OGPEegj1yu2eAKsycByG5oZNZeBTFdyWnMMrSdfO
4j1S2sHePiRaFzhS0YhAw5qUiLSdS28teunFolBzDc/lLoyPSC4oN+e3HlyvyO54
lKBFs8MHjterFMHJPyub+hBCJbHrNuGdVZPbBsAw95DalPsY5z2GYmkpZtS8up7k
9JDpVbLPBbUr1YcEQJdK0trn1Abtr8pMDmlRuWZ+eVJe8u3w1EiDgZek/OVEEqRN
HmLeaqOhgkP6SioIZR5b9f5HKEKbBjmyLqpnVdggIBelrKXoJQHDVo3WHCLg5vwa
KMDKjy+EruOShfb1XFsM1yfN2X0yW7Cx8R7ZCOE5W0PGoILdI2xpalapO6mRtNeG
XyOgcbQ+Wjxunnw39SIGmi4/zcnMyzzbAn//ro0tpqUz8D3HGjOzJFAcBqCq8bOX
mqRh2bGpLz08llGsydIn/lDgBm+MKyh9a3ISkAq9+2iZezD1aRQXPSJXm0PNRsMr
9/3nX90fCCottA8/Xj6COEzP1dqxOSMoJU6PR2esgp7PcrvmTG4LUdVMlOQd0QDb
xQuJcisikdnf1+HSc8ShI5y7Ur63xJ+tQimJHzGm55E=
`protect END_PROTECTED
