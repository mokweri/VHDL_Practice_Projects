`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OVk6oO5sq9WNPeKGYUexPvfgMBl+dS1MZQJme0/nBEBt8NxkNXxClyiOyP2ywf0v
6KSoWIESqq3wakRaU95tbVBBX45+O2LQ5Ul6TxEzdWDErkJAvHAIOOQEIErdp3jE
eAXvqNAmjJutPWGvmQM9EyYBBWAJf77d8EYF89Gt5bL5x4wBquavjEeD+8X1sOvd
nYAYiaIwyvrPVbyo33sGLBDQkYqnfx0Z/CoMJsQULIo2qSxBYxukYXikbw+C/7VC
qvCDWKheBeLewCrofQDZWMIIiEnnr8Ckr5/q5et1V7ZNdZSmzg4+FTT1crT0H6Zq
ts+WOwRC75PQ5jzvFM5WiuBu0cEKjMtWyJEnOzjvhWJ64nDy/8eiFyQ0ECN3SoDf
jbTVKvC7xCSeZAXfYs3hTjorreZywQyY3hMIeAoLLIl5zuHZY1uAvVm8MR06213A
N25I1gUJN+0dHDZWbZ+EYkyP8L0WO8KRB25BbhEbYUSHAL5ji3FJswv1OLp2EDms
gbTqxd387EFtatFlT1RTfAIgErUGHlGiwbh4N6DgWR6Sin7AqQ8OS6BdkyzmD5mT
yJbztW6fXO/NMJ4Jrmz7TkjmoAf5Ctav3zAAixnfgCzCZv25QmPq9sPPX3n1YVZ8
fjGOJtQPeVQkeJt7ZL7Gi2U+pOQndLst6/x6TiCShWZ+AKvFzg5wfKvfUefkSDrn
Ooiw6RGQ/ONvHZe+nOKUrOtjN/6ZAJLGAQPQNFJ3PFTkvHKhC8DQbhre3gZn15UZ
WxCx16xMoLujDpKjzd2CTBswur21W8WCmoXYMd9tuiCz90eLreP49xuXAa4OPMNg
AQBs0lx96QetFL/le5wlKwGiI07Rw3Y7b1VedIyT3kt271PaRMhZycjhuG2HMd9Q
lp72FPNZBccWo0whxZjkxP2jtsdOnhf2DrL/MY8hJvR74rJk1Hrf5EGC18/Egvp+
w/FHsC1zxUIAJuvlaeAltJwwfC9rcmIfIUaLvbw/q+sFHc5MKmhJwBTy2TBuiZlh
Wr4FRe7gV2s2TqY/FmvpTghDpY8ttioobn4scsjCqsZSGtMnaVUxINi6D7AgUdrO
/6rYNHfFYKt4Mf75SbDyR5Iir5wYA8RpJ1R1UK3CUBoWwRZ9bJUugF4AzYFiCZql
S/F6jNdoFcyXIaTEPDsRZeLsSFQWJ0Hu4KTkMFUxhMktl3KmGXiWpsdol2pEA6gk
C7zUZ0OyrSMyORu6AWl9k2Fhls8/4WyOstNKP9SFs6jI+pBntizbE34UcmnCb27i
J7EkmX3fvAphT8CEHyHIDmqklwFiTJ/BQ97xE6DCV1VU9ABO3RjSQ6LSXlbQQ6sq
Rz9kbX4+stNrt++LPj9SL87zFVpiOFbNVTZja2ndjLF6kH6Dn9g4t7EKjFIQViKI
6wNzcbQvkuOOvp5GijYGiVI3LxGK6xwljicJnfMGFwz/DwG7GRLJxqPAdjctWpiF
zuNqy1HJpN0TAGLNdP+gRV61skUspWGxxo9HVa8ybkY11VIXNQFaaPQ05rU67IUZ
wuWGS3d2VvUr7tE5FmcrLmCHD19QMpaaAW1xg5KtbGV8fx9ClLwMNY3vb5N3VM1h
Btrnd3WDI6Svu7VMwgr1yyBB+zMMTc/t6Ua4ON0IZYXlae+RO+pZASXGTPY6V0rQ
em26+fKnCLiC4vSVktlWDuN+LkIeLZ0pYZHLtKx0mYQDY846DI5v1iPl2EDRzzeW
HOB5Jqbb9LKIwcmnLgWQA8TI76hAG6SNHqWwgYkrTO+nC79/9BE8QXPBgiyJHEtl
0e17+TeQvqAGnBUHPOYx2nW4bFUlsb3C9Yrz2dO8jfl1KMY7S2hyYAd2SS6QIHML
vdW5COYYv/Gq2pQvWk/S5H5XjKnbgD/UD2NVqoH6CaZZeDuDzUWXUbIo2e/vInnh
QAQxTOSLjlScM5wzBDAzxomsoFkEHhGOn3+rKg4YmC+e0RP8/ELaLIx+kVpFy56U
tSCPjRWyo2N1TQoFHFCLbLD8diDJYQoLW94NsqzAqwFyYFuLQbPo8iQd4z/Tu+lY
h/KTmw/yI8msmXx9zYenfZdvVogTW+jlCRO7PvIhDQf9DPc6cHtWhEuostjTEhA2
aO3zpcV9jrTfiN9E13qZP3nhtMWkioFiUao7BSv4iDgv6pjlIXcLy5ZTjBF5Nejg
V84KiCzwmtxWXwKOfofOAkF2kJ9vOS6HVd8ocdz5l3MRq+gjBGTuehDBjB9iQKzQ
n8Yki3rf0KYte2lrAU8Qs6m5WNNRIk9WK3IgKnbY3cLloeYLa+4emNZPB75mlfk6
UIOJS7A6CQJm5gYyCN6vOecLIdhGdHTCyKq+C+9tP2PJW2715V1q5/YYjuNKhsSO
bfe1SwM0OVHn50M81UZkHWKCDqcS9GENpZ8kxt2wp3osbCcCb6DUc/1b0l6PgaAs
vum5mni42BlqBk0GkYKIaPlA0mGZ/Jxi2Vk326o3H7xnjIR5seI0HvLDu0Eb0mMn
BD1cuajO1yUqvZgN7hXHDzdE0ik0ELGloDQdmw97wNFLbHZzSmkl8irUnUu4PzdF
gW4CQvnxaioZx/+azqxskckjiagB0jutkKfKlPGUK53kKhGFBeON8MJ5Jb1V2Kkn
ojkleBMKJ5iKTyvNYKsZgOxwvLS7CjI9sdCpymAHv/ngnPnwFpaYgyyTA9vvDOW1
Zpim7kLUpJ9jK91gfna9RKXFNKDDe90vT2XlHfQ0MOCGWIvekZ87mZ99Y/J54SM1
pVTwyoKvfvAIwgdVus09I+AzxN3kM4hE4DTRR5Nzy/HQNZCeDqxxUStymw+UvWts
sluTM3eY4jWbpSvGZ2ebvcpEzfk5cagJPuhiivwbZX4lNyB+p1XseIzfEjpzUPPv
v8rLgv3VGHSq2c7TuPIFb7AEpCWTyWPq67sScjJjHvSfC+AK+y7tRnGYmMvXdQ2r
YRKbeLAkO2SPYcs7VAPCftfyi7Yud/l5XtboCWSDEtrwkdjnPJ8bQ+45yznrv5oO
21DU3gkzzveRrEzwyAKYq/l2ZBbRapvujKU7BnVYEEriCmeR6FY/5w0mibo/z6De
cZsP+fjOd0r88dwD+qTcfWqSysaK1RYlle89UrHwtM5UTwX7rPdO60asZpb0CIeL
mLz0Ac1KNyIpEPuEN8MsrLEeJQoIXUIa7Du1D5iZLTeYGCDdrxDXLFaO/3BK+uux
h7ia3gwXuVHaRdVu37dFsd/YeBdFBVsoVcH2moeo+o88YMMkhegzsElhpFpCGQmT
fefDXP9Wf+ujaPQCeWgVC3GWnaSQDu3Ky46xPcwqLTE7T4B78qAdhjuaaHtFrf5B
qrQD2pLrAWcSzXUn7ssgPEUgOPXnh3a5F1xmjhSjPKm15MhPQl6BwmE1PS/0k9Ra
GXxRPKLuBfWVScQomVYwhRbo/Yv+XWHQ4tp4BI/uoahx7AUZVBXzB3rbaFfgJbUk
Nui/1f1AEVujjSFI8LyOvSBrC/nuHD7XraewMU7+hN7TkbVIlKziO7+uCTXftCtY
mYYoB/cOt0zS9BgGOkAXdyO/3djUpBFEXPv7O5Rc6uRQAYn4lFVlQuQ+91VWDHxe
JkjslAG+s5ll6HL7iRb8SY8NIK5bdfmz1haeTRstUAvA6A36O7bK851Z1H3E0fj7
JdvKnJGPm/DttaSWDyk3BFJMZkkB7uXDqg7Sw01ayHxGH/t5MRNI4N9e5SkXAD6G
oMbbNC3iRN/UPQEJ4H8JkBv0pESeRUUmu36d0Em5ZpWPpStcrr9qQkn0HqjhbKbP
K1b1yenr4dN/mjalu6Uz6f3RUUK4ShLg/hCaVJb/Dm7zZlJlNLIHu7I78I2vujjv
qINXjiQ80OFCC/qGdLo8OKqLDtPuyxYr8dAL7lZ4/Jj2KNPoFqkKhRTDNwLt1W80
UN1mP84Byag5F3L40wKzq+W/Xmr5q+KHlHnqOShemOt4F6rr5yF3l1JA7BJrJv/F
zcoh4I/uTP1RCehF5ebJFX7Snt4Co0A5hgufTU7kGzY=
`protect END_PROTECTED
