`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxVA6zvmAUvw0d8LNfRa911/csG+coSc2HJ/8ucathAhaGkEfNVQIHhaYdhberB3
ZhbMGHyAZZQcNNjXeVOzmH3CIsFFIc4BH7Uhn430HPll/3VDMU20tZtFc8hitSnt
fnWoSJ1wKpsMLhSQ03iwrQ4qe+XNq/CRrSwZ4F3cIEL6O7NfBq/Hxnfw/HPsUXKj
SBvaVrDa6FgiLenRioYrwk8eWrIu286tJBDBmusob41rq32qsnL4dV/fZthJ133X
C7Q3t8kddyAcRd/602jspRVqqgKmHGW+HSAYcbZn+Gzp6wr1/9faZTcmzGwc5BHs
P1XvaiMxYLJj9Ez26D/9z+edg/qmnlX3WL3cxuPULMWSQsDtSL0yYNSZuqCeEy7b
zBN+0CIbeLZjtnCneXvZ0sjLOiT7p0VTNXrtaUkiezax8f2mPufF9VGA2GAWJ6XZ
WBhjP1APjiC1pPEvG9/bA+DLSQEq2DKJjg+EAykugIRyV0Ai8pex2xPUK5WGQC74
6D9vj/ma4FeWIkW/u5G9u37fu1wJIL8gEFjDdIueLHoAU+Ti5dGjakOhvWLmJoz7
nEuGlyS35PDqKVYL/Scuj5rhbi8YpCv1byJeUKyIQW/A1cIAnqPFJdjaQIrN53bj
+GGYvoJx+ENFrvvq5lTv/qSfMhRb0KSGg8cQWdlew06lAm0hfYwOQ8FrhnX79umO
dOA/1Ny2MygzwlKbsrPoNLoVUhT9YElD+oxG0XoO2grludfAtLkPaO7zl7m3wFnT
dTccAICX7oI/gZsxe7SUau8Mi7Xd8+3veUAl08h7x9FsNiDvBVrdA6Zs78UgiZg3
`protect END_PROTECTED
