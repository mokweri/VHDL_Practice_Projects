`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QoOyCiTGutdgZJny3xjECUy6rVpSQn3Tra4QsnvuTWwwa56eyQUy46IWWdi56XYj
wIKRujT3m1+4kXqhVCZqvDGMsdt8q2xW9rmxY3wP9+TpNwYJmuoXV2q1fEP3Kihc
pjMTjGIp8X22L3TCGoNYO3B7fclUM7N08KbqO1oixqmJDz0NmGMmLSiOuAsmti+Y
hafUtX+MawmzgDvuzzZzi6MHzkXMKmsyQUyS4Wg186yW/ZjwVzkkohLnqYIA9fJw
WXb1VqELOhGQKE2qXPnxgRMdp0ydDkJ+D82iOvQoQaLEWq2e1fsFSdaSwsdAGGYX
OAQ1xcSZEak2ImENjsJiEJETfCPmCewl+GiATRG1ECfvPCO2P7av9WBGoMDDUobT
d9cBcxxDHJT9SKjyaYJyXGw3sb3vYlkTuOOOKhfcAu5bWud8PsU7Yl9aaKnNjTh3
JSioHSAd38mjw69IfiLObmmhKuJEx2XFL8FF62uY7qa6GdoSRvF1seABpoliDJZU
ieHo78uThEkXO5qNguLhoAgi/YAmlHn/Qs62D0K0HHcEAKYMMPjdVhrdXaTFKpzi
Stul5wMWk6XTILtKhqDFU3Ztvpc2teyu0I8yN1OrrE+uHx4XKRIMElO6TeNE20kc
RP0wqSneM/naayfOMS0ozJhdH9eYon6s1odPoRZzXMYIkBNL3RMN+P9hmSXjdX6W
vn0k/mWSF+TKLs5VMn5YoWSLLeU4Cx4Dtgu02Y7Ci+PDWOVbH1NW4Y2bUbwd1E7x
aGNa5XNCfNZ+l0kLyrinoQN/tuTTmGpV9YuSVN499bd7fKQTxxSA+S6KXsRla3m5
P5p5crvC3a/erqfeynYbZ+Y8HJNDzwXDv2lPusT1pCdOeGf0P/MpC7+djR5qLavZ
6JJ1ZIDnBFXfU7G9iRR2hStcUhxiNNib9UPMXBHbq385pyZxAGBfW5pV94iWKxGR
z/FMnn23UOaqw0Ug37IQe7MrK6sEdModV5llvVR8ndIa8uvp8m10bqDrwurnDyrh
lcDbvBZWAXPU8F79LO+aLGr4PgybnT08CM69hVgTBbOXUh5Umvcmf0HlsYCETkFH
jh1JBZLIDOTOrQP58SmDHCRHSZzfbfNUjRniSLngQvjxoGYAkaPpa9gHhO1QYIxA
fLk3/22lhxo4f5dAcvi+FNl5Ts8TpE36kqpjP/Bh0+XzB+N1qqpa19OQo+AYAvGr
iYN35WQPTLbAPVmb1gtSmZypTtzwtJQZL4LHkYVHXD++CfMVXx6uRX5YNbKvgtB0
BUxR9oDsIS0J9jLk/M6E9B+hIDJMVIVEYhGyYlCPuiUlYgrHx7mYPYkClvpWnlF4
9eqzDgdmcNKhRjRMmF6WRZpi0BCJKeqLqQR6NivXq8qzwNTnjS+ncjLm7TrW0VS5
d5o3hFdndSWw9hbYES/FYFXDx21J8cRZy8L5zVn1KWBTZjoF9h83tS/duYL0XVPi
MsSDiKg8X7mhtStDHSZXWbnGKYvWyCYVgiTKXOcnuyOa8xIts9JLIJX9CBbJKhFz
qs4k7/Hwf6+4YmeKDAZrWL5VSws4tVUAAOep3Ps0Iqm+BHvwjX6Eu3R/qzW6TbV0
ig2Bz0AUO0CAAM6ugHOzjc74nU0kAYHKojmwAqEsvkk=
`protect END_PROTECTED
