`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MSw2ZjRh0s8ikiSFzIAIpmLFOT6wKeGhorn08/KojkdtNPD89FjiTGW4UlGmVPem
98gA7u2n9At0zyrl309iUQxK5XyMaX1WqccLPxpSGG3JYAd8j1NQEuWfLNL3W+Ku
Cxhss9GpBjE1QMKWO2DWFkAPWyaJfAl8+o8/kQNfJfeiyKFrNOQGKvj9xpKUmdAU
Rt+vPjEIBvPJR+X/F2qtg+40nvKRe6MEcLpHZIDc3OUm/kPxRYa5sQQhwl9ahHII
cP6yszACDzKI83qtN0iVZlJbK6tu3U/hgU6NmhZWG+4f4DAECk1UiBbAmiBWlVD0
D9FqwyzK29l9nEzwE7VEYoB/eJxiXgVnRbMN0OeNPWk/6XmXfASFPaBQ57ZDlbJB
KnY0UWtmiD3htVzu/+xJQ2ztQNXqpfyGL6miRy+hkqSX9NX9AOc7E7+AbT1F0HXl
2+Seo+D1QeXcHq9jRdoDZn/ZTcSrkeyuBrjXtZh+rVj7GGAJA+lyWBXnIbTC1uNL
Pap+/VGE2t1SmPheakI+SLisCkiXZQnZ8+tZ3fSKSK7u1EbEL2jUDCRwsKsaJ2ez
Jx14DcPPeDdtu0tpWCioCIn2J+DCIilVGmvzbPQVixrBD/i6I1Gjst85B0HEqVBH
AOQ76P+Grf3kXvReCq/QPzENBGjBo2uXgVeeldg+ndO9aoLLz6Z/UVPTWjLJcMxx
+ebgtu3Pu8KyXSTbWIyNKW3kLWqd0jab78EzMb12oh+JPtrfwtYLV9Dj21cUIQvA
9EjnAl9nY9JF0KXwyYmB9PShtPBDmSXiIplEB2QN2F9HHn2Us/Hq6TxPBKYcvLiU
iZuFZuo0PjZkKNt2xriQK57TPgXf5CVC2XVxxx8eBa9jQy79vj4O/O0GclfEhAmb
iCeVyVR6jPonDc3kzts3+A8vmSEaNazlF842or7ibOeBizAVlXIIv7XrCSdehRfK
sh+YU75jVKNepHftfT0t91m+by8jKg+LC7BJLu8DcFSvbniMdpXCV2DeqSUsmQi1
e7F7hUF0ZrPngb6Ji1WDUek+fAA64Jesat45AzsaoA2ebrPxfag2OUIUmCBDfhic
+Kc+tVD/JJYXw45qtHI5HQUkJBlWaeYiIrdhDhvPqx6xLgIPLxIkOOCZ2FLagc2r
YmG66sE3Ljzipm8848ZlU8gYjTUWZFWFzb8m2JpU9NbqDWfATzIlmeSokJLWxSlB
V/PKGGAyMvizq4u8QVbunXq9Z9ToNjqEUCU8kDapjM8te98LxfXlFVmqa7l2IuiY
oMKpraKwtrKHVIEU66inyqTSxyxWarYyRe9JGfCGp1ARtDsUkCVpL7QcIU1hWlOs
t+Chrmn65WL7XFGd/N0iwGlSuP0kiunqLA66XrEYdLVVTaqj2eTBqH5/A9qQ2h2M
U8lqiabKX/X3hY/a//8wFoSZpWs1gL/GSf6s2k7D3aggbyiF+dULX9kkf7ZZWScv
0+q7U8DCec+2DzJpW4JFlO07KowpJBs3TJG/AJvswlwPZ52zhp4yd/0FNBRRdpIJ
zFPbO8RC2+HG9a/vpD39lvrnKqA8G3u/Fg5RmCyuYTiQQjwRsHW+Y23AoM5GkVjZ
Yb0puQ4K9wdAvcrxWGUhiv91hSinwyF0N1JkH7IaeJl8GR2sC0dHGr61GndRmsSr
U1ZvaQItCGBRtX1qPR83CDH6HS6Emp5j8CpltCHgbOJ/fSenFa8snHGp+/wN/1t/
NdbU3MhNV34KLM+7sP/Xg6fcc+hhhkwA+DMldusxuY/ie58ZISR77e7H/3bqjT7e
eDFC9h4YpyWpqeY9DrczSb68glzPJKPxStsQEteL829iZZGHH3ZOuCjBttroCt/t
o67QgbjjDL13yfeFKp1TemdSyQYFs02/ADh3IaGZkF0WAJ4U0Fi69CztJNMXCQTt
Bys/5TROIRWXeNK7peyizIRzeU9vGtcTWAHIy0DBA4xWY+vuYRf+ZTHsZYqUnbb8
xTqezl/OWXqsSRZHkJjnPkdxu3uyrIf3+e/BLQW8gO5L7/yzqZrZNy11BNxhWno8
X4HyWWwZ7TKHlRdJsk6CaKEIMGxrq51xJ3VWCiNgQfwxTwwRnd/soAM41GqXXXnO
bCU/eoxddOzuV6SR9ibhJ+xY/jcJL4HiDPreuepOM8i++XOYmIYpMIFvMDejurNw
5Wsvo3SuOY8BKjfsiZvBiCuDEo6BHTmFpUrsDqJMVdwkzMsH23mJIgDRZV39X9zb
cnpqOUYfvrpqpMt22lp68eWvR6TrTKOj0QmFDc1h0c2zzmK3jU11E9xCv132V/iW
zIfOWaIpHTkD/shuNxrryQ8GT1su5T/R+MskZODpX2AnEjMeee164liNlG8RxqPN
yKljnYbQVx+5Iu5rZQ3FB+sGHEfmoQd1Q+CEkwVQiWbAhWndVL6lu+ZCK+vTtuKe
vGopru/S3QdCcK4ZfCPoT7jmzbknkXVTFvbcSJX7nCqpsE0UsYVXUqNCrxZBHVso
Bb6UuPAcQBeoSTEbCtJnefGdlS+FSrSi/N2MND5Ik31S2+ieY01cgbNY3j4OJPW/
yeYUjl6cCmnWSVT0WTEAt3ZyakaUJ0dtMcw40gQVYYqHDXsSYgSdJwpobgJB6DC3
EWCmSO/i/9CcotIRzSHm6do6v3Pw3ESmet4VQTptO7bueBG0MyD8bTW/54s0cbGU
XqvDP2PX1nRpP6QbjuX/+BgYl49NQ31AYevRB/o8JtuY0c+GVj7PcLUS/xpC0OQx
8hWIPP/fWuJfTGzI/KHoBqNWvzDFrrYnSRxFgQup+hrHX3eitV4eCR+5NnrifYFL
pMb1IMg68x6wmzHghZIkyd3LvTmy6+0FmcESZeZ2WpcxfTf32ZPeO6V7QskJybkP
1mXEzWzufY86cnLfTezuyRMJTZWPmZC/ZOhaA1KOyBymRkg5Dn+rlWNJf8NaEAaT
MYLaaL1QYHMM7g/WnmU4RaOINbt8oYpdRbQQ4LZLJhkcEhR5wbqbjCP98WT7emYo
qSUNa0uDRwaVY5edHIEDxrCqGPTp3hhzXiaa354fCYRLQr5dGcuIMKIpD2EH7FBJ
ZalRRy/7hft4RsSwJn+xK7iCrW/H302MxsLPIfpNmsT4YeHJmcZEGq1qsrMUhrBK
C4DxnXav9pnpoRcIg5FybiUhSFMkaIR72wY0VBgJmo5KnK+viJ5nzH+kcVJbpzzQ
OgQ8q9CW7IbnjD3FuaEFhqE47RnYA+8qToGblzb3qukt4BB79IPGKmKzX7TSHans
zHr+QiDFWTgVZXPjHd6OJWYWAZd46wYwQAKb6tBsYvbnYA8Gl2lWjS3309pnmkVX
7VLFi4ba4RR4cq3HK9whv+a+/LfaOW8Jgy02YpgYqfmGOqEIDkCMJ54XAL/CNbtY
xPU6ks200UKT3FbkROJG7s4mkgrUcMKsXqbI/fO+iYq5sRd9DRtoFEWnOZTT7kba
Rl144BujNRVGkBng6RJdsSzNMOhqAC+CQBl1PjNuHofYzp8jLJJpz2i0f1RMxdk7
P2jzjEdlzOd9Afxu4jDwLyTiqgHdS1pSfiI93U9cD7E8LJrUGF3Ugi3f1ZO+qJqE
CnVM3KMwZxaeTIopBVpOF2e3mZvNv1TZl65AU1GF5QyjirwULLX4CS80tIzTSIlM
xNVvgVmp3AnLCP4Sl8dsuG+3RKktINy+fFfP1qpL/bqntrKX3je8mOpnhZMX1UjJ
ilsWHn/5NINxrWnQGN54YirZSAyL2OeEhak+CswLCgjBIqeDLpCTL4C43BzG28gB
E5wBRu2i1v2GdKYFjsoIYTm9523aE3fh6QkD+ri02tEyXZJ8HxgmpWkSPjq1r45j
Yv0SgGPRalMFEHUejCxljHoVtUC8DklRX7NEV7EhV6VaKcAurbDBaTU6N8J33AQq
xPv50ohg2UYPWhp2MvgYVEF/0isWAHeUNeIl/LvS8G6z09c6uEvUGblRvyQs0sv1
XZDwTXmJs6UGl/zGTe1wwSCKXylZsqG7u+s7yNU6BKZjOhQ6tLKmuLTHbC/jfsch
sP/pSm6fhMkfykxgXyMRUgsDv3VowUwNGDD5fNQN6wtAGJChrVla8YVGtK5xPYrH
gVef6bLafxFW5KIlHkSu+2PKr/fg0UYjV3FnEMvZ3Jikqbz1ophFTSA28beNPoJ7
gOki6xIbHrIXGY0nBhPknLKeuDPmtEPQS4LdMdHPSmsGRhLUlyYy7+Qy2ronLNVy
mDT+fLtpYTr6adwjgdvlO92MvLzzrD/6FHd8mnk193DQSOzBvjeHgQKBQSt0Q7JD
cHy8ppo6QkDSpUjgLbKyUyvLOcTXVTi1yHqETSfRvOY3HjCDnLhqIm5UUUbVNgYj
Kt0lL/Dcu4SE+rkJTFtAI4a8AGH4bMvvBeRUhtPHHp12K9g1HVS10WrwkLWoH8wp
6Iclwy/G4k5vwY5YPb/S9Vojqle76d+S3E1PxA5DW5AJ2cZo/D58rTBDStGOPxHT
jrIGKgkzzRKGg8EhBSLiY5ToFTFmefgHTyA3asDCTiLMO/B++j68PRlxEu9TSEjj
ZQoy0jZPEsaa/6GwytsojJ7dYmkOAISZdsKyzcU1J3e4ZEFWO06B7wDt3h00J5Pf
g1krUaZ7ZsfWAFzeO4ES7UZj5stC8w8NP7B7SeUhcZJ+JRwXkYdvqNhPrI53eG/b
6JQc9zUQ421rxY28hfCkuIPhMN+zzAAgLYIVhFO41RtF1X53lc1BJXqBeZW3acYQ
OAWuHqdtktOXWJIUQNXT06bFlXRE6UnCSkma1ZzQcY3/nkvQD1TAt9NWdDKpQyf2
+7z+1mBPWOJHVl6mnqh8LwBd7hAr1IK0NTztBUSdkzeEv8oKVsYlp22Gm1TxMVzl
3l5hS7nXBfc5tMTM8BZV0l2bbQFvN+4vfW+w2ul2JpMPaAkMDxO6Y8BuvFylWLFg
6m42/PdQngDcNOoTKpnsn6cXAdR8J6zkMGqRl89h/uatHsX74SNHjdP8mGTI9XyZ
SCbCGQEiPv7Q9IG0IB4tL9ADLJfVSG/G5mwBniLW2UEkU5HSaApVA4g2vHBOFr3z
+QoVhRuIJjuf6dEdfm1akgbZ2vH7fuZyGh29j2fHrjZ6CH2qLEUr0yEs9A0emuy8
ICbnSIlkSjc4724/dVCMlG8nTQUZykG8XEpiJVV4DGtC/XPvL78mXzbqekBQSG+y
oX+BDrQu8cTOchXbPg4xC0Nf/IkuMeYtQYgc19HdCEjMYIcY3kBvf8F6w8JJ//0Z
hMDlljZni9cTLXlsEQlc1K1vkIqgePfkbwdps88BljCixx8OQkcdwRIj6NkSzIaC
VV6nvVKYewRWkHqw6wpzGyeELeDKTIv4784PYLdsoJxDZwLKcAPWO0m6BH+ZMDu+
DPFoNCYCk1AL+OpvBPV6+c/nND7y12emYnhG6zYQK/Go7KnwPFXfaKqO6F/MpAnj
MS3uvVMr7Sr+lUkkRD6gCW4q9Pppy9IvXFcUc6itc/WSkwLnIHghy9cmE2f05pp5
uahW6T+j8tMFFHLTENav58g6CIOmyCptiB2vgtLqzACSa7T4bgUn3YH4b+MtILyO
OHwyosCkVWwqDbBQKztAuraHAmdk+KKq11Cos13IR2ejfpy0b7sXeBX2detEWKzO
K5kHrefVBvtR3HOMcXbGM3S9mfja4rk777alWIuFUticxWFcW3smyPxvWLJqnL6Z
qFGCRM/ayCURXyrlapVuqj/Y3aoi0qXmAmQMlhVX+3XapW1Gc6sKgZjjGfbUXk0b
jncIgjPv4Bj7nPs0BBI5mNLONTZhS612ppscIbEnO9ZkicsD5JSufgFlrORg5nSz
6aX2QhVMm9zKXSMl6gow7jImNop78cHLKFczjtmKKfpS1Mr7D9ItuiMexSMxcI5a
8MrDtu6NBMwPUJpN2Vx/8VPz9deg52eUUFfqMOErObQfMW4QTu+Fd0AXNzVy4WDr
MwLdzvWgsYHW76NyBasAgSpFQiHeklFRiQ0wRi1SYNU0WSAK2OWTcQZYeHaZPoLW
CDBKnNw7VDcoV5V7Y28NTKZHTrzcO4IZf9bRGE1ZAKaqCwocfmRr2qrZyqZXC2aV
fAMjyj6m3oWpl9giTavqolzqS6/pHHgk4J2wWlc5k3Est/pRNMz4LG3v1Hop6kUf
LBN4ouo4a33XwbGwCm+wVzrRpY1uvZrYpzNMWssVzPE7V7HiRkS8cV1fmDEIhhq2
zOKTB03NCTTze01lKw05pPpN6TrHPvnqo3Xm35t1NJNgvrdzXKaGGtgLBaRemuDM
+50YPnUXEvqV46ka4ga/LQ3dEt/DBc4ES8RD9I/eA4zBypdVkb3H+7NwbF3qUFp9
9XP8/OfY2xWxTznGwDdtbzJO9+M35OMe4F1WeGF7gzmGP6HnH/ssllGMsL2rzLLQ
bDdgo47chsodeS7nh/yGm2EDerc78g/5UVqjbHBSj7kwGAZ0zDeKjmFjB8u7D0QL
TxPOSsGRrqlAw7FNGicGEMeSjMn/ZMlkAKKA1gIb9CMD0p/Jdnla3Y7Xob/vPHli
cvhteDjGAjln7G77JM8d9P6gQ869B/+xBvXJ1N9BY8o+1E1jNhflhdQLu50BBL3U
y5+PJytjuZihwIcyvV15UgbwMtBmGTA7h2FZTd860flQsW6VtqzuiDJcedyPc+Mp
Nd5EaDycVNqXAy5/1yiAPGjg5+sk9eETWruk7JJSE3XIua3ihp2GIAXFgXstDRaF
LHu49XLlbvKfmbOhfvB2TNigDAFaWaAzx8iCce9VJRLOVLAwZoBSSyKEBAZNoQSk
xFQW+h72hQ94+t2kJeey8C9WmdSZ1mbS70hDu8Hl6W5pNekP9wM4DR3720y4V5ti
pt1baqvKYheHwpI4Y+zIPyguGfpPDLaYocCJt6AUjIcCnD4Th+sXII5x0fqThWxN
xRX8FlhmZeAEyc/OukYL0VEvEB6qSP8VPtNfHmrm3LYWfpCwxZxmrKg4W5dA7w7Q
lPWnRmQPQBvDQ0gZ13Or4G1yiqm3YgRW+6HOvDvbVvFhMs0139hUN3HVGdSJx5Uz
fueQfId5zFkmT+c/5TvNNN7SQxVujwMn/BZxBrE0XKfn3RL7tqlPxUqrfbYVwkA3
+SQNagu3uMWp56yjewTy+CTNgn2qUS2El7NyAsoqhKNpL+v0ahRHDkYl2hFZlQS7
3xXVU5D5RD/KQaHHT5/aXUMP2+evGkqAA4jNcDdf3sfcBTYgCDLmNpY1AiPyAlQf
X57+nq/sm8HT4a24su6rVc9Xn3z56XwvgnXTgB8BsKcvuLaFByNxIVOrhLgqI3n1
ISUDoMlBubXzAuZjvb0xV3zmC+nFxeyiePA9hNSNywNSbxGvyfDEWpV0yydQolSV
WvSwhbmMTw/GHl7tPIKUNmy3KI9zcBoKZ6ds+VuoE8ruWWpBJzuef4svKBbJiE2m
nEOqThYcwe1UlKLKMXa7AsSv9uRSr06P0RUrFze0b4WAmR7L9bjt83sz2wD78tk7
yhD2DFc2mei96WBfa8IUnfeO3XzcrEE0S3A/ktAOnIEUkrywhJbdSK71wSW4h9zU
eEH59SMyiLn9jlEHh2d9to2OQWN4Yvw/+Aq8298LSYbdadAqMYa0gu3V+DBt2hzG
Hycqsx+5E8stpWDWtrkNYrZDm2kl8cca6kBrvURwehProYVjG9EZVNifr8/qmP75
YgornIRaMa/jk0yUPmzzuXKwcQmDNAVD3MSHLuy230XRUaUfqNp/EdDjJfE4wrkh
PM8ICVJRvHpzA3XfsfC1dmsP8y34cQSXLYkAEAKwKfeej+iTeHVbdi/gOCGTcyZ1
vI6URml24VXxxV6MWcgPtXgO6RAWuyvwvgKxmVi214GWQ5S6rHcki47fDtFwuknp
5HdBU9qePxBpKnKZa6uxVbDCTjvhDSwQOV+t1DdZrSO9oxuW760tby9b26OGlXJN
xNfB7+WbLTaRbQO6/xx7XbdX/VGykaEE087tXwyjZRnjQIIuwAs4BbA+Uc6gSJmg
le7Zth6cMi1p0t9CZxzf48J9soGZ4VBX6NGhKRuvy/qm9sNve+YHOMvCrSTeTf5j
Ccw5Dw6HISJOiYtXMLnWvIv4TR7RXUHbJHbEoM5qMq9V62e4nPE7g2LBiAhBdtsA
4cDArX35rrt6rx+If4tLakrmLoiVt9A8s8yzU6w4aCvctbpZb5ETsDBMCty8bx8C
2VmVogAGnX9OEK+ne9Q9O4V8xM+j8jZ5S3yiq7F7AsRTMHnQ5Jw3VXsmLQL/L4gf
FNl5pGL96nVqgpVfe5AmUE+nR2YCt3Ta+dWHm1S/JSJwAZHXwjboOWYt/Q8uy0qL
Rq6Qv0N9kDciOmvRCGshYEGMdnFI2tPhMyKWWDsTg6Slwo0iio28hgl0Wc3pJlp+
+pR61sPx/DsWqH/X7RohNP4JJHKQItYO36Au5l2FmuUqvWswxKBT51vFh+j0bKJf
eWFnzfr22IZ5Q0kzrRERatatdmsBvBer/zRpTYz2u6WXjLZaJ7U2AOx114MGtJZO
dA3Icr9y8SZfIGmvZAKn6hUmlJNNkIhY4XfDFH104F3I6paMNNZyAitzAmQdQsjQ
G92eirvbdD9hoHhSmX808viRmNc99h9nVzE85l/di9amxZaTRMtW0NHtn78ssgvF
zoWxGYfq0mYQrsDIcwXQ7WlK8NzBU5vAgXi0Q0FLUJl1Lt7rrH+tglnORtWGWfnP
cwWgcG/xeFdMyzbkVolKTuRuhxbQNfTn7DOPLXpAOYNLJn25PZc/0T/1tN+pSa7P
G1tb319wdZR+rG2NPQ2tv0Pqbv166E0Ee/U09tOe0EIuI5G3lMrT7eW3wHfedWVc
50rI+nIRTEN0TPYPDoi6WJ4rrNaYF59JerWwNGKSAoOwtqhtXTnhzzFaAnCt5LyA
yYA8Eia0HHsPTnvFp9V+Ig/kB/VvBKXFvc1AmHibBaWxOIw5iupPJP7sglFTLkWk
zfRdnfSaAEOBydb2xmUHTvguq31JvqLJ6j14aEjjnrNMKgqC9PG+viQ612MHBbOn
EEM3wV4nytdrCgzJsWm2Re6gfKyyIKyjYOtdl4sXcs8w6ND0yDKpCAVxE1enHNzq
65W9IzKEPlGZ2M0O9F1+BVzzkxSux0UICT3oEPujWrILo3W4XALihXS0fnX+UY8O
NPYDDTCSdv8dOn0spc2q1rphHmd39NwSwchrzXYRQbynijIpgIbncNGMcemr68N/
P+2/xrdXYasfIXJg5q64WqjOISHPUFT58jFVZeV7MyDYs9fcCUaZczb+xwS5mVIG
pN+yvvtm2jPawxCWw+BOc2UOn0LrouwtyvdsaoLoPt3D4Ap0rfMlk+y2MLaA9snP
v2Pdb8+q29TKIi9mNVe4fNIGIcT4f01/FRHsaY8hC7izU3uU8Px1lhYXSUCCf/jW
pZWixXcezUwzL4GHKHlan53jSswAzNZjrlsBwQbORmDgjbcesnnPDMOi47l031W+
af31xrxiH+2X35+VBuLudrmiw82ul5XkC2BlOtXiljcTA4/iwn0q2bb1oYGBxVES
CN5h7HpGAbXOa1fmrc08u32SSlwDTTrWcVpcvSXOzO+UOwWQ+t+Qz2RLb8lOthPo
Hqm+yW6COSfma9G8QnXU4VViP9fURUyVltRZWDrMFeaPgLTImbHUyj1tNdoxi+kX
U9RYmuSFxMmGmIxZPTnLWTg0mwIwXQ5a7haVuGkK2wGm/hfvF+SQKQcbY2AOrNm8
XwvGy4ga0CCHATAliO5GfAkeQ2QRGY5lLSq8pWX8aeZG2kkv27xrkz06VhnOOh66
HrXwzD/9Vrvzs8UehR52bu3KNtj/YDaitCu8oQEcKvUfHXhfsQHLB+IItE8ij0e7
cZPGnJgeDM9AbFBHLesWe1Yt3by+M2XedarZdTbxM7mSlPrxsDvfY+O6jtkOrLpt
dt243s01x0z7epV9uh87hX9prmjRZgAdjcJDamWk+XLlaUacoROLMDXJ6KPAHkQj
7Sq57HJRc8WwQXB2UwDhLgrgcZKMLc5Uj3seP5x3E8+DT2Cm0Y+gga9PfTN/e9mK
ii+T21zj4LFQhHdQG/zFVAkTQg4A9i0jm7em6w7RFsVDb6P5V8PuZfi2vIIphhbx
IYAb5TCyx4qUEOXpbRUQXPQ2bJN9ImombIqq3FE1KIAEZsRE7ndIzo33j1ws/BoH
/Zf6A7sJpr2vpuazqpZ5Z7IOHRS6KeYZURR94vSuvPGBwzINeQm2kj+ijUUTD/bm
kMj3xq1DmGC0XBeA3r8YPLBNoyAUQlDKs9WWb13H3cRrklbaCbh3J7UlO8yKxBL5
2hIwY1JTLpHRpaaQHX2acF3NLB/2b/dGHypcqo1Fz3WSetBDCRzl77zOvYf98dix
FWarK5mz5UPfjbha31quELGLiy9NwAwAa6mCM+0h8Ey8cuM1LWELmkpdyXD6PaQM
15vtYGggOr5w4Uis5KU8Ah/CyylXvD9arHAwguz3u1leBIhnuUEapGTsED1upCPg
h0ruND2dX6uECy42EUQGWrbf//gchG8PEFSmFLgR7+xKVQ6auXeTbiT1vbyNgn+D
fUhPzQyUlE0hAGjmg9cvaJsXNq1EFTMZZrn0352+cJP6Zg6CwFP7GHuX1MBa6xh3
VLgO0tu3e4TA6GGzAGnsbl7HTIK1Gxc2LWqi6IJNJ8ZJyl3EOInPwWf0H9RGHBEF
8m26bjbABJ3VcKPSq50sqMbaD1G+LrhCwGVzsvNiHYd3B5OYwb9ySPsPUYbYuvZb
RSsifBThXY2C1NPG63Y+wkCXgYB2qI/fROYdQ3OShocIgetDewEBsnn88+MIFHXm
kbcD9MrARQHFE6UU/fnn2vBzgFlQnZ/eM5NWCkuBYU9njCpnw0gd0ycK0RuGif8M
+njKFZ4ubGfN3wbxTQ62zzlr4SO91Di2Iz2BsBMQy0AUq/hkypBwvu4cUiAj1K8k
Ze6aLUFm/f1zQecOiHL4hJ6h8EJIE47e/mFdLt+1bkmHbBwrIwyfCDGmTKmixsat
D7w936ZiWDYp4H52wR/bHkROyY0nan6dfemZhwRiuVkSpXAPy92quDYZjpA9fyv0
tdKoGJeUrSDem1sig8nQ/nGuJi1lsYEbvofu3KdqwPuWlDbvQAKLYqkpz4BFrnpa
v9Swd1qeh9264kdWMaz9irYl0MIY6fbwUs0piSP/sNJ+ngbUhErO5+c5plWZ3zmr
lFTx/ZVnN3ltZ8OGfJe7t3R56PoEcLVJ7MuxjLcb1sYWp95bD7LmjNnMMtUFkcPl
xNfY4mtZ+8LwRKWzRwzdy9/W3O/msUcKsaipwDVfVmIJw+D950EVcxnvLWmRpKc2
Z62joMF4O/dxixLWGoV5cWGcJ3Qy8ztRMHn42fui6zsP0Gvs9fccrJLqYY+FmP0J
l2yuR3YibTTtXI0AvVaK0DIMdEP2NDPi8iI6L3uM7ASnUxRcgbrF4eessANQHMGC
zU3lfyvnC3RPrP4mVBItLTT+DPqR/CpEOS2R7I6oE6W/HcGBD5En8pwFSRpXOzXe
3VL/QDXrKNhMATKkmdpLmsfIj1MiGJXql5A7WvD9P9nYpq8DFhQjPHoO76ZBFEaj
+ZY8pXWCq+0O9hHP5aZPMB9Rmr71X+qsFKhkdkRv27jfTShwNzBBmEVu+nG1CfSg
jaOhqCM6PbkMKlNdg3a/KyKEXxQVd+rvdNIL2t1DKtSp+3a/YSTqQL4TErw+VoFz
wcUKy79L+1pHjBE3oAuja83XBB0VKFUWNXwyPrD+DytdSXcV5BMWUAUF+mMBAQf1
XOqh/BMmWmOhS91oz9csmZPGvuH1o5hssdmnXeyyqAPetUJKVqqlmmK9qlfPxRO1
LYBcQ/4Ei+a7MhaLnhIKiJAFzfHt1hJLrzZn9IB9AUYAI38kTF1IluD33yj7Yg6Z
qe/uLvI7wJTTKAYqavbwl3mWWMyL3ycJQHfjllfOXVTJ5L8KA9zOKf34wn3dBoX8
9Vv8AKLKQlofIm/YoBolXz3KNwPnfmR6rREPz2uH4o2JZbmdficnHhECEvsOoUYG
IstkfLsCN7rKzVzQDAM3Zkp9dmWUXrp4OaPzAMb6lvhrpWPR6gHUr6NDuD6xzsV3
t8I9a7tXdPkX32V6b01gOGyeBpTbcWl0mWH0TXo8OwXf1eXsfNzC/0iwK1ovJ8rO
rlNvkyCveOmRvimE3fYuWs5almCHgl6M2KrMiEjVCNaYFn5STGaGVtFa2m7RZbWd
Mp+Q3diK0MK4r3qtslljwTy6DOn2VqpOy7oP7xA1wSjtzo6VwrBw1lmQUjffTLpp
z74bdFYvMrj34knQlHwRiTBk5bHLiCiuuIvOGZsM2UQXhJhquvvzHaMQDoqBUXGf
vLou2wjAWGJjpCRjwNxYd3QjHt+QPEaWn7o9NvncEycgnyQvOZpwStU6dDGC6eVZ
q9D+VrpeZnXOdeUL6dKpnlvG779Wy4pgIFdv2eU+hPU7VKPZdClzggQuzaTzotPJ
sc32gSUeqdnYcDVedfuSWmhMfS7BlOR6nv10+EY0iyqNEzRf2zsnYSIziDWIhTeC
gcxjn9a94jIAYPB+fxNSaRXg4UmH39OkZ5qpcGvtI9wB1x/ROdreKaT0azUXH0AH
7sWcZiK/ll2A83N/j9NGbn1lQwTef7uW0tVGXUoNlaDnvKfxR3hwQNuFXyCm/cbm
AX8y9wyGqtd7eEWyFkuFYdznwYsTilDMb8Go+5od5yo4joq+O9MXNd1Jp/0YjbK5
QJ099fWCrz/LMsQ2y4JDnYCac2TA5mnB9AFBPEdmUFkVL7tXHrFsJa90ksq10+8t
N+EnJ2fsRHV8ST+/7AfsP0y+nA0h2CIwuIcVSpGv+0lltSAvA4zuFAqRZ0eKSZFC
r81z4lFEKqmfhTwS9Kx/odZz5okmeEeousmp32rtX/0dPsPIPRX3+KIKicWXAgGA
VgyiT8E7JQZTTiYtmpHWyAiSLm/a0hw30LTfaZ2YnV1N2ZoC3xegnZH2wFGQlIn+
2KOrVh0NfaDJHxwHL4pi4nQrF9lpRUrJN8o/+edtG+3gu6Vj/PKUopEisjJeRFdB
6yi34EfDdhcL5ZcpDzwHDjUHC59GspQs3Fm4fES3FVTxl69LPES8cCMA7tWgaYT6
ZlkCXNGekggV5N+BenPJnYPt4bvy+izQnjbKW/tuDRfj216cwW8/sJH3P5SFyudm
bfb7gh1gGZQgsdX+jnEdPRZ7pVOXx1n2qjzJ+NVzNtGFav8+t9SS1O9Ih6Q6LKqU
LrQFycFVKizv+Qxcz4lXfmNx0Muj81hg7ZYdfyGJWC8wBfkylJ6q4Ny7S2oKn4hU
`protect END_PROTECTED
