`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qbSZGynJNCxXeuPg04MI3v4LvmbE5bYF4mDttIuf85xcEVWsnhJyfzoadJdehmcx
I0TjsSvG+ap/YMR1ykU4LXvzeKjDoFlrOkCspqHkN2Nn7p9XGDtC+j6GgftIb+6P
XUL4wi8m4a3nBGcycWwxcVNSySmIhjda+pCA5GY6naPbwjNu/8FvDDUcIn/Ib+qR
1eVulpkuM3N7YJQGwskNAz1D1+JQeSOvdfkKfGDFyVs5QnzePkUAMSSP5s90fMe1
k77dXtgT5/QpTMtlTbigIn0JDXjtuQNV6a4in8tiJ6thBaarWitNTlU2Bvd0Wiap
IPwe+tkzycyrv5/2hdV707uCzjx/VOQbGAWyFscYUuvyB0wpE7Gc5x9b4/luKhEd
S/z5emgylSRFxpwGkSAX8DFK+1Jx6tm/fo2NxZ6QIZg70mJtaccaep3IAf9utoar
oHznTKmRb0ZkIcSxaAYcIEDM5QIgIPQiG+XHC+4EFbMCH09n0LkxlCoNerG2rXjw
CJHuv3MoYDexVJFXAzirRf/+XSsGxMFekPWhz+5ORnwqdsRcTw5a3HOWFPF1/67W
3y2V6cwmcidFof0JKnGUvXjv7q+51b/CIeCTpVf70H7hb+Zpxd8xkKRDKCj7PCiV
PKqqT5kBEIWZFY2kAwu3zaq1+6DfZSnAqpEWHxDJZN/jZP9xZgHjQ22GqQAPMzG8
4AwjIcrQ43+S/G83JPp1voGSw+Oq4oDsQ1SyxWZpDFzmPVLWP/Rj4TjWHwBi7JK6
p/sZGu3Qk6qIQtCnaUv7mk/6wys86eUtF3Vf3dTvydnzchOai2/DRXArxox9tH6j
vtdryn6BHKITY6SZzWSXX7LnK0FO/JyoRlWckdypMt/ePZIeqrYieShYezAk/0f2
6eslCAUmDBGHCzrMxnhzm+LUHZiM0mbhZvJ/XWZCoBsukxS5D+R8tpl/gn+Nrkk6
0JigqAJysLT6mRYW9aY+8a8TrnZWTmGwxyW0DzImx8ewE6XBWCvTyw/DOXwC34OD
e1uZh3AODr0GLMPWsgo2NRuRHAhCxTVvgnkFofTWiOuIqOH+bCn+jS0fcdVmvkBa
sREFdB0mmTDD9mgWxkgvakmEl8E9iTl/iVJDPiXFPb2EtvhcqYCvcMBLQyO5Xh3c
BxKegwxvAcIe9yQBqomCgE5SSZjAoEn9NIcfKvTTAors+Mgg8tB8QfbGA1Fg/UNN
AROu/vxqG13FofPD00FL355aAVhkELh+nRqIEZozEFD+G3RAhdhk1HFBAWLBJSW2
FY7tZ+mQmKobxB25xdgHkx9aeWZ1uZnRwW9QIowPe5lXUH8fyITa0cxejd260BcX
e95aeX0bD1eMu2+gCLqBS7rx9qCDAbubNGJISh3T/kMVEik4VblE9fWi90IS6Jt1
m+QUkm2NTJTXVwnX39/5RXEY6I+98h7XVUjN8p2Zp4fQqHjNi37+G0p4sqPyQlYX
vwtH/DL2IURZrkZrc2Ldv14kP7C2uEK33LRd62JD0Kl1dGlROweOuwd5c0cEQ52y
JUzzdvzBMrBRx33BwNaniLa7TwRzMlSYwzdiRa3dkMMtSBXpSMefwdMh/pGgYTAy
pJkNtc/j02f2xckw3fnV+TqOVUQ5Xrd9outev65KQTVskKGjx//NeAwyP75xdrir
E7wzk4wrIDt30Xaw5T9j4ATWpOi79POmrMYzTSXe0/DsauyUhn0NSLwltHvth2Rq
eG+qcBOZzBDiPC0M4nwmiJp9jDyzHRcT04HyMtlU+oAzMhkrixNBgSF0Gx5KZn01
YpW5UKnxsv8/Nk24TxD5tao6cXB9tP+WauQwNMJ5HesyN3X1wbX2eYj+wbh+f+ON
xJxAOwNprY0lNXcxUTqx1YQXnCAqrrBM8agLJNOFR4LFfYkR1fxd15+nntPK6xG3
L7v0PaJAMgLbqm/CtLtQyS3a1BceutmXKm8r/IN+o++bhdt+UsNhce5xnIlDaFtn
WNBHDeBi/6g/mn63oSlP27BgvLHWJCMQA3sf5o9jTNZe4f3WQ4RUsULUjJTtM3qD
XsIaG4ZHgPc4LG9QOEQ0JoO1YPcP3HpNUnSNAqZpoeaVJhPnWJIWhVJN4s++UPYJ
Y3R7eclAyA8ZjiLoiQXJvSQdGeereLUV2EU0zdiz0r8VyrcMzcHlpEb9t7hYAXN5
pn/iRPo5w0pppntRjNkzp3Ts9Ndtfo219flthfa+lrx/EKH9OfKMsI/gr9YgQTqb
kw+7qIwFD8HfXy4hS6pP+WrARToEbFyKpG75omVxuB35kiLGNPqpN9Hnt4SiG4SN
IvUS7hXgUy9yWg7HQoFaorlxkndTmLQkz99m4d9BmaupxIR7i9rjdAnj2fkANRct
scxhk9kSfnlJfet9Y4kAMMWmzsAD++cszSyzKJrrxfY57ZNHncYletQgqXUSwyi1
4iKMYuE9F1Zm0kM+3U2zDuHoUCjBQsI4pxnW4wAQPOv8MBOBPlJzdXd2ceDR0Vav
22y8W5u5quBFIhnQXH7hGNtsZcmJLtprCMVJ3dk1ufHdkwtEzpu+faFUJzdhbvl7
64X0Q31sjF+6BJ1n34eazG6fDPUaiGCg5c6fmzcHl1u4sr6xtGzN1tRm8M9mmgN7
IdpIxjRg1N4EjlZ8ACC/ow==
`protect END_PROTECTED
