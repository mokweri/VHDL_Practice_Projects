`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/41oPVovqLSTtK27BCyHk8Y137dqWle1KYa+UqfISwZy/IoT6RBI+imRSrNm6Xwf
VQeakoyfN4Z3LodP3mIxvHZffMb+NdIS/LKPLZv/ohpzs+n3GgRoPO32NCSZH9oo
LK+fuSSbJla1bi0hllf+h5orjXqGmu7qtjbQZ5Ns8YoaM493P6j9fOSPYMpDpAER
9RbamXO1NeZouvEBJfTa5+kiRDnCbfbd3Ei5YUJVSyMZXbfDdWk5Khnpkr787r5X
ZxV65WoR/xYvmHcRzJFSeBZ6AF2xTRmGFctuT+8h/fs+/QBPUp5ZtOtTaKZkTcQd
xe/mWcYQNITwZzo0g7SrTIhjk4Jp7DpKTkk4M7R9KuQvjo3N/4zRFiBxLDUUyveL
OnUzjoipadnre/s9Zll2u/khZsstaKunLaUDxoaT47k6gB0eE0xN6dAyXM0OxsgA
xJbsNtR/FGAzjpGweO/FfMiLxpI7zZLQLwjXZnpsJX9EuB4Hst3f8RFqGkYCjjLp
/LyLIe9oZ07KC58aojBqPqQXuHnTTZ4ty8gWFDkauvyYk8B4H0MQvZ5rYzHCDabZ
WQAn7aiosWjmF8lvu+HNbVqJSACG7CE1G40VLdsEpSdfYjWL27kbMAGecLS9SYZg
yVmj5M054u9iuOslffx1eaWH2we2t8MPUq74qMgg0F/69GAgLEg6bCSgPa232ipG
Erz63s60Winn9SohGCRkrkVVGEZ7p9Srre59aFXVFvsSp8ogNu01VqmfTLQbHCWa
aLEetSyFcSuL0STpBfyiKXNWDGHMQK+zNi9XUt1JtxV6AxyltsvAfuNPLAg5yL7x
sww2nQkqhLAX8k6xlxCsnuAgUMpvTaQfAY3msu8eymW5PAi/cia9KWdT0RzN4mkU
uIQJJlP3W8EGSbms8UUUHbilIsbQcXx/I9e+UH6NYoVueAQqoQGnD4mMgX02ckVi
H3xhCw401w1G9CxL28LMpFyMRovReJscvLLOL/OeFZolWlDUfpg8PPLW5PL6osvo
yKsDUE9SKdM/18/UWWYLzhNJgkJXdBivUJ6gZMJiUdZJUnlqOVkmZNvMBvw/c8I9
X8jb61FW+f8ctL5EvzSr23biLv7Jw47pVsrrK+io3V6BE+urMv/GvSSAW5EgQSxG
w3Oa2dPmf2zyiiyIQ907tiqsTAjpODgCrfUZlbGwVqxJtItII1cjBxxzL1WBCO69
MCtb3BFM/wCmtgzReJNWcd74uHuMWKNEa1nLeUleE+c44VNWbgK6s88L/8B3Pulh
`protect END_PROTECTED
