`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14mXR//EMJ9uXWEnSHMifkUQPQN59v+pfSu5xF0IrsTKNxYcMkCRpwGU+7s7WZbx
EBx4ckMYXMD5aAGd2GH/zOQ3lZ/GzAXwXJThiaS3juw6WgF5NWtdBNJm6sYmGb7B
OJvLmBFVc15LfgJ9UxTNo739h/qUCXhjHhqMSHFnYgvMXGG+9WjF42df3ohEVPMh
AzS+WfbrYXq038aU6lkLgh51UQSChRrs2pPN7n5afvTHkVOi1p+zKLDEyqKkhj9e
WY9AYXMFvniMs/VSRHUv+pHjAOvpK8tXH6OqaRHwoIp5M0wk++EOIcq1Do+yo+3N
y4oLOTr6dAYokfCIVunYCmyXbX0A31SOiOfOSAl/JmpOE3Z/4uINOsBST58YO1Oa
gTLXHEpX0L5hfh2pN+eRs+Vb+3PNJk03ibe3Kz+zTs/fH+RiCViInhsEQ0k4Acig
rttw+/xZ0OSyw3mVyjcXB8wda/F7oWWnVnWXN1YdggAfuydHlakacserrdVDlG7A
AE+jCH8yXg7jC9zaVy0f3XCKnHFBTDj6DxrI3n96WIGt7fHbJjdubSAXmQ02aMbE
nEALBLy2QfrYOM+v+csG2mTYf5qYyqGLBNMMbLrWkanTGtyz1HGV8ulxnaKmc8H7
vNfqpFJF2tEqBhMi7kLtFo7hmNf+8zyPDB4VOjEOJdpl3UOACRje5mYIR3GmoTtM
pt44kadyHC+U8cOEPTbOFrUSDybLU+5v32ue55ZJlB1sJR1sAYbkEfsGWcEhbK6Z
XWX9teMkkqZuahYcpjEbcwSR0NkDUQv8so84etK0GDnbK37IiaEU+GAC6hkJuuLx
42bhXqRvucmdWpk3E9mabZ2TO+rvkGULT42/j6x/80sJ7WWy6ZUgyqr2YfeIzOPX
XPnEj13dbvn3OTbwMoqWGDNOTYpIWlVRbmUU44x2GVWb4FGper9UotsWsCFEsOlH
ecAkwvlUiYX/+Bso37twCSyFp89oL31CKbgOeXcr31ASz+zSh3A5Zug8T7LtNJ0Z
BW/lVy0hHUjqRZ92AiEW+dghta2S+GczcC28zlBc8ekLLLBCwsgN4LMVGNylBNnh
3bUncRM/ScRkZV9rt7vCEMWP/TD9wolFfm45jrpkQHbpPDhKESTtySaR6mp0vYf9
HFKlnFkeEUfgE/R295sDmwnZ6fltt5Uczsq0316qrEQFdkMpAYNLhCCFH51TCTIv
KTWLe4zNEi91cn16j2dLiJOup3MFjJJXTKqhgxz3byeWeDCbQOrbr0G1riVt/sM6
+Jo9pOBjfLhBl+wtv+O59v7nObxK6KhNfZXxUw13GCWGaASZb7KXHZuTpl6g3lTR
hyrFozcF81CIybuXcDF6NPfyC6s67wzUo9a1NdjVa7LtbCWMsMuOWlTF3xPYYbri
R31OAYJ7JP7dgTRrwYjVoGRMG5Uy4wjCztZwZcPV6lboF5HisWqOnQy/WBWDkhIy
mHe+HN5mZWP6fIDm7s3nUloEIs5EhTa4MB+/Wmsaxr11mAWoNqyS0qPwjIg9VdMs
5XPCQS20JDAWX5cDPCA+MDmKZNuW5AvgCYkZHK8jXRsGtINuoDho3MUl80BsNaXi
QCx2a1YKSOrOock42tpLSXaMDgK712Dl8fGXU9IHXvnYZq0RqetayIMqCyyUqkJp
963A4B0iRcYboia41K7jmnQnkFlsqeW7Mc50abBCLBV+pE1QNRrw9icffu2ygC7/
bDCV4rdkLrJTDTUUSo4nUhUp7cQGe/A63ti/yOcTwH9b9XxeCg3+4/h4pYaNiFo6
jn4sYj09/bOywhEZ7rhKP4IfwY5bYSW+6oJw08iqtGDcqDMA4bbNGGuY0wo7vpxv
k2ESd2qVFs9GPClgAUaTHNdHDrH9DFi70f4MW4FkQioeu94yBoKxYHHH1JSqZpg7
1i2E9K17PjpvDfjVOMW0RNLhBRkqPmN/fkHEWhAoJkXeAq2IYZcAqoy4g9wU0/KT
+9vSGlXaPH8qB/nZfhedlf8krCkg9OjW72PavjE6hyCNcSQu+PPwajNgua+Gm60D
Fnme4YTkk/5Nnk1GHmbKhPS/OZdlWSPNHlo6QPz1BwylMrZcFOguKOHtWHecqldo
haIrH1z7pk3bVaH8ATN+E7jB3xSXEiub6y6gg57VlIa+dVps5Ne8Iq+ssHCDH/DY
RdXy06NTnIwM5LKrzCfJaicagUUfIRkszzkXaOQc/aBof5NdHKKCT2WQbM/9jbt1
ZlayNZTrfFotYl0plx52VQ+z0KuEvpwCxBBmOs3cGJIBeGc7Ojy3o7Co8B0GsrQ6
C2YBRrdUokk/hsPnRqAdgA94iSlFUXnx2rumF8TN8lUgPsgh4fBMNki881YM1fiE
vHDOaNhb6UxkAjKnFVO7mQ==
`protect END_PROTECTED
