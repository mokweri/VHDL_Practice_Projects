`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FCcyhXcpqhDgyURqVxfEd6AaarAUuj4kkXoYxPBnVg3MmJz6CwpMC5BtDx1/Lrfx
qrP2F5lI44E+eejCaY70BQxXj/iAhwNydJCWU4jcx2K10oHHBFOCxMWsOWYNaKrp
vlC+vt20mNiNcIa/Hxbrptkk/oaNrDQkcWrjdPun6FnHRLRwKwdmjpt1DQYdFU/Y
eImhmxgNbyX5qnqfaPHHSBJjxstttDLbg4cF4kCK7w3f6ceV8n1LFs+7eEVkLeb3
VPAzxdm1HlDbr2TEWqiAVMwPITVCSH5zDXDU3Q6YB5TS2h/UshEmpUZHv77bTNB9
/UOL9mIsPfvM8rGpAET/z792iY7CEwkbaFuv6vSRFwMZA6RA3OOMJQeDNyqrUgw1
MwYj2pF6kstZJ4bilG+iE7ycRjZ9MbO/C8J5GFDoKh2wRwB5G//VeSExQOwzYBpq
ZhsFSzMJbsOpsORKAP3sGRjZQZeyCRMAHmIlY7lqnGdyXkwHV9GE6pvsT04GYx21
LMhvAeHP6fu9W5belZ7invRCE9ePEm7UpAEnTm4j8irTyfCFEJV69RimX8RQzmDu
5IgmSMMpzf1Vi6VQha1kDcOlqw/F6rugEpqPmQspmZeQPbTha1IYtqa7TVKexxsR
d9qi+9LLvZxuROpCZGSdsEcsjhPcBmOegSUulutmHwflSoCWKvkXg7WESesbGerS
SNyhgQDQ2CfUT7Ps1DFuvN0ItHhBAZUlaKZDbzd3rhJNkAc0Ca8e1PsgKwHP/erw
0gaQWAtHOFmWgk0bjh9NKgreUVOKCyJzbLNSPa9Bej6c5AUmDSr2nsC8BMg7plGc
VtJBPLLcC0tsy51j7o4KpbSsVui9HIQC1vYpJXq1t5OCW/iO9zrE7cZjUsEURaRk
9UuN/2Ascc3Csc47r8a+KGvw4xPACZCtiO4uwgaGrGT4aKpxEwDV56JT0COab3bT
XC+k2TRrPTRtdOXuVwIlIFpVyEXZBuh/86iMSx27UOC8S6fqCY2FG4fnM4cHITt8
w69cNWxPfzl3s95qqwbDsUGmyh7xwX5TSmtrXg0PljEcdJNWYnhe0a6fqX0FVzKc
ZKXp/BK2fwykKHN+jmcWSDNhcGNGTglvUYL6UDoDfQMJWAR74YLtS/Pxfq2j6Lfg
Hgg6MQRv2XrIcdjA6XZwtSuew9G+UxecCJtBHbfwO02QDQT5thcmKydagDW+3VIH
HkOVM47bLu4+jIY2P4W3SxnKTFud7GmoD8+0En/Pdudl9faq5t/uqpdcXJ3LWEM2
m0FqaZmfp1tdO0Y/7ORcZiSDHi1uLxpvaZbvN79CXvmQb0hxNV+exysz1C2ba1ZZ
FnmEJqDc/4NTHihgWgUoAyiUvjm7IJHcEvqbtozCzd7T9ly/6b2k1UqtZRgVr4u3
ugYFB04hhj/+tHSbLqkymYi44HicttnCsEQ8LDhAhx+YTI6MTOkOuXGrXv5ogth6
tgj2yz4AYnixryzkqjgYlsIrv3pkkfmAiNpJ6zImvyetiqqI39ZPj816NK8z1sTk
hMtHUwkovQa3Y4tu4ZRSvlm4fVc9iIRTLJOWcj1SsCQGI7Tgu72goC0mgMFcxBQo
jWSRnErYaGlQZYibBHDdCGfn3WR0stcKSOV0+ImmLUbzcQ1riXUm+AryoS6rHowS
Ba/EZqYzVuz0/jzZ73YzbxwHR0SVMYdN4GNwjJnVA0JbiQFzC6TaKpxG+brd5k1+
qIBuSkUphxmJaYuioZcp/R9mo2VfUPqEt5Q+3BW13HZCu5O4cS1OVbDBaNYL2eYw
szYUdxITCfjGUvZyjW9tMq2xg1AD7RPLedrDTztMsc+pywxXj0VEjqztmNRMZClO
CP3GYnFhEQHXJn+bWr6Mgj4ega3p2fxoLRlgzUndQRlUYusUMaOBARQkXri9eSVj
S9l/IzOameamUzqs6z/sxHws1PBE6mFojaWMYD6fHZ6pq73vHuS9kE+zY7b0Elk5
gFzmGMD9NvZFYc5FYsMF+/dOlxhXg/RSAROmBepCn3ejow/4gCwSvLr1oDRa+3sb
wpCYmj4e/GMacfRIUEY3G+h4g1mt25jUimmwLd3Es7iJBkoT7ulvf/HRm1HiOZ5I
oRnie70pon63R2XneD4VnOMGSgXZepPZRjCrvDWQ2ez7MSbSYFIfxfxbhJli91wn
ZdDmoF0GEowepHsvpEkSUxXD4RKI4Ty+Lf4oBnOa46Y+ehc0/4FPsre/mvbyvVkk
gg5356PboVOjLkqvvk1/XdZTIJ/5/rAYkYZrmiS86GSWhL9VnpMy7eeRVh8r5aV7
kmx3b+4n8/xTjnFhwIHgLDwb73NxJmCY2+KOlE7oCcRvv607hTS96WicA0MKIhLA
ZPDjdOJFwi4RZndmxG4JvpoC799hNlS2ygQfTLCLp7MgyFajPmehWZ4crYIU/rY2
jQlX4vyFUsm4vZzXPw+vnmXJ6qQlLv8Y+CkrRLqdM+bgar2JoKpSxam7ozW+Pb0/
aoG40dGwvpyYVKya1XCdcO0G8Q31jpkwLU2Nn9eLFi/o09XKS9NjSVSQ1ZQ9/4wo
d9tp1VhDdlwOVe0a1wQ0daTSGoUYOOzXDalNks7o00l5QDQJkguoszW9d1rJBrgS
RGetaQjzgIZnEOJ7moC2Wag7VxdXW62UqED3+JTZE3EgPkJZ76ijW71I+rFFvCkL
JPTmq5kOHtvcgbbJQCPszD3uJUOle5poPVYzLrBzxuf22oxM8+44cpLdqXMakuAA
hk2wlOqA6bkwvlrCpMq2WPlKniVU5rplEkUOK+lzxBxbXTTBhgYvKnIuPN4cyolF
720OpLG2XoHlL78x2Z8p1u8ed0/LIMkiKrL7aTW5+j0BcU8y/LkymYzhnWX4y7Sh
c0Kq6twb4tesxSjxSyLeUbax4xTEo/NUo//EVxhcqWDM3Daxw4CRCQm/asUnYUB7
fsj5CGXdOe6wBnC1CLq6R14PAL6P/YwMi3h6SVSks6UlscceYYLLe6IeBiMYJa/G
oPrZ+g2Wgkais7tqEfgb9B+kJk42LIZl2XVrshLKfLDsbY2JixzDJNgIISWmDR3V
HiRAWJTgp+IMmj8blKNKmhquE2UwRLKb+V5ovSMJ3jis1hAbccJnSY8BrKq6TWsT
RydZJWu2AUcOn6iVDpz1tVHKmqE0Af25KIZVf/vJch3S0nCbyMH1Jaw5P3HkesYX
kA6GehMRAp2eaellXGV8Y1G0EtPtMZiIUr0Lctw6MHqsudb+leuz4papaaeh6lpE
v6QlLpg1jYr5gjdCk9VCkNidYZdQERqtPjNr2n0G7jKMAnEb98jwefviGdOTGLqI
GOISztbBWcfjeAWsMSm4a/qMtbyOcK0YSrlqEFpDpw49dwp7XfHADfMK4x8g28WM
n7OqU7Yvmlc0Y3lGX5iKMm8yiAsYQt5+EzCOf/toANU2ilBGmXdTev+6DGVfFMxu
NQoYemW2jl6lVuLBsWEyMWhHS1yLEUlCs2SUSclClj6I1MrhD8hNMFq+KwD1GzPH
qcTRXHIJrIt02zcT/u8bkMDE7KMhZmK6QTUgbiWRJS4ZI+GriyEvnmGitco26iEz
Ibk4qnfxn4eF/OmpMt+PnYun2+n/9ety2ukBvPJC2vOwBcwIGcogOWKKN1QqCJtg
UCTnbz+KnyxizPRXXnfZap/Xg4ChsHNh/b/+XfvVXX6+1Grn9lYYEyFfZTEfTlP/
9bWadI5bQogckwKAj5FI2EhT9/Ft2asOXNjEbGncuuUTB83f4+QL8G/QeLBAlCrV
B4rSWYH/Ps0gvkbLhqvcRESlf4IglQHGETqPqHYCZ4tVTkBGI8XDbDBZXPrtMNCr
xPZB/KR1Ox9/cm1m4mpNJNz6DRN/hpoUbPJA7i9h60vMeIxO9LLUy3mB2hDFPPIO
Uvgo0MXjwoxI65wkUzooZzG+cTs9eN+6KAjZPBwYzEFGZhqxi5GogYScePw7i1TT
KtI8MtTiAobvo2JkLsTgAKfq/kUC49JR3RgcxvHJin3h1CB0vMbvORCDgEZcG9ty
AejcsJ13E+T7Z18FyhKVhfRHx568eWE6WgquKzlXvNbjiKo19yRqv3uLbJmQNbQQ
IbsZ0Khmqak/JVe+W0d7jNY6B3EBgUrMKxJTXzjPYnwFj87hGieT8VmFQuT/lP/P
uurNUrUKaVphHzMd+jNwcTDAX1beB31Yj/AJ2KBlfHtGJhzJ18X211yRhp7omtX3
gF6ODCC76YR79yqIpBSx9W8/Hg8aTH/zPRyusuuiT3FTxKIuaSNiQk9/q2z6NW22
cePjT72SBIgWnicTVGgJdWlOPAWkcZH7w8QQUgB8VaYz9rStubHyNCIjme40/9tF
0J/QwRaksoGzqQTBru1zjUC2VRQHYzjjGToGfwKiggkhlHAaUe9gA361mXantPK4
R/H4Jmk4R75e55dk9diJGfEDvyCYXN8QZQ1fdBuosmiEOJXv7+ECRjSdmj0+/a2O
W7m8YVTKlY/fsnomy1axXMihPTW08+apF7rLV6j7GGOZhmTOeqIcWkzW5EE9z85H
dbmQj7aRf+Gndlpi7QyAZ+7xhErnnko1mIWHUOb/LmSjFJ/js/cVAPa8klZ67LVs
G4k6lwcDQj3fcUxlg9w9MoG3NOzdhiK3ZeZ4W7MZJClF+Q/3nw1FeC1RM3y41zoz
wfNcbUWCQ9OfI1ZXc8fdlgc15udRCF3vT3epmTh+UBw6QvECr/5XlLncb8VVy+jk
6yhLAEubM2ejzlHb6Sb9iXOKh/7q84MzDGOkSYdP7mLk6WizfFGhyiShTdKY/g8k
0lS6IXWoZsKeL0YhtdJZ5WrJADB9uO5Ud5LlfTZWB8M/Gb1fgQgR9MKRzmmRC4Jc
wC1GFY2Yt5yrvTBki8kFUi3uGFsxomWYDPeKymGbFknO5G9e4hgh/a7UmSOsG7gl
048lHUBOlLjwAn7zWdQyxAHz72dE5GnA0cq0rrEiHxKzbm0QWJZdNRr2M3vc94lk
uVagmFsZR+rZwi/6d8NtolEFjMaFthm0dPBJY/Dwor/Hjf0rEzFD+JEA1JXKl1Zn
nfsZ0szMPam7tagiuKhyAz0j5frRuQWWie4LhTPrAaFsfFLVx0dHd1AwGec6eMf8
fFcjM7ClFK+CJLDaQmZpsGcBG5WX9o2+pm5ndjX+DWshG9x4IGV8t46ccDrCVCxG
/r/Qobmo3sgoGb+4YdwYICQgQ0H3rZ4xhQFj6j1oBtbZa73ERxd9mpG/cV5tjCyA
JHorl+nZhP8Js12062+sDO0yXMTQcR262S9ML8cTvJW/anOAm+OWW/bbjFptxvef
DwoCuoUakhmoQOpum3hvbxHvKKeDIZ91KNMqNstvaitKw3UQt2GaDn5YtY6rgMzF
wAoKZsl66eI4xAMoXGWhp26iRveON9o8JMbR4J2ZUxfp226g41RWQJGkG8IHltcf
bATFmTxLqK/cfuCQ9cA2MBzlmgkhf/zu/ZgyM792DjddMDl2IqKB7nLmqx5gpWKm
KmeySI+GT6r8xM9w+Sy5Z8Ties3kblZxjjwGhti31WLNiAL4B0SL3BIk/uiNF/90
XpjaMxnhvSSlLS9LtFI5CAA5uerwSd8PksKLDmonyFfkArhT6RhJj/y58oBR4U2k
uJBG8+B9kJC9r8Y1N14WD/cQ2mdqvVwknegI7rF3Ib95Sr2NFiCUP1jBjoiLO100
5EBhQ8sRLOMmmif6t4UCCPyq0p4FnftnNMxDEclmaSJ8LZh7yH6O9GUnHa/I2CGL
u63qF8QWDmzq8PmEUl0ZeMNPwWXNxf3qEUnt17fXGZwzXrup1ikijx9qN/ggfcOh
1bnF+onUWsZCiPsTOTOlPQ7no7dq5++0brW+7Hc3cOsQ1eEzmtFa1HgWlTtBSBk2
IE/sZp6mO6BRMaRC+gRe0DgPN+g1RVirQRv8QPZ0lbv5DGE6MS7GGcGuvzZZ4Xd9
j9HNKwb1kqp8AVXYo0jV5KkF772GBhOLYJK+6p9xR+ibQtxXoDEhcQX5hnuA3yh+
l5ivA1B9FbTc+KhYdjW+Rw7UHCfn1U6vnLsL0ziY3khQ7+EAW6vpcp0BkymakGjK
w+EbW/sVNQh5ozbbs2xPPXM8dzsNCMjpG2V85f1gxPE5KPUUqOYzMAQgsFPLAdYU
16F1YAqJbfFuwaUfmXI7QANyoBjfRaEgnLBiSsFJidmtsivtr5weBdfTUJKY4Gm3
TRj9WYta9piQeOBk1fghjf85Q/o/15oFpFuJZchAPpETSeXsKrb+LDMnqLIP5TnC
WjAdWU+h+6AFcO2G/gnD3SLcKVH5F/Z9zvZPiBLqF1UToS2IrdRXlrFLR7BLzvrv
SmLvkxA1TmjvyCRVVMdppYOaaCN1uxUOITwGxjyR9e3hwGq95PzFbovINAd7FxFk
vAFlP6MJEm5Axy2FxZj0zjxBcnqpzVBrF6driV7SlK5T243uFjRoVAS25kZmvYyu
HwVNRs2PrWdQXOVCnyL1rdIj4CCfpCcPZ/OWa2B2Gr1lCsNeK7N+czEpebtGLcfF
MIwnzEFUxU9gOQwqFxR2lLeXdjwA5d0eUxwbaKnAlTHgxyfkG4XjI3jDZC7bhRlF
HHKbu7uqGfbtOmLdhf8kcDU+fhlkytpEpHQr0gR1iDMP18n2QrPcsy9LH+YUQDup
vRGXjX638OmfUJNsPrD56KVaAvuHtdNB5jKhRvJvw5dxmlWIprTKXtHuaf+As3Jd
Vg/6jTuNF9plVGz+KjuN+WYxMn8u4tXUcygw7Faj34Rp+etj8WkYygEVn8xFWogV
phU9CefehUdrwvqVNrEsP6nJd0h7MSuO/f8N22NwfzrawbMBhvBXaruZp0zxU/YM
IJFoNYJuYaq/W+Eed715OUJiUQDEpHFhk7U5BvSYlp8Q+JuMAv/H/PYswPliZSh0
cfyRprW/PqQqzoTsrvicpQ70A0zBAogyg9I78sgD6phpCHVXc44O9te8WYDL/POw
rFG2xNDWkaeyv/e2YPMYmTN/bC+PgBCvC++j0T4kP349dQQpktIfaae6QEJd1glT
RY6m+moJgVRvxz5N2QjgAwPxFVW4s6wOJIZBHgCOESPVOEj9PGVJMxObHDO9ymnB
n1WiIuGRsJBB9T80SvYCaiaZKFARmAUPnsjiQsF2SEBMjoi4rpe31ZBXan/WeHmV
K99z2jojQyV0LXzRMmBq3GSrKzlYqr3FqlwTCQRLj19jSTGLJqEpJOIxqxMi9wa7
B3VuM+5TFVX3j64FzQbyOfOv7KaL+TNibva2NYDZizfVx0LT3u7TRLo1Cw6H9Caq
Xm5+M9ONYIzP1HZ9HqN7qPqFGKrPb4mT0m2vrQEY3QaXubKslxr867N2qiChK+h8
S2woSX/lu6IwP57NcAefIQkM/mVHSgMGOKGnXKNVwUXN9cRPGfc1+FhIzsxtrt/z
Dm4exChkRQRGywnbkL8kh4UPgrs1U5vh3CmxOSFowxS7lgwR+yw1T5RxFvZ5fMTT
H1nsM9vqbIEfHNy9Xw4lBDLTUATLO1RAaVLk1sQ+iERHlmgwG9E9nRlv90Ax/rr2
Hmllh4UoeQhzRDm7AvN3A+SHbl/FbYORbtD6Xx5qaP/RCo6/6aaWmymtkK9+fCmo
J6Jfq9NL1jWHP2PSJ5r6e+1J4fMjlbUImYRBImzCqRRKlYcvxk8p9gWMZmf+NM+m
zIH3a8z/DynhaRc/N8lkv0OmmlNI9eKUrDCHbR1Yr0gGzTSxroao5XaDnE0YbJQJ
uyBLL4XWolE65SchTdEyu+dBljyIaXUZT86bBgBnAu73IQya8tWT2kdVlMEap5Za
AWMGl7i5Zgaq0HxHWmHWczVfRPSdlIEEZU60MzXvkBtjZ1FoZwEN+jYaFFIArvzK
uL5tWWh5MeLG0kWbvSVtT8LD56eT0MC+S4PAEihpKA1R4L3ifJI8FbdPmvWCubRL
WkDoqe1rmSWBQorEZfZ+1XWKLwrZLh67FazvFlPl1635mqFpj9hhpegVRRItMHLO
pu5dSEN/2ZNzp6mua+quXw1kqRM7pXhD+dnZ+XduRi5pXoblEiLzByElCzFUJNsm
683Y8qceS6ePz9wLRD3ObIWa8p/bAqEG6h9+uPsTQnmh4TmvMyGVn/DgqhYEaSgS
uFFn8eTZp953WdQcQDwoIjM+sD0dm/falP+cF4qVW7gVPlKp009g8QW+DBuZFPP+
jcQZknqWpSY6s2/iwubzkNCrVFW1RBTd3prX/DEc9wMKZ7jxW/bokTbo63j3e1OO
/n2e+JRvkezWpHZnn/pzqHmp/lZPzwFbOMyGPMwGAfCxNREPrAJBVBEbWQnK+l0H
MBWIMil5cIivZp3XKympAg4ncHyVWQb3uHFk/eWrHIRRCQlb2uIz1zdsVCHFA2yD
gbPBjCdbWuY6niMfFhTgLDBhrpVVtTLFqKRVnWxDSJxK6IBN0JI5smDAhXA3hLUo
/y8Ccy6JBiqSR0ZAf7CmWJqlJAM1ygmQKbCCTaHRHxxjmtCLcv/Dcpu5oKwL+zMl
bW+9JRXD7D61KVjzemIkASNFdPK8KZWbgjoLn8tZu4vLrNMSE8XwJOYt1SaLLk5K
XkkuQ2oP5gkCzj7T9VJVVq09cnypFeRvIBJSZSESD9rKn7Oj6Il67UsAknZ7tzbK
m7tGE5uR0e62ELLoiKtFNNHWVlRICnfNpuhPlAfvlk5JI/tAeSKser+VSF/Sq3fT
jIz6hmKFUDQFiE+54P0E9Sou1bA/aK+N3XvyeXCQObDwHijJWG+5ayatkBdab43M
bOP8NLccLA61Dkoik+8xpsGAB3w5URZ34yo+XdalLoc3f4FYrtCRi7kyFXdCw/c3
66oC76UtGQcGnZ4Fqbbq6aiKZRycpZkwiYMvfRnIrjeL+21lrCVMSnJAf16toAdp
h8ahZTE2ZJht+uyHmog1BTAZ1xPMBCNm1Xc9eGV1QiNGzWET8xzrPJrDH1dwY1Uq
nLre0ij9aaelexSrYyXhoUDjyJgbXXPbAij40Qt+5CmP/8Dyr9lfsAvDuUzwO6io
qegahLaDAlVhAnQ53VMSq1VZ8tMDxtvMbOTGqThXqCh7YiWRAiOjR5m3D7GtgQHL
J/WYxob3Z4qum2GxXZinKsG2B0/hQnYd0DFgXHYucfMn0v4zVg2bhXJ4hJDCM4I3
huf2pD8VRrkAzrHBUUAnUBwkBauiOWGeeUGjIBRYM24vkk3qEayKNZES7WQSguHh
hZQMMpSp6/K9ADb9kf33qWcbF+yCsORflEUscEHnwbjygsugSH3Tda84EzvAKEkl
OQ3JIYZ6aA4QR09tbbxyp6Vdz9SU0cqn4dvA1IumbJR5TBe5eoj/ywoJ7tv3XHPY
A3vgCVVom2wUq4islUgS6WzmZQiEbsWDYzsnTjV1AGbZjvisrPP2ctM3HnHfb8Zy
5rNlqC7VrbvkKMiOoFpmmNO/zdPErj1gf3RH9h9C7VMzAnVnv+Xd23al9D2Fc1/q
8lXZwOETYItOZqda02d9yTC2f44jKyrtPltGXyaToXBgdten0QbbShYhoF/A0ElQ
KVuSKk8FCFoNA4cpDPH+IX5tq6aPxfNRujqqbR7KPk02i6xPjXUjqCx3qpS9QMxP
GDcaCibw6l6unL6SAoXzmd14krJIlXcsDxbOX/92/vhIrVK2kq0NL7PACK7E/ENQ
zYmif0yMx3B7IeQ7rvFHO200i/rNQKNF6Q/GI9IDemat5rRnbpYHI8HwMCZr7HtZ
pc209OdnDcyj1EWm4+HThi3CyNigUB76QReL16lqBSCNpu5izYg8vGbiteCW74Ci
z6GQvMDdCXXtpO9vquIklyZSktoxUwkngYZqjOeGoU+/0dFcz+shqDzZeasd6j7r
dcZIYoOVHJlFy+mge6B2bY+lAo9NuQ3QEwqhn9x9MEglr9lImdZxSzpgug1PpBcW
f/WUHXlbAayz+LGU/lpGgDPumpGZQImzmPDVsHmz6QKXtAydfXkumYT9AcnEaXOd
4u1RGZi/+eDuO2xl5rWXWj0IegqaBOZf1nSOO7+x2CxyDXmeGx6YTkRKUbroyrbH
tbyh9XvbCQxKUWbD5os5OHizPsWQvsuE9vqqfe6Z8vWMB6NI74+41Cc9ZztwmKdY
qTJjJ/8+GxgBw1XR9JM1PbNHr40OUSyMx1t7ApKn8MQfl/EaVgtFacXSycmMxVGB
09VxlDiFgrKRB44/oANGcP63SpkT6mwXxFG+7Boapd6pKTHeaAOeyK/ajhCvaeD5
BaS4gEUNZzEqIkhq81LL2h0k8eYBB75870pyfRQLHR5fVI9ss4aQSrF3hul7Wgux
YSkV3KFNJVHRwWAuBZI5/P6zwk78wYY1uZ2BFmb/YZM8NZ/FArtIxsQxkCY9nwun
OmwWs1sLZlT7Vg9UbWeN/AsN1E5qw1seyxJAkuZIurtvp0vyBv0PvVzlcTZX/NcS
cF7Y4DfxnZzuZI3zpXwhIYCkRA4SjpDjm9xRhkxhK51GZHN8sjWEXekVXnjyDV9P
eQ2sM8Dydrd1yt2VdTQkO//fo7m8rJNW5JedbFbssiFJJXDtJCvXTJQDQLNsnznW
GGyx8jMLKlwqf87ND0Uj2kncMOr0/aRVR378zEP6fyWAsZ8MSvNMAwysZ4iqG/QQ
JXe5A+NGEv6cjF7RR5iO6RCrEdyRDRnAvgBQKlpb0RWlTZU1OAL35qyz1KoMN8Ki
Nks53q7X1/E/aD6y9LhfBEzitXTmzgHCIDl5li8jRbMuwwbxvUMxDpLsXcHBy788
bzbNXT6JMWtFJGM8ulDSfTg9pUNQTYIH+JWAwoVIWco27mPV3pwQWgaPxy1Gi8f7
gjZiqbR/6esE4MOGIvurhdIRuNDaHElEcGNr1mKbr7AHnJeA/PuZcVK0QFlDLLeU
5CXL85S0d4XHSXcmQbrCtFg9N9GiqUHo363E1GQ+4BZ1dGaWfkWb/dFV91xvUapF
m9rGaY23hXOOGtbLB1bL3qn2b7Oq3NO3IhkZrB2c0bNmCLd2qVe8Gt+a5+6azoBA
gf49cmzM3X7s3k9EBJyA8cXmeNTiSy8lANy4NWs0veGp6ldSOAZ5bbKbQk+16nPp
lzHErzpFI4pDnVOMKqffWhUoZeaUgsRxvJwixHqCkKwPVhK3GVn5yx/2EIc3x4l6
f6NuDvQ7gfaVQpi5hKCOslsaplknWNk/dVvh7vFvT7+VvWZT/gglLoI0yMjuN9J3
W+f0vFSGpQFG95z/kEgAviEdekUDlBnm/FA9JddaJ8tXFyJ9nyYrysAFUEHQxRDK
V470bwUnzJHPjeumYw+kss85KuJm2qwKhUSd0730KRuX31bDt2Feb92Uv6iS7JAz
80MVsX0JnozRNsGNtvmiRnq9N5c5DKaIjaN1IxrnZ6Q2wwsUBzba/DD2S7M0M9mA
QztoHtxvUbwBs2MYgwgSE7X19bWv7sGRrQSiMuNAWfzvh7wtWjcoN4Dc6BMvkRhn
uYeqj8OrbLc//ngHHpLFRl/PE47twdfQhkbZjGesYEpzqs2acO8uBL4sW8WISe2E
S+bgfrLaQC8L0PwqJfsv+GrFJmfKrvW8U4oeGft1gvqZRoUH6vDRTzTIfUxMPO++
3sgLzByss1dbrQ5QQ8RFQ24TjBwwKojnMR3rXkAjAY2Lizh8Mx99P8fWxTdJcB/S
d0q6SpMgC1OUSOaocMnz6m0UiiC9UKKE6zSghSd5Dd2Are+rNS+7jyGvsR10cnWh
B5MJVMMj+78q+W7ijM1ANkkurrcbALkkUC3rNbhErhq1qqcqpS+a36W2YZgOHt0l
ExLBy+IBqM10BoZELLEHl0lr37w+1/5Xy2QX5Yairp0J9yA/YqxlXaPNS9MzV+1f
vrgRfg1HmEkV1AoKw+J+nTGFpNaNLMCLeVXur9c8kWy3/de0BmO3azDZmVKfPNvy
kGuNAhxTgdvwpgRsQ49+Q5Mkwzb7SX4mDuZw1fKnbCrxjtNBB5JFZi43ZRE3PPfU
5aIdpehaHPzkCCE7XE7/cFbSam6tUzY37XSGxR6ohO5CAFVE5GarIKZbQs/SKwaF
Gp4ZJC3we410J+VwswQO5t8xVWYg0QORHpRSsC9rVYgQtkNq/TmoXSoZe9D3l6nZ
8YD/QRTZieHHr8C7eps5wanCTQNo27c7rMpRja7pu9cHhhbcAGOr4Chu5cD5iY+z
/vi1WvloPgBXInesLwcSY6v8yvT22fz4p6lbTmC8jzFq4g9Rqgfv43uLlhI5czPW
BD3/5iVkGPrObhLtKeQv75GXYAvw99APcHG/tY5C7iVIKQ3kzwAnAWpSsPELk3k+
SS4jmZiiYAv/NpGpnoiX3bjs9YessfAcufHLzB0p7K2w6kdHsbLN7T4u8yG17ixk
AQKAtH/5CmBS7wTlHKasgf++258jritoBWbYBgKYcIVxP2iBFkGS6ndl1KNV06oZ
A6adxk89n78YxVcwRfEslxtUpsLStaHuGKTc+yEQ9EwMylMpvuuZLr3cDg0OGI5A
s0JuGy3hNJeocwEEm805s2RM0QlbMDDUPS2ZYOOtp7rHlqKUu+PDEoaXD45kq2+p
efrjld5LLSYtvn+JFoN891PskMWo5T541ixtFoPM6m3Z+UyjlTZ+IKOkA3CvmLcd
4E24c0jv3kZMaEbEX//tNKUqfdi74QWwWGehzi2qhpV6EFu2NdTYSKVoTQsdiVcp
X2Cbl3CNYCBVawi3OEOX/BFQQGhuujDlcX1HcOqT1NS0cQWbQD5L/Ou+UMJTY6bT
mmWLnrKZKi8GKDiftuWZTCb1LKz8OTal17VN3DP7J5NqFwPjgiU1Ev9ecBaqEUt3
AH7FlnjyOXY4Zf0cP01BMIduQd2S6GOCx2kUFog6NszvwVAWQ3qxetiG/695hd+v
Pb+O+vFMQCirIy/lUu/tI5qAfBvTUq5HsNmFbyE2gZy2ODK2Cc0fKFc6Oh12e2t+
iy2inI1bbz/v2mZ73p22/EXhwa+POCo8ViGf/CciWORWNCUSA7yWpWS8+5LD36bh
wDkShemqZmQtMJnH6C1BY5Kde0wI5xOymkPzBmN/Raj6PPcO05rINIW8MIWmExff
L7VIDmGJZXqGHcsuJYztRCVy/9MGEArTZPQSCWBaav1NM3mjjGTAEcTmMCOxL8zx
KUHgKNG82ctq63b73ZFaOObScNdR+YpMEFUYO2p12XYExkKNzhAgN4rmRZW3kAVu
rYWmqmuLzXgsMWpGQu8UGXSQpL5TUPDYFk2qAOkqO4HcJCc/PtfyZzZpLFChXVse
75w3hzkYU6fJllTGxsdVp61hc9QgMhZmbJuu9ZdJoPCG4S8EdOcYF4YS+GLhRFwf
lw9Q/r2uce7T24QCej1PdJ93tclKbrRIPH2iwwDe95id5BVZ9RkvaYwckXCteMYf
qUIJ+O2XCGvV97hqswTQ1Aos8qM4RFbtyMOEbCF/4WMHrHY4i4BLcdxuAY2g1kwk
+WyfoLjk2z2yV+im9VlXb25d4lsN6qASv/K6L2W/MbhGie0EKZlSPKyMeFuwIvYC
DB4BeRK4NzuI7mD5GeQAFxW0mQ7GscuXbj7IgrckofWaB5AqTp1XgeZ4XO9qysGh
GRmpXaqi8yeh0OcNp0qxioS4WmAK6MUQZ8HtfnYkYpcFl0bjjhZxKSQaTAX+2ove
KLgGx+M4H+/krA+iSY3zwSVMTRA81s/lWY9yrJGwibkf3OGonCnTj9fASJpHfy4o
jLhLhquWlFllBL+1yhPde2679aArNUyS30p+8m34NvWM9Wt6T2d8BOvmsnejQ9vs
o4Uz9odXESFc+PjJGwu26a9L2hLwiJh0OzJsRuTjZxbzZqF/bdzo/rGZV9ezhycF
c/8CJmFuyMOr0xyZiAi6gWoMiuYVH5MtfmxBk4kS4Z0XmTn+2NG7TgjK/XOinmPU
JgMRpf25ONxzp22SGyt6sbP2LfN4NZi0JQsHrSboF8ifvJCms6Lk4SqsDr/KzZKz
VUPonJPLMYCfqIdjyalxHW25ZgAzvddSVhYeEcBal6uIpfHMq3Ir0kf0Y3cEIusG
lM8xpbV2nLieoEZiG5EP6Ecf5mucJp8pEwNMqOMX483Fo9inPdSbXxqMvWPtCiu4
92hesTgrPnPdHQZX6Mg7W8/A1DqtuSldvD6J7d2E6LYSWf/62y64RGylB/2fszmB
7Fc6Awzi1oxGvpj75g8n299GMHqR5Y1HgOY7CV5ebHNqtsZ2ys8cjLmfoQK1RHbc
js5FHwyWZDuGXvlJZB5x3ZW7v7QroGLTh8LgRfAyFRwP3qkdff/hKHuqkz8mUveG
uTyQXQUGRBUKt4uC2S6i2VQLGLKHJ2LaRLtiSCTRITQ98hDkM3USChG7HKu5x/d3
LKWlFt4JhDOhlhd59/7jLcugrIAuN0D/mib6hC8bL6RZ3AjmoXeylk1q3fFHoVvp
37/LxODBDrzbMCLCnzQ96dsoeeKJ8zpjvqD8EN5oJPTsQJsshox11TARe4wTbCIc
yU04USTBb8HvnxsPA/RbIhH6ddHt8JgQp1KZrVAe9zHBAYHSHghV0bfGx02kwwHo
OG68n6YnrmdTO+GBGNVNIbuxU/KilwWT9Ij4aIkb9LWKyv4y2p45kxo9FeDzFuaP
VM14yFjmbm9OwA7CXjvXu8QYuKb+8i2J8bSk82CVkpSbwfXnQJHlV0VCsocR+Sp3
v4FKtbe9rZOHYPb1Oa0iZbB/VkMk3y/1IcV/c/60M1zIlR/onpJju+fPcISj04Am
4Gh/ea9FJeEkmU8FaZ2UmFUC+KbM4QiSGuhW2uh40vehizWPh0KsTYGTo32Ckbr4
SSQ+Pi1JmWnF7AGms2jywJjJq7XZtE1RWAzGcuSp4N3jbsla4bBpPbLTHhwMME79
TVofb+/+pSktx9GpRy6tsKxywmhA6AFMERMxDoxOxFDgfBtEOlvrLZrEktXqtO9d
rK8eOsnfUdn8B2arjRV2qE3AW2LWa5owSKLoiz32yU+ZdP6+xM2Hlqv2B6bc3CNJ
c5X2AfTHximbQ84LsTi83/4j7wsjy1R/9Li9sBCkeAN9XTnU279FM5vn3MVGsm64
wFITD6Sv9wZu+OyN9QoUsCceV1USkZRegchOaFXyxt7+7pN3eZt5LNFte1ZTVZAg
q98WhUjmtQQty5lc0/4NA94/GcjvE08yVhdFXdaiPwfHU93if/SG9KZVps3rB2Jh
904ug6j92R3LYCLCkE96faTAggZLnrfZKIsi70OHHutQo3OqEIO8CYxf3DJljMFZ
NsKIzLZP6kYPTt4NI6KrevlJ8n7trSlradIivFNJ1dhtqNLzwe26FKAt6rOCH83+
D0sjAvcyFAsT25mQvAtKdS2bmXWamnbvPha7b8WCkCZ+1rKl2eM4KMy53r23fkWw
xF6RFJd9VyGBcYmuxCgBOUevq+w6v/XGMAeQjkULMF0VdXc3pNobwp/WDbO2At60
xB09LlTXmm3m4LZj+VJFe35YkJxSvzOnyns1QHwmmnNJvkS6KzpbzqClvqF8VIdi
fO0Q8Xg5H3V1n1QVu1mULbZrhzbTHTpNamXoDF+vkdr/O6qO7p7oZdsfJ7+ey3Fs
pQsPCam1QqY7cksZLpvngMlvy0sp0M+lcvNP1buJPzn/0kDumdYk2Vp8G5qIzMqO
qyMO0XzFVnrPagP4boHxjI8X3hrIPzSEsfpgyRNGJeFfbl+Xy2xH5p21cArWTLWV
OaYUJ/S+70Zis58L6L8nI2x/d9IiJVQg9wPBUhGvU9eY5lfcF3hfFDbYvedg4hVt
mAomsr/RqyQinRqViSNkcZlxWda9igpxWrAXYFbjDIyEU65QQOofO8WrMp5sRHt7
vyG5Qt+dU7vZRPrn/W2eC9UjSBQxMicmxqTNjsAyosOo/4WKCOTzpfE1XizH4ZsK
WP7OYU01/w9/Da6p5MeerPejSrIFioe/t19cKrcn0VnyZUPw/Q0bpTQkIBf0lFbz
GKgPq5Syxb6bZEQAx1zG4p7h3KW5yOwciZRAcfPbz/nc+D6ybtQEBp4M0TU3zmlH
A44Ea3AvZmMOr8QJCYoVqP/7fATr2XAO2R5KP4MZ1CL4Sgx8HwunGcd4xKs8+EJO
0ALyHtXVRmBFGvshVvBNC7j2rbfogWJQch8LBDqn7IL0GfS0zCg+MKF5psjXnZbD
AgocSte20EExDFc1NIxYd0NhoMd63NTPcXif2lfnkfVW84HtqHO53/6aemTBImoS
1YnQWLGFRSp84KeUJ92gwwBqx05sdsoxRhhZH62xTdrbbUx48HmyKaXmRVQRX1t5
3qK7rA6E0ewSQb3Gg3AbblZsHvQE51GpcRjCliXQSNfveQQtHYbZ7Yx9hS2YRoO6
BSEpFOEq3jDj7QELRjz0iHN4ks2Q5K4PqTy+Jv60HJ33wWuTcCeBsc2eQRhhJkKe
mMSzj0tHJNBE7Ta4X0C9WrEiXWm2LT1/ZTDxVOf9Eh0ye7Sj1+eQwNdSw4TvUlP/
bWnzMFsJY9IygVCjgkYgyHamIvxOMzZtQzPXfyGSZiwJ6mp0SaZeoAyzPWnFYEGZ
bDdyzS4wo5NgbU0C3LgLeeQn9CGbz3BFyz3TuvNXq4eybUlSFBydDfIyziEq2t/f
8aweZgKZxg1XxZZJql9ijfY7ITP7v8a5fYZw5gNOZbSVkDF8qXVocpUWXpY/8tZ6
EYfQZ+d9LMtPVIXYfhINpGmg8BWQjz52Q/KYQmUHL5Hek02QM7pRUTjxD/wXI6Fw
tCqy7JB0vDRLZj46JXWDVrlzzGw3UBsMZaPz4A3yjv92c/+Ol6rj3Ig8gOtP2o0C
T2QkfwrILWzS+RVEcYvKap8VwK/PDj+s9cLp9AD/ws5eyGqwi+Lc7tAkJawLEwtQ
GprsDbeoHmCLo5NpLnsBmnfRhL8ar8JTOrVQD5f6AwJKIq+L3px7D+2db1FG4kkX
BJsYLptpI2rsA2QuuKs/uK4YL9Qh0ffBSxwC09KurhfDsbepz539jma/UfewOciD
Eb1pkSzqHHg2yXhaLZPTQsxjruqAn3EjYsOFdzzQP1p3jsWTThzYjAlgtHoqWAFY
rAZasylAIsvNnPyLd/wK8CDInsSQ9/BkZzmUhNBXP7txWafix876iCOmj1vGhX3C
5763bXhc+Ik6xxIBRFZ9wR0bcYvYaEABo7lnC3pAofEuqhllBLJfixgfaDLZF56f
4/5lKO2j0xdCQ9u1rW936rY+WjIBfz8dTkgEhU3jtvLitp+d5A1D2RhKWkzNRzgz
kCZbqJKDQWKEq7vTzJOTyzWnBQr9lh1lBB5KDczxTIk0fzmR3/rHO7xFOzd2sPdf
xkn/SOTrimNdggEKrapEehI7ZHIpyeul9LUD2E1i+YoycmAFbr3iTR4ycyD/D5sZ
+OOqcRwYcxwMIjsQjR0FFmlSMCfTKqWwJF/gVM2Ntrr519JrhF8Lczx1dDkHg4BA
w5M9pRbutSg826n7k7XWdAHCv6pST1rfQ707B6jmr8JGSbhHL0Fywn1v1HURmYsZ
EFJfEb6/Vwv+ZTfomB+hn4quE0iuddtrPW3baLAjjN7QqUbzpIw1X3E+UqTrueO+
l0ssYerUxJDlcdGFX55Zoj0TumxmaRCyfMNq4F5fsFWSZnJQNW1wjMNn0/H0aqQM
6YBo7qSQUUvR5iQug8Qgr/i9398h395WHC0yOVE4DPz+ubaFv2tM4K6UAMjXFo1Z
d+9mDINsxNbLrJmjVPUzizAtnZO6A+g2Asyukt80CbBcUh4+7shQRwtCjoMgOMQV
21jlrjOsf0/lGahWCVBp9QUiY6YFL9tQl+OGZBKmbMmg2Q9CptzuDVQ07DwgwRUw
Q24piwV4IyfbBNPWCoVLNkjbdWaDkkq1v+sIeddC4ETd9JNDIX9Uen4RxmLnWXMR
CaBvZvxPN1C+1GZ++oNhRQOfBwN0GcLbXdejBHFLKbS+0cRqilKiU1ATAj6Q89b0
S/f1mqb+WJ/P/vdCJzvrmy5iHFu9zdl6oNuLjT4W1RRoVpV7AWd4a2fA5hhPuK/J
E/svDUQ+dVG4ii8nO2OlGc7/DU0xSh7BLDLroBl/ScDuuenLDqNH7Lx6iggaWjpO
HSmXFRxGgKRbbcapD7Io6LnMgoLwIpMEj3v0aKfUqhNLpwj0derfdrnkeOZtPUAZ
z4wHbyFaevS+uhN6xhxnfy0FhFRU9Jo6pn251f13Mz6wJngfHrMq1c4/cTOVNsoj
Gm3vd0fGF7VZJ4mgLRmcxODCvzUw2NeN9vVehhyl50jgsRGYFOKkPFuNWFyQq/q0
nkcB9ZxC0zhxTct5xgA2melNfRv+TOyug4V/g9sgM+H0Cpd1OUO9ugoWYXFm/rAR
S3lCa/WNsrq9rniljkYn3YdNcWDRCS9K46KFgyn36u0JNH87ymwJMYg31NcBNDDK
TnypR0nDlkfTTs2UKF+6wNxFh01FVTy7B1Qfz7X5i1208GjaSsRZw/scRCLayeUX
WNNRolYo7aBmM+YEUbVJUtLXWLoSVa5GQbDlBeWUiPdxdDiVmhYlHtsSSJ6qZgfK
0LhJuvwTku6UIDeYB6B8tUe3zwFnJjQZH0/5uCPfcluG6TKg71F2uFS3oFiD/bqe
NvK+ktGebWAodV8Ew71Rhr6P+mQpVF6VyHq2yMBSGlp5airtP2U/VikxpQpanGDS
RAE6OIRfW7MbLvSBRYy/VC33+nj0loUG2CQJSR8uwgJm/gbf60X9D/Vp8DNun7IL
X6DtwOUcamGSDqElWz/X5TokXX93dh6h3CxGzmkScBq7gvqS4Tw6CivplfBo+Hcd
oBl8RllRCRFJQUhL3mTzX0vyB3RC8WaoLzrubGSL20+xWbmrTFTqQ9JYbYKrLHTX
Z/ekyEGm5ptMOvXVe8j75RrYhfkfvha+IN3t1Z413UUoPuZlB923X/azPV3aVbCj
wlfcFa9WoHtZsV88ienCc9JCpaGnFNMlCN1hOvz0G70TSFanzKPVexVnzBCYwPYU
YeFJoEtxzp+/+pTIpcK8FjpujlSCb/Q2ggQhShrVjUUTzKgQw297jiXKLWzvbfXI
zo6Qz9zDPFuFjBgRJ6WJDDEqc7alZc0qe4/yvpyInw3gx0vao2nFEw0DApTwlbXI
RS31Xhfwq9Zogl3jEgkKa55hmFxYgwKfmIQ+VxwDJxbCEA4RwqPJDAeHkr7scUro
0hv52U0guTrcwIHPeMyl0wYdG+a7BhKkmGu0ema5AAhcc3uyxgpP5JA9hXEX10TM
NJY7tlT9L6oro+zJNhaOdBIhnxk/sbthAFQtcf537dcjdh3LOm+JRT882l2YjszX
HHa6GvqIn4MQDfCT4gynTMJX8FO4lbayoP3/3FDDwymkv+FT1aufey+ckeqcxiSa
M9E0jIW3EGcUlVEoaZSpyHGzx/duOjF9o6ylUxp/mDKSBoVVmaeOF3Wud6UMrdwv
w9pSoksZ1ZB3B1lQfE4zcQ4Qd4szBHdJeVH0ARw76YUVKNGEXhcliIItp4ZUnDoE
eunNy2c2swpJfOYS0M82sWdDM5vagrfdVMR3ZkNs+0XUiATNP/sZXAJ/nYOttVSY
43jLHPLCDCtbT9c22EUzZMtHI6fFPWk3BWX7eJB82NJBrGjGyPPdS8toWnv0jMoe
9XZwAQujKFQQe2nvUECJMeqaXaBOpYIdAyviY7fYeDfo5gKnkIT88J3JMF5ZpgyY
Cm0OOjy/CGJLuIYWlViUru1SzmrCyeB4lYx2FiUecsLKNXRfKfF7A7FKZaUDdcKo
/9wg3a8mTxJTofwh1tDCNaw/1zqGC+XNiqprsJCKTFA5Z9eoL0gtkPePODmMan2d
owrGO21CCb3gJuVEpgqTVj1yYdYw2kazqwpDEH8ljiYIAVTvrLahfQaTA/l1M9/N
mZ+X/AS0NhOiC71OgvsPzcO9KzZ+fEldjmUTOmETr/FIFy3OIsjUj4w6t9+rfOXh
+Sp8fNJpRuhfFy356NzPFj9QMufoS0o0F+7rtqGT0GipgL1DrC5mIOa0U8ofYz21
uknpRofo8KA99NF3uzCWR1zODFGbQVtxPRLBsQDZNyARcR2ZSFvghNF/FDUMmWns
9nHMV7LmECKWg7pLcHlX38XkeyCbUmsOFNpfZlFSlH76mGwAyVC5iPOLTxTZIR/i
Mg/6AAIzgc9JxZIyg+6pGzgR/tsNPfOYqXZQf/BdIhb3X8tcpnr/mUj+XWcelI9+
qNE2rFWKVXowKxWpa2g/ZPVd5eztcp6tDrorFC4DjsWUXlteoYmYfWJwhlnf8qNl
ojXK/KmNkh2nIGDQfHATtsOMGLHiEbjmckFswbEzPcwj7w3L05KA4+hzBkCo6ldt
Zrkua6D3t2mQcqEaRpDIyZWtbcq4KsUadfacHDvh2JKp2Ckat5BJYeA1zj8YC8Y2
xz1yHB1w/7qA4d903F87wpUWFJ+7zHKcvhNr7EK6ztvDYkoEAtCRff9tOvZbDrIR
PcnqF9aYSmHJGlO+fyZ9JieVYopRjXSki8LSgy9y72Ownhp7UP/XooqzTseZzgkQ
yqzfgXnlqinX70hEBT5DcdPOLX/G2NG0+eYr5AuVlUSQ+SC5SQw9g8X+4skk432z
SNwYw9KR5vSDnF4Eh7aUg77UXlq6jOK76N50zfAn1n1u8FsMtPcpe68nN4XJPWQw
6juafzS7TovZ+vr3vaa5dU+gCPB/tSDJa3OCltj2HPevM9ULCcsvIWvaAM8CKrix
kTbzt6xIcYnxIqmQE3XVfRGqudT2aclendQ14/9MWAG1tnfZmDh0j0MbyJePgyhU
bILLh6kS9kx96jUYCeYkFVn5YRcHhrb34UgWD9QjUG+R7VkrlfXS72YZAVCENixv
MGASeMPsBlTe++N2F12iJjB24GTVNsegExYIwnMHpD+pTzGCSsQGcVkmjKqO9dgb
Ud5OYrfmFZ5vhWq9cK7Y1bnsreMoKhsLQHPXpLj8MTmOFJTQ+ycQbitV49EPYXqO
/nDBqMzGYTxkYvljcQV057sYVwM+1P0p8U4c8UlFOhDTJ4WkQgRexdnBgnZ2yRAE
ZHrKXH2wxyN/h8e4LUYxQAdBZRdoYTcPyxUnrNqTGkjhG0ouBnXTucYqR86giX3A
3kMulzljgHV+3NeOznCfbFa5wctUM/goImKe95c+o9OChV3f/r3iY/uby2i6pZHf
9DY7hPlIypEYxcQuWFvuERXOCUE8WaE4rZz0aKWypWgUwiWRqCeZDeaHqRYrf4kG
OP0zq0X5F4zAFIIBNGfR1JB7CaJ1donee0N+tqmBShgWnLj4szV46lSHaor483/9
KihzeGY5+mPwyg6nxJIQ1fnb9xCVvyk7jrkhqjbfdDZIlerbpm16F7tiGUaRYOL9
eIQCLSHmbsQU2lyUeeyYacEL3h3MCiWsvKdiw6+PZ90pttDUdK9SPda4bEyfE4J3
R6AinJrjWuNlAdfzaiOq5n7eJSjhqX1ejl6Zk7Xoj2fOApMe3hjY2tvA05JY2MRF
sJ8CtuUS2MoOkPNG/pnuxC7kNA55gMfa+ncvdAi8Tr8Td3Gfn3bm2llCRH+mEauI
UhiyAd6bZpjicFLN+rMKj86UPOhLuE/hHrxoZ0Rztwj9BuSftiUWkrfjBiihZGAl
cpGSXEBsOJC4fEa3I1JVUVxWnhaP0zuIjc7jtRulZ4pD8bOh1XJL3wsA2TWHuU0X
2cf0/PzCmUbLILvNY60D/Cn/f2LDUlYAZWI5r+AzcPy183ev/siJAS+PrmLLYPlp
S9YUS7C8UtDQU5xlyt4RE4dY8Na5/xq2Xa7WH5DS3RbT7+jQSK1Wk5wKFxGilICP
DGdLcSqcA+0UMmrpN9udkUsGmi/zHWiHXu2nySAS9kDMX4mDAMYS8f9ekU01Hj6j
p+nTevlQT+CKnCaDgaO4GxosREyG8JdZ5NDVQSPPsaT2105brSUtdbAHFDR3VdkR
TOwj0kbIiXDYJR6wTYDpE2TBsJZjCMvPF4wzXA4AQMYcuO3p7LuGqKv2/gMOj4+q
kSSnAEOTillbiI9Mvd0u2/vI4dh6qVlsUa8rk4aNDnPSz9uWeEMQDVTs2Bc0SPXN
ZwYUNrWCsSWQ8gEkMVryNbUm69Rw2/zfVh6rZouk9M3g15UzEBmLvXfP39CJp/2z
fafr2DfQiZeQxzZgmdqooYBwHf5m/chuZEoMqyJMQMzebyjM7WijyYon/tghC3Kx
T5BP0QzgoTAXKYLKUIx+KN90aNVKZmbuUb5soSL8PuRUyUQy1wV7Gt+ajexRHxUK
rJfzrpmd1dkHUgII0U8Q42N8PYwDY6/e9Bk5zmk9kH0d2M6zSp7lv5w8KPQvTHey
ROwPhFTo1fKmWvUhLZulh5TSedRzCTg6KSrrTw81tYQd1oYoQKkiniaofiCYKM/f
vaJ0NFPcRYvT7IewjmXFJPxIrHZ9P6Hdvl7wg5SumkODanVVtY+81wdRmE39rm+A
aZbwd0mLSd68Xw6DnyRWmGj7rrrYl24Z9HYOaJEM3mRZzXUf7wqxcXHe8YOTQwOo
OdXIO9IFlJwpo+9bNK+LGK/1jllinex4Q7PR/BGOOpZtJBN9pH0XfZ8oodcdhaNr
wJ252GvGFu+G0iAAB4nCjymEXu2Tc9JcyE76g7hgUQYRfj30KPyTUR8RkQabQ9Wh
0cMsBMAGoi00t39o4kHbyiEYScKIbD99M1RXFjXGITcR64fo85LMpMhlfhjeO5R6
jQJT3TS8prGQnRpJZVleNb0NQdxemOzJ1fI72I/lbSYNl0Q7dGCjN2zhrOgbKNit
HCz0U5PhhVn4WBxuS5KOxTplShJYMM3yl0eInDbCfpuGsQmx8B6elPP/yNIWdiaU
mSw9BBmU0jPITRjdQNdm7Op9wzSNZmU3CczN49rtMx4ce4wUSP/lIY8OqxfRIzDt
COmQm5SC+0LBKg/7X+FM7p/jakZsgPEB5GBtPxQaWwERcyLO07ljXFEMQZ93GNlt
/IxYa6nfSEAiNz9OlT5WbL1RziT3hkS/2Y0LheAs4cn6N9LTb6Btt9e8+i7ZdgKo
8+y1QDVfwtLgKhNR1+wgrdZkuqTr2LHXfxSQzme8CRoxVEngHqOaw/4EdfLf6XBm
XyrpsU2ODGpDCYf+GIwEDcgzpKPtXZT+FL5MnQ2t7NtmJ28CTyLtbWxdyS/AHH2l
AychOQb6RHpkWti6ClsJJKGQzH28mIUJNSQWxmgk+gD8RX2cfu4Ct5BkAj4r0d6R
9iIg6DfHrNLu6eZ0rOERXUJ+TIR2Xv/gvtrIlOg3qZ3GRH1y+lmunXBGBxhS0Vgv
EaPWvawKlsN2hbGorHWbP2EtZh+BbQzIlbZoQ3ZctzCwgrls8TPFiRZjSeGJZoZ1
0W6SKOpXkZrUV7vsu2gYbtR99AQNwidEMltQRoM26MjPfX5sf/EB0yKS2A3uQ2d6
2O7t5pa3FZTyPtLuGI83uney0unRJ1dVakKmwTcEk+DsCmJCGmsbAoCfNG5xX+0a
eLdRaU0aF4MFg0Q6hmFvcAa8ffSu/k9+HCig7m5mrEbMkJazC/Ue19/D+26OBmy1
EinpGtXmjSFM1f4XzMXFHRQH6p+CAyEl9WV40+FTBnmuq/g15mSnIJG2ll3YgSM9
4tunU1SBLXrWnEBA8sjTa+1iAESvKwQrlxYbROP1m5I5H2sEmSs2zZf0f4Do2tvN
NftqV0CiVLvq1dWfMHvQkiRRgYD+Ol3ov3NIFDvhTLIJwdonZEPba75TfzDXatcU
mt38cG2Hg3B5gWz1XPjkvt58mrrkYNw/KlNTHWF0Ti8k2BrXQsLG4GxwrT2xUnrN
eBI5aKb9TbvlNRAM9awH7I94Xsrz4jorHbuzlQW2Tdr06BFRPCauGGX5iNpSkfJN
Xsi9JbbjYE7T7o84Ngya9Zv9XDgin305HqjEBBEf9ao2QyuA2FNScffWxX3XqYhp
6a/9Hf+QLb6IvB3BFG5Ugh1aoPgNMr/p/apKu5ZHS5VDG7Sz6a59wj7yeU4mirFa
oq/U4RjLplpk9cMIZ5/V8W6mEbOsvV5n+g+Qy0Rka05gCpsBp+ncTcV/Y1UtBKiv
2nnw6M4oFzLxnxBEzBAmsvlF87gXbw9aMZYwX6ImVL6S30ODr2A15ckOZir02p6f
R/2m6nqvMcHFPo5FFVIe2RXZCGXkCVPA7de6RuFlSsA4LHAYw1lcqGtkIE9nLuGn
aa8HqHgJR4SQ9xtL1M6QIC9oCqYic8ezv1lin1UvS/3A9slnRyGTaJtPhq+WrNL8
BBt8G7yhfdF2x2gO4hhGPddwnAF39D8u28S7h2S14YBfiU2ZcLtcS+ywjodDS0xx
iytOcW+qV7QVohdwnxukqUth1xLNbOyMoiM9VmLI/D/z8dSoaVNHPi3BISFVPBy1
vOmO+K6NqeWudBMAvMbJA9iAyDkc9TShKQ2wZQ8Y4s4LFo9gv4BtTW5mI9XfGEBb
jQKksmH9LvYKMloe0OfYLJq+oIfL3I9XH9X5XGskdcjnynFRBw+5aCKV7gs0FD6u
mnaRIVRUtwpzIC+2cPoomrh31E04So+q1axX5r2BoGPMIWzIUmalvv39RjOAy4fl
USMQFQ4osQhdb5tDLp70DxUuIAdfsEhWcnWU3sedZFQqcLUTw4lK9yGMCzQA7GVj
6+7CXZceT0uJfzTl1HAaM/HpVwVS31Umz6PiM6TNxDswl6ZRuUrBf5jFevSSrBzq
yBycOhFc1f+4gmOw+3vU1rYRy05ooDQk0dytGmYot/PHe/vlfVeE3WFKWt9FUeLW
TkdBEbknUNfz/iu/H1eBO2bhY8/NhE1Q1EkUD51oRWNyNxdf1vEi/V5YxWqTJweV
tlUsv1Of9sgrB0kdAZ0+A1CNS81nm5j4Cp/sIbYACR9/hfdSaeI/nxBIQ2flWwYc
cl8q15Rq3usjyVjTG/sJzXiFwwJ/yXkHZA7ftDuDvXD6IdFSfhvSAOonA5+83GUL
rdUgdACWzOI26UVYJKR0K3pFcNZBvOECuDSqo35jaDJ1oe+JmXNfqdHKkgwHvzES
U/AJlCKiY4jKRwXgBQnXse7ca6ksb94YLnFP+0kxp7tWMAevKYZ0CGXheBdviW5H
OvEYv6XD5CNSV2ekVVo2+LV1Y5mCLJwOabWjX9Ev8ileXS0uog3syWp4VfAV5po+
N6VVqWOzK8TejTqKHTs82jHsjA7qIcJ6rZH9dmeCEeDB3ZMSFEBqV33LGSR1FcRB
8/DzlS4dHzWtwS08O1SzDMFW8kneGiF7552vhPDqbu+zRDX1HQ7uvP1O24HVNWj0
8KXV2T5sDxKTavdGi3DhcOtSxv+hUKj6SF69M49uMsrgevaL/zm8lN71VCG48Yqr
koOMHdXbeNY37df6h+Cwfnk90n77LLhql1nVQLAbvM2oUI/fLmxpTXgz5uZcA9b9
Rzd4tIScL512MD89ctiYeBkJTMzDfQwTNSddVh+ldIaEiZ1E8tAWA2IuWqr/xAsh
se0kDBM3SJyTQj5eieDUVwDqKAlR1iesqdVHUCTZWf5ZbVYaeHY4sid+qS3ya6pe
8ID15gNY5HbouZiEdjoOMY56tgW/eQ3f4fp7dz5fOivbMkcz4eCSZEDm+XYxZZ6E
xe5r++HuZa9gDY1tTNpM14qmO0yKCnpuo9VYUJgWQwvlilpZB2rRRLXCy5uAsaFZ
Fj7MClQhm5VATnFmJVgyxQXWqtiwC1/a9eTc5zNfClnIx0V3k2OMGgVDDKXPWmRw
NHCYjN+EBzxuoZnl1AP5YHfYQhD7bKSZbLATCf6SP23EFXnaEN+xKdNldtf6IP/1
QT2tFgIMq7PI1izqmGr1h9AfW4IfAVbzVifHJ5zfK4WWEppyRxcuz8701WeTNY1Q
UhDlux7KbHdj3rIRfshTsIw2OptI53jQ6I03I412E0PdZvuW+ZjWqjXrBSXPc1kB
FZQa6sqkJBGOhwmdaMDj0v9xnZuMaQsPPNvJG2iyNfUBlioqAZVSq3T/Cbmy5cpn
d2qNF51RcohUpoe9zI9yDl5q5UC/5leNzh5Isls7rjiMkxuBOhYjccxZ4J2tJ6UK
qc5yy+qzG3sp3EPI+a65fM8Gv4pH8AIlo5gdAwdXrZ2YYHMPzU89J46E7No/nEHK
3Yb9fYZ44sSI0TUlMf+xtCp3XDDM11GleSVvP1rTIZT8wcYDHvxY/XR8Xt+CoMJj
0lpDw1akWH55EeH/4kUOIMT/Bg4+elWWI5VqeGouPiF0Co5/mNvrLajOchQdHbG+
aJF7VkOYmHVjaUL08JKbvxQANZ3ruJfm3+LZcHRxi5HTF+zcD/VXRtvcqovGvaoM
Dpc7IJGVsqklheEkpAPtHCJrYmUt3bBtPZ6gNeMYTSPT7awofxVLeI1mTyeXeqVk
GCPGw3kyRykF5Ooiu8NQOe6oKliDJtuh5sT5kDbNRqPiaHN6gfcz/B1qFIaSsvBo
ww0LbavprTh/XtPipVkK1GnLDGqTVCHQiCJJzIM74vB0BegsIt/SL++GsAxdkOcc
xqQHLwKU3whknV0dPYo7GCuhsgo0+ReGNrFw3TsrGvvG/ndZDoq8pv+eqOeuSiSm
mZtIvlJH2rsUD7keM9n7HHRulnjJRAyR2yqvlRwu0XQrrddyzNE+uoexqH2Ekck1
33F+VwYZ0ETKMseIqdVEctlRkpi9CB3q4D3rq5QCMXWCG6ujPwNNKb1lVDAyREOr
KXC4p69KNe9e5LP+iuSO9ekfg8N8uTqJIWPL1NGhjYlz+FYZACSGrr2X0ZGE9oCs
WRDfJx8SQzET6uiA0JLu39+DkazhimwwFPzUVsf2CCway2+y6NG4YJjbQZ2MGFsf
/sw23OEneUQ40Tft85qB+MyQsp5Pif3n00/wBfGpsMLmqSmccvfPePUFEHbq25Jx
h0bVLEbUfzThQJJMnqLmrvF5xvrSS+0I+yuHLz0wbIK9Vh3nRCwffzPwNDyxGSu6
gVp1TK7yCxdKCVZntAbJYQiGdYUh6lPP5tvF7LT7FVuDIRWiO3lJB4wpA4ksN2nt
bYGzVgp5LrtkdNzl669JV3zC7gSA9NJZdSIRJmP9xOOWCtvgbx6JTKKQ/qFLhGK/
nTPZyMUm5XuanftLsVL+q8+xdsa0g8ZJicGMS3t376teS85prZrZ0e1Ja8sM467I
SvkPWBIXbWcpXhb3JsNCCGbmOrlkhoLHmJFWTHMHm2iycgSfDFj4ig7FnHIdmQOf
MMqrVEd7gzh5oCTjM/UIyi4GIcnXRUTP/yqyrtpEFamwb4rAwnJ+ebPPS4MSSFcm
wkSfER7XMtAoqRxqU4AB93dtrd+CxCM4/1F0N4TidiLRjNZz/5PFgXr05jrrt1FJ
w3dfFt/yxx+fjK+AiC1UkvnYMJNnvQAYB2//FdFhNb8ABipUEbexxZ0W0ExyK5y6
OcqUh+HN3j1OAL5Ebrh6qOsTw0foOAm1Z7nBO+hOXKh5dP6xMo0fp7GuU7ec11Vc
yogRDec4FuhrEqoCFFBOAY1dBrwEkDOK3R3HsTdDwvotGyZxF0whinANvYdo5sx/
jHhaqzjjaTJE1hKCTLLQ1DM7GnRBx85zZZPNdE13H/X1uQ0qwr7RT4mkubUvFyQ7
IN1IBu4W1srT9nzjc11CRLhf//pRFmPat38uruy7MfRqM3I+f3/604a5M9fAxBci
wJidYbjBLeHUZzaUoE2cfYm6aWKfIR4UNWaRBIejjUj2e5brcZ1Pu74smaFgYV24
GedtrHivJLIRsLBZdhaRTwF1+mYoyN2katELMHnSwUB8VsX/CPPUoxIgI842H+pX
h+A5EveeF3NYvKfeenNqpGD6M7UfjpMJObFHcmLfGrj9WwKYbwzJQJ3MFvjzXwSP
ObHfuERqG1I+tVkilWwA3tHEQeAcQ+yyNvZf1jta8+KOIWO0XROBkZ7xST1WpgFJ
+tZLvi6EjyaDn7M4isBgAemykfDmyTJxMuvR0R83RFvQTcuuB038tL2kf1GWzX2R
Vhpxoqf2FSKzbmHuOqqrwiNRT+jdDe+fthGTR3JcRMzvWzC8ehF12FA5+dGf4vZI
jHWMsNJkpcnBzRzOjqQE7CwV0bMsg47Cz8WV/rt+xT8ldeDSd+oyfUeDKhRTfc7d
oSdjU/FwtgnuCDYaou/FmR9DPjo1dU2KcSgIsSoebdWCfYJgli/2yztZ7Gl0bJf8
Yi2rgxZQBp0utN2AWEksb9FHIwdR89NroNZExtNoP9yHK0zF5Gw9BEf9grTUaKuR
AKX4x7ukE7lrN1lwlEZmEP1V2U6gAOm8VWGqtWli5i2gMozEhS7Ow00RBNLm9V+1
nTG1iITcW7D6Rnhpythu/KVO90qYG10FwBYGvgID3cbDNmh8J0m92ptIwY8abWg9
PlB05iUaGBMOmltCe67xrp8stUoJWaPPJyLQ7nXl37eO6B75XZuNhGZ5j9W9Ak5a
G4AYBGhfl9d1NwsgvDxWYIEkdILobjdU2+6EcugspB5f8IASyel3l7+FXWIFckFv
6g7thuRODa0wtJhqMgax648ePk4MpAsdra2zQri2sFZLoKYR7O7T6BOQ59bXaeFC
h9vWQZtVXWLKtNuKu+z3FtX9KqUhIlrYNybCLjHNde5QpFQ1EFWe8VyClX5b1FXo
itpdKerlGcK+4VMtB1Zws0cxQY7HElVfTPudw00xQqNYMJ4VPFKlMjU3KXKYwrCz
9i9HqhRc6YYYQxqko05NzlYjP6IoLS44gE43UhDsAOqwhQO3eQJjyPIJ0JZdYqcl
MuT7VzwzXtOQApt/pceLVrnq0Z9H3RbdLm4Jj12cLonC9kAoc4JrRVG2ktO8VN8l
mxRIlupkkWpvQPE+nZImRbjgG1CV6+hF/ivJO2MkqDppXKAN464jSicLgwWuCaOs
qMc0t+0iprwFa8Zt9i+XAlFwIedjw3Kn4ovz6nj30Q5kNhs34rjcfHcH0ocwQNTv
HRsC5r39RroBmvqDDkOAFAxJizbEz16NtItw22GjF/kokqsX5dV5KUZhJgiOJo+7
MfvXysAu/KJjasi9eCi1ZY4Xk/52EsdP9N+V64g1UO7oLbKzV75Ykz5MpU/WIbMg
kMeXBIpzaoQGnDJx89Ygi+4spmQSk2CWOAXj4jIW9UckhH1kVWbsDRI9Sn81PDSj
lIMbFi0c7A6iinuaGZbh90MyYJZgsyHpU0rnZ/tzEnNcCliHvH+ECD94hyo5O/b7
Mg0BB1EplTjf+KEaW9Nf50dj2j8z7jsEXxru7IlSLQrln/MwUy3ICZkYGoUcr144
DWnXsG9GELAfXHj8/+3k1558Z/gs4xGVAGRgudwKn/J9vx+DJ/BsR2CY8/F8anu6
8s3K5Y3VOgHo+gQDrvIYSyxBK0M0zXK74F2mAm10rY5g8Ee9TRRvWZqCziS6wYW2
ZSFycYGhHNv/z/bU8GLTA8Fh4OcHnZhJ5MpxHhN81vnOTb2uu//5chjilctvA0Uc
3ESDfxqKY1IPIIvWJ6bT1eC4HUj59IwnRnP/a3z0i0TIAVWW4l7AIGNNWYbafLX9
wCGps5o7BDm7xhn4rjF+A8lLOUwEz1DS/LNxbl82xU6+QFb+aCd+HD/NhmRJVyRx
ZlXgM8rrZBsuwbZn6LVLP4j88XWY9wWGwyY+GU/sdoKaJ2lL1wQ5WFbkSD7gjHll
6ERlewOEOWzIJ7+m3P+NC9vcjQzAM/3jbG2RTYkXJP+0DcjA4SACcGzcXRao0IFB
oSKhVezgGPZz1JA5kRo8nLAeazfcS03SD/gdFoNKbof73JFAvIgWvPygqbjBM8sQ
/OtS9iKv02nypqY12K+6SXR8BqlElXNNxlnWKOf4M3/iIU5dkhEUTEDO+l7z4pse
Thf0ei2nNrmMj/TyE2qeED42x0j55dBY+6yctkYJ3DYg60FZTBvnyMikEb2OhYqd
vcO7s0n1JX4hTpXlycMddF5J92xZpKKBMLpEXG1oWXkiFWUNEXfqgSPYE7TGCYMd
A2F8Ag76EMkes/FKSloZ2/c0AkgHfODMUGyga75+uTNxphlaD9Htr2gVq0kWBR6A
173j/p7on3xbyKMlnfXV07dow6GZJx6jm+zn898UZS9EjDxAuM/NgqjUIlYTxF95
KNqD9JBfVP/lK2qHZZB16aGtGTCaFapUjGaORtK+4RcAI0o4+jn3JIyfKcbXLZcF
zESXgG+Qlr6DX9g+gk7plUkPAisyZRlfE3oKFBGz+y1guDMLJh950R2AFgXftWrw
1wuPVLHvQf+G8cyhR+kijkgYpfZVgdYJDPCQFYyB+my5q2m5Mh5phBLMB/FFZopd
IdVdASyPw60lNLPVUSypG08Mc1rURi7K5jW5BNbSVHwKNx5e3s8urBZHD/TCL+k3
DfKVmsz/WtpYrZ4naRlUU7xh0ZFee3lHg4K7opoRcNrs+E5UBr7sFUEGE8n5sVQ9
Sh85waAXaZvXIrKypPS5ihPtCu6eNVpeuksVOirGOik8Ka3+SRv+WLa2p/MP1qpi
ZrZupaLJv/9f4FJmXRQHXaObQoMZtVbBvXA85T74O16cakjUC2oPdrLVdXDx01nB
fn0X/Qzs0Awh9Q9W56ou8qUsuojWklTkAaEnNf49Ro0s8wfdMenmIhCFXZMzRYcg
xfgPuYOcOPnqw94hxO2bHeWTd+1eM30YozkCOFlb8F6r9obansPn+rWCgY37jCA+
eHMJXWUxEg+lcMOoFsgVwLTy3itrVpHT8sBm2etUZ47r5G9/vAMyL1vQsUoiAcuu
v+bWlCQJUDjTg6PfcTMLoFJYbvhFKTVMCQ9R6oK9hYZBKGcu+1d08hjYTD06BnEQ
22PjdItOWLmGo5ttNxlnmM3PHN4gkHE+Z6WH2kYALSACd3LAjAgHq3lQ1D9W3OTN
INDQp6wzTJgg/zUAV2RTo9wKJtO11h5hdmOIZdAspUst7nZXXIeSn2yUJGhnf0nA
EYwmohScj0aIM2Bu4cioRVfuQ9mEvHOVWnaGBy2XsJ9AXhOh6MD5yE4UzCr6/Rui
6KYbuLiI2yquVenPqXGXPUl9Qj71iyQbkBi3X1KrkCNURD9XSkzwE3Cjyjb4Txzb
wi0H3ddyTij+n6i2iZ/yiHDgpOOwJR6GIehmbzeCP2XafAjkT6LfaiRegZH0vKDM
3bWw1B0OyBBq1nXIQklmnfHXaZ7FWy8qu6uhDWbrqP8ThriB8boV5/5MSDwgzWk0
Zp2ILIDQ4Sp9sr1zB379wRDuNkeCv1PaT+ex3NYxElAySBZzEE/6ZU/T+aecsgo+
Qa+LDI6zt96pW9TPlAoTI6r3alX5wLRU0xxsIEicc6UsOSNX8DCNA7PqezI3MHbJ
IhPq4PXjfwUu4OhAiZHy84jJka7HlvmEk56+jay7wt6pj1SEnLxEU+mWFFH8DhMT
SYr+Z0STB6+mpGSrk5r73ShAr7sn55PLbiF4frHWkzvoQte8iKI9RvgxS6R6VcoV
KcV412JIjBDomGHv1VoWg1G42p7sQburyHekWg0CBnoWlbMMgC6T8hxVGbgClRHH
j7TGqikLPipYmFirkiqnWtncp3ITW0XA5hZwFfi3Fe1TAkr1gw3Qqg4p7bJas7ae
Q67nobnYf6ogOC28HfaSvOa4aZr8mS9zxiCwpr/xtgnT/QdRx/Up4mnUZj0RNG9N
BcyNW+apv4E9kQvUZJQF6pACcvB704wpl5TervMkc5uFxPhIMHMmBE5bZ9H+HurI
X3GlK880zNuczE7IMqoWSGOQXWN6pIsaWdNpohM9qj0OIm/FeouHzuxhN71mzAoH
89jEuoGx11eYd9MQylm1b+OwcyDXGJbTSGderc3LNTrzxLetQxK+DB194/yZc2yk
e879mCEfj2nw2zO6rqtRNII2QpcxTXbuXb5/4suMev2U/Gbum/BAfgLA1ZZk6U0H
trOVrfICgNEPa9BD8FXqESWyRkSij5nDJbGo+txKa4tji5t/PPluGTRXdlaQCG+F
Z6bSBUf5TcAwFHpAYp5sbrE8wONVdE9jUOrVhqy0ULIZYh6QO/Dk6HsaVUk+/cCn
+Zz6rW65Nt3V0pWmORKMdAbUXfM8kHBaY/rh/0AQmBWM0Y+2PFNrOmMN5PfMwdgE
fan/iTM6hzzSmMIOO3wlVX1WwYfeQ8mFVQd6/aYVo8R3nY37Qp0V86MbzGQ6nptE
uW03bqvmxlVvbCZ3dS6RbE9zWkIKw8YCWCA4T2B4BJdhFY0+U2xOB3VVnGjQ7D4a
QnEnns8vurwFHneqNumM0w/3SzMIbAW1Pd1QvKbNh3YCuUUDG1XuzI/gevyFQywV
I4aa1eYZhhj2F4sG3DDcpOqaNn35y2vIijXdy0nG6ZXTConiTxlGRJjP0Yp96XbW
PKIeLRk6KGtaf+DCSS+2cIijQAT9o4pFUHUABl23sPpwwzYTQxHt3V2qpr3hDrJp
Q8vTqfwNhbsapf9sMs4sGNed1KxBOLa5A05sfD8JfG/dhsA3XmPrxgiNf2h5Vqgw
zxsJ35YDakPhmxpIGy3Ll+/CvGULFuXUeeL11pRIZIUCSTCL20ujgVn3M9vTZt3Y
2uL2UaZGK9pAWluSJKwX9cq7KGxpaNskmN1dmIV5OyIOE2JkcVilHEn72uCOVj2F
2kjb68G8UzHJ/DrETC7OSfdY0AlHpwMOGHBZWh8PKoSfgx2W/rfGLt05nCbZWC7b
H9yyyJ6jlAYu5/qrxj6+eS02oxEclhSCvVAjgyehdaxYaRXyJNZSy1tzzmXsV0Bb
7bxC3sFjCw7sa6gCtIU1ySxur4dPEG4bI0kDH6ZzzHdEspVJYphnNJUJhpIfJpwz
GEt3Sdao8Xc3Y3AgfuE6txCjqC+kq9wC2FqzKqGwUrAlaTETUPaxsKKIwBTPc5/p
U3EYZcW8aHTPAE4NEC79r7xSBPIGfxN0nmSZXZ5KIopke+W+WMGtTEA2vW6vv4Xw
Y+kGYVvXoeTVFAEDhpgU2ndNgywP3wMEdcy8it64tZREc+sTXrgCcvR7Rf4YU8nr
6HMagYyJmJLQ6rRQrWTqE7LPT3Afl6W89xJrGS3x1imJYFbMn0su5Symv7cJYTKm
dyKILvMG2p110a34gBtTVBnYUEthPyu6x4hz3sRqUelO8dEiKXujyScAFg9LytFw
rhbtbnJWeKURkw7tF+aGcEojISE8/MI0PjzmXGCFoViQcthW6y8N7E1AJ/hOhKtP
sJFLCgcpGZ4yyVnKY/Z7RyIGCngj3hJkbuw6zJG4L2bOz1BWBj3Em/uh5bUwZUnZ
9K7Q+TEMX76MZRLu0svICf4F4EKxauYfFWNCd1YxeiH2WbGVSl+59DDgZZ373D1R
k0iCIMvsCMJX58DFDgQ7+zIpM91l75pPS3s7XJe5BfTMA/81XkUAl/FmGAjfCS+d
+e6gj3+bABHsoBMkj5UnlllOtaBFHSv3fXXdx73HVjV+ZbJ9qbsAssLyEOdnqMOZ
/6nvficbpWk8sunSoiUe7H7ljDS454sEEe9vfccKMS0WwcujcjmGBsYAmJGAbDk8
MgV5jdICj7dkrW+E6ve+NnrmzumgGx1ZP4EjWaGLypjW1ET73tDbVp8UkDLQC3/U
veArA9B2gs0e9o0je6xkU6k+OpAHwXtva6I5QbHlZh4b2KIUhi8DeO93n8Gp5xMz
NA3+YTPspc4G29TLInzuvF0MSgD7hG404n1mqa62OPQU5uayOYGAA6eDQEnkUZ5K
TJZ/kewueQLtTxTZy5k7HxVXagqMgci3IOMRAlg63Kze0AYTQxVC2JWvi6nU6p3c
z75pbvjoKaukGFvskawIUlJYbnW7zUyvjcRsWsT+PvxrE2eVH3i6ho0/b3ZjE5En
N/B+/KvWftW+gX/Hsb/kd1rAmVE5Yny85LXpJ7jbqpmLwuMyOAZn9p8skSNZ1DTn
XEqj7jF2oE4gkMhFiZTREwM8dWPCc0KYeMlTIz8wbeVaIFEQbCBn+2fPsV6qMwP+
Ee3DhOu9Ei4pYP1DodFJFnAwheVIsYz1pB2ZRlXBghDW2ytmEZzLEYCL8EBmIviu
beNf0jdsj8JegN5xZaJeAQnu0I/K4fsfet9Z7Vv78I+19YeyK5dXp7Hk8RawRyg7
vYatDWRh3Re80yKYLLvwWIMbUU7yKztWUQIrfKGD6ceA7wAjZY50oekkv6ghKSU1
IDx5JLaSQrkaKfylnKsoB5cwNusaZK0rLfjGKz+XxKTZJAXic4IDr6vbODONxZCA
XQGWjf9yW2yy+Y12sdVih+hpKw3qa64OGdchVXQHK4vPrTjKM5bat5Oknuitf9OF
kuPHB4/naDMtYMIk1J3wuFyvFHz1VcRGZdqP7xyD2sElPJVmx6AfalfwALQxqQbr
/GtxtEesGLkE+WiqKgm1eyjELcd8CwN7RiVvNIHwlT9li/VjFReTzK1MQ/AAqBec
2aWjWrICn2j2DMFdKhIIcz2dyCiMcXeP08sH7a9vIK3ZRxNnsePrdvSIUUR0I4Ro
CL0gZxOauWIn3gOk9oKkprrQxWmtLSAom8JYStXwZxzzSvhkbnC4NlKzwVQftKee
I48Jv3fRP4wi6k+Eh94dbyE0WZI43wg9Q+7CS5x6Ca8CaqBEtjuwdaBEiKE8bZjw
0l9pfsbcgkQ/6EQwTLAYgzeK0jK0Gi7CfgE/vypGDF4ImCRVgZjt4AEOu6ooBK4h
OhEaOqF+Pu9wyRftV9pjojD/z/kAzEROsJNB9aRrOgCDuVcbxhJ7XAFqLz4hZbr6
LHEthJStOdmmmxkeIGugG70UDyN+W9bBM4pz68qXIGxYyU4DeKFUIJe+bKdQATZk
TaNJIM71Mr1j2IiTRE8ogzX19qodoUQL0I2TRAxEuI20oNlV5gnodOUTv9RBPt/d
jY+/NuuY7WVnHeW7ZXiZlpHtMYzPgAo7kwSfk9M8TKrzJwgPGxBT9aTzrEvlSc4p
phR/UCuqNHtbaiOn+BajVC22AFhV5L0pyVyV2mPd3qdNS0t9SUr7T/1L0CqDd7j9
72cVfrNS+UsdIyAhh8NtkKb2OgBcF5f5gjMPzT1TzKRAZ0iPaSqruxsmhCVmYP0n
SCQCaY5WTHO6352gZsDCAT7mmcNTjHGUw9WzujNpb+zcBIQ8ksllrOZW+JehRaoe
rYdVxRd0Och7p1oiAF0OXSMHRJNYc2Mu4ZItJWq0DsY0VdDd5uJykzZ/QKW+tRif
RegUASBUhgUbAFPxWbR2Nj59weMqkF1vwmIEbmMnerKb2f/liFns4XUCX2UV5Hti
8KUnHNDQx0R1o3aGaKddx4x/7TQnHncOhTocH9Yni8X0j7YuwbkHRNH5ymkczOsC
MuTpnlGX8XZ8IlQasGN+3C7Zm7fCxvtkCa7MaXCGp1KQktkvXU7o3dSLDrceoX0l
TY7WK2DVr8NFqu/vlQ6jG8eRMshYesDRthQ7M90Kiuj+/AP+EwDxcug8yWi2VA49
wSQD+YMxXg4BQbsyGjCUVxlhiXWkHdQRtiIKkh2nppO2KcJJyRqu1kdZ8oXHW0cs
iN+LMDhfFprfmp05tO2uMD1acxZkAt4nQtePCZKCH3U3XEzQ4aj9gw5IErvsJhFN
YTnL5TatLACeMiNhzWP/FBx0Syt55hBetyVB3Jnyf/BMVUh+KR8qLgVDxx4kpgHh
Hpfz+X5hVNM771oq2DTVQyNG1POs2+3UYA2BEn7Z96cle6Qn15ZAgFAeWS4tLj/E
TFg55dTGaS2z9zk2XOdMyo0+SUlKGI47Yn0v9TrCXYM/+2h8cx8G1psQN8AgvOHW
+V169mrXPPPEQMZjm6mi9IPNvrITKincZZIDOZcDGbs0GxjsEAOKK/1c95DK6wtQ
+h1w4FbTse22FWzu8RErDG4GD1PcnTkrRn+XYG7f16we1YArC0dAFNQOU1RwO1n4
h/SaaRZeTNNXpmlbovCVe3VaTSFoKoFAa4mhdvSSQZ7PYUKE/qHLZkgHMQMClH0x
jQWMEFx6eOImJ3l8RxhH74XlZbwMrLxQshZRR2MsV0/pNJW/zv5ZYZdRLo5uM4pD
IP7ZgSZ52dQVQnLCmmO1RVAByc0LMWdtRg5K6QQwQ9zheLQ9Ch3sl8Sr0Weifi/i
H9LfbYq/QPZ4th6uGA1p9+8i5Iy6eNF0U3AkNglxWd912INszIcDYOGZ8jd7Xbic
0AHqso1f43o7G9rJVb0N2Dx811vFptc5zzoT/8NPTd/bJSymSwkr6IRPq9JVOJPz
xTuV8TKCp5aaHpcJvl7BfdgQEGIZgy9tQs4i1dBGWSPFoXU7AhqgeNKspJBkRP8g
92mkI0Nkjnul4/49WZ3jqVOg3LFTcHKnwzSY+NnCiWlmKpX4CD/GOOlBJxUXKl+r
0zohXo7CEclUJ41UDJoD/NZyGMp+Rv5A3DF2mRqophpKp94DP/javfcDFwCtOm8w
M7zeIppEBrd5nbyWJaipkn1Mfe5/Kv32q0Wadim0WXeaYrr7SCKKzOKsgqu4GpMp
sa8/NgMagpuKfJArTdbcd6uiYivOXxyT/bndY45gxRnxfDsDC1g4DwKRziicC0Kl
mW83wrpC5hNq4Jc0AuiQRHomJD6ebyT8aXX2CURrH5u1Qn6lJ64lXYv/56XeCHfM
wXsvMAYkt2MO/tKzhhq0ca7mHphbP7DqUlElboQvG+MdVDk6DowWAHG19muQ0Dod
Ej1JB4cMmafzhCasZKQw0LjAyE2m+eDYHHdkCXbMOKmFcqIyEguAwB4hXPny8+JS
qA9dtatxDIK2Ys7VFDOd8R1BapaaSB4bNIum4LyBko+F2ABk/O6lsHKKpFp4BzTe
RoNQOrlCCGUga5GJcOHUBZnwJaJKhX/GRKwpIOKoD08UNTvSXFGQEd/Qbo8iBKP0
Ez14GoeeiiscyI2rlFCmxUR/iiVsy0Xg5JVHkawfbb5bqBqzKsre7+i/Jjj+/T4s
N/zlJMRAVxs5+DJJorOJ/l0hFHhpyXjiN1llahDq7huAeOxlmjibnNpPnZdyqR4r
SUox69tQm5H8fi40lk/bQIlzmLBILBtQydMUST6D+Qb9HFBGqi5c8MxPPnK2hrgi
uCYA2GSYWZFe+7PeB3HQhI3swu3Cd4ITQBaWaSTt3fcmfa/mh1RM0AodPHlJaHZv
r2dvK/lxSoRnCT8toGQLvms0jGmYcEF19Y6h4PO10UBMWK83BwP+plBhTyJB4ou+
pGS4NmSkUSzPwFr1M5SbPwAZHOEJVMEMjBzOB/5egk9zZpdbUjN0EbWe0CvuqaQ7
6EwQYkFAjO7qqs6Si9OuBbmMfg8bOZ1qOXO8nGl5gxZq4sRhJYq3kGvu/P1oSTyp
5pOGhmM7uny9k4taUKLOCiOep78A7R52Q1z1lNOWZhmMaDF1oQLQsrXLzyj1dvSA
5fW3obry+g+cjXduT40AmbKz8F0OIIEzSx9Nb2tcg3Y48jtID6vznDFg2A02fkAE
OAUprz6y3jRMs7AJHmpYCfsJQVlDUd2pg/QafKHny07P8JfsrIYd8H76e2yTjG6l
EYZKDFEWNLqJEkgCd/SYzaa/s/g4PMpHYqN+6AQKARqVYmYLOzg6EPjwsotBPTX7
9fuCpQCkmUl78VIzeCBqBH3WnodM3piCAhW0ep75HCjxKLl0j+QXa+fdKFXsM8U0
zTeGmtdEvCVEOjZKntX8+HqNWwexOWqWRXgPKnNiFDLN6W1EQO3PQtI+teYpMbEA
kl1vRfzh/1IeR+mL+BDGDFLjNwtVQq/cfzYc+NDXRs/TlUMIcRdwv6+3KkdMSRSl
Sn3jeqz3GxDXmHiybcaQVwoXTedhmCWVMg0u/VgWDTg7VG0tI/6juXdcL8WDutHj
i5CYa1ES8NJEbppdWklAiyYOmiuPxTn77bdqxuCHLfRlO3yQ9HQtAM7FinjPqHQm
JPGbPylpH+UrgvVdo02r80VkxSr+o9NhsPSNBCv5MWSZJPhEYjKvQRNRhWK36Ll2
HPmKC1xzKGxDaH80Xnjxhw6atFG+bQxrnbskQT9dGGXqHngoJ5L0YrpH6Wm2CUPU
Gmhpb3oLKbdweKX1KTb3N/ck5qObi5Q1IJyTR8N2goMOovt3/HpxssOSdO4huIcc
xHzCis/bzgr5M1V3nSfLTpcWJVtjvZ2rC/ZFuELcjAEyQKcOVafMF9AEI6jtoNA8
TZPy3xnBq06OK1q6WdDymVRGSqZk+CkgCsZjXecMeb7IHLNhRjEfvGUaWV+hvTvC
qvdf95mUiDroLVk7KJzJ6UxdG8BB7UuxHd7zMYYRXr6P8CLSS9C8tS95EcB4q85w
RJklTveiiyRyj8dCUgvfcfvkxRlwHkBotjzQ1N/mOaFjpmljXoTD5MrChlRnYWDX
OuMYMxvfxkDoghKPMmpZWom41vU/DTu0+gnihYKh+2FqSQzdyvS7s4SUT8lxUDdu
1Bee0jycPL4FOBg3x63tOafiyE3ZxtWbDf4kDBGmyV2atjbgjRxeZktZInZMTZPg
IEoBNDv6mJaOfl8Mo04bXKNqSKGdLZ8USkAPul2gPJMwkyNas+0y+o2K4C8lIUQT
LH4MKoEjUZIVohiyy5x9E3bvYpYXW4OxHAeEtC9Vcv5KVvvjkBbBogSYsXNAHdL4
avcIP4HkpTWt9uG03zaC7bHlTlc6jjE5VGBY2ECeEG15Z0mdzcBmR5x31mWNoZyI
0nFdwHFWAKZe30zKxFErOhzWJUVBQ+5yMdjNiQytavq3ruuTerJFK/dvokeuaQWU
oNRIqLKP5wDcCBOu8WfiMG4fiNlDucWquSqdrQFcXFR5PlT3ch34wIZNV5eGr+b4
JzlnUoaxzJViUqQsKrVCfHE/LheOMz+jeXpoRqKyoRWenEK0abVn4vpJC1a+bil3
IuXm2xVRykUIUlvQDUxesR6y87R7OAQ4vDzoazEzidWCNLujU1h0/HFX/VipK1TW
P7WQ3+Q03WmvXKIe2eBQeEX/V2O0yWI20G06FqYTXEz7HOzI9wSldZTRv8E1wynE
+SbflStmrCw0kViW577IQo3Ih2Ngrj1cL4JcfOV686yf4zeTAqGizU/EgfrZS4FV
WI6B+Fmf4Da6/lTr+TwIBZh5KiDAVQKx3FTiem2P4Re5m0ZCSrJpvxRAeuQPqkNs
sVHJSraOajA6ktKdQ7Lc7grHynlom0mcdDV7ZxvGyzT6pegO9PW7oqQqzwxGxNgd
jzcmg9tOev/Mwcx/VuBl+k5GIb5IFGiHPzzO/PKgNlBUTjUUtmi623MYXXEiQgga
O+0Bv+w5OoU8PzGcflRovZ7Y4pXUNvl/deR+bkEn+G9JtmNxor7BxvhyJ29v5cvU
9g4skSy5gO17a2TXtaOsx2Obsu777QuutKswM7FP/+LMGCumoLacIBGxXHPIo//U
baDCLfVwXS+7a5ClJawsv/b+hlKcXT6SKbArLGJRHcToqZ6GCuVB9stcGQapfbxx
SDg7jlw5Up3zJoCIyVvGUe7Rs1ww0+HR9lmyjP5+iwPesE39h/r3Ao0p7Zw2nog/
Ahx+V3cmkba/RQyojlcS+TkDDnTghPtt2Ai7y7znUwvbckT4l8XaEwtNAJkP0XV6
10sCwE1I0qCNpV/y4kiFpuqKUQ4IOiArStB33jYf+ruoZOGw1LLBbNTq9H5f7RhT
cYZWmpAIs0wKoLHr/E4yiY36cRPK7qYxq62lHrv2PHB1JhpcG+eN+wHMivRPPf3M
fE9RFYSD0cHdtQSHPKbUsFogpKA0CcZM055zYMaYvE5WneSoTBCZTjFt9a3VkW5i
DYa+bfyfTwRzs15RnM1L8Gh8/CbFeQKJrJfdYHJ5p6+dhCy94lg9ct6xBKi6pO7Q
vUTMy42V4lpSTQZiCMe2kKw8vk/8D7YgWhKvGTo+p2K/QuxpnNkNGmxHDXE16/BS
tdy6vv3y3OFgiEGdrQKSy4a9EICzdRhJgxorO6L6WCIjcZlVfqRpHmW/op25/FV8
JYcMYkAYtBiy3vR0ubqxXfDtaDZg01e24o+jETo9rOlxKmQDC3fFH8UvrRmyifUn
NkNvrqRm6JVXyRo83fu+Rt8beTsG/b5hKz3sJ/SjHidUorirKgZZ58SJ7d//fHLG
48/KD4sarZCglIbuG6JpfHv7MrQh6qW9Wpgd2XJeClnas5ndIfqfE451yqRl8VeQ
lQ0VkcPkI0gJKv2VcIPg7yQnuOtNaHI3Z1tR/IPUUFn9SivAhD6QpNEoTvoxK1Sj
wymrgZdpEJH4lv+IjjUo+Rfekfxgy9WvTsK1DQvA7wNxpcBbOCT9ANgkt1aE2d45
wGPfJXaKZSHAYoyESalgVCHmJ1PMbuWl+8ZeOmzLXzQGIqCV0NPV4gNowQUhkptJ
jjaMf22fO3hC+Cv8wokAD/zjMXhRyhqYeZshozDWcll7P/D9Pm3WKW42NPQMASQg
dUUTb6AXw4cKjj66LdaKQlwlteQaHafG1QmATOHnmMCJwOgG7iyUHFyLNfUPhjuH
BrT365zdav8MhKSeCa5AfjDdnE50ccy2YpcDsB8TGziHcKex4Heo688K1MalQRSy
XfNT0GO/n/atTt+RgAQGKbip3fvsJ2sFjpmQZQFMiy61vM22MOUMty73YqOitMu1
PCmNboTaIFGtb2gVeLHAyiYKJtPzl5frOVoj/yV2xbPi903Wmzfn+yZEM4c2PJ5N
RTBziBQM943G1hWKlAEgksxYrPqqg4RDSiacFSX0hvY5nIQBI0KZVHHOmX083SZo
/iLpp7hfXai9iilQ8qHs0SYjI0WkXJLcO+ikx+IFtsdX7gcqUXAlEXHs/CSthD2P
aqIb7/728H3qQ3BoKCLCxtxWjdee19lEmBYPY4ABmxRlRVN/bFuaAqjz8MFlXsx3
e9TNsEG7y5c+DUgMME0WnO/k5FY/o2K6BnqUOsI3BByurxPiNAcdLeSiC+lrdKNr
Kj1zkOFgPkEB4Nw0n24RgZjD+v3t/X197j9Ow7n6hhgedJrXfjeO/73EuBPNHyac
xtNzPGoMJjgWNK1W9Komf3jqtu762RLE0yahF2Z7u3ZpS2NadB1tfCaKKtAEKu+N
2IOZ1xOAK6ZOqIq0NLYArzQK75T9WTnraR6K0LtZ7Hg0KFpMZIXotUWgmRMFyA02
s3sM06LXOwO+1RkYx5O/G+vfFYYtXcLnQDE9gXsrygDkXQs6aZRBiRElS7+UXctT
eVQ3XN2SUw7JItDOkEIFzgW9MbE5BttvzlQ7megQyCss0HTmJZ4bIgNf3j7JBOii
h5n0CN6tmta+KC+K43dL9e0jGXoslMFaXlDEDApkgeX0vRn8vGwt1V5kEoAJrrHt
3uJN9f3oLx7KSOYucbvQqxMS3NE2en7VWG3Q5N1ZSOcRCI4S6/KYG/pLpDCpZ+V7
rqQt4hUDWDNDWBUO2TeDgU7IGKoNTeLsn5Ls1lmGDbyN1NGak87NZQjOwj2rjYfR
hwd/Cp/PaLFwDhXZMfcSp0vNm9N0VdF3TL22WZIAqv9W4uI+5xyhXseJzj0md1s2
EwKTkVyNGn8iu9rNJsr0TEtZhX8Hd23iXD04odDm0dhhisYfgvyFFEcM6THC0FSc
6SyXFB4Ww67gnSh0VGN9iGmaCDPIeQqWDVcC+u4Nsspa5Cnqr+vF1c7OmzsxrRdp
YaX6onGDGwvNtBoKBU37fyrJyFRYxeaW1XiLa6/p5Uom0sc2D+ztS9Ph42iSLHZi
ltNWpX09tjSbbG/zVHo+st3SfGdRBbDHADasZtxminzldcX81GyjRePEg+DnoVri
TXdMk9NJnK8waNJLT2FYDfzK0IW7b1OzHihe/Wx0zBIADRQ7HlwZVgPo9Z2jKD3u
La37ZtJfXYbWnWGc3836cQDJBl76eWyIzBB+Ce6lQD+MzVRo4T6Sx0BYqAdgM6qf
KGE3gJ59gQScycfU8FzwdQglaWJty2iNFmYm52WPCrtCTX3DjBBDaGpBrNjpEfJ9
NFIHj2/8ku8awBjo1sf3s2mW4qRExQ5GWua6ocp6PLzGgYNGQsmFuL0eeyeWVIBV
P3rCPHgoc1LaG9coKMdZyQTiH7HjTUEGjx6NkdGAFDgl7DcQ4buXVbd7kouf/Oeg
pdGMf2IALVADnjZTY4A1YCaZL1Flieuxa+VpqEinHJSRpDY0JVxYTkvOXZzRhXyd
rkE+dozOW4UVJMvoW2hhhp/4qKycX6Y7LnRTVXtI4xUtadunV5zhFDyWLRA5gV1G
aliK53h2lOg6vq59BKh/bdlhAZSTsvk51hmmRCinUqG+66ps5u+gbGBdszPO1PND
dCDnE2+3xch+hnSx0kqzohsCLXj3tDF/z7jpmxVy6WZFZLof+75+2go7a+H7xd+F
CiQe7drdE2M3bsUeF+7miUCOYPssh4HxkAAGzd1MPX7pZdaYG6lRXgK+wHnq915N
LbP96tb38AOt6rfmX0HQW+ZOs/fnaQQwGk3jvMD0CtBZKOBCv25BEuun+QFAPBZj
C0Bc400GNJDikkuhlc4b6/1vvk27RSrZV6nFdjJQCib6BlSECLp6yH0TMLs5LHGk
Ihd7yBWKIZvnDhq1NDFpa/yRwopHHPSDRglyk1aXfCdXmKq1q8a08z5sEyiRepjB
M9jlvJkWV7EOp6DYi0MMfsuUR0Q/53xzgZvg2SYEoaJEgknc5cIuF5rUGU9WLmN0
D9X4Dgw3Ef5cWPtFuQCBFZOX21WIieFUQ+qD8qFQe8N94EmqVXC4zRptBwYiUIZN
4CY3p4SC/0ueoC5f88ANSCceLC/00yEC23ik8+y9LW3TYMDWSZvnt1eRaCVVID9q
Mbu9BHFt1/PEK2Aw/r5FIy8gZo9O0OWxFRU5j2qHaRioVZKAuadc3F2G5LZFaWbN
t/r7xJWEQoPt01AdcVE5Sz5DNLH3AVD4YlXiR/ljV3j/8WOY7CSxvbB0KAO1+IOd
DQCEU/WSmArUbWLi2EuLZS0en+lMg7iFQzkpAR7KyRkk0idmR4skqHvwFXen0M3B
t/Zp7Hk8oPs8IGFAq43qrdiX5TO9sVZUebatRPHJ6Qva95xA/mcPvTIk89Yzl0kv
4W94YeSXEptnJrlgH1vuFKweX+p0Cr/gh8Etjgzmc2cMPhYHWyk7POQ0/UhdXeep
ZrnFyQcM3+pA2NkAfZM+lvWeueDiMdfYqtOlqGydAZUYqIoPLJ8EkFj9qAmD01/9
0FO0eY4FXUbUv34IAFKT7XzeNmI5XkjWwdgTouXTZO2GzENvM0JflKWTuprJDsO/
UDzCpzehzkcZVIPzO+pgJeB6qe5Q9l/QmmQa4+AtcxVXn6E6a44lhjqxX0HPp9s4
HIC3q1wbdWkdNUvUDbZ0zlOldDjNa1DvaXZajQf8m+naWt+foYa2TIq8NkoxhKqV
PAct0zOVOO3as7F5/wlL2czPCWsd1PNg9OoitNQIKghzFzPY1OKlvpPPRzQda85a
OuM2gSmvkI1IQbWlKHBvLU0CC15j758be5gSs723r72tsObyXyh/43Csqjl44amM
rpVPWmuMKj9oPxhvyilJf5TLoSYwve4Ih116Uu9pQ6nhd2NP7zZPeTwb3M4oTZ8f
V2qkegUf6uauwnTEo4H2NGv/ef9J56qthvTefUMMbPrkkOLudBx9HPoVOYsy0k7l
QQ7jQJK+eSDV28ums7Q2bfpoIyUkWD8OAQk3OHUpeEJaNC80VbnpF1aTHWHZHE0v
8x+qyBRhhIWEbKvodp5fZ8EEJ7uiprEar84J63nwEXac/6JBM69ok1H+p617sN6U
NpfB0gvMHhPTPE8hfOpFuOb+hxSPWVrxgdGZv8nYOS7OmA8I2DBfeWpxZKqtAUGF
mPcVTfZKTXQpCh3KT6/6sSsvPTDm/MWG1D6tl/e/dlWQAaXo3klsXQcWTr2HBWhI
5neoELiLUHfKwQOYfaRy34E91vSkAdg/lFJ8pyz6WicQdvXTxLY4BTGmxc2ROFI7
ZQ8FmW3xtaCNfmwlPjtswWEb5nPbBRB0e5cuV1NKzopp6C9xkb9QTMvjtIiMtA1y
x9KZd/E+vMtEU3+TFFNvOpeoTPHsQxoIf5tgLZB9WU4GKWQD+KE0IssAzg3LICJL
DubPEslm120CzG+78rsWEDd1Sa2xdYIvNlitDGnFe+Gnm5AaUjyPbKd+fEtu8Bu4
fVHP7FnN5Ixzwzo3+Vb6wFJEWcqIxKBP8kEdebzttfC9id814j13VU1MRL06sUsA
NbGpjGkyiyzm8eZnYp38mSvgOwzpO44J+4oTcotWn7ZF0/GIxIIykIB8D0ckDZ0a
RKvxGDAVr2O8krVruV8Vx7gfsRH+B2oSYtcPiPD/l/hqBI7INc9gbuIpdRSCkdYK
NgDRNito/3fg7EuLHSkV0h+JqL/Yu8jnJaLrdrjQNKnpnf80qLjJpHt4c9fUS5oJ
TsvFdBqhqpQySk2zmGUJNWOfBqswj8aKg6ZtIBlfkSkAa1Ir3gMRfcJxq29stQS8
BSIjsJqAblRsmNXE68ZFgLCtRZbnzaHV3w0SH24+Gqx3fsHO9cGYALIxLAk9LgED
wIoT7WoDuE4tTZvf/uIpjp0TYDrFLtCaJfa8PH0uNFH6QEeWbqeP2dMEGrci86hI
+W+EBCVUZrRXeSIIdpgl4YokJ+XUrQgkzVUoGJ3jaK+Ug8BX+sqFTguQcoAr1mUe
nSUn/hReGHHGO9Y45RvT+lp3s4jhh0T3QF1tmSHRPwizVuIAghXO27M0Q81T6SdR
CNuiEQwPMaybt7n5NLNctrd3G1unEoQkrZWCCU89m8ecWbH+yGXrpgE+llveoiBM
RZ2CUx8JpC/Fzx/FipqE/C/AwmW/4hNnYf1IkcSCKgZFJrqezygGPM+tqeCmD1f2
Y8d7Up21Fw6t7BFmSJdlBMhu3m0sEObrQhwbMgnaLcDxvZrFPw4+DOna6Br6t8j8
SxTIDyLlnFF8XmW1NVVf92bxSl4oMnW++zoBsdiBi7JYTeIgWo1fl2k05WSU1T1r
ZyQT6337LIszcAdMe5qYkdL5kMXd/RQO+50J4J8xk6fIk6BUnAJ04AqOMZnbUff5
4KGxusug6PCBU0mSoqc/bNWFg62wSCsqIutc/BVILSS38ftG4pzG26PGl0BZJtSd
B2YD/e0FitvY9IeH+MrNv0uBzpmJ37OBeZnMmsO8P55V8Y6FUcRhrshWggkPi252
+XVOl3v0R8O9J91dPHP1UbMlCDuZbiDOTfSYX1dp6CCvt9bgBF01sEGxEEVmIpFD
a/4biZsrHlYjIT4pOewRaEwLDv2ZlBA75TScHjF8kch08kMEPwV/uKxc/7L0aP0p
q07uHl8p11wAYuGKnKJ2eGmnISn6cDFWt0QhpKOjLFOGbM3sob6w0zOBeSXRXCrp
Es5U9j10YcQ5Timb8AcNer+ICxvvjSyvi8zDklWfl7RuRKp53THInV83ZuzkOrg5
LHLfhEM2O4CRX/p9pnTrfBZWFtUe0ggHGGVb/aqyyDL5PlVTrkk1w1cLaIxOhfk9
G7+x+5vOzCz+QbgboSU7M0vpAVxXVb3+Rd17WoK3k4wpsCN40gyqeNi0eeFqQ8+j
XPECKIz9uMEqxJUblcJJgg3bwxNwzyZLDg6AFeO06H11QxxCI/1aHefeLjNawjOh
CHunodjn36m6nCo3P24D8q+oFqVj1PhHhD8FSV6ea1Xl1QdCcuhPqoHQ98wbAXgW
H2PvWQhJnk9ys2auQs4O1TdfcsRNp8tVwlt+kF7alpuwIB+gUMJAcueRbZQKu884
kkegLqxZYSW1xj0I3XLnylBChOzgjtLLfHPzLiSnBatqhq+agl0mmAyqS6fvcCoH
bDzlHIfK0BKuyBMOeMjj15C863nJ0u2ouNqtLm8S0meeDFgLYY+AW3JK0ElKuqsM
WOZuLzZ77TjpNa4c61HqGnwaK83BmHB4OD8Hyweo6Oi5ZjQC/VM3rvSVtOoq/MV1
mf9zBngrJYEO2uuJbB5tINUp4VXH5LzpBRmx7gWRpGhJ35A0Tyxk030bwkmMAtBe
5y2i+tf11xjzIxwmbzkUMJEWWIRvo5Ve71wJ3DpqPegJUyOPDiohLo3urgq/ci4W
murOPX9Ctnrj7ztaUoC4nVYh/fbwp1UN0ylwOzxYJZgLVgW3e3MHsxm65tXou4mI
CSQGqKYDObk5qNsTdS5nbKhozZmSzxIFkskIBek3xyD6mwPdbStOX7hRR9eAMlVd
4i7wqAn18zBtIPGZy+WHT6hR5VewOz988FUfk4YV0uIr7Se1Tbu0768HquqUQLN2
5DKAsYggf9bdPZA4tQ1z3m6YJtD/2HRhKDg4dfw3WjQPAJFkQjLUf1jcLXGQaZ7N
misA5jpjVGYKAWBBCsGNb4fQwIOeudEB4JTS9/WsP8hPWW7wQ3PddMq29BL0xUhc
3MFllJEVBfbJN7dxWGzOxGrKEaLWMbJKg59UuYhCfBaBUDNp1hD/gP45TIodnCfK
auHHx5RDtToRovs3mSJvLR0wmTWQyviMeoHPbbIOqgoOtX7wU67F0kB9PW5l49Dd
EKuxB/EcJcAkigicnMF4AdQ3tyk0nG8W1jJuvZpTZ9AAoAhDxg6No+FNAsPiSc0D
+uYdkgT+pYnSHB0nONK2mWJv7RIP3JdAPFJ5mK8Jj5+SXoBRdF/Kx27CJDeofTll
bU4bxosd1oVfzXDGLvwxzr5txHcLVl6MLEmeC7mlQBQNM2mMIzFBNtWci2MiKdVs
yBGjV+QRc5ofMUgwfjQgWDUKXZ1O0K8i0goh9OZD7iKi8WcHJ5O1tJVrAzAJeKqC
wX1WUzQDEgOYJo0FolWsXMPEfs8lTYsARGfMUbbNznPRzO7oTvvaBJPfGa0bjwm7
o0FE9nd1z6+rdOt/MJ41kJmfTjmF8/4BCaaZA9px3KsPjBSsSMbYLgmhXLIky4BE
QxOxeHkNzXR2V8DHEPrlhwq3NNwXny7AXDeN+aCTdzGPQMKCiBfWUkygVwvyK3yK
gMQewpNmecnZNJFiRfnJBqt5iTbCP4xOBGtRTsTuQjKKjV8WLmturK1j+M8LLcSf
TXe4PT9NUt/pS2H/ZqhYBqJJ0BFv7Io2XhMuHBD5D9kfoTraY3pNzTdcdH1LvkQY
B0EmlbRUMpnswmvUZimr4cQYxE9OhlU7lJ68b2ss3IVA0TocEqn92Kpkr/BAq6Y+
8pCLRtH+MkR0vOFXz9ee9g+XskBmIjMmyN8I7wY0vXzVw5Rbp6mX4VozMvlVBaMv
o6TiHDatHBXdyf0vU6ftM/LSeNPPLB0Xs67I9v9Lzr0esi9/nkFBzozD952v8IMm
Jk1sX53zCVUajx88zzuEemKs8XehFQ3sKMDz+CoKCxHp3tp/9Jz5fdbOLafCwc9U
RnAd0NIxijIqzO8T/cCZd5VQnCcMc12gTU0iilebLfjyfb1bwcCID0MUCBbuV3sp
tiePW6a0C5NsHh/sUSineuse8R3C9rwa/5FLqnLwnmw1e7n5JKoxuqqLe2Ta8p7X
OwwDV9wgoBwAFC/aXxfYpO+As+wxUKAOIr87Q8gU55ejN0OcXd4BYrNtLIcGpcP4
CCqc6474oeDV1QXaXki9OUDun5ne0pwtEN1bqFJrWZwyRo3U2QLQ2muxVPHaWxTa
s1lX7uLcvspTzs/XGuGkW6lHkNay7/WHdn0gf/M5Jzt79nAlL9AlU+IfKgd0KhrH
IJDZ0Fdp0+Y9Vj/i7PEXpMQb4Dqj24axDmXTLY1kvc/rDjxAQoOK8JGIsuuzSvR8
E2nUyuuEZDXtYjY+T7TbfIOqxAM8sR6URo3CAjmWybA7QBArm9Tpv5uH6IEZZabw
PjG2CUM5x+kLiVtk8sRXxaxD+CYofNWmIoOaw95T6145M2y5KrQJT59FuuUMBsdD
MI/hs75GqLo31T4pwUZ5Ij6t/3djXdLHuFu9rptIgEIjmFh4d8BEpmwU4QsMRHwF
Dgdpd/DbHX/BP+Qi/wFjctsfFuyOP5DdfVWlEB2VBSh+5A9LZRyPro8+KpqZUOOC
1TmkDbPEx6w4QcqFktzHZqoGDMXnZ3SdRvM0p3W6rIupIDhxbRZ0V4zcq2clgiM+
4JRsNp+pfnnNiNjpy1aCdagNYZW4eBjrwDgCC2+E1D9rsaApwmnO9jCD/XrK0Ghd
d2VnxOeEYJaef7YPBbAJxTlXfZs5FcCC44OYh+t9/ZHiUbXED8FRQPr0CL7WI6aC
hocSk1e6e0VjYdwAcsPAwMrLQQZflU133zf3g4yDXAuOG5zFZ3GB7jNsCCcIV41+
r9rDb2gLuxPxtS9lt9/D4Xztm6qZoPIsOQDNvDG8viYnaf2iD9WTmHYtCU+GeCYU
ZAmFfVY3IHdtl6qOjXo06thbCFuUkQt0LJV+x0itSjLaJTPT8D8NaQIHr6zfScY+
9hbnKkwJfqHJgzwPBvVtyK9/r8ke0Ra7MPlPdHZyO2+oYqdOxJIEP24lXR36akyM
QEvBKE5pGTg3eaG//iLW2YPVFicllC/p3cY2V1W2ZCLDsI/gUWp3T6HTl7oPenZt
EbEBkMGBilHEa048ZTsKnSANzziNXA/9plYMH3CfFF491WCFf61h9pcGOMHihym6
qea9XOp2FoXfiIkZIMpEvvuv6dnlgTdjhyAPvruWd+6d5OxD9whRfsVb7rkXFaZY
9z5MHpZ1mLZTyZESmXNxGlq6j7QPed2f1yabpw2RoKwwInnAnSrPk2S8HFxR5hnC
zjFmerN6iV7un8KaACmjxoXUT+nKy3/vVwOR+AouVkiNrSaOQEWJEnF1ikrHTBHT
eylpe2Qqp7DEHBPxDWmAQm0BvzUJIaCh2TFWkcbPyeHJzsUf71b2iGumkKigFFKe
25ehh4LFxsqLoguS1aKxPGIyL4SOygh1iLEE8kPYy+0xXMm4R3M2kQosBGBT/TDN
5Rvp7UwUAYrLfQJGlLO1UKguyqWOR/fXGuqfr5B6Co8+8G3mLsxRvCDOjhKFBacU
1tDMc2ciKseiRBi8QWTpeHjklxPRwAYmWZQOIlNeLuCPoiWbFXx1p0AOq0vgRAGp
DQQ7RJxDJJrTfy5/HnNoyGng+hI5uIMYXWIqUxoYO3QmaU6LC+c1SuWlhg8LFCN3
Yr7wG5qcT4dYiroDNPm4eXF85A29fRzudlUMVlsGFTsDTUQ5aeTz+/dGqPKU8CJu
CQ18DYNg7jRsLg0X368UAJKWuyn98TKGawuD6ebaMWv37ZTAeKXqm+N6LOgKrIWG
lPdV39v6TjKLMHexjF4NaiZd9qonAH5s6lPDnqNlBmmGl1DqjZaxIwOpyN4LHE6j
Ci8YMaE3405fun/NrWO6VG2dkizleSJ1MCAqkeYhp6lVjPx8aa4b37RdPSuM3BHN
oi8w6qGIib+EVFqlTT9Ncr4HwoL4I1z39DV/ZWQ2/UKb4UUzewJtbYIkFgp9CTO7
Q9MvQqVLODd5fq93OwkRhEQdjLkJNazSVz8+5910u9MJzdYiCTX6v9fLm7bN97OO
Y7rj1rPPT6SB1eUU0cRwHpVPcSs0wpFtdgkydssYFmWyBchWsTOu4BZA9SUu3Dkt
gQTAI3jSBj6FJ3htMCXAV8KFLgGksz5/h9jxi/M1MDPuCbFwqJjPB4i6OTRProxq
BninPdAhJS8vDE4TcvRRXsREWNghGIIpDeIl76btTuy2t2k2hAMHHRzvmx3qoIWq
EWMfqKVWzsSGFw/dvonK7RrWzif/12DaZT/4KPuoyNkpuGTskPO+xcP28csGIiOq
PW6ouEas2DabKgzA1KdhwC9Uw0xM+XdrPEuNjCNybX+O/cS6F5X+MpvsepKnyrmU
rI5uA3S9RC4aZwfX8pl2LCoFva6Q7L18wEfNQiBe6UoHwT5ZkP3smdBm9qX0cLyQ
6aEzuM6Ig0bpG+nJXYtxHVlBQvH8NRKbkSmqeRpsUSjBQcUYy/jYbWgO44bAbh9C
G3bya3dKYPjlsvX1/CP4DqBx8sngNn4etaEUPHTZQjvbnrbc0f9xtWGFuQjZR2GD
uZo4VtqT6jbRU60fJfKyY97ZRRIbzPgqAWpj6LuToeq6CT/087/tirLpg8WUIw97
KValb/Oxw8pJnr8co5hQ+vbvmxpFbhXyAkACOj488R8PuO4xphcLsTHQnvdbUZy4
4u+c/eJgNBvKvETqzBdvXMvKEOgZgbHkBVaXb29UjwhJ+K57MWqIiqGL55wlrwKR
6e99Max8drmbhdYIJVSGmQc/jyT5lVotPSrLPEv/8FZYZG7caqe2tl7RJfBzOb39
A+Z1z6FIWcXrG6iF5QG2PAHl3JxZl14peCDPWIGmW4byQkZVvV4JOKkgFMxw++o0
6NB8r2wHjSIs8vpf7FmLZIeanKOzt6tq72JxzYgc7XTH7Kiv0AtcOfylNqg/wA6R
pQR1iYEC4ss1Ao7iKC7XmlusU5y7jbmt7b7cn2K0br7xNhpowekM/CBPOc2KPiaY
10pLQiFFh0wI1uiLWLiY4sbm5Le7M1zazKjXzwwg3QizACJQmhDsNaLxZbNd+D6k
SJhsYTbrkr86HDcDHSwUjqtMqlzt3mamYmrYltHi2v4LteuBCZFILuJT3hjaIdgo
mxReHiLo3AGbddIO1ozuTDpRcjHVw/qAoQSVVXwtdT8sXWuPa8dTtWyzyw7bMaAg
GtWE24aTYWwVx8ynvWfncPP36BzIyDpsrwFJx+hib6AnZWMin4oBQSOez0M47PpL
/p1pxR9jdZNsRSPFcMDTdKS6V5q6UpoYEVbQuZlBlg0suT6+SGkiDiarrhYY6o3N
UzAdCi2/JuyLKgy2q+p/peLmXzEXWVcXngyt+tl1ZZfplFAw1n9M0l3z4Zs/rbvo
3qNQDcbSU2PsMECvHXfuT7L1X/Qww/KLGUpH/46+I/jnmXFSceV9s58qG98ubqmU
pp2uRI+04WeAYDnMEGP6BlrTWhep6Ges0T+65TYGcM2ShlMeOCciVF3mpEUTd8VH
CkQV1A8snSy6jgXI7Vsoay4I03f0ubsrGYuLoTDFsPSnQSd//3EkxwGpSN/VfzSh
fPdlcZIsvxDW6STU+4PlmRCCi+CUwJrkE8DFn+vMbozQMxOXBVOinjATG5mdytLe
OgedcWKMJ1o+JZ1WF1Mh4x/RFez171RbsfzNZqU1xdAW6T0MV73IzRJyCTI2K56z
jlJjaPrGIgOI1JFT4mgDk3g27oheFLdbPBpFgzfMY/U0PYXtKXP84q3Czc4huhBR
emiQuVMgdnxqrYnRyFKvrZRA9kxNfwGzZabrRX1zG7s+xo+9OBC/1GK/l09+uar/
VLEsB9fyRzS++gS/Kwkd5yEwf0VnxQiWelf7tcvokTsoGPteqLER+1eC5RJ/JDBA
Mnja7SzpGuOa8X5VP0GlyaswLy2vIdsejxLN7beV68njuz5xDfxP5dWpLYktR8EY
g+MIANvBkPLQsfqkOaGIKGPLtr6TFQKeQb2tAzdTZ/s2YjpyoxD7z/APtIR7PArP
xoMjVPsxhnXgqo3XVlUqYCaLvfUGcNfxLqVB7N9O8x+kSCjiiwASxfHmzBP+pwmJ
6gcF+vUcz390XVI62ny7Thzbu19lKlK/GLpU6MJegA1pZxlXAxw8GYYwuL/gxTFw
1jAhLFFgPzG7qS9mfGLlKGyJhOlwAeXE2FnUIGXegw2UoPn9TAiW5hjXytU90rv8
MRmFFXTLwfRhDAsN/APdiJaK7vgZKz5tqm6NoQKg/OhylbYFvc1llP/o9lThcuvR
iMUQqYpI5uUi5s+15HTmwr4AlqM2DyJQaOJQomm5IVrCG0VEUXudzFjodTeUwdoB
5H9s5MU1bQAw/Soi/PrLstpahv4XGI3kQqrDjV10l7cbwq9+DRUa9lto7tIGz3ah
eX2/inQjSOpkBbURIp9dooDgAipsBSjOjrWmLjeV6RoWprgzDH8pSrwndqsankCF
CrEBK54NuxxmDPUKMtyMacuPff9G8ia3I+DiHyvCGSB8k24G/NhPyTh6rW7NUwdf
U8+NVGvisa73q5UXlrlFpqeJULlWWm1dmGiI4pOMoQlhI/E7Dt+PkjXmJ+ZHUTP8
jyvvIXYsaU9NQLnxXJHeX5D3kVYlWAq6ziFfwczUbe73TsggyBiKzOmVkYCgqCzW
YwkH7rkuSoF1toCEets6t80GEpIRPic69m0P4NHAr3pEIyxnV8APLlf66u/ItoDN
Bcw0nf5dHhXoU+SjOwbP7DRWtuBR7KKZU0GNnwgNN1PNjU46dLNqEpJkcjzoU+rY
n+BUk3XOgdm8Zw8FDxNOzFy+IgqxWN8ixuSu+Up8DxntKfsQaUWSVL/xBragwbah
xaKZ7MSeZXvIEXGXz6ZXOmdw2oIDAPuaczOgm1OU/l95X3Ct+2ufUuas6Phkl8vN
jYZQkM2s0pOuiWZlR2R//3lyuKhfXGhaFgvKL7YW2jXKAZ8JCRP4PRk/YXUaIRg/
7vuLzW+Q+UV+L0vvcRXe657NtkDnMBu8hqWclYS8Qlo9oaCHVvFJjewz01R/lqH/
RR3ASlcyeZdURPYDMiHxlYKnYB6cEs3yy/g1TLtEI9EEy+71Ec6XvFK8iXzWG3aa
a77KcLXnGYtY7oazuIqKlHexNSOfbrzizHgHkvp2uP+WpcrDd4huO1VWT0iwUBM4
kK+mssmxewWkH0VsErUe3wGCxj6tdkEHSctk0sgfRsVG+Zqp7w0qqWSDlk7l4YtP
tUKdKeonYc6MR2IUsU8tT/zVkcodNgJcYn7EmZYXiE8BWBgaFkwTFtSgxspmk/QM
UGB8h5ucRAiKN47phi+U8nAup6cIYDI3A2aQSAWO4+WzBT6zV0S5W0kSVPrfICY5
AqngbyExkmZP6l2YOTlmfGN5t/POTO9tVlns4+edL6oiuemEUBFcWAUgB8pRaEpN
G/MCXzUkNA/PKfaNhbE6htJV1GF9raM8TfmXnKj808xl4J6bUok7afZq25dbgqHT
7YGhf5+PUOXyGDTNouPzj5Ewoz3Xl4BupiKF3fasURlmf9dxGwIUrRyBDp8qvoiA
VQ2AKsaRqTarkWtMqRI8PuZ21bUqxpzHDOhi2FhEExyKPCIWGF0k7lbIqF5x+eSj
BaLgXdCZksUIUt5Ds+dnN2sPGVJrCyhbNH//Ji4Nn7RdFQYvKnUKLw8yg5koX1Bb
EeYPC895o0rGJQJHBEbD/ktprYRVSwQk6kKMzw76aFBMSczebSGJzcthKCH/PjMl
E2Tti2zVAe2zGR0NDOx1Sb7ijMGzVRDxY5D8xNuWk8BnB32o9/xPW+mS1lWuo3gI
quKm7Qi489XcCc7lYR9HcOBD+7dtp6D8d5fOK0EEtjWwTjgqYg7mAme00DJjQlBa
uGzizg4mgd4usSbS1FwQ2XiHCU6CiWcg/uEqLAQ5j3EZ3rddefarMo/e+rzJjHLE
i3E7Gcgzku24UY9MpfQALJmjpzD1p2sq1UaRhDE97UZ9ZfRvMHcAlNzklonA+YCH
ijRNvUh4Cl2ed/bCEgHx+Mpl7CUcKjICQ8gQnnUak/D8CMyIZonmmnvQPP9i+aoD
vcgvnGPxZAe3cMut40MQ/wBgXvvDmTzXwX+ngEQn6UV2aM/06nlenLDBB4kiyFOK
TPXz954CIGk8ZNibZ1Uo3hzC5Uo+0Ou6EH/phTbH6zwV+ZLHairQ38MKr8s57Jep
T11JVWwXMy0TV33Xg5Y+SsNL7lEubLCjm1rVQ8byPAa7vPLuOc41mnKsMY9MujXW
2807LftZNC5z73kbEM2nlyV3XfxIP447HBIB+Nvr1pZduZqkHR8/3aqTrHyxM6GA
In8reZ6Rnhh92yQfSwDxQ96KJt+eUXTZ3ALk6H/0Gy/drvdmIlUjgbNSdLCY6R85
Fc8/J+NdwVqTQNwyKDLNypRiB5igL4JlxoPvttQxQmxx70B62ngVU/RB6V7l0vHs
ZmHof+nWMYqg7SEbcGxdVcLQvq5uBci3nZ421mwxpps/4K66K928qn0fq7sAXFpy
dtIGUezBcO1B+AVTzjlUZGnhwLEHR7O3RL270Qx1fBXxh5zdWITQ83yxaTp3pmz7
oOIIL2iSlU2X5bNgO84Y+RjL3WnGskK3RvIffxx9Y4/WIeBcJKy6uu+lARyvoRHO
piRn5nA+ztUt3zD5oytfEvEg0rIW3WaHQL/EB5MuJmUgEH2wWaysA5yHEuTfaQd1
zR88Pyz0FgA0tvpkvWlAfspg9XuxwOmiejplHfPfKQVrp9QiA8Jgthfj+vmCuzZQ
yI5FRYjs4GuvJQ9lU4hABCj68dmhHAETnmvOYFLq1UwXOTJPL/J26Ecy+uX7zbKs
CBdsoNFsJXS+1aGpGM+XZXaIp8vOwl6hJVe15YJaTAmgiUMBtH0yQ8bwlTY1MYTb
teOOwOAuGArLYQjhL9S2ewZ+E5xczGBYAA4QfwAyCik0Obi9TGqr8ToyKC5vhTWa
JzwGLfqIffSo/4PDoXYjn2BucFeRcg38UNrwQVnsBs/yAzaA8ixZqClhkZl3U34L
CxTwQ1u+CIHHSMYhRtcks7oqaYEwaxhFQW/2pMlpu42h35PD3bOvu4tJ4u9ERD59
/+4ciCAbCadHbumbDuKKcG6XkAYdU3+lo3sdYCO9AfeZvJ7RAEODi6FO8wfOKG09
9m1A3PKKXoY8qnRvBCg9laVNxHBzJFmgqvU925oJNdIhCiY1cRXN+Kb8rONWuuz7
dDT5hB+Bl+2OCYg3p1V/LjW2DxRODAJ0+eA/8ayK7on3e2Lrm+KaOgHFzX9B5haS
VJZ9HDMiC9t+7RKS6iNoSoIxdwS1mIW2CGwmh8Vhi9GGvASN42H6Ig4ddFHE5jgf
n39eyTWPBZRrWKC2TfA3AN49Llci4UH/ewHfxZSxie+HU/D6uXcLJdIYPYsMpKBr
74yZYGbwRFe6zcvnn5i02a6c61nvtsVGvAPdbjSddbQDRIpt6LI8lX/2sa6vwXLz
TzYvbaH0ftlmik3X8F0iF1VKc+cKSRfbVqpCf/CvFBMJh3zZYNLsg1i+wFyPHkpQ
ey6HYYGw0NNr1qTRYWtdSBU9Tald/nkesZD5sjJZiZvcYOy4d3hW1Mi0JWIADHKk
YGoxI2FLTa3ryc2mRub0x500kPK15Fc5vjzf1UywNLq38rvX2iKHpUjX/ZQ2FNte
VtkeT6NzHpgApk4+4lrBFbejMiBa5TChH4/W0q4oTieI79zr02JI49dZI+e2OdYI
wJrPiECC332SRtTQj52ZMpdnlC0nbmDorTU3PpHOMH0MzqXwAz3VZ9B6EwyXPryA
C4fSUqHwrjdbAxHqQnwVXmCMkS3eDBeGmc2G/fBkCFGvqtOfWrAfUW7Nkr6TAWSx
4Tv5w2fKe7sZAJP5v+oqTZdAX4K04aCXMsqg0cd5kU2A/VFiwOA+ifIctprZGMaA
CNAoAcjn2W3fJFUWXyLEjKM20W+QEzc2lxpEbf5w5NO7VQnDp5071Mpwpszi3r3S
HAUReG0W6U9awSSkUO8+dVfjpwxsbich6nV47M7pNBj2xwtRJS6cAWKiwv8tZE+P
p4dE42G9FMgV+FF+aIfPdKe2rR8EXOGJxRyDFQULYrc6CRsHTH0t/rHWRsvRpMUf
4YL/LvI2QBf6gjmxg4UwgwGeIJxb+jNTd+uAQO+qTqgq0po0lqzsW/6MiXi0VagP
cukN0sIogXcxtRE7ap8mVj2Lz4IW1coQvphQ3xG5v42YEhZYivDCLjGi56b0Bkip
HdRxZF0tT0RY3z9BiZVeKXqm7vS2lu3bcLgpcHBwBKLkQKttJ+IIiEstwNqk5kOu
IDMxWlrepTWrxXNcb2CqhD2b8aB9nQLaLISlCJ9G5eWsDfQMhkct7QOZG/a0knJr
IfSeeyoBD1xXwlYzL+aJokU4A40P5PWDGtb+X2W9cgBjmmeA2yRwS6boP6K5x/Tr
k1lMN82xr4hZkDA//uSziU+8kg1YQGootDPeQec8hPmJL0c5LEEz0GBoghzLJlIr
qpK5v3HKZEmNiNbVfcu00IKSXYoC4ZsqRLInobC2/GzSDjxGJ7O6sCElxWtQoSFg
Hrkk+pw0ThYJoGJpUUzMwwfAwmr1TtiuF3ariho0jtHNbRoP3pvXp5zmvH1QO9+7
gTOyLytgqqw/SOd3Do1KEMTTWslCwtslDZkJ1xoTJ936MWUBnVvxmkN6yg0cL3LM
0n7YlE8HuwFnBfLtaRNVBY5pDvbX3Q520Ih9aBw5Db3FnfACXaapRoICk/0ICJAV
ezKHdwsb/E5qHEE9Yk3HsEWd/tntDfN83zTKaV0fNTLLXUc7W8IUXjNEmTZZN3hu
f1+RLjsxa6SlSzz1Bti4YQNNiYc2mEFLFFCNhqHh97lkEaEOSC4jqBFX16OmiCFo
f0N7h2lHwfzNd+aA49w2YRCLzccHuwMYVKSz94cUqod1EfzeDdA4FUWX06yJR9x9
nFw333UHk1Pj9ASyYehI9R1Q1Y14lfGjVAcE7t+EGa9vLX/kdwOUFLR++aY+7qvp
gUFD/rFqK7wXyEzT/3Ib6ASUuKL5Kj0/nS+T3f6ylr4n/T/L460IOftZLaRjXUcD
sH0n8ecL4YDxelBx2y/9UDUEplx2a546u/fRG1Mno20U+x0K2VzO2pfexBIhylms
YLLJExKNRCe9bc34w+RrW3oqM91RjK4Ngq+6d5pgV2FYLQHCNSbbqeBkKjJ9nX9D
xnSngoMznT0lmwbLgHBAKbVf5/OK98bGE5EyCsDd5gUKp/XkzOsCf0IxCeRqj46X
FN1GFFzdCh3emR4M6ZsTMe3+Xt481lS3E1/Qf9+eqmC/BU/5nFW54LkbnrdnLBSo
87NFtJ+thJZGIOUmZVfexWXQJ36YCM+/vO0bDPo05J+RYJDwHco0Z+32EUmi4ULX
PqH5rqSogTlONXIU3b+/9eGp/LxzpY+VXUspAovNgz6y8MsnOeLPWlivgmAiqJxn
37VtZP9wjSSwTbwzRq9L/6bH8uc+MbGfDK7fmYakKw6QDFWInITx00Yr2MVuo7Pe
vqdl6otM84Pgm/E0SRBDI/IP6WyWn0T2Yeox2DTc8jHwcjRB7tzRHCHU7+ypY34K
R+K0iDO8ZvmuCOUMnitYV7R8y+GLotRlPHIF7TjNq6SEe3o9G1v/IEM+zxMyRmDl
YzW7rqRM6zf+sWHVbwUZWkTb4alkgvTu39wW2PJKWkXPg1DJ3ib6xaygeQckmNlD
K4VjVnUBOBr0ph51VXZwqfPtAVXP1TmXBUIfYAXlgvdiiv0CLiC/xd1f5rePqKXh
X5bLTpBgEL2JS+tKqUcyuRBpaUTtn5SYTYO9DU5Fp0U1wy7G2Y3Y0dkGuQo2nfOF
p5gs3gA2igXjFBD4O/qzmS94n7guIgqFJ7ZhCKkdbgFVk3LcrbCDdSYhEWoZfyef
IMHSCfp7Idaqal+IUindwb+p8s8tzjGuY2EJkIDesoX6cO7Z7aX+oSTJLIyCCeyN
52fFjCpcEqfHXRoHiqNnDCp8d3w3JX5kPhvttAg6mA0/yPxCVqF+rPR+c/cFU1LP
aLRohnO0QInZIENo98GnEZpINdBzXIom4dNLrltpjgXz2VH1R9YAevffASA3O10x
6dfmOAu1Fa/k++/iC56yoOKw3a1io3809LiRpGRKWgPWibdI3wC1+q8Uw56gwU25
jwqTvOEbdHkOpykD2kXBPXpeosZR1UpTolREGzbH2ry6GxjVglmoDz2YJTLr/sNn
X2m3TZo+gfwblNeIfzUlstaPpUXHojrOsYGXPfZLZjUoux4YplBzjR+lsmYtTQQJ
BRQUEWW1As3cOBnNw9yVOYGTt7X7Zm/muXg0GNyByuVBEdcQrl+dRbLTfPQny1kH
Qu2VLTrYyhN6pfWV4b3FmGnhU6/Y6JV31malsFdn6cWtkmoNFahfR6bPCn/iynFP
ENcmpdHvp6SwRedrdk7FdXBry/9oq1T/AIeQsgjCxarrwwW5MlqhYxNxqbDZ4lv3
qBMR6fLIZhQiFlkdI2mbmy/zX0FJPvMAcVaj/kDS2pSeDEExuVXNxaAyyxJ+da8l
uRoFc80RPrtHxuJRcrx6Db+KH0JRxdyl3lBQCohUPKr4islPgoojAfiyPQsl5wa3
JTiBoXXAX4ZSilQ/0uiA+wp7skIh4FULKiSGwkFaeMignM8smqVSowgIUH08QmWW
NJW6UetE/x3rdb37AKCtqgyny3HcFFCxn6i5KFPv4iWPRC6PlqAdU6nD90iYiohL
f2qzcUY9JfKP2433JVCAwIaiK7WKri6qqIlUPw2ct4KewvzULvnmMUY2n0geSpJ6
PCNMBH8jk4iQBBdyGGluQykObYgzAMBuum+BLL9nUYK030W77iLu+5ylOyFTrosC
CxpfwoXw7jyNgzjH43j67cbvGAXjESMOpsdEGOVOpakYG35oooSEk0K/MNrbYQHt
ITZVPpkxJYqv0kAmkTXzK+iBt3hX2NxtdPGfgcgw34653u/lGhmUyOfgBGvfLVxh
Li1vHcTWkXXvAHWtsHcfKhcKUv03q6LWUl+Kmhq1Fvdzr9+juHyetYH0UdLN1Jm+
T8vej9uDp2/tRr5QVdCQ/Q+B9iOuGI6HDR7+10Ivdc+UDKjN8i2ejEzpugXsSvGm
cKZuz0HZWIHKZgrhR78c8PbBIgingiMdUQLLCl57YnSCsxkwmGy1/oCtZxvpY3zQ
rRA2Dnt1Xv+Pz/spbQSWyuyQowA+XtOmseRcYzbX41BbfBi2h2/PhBVeD8SfHPgE
77sULGASpWtcUuquKMCTp0ArMWXJ6WbJrZwPAS2cek3c7S+vTeGhgX929jpESM14
cSSnw4w0NVluGh3Gv2vE7IZG6y10CVp0jxetcpzjAtzcp1G02/zY8OjmahNBXXGe
GvajssXq0M0BHRvDtbPYv5YukEhpjdCA/A/GrWlAiMjXYkAO8t/8lkm4EDrjtzwE
ivnhKOX2s2HTyr+Ubz8CxbGXzyJTVqUlaRZxQtkaWa3qMRoXKp7fdUc+vNnp/4UT
ohAucKdWdxieFix0uJMeFZ4b0X5zZLOIefD237RPGH8xz7SJphbHj9GBnbWoy+8G
d1168jGW/ovrnUtuvTVc5fP9ogPU2MgeEjHCPFPeOuxbi0pwYxKp9i0XWuHBdZSq
4XPe3Et986fmhw+e1NHP0LD5CqWcNv3pLWStHV8baOj+yJH1sW5RbxoWID6vDrE2
nKtZAKhTchYLWDNVz490uRlysnaQhFgQmznhKfOwxURQy2gWsG7+0rJLUmMxoarK
uSPhAlkf/68rPFMKzNx7a9/ogrUJwWNrzbiNzT0BlPobk5nFka3MFE8MEMTUfvld
akO13jxMeb7AtBCFlS029z0QRHt5EIa+U5dUV2xjBTQdEgNJRMzOnuenF6vHvFty
m0ODcU2JC4ZbRmMWe367sQ5hi/+uFCiZUfmdWgUF5dD7/EhKS/E/SwPECI6JLiLy
AWxfeDbZgymz3sx2iuyFlKQMybyzYtZEeHVvZ7u4Uy8f9DQvoEJjUQv5GgyH9rLO
WWMcsKY/0a3ecXq/pWH2QTXL5ojaSa4GJHrcOBbKGyDj6CD6GUJ5Ai9jiIIGR3Nt
Ch0Xk732eHvHMVwUJIGoegbD5A7E5HKpVwXaIpFdzMUOjqS11bXhtYClPxeT502K
Duz+h6c/R7aLv0jqqkTgcIdGBWKTgO0ecPeXsANGDgPhoTtsX/0URYUBvmjGyKPF
9hHCmXKQMFw4znxMF61h/dp9g8AuDyQwldj65fnds6/j3UO6SzJl/sVFPMlcLw7w
sl/LOfADupVUIvkrED8DUBKbuT/urSZQ0yS/IeRgTJRmFEu6uRfeZghfLAUOdxmR
y1xOfk4E8ZOJY6pqRgzyCJ0ZU3aRJ9RItHnZc2HvNum0JK7+9t8mqU5+s55C0Bmx
ia20uCFls2JWns8KA65NHpsnfbUPvwF773mfG2YIJQ5Yg81aqFpILq9nn+IcNOLm
5+HVFVkEm13qzH4peJIG576GhYkLR9DiaEkcJBW2Qr3dsTA4WxgiYAU1A8S6bFUN
LXRDPzDyeq4tPPqxJ6ZXCVJTGfca/UvK8H8MPoSorfEZbqrhgRHi1FxJDDS+qAh1
GD0mgEaMqEWu2p1e/iMI8j4NVtzodlyQOP+dM4XR4KD0LTsP88GK/JJKvA9oBTlx
qj5Qsod7fXLvddloqyWyOah6toxKDg+DkOECMus1hLpOx+ktugoB9iK8bFLvAknW
oS9YZZZxeu3QZbNmchuVIvFxmBx4c70fbSnMJoRW+/lMl6jiD6dEmnQXckJ5mHCp
tJomHN0E2pDLvzB2gKAytHNZw4Dc4QAZlJVjwqKy8ZKcwX0xjwUoCMCrszZ1G0OB
sYnw0p360T1L7b8OxRFz9WkP1TP5uJb4Or3DeqGLReCegnLAZIXzLGJfI/ftQstB
iKb4e03NJbEOjIXMkg67g/xetj6TkjBOcARp97jgeKugIFfruzyEiU9uuEUTEWpK
DyAVNu67n53mEKwYDnDCjNRkHtwncdqeKVy5UwWMJ5oAytzA+iL27HzFuxgQ7JLO
5UNnK4CCbf/+P010hHEZTuJSPSWr6ifKZ8/lLMFm5jKJOnQ8/BV38p4EI9NZ8xdr
JjLXwRkb/hvrzZbIEqeqpJqfruB3MoeLSj6p74IZy26zqmMb7ms7WKXlX5Vfz6Oj
eyo0yvAWVCCczdYmBDNGDP3PnlIjKwFIjHtDzN2Dsn/CB1yvWX1p/CnFm98UQz33
6D1RPrFf/Tw1oCepbwSiItDOLrOnblQNGofsDmW/qzktungzb8eniHIJ52S0BT3N
pGwslB648/ivwOoPfZETo7VZg2w/noYHrIgwUZaK94b/wA7o6HERkAgSc7ZyH839
ePTo/DMXSH1E8w8w+FArelnrrLjfrf6mwn00hLxriyOkR90qe54nxvdBO/P90BBR
gUJF7/DAa0mHBWL1x8YZCeu5sRTpVIyYy21m88yaoBoxzfRq/FD2s+yOez2DYLlR
exs+k746zHCn5Ns+M0zytWQJZI1m+2XAgzyJjMrcIotJ0D4p5ip7ojPKLAqZEX/6
uc4IbKolyMXBxwnBsJ9mAblmcv+hDeIsHxvXIV8sbx70HH6YxrcaIKa4A5KHHJWV
vdGuKQDtoN6UMrr5qU0ANAbJ1H3SrvTtlxHMY3+zerjaFXEdguujnNKxQRkwe+Hn
8MpVNUYnpYWvFLbjVkN+mHQBOpc+EwR3a+Y2/bi3SRdszntDjmHAvfvSFwJvwQK2
Pm7uFCxt92PSTC85OSKrZo34cF/PxdgRQMwPUuIMbP0mD9LFmm54eq/W3h8zQ+d+
Ps47d/fpvWtTRXu0Dty9OoJU7aLvd9i0ZBC1wypGzerWHYhJbyqxaamalh3vOMEu
3gSAFh942oNBdr6hSP0Y/kxNhKs9g1Jt56Rian4yzPvsjdPwdeYhXN84kqA3/B1O
V36OTct3ynXCFxZhMuOxhKi1UBBX3rS5e/VVSvr8cCQWfTE1UAw2v1oYHuTgvJC0
0FajkPl0Pnzwrbckgm04ewGimhOtYuY/ym2Zg4ows27xSyu5w4Dojoo1wn4gk+A9
qZCP6jrd6W6+UGvJiKgrK6YtSnoal9lL4RcmRLMB3NNEklzmPRdUHGA+aVAsEGIg
5SEucwXr7hRdp25zsScXDpQClN4s/ePZW0PaD31YHi3ZFVqb+kNI/njUVkQ8WF4e
t1mFafEMKDYORrtK71dejbeAIA/l/kKEXxK6p9hlp54tUErdYORUxaE2BMjK/wSi
UVm9+ac6L9fvKB1jrhvc0Pemy9G51FcRHTABQ+g4lvE85rSCgcd7OTaL9IEKFaeB
jFmQowTH+w7aRcL1DDmcW0L2A278DRsa0+dWAJ4XjX0QXlVKVy/e+rA6DoG/J2iy
mKb90CF0u4N0zntfGRRPu/AhyhkZnkIgo8Rgw5cKDO2MxqYCBdMSks/7tIB0sdi3
3+9skyPT7TVUJ9Io9fJeF8HrROZqsSlNmq3EN3zHk7hrTpL7gxdlqKQArt+d6563
fhqjSnZLHlASDu472wcByNwyGtpCt281dZal1r79oWinAvgcnqqs6vEHLCE16nT/
misT+gkmp+4lc9yXPFtdicIKwbqVbpLl7gtEIEO5cMYU3mDeg2J8O+6ghMz+aeAF
GtGzmFLDagIdccY8uxb12x20xX2yNq0bRDW8LQ7LZAmgrGhSv+Cr1fNP4bwpnrlc
Oc2vYNjjQOwxhI66qUGLNpx6/omF4svspo8+r6qFKQePQ52+Lm7Nxxy3MhuX4tTU
U8wNPnpw8Txln1AtdWwDk8nGqWKybixeZH8f0rHvHoxV319R/6/lc/iC1TmtBEC0
yhppGGHszfVxylWAvKyQx/S6iIP5xTH1KnaWD/W83RT9ATilezHpvkELHUMvnmFk
jEFSq3s843pF9JqrKOIgAfK8S6/rjE2nW6EH6IBe5wOHeveoyVPMrAy+zk0JGhsJ
m1BRA5n9VxB5fiC4d1+YtD8bYQyVd/wd/5OVKRKAcCdvcUOw/I90FHiN898QlfMR
XJn3ObH0qYaNTBC63g95aDbQxq3MjDfRqZUnzkZxElNNFgIvFmOhseq1hA8CPUDT
3+H6SOFVmrGcd+wXnV2+M+c++oLJyVGBCXk0YsABalPPtIv5QmxwKr28ySO/3uF/
b+YkC5xUuItt9CeeYKO35PQSzkQZZDaGklyKzisli1K1ilg0Ay1JokEFRd42d7ty
EPDUuWkz95xr02nZgQNVdwzQcpJgP/uf0Bu2dD3RZ0XfbaVZia0VLhGafkFN/J2m
nDixp1PZ863ygCVcyQcJUsVXsUrA20abA41OMa3Nvu3pB1nueHtR8Agv8niiRaTg
yy168P0aAL6b3aXthgnJIoP2XABHH5tqRRoOCAzluWXjn5uXq5k9ScU9M+cJnN0R
qi/mcx4+gUz30NatS3tsJ9NXjIz122bd+PczQRgJNZGEsqvfOat1Jy6F8kB9MP6f
MSV/07NX6E99DNctRTyzZq8+7Cg+8mFDgROR7Pc798FB7k6S01CLEQO3cMQB5atG
/2CdBM4sZzMIk3+9RITdn6u0sRKgm7X4qyTYr4ljxsVGsmCaiof/oBQ6unpSWwM8
6f0iNqOQvo0pQyst1s2nKsZJM9FthVxywCVooV/6qelN3P5ANFR5ZJnKfk50zcPZ
rgnCZpOC7gW0lTLhmC9NY5CrvS66zPRSpHuBP1wGJJBCVDThl2zw8zNVMI982Rr+
dlx+3uNyDXOXuiL/WhCb0eIK68/UT9fXSms0ZNgJSHvghpW3CLOBV5ooaLTZesmM
X+9AhF9olPWtCCd+qn8G7u36qMtoRqpX+XGGzx2JQrwUnu9gSDzh5WWQDTfPDwue
bgz4jaWeLVBOttV/dbQ2VDyJVcLrKDBlkJVOcr5bFKFi2TsqoWDgJYqZyl/4mjvv
EVPkV5T2Z/qu8dO+TWrxO5TSs/nLowLiGX3TYO+cuZUZ/00sUvtK1MA938AupPbl
5E8GV5yXsyDABXIXVMt31iqK/EXGhu+d1zcaUtfrImuiWUXjyQktE58jhZ1TWeeO
MGyZWHPQXXOLbb/MZmz2MClYndeQrltB54i52jHB3KKewLfJWOGmau+zzjyl1uF5
1RYwySso/cv736ox/WHK6u6lQxQs+wHh72enTfb9Sg4TxwsWhZLgh8D7PZlQCpOU
k/6AFmSc73a7H0HyXeQPQ1o/aLdrIMW4nVeFH74hAWppGMUY+mGfPeoGJI13oLrX
KlqgK7MtNmbRo9C/D6+aDGh6B1fWbQ9YCVKFuV0ud41RkyKvTC2eJuILw+jD8O62
6Y3xiTVaC5QJUQE+4/lOFeVYMIwbhfQmNgmQSeqxbCzAxBRzDcGzfOSV6m4fbATF
9ajG58IiV2KHe73H5bFSQGIbmNpgbHHR7Ea33jvrMkgivLiq9dL8Wcf6kXuObcFJ
E0BEc+9z+wblcWKNql0s10O0YxiDzASEXLn9f8xW1cwle6T08bKbOED4mw/8dDiB
4gTiDDwq4EKaL+A63vOVI+EqfVgZhGy7HHY68hpQvd0Bm8/IqjLZzGC8vijhVoie
NwSiIpTPkSr0Nk8sbZ7cvkC5Lb3fZd94IvTixvGeLSWVGZiJ1qB9z9pRfaaKfLuy
Ezuz2a3fatgRCXdlxWGrlg2C+0mv447E8fxuOpHZl8FTm8O+XL5sQa0Oi+HQk75R
/NwoIXfdoBkvQtncccIJJhbKDRZAXNUp8VwQCg1ShFhZXmrF7eH8zhP0b93jK/cA
fczw0yLIDIe1oVaHd33XJPjCiNjcNSqSM+fjv01OHtadhyY6yp4HiHZyFd8Hj+Yj
Wmv2H2y5ptQEws2qVOwj/T0M5GE96fiHcUEyTcCeMU825Oa45vcwRSYHOlDqhO2w
oxLAdW78kjsaJaabn3jb9YABToHGSVrH9ZMV5jJw1V6AXDlFTCVvvHsNOqq7IbmP
j7YsYwFHhpUWyCo8sTLh5HHFQjflNOz8Y4NXJ0gmEW7L96YSoyDS4o6AxQHABzLb
tKvlw0CMDldCWy/CT0kp/8FhkrLxcCa6N4YwGpRWOZsIhlF74lUJiGRIREScGQBq
inN276106qoLXGKqvryzugn89/Ie0RnOR5xy7f2wEw4sqEiVpu/+NsSj0XP8sok2
NdJ9ouVRm8vUBJoi/m6bQk0oIr+75t2BMzbmdWEO9WL4EEYRaRPv4FnUxJuAmpP3
h5bhAOvb7ow244rXmVQyzjPazEhkUb9Z4O15+Q9AusFmO1PcPbA6KUg4HL+OHIQr
e7vnlXsAjoeixMeSVc1qcsEw1YmP2AvDrX1oN6OaJ0Q7DjOADW4AGSBzNvY9htre
4njbjlqt9mup+aK5ofBZPDYm1iwFx5EnG33k7ZoD3n9KC/BP2D0ts6v+uh6gY2dx
jn8Hc+suSt4bsp6ln24gwRtfnn3IbjiOBQlINtAlzWaPZJ/LD51fl95USgHYE8Wr
6HoxsfPbWVRCBmWUrVS6Tq/p6tU0/SrtBRgRiI2EfeDcVSn2Vkr8hyELJain+8mF
OZRRwgHQOgbVmLGnsRbnZVgrwKrMQRUVh0YUHfrs0Pjf8xVlQgfgEfI/DasoCHMV
ZwYgL5PVYKRZyOIxE/ByzBwfhkiPndMwlAB8z5FhRhDaXzE7XJFoVcDsSG6//zJJ
X6pgq2X/fq5kCf86CGiqZWdMh1J2PFkaMiGGp5bia+LrVDjwTfZ57zkRYlH4PbRO
uVVjahzh4Q1jQoeHMfytnAU7Njuu1nTteV4SaApmWBsa/j16leegkjBEU8k5Thgq
5I/TaGRDOnBB+MhTNlUhLtsuJokSuEeIThRC8YV/bChEAaxbz7LC0sC5uF0NpSUK
mcXu7PRwNx+XGN5vGF6lbRXwhZuoCWfB24mWtPH5dsZ4496PUbl4+Nc8LblPHjkh
4TC41SD/XHaml0cwWEcIes7dsWDcfmqly4Lc+/gBLDtfi4rF6ozKYubV06P7MDZ3
KqQQQVjQLE5lA3ErZMPpidUakT7GsgTSMeZLGscYWtXR0lVqvLfMCkapDXFwCRdC
uQIwQRJuK9r3IhqeA0tnb9CA1v3yAw705bTY/PxSPRyIdlCEzDP93s0Jmdq7dNPL
WbI+qRXlgR8nAutwZFt/UWEpZ9FszNx560ZYQXt63rLQKvUjxeNsAj4CDXXvuw9J
UqObgDYWS0VEt6O20usRpC48CrdGef0MpPWJOPuySqCVxXQIdEI5hJVqmnwXU8W8
jWQpw2bBWkb2YyH3x4RKaquygk/roX9xqIjyabqMcE7XZ98HHURepEl7Y/G/AGoF
HsRa+jRhUS/WqaBXFJobJqUysbdXaUtd0Y/OKHBF5HqMQSXtf67KQTqArkWCIIRO
wUsMN0vnGoFJ5CF5Th5SUWl6rTBkLU4ydg91UoZ4kvA8456GUX9xN8vzx+VcFCFN
K4f2efsQkpHK4UNPwX9gqxMHZ3ao7X3KS7GVLMoRTOXbem8i3Skap/jLZ7xecpS0
Mkl1/vvaDER2ucYMtJm/Q2SWYzn99O+GxA5BK+r8ZjBiUdk0fTNVBg4FrJapWmPn
DIWKQmLPv4sukjwrq+byz884geZ7UGE7Dkvp10bwqJvZbGBF8ZQTa2aIVyUPRFEd
5kCUC0DdCw5Lqt6iU2nKvC5hxkpJSIa3xI5K9w0E5J1e9saTPFm5PBAP3bvkRM59
LNre2hQv6682sH0U8tcpUdou7pZ9Anip9teSI5plKJYiPgEGR5AFd1klR95c8uTu
uR8BithXYteTHxuxZZDFOHm1OSr8mmyF1pDWlO5WsXHPPSEtcZ9o5H7hAF3af2ET
oWyy6CzLV8P1Dxj0285lGLva4Hj0BVwyJdASkW0KIasKCetczaMg8xXi/80cXmEa
Q0oBcLJDsdsyrPS/7hYt3nflKsZmf2j7uzbScvZIVQlw6Y4vFa+a3xU1GBNmroTq
CPOJlJtq1FKsQ0iTxXL8e2Iw45HQwlANvAG2LJslwNktOqwh7kfFbaLth05jRFJV
wiLugLTCZhVqN5rKwlDXVlzjm9edWPZeIJbefD9CscIYrlqjdHDLF/SnzaI7Ibhd
TYEUCBj9PjeQwZHDMEY2KKYpPhoGsFfj1rwoiwLkmsuv9yansHCBEImCQTJ1Bm9u
TVEL1TkElpey8cJgrepZIlvuuNJEpYrFIbE8LkMPonPMi3/vmsw+Jv6miBoGdmMV
sArVe4i/KRQdQxvlUvjrQo8rcb4kSfM/AfNW22wlDd7sDLevzjubET1L+hp5j2fZ
SoRxej1OLL7z2vE+1b6Luh1k+Z9UwTnBv7Tu0e5mJHqmNwPpUT0nRv2cEnidT7zg
SIVVemZrczrfQpT8thgR0FzNGjbbPzhXUin/MoJV6h1Z/tza8aQJXLL42O9EztxR
1omVEDXwtISP0QcWBGmcQEyUgzEfSl5xEk8iaeJLN8t/XQE2/pv49uF9TbzXQQFT
1JpAa0Nw+9dcCgknj4OMqCU6yXtMnRxvSHLAyVUpZUP81BKxd/0/6tVX7UKP7ruU
nAozQYfSNHKaArKrIgsMNRy0mi4QDK+uus9CtRhSZX01DcVaoiFmAYN+ssfK3AAj
fnAeaVaHmrhd7CQo0bS01xvqY0rvCX4F8dnB2wdl9yOzosAwW4FlrsQvOcjAOW4j
94X9iKsRCcvyMAKf3h2x0brT632J/7GUOvMS8go8kR/BKMJhHkTOh6mJOuV5BRHL
MWTvBhTC3mwRUXqNSgOQ57dEFGbD1t0asZrv8dl614qt1ZPZms9MgHYU9pMixmw7
teF29r6kGscauZhBRsToYKYT44Isx2SJGcFrQAgI7vikJJOF8eaDxmjlXc8D5VUf
468VWxoKZFco6swHuNGbBNNXC9nh4rDZw4qNfIiifRK9lr+UDm6rvOW+FnYEpFEZ
Mst5XfJYL+c//02pOxCv+AgtPnO58sjx3NKYrOujXcCr+2FQwQigHxSyXQaKO53Q
7uSRpATybmfZ/YpUJ367kSqtG0SJ53jvFMbj+YalC6ItmPshQ68MIcGcfotH5x+y
z4hV5frmYScfymmz0i+WzFnQKdvzjUxPDtcqei2PPzcVMcqQ6FYAA7sN1jAuDMoq
krFNv0Mu6XKm6iKBiocWNdBw3qISIrgM6+tiYqIQvpZqfgN5FDJfjJ9UzWJ6Z7e7
siyPt8vdhzXboC2Hkzo2rqngsZn1DNU8LxoJkwsfNN9sBwFYrfnKw0FjjMw2CznN
D+vOsDK4Z2CS6XLa1Q5BIisgnflqPhh57sVRuP5q0nIWeqoVp2qaioEDqTWiLp+3
vEF3+/2UYu/iaDdHpcKZXTpVxXNouMYdQNxhKn5w2ZFHPmqixb7A1HVzToF/o9FY
4IkDCZfSJNxcnMY2Mr83nSBwUj7vay+8ywLJYBNi9yfb2BaJUdUzW6ZlrotqwkDq
Cwk5EXblJB9zmQ8jtHNmWPw1b4D+lQC0s9MqeWzbkxN3sl5xlOgp+S7hdjP3KSBz
1ezdWuwg0UNm8y7aqEWyh8A1VgEr/pM3BRKRdL+wzxkDdcdJCulfz0ncQiO7x+5b
AMlH5nowng1Axhx0HVY6hD7ntU0MSL7DA0hvulALgDgY+fGBmOdxkDJpDfh0wPf3
yw3PA+qpATDdDAFD95JX9E+f5g/SS5nJf8016cMa943y4DDG2fAynAkVbTG6HnjP
KV1PsvLIDijQR6be0lUEkt6ZKLQEAX7scEZaxXL4Vq2OX40Bk8+51xnfxss4BsPn
dQd+htMOnjg4ddCnVD76m+GBRtJatSG3CoAVHM92LBi2oCbwaOeBABJnLomlNnKR
IcUT76CFqn6TSj+paRZpHRSzpPLAln6MSFSamYGnyyGFCE/aG39a+DZH1nFKh6J1
IKc5feIEdsHpnvKhINeaf+gTXhyTTfoNE347kmgkm6Xv2Yj8pBPz/OZcHJCT4HE9
M9g2frqW6Yim785xgHbjldXd/lzkbtyVuPR/OAZAc+KnsWmbBl/vhHeNMiJ2suiv
IoH8WBYMVSzPS2PkhNiwGe18kqLEu3emPy+iYjYfCLbYQn8VhMzXADl2OeE+aWAO
7ayzpsz2Qas3mxuhDhVuk+raEQAm0xF6LH9F7j+hes2FYplGs/bjs9+8dW2Dr+6e
3dS5ZCx+v7bQJ/1cpeo+qulDY6qb1dXgZrVELayJSbo2LnMMW4xnjPVz6PFJER9M
W5cCksO/TIP8Frac71SzpqF2NufxQ5chzg6VcIWnyT78iUPLKkQwGUzV9woj/sf9
PhaX7F/fyCmOLtFjhTGm0yoNciYUNZ/cidLbNaP5eGCEKNFC5oZzNOMo7LiTA0FJ
r3qP9F6JLY7qVeSloEpYKjqEy6JEX5h4v0hejsY/G2pEcmkwt0HbYXYgLvMg5Mrt
KhPqXUnXFrI4TzdY6DN1GRfqBDVLkQnPjQh4LK2qsYdRRL/Obx+XwUuWM7Zh7/UV
hhZAwGSKNm0WUwjq/r8o+HX9/F6S03G51OVDnlHZwgIl8G4gH2QBuczH3mlqV7I1
TXBDNxoe6f5Swoi/OCT8W6ebwqVxe+Gu4W35eIUk2VH/ev0nuGhRzHtihhIHvESi
WPXMOAEeoENtArxUlvy3ZPtSHeKe2QG0q9KVnoqA7TOT160f92sRmcgG7Pm9JgcY
80mKV4M8kZQUoetrZTNsvsmCS1stbwV28jPasw4RD341xBPGOf3icvEbVHHe9/d4
WobCQ7RQPtBHOOxUEjn2RAPsMZ0WoNNMtPNYQqaZm7TPejkTCSVV4GbGQI0oxQQL
0rHJOEZLRGnvUWGn1I80sREoJhkWCn53kh1nDZp52s5jE3BGIsS/h5qugSO0Pl1V
yBAIf0JxfPwzzC6RAb5QP8DGiU9o1HEMGH+vjhT54S3oAT1vtNGikyxDaF/Hmc3N
eI/PXodrx7b16JyACJC5zUaLUPp/ONYQoPuR1fujjgGKU7qq2d2NDZMyQTpHP8aw
tf6CUdS9c3GwEDWMAcAzIOA2ks3baQPTuZriAH8Rxya9zH1iAse/hDiyJW1FvmsV
x7zSF4066J4547NFerJeowfZHrfu21qeUErsl6rd/QnEsafFNcrwnN770+obxHVm
h+VhIf5xVAFceDjVSSVqKk8e3cXBzFH1XM2LxeYYHdXudCRKeSWzvjB7t/c45+D0
cNmFCOdrpCmH+m1OGJ4O6vFMOvqlqkRnT2oYgVxq7QSiFWeRQNDvQxJ2n+XZD6Ty
d+NTFTc3fO47YLhQFm/9I2gsON7aoAaXzsRYaVtGmWeiTuE7taPfKpGgHl3ILRMt
zzPxVltOn+I9a32TPa5jfn2d7u59asrl53WiYat+cCF2C+nz2ADVnyZBuTJgBSQ7
208l/noHHGC6NaXxTBuvvSCueqtB9woGpECodPAh7XZj+uqT3W6GrFFs019SLW1J
OroQ8pPhF9WaM+lWj9svBQWA7u5/yu4YQYYIbjAvcO1qoDWQmPn1vVeGAjIVIch8
LTm/sUmAXTPFJUOK4SvXuhFs+8nEUDlHhh8NSYeJexEEluicgK5qPNxSkEDOPWwv
vR7ji6t70Cya7jUJcv/HoOOQAIFHkP6wwgxdWv9wZxDIO6kxRHZdaHcYQoMmQnWp
Zh7W4/IsVmt0m7ItLDZw34C+dE6QTG1HrE79147+bWvOF3Pb0iskOUM76JVW3r3S
39K2T/egKStK0ukvl2Nch90HCNS+CWG5n2yoje2Bw5stbhPMlmafK87upGH7aI4f
UHS1B20U2cMOw5iZpYsY8SjmJa/+0qlyc/lQdyBEdXejTlN+WVPahoa+wq/dzq78
8ZcPJQZMnlPedcqG5m/37YlWBix2MmHF1p3+uZEO987e1MeM54uvWIeJOtHzdNen
fxmNAaWuaC3nyJ16buHTKzMCzulTFO/ds2ua5S6cKRgYX/9e7JLKO4MF00Y9G+cs
bTDjdCylbruIwvX5dSCAyQ+3uis8RzMPDYKuHmvKYRuA0hcpFQCJsaOEa+s9fkk3
bKsh/lxiMVGdef3aSPuJYGdjQzE+CiYrkja9T37GEAxoz65c1/R3rZUZYIQzUziw
avnrFsXWOM6YNI01UhXH4zpvnH8sUebOYouQwEx+dkfhGZdHmRGVub/Mh6nVRDI/
AHUQbGVZUPw9ExROoC97RZsXzIn7c6d154DDSpE5ihiiVsL+flBgpukUQxuX0sts
SiiSLOB0EgG/ar318rxXTr/iVsvvcNOsWrzGXoQUXY63pGbKO2+IUtj6kiAwC2oU
S79Ht8gnUuCtrfqKqLpSE17DimJaTyW314240Z7ryuO9tsz4ShToIuWB/WKLQTRS
OvjuYLNrGGOTcMvcp0V5lkqJBxQVvPdlr0KG2A+N1s/7iS+tGxqnGkrsTd9DmCU6
n/yEtgZdlzrzwna8djd79KumHxWIVyf8Ag+x82aCfFLaD/dDNp5AiA97H14f586t
A0qe1tBhkIYrEuq5LESLzwz1NxB2gi1OnizO8cf4JrY8QSU9tAUuzqZ3JO4TLZSa
jStg3ppleiu2Gk8wiQ8GFbvIGEYzSxJ8xVMaoLYj2VHl5qJynhCznciju/aNXnTx
tpAtQErc6oOyIu9yuvGiUPvrSJYuqk+q7Bi4QO8r86nzoFsIzSbe67jQF2pGtSnm
YPBMNw3k17MsOK93kc2Ivhzha81Xjl1ggUoegJOStkIDQ33H1Y+C0+/kTVQRP9fQ
iLX8Pk/5aAzDVqBW2x/RDwFRaflBQAYHUXNuvI6enFjV2SUzxfqq93T3tdswnzBJ
1LazuAzwOen0La7/u5GowYe7uvUgxlGQrvotD2LWKnYG8TqSC53kpjeGG72aY6h9
tLlc0Ojg2Qg6nsoZO12LISERcRhN8M/Rp5vbj5pwHl2xaayxJMYr2v/xO7D5AclD
4hIBrCnk6SZUbRBkUZ3YjAhHNsIotZ7L/mtRaUQYFQ367Ifk+kvgbyEf7+dmcwla
RkOTSKpBvPYLfWn84GEIJMmZUBsVn5Z7qVDcCy+Iqy3HAgxknF64UOcs3nmiDKik
/ypw7hZw3bdhAIPajSHITsDFtRt2Ce8w1EeXcEh2H9w5MIijXM0jgTLSIM3zMh9x
gnYOxY19N+2bO0M8Td6JGwL+bGGDWspw3nKJLF16X0VjfI3LISUGO+KMhfrYUAj5
a9mo9c5Ev8xOtDeST2rPxU7oGpVmNMSzMvBnEYlAl11UoYQJp9mV5MQjiBZhpHpJ
6kLpqwJ/pw4Rc9tyGxIXcisccapmBZBgo0fkx5QpVsAukajmotj+7oKaKzhZVnH7
z3V1lwAyjJMATcxBHykomQzNE7rR90Ujcr/NDtxLqsgp+z+KZ8Ty3TtiW9DDQeLR
z2WlB3tXEG7a3FaTSZgi5gFFA1xIMm7BbaZ+LIythtUH4PFUH5k73lPLUc2hkwBc
R4gef2pouTq5iFVbXfC/0plfXsP5F9BapyiSoDjNBoGrUvyP6jWXFEkzAr+w6SKw
JoCOIHntei/3sDbyWCy1XTAAlimU9AI0uWPJgQcIDNX+5WSIL6+8NY4lNZvXR0OU
TjV1Ww/eMu1DU8oVzRrjtpZ8A7SKWinB8x9kAkS/7BvFnGxJ5q8fCQyvyMl2/4Yt
skAOnMeAUw/DyTIZQDIWLsQwJrYAUxLK12s5gSwg26AZ6Y1BAGy0GBSRXnrJQZ39
6GYSlrWSRSXf3cZ53yIiNafBWiKBf5uWhGAWd00W+TtbW7ko2y3lEBpevV6rE9SG
KCnENhkQkjDLH/Du1tHVfzIHJfQa++tAXhJ3I3ZIDYDK15dnhCOPI6LethDYQP/x
JrN8siUqQmB4JJpQZGeVnSTboqqgHQMIIz2sItqfajYv2rZcf97ykVbu+JHWl3vl
CGDiy58WiD1GnhL4nrFVRFhhk1Jh/IpHheGGQJ+CxjZMPQ99XcNYX3E7GyrZqCSd
IER0UW65tveTY0hALs8Yme03My8wjbybzXohENUT7WSdzM5NrrK8RUFrST3IFrdp
zcACpAG3gzZFmeiOodYUn96oYdrprDOzTVChCJcfcaCERWfjcwhvRYuc2ot+k/Mc
IPHEneFxZ97LqYbiiz+jHukH85XNNT1ERr+5QwSJ/HL7GrJNpP9X1BhZgRv8P6yt
lNf1+786TI8meQI7THA3xBNeIuI1JBWQ4pnkfyXcLzgiINWXSZ+F17rsk2y+Ft3f
9Gr0A/hzWU9I1wNP/5v+fem/YpVIjGa9Jhn9M64cZSVTzcg8HxyBYvRvtCkJa0kq
YOYYjL3xK9Lo0Rc2efB/TF/c5nc5cQfE9idIa0j7VGgcm69C4EYsgaLPWRNLA+iK
a3GacK25+Hgv3ymrWSkpLeHQHPI3lpZ2Dt72Mn5oRW8v/qRgTEpzWNUBXIghYVhf
KrOLk3GMkEQ90zzeBq2OYSzf7EOXVAgWCRuHa8n14CPVV6Mk0djcYOZfeWVVQ4AU
zAX+HBcRZbxLXJ3K5CRMe0zOEsJTNr2o4oJDDS+qTsbmNghLMxpZ49K3Zw4v4IJP
9pc8bg/xzfM8Ge9YgobvcNp49dxem+ncpV0L0ca+KlgHFhAsf597U4Q5kjA8Jhyq
elp3OOdXOxqPuQTxoRPfxulirHweS6XSoIjuslmkqBbFPEcjIKvyF2dftWzKtPGy
YNBLqmPEdXnDv/uTlnKcs5Y4XD8RIny6XCJ7LsUkIMaAHedzY4ATz06VcYk8aeCp
IAjb8a1raYlycXwzcBoxABgDS6VKQNsXnqyO29vTOl1//CWoNTC+WINjSNq0nXrG
pet1wWPcVcVs1F23oMo/MmKZSy2IZaTB5KIdxaPrKPUdiTSMtFqiae0mi/HYEqI1
x5ovjscEm2d8QWmWM0GdaImd827DnkpzlBMYW+Wliz1XHBwCieqEFGqKyww6e8Op
mSzp6JRBBKUsEToJprhhKNOybVALeO3vXbvxIJ+omiCJ89Usgwf9YSTm8quSBRhL
EqwgzFHFQQe+gXgMAT3y780QOVYoNZzjIJLA9+24GCUL7xJ/mNl83SHKJ/wN+vUg
QXeowu89AVndcXCaaKqvJsOzYVWAvdGA7zrbMcUqFA8VL5nmBAxrG/qbZQ3tCsO0
SZ9Mu+Qgt3TZshq2YIlUdfN/Yw/KwDF+9KnM9QChqX1irUlO42u0p1rf9hq62u6P
ZQX/JjjG+UYdKWg9Q6eYqVf6xYnKcdUTlUyP8oNN14EclZLebBzzq4xOM3Cuus5T
uZ01Ll68xU3MVwsdanopS9djrqHrSGqgfAV70+gOxE/c18knf0li688Q8EYWNhtp
5syoyFifodZEh5APsJAvkDIt0aSmtKJHuDgGaSwi/cuax8sn9/J2sM0URsOGEKED
V91345JXB5tkK1DQPcAakIBzlm9bQAaBq8/xwa5jpo072MSJ5bWPf+BorSOxpbDS
CUhWVJ3jzJ8z/eN5cMYJSSMWuIKcAHsg9Cwp6xeH4l9/D+VxQnn/jVxlhqpDXMWU
J0FbSAwAkl75Gfp3reoBKaIYlCy6tpEwv+ekcEDcerjsVMsSBkdI22BjMae7e5z6
j2R/l8NCavFuxwOJTGEY3LKIs+1JsP0MlOfyHf1zKyGKCA4ZF+lJ3EzxMg3e5+ti
gugA7IddOE9rHhTNHYCFxkwEnE1hy4wwzJKC4WOm+twwSV/kU9coIH7voYH6W/M2
w81hNbAYUXFH+EA6C3LPLw1id48tisDHIB9X2u0liFxNyrEHTw9ZpSND84IqFnCo
a3gFLBGlI5HoAVzzcesSV1LiVea/O5j99goLK5vu1mWccTuQ89Am87lrAPr93atc
e4Xll6FBzGBdg0MRiAuRyG0+TD9AjWolFpYLfWeefuZlRbiSrj61RxsHlwr9NqiO
cowWBsOtvCaVb2DjHrl58lRfyLDNmLOqY2q0NLPx5EI7wBMqUHPiF5TdRYVgu7LA
/ovHyNXVfUryFI9g/JfOsGuSp/cgj2omJ78T9wbpMJttDV4Xcu7L6CfMEUpzpMO6
kW5ZwvE6O1qoxrIyt5KWYJtJJjeuINHB8eY6lZdi8n6ZIvFnSUPH94q446PLPndC
tl0h5XoO2tONJDn+4mQCIzR8H8PzNDS4zZbsk2q/9GFFf5/lGiSaqBV3y4fT9RCx
865WEOhpYyDzitwEP+ITEJH+lPKtWyB2Uk0Ez1HVYR5BEsesYq5cp88X62v35n6K
CqncW70IxEOtON2CgUr2NIKTv/PdJLXkJG+/BdnWMnU3978OSfRxdOTde0yButeB
zWO7Vxgz7EB86uCzNKeJSXoIKsUJEjI2K52LhN+tvPTppHK8Y9+6rpHQPHxZDGfk
8PZnXJtnv01QWdgI0OFG/JndLhQqTJvwIudtxADYOXI5ar6DJcJcg2SWdf/lJcNm
E1x9RCJSZGzJXD/TIh5XwIx/xeH5IjcRON3z8XlpqKurNTzzlvwZh4QD47h8g1Se
fD6WUsRiPmApq4We9/xQllyMyviQmWayQe8LKrrLDTc3W4RWB42HFSrWue2/Ln6N
uDM4np56UnqQD/+PkO/DGgXry8H0b3WV7p1AV4n69cdDZeGQKAjXq7+DCoNKqFzo
m+Hlphk77C2m7LHVQbPHe4BN7qBKfqs+9ofIb9nIX67D6J7X4FdLuBLdrpoJZgNF
5Ktlbb/vKzTz5GDSKyBMUYyjHGTVuAJn00G8EtCJtn+IADwnPbtUYGM97a4HQMxq
JfWHIF1mB296Mvs9zKJmeiKBVnnJYfybnzDFL1fEVt7+CY2/EyfLomL+qvTeAWrB
ZztxJYQV9lYkw9rLRbuJ6oENa+2rsm9SoV+mfvITZZGW5PBDuBn46qX6J3SOunqQ
o7Q67uhK5DYJc86lU96Jeu3dbikNJyO8s0C8R2y/+UaIg15NvHapigAQRWXeXCjV
N1j+XPQYlPeTA7g/Qxv+szXnSKt0tRnfNe84Kdt4InvR3q6uLkK4T4+GSWSM2NjR
HjxY0CVZQ+QZv3v1nwseVBpet+mkDebsVYYl2ZF7HpoVbj7NclyPXhEKsHg27/sf
uhvNMdChNnG+7/RWnCA39uwX/1ZPrllUUmRWIRjOEfSPX4n+Ll7ZCrACoMQVwF7y
pkK0+zAvjiTxszUpzEVUcT6R/lN1tsDd3Y0HtW/sPF5P4A1uwY6gVsYks24Nhc7C
S9fPL4Uw2HhzglGNM04R7V3fezVjhAbFOc5zrIaqUe7Kir/V2LS7+G7LvIFVdfxL
DXKAtL24EWaAZ1l67l98Heg8bNSgXd+W9AXtqDpwkug/btqExdZPhQZ3rkNOtbbZ
ZAq8vq9cG/BYVF0vgnk64/EXu7Q10MYRgW+dkuCJToVdS1CbxradW69fcZPJom8N
cCyH6LbvDPzTO+LGCQloxTfvyxtc6MpJhYtO5vRLx3/I+YiX8PB1bAiJtrneda8i
68UN9w9iKPKNQhtdFidD3VpS8hd6z/G7pmLvHSKIN/kHsxanjxCzJVAKTFUl6P1H
TRq7+/ntmzNbnG8mct3coyMz8x3w+1UXyjnpkIbXvanpVULKA1cBsI82xce9Rxl9
YwofKytGOxl5SBorqc67j34XHy82HftX5xHtlpYFg0khZ+3st2tkN25jrywVHZFZ
9RYm5f5IvQ3+aFJv+zu7Jj0UAYdMGBX2fpCQaieqBlwYfNnokv50McujBk5YYPRf
7uEx0wXGPcgUnnIF2zucCLeiVDnIJZZVh/j+Tbk3xsA41oYg5t1HPXRtB5DNDZDd
/oahnWPoFQ0V4Xg9a1g2DSanHGDoOydnzjPj2M65PEBmb/9VKCUX/cW3YJJF9Iqz
q1HGSJG9FSVi7FSehjznL+vJA6WR9DsBkJ6TOaZPqC1QkIDMM1tzPB5x1vMYsnha
pV9dPU9j6eeLni4Ay3lzvLlO7QsjoyxL0hGBgrwuk+rCnREzZNO4F31NNdHnUof7
htl1uVhF/4jx6Yy80NsNuHfAHeTJL9zXkglGM8jb256lDhylTiAuZXVkptfdhmmX
iLkCYIhl4I/Ee2bYIVr8e04KaeWbE5y0wW4JSRNuSYdiQv6jbI3gnVBdzlES90I0
uxMPRgsx3Exp1M4OzSpeoE7NPdApVEAsgOHGDmc2zlF57+PCLd5qijXk9eCwD/DK
aLpRxmzfQRQTFa5gj8bpz/Mr9b2JXnGk6EE/r1/gcFmvCmdpHyG7XM/hXXvKbcNa
Lkzb8ZGj1C1b4uhDklzN3QuXf+C4uosiNoEgZEImNw3RSPQhWOCO2lJ2FnfRBMnH
f8xz93BpeXJe46t3xhGCaxU+MPb7MQIw+sEd2ygJHJo=
`protect END_PROTECTED
