`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNaQEYxvPprFi9JfCa24KI2iHum6sG1TZA9BqFCf/KdriQEgUbG4h8FeFW7uxhtU
0RUUznVK/n8lY+WZFnI1ug0bczaCXEBotI5zEmBMoIjZh/3eKriXtwDpoHTeRjpf
GyztzJr/4XIqBr+BMPHp3QWjdFp3EA9fydCFLXQXdWil6PQ8+n/+cEaxq7uN8u/m
j0MTDerf+/ISh0u1t4iTbWu/aCsRBiOCZv0CiCl1xX2ZviZM7/Mxlu728g+nA99f
cfPAqzaL2dlKzGeAm0O3e+DihF3Y0tou2+2UOugl3CqlV6+zQAYIpp80GkuCjofr
Wx2cDNFFqt0Fkt41kV86/QBp6Ueut+7/JrATBdtUtSmt9SFRpAOfs0IHmox4xXCB
6VMef8m0hajLy3XN2nkpXS+kuVdVjVZYfz3zqXeWc983AtaF4AD4EWZNikw1NPNI
IYd8/in91MqifbFDRoPzQRR+kbFXAH3Sz0kRrPtaNcksvTIXPG48cCCrqb7JjXx8
X+xVv4NeTqna+6ONXd4zkK/jGfPOzLEYwYbahZ6l4FMRGZJO+PlA6ETddQ1y6d63
E094vGH/Ju1nyOBCTWWuXZAKFeif/opbWxdl0RT9P7EtLvosAnB+ux4aYWxBosK2
ML5sHvP7ZyMdNxpHh1O0WLb63WEIbuUPSn5bgpNYV7nvA/vb5BOIW8NdrdijF753
nBgtfDZwVMQP2i8etKGK+vQ4ZYfgAq+5EOvbR8GNg4LNTKtqoL9lT1k0mFCtzeaN
T1wg8GVQq7H+eoMZkFYSXfI9c+/gmzpsH2K+OwDn6miBInI1UGimR67no4BkScOG
`protect END_PROTECTED
