`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vA5zKSlcIcFgNPr7qQ4Fxj0naRX1Co65jl6V7nB+TgIHBMgZi0YQvaZwtkp42HYW
ofChXeoYTmLMJkb8NFICbvOjagevUxVtUj8ehbqOe7JF89gaSNIVhUG7igqYAkMj
knHS9YlvmBqGc2jmIYq+MNqN51OgMUmDfhskaq75zvRxW4nQt9fPmdDm2XIv0WR9
oO/11fujKW8C9vLHf3gTwJMsULKOpMM/yMTVqyQmxARMdFja9T5fWE+8REhABZS9
j/JcAieFKOa66C3jRhtTtBL531M16FQp1jdIM8mFrJK8Lwp6apPGWrVTf2YEkauE
kA4XQZFKD/S5W+EqZ976ntVsWT+DVreKV+z9oZLb8Oas+DPCbXDq1jPxaJHHCL29
KgeNPfh7dgjK9jDA6/Zetc9VsWYSn8ZWjtghwfca+WjtwM2w+GDnlrkltf9hB5Bb
JhTcnwPqMx/+Cvb4vmm7DEy3PT/KYFm4qMvthlEFbS3EoRmCeT5/7ZYLdHde2vH7
28rTHiAaPNKaazud9wpkM3qcf4V8VQbE1Fnd2iOQk/gY+4SIbzX3UmTj1w9yT1Ln
rBsrPNo851sX/4yPs+zQJ6ZItKMvHltkOTK7dv6b5/kBppFlwwDjNE3XW0X5Vfw2
dqjRmpY5IRKXdc7kgPJWbJ6yr8wqkVhWeroQ5rEudic+sS7IIgdl5/WjhTCnR4Ro
73uSTgssuH/un8KAPW8p9bixKC/Xl6Mambk/aJ1uCkbT9Y/ipARzgC/w1EE1beAm
e+8YSNosJbucJ4ANK3gVLvw43ymqX/u4RRKdoMWimpmjpPSYr71k3BF8DK6ZfXhJ
jHgV71fHbniP1LQFM1GwB2sxwkOXGLsqoAq8YaWWlT2ZftasYYX/rDseE1mJ7236
5XNGpyysxaPDmeEBEJMHjmSD9Ej81qR63HR4NV+gnE1F7gDZTex4qekv5M2fnXON
3lvb5DepMArklczluC5aeRR9/d39onoRyVrbt8ZNJJlWE+AwP9kuDrEo2RtHm1im
mcYwYuT/OtZjrVVKEVWAmz9XkbVa8g5F9UnrqxZpvIVoDt6n+AeVzIz2EvM0lcRU
+Y/8Wj/IEad7VA8Sc8XpL3FzeEpwagNMYeiaMRrEeHGZGp1XysyIfW0ojCr2gIlo
Lpr60B7Dt4UGplW2wd5N403jRX2G+C0pdatfUfemd17CV++KC1sTwS3YcRYSL3Yz
aqKiMoRYHd2prRKxKa1YdbgUX0GKTMQCVOJJ2+lX7QOEsJDiNKwLO+pmS+4zC0Cy
f1Rie4CxF1x0M/ltzuUgKV8SffmlrW7pjFpgouC7IhQZfnDLSr61KckWi2ZjOvB8
weJ4Fbvcu5xZq6j50tHaXjxXCnw0M9usMHw1XyEYS7b7JQs1qPnk43DUnIgCFdP9
lFsn8cjHYsOcmHqDg7GOfRM4fsdtqmEHPLi3CN8nOaxYDFoW4GiSo8fY1sKlZ5eZ
h1DRT0VCXgqY+WLADiiTqvr27lDjJtPeBj/ZVPD6z71rrrSS3rpq5iR6g0qYUR6p
yDPFkJuIGHQvb4lR7pIcP/N3yLLWXz3G+8NGmMocvsXFjQurVFbtsJgEoeAbu1ew
9vp5t0SwJNxhi+A0M3u2BvNbXsLWUNM3l8fLJUHmWAlweepa3HzvWJ16r0i6obhO
BlvliPsbLHF4XHwczvKnQQ8q/IJgYJYRtnkHkxxG8HVkPERglSSbAbjGsfN7QaH5
pthYklbASobdEV0b21J96LfL7GBQ9UXvWzqtUnncC6XeTXh0D/EaLpBK5tqyeE8G
rHJWPlrD6JfckjcuAo1Y3hPtkkdt0G4An4AlX6FICR8qofwHtyJiKGCFwXx12MG8
zxKpIfxVUxoSVLgEe1JoYm7OcnFS9r45AkFPRuJPGG0q3lxvDcmh6RdxRfbBuYQi
k4IiACEsj4awQ1Ws7fbNAQKWWcJutoJLfbELc1ygOuESlsRi/SJpJxD9OiKwAVHr
c7gCPumlzEWW/MGFuQ1oGY3cGiYFVn5HpCqNtDoyhr/haQDER3laknIZbeWDpuPK
y/K4CUgnUQvcWAittH19WomH0I5wy6zzTG2UI29SBeCRcu1UkHVFcho1PzzPbzSd
hu0e+Q0ME3ElNDPvs9ICXrmUd7sdxuiZ4nfVw6MOgZ5lEZo93v9kjRI5B5V0+bvE
62hR6NCBz8oY0RarOz/ETcLbJ2mOVX0xxuvvu32hYbfzF4ixU8flphLAI5f5f1X7
4Yk5aX4IIbl68Xah/c+/oo6vcDkF+gic4ww4G1d8YMksPP0mhul9xWK8lT4CHsdl
2aLPjfuyFUj07J5uckxmSr4/KwOJ042WpslQoDrE1MFltSx9uGueJv8lv431+BQD
igAR8f279tAbfyK9KH9J7xxVQl+lx0cKPX/h22Mx8ea7KqQ2VycfAJ4OMTrPkf16
`protect END_PROTECTED
