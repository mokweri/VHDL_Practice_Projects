`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+MLqEN5KOglJE4dgnmT/B7iS7SX8k7umvn2Qpb9DRzS+Zr9H4ahExc7auSdNfIH
TEXGT5sM6/S1esfttmyiVnRxNnk4XzCV6t5J/gGkvQwL8gWyInxxnbA5Z5si+YgG
7A2G3dFKGoWB8raSg0II6ijj9vcyHq1uJVNZKCtaGMeBn3Zs9mbksyElFK/z6u45
WZUhztPUChiee1jLLHVbXeV0M1XxzMH/Puw9cSqWrqs9W518CoaNWsUpl5kNn1RA
5jVJATInIAS4I6n61nq/JfRvQ+eAQiaQWYMBrHwOu+HEv+WwDf0l4ZCM2jK4nY3/
nbhRV9oQvic+Ek0xBfYkMtvlkV8o+B3MWZN8VrF+nCJC6SWuqc8syeeAm7vTZj9W
V8M14QVLr405vlhh5coRftWRmI6anSMgaLSthQq/Cg+Jsfj90hHz86xuru2qhct6
K6RVuKmcFln+C9/1AoFInlSlkt2UsRcKmfABr1HsYec7yEFJfdg4VlrQ8wq+anXo
CXe47bp16DqFwLFQB8sKXAC3tbK0tVAQlQW/lbS6oK1xgUGkhOl/CfgbhRSsmKpr
Jz54NlLR9nzmN3z6ivmPzKijW30iv3gH1dFWBFwE0quPGq6PVmamMFw34M++lDRm
Yc4TSGl6TGml3D4z7JeJve5Jlp05yb7+NxHO2IawzN/R8zz7apmFzjuuoEuRAYxK
wwzcCiODDwyg+q2hmX7ffCypBcOWH+q4JSM/EIrZe4FqBb+m1mnAWXeLDZVyvRtV
FuIMX0Fok0XzzC/yHTrnoio0EYjfmhbRc6hUJ2n53AGYFryUWPLAgL/NbSjPCPJh
sYznJJvMR4AcdsN2JrB5kpSEqIV4w9JjTcaQOvrYCO2KHuGEhV4uNOoJkLYrRjzV
b2fMqm1OFkFKSnI0dBqkXwJC66R73aJMUfre2NqiH0i27BpgBxaciD1JLxBmyffA
8kY2QwOxbDynXfokz89/btXN+72vMwvhbC6JKdRRbbvAtJN1nGOZmRR3wlFixeEN
fxvqsyBNg5NfCsnwKSTXX2xuQIWG2MOYBtakXWT6TOIahDf9k1diu82kus/8RMQl
rpZCLtMHZoK/8t6HSLKMiHKVArYWWpLONrZ6JHIyUITx5ePPzO9QET9A+3n8ed2C
ThwfW7RrNeYoA6KemWxzF+EKZlKioDDE6/Nnk1JyOETu0Lr32hRnej2LZrewbliH
pIwzXJBOj/DXXFGaUcOT1kpCSUBrYSkXIm3wIYJD8qcSuYnpFkezDjYOPbwC+q0m
ybtQehZD/4w8QeRQYFmrtwjujnRWrXFkGUzOWmT1mrOwmV5hI/GSPtf3oMjtVvKO
PYJDOmsQVaz7Bip7Udiv9EVHwCNvvlmWYJG5YGnbFuuUS96Q+0lBR5fTcHq8Ppsh
OapuMKj0BEjA47AuTRpLQagO7f4gpLcNwnn3/9oMGoejVMzjp7GQ4Qhq72+bDmYC
yEdLdb3dWUoZSsKrUkAZIDs0qAISzkvcipucF/Jb9DvP48RSeY//bMbYHaQ0kLSs
uUyrPD5WGNvkFz+vlHKfN0g2ROmjpIhgeMDUkmWeW5nJdFqFLV920vNIYLgsagP6
2T3x/c+vzdgUZA/2GWG7WMEc8D0ijTEWT3FFBIRjK4kaHGOLnuSv4mTuyXMsJn7a
4KqGOzqcYkcsNw+ihyKPHXZ7mb6Mo28YqApPiCoJ/wIIPpcDLA+nCx+Ap1HKFb++
6HH2hbViCIy5eQaeRobE9teerLLDYnVLo22HQM3751P2Gf66lqwJKCNGFgS7Eixb
zflfqnPbt7stbEcfZVqKpRQ5E0B+Yf6I3uyoG/p3fEE7YtXUSRNjyvSlSqUMUMMU
+FXBt76pzWK0aQZmqFxf7TC5k3TSfIDENxmsxuDAklTWV2jPZ97dJxd9+9oi7wSt
oAzIArX8ikkK4Yq61gWO7mIRtrIzsWvNpDXRyjpmhrJ4JMB7pK3NbEY+v/JazW2s
Unflx/yndGo8f1W6F6/+KPCnF2Xcg/eU5zmbM7Ihu2wad2GqJYoJcqywlvUwqTGl
q8VQWRgm0PccsquDpszDMX3uBD3IEg0fsR9POm0opBzTnR+fFHdGy1JT3afqDvi5
heyKr+EuKY8aK5UfCqDMzFygFHpCRl+g+w1uQfYzUJGIV29YydF1MoAT2vtQUe0I
KOA251IVDaJOsbEaUFJn6NTFpq5u0W5Paetu4taIEOP0x05qHQZ7CznTtIQfxG6f
GgytRkr1jD/ZSJqDeoRXqNB+DrHkkRU/c1JbyVd0MLkemCX4VD+t2M5ueuWDuwMI
bmohJOVMWF+8PhgxokC4MLA/JKE7oesw5D38VwAk63ytXtIzuc2CHovxSHI1q+q5
guK6OPSvgNEEMi4/3Kn6xF+PF9u40fvEGuiNDIzwb1OrJxTO6/bzJgF8I9PvOyxo
emAMCi4v96hrWJhQJH9+ORpL0VaPVuWxLqAEQvUVVLycbrtf2ubEn67d24cmK2hU
M2YQcRF4fCgSWvEvhcoCd8WpzUEiq8WJzBlovibQgvpws/zpzEinoYLD3keQDTL5
7+fw63R2STo/gnLuvMCUvlWBfwJUl85Ycf5p7xGgWwPbs3Gh86eCvBPxq9nTgbma
wKGFkkweb7aPWyFJ9r2uCxHklSj08aZwXHibk9SAslu+oKi2pO2awhbrThHgMegP
nN6mfY8rCoMJgOq597yelVrbLqUHgaG+Gg4cNwg9wn8MxNs2jJ3HAK27CjjHbFBv
rRZRahmgvJTCp1aBV2DVggPhOmL5FOtTdz1hvJD66PoSg0Tkv8FdNFInfc8G0+e4
Mnq1ECnxXvpnLehhi3MhU7PH2oGJChaS79EDKdL9ShDdywIYDaKx8LAWLxsf6Z0U
kjzDtU5Z1/0cfiqyO3CRXw20QQVx7uOj83dPGV903FLuudICrxfelkMD2/Wk0Mk7
4YtTqcWW06SpYh0/cForADbtNXYOmZ5htsX0FXeEa5GnMKX+5ZVUHXwx32R5pH8K
p8GrPBm9mA9eRS1HCJSesFbjCbvIlqeQaHGqCmv5HS22yuJS292V+On1cu45Xpj4
YC9qvxNaRGy7OAYy6ofLzQJWVFNfrKXzJmgjMuVKuF7bERzqoJVSF+cjx0ei4gV6
qxTOFMzmxRx7yzB+p5wy+I5OI0d3s/OsOtJmz2BwqLai3/bPforuZkoTvLu9XA4U
slwSiOhGduxzA/af0+DAaWiwONZ4ZzG1qeQvHuhKn/f4ymtwd+GS9CFUnEaVANnn
iU9H/hJ74Q81Q6iOnI0uKgrCr9ehNmBiJ8ROKL4kEktj3IugwThFisiqUPVmHEa0
6EsqujZxivJiMZhQgntR0DssYzP3kVOmPTBBE3YaeQ/Al70ccx59BagD13pi+cef
MsR7hEBlUIdHKGB+Tph3owaCUaSo2Z4+gEcz3zS/v6J59RdYjAKi6IvFYgOFQ239
ilOc3W/GI38qSkBjDs030CFE+VciupgzwCuDnRLBbJTvk2tKIoCi5BpL0oxYwMxP
AaMpCQxoOuf2xivPCSN48K0Wp1lnnYGjFR8CWOqSP2wxVJmmmqYvN1KYf80Dyuzc
DXJDjTvN2dqXD+ukftIQQimjOJo9psli13IZdmJt1tJTuplV6nJoVT2HQX3u4MlG
cwTdchclL/nCf25CEDEQEgGZfTT6UqRBMUorJKtqbCJkNCVEc+9Vcejx80dhWR/v
6EMRwHQWrdIuGeVohcFywbByzWmG7E3mrX2Euc8a00JB0N7FX+DegBfWdBs/NLVf
Pb0Z/I9WGtPswrKYTVz96rkqgPyjsHhQWXoZyD0bY1/LQ3VODN3ohVVr20fpSWlv
fMZIPj+QKMQHz9mDFaj6qI1B23UcfMB9f/fv5kUGelZaIAfBg7Jjj3wbCMl5IvBp
u37Ty5k7KLd5PEPtZslw49CvyJtkCyDqWuPF6uD0ZHqXcZKO9y7djateSzbUzhgn
5RElNRoWSnztHEh/ZC1mO3lbwZtlerz/B6e8Rup17tTfZIORn5tCB7nOm7Dy6ECA
Uvp58JYYs2+edMo5l/Qax/EUUFCmGpV0TyYwhb4YKXiidurwNFum8zLtEbrhiL1O
MCnyu3VDcwlAa9zyT6NGLli4/pAJViFhGQzk7hQOHNGQd7FzDDBAwU8qtT6XCH5F
FlCchRGULs4LIL0QjKxJhw2yhpOb/h+FRqC3s8pY+xQc9UVr35E8/LjQ7XSj+Gpq
ZeppKyivGXLOeL2Q/TSoDB318hzvRwRKCCe7k4OxmQs=
`protect END_PROTECTED
