`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cD+GoAC834EsKjCd1ZnfvOi51i4//oeCbABNoHG3yJrrpGer5IQXYYxmPzq3995
XWkHyMI8VgxYlt+CQ+AzfDS8dqfZm0buNVkcI9jriFyv3V3ngFSFWyOZj0t9a96S
9aVrhl03BKRcgyuiWBUq170S4tDnS7ZRtlwJcRFcPRwsHI3kjXrrMg1TkXFY0qER
S0wQdPhAxYgF5GZJvJ7wcHey/xNnljaYm88Ootv7tG1G3+pgKXPHEE8fU1pqaZN7
rXsMynmw854/BfsIOUf96t065ErlhZ/kQ4++NBJX79Upn91cVmXBP+SS/Z18uDnC
iiwE3/MU6RqtCY1xGwdM4PRaf/UqyxZF5iufpgV7jqS1l6jNgjci8h4n+M0Ffd43
mVMnI0mmI7qnCOqYBdCoJWlC6HwRSjuFUXiBPG4uzuC6+IRztrHpEOVw/qy89q6A
jRBK/vhrFpYURLjMw3RgFCSBdhojwZ+HSyyoom9/NASKG4fbUS15QJ+Z9zwlt90i
fb7BwHytjQQCCh2C7I+Wc9bVk1Gnh48E6DNC88aGEljsgOVZz+pqUx7A1+UgPb5y
pDoD0aVDjblNTQItslzGe0IQc/Dzlz8a0ZB9o3KeFFjKPeMkFiyO/kcXfPJ68feA
XVDqtEroS/x68xHbSXwlUCZvI0Vj7hkLeo3mxPNt2Jj7U+6Ye0rIDaSiR+PzrT3S
kGcYsaZUNLr0b5dHR5nCXZo1OEmzSSFj6Zz5kNYYHLFgrTLYYxi/ydUPw3SAN8Wb
l1pYy7LOmddfpoe+AcGwT4GU7nx7eZeMJF8+SHy+e5ro9EPkzp8h0sCLOj5v749X
u5e1zW6b91hegFIWZvtfte0bZazeIyNO2SYMPnSgYHTpOsbC29fB0wrOa0Km82aV
bxQdQgEh6ZH6z1q6/TN9aFXitz0IkfBW9q4KdXwtarYA9icrvuuc8ojDs3t9q/S2
RGsR8N60VCXWUmFcTgpETOLUiz2fyY98d6iZ/wHYKR3EIEcBH+UH7uVewXHYz11V
o7dPfvk8I+b8lBpm3GLOp7jLW763LS6Lc5sMrghBtiv76TKjI7T921SDBPviQ0Xe
X10eka3qzO+4HjDVKKbx0m/7nAUaqiZcc6SbkzLG145CvYT5Y+m9WT0ATBZXh4Bz
J2AL6g+x8/5CSR3MnLW26kclXI36lMmWbY0e7TjZ51tvTYTkLxayGSVPqW2LTv5f
5Sw+nX9XKKdLZlevPs/OYKFjfaAwhUKmMTfsbw1R1I+Z8PrejtCIgqbxau1lS1XJ
S0iQMOfs2avxXPtexMMuGNC2bQNc2SlLjw2hVbKyw1OAsQe8aJklT3ibDCjgzO0W
z2dPsxTJvrGJWrVpoGpLj1WMU0f5BeUU+RchsnbbEtRMNb7sYDmEFo7VePaqH5Jk
DzG5W9DwrL6SRhDQH0MJzaVPdeYG//mVjNvU2pLoYA3DOSYvo8V4kkhVzlkuDrb2
zuIBCvDMSw/qSO9X94BCdeO1JM9yIZVODCOKjm1JXjqDLWJBQxHqEeIbFTnOrtrm
wBhrIz+zPz24z04d+A3I2+HetjU3scKbbCEye6PXclpgKKBIMsIfDemxWUSaLcCy
6VajBvcxu2TnsX0482xOcK+3rE1ydMZIq6LmPChfFmmB0rwWz5QytvsOiENq9iqk
fwpP04sujXYkEsvMJpAl/dmWHRR7XJniCdJZ/sY16j5fGatyQJRlJw71RMcGLFhn
2T8rO4r8nYu+PU/dPMmT0w4K7F/WACwzjn0XjgT4hgU0b29y8bu8fJ/sVlYfh4Mc
wRxMDAYnqpm0pHlEntPKtHohJdyQjg7pFlCYMBIXlutm3NfdvvTV8A+RYvdrOEVg
hYF0n2N4sc/wKXHb2e2yTozCUpAzePTKS+TXONp7CUfkTf4A5x6KOvnOetJ/Lovr
X47n0v9L/njsa/+Y51RNLehaAzw6/M8zOzJSMiirue9ZTzplGq35FjC5N6wKL5WY
fJs1LvOM+9g99yGTwRpPRoBrLzHM9DgQiA+OdGqZQQ+av0HotOiX28vxXaiWbJ3S
dqKjYtDdZPioNOBR9giOIMFbFBqOKeZaSIPdj7+hcAVARsSuV7rJZhGZ1XQzKhBE
MMai8/pPnvT89pRV6uVvDWlA+mekeuIL42AZ4mpv3FP75pwpLqspxW1N7ob1V703
sU2SegmzCXNm1y4ZI0ilELSgCsjzyZf8XpofTRRaJ/1pPcpkLqlWhVHeHnfYUD5U
mpd9yn8If7/o4t++lQZHKbCWbif9E3wFMKg0aeEkJuIEjluKoVO7oeW4y3zM4NY+
gXnMl8tNFqWY7SyFijWs1OU/gXpSHW/89zWsXo26E45tES6eN2n1KFJ2Qb7qIBzM
pS8qbnw2aGrcussMgaS0JjTHYMZGm56DE1P/cCfyiCRqNV19Z271BlcXb5Wia+MD
X/3w4y4TRSC90a5KSfziTuvavYFX5kFLG0M/JVZYnTSBbjt4t6zp5nLQFVyYNHhy
P52uLY0VVueJeAP5KpWzZTPgH8dPujny27bHIvXsItqkti2f5RTk9CmZPTS83bKy
/0+3p9csemV205tlnMCwEn2MDRhkcrXwd/Ri8Fh5gLNJktZiQxvOV3GL9ksOcL+j
f53totXKIi9MQfcucOS/y37nuJPDybmk44kg1dzFhI8VAr5HmgBiVPJSKIovQ6Fr
wvmfawXXqPtWVgm/c3XqOgvDBNvjBCd3cE7Q65RzD9N1d7Kx6hPMlQkSyKde48e4
YMpxg1PwCj26tKuQfPZOv/MWCBPIOpz8RRT2MtR30cECDI/kgxUoII+YBzd6lQW8
o47glBaE0qhN0LUf1jea/jbJ7Qys0cIlRlVtQuwT8hpKh++Y5Xq2WTO3ZfhBrXxL
hhSq4blLQRvfNo8XFnTvGsHhx4U4WYARWwW3U5ZItnByBvMTtRnpd5QwLUuOoYsE
9O/wqYXACgbJ57ACZFDpNWNrzQ7sU4wvTPUMTfANKooFKtZV6MMvAHAC3EGG59Rs
Osh/S/xnXQMY+VdRsqbna+Y2ILK5Q5lvPx2BO3uGU10qUzkKz1XtuKIsZl8fKqZM
4dDVeuK2HbVfiFa1twq0iDhA3RAvLIeUsrfQSoxXN1iCBiLXlGhPMMg+nDQewgU1
Jy3AaCw8ebn4jtLgLuiV9rVyKxMRKeDekPfYWMzk5GJHJdXB285A6C7jZLaNPWa1
YO6fr6lAAkznsfEAxtfAtRYQxnd0o/L3U7s8AID82MWSUoccDDvCMdeljHdSlrMC
SGy18nH29DwFDXIRcY3QuV2Uta5YuvwLohSdrcJNKPRXqRZORviVOD6l6kp3WRs8
M+ZnCoJ+oNrgwKhdYMvTe9HImNmiffAMbbGknayfy1moo/+ImGfkrRkMTV+L5vj9
hjjS3kG6XLWpWOkKaMw5etMmxTmcWp9O/Q6XzRsUOtY0yf1hhK07lWQdXgRxJ1Sc
SyIJCp4JfEgK/CgLE/NklQTnkGAFWfv4yZILZdgMrOI/FS8Jjq/c9B/a7zYjJ+ma
oT9GFBC+frIXXd6hNox0o9av97rXL4FMmqiFkDOHWD07SW3FQXtsIIcrH4PXzWGg
25uWAF3qPzCiqMTnM/abIGlTMGM1gtkK9ty1H7PJugCBuZR4UasG8+6UJWZkxIfE
VPRVAUAumIruoBGRaiy0L5v6W9nyvqO4H6DkP/Xf8CvNghJvrpTM/wLmmcc7FRPC
LoPLITgma3ksbtZ2XjBhUH6aVdKChk1QaybHHeNieM0R7Urr4y7/UoAizwHtQrVR
qeLV8uUs4C0muXt/zL845CYwOW1WdiIFTRTxLKoLKAM7JyqK1uKnBOYDVoS2BumB
UNGc+SJ3Q1Y/uONnTh8ZbldasAM9+NGyMcqXFjg34M0LpE6h4lvl3YMTmYiFTUTn
kS6SB+QIzpft3v71UXBO3A1GjtB3ePx2FxaFoBKSdWvczrrkM/rmu74M16ltvaiG
hlh5yNkecALxSFDnqV73u/bC2F4e48n5m4wrEWbQIKL1AS35n0KvG2ZP3Nqi9nx0
rsqnYAlkQbDDYpDAOIKp4RNTkIOHtckBG3uflUaJcP+M+Fzmv2Fs5WbJjy+i097J
AkeZL7bS4GWDwhGZNl4aDtD6JJKa1g6n71+LPAL/9pRwgTm2/la9Foomgz97v9Wg
Znv8ellEiZ/0q8mWtsNfsfOgsrdZ/erNTF1yOkZue+viqzz/xQxaFYZdruqr5Zln
1SV/CSCUnOBHE552zztMSqAaYGhMPqt5Ydd5ompS+z0ALRc8vD24tTsviuKQMuzQ
9Ti9ztj+JyA81b+uJB7jRCF+mGBDBf4+Jb23EQebmDsDwVqmXlDl/deLIYlxvYZz
sfAx4c7RGVaq6NbFcXRLiQpCj/VTXHKBLnyz8s6GasTJ16C9WF+BqFd9OECnhUXR
V5CbIRDi0yIm5NTCer4zE+cJlB5ObBq4pp6bBQtVRevbQGxdIJFbm8oVgq81M3lG
ysoPAdbJl4ldJQOzEW5e2I6rrHCQQs60rnE0dWXAG1ncI702cRhvHRzn8SEjPcZ/
QuUgfVu9eF0SGxMBZdsXxsS7KzoiMrUm2s3WtNtic1qPE0F9+QeHcl5Oi/qVKEKA
E8gvz1Isak+H6AopLA03Rm/MUgpAyh/v1zywtRikBa95Sdq6CowgWQonHukrJfbt
wUgFQMaDthTerg50OcIBCzlTa1mHId/scSZsYUnrN7qI8XqCYZ5bJHldZGB01cB6
zoEjooaA/zKfu+yMNeO6ocm+nsiMUl5vxircRNbkE0s0SiGE6ePkgouyqWlKgl2Q
e2jw6VyG2BmI/ZOY4UFlJ+Kvh5JVT+hb6wdCUjTc+tmLqUDrlEK6kQayDkhg27Rd
z1Gla2t/06Lg3MN0vkMh1X30CsO4yR+kMm9dTmqkmKWt4PgU93gd+Lu6Jnw1aXE8
7+IlzL5BV8fNHnh+aL92cmYX8F762EHZen+XQ7CSpIqGOVMIePzYPUMYy56NooaJ
`protect END_PROTECTED
