`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apVOAPFrv7VBaB3zznWupLuW6kPdz13wgyifj+jIvoawizggKh22ycN/jDGzUPr3
G8PYbAX0Ok7kRApXxNYa2afSVAl/f6FD4m+QHvHhVJtHjaWjyZiPM5ADKR6q78TN
G/yrmZ2Z9LbwT+IUCTSpQXMCWeTYzmTM6XgyeurEp74S3Ud6hUaUTUTn0l70Tuto
jJ0koXdBGlxruvPB/05lPwia/g+dWrKbRm7LOH3qSFvaHg0BpK3opMvwZzECuC1Y
yq94cBaYlqJdNT8wffKkdpsMgaLK1RlkMHMVtTgIRfuNhJHIdPabSYOwOk7r+cNd
AsOVOSKgfG3MT8FPN2mtAnxKbZAm4uyZBjG51oaaZ1ef0oaxoJdMDe68RuMnuxsP
TVKWCfKHAPCPC+IkC4Pd2HYX7BOCs2jqwt1igpcE3PvSniyPvxYfFAOUKM5YRFOM
EuY1IMDsYH6bLKYrjyoJXmu9WoiJBlxJqRPqoDYy03+q463AZKwnp1YkeE1e+7in
cn6xpDpJdOrkFnifvuZG63GNGa471+Pw1N1ohPiSyKXq+/E3rlvCSfSi0tnSjpd3
Mauhhw2+Yg2/7kQ4aiLKt4kvyB9HmtUde82cKumAI63JX/mVZQqxdLMPXF7n8xPF
kwu4ayEcOj01nZy7cD/meybNsAn9Vy2KqHdnZzCU045y9h6PWNCSUU/YlvIucjNa
KPlHdxvMIEGlvBEJy/qgR76HWwnB1ZwfNqagKeGeIeNE8KcZlxIsDVYzr5gG/xbg
323hhekTyVlPYTMFH4SSoOCzQONAbUGPHJn+cpTgwmFXHA7qF4yR35GvEc20MX/a
UZUQ4rj/5pbB6TEokHoCGEhNxPXRPCJ7j6pzp9vXfriD1bdJfjJgXp+59xNavXH6
xke4aA+wHQIAl+4jS/bEkbpL96Igx1GuYmBA1CmwErM/wDQtSkxJoAgZ60wRao8v
Yp2RubB78vIqgkzYlnpdwxEgYPO1Uh73z/6DC7eOeT+a4Aqq7S33+NGPVZp/AQUN
/rMf3aYW9qgdI1Wjm+6mlfQPkBG+C1feIXbwJEwySw6apcv4dXVc+b6JSLaklkpx
d02z6bTaiCpdk1wYYq3ssxW7wABrXxx+0CCekNjUwOWqWUqvS14OuocA1UsW53+Y
YJ+kFinHI+PpNJrsPUwd+TKoYL6/kUk1qAm34Qzq25Mvep8QpytL/fqI0rhPuWn+
tcU5vEINW67d/6MMYGIi8mq725Qtk7A0JDU1+vlx0V750j8LbPacQvGRLlOn/k4A
zuzXo7DNGtsM6JOrlgPcFwQoFNHoLgS6Jz8r4GsVy1hoXu5YVPFHzKoeBgaHS9B0
NFuQz1DaBUiMAOby/6viVLmnaCx0RIYT3nI/AtTWg6s7OLxOjxyssR3mV3clx2ob
l/5HCizq/1kinlaArOXR+bAxm5r0bL6xb/wcoX0L03DGWnUDrXOeP2S9dlrtldbX
rZnrAWRT6Ywgm2FfWvJk1CBstZH8vWWAwZw07+T7NQR5x3QGqoTDChUtdSSAQ9kP
Oa6yfuCdOli8cDxZpAtRUG0ZlLxmx7eJGZe6OaztPhFSJ/eD2fCWkaWZw2Kk4H2D
u6DoZ/M1zSAz8CBtmswI8X0C4y+eEr4ktYuG3ljwkt6OGkw7xHXvvVFsmFQUsysG
31Lv5849WFIKCc2QqVIq8rF5a5VOmwSf9aJKvGkn4lAJDf7RkSedtgGMf3F8SBJs
rI/W21I/1A1dRHqhu5IHznwF1wnbQqUzay2c15QsRb6W8CXbcSZcjcmeF30OIOyz
2EIL8z9qoD7DkFjmus2nZIV3yLiDGesWps/AhYldgpPXiyujwd4QDLihftDHbfzI
R0DmBCgf2aO2joqCAUTcukCAoVbtsPMEQblzXXNNIfpiNDZz8NNxQDCYSxpBdeq0
/ztNbNxIxSQHkC7PABYkGr6uI+Y0NKsg47UImXr2kYDynaPafuPcCRqK5w+Hyy0p
zeKT+sOW0LPE15Ve9C+75i5HHMRkD75aOwzWPFuLOWRZf70lTLPsoErFd4V8vVG3
sz04PepECp61pjPE21oMavc3OZKSMvIU12YD8qQN1J3w6jFbZWAKvlTeSnV4C8Hw
z7uLZJT9kLaJuIXitAS7jnbv/5aJNxHjyv3oZnEvxAzegReCxyR96pfSXqhhzIFo
V9lBNbUv3ENKFipGZKTOsXwybQ8HOhFdELWS+BuNgnXkxo+SPU0C9UcDcnkXZzgQ
YgKc00f8EwUuAT8nlXR+1He4Da6VmrkLXvEPAIbc+fhBfRp6mM0N31sXcTblCO3+
82Fg9TKU4DQhSOAjrssxnjJkdVVPpmwjlyfcoj/uhz+xofJq5kI+374LHhZO4SRz
Ib6Wq4hkBS2G64WAYBM7ptM2s2+zZ5kYTC7k6eVDHJBtF3WlToycyrxFFocYy1GD
k8Ubo8+upvDd1nLEB1IgMv9IJ9goTiaCNQcZnrnrj1LQX9WfKPnbuG6IcUe6xrYk
D3VebJ6cZ2UxP0b4CPPHjdTwxYnb8rM00E66qIp1UZzAQpYZZGOihM3nWs7NUxB9
TnunQOvlHWWmgVAyRflw6NccqcU36I0G4HCdKPQ874fvSjAn6W+R6L4PWDYdQ8DV
rEbQ7Kk5faVnaJtTlGXt4SY199lXAH0tLLGylyYKmzY5ckempwFOJ2JbUFCf92P0
tj9JR0xFnk+S+HVIJXZabW8jtwg/m7AKD1HVzh5EWwGZ/D0qYp3FnONYg74HKWk+
WlrMFxUBGtcng2Wz9FhpT2Is87fho1Kyo/aUG22PRfnM9mUWhQS6BU0bPDsfUu9F
SXlYwAFmz/X59YcQ85Wn1tOf2UBJ/EunITeuXCCNjwaYkWS7G1Fq7FtK9f3Z2w1s
qdLVwD/mMMaTYY8LWpDdaSgf52DUjO+bMRuDRbBUu+aZxQ1qdGkgacz4Ns/qm3eP
KGAYNKXXwBvDna1hV0H8GP/aMkr9JJ2b4jwuceOtJwkivA2FLrxMORfCvUDYTABb
Dk1XIcTo41IV4Z46Ois9aGZwN/XbnC4ohWK5JAu9BXhUUWooSe9fsKUE6fZKLcdu
h8kdnLsYCoaiz4K3DRmC7FrG1o8O5VjUQ5KEytkc7wxxBlvT12JTp1yxtbqLtZvg
L34a8b/W+F173LU7lUHOfV38IVki2WKcHOvAvsd2nEtESH8VutRmXIcUVGTsKTf2
EC7CwiN0NszRxWHtyEOUHlRCoJfExPdkbeAAw9lvI+ry6VKJLsQ1cam2Sff+FYAT
8+BfLLH9qK4PhwQRwlX3LbYd1w6BD4/s3FDjTwUJpYKJFixHIGqV+xpWohGGZj2I
CZ21XJvex1DTt8f5dClAoeOkVK9EP/bQ7mZ+zkUXFfT8C9X/z0qT2VoAr/cXslkw
twJEOWCPDsIW94UjF75Dcz9g5YPukPBKW0kVIE2KAUCe5PBDs82yToyZHv7tCA38
M7GNNJ80h6QywJXtaj+/hAAP06uDq7LjPYBvhrHVKTpvJzm6GlQgrwBh8nbgctKR
WABvL+VGNBsxHUz/l+f57xwsNC5Bxcs6GjFXRkRbP5Ex6fNMffjJOT/XeZt+A5FI
C1ra5dUI0yVE6XF7ChzUZYIQbjfqvzRsanxp0UMYjQOYV+zA8kdnX6EH3PL3D1Ny
CoFdefao792d4n/pp75pL2Syi5FvfG8j5fqyxqNNjtviTlQ7g4fuS/IF+ryh1bw4
mX4fbt6U0gAmeFfE3+j3nQvuBhsHbiw23rEpkbrWfJkBvJWvWUbCua+WFscHvad2
ToZDaTgMv+U8ropnq6s1FbBuahJZhwKoYLqWpPoUs98Fge0+9NsTp6Uw5kxnL7v3
l8EQm3UBZnQpN+cLhf9fe2L49yS+aFv+BvEiLC2La5ZeBX3SbZ7ayy9gd5bWe2Sy
WjHdH9plmkvVKDuY4EdzxJIQ78W+RzjkeIVbdqUATB4xHmxua/MzFRQgCXeU3Nxk
KOS2b+KmAe3fKLAQT+Zkcd2bVfxZsU60S3AkpyqyzeOxilqRjg0E6LbEjRWSUJSt
3gtORMQhJkHSQyTlIFQxGQSM0q/SCGDGH+CDLnMg7GHuuLg6fmFZ0phDWoG7t4rb
oG6hHy1Ltctx9xevVWGzPm8pTlMeWA/Y8qu+1W7ToqQ/p9bOXX1xkdjmFQn6wpo2
58V1zbOxeF3zX1zHNbDUqWjRgpb8gEreVrbvnQw+px4SyDghEwDiw6XFNaQhivDn
9M59HfDt/TPG7+Qpq3Ha76rFI+135zHmFk1VwWBMz4oBhZozFuQ2LlqlbYyUz3wI
o/L4qwsqxlMDftRoRa8T49cKwAWO8D61uZFOynDrxdi7zmd3f+tJopwVK0KS4Qfc
kOBbAM6P+1iaWyWbJRTjUDJFPOfP85uIzbAEiNSlBKC64Fi2a6+A4YHuEcRAgjJh
frnWZovrhpH+DM5kOn4kZntRl0whyDjA0y5/3OXewDUOA0LfcjdnXF4sskUwkFHb
sK3hx3WoG+rd4DYdAGqsBwJyKRu57dCjiuwOcrJthu8mnjLGoew2lDQ0ZZZV3mx5
5Xt4LVVVSqpsNW/9U1DmWjBhVYl4eB2VR3z6Lz5oEysTfjfmw6R+OfoegNdruX7+
Fdl8lGyZtfxyx22aR3i1F3C480n9nwj2v/YQR5CsvFtYjX/hadxMqHpC8dsE8ZdI
ftuv8t7ykfGhPcS4+cOT1n/o5mhf1/0Duv0hyhaztx/eT+Ie/owhJL5jmIYK46jh
lgYbaHPXiMMqJ36tugARFQowTXQTYFkfamr7wqRwyQKjTOixQLcMliwAzeJEPvDs
00Gs2C8Qc3j4SlEolqE9tRuQU76LVI/mY+LnPthHm2igtBs33tbkMtk4q4Xp30+a
SNsRAwmFUO2yqOrb/KrapN1BU1eEpnEIkpNwYY3jU1YBpRD2UmthjOWYolkC8Zp5
BdNUi7BpZtViREfWwpMnw6KeZWOO6kmfPQ1X14PFq7wY0HTcq1h416v/KKTQth79
9L9fT+UFGLZq2W/SDsSRZ/qxAs5DEzW+pUcjhSBo5FiPbDzlEcBQHShIK6EB/pHl
JDekiUSJAe33EX0WB78iuHsj3pFV2Csz7LFgTJOOeVn7hzMleQF5B/TKmNge5q8d
+PzNM1UmJkpZ/DJRMuhLUxRNgAS9HoP1dnsvCxU9RY3AjdbFyugUr2syB/r0BW7g
y+bEMaNN+bBUGZJ2lgalriPEqgiLWZdjBmSYoQdetrMl01vejRAnGpCpBRRxqb9A
l21TeWOHzu7B197QWb/4OBDmZDKfxFZ18TxpMWKmW1GBic7oBsEEysKOhjW1Eqb/
1Mp1eL194b2fqzoxbOsKkwJCgyMLZsgiKyvuUsZJEnj+OlfBNIqsuRZrwNZQLejR
FjTtPeCSabEPEXGSzwLr5QSd/nfouEEu1XsAl36OfGg7bq20ysJewRUvZWBupZRy
+s34jqBN/U9Fmx4rIM2Bu9Ctg8VzJOPc7J5cSu5tqHssKrSY0TXQFQMEN5PhOSsb
WtNRuqf0xMoTp0SCuYKE2q/F/4TnhOXlvtZBHUfJfu+0gN70UyVVR28dZC9Fj/2g
kDnFKH3jEYhZOPMD2yKIVfEYVDQ5TZRPjy5sf3cqOu5N4BJ94fiU8UbT8481qhed
eLk9ptgXQX57JAt8F7dENwAb4fSOyR4gfdGfdhtsnOfzyysUZaetqORSpXHnuM23
y4ut//OmEZD8DNmpzLbh8KkecHmom+fH6gANnwUppoNo0v5lHrSSJ7uuKlS3BOTC
mRJy5IJegajS0A+XJ/nrFhPsP8Vr5F/iLOjNExQGNOGek6ptgIUonIKZlxLhAq5U
ugT+0IXiVtlFqbfx5zluL47duj7T8qZSSc7fhWNDBEBP6DoPnjeijLMGWNBx2M7B
C+KAVgI+9ZRaqy9zsPMidFv4SAOoF0sCYiwG2P9rE68Wl0TJRdqBJEzCPQ55OVzM
l/0aIq0kTsdwwl4ACk9F4JLj7tJ0s3R1vR2ueAiVLZ8UFisw06Hg5G2axUR4DTr/
d4TIM5VG7Ny4by5vZQdlg3jv7ePYu9XRbBw9mol2TCuju/Yvjmsc7KorVF7b/Mh2
1+DNb6Gg6viXQ6LhSSmvfojaDm27TbTj8vnnC3mUHRGIuSfZPeEAyJQLtutSRctG
PGQa6vWL5ck3skSrtoBAfF+4ixWAgdi6OPLjQAFFQoOfNxb+ntFNpgAqKIe8HBGl
bPyO1Em5tv/l7TMWLEvpnvWEunERRhOIqIuwnNmaFwFtUuQx8VPcw2CCtvksRvnA
IjS2cIyi8Lmec6W2L4XwQT9K8UrFyBlerydmbTaZ43sMIIfzOfgylLkTZMU8xlqW
jmpWd888vBQvrYMaDHroG1ibmQZiOC2tv9qDA1zsFMBJnwfLiEkahnDPfH7FFMGu
oaAHZsx4xKqEEcLgcTrOS0pbbzXwiv/qQXLRqyz/tF1tlBnu0VOh8SJIQjKXYTZw
Gzw9MKorGwWwX4/Sw/3LxGi2qWOFghgQ0U6Vd3ef48QJ9qBsb4ppWtPjdO3wHQuf
Uue0kw15EZR3MJV6T1CyzvendP8Y1rBzOHDkUcXYrN0i1kVNP+a8WTZqq/ZrLT8g
Ma0298mAa7wFULYacZJ5LXuQEcRQEOXrr3VPn0sXpw54UJab9AjNUBDSHSZqWH8s
j71ghBk4pz21lc9VRjNAOBEqcZRBtJ3HdXApNd8lhBSV5e5XMORuS+wgn1sNrYCK
l/TFSWhBfnAJhVEFwYhXcHOAy5Ow4TH2ZPhaXWpee0wAWiBBpzStcthkraHQB5ri
5XeCSA1dDfs0VjuAVO4bz9oYn3FudVsN8XdS9z0xxSlh5WAuZccFGUEUtwA7mbhL
UqNOd3XdJRwUD9OOp2iixcPMqWRVAoSvyrkD1y2oIcymlIjTa0Rki+On3TiJr2yf
2z8hwVo9ca39rW+RC2PLcZj9P69LP4F2i8Jy9drzQ5pmhPeaRRVCcXm0EXaNadjk
rNghX8MUhzYO2131W32OilC7MrjTjuxFhxNcNd1EnJdoV79KEcCaKjWqaTcACoWx
hW8+6ZSOCaw5SyYcYJ5u30NQ0cCn4jAVaxprQjPGUdb5fdQoBHdApYvYn6Xz9f2k
nrCJNI3+E9j3OOuMgJu17nfEq3UUwtD9egzwLFwQ3Dg30KGSBIDfd9kIGmoFkJlu
V+sAut9RQ3B/Pa+rwSAqDzm/Xw6rag921K+G974SYvGKhHG8lZWIUB+bXWYTmr52
TpFslyn97lzI4X1yrfkiSZ8Gl8fgEy6A2XfYPjqAVeNPJAhVpYDzO1tZq4OnL4Tp
Z5ubKFfHuaJRqTj6QYuw8tChqPAmrQnGKbUn1G0VMpEqrrHMQcV4yfDWVCPvqg1z
3b6oWfWi9RtMguJPwyPEcq/RiLK66i2F+5iKjkJ0padwOjBnW4fLTLBirYg21lf1
tKCOFnaDFscfSixPq3fbUVGXa3gQLTB8tNPEyBY8OxHjeHX/SumUDsd81Se2etQJ
YhJUiY+Tv4Zz/sIldfkBr6PwgPn4d3pJzkZE/0XE2hc9IfygbXJzUwMyzXh7/MYM
Hz2HxcwNVlORpgEU8FHHxU7m/J6std+rCe862A/CTaR157DUTXrfdgKKeki8HgXr
WAdj9zQLCxhyVjQbKoD+iLVvOrJF6C9WdqmYabP6RU2rIId4yuoKeY1fQtgOH9eH
GJLgfZ+3HUnWqqDKq4HlpJx3gsJF/PmsrrygYgyC80R73mGOFcFlk4yW2mWISBz2
uQneEojTfPJmambCe3I3V3tEfzYYiNHPe71zguvh8YfKwR4xaYBNWsnBzLMybnUH
lY1BFUA1NDYOuEtMs9F6i8njKcRh53Bp/sRmY1+iisItbT9pLzohkvtTgIhx3+5A
Px7yBuavqJkq0vl7IynBkfB014Rc8fp/LxlwktiDUyXSHXD/t0JEiKPuGQ4ERkmW
w35tpSPiTYjozz2gdTZIamF9IHGxHPJ6K1+QnPV5Qk5v4e8E05qRF7G3gegRMOGV
gUZll/nLZ1wd3wnJ3xt3+Xkv3ETPJFXbDUOkE5xv2fM7EKLJ83B/0KxJ6e/ucRkL
TZP5a8vt0BCAMJMGnHcNAI7RsuTSEVCMKwWw6HC4/L93CIbUaLms3Otlc2IA44a2
8A5AP6/ahkd5ORx3ZFe5KBhJMkJXP9/Kniw7stcrw4/FQBdL3pkJOSHCbxbvA3WF
sct9qMSRVrSYei6TG7yOEHsjQPctg0auXUbS9LLMiIiOb8rumiO/uWiMnNSl8dDB
Wq402PpWKVNt1GCTISHOujMrf6x3U9PnTiSz/kHTH6xtO/3gJZDEGxd6FQvMYq/8
ow0KEkSVxbNQvwXMKtUNLxAo/r8Zl71BxupYQiqzNzHr8JKCD7LLzq6ev8b2cXSA
l63qgiN978S859QUM18WM81DINNm47KJ42uYFPx8lVmbg/84MkMVaICOLGJgmBR1
jNXVVWaTzuHqnKSz/s47D+gct2zgjEERhhuZyVI5s9+EVHBAGYVp6bhTH7bme1oj
iRCXcZa+Zs80X9zXTcVGnimzHtllsQPiLEfEk5yR57R5uEj6zlkydyhy/g0kvIEX
lqzyySc2h0MjMu1p/oxdsehgzxALjiz6w+O6C67xUnKIo/dpPODoJLMKQns6+wu6
msybyfi1344PsvvKFxHhqB+8xI32IdoAWD3n0m6M865Ha1HGQ/9y49nOsgKGpZFg
W9EhU7n3YKLvirg4NpB70m4snuZ65f27OENBPmForozfw5SaxEeDk+VNx79jMu2N
u0YIgKYoNPAZnDPzRWSkKTD1Urf6+8EhOeS6ZEmdxkI2x6nGpwx6CO1QmDkT0eHm
UhsDa/T6ofr19b2C3Baa2evUMsyKS2HPylFTfVQA3nPFjb8oMoSBWROTSq+TNnyp
GRgysCGqj1pvZZti0fVYM7GwJn5gz06b5aASLKKvc5WOLAxOzoPTv+sEufD8QqZQ
E8YlQs1xX14C8FkUntknM+iGV8IUD3QLdHQaorHTwDywiIIUKBIT5l0npF2r7dxN
fIqRVP9frU+kxjOeuh5s9O4CQ+lsiv834tl7J0LOHPb+sGN4P0ZYPrlCXXG9npNf
cHaj4GY5EfbAbZVntceYN8Q3RYeHQwtNnxX9U+ICjYgYVBaWD94xSFEMEc5LongH
SHmeygVUkDGKT2hIbLFWsjRP9WI6dFbpaP+ufB9EW89jfSpmPEVG9W4ow+1RSkgo
CGSMXRNKRkZm2TtvOt0TAsKPNphFjbi6+oAhDtjTsduDRw28AF7Ya4lGBr6u5MOj
Gbg7buF/W3mxt+CfteyytB5R4o0jPJggvGW1b224aaXXdQ9dPAJ8KXvoYiSVpY3J
+8BJoYqnnsljPJPtg3iQ92JAd3pOjzaNT+lbZAIMGbfsAO+KEl+PiQ5kdewlKQub
tiL6+XgKlxDmSjAUTAuo+4etkhcNDiNURmetqST3101Ys3Zd8lblDF7cjU9pMffl
wXEo8jNQkrls7bdG2fcpDPcmKnCVQCfZBR/dWNilV5zmkAVaoq1gvYcqr8gdIDvQ
QEcXC+azPTJRtShusZMYDMN7QaNrxFsFs0vhLxXe0oflAjdTe2uXUNytMOME53KS
1V4CRxbueHkIzKPmDKe52n1Q5Y3L3KC43jA8266upGGT9AGd79Ag6XeXlC9eGB4X
brnuX8pctDs4FYl2sNtTM8bdoUpsyRNsHZGW/jzpmZHHqhAIIB0TT/5LqUSXM5v6
eAyP1YSTvA1+TdLc8udVo4d4JyrfCuSo7ghfffSMafHxzQgaPT4eBmgBuB8nyJwa
zDvjOSZx/ZxjCrDPMcpgjIjEi5OW9uxs0EoKVMNEmsjMq3A686oiswUtyD2ihtli
JO/dXNphkJ66qWFa6mHNcV2Lt6Rpay758wr7zWjXOU5O1I3tQhUlB+KQaUGXH/yA
0SDdUllkqj+rlHNeedmC9dSdcd45HJ0sFwY/+PVMBfweOnFT+UyW/+rdyw+SpA4o
fotaLjen4qtRCKEgNw5a/YIqUdaCN6tCHR0pEfNGhlYcnvejhwYehYBsIpQg6jK7
wJyzSbATKlpyaRUU9XEHm5QCi5eFcC6Ry5X+JVgeXrdDg2cVvNQT6KtXmIX3b9q1
Z9s6luRJe/EYY0A1+sGILGhyi++isxflMCjsDfq36i2PdKsF0JIbej8dVIzJ42Ru
sWP0yxbNpi0ka/VTsU/+R7Rtrneazwlof1HQQXFIP4vAjfUjLZrEDA7vNbmop5LC
bQRHw5diPnhydSd2g1Rp9/YR4bOiDMTChaeNEIU3AeWn6jBwoDBL6MZCr6ECkZOn
WymY0ucSHEe87ytkAU5zwxb+E3Qmj/uYf3lNS6Q2WrxuoPRhUwJ4EGttys957uzB
/ufmZLw/bV6VAdVWqLA4dHAYHRWuO7IFo7GVtE5UckSb0cWD4v+Zdus/j4RDCkuY
zkW35qlBlzW93SIQfYORlq0iN94dy+2uSLrpxqF7IcNnhF1NlbzGnxqFHCRqjSca
mCfU18AMlHnyWUZzmJ4wxCBq4wUezhNo1outPrrD7W9yMFDWFNzWTc4GjXKn2u97
8KWg3ifGDxRgCAx1CUpPw3XOdU76a+cYIAE6LaCbs7zkKNgRtYhiwoL9DQrC9DOl
DzvxvPTRUUp9IWXEX599BOkICWDc37huXNymCjTKFlyR6MfFHfQzBDAgvBL9W7h7
DZSQHJ1U+bikLuYiO7p8UQCKiIdGuAJyoLgKflcQqkegtHR5dw6+p2EOqzOxgOy5
L3I3KITrUkIX6Vg/ScSIyFQFyaT1OK+y7nyqf8ipGthClZcaVTHZHUsbALwoY7hk
2HwIQiVAWPNOhk3k2p8P1ovqbd2T/7rJY3flca2Ym+aP248z1+sBbOdNERX5IY1u
/DJgXpsGnEDeIyMo52muM0TQ4McFO/q+ySO6dY2LhLgoeggpEwaSHdToN1no+eKS
64120/EJ/I3Ft0W4j83r5VJArvQHXelyvZ3Wl86t9K5M5C4YvuerJ72dwRZNn4/L
iu/YTWJgWc9cXIaylzsyQZwyTAAZgrEsgKI516bZuQR55DU/EcDOfOWsL1ohElwQ
GEqWnz178/T/tvcvqTbgqk15PRE/pIC+C0/b+1NXDeF7HUIDK1fVLEOEe2RBBDJ6
vM/raGX4t1Is3kt/wpXlWRvm2y7eqxgzA3QcKHX8/6lNvqVFJj66njOYTe0nkpCZ
NT2p2i8b0yBeFCsEV8dSErOE5z2+HABpizFZ+UEBc+HSIvMlqmY0TtuvE4ptj0Oj
LbYD8yz/LC8eHAdbZlPr8wV+f2z9z+pM9eC8EKmx8I+q/MLfLLlfozWUokMfrPHM
1FVCGwlPayZQUPi+vvd0yHJjtAGJnt80vnyf8bObxmU439uDgkx0ew6RHrbbmJOp
DVb9drjDgAZABO5pZ70TmxXWKBNOZa9HtimUujKr75BqqZShiF5MGt9NpSXBEeFJ
vGrt48JpSQPlaKHf0/5X4nUKMLfpkKUhV/dqZCGUIpJyhea76rB5c0q9mmLq/XyE
c3QvhQwS0aWxG4FvcvTLn+y6YLypALfGW9aGmPbdmpaNMeXr5AvW45DSn9KI+RgQ
XCVIFIOfyECm8JQlDzC3id6/MClGD63UBibMb7EE1kNNz+tbnpWexMDISXY0wwqf
XJS7eOsINWACmtZO1pCHyWmJZ5ZDgkYuxN1p2QfmYSnDOaobanMlrLGcUoXjwqBk
w7Oa6hPDtUVMgobrolFiAugAHHssUmgCNLf4LLNoW23isOM9JdxEYGZA0KfRgjsM
d2j2dLMC7eEndx8LUNqs830eomYeWityKkQL7JUnRb4Vmo1iMu5xGoZzLlxasBIV
pwvB3loVdjNE465MsHWAC5f3oyjwSxJgwXY+ast6oiV9wCrS2wozcdTxMelXqMX2
ZipsxAktMigVtTln21Tsv98gGJoR1Ex7I3aB9Ln3/OWtFGT/94p9V7AfJjc5v6eq
AdBT3QGkkfpo9ZTO3ySdIuHlFCu/7F0MnQGdPc/ebyVtvIDR2XNgApGi5fADCD4j
H7iGqbh3+BBH76fcTx3cfTpeZcJIdLc8Cah8Hzi/YbwCKSFrLPm7k7T2FTd0O4zf
0DCPd1xMQsS2tlUZnEgSS5KqMpbgemUX/OBx1ki7Nc+D0mU8FfL0y7v30jAWqn5j
H+H9Be5YbsexdCx+5uCD5z5ZMElh1aV5FGYbIJFTH++bx2NPMz8ag06Ky0Jnat0F
KYUO+LO5goxsmswREXoS5TUQCBCViMdoMrCYVMx4W70RSPBHslStNnCJpwf1NFIR
jpHDOkXL7fpeqCapIuQVNylxqrZREHZa+ZQpWhZCYoHwq8PJ/5YIYWXFAmuvYQN9
lm0gqd2TTkVR6fXrTHskIr9cAF1cl5gfT4wC6AYoElr0ifSmu9RIFCrRm8JrcVG9
TMjtRm1pe8cBurtEtkmf0rkFYBahaJcjq6qbmuMmcbh0cRbo2AEuev9fUaViGFPf
e64oSUjgPbUm8xRvpNlZhDtiRU2azb2tBv08IzxQVlacLnsa3ubdcYrTHBfnokyB
GcvnBIL5U1zZfqz52rtVg1NojJ0pv6Z7t8WZmW33OBfm7QB538MxsbQEraicpg36
7KZiIs2oR7vSGOqh9JA/7dJQV1aDeDrnp1NF1uPBcOzDeWSI3hJ+1Uw2QrkMQhxP
QlSqbHk4ZiUlAEXB1jzl578hcSXbaV22ns7bR2DJ7r2l8DreHYsYTdMRYgc/5C+7
4Inx0W+3sfod5dDspoNtdLTXh0wkqPyYYHnQfCcLYQqgTnPV0Fsy0a+foJTIz+bl
NiVw2t/Y53JaB6/YQpF1LyIT3qtoUxOt3si36abysODHOayr5Khlggwb9TeXqQUB
HNdFCHC9FMe23ou04y6kiIJ5I09Gd01UgCFC9bq0uoTjRHDq6dA+pVICSvCqe+74
ClhqiKd3urGKx8g1lh2RMC4exWjplU5bEhYbxT30Q6DMb6gErSO6mACMwd0bZaPC
WaoxwheNYpnV1kKfWGK463Jo+gYajXdiyLxlzxN/BoSjCBn2P7xUsx+2hSZlxMZC
9fEsfoT9oWS/Pqzt6muwCZDhtBAmelwx4Zo/ARmdbmLSKiOQ14BrO5DYsdM+wWMK
4yyPT0e5orPMG6XGE2Bq/SfsASvs0C8bJ5NRCZ8ROivQzlbaBpk1UiNMDAYPT5Lh
kY1wZfsF/2vvoxbqdWdmmu2d8Wim8CsGf3FoG9Y0r6CRzXG7tus6xL9HpqKNIR9k
PFHLKaVovOSR/KpcIFUpaT+Vmo1t611SvtNaPGiofmoJfFo4CcYtq+oxg9ZSIpkL
z2lbTJuHxYeM1znQtVNoVNewmYAI4oRRYS4X91kX2EnMsJvUOyIY/YbW0ld6DtrO
Y7m2sR9BXqpPJrrEonNubgLpgoA6d+u1d1wPZRiRovpyJ/pXfpX/V7YnGWqezhcY
1UpSove+PGQoefI8WuNUgaN4FfGTqg8a9n4KWIleE/ixr8ZlXqi/rxUrQHuPuxcC
Fi21nuKtYn5dns0iMQ8h6Tn+t3RikPY5Umpn8TVt10oRpCFByIXbYPUGoypL11Ad
E93vTMowOcCQPb67GAD1dTc8Bo03/V4gqdT4Q6lk693H6tjTsLZjgxpyfddfVUcO
mv/vZsOZhsD11lB6NmtIbjAR0w/hb9Jqy/BnDHbRaJoL5e4RnJPZimEwmvdXWekL
DIjHy1ajTBdp8SIcRTaQJzjmlrOrsqy3s89ABc4pXQMkkYaY8rW2u2IZ4jbxjcnZ
sNf88n7fixMsA37bnfKHo99UxL4oBP1qBug5vXZGl/sxej0lzCdp+ZxskEkApDZ6
BcfTc+tJkOG2u0dGcL3/Q0mVgLJyRxKPrhuBRqMwCc54VwVq4exbTDmAggXDbjp+
xxweHyku1qQT7cY7qOhBE4NPBOgo44WyYWTYnVyHJyMG3oe2hfNOgtsdTaqIN2U1
GG2IHu1TrhFWPgZ5mchgXUleoj1sAmmXErjbyor8IgFeDd7KxBBQaIiuZG2O61UF
I/y83Y8G1fHc1OhjGhy5z+txdv8vFnv4umQhN/Qk/ubE/yoAkOvLlQ8RiIG9EyEA
aszClVosMzFoRldhPIJ5AP8lFATsgnvNgIhqJfioCtA2mmvtPSL50IEK6BNno3ul
s10WuuXt75lw4d5vx90NNkemuLeExt5ZXGgVHkOgTKIlx5aA4lzWHqepu4hFQfL/
P5RFjRmratO/dUmo5sSGtwVIGXu9Xg8RbJnzlafqbS5mtUAoWtS76+wVgzDXgGmJ
ftCUutb2Dbay+3FgxzhuqCP0L0b+OQMEx0f9JnM/LVwCPue0J8yh0p7oMJoylkYJ
Gc+YF/0n+YWiAPtXc9Y2EFCo1m7S0Fd4KchPJX1eUj6OBPZd6wFj0WAiUMae1oVi
nV292MAkgVSQ4GNLwSyJxziD+mvX1doyqx/J9i99k9DB1PhKiZPNbN36JKK25bv0
kK1I52QkKwXCIoNI1UgVzhEeUiZr8p1jA0+VILQtSbbRJAxwL9LULivWvhxdu3yH
9KiQGLsUdM2fJKlZboOYTSPeebO72OmDWmVad/EvDv2WBU29yNQYq/65S2nmA9WU
oYyVbtumVOhL1igbJtfIxLbwPxCaI49WYWMtI1m0gjQY/gm/8XJGgJ1NdGXt76la
Mz6TINoxeTdABsHjjc8T8OyXXfFPpLRfl+TTrRpenQwYWsDG8ANTN0x1u4xjCoEb
6hQRo0byUYRh1NBX2bZsbb7wFzwelretODpdVys+MF7de22CvQlIiH41Xnf+3Dh8
HYgC3G3kWywAhaZX7A4MzxEFzTu6mWicJEmggZg4n2akTgnP0lZEpMHL/iIFETs1
Keq2d7DC1VBfr65azd5dqFIZM9qCukwyyw5mS8vPIXpEwSd+MncuhtujGZwI5dBH
s780kdSNq4tNSoTeZ9sVJt26uyBohesLZLcjVI8BsIwFnV1WaYkfnDp/5O+stRfo
GSuMDCeKYPqHQPRbjQSOkwTT+29HvUgiQ5FXsHIIyuc2rjd9LUyOGNzmFsNrjbjE
NvdTSeD/PGqSwcogXriOpUweRtSRDgWNj08mNrLQB1obd3kh5AZSiGjK3z7XNg9k
KTruVYpeRuynt3BrnsWqQnTM5Ebn4Q0bY9amKqg7FPb1okKNRoIuASSsKo0uDzit
NajV6YV6udhylPAa3jgX5DvTPMmHa4OT3iJwEeRFXAIaZAktQiwY+0ND0YXwTvb0
b3bVkz1pj0AgYJpU6bFb2y4nIbFmPc6dDSfZwrardRzDkErhH/1ljLvBdR06Urig
0E0WpF3U3dQnYV3tagQ6j7b50fyJ+QRtHcfD6tHjCFn5RarTtDwoENolPQMflmQB
bLVaOyzYp5d77Iw+GsjW/o0ENQXOxW0mjcbAc5Kkekwb4NoAH4p7v9lP6HFVKY1W
CkY5w8/upcGAWuWnUtHVjf9yipNwid1J0c/zBQoovpdCCfkJO32ov0bYJ5uNPvBr
DUHW6xF7weReHz3zNEnfvhmIzMAFW28zV2efKauwn9euMKYVYRYp/S/I+TfcCVZt
ALEVKSyIBo8/TYb6QYg7+m/e+pcdPMo5k32N82TQneHujy+i8qQkeAU93fBUQNUc
2K2BgNbcJG9hraKPYJRQ13u+XtA6cBrEBbLYNlTJ7amiE7z3nrpjK3Q/g+yJUfj2
ciDyjAqFi8CRiGOV+ncJfsB6MERBNE6QPCuodBdcfRa4JkjM78dRbAUvn+JUkVq1
GoNLpHbm8Ox4nX9dAcqs4S9jpmqgdIhXjXWA2tFJj3AkVYh2lPBPqrWG75O7vhug
9i21NWwj4jYI/XPr4GWd99j6xNkHmW2Yhis5UMGfHZE1lBRdpftetj54OTdBeEVa
5CkrGQqU+m8v3KLciQadfMcC9+vJLKcalcNfu1cxCIIq8zJz3F6P9xt/4+qgII9d
bxpwJ7lRI+hbktfjnPJ6NyWdMZXmI1iXEd+vGpLzjIjBkre00ZujvHSKWZQBkcAO
TQLUdMnMZ1tj2GBRdkQXiEKMkgnaTtRK/lK8v1iQBYwLCEsC47RNJFpeU6GEvwwZ
McOlNGihwdtbB7/12o7OrnW6s8EtACP4P6N69oEktlNc38l3AUyOLTD6Ts6lXUYy
plHvPFH5cz7tDSesZIUDNVrD4dFeSQagTRIznoF7gVRi7jCvU57PEl+t11pBaYVP
Gue5+QKe/XNlaQ7W7DyYbm3uPkrJzQuJZjoOKqoqj50ZAusGOzX6gX7mfzrG1QAb
PCOQkmRQHAmaq8dxhJCeiMdxpNFnTALle2Xc81zTs0AssxatIL4lPmf6MKfXIqut
b91IQ2ZXgJGd/WEAAYtGnwuiDQCIKxkrC8x0YJWozJM+KjiA9YyVpbtdJZRgCONk
W+H1UtC75rVtLtjLMF7x6RxdrcIAVUVLTs+nnmpH/hxEnWCyFQJtWxMlD3J/k8lr
evJQ6ibWn3bcTIlr8BQZ2EnL7m/N/F9ttJOZY972Ig8qnZME8TTPDKkYOVHRuRbZ
pkdLIRBVeYbEPj7/2Rh2jMdwgZXrUn+AVL91oLBwaOtSrgZYEBmmI2HU+E7DBLZi
7C5lKEXJ31IC4U85+S7HxGNt0S39IznDArm4ozuF82nwDvdNJOvzo6SGEvWK+shi
AleVC3C7a6D0n+LkU1CTZrAb9zxSo4GqIEd+pfqaXw5ebr4FJiKZ6jytiKGlvkG5
LveUI7Ns5WNt7xRFM8STudHCk1a6KaLhVzm+VBu4bt8h2zv95lI7K4YSrlVYTGEp
7Nhadi9DAluM7Wfz7TB85JC1+uPc7PzDAmHtfedZ7kfvX94FNYNk6Oj/fa7QrPr0
n84W9fMfDt9CaODyLlvUpMeisywzV0vNuIqNbyPRxrpS2eYQxNJbVrvEQmboWSsF
8gew6ObrmdcR92UeFW1na2MFOOckhYVMavoHEdCTE/vJOuSGW4R4mIvfcbsONl6V
jjC3kfVQkyjlUJ/NY4LAbzGVtbhpxV0nqu3cwsqiA37dzgcRbYL/P4TtG53Z5N+v
5PLAS/bD/nwn6J/jOhLJ8ChChg7tq6zKBxnfbKLHSAeZEY6vVBS9U5jPlN95e/Zm
n7fub3crgwSAxwFvb/w0iEpUCcvwHZBqGRl1F2xTRdJJUO7tLvzxaURWGK0h9ZED
bDGzYcUEeb0JNyHoNnM/v9NKSGkD/SAGJZZQDEyhqTcrD9TzlcPXkmK6ifabXgZ4
HctPokRggtA0cAqDJ1iblepAVRgw2cR8E8wuuNDKSUUbHg4/UUN01At5FNqg3biK
ze6shNs+zEFEzRAQi3aEw0S34e6Jl8WPeSxYtiRiizS/WCDu2q7vWi9q0PphfhNs
/c+ZIAabmO1EtcfX6yoW4ERBCDFYiicqghNDA3lV2hk4XJZ30GeLS2TUCa2sNH+Y
2dRkqmFUEKa7mjrxKK2gsyjXUcHSPEM9B1R5vB45+/wNfH/nNrr3tFwiuDNZkchE
IasYDaO5DZDkW71jBn40HmRNwWiErhGcbzF05BD2rx84Iq7txmS8GBacIWR+RVbO
NPQK5+hHxOW3P8U/shzvXQ/srjHr0rtZHp8J3GC1dOoaeNCTF2OeAIQcjkPSUaR4
kH7Y71ZYS2Gx3ZBAO7AAUyFbOtVGbTEIi8I3jH3SUezOaJw0EPP54kh4icxxLh8k
3YhocGi2mZFgjn7JoLBrZI8plytZyG5M6r6L/dtXz5xbIwYVWP69oBR1YtfRqP3D
6sTbXF0ekZ32rJM4OD6YGVtAqhJLKZKUMaS2wb0WXG28mR2PgVDv8CDIq2JzvkFO
XDL3r8BcMYKR7QZlLGibr5rIQo4dR2WsYdJUpL+/x8rGLojuWHXQgGIWbd44q8Qz
k1cbdqGkZmwNH5IhB0284LcIJvY9doHX/9NrWa/E8gkmPdfddfLoECkks83jvr++
n8Ld6NAs+5CtQHlC4b+DGETHGLu9+QXNSnm2Q+K5BjNDtnFodkMtL92Q3/fmcbFh
sSR35Qyv7FN/T22bFZAhy/gLHsIW3MjMaSOpljftRQaLhzbA/WOo521REqhpuRA6
ZWI2vCk/xFBWgAkZ6qDNFI4felvrtkBMBuOE2MO9J2eh4GfaeTBw/eH+WYSDy6hN
XtHtZjP5xMrAA7d1Se9MaX++rD8hUmb4jUDNGLJBqfvyNXzdkdMICNwIQtSLi3AD
SWrPgUMOe9O8rbX3ZE+t9gEOqUi5zCb4zGSJ8R8ZrOWJgNE/CyWbyMcZjT8fInmF
ukU/2pETLPvdjPmeId/3zet+8u/1qdK9oRni0pvz4M5SeoVDEZa+tYmQ6ErmDjLX
XA1ajrGWvf4bTbEKRb6Yzz7EZW2yUInw+GUgDAwrhg4enF28RpdUuY66bSCewmRl
E0nrp8fQoDDHhloFkO5LhWSwnC49WAcc1pAkX63CvkWA53I9VVEVbbEL815L16MG
Nn4901B23ZMBtWqWgK77trO/Tz4XTSdR/NmHqKwl778HulUvyp6Ez75TJ7ZlkGaM
KvDZwZZ5aeoneQKi++LNjFBLmHOIt5zGEZhDqC7FxbIbqo/EXE7x5XWcu2djU9YE
PnzK3VBEPPiASTyD6nBe0TOr7qNnV4AIY7qfofe2nMP7nYNyXTdIyWI2dU93XF0A
Aek1/8bEdZoYN/8qD/rIY3s2gNUxvOe0v/a9b8wc2YXLdIwDzJADK5lCpS9CN9Yb
hxp9GrhCcC1jgpgljWigSxjRsDWrByEqXmGn5QRRi1zSjGqQMgy1LUaa1SjYZoMD
p0stRn6oxW9aHFXR5vaBaYPQjgadk+VndZdqKQaQwfYbzdttob0fwOg9nHEF82Ca
t4vQJJAcEOtzivGc14udZiGjh52526YkNg9DTrvmBG50DVtMKsfR7qFS7J/83o7D
5M53WAeVlY3Zi2lofbLl+FBFod60c4aYvUXgKKJKeXtpFdAf49NEH891MhtMgd4F
7dXoimxbRy1y14qzouDz5SqakkT08KGd/WTWSSKjJcyr1bpKzm2vpnsXLoDoj+HZ
W8yMyW+lDxrvKwvhllSi0rsTfZX2QkU99ES0kYPq0OxJozZYuEdjgEIBplw/4+rA
VuPNDoq1UQEz7gHQU+cOq06XTm5zYpl9DRUWE08DsoMjHNasR1RPGR8Q6mRRwgDB
LzHHXlVA01hxfvykiszdj1bfPWPzm85VhMePmxQkvwTwc4kCIxNAZht6OMhhmdNl
SP7sXWLJvgnxMlw87zI/yixdapBh/MNVbwk0NYeoN2OyN1CuTf6SpJoNOYX3VPkg
BV3vQpPntC0D0cza+xSh2O88tzd6nQHcHpYbw0iKOptH60z/5fG2D96hZpDBvuxk
arQkgPUD1jHmCbgjzxZ8/Oq3D1dPlAYqNtrtp5q8WYX+XczuSnGcUyYZ2qYx4l9x
Ah6rFti83mfkyyQ9khUsxBMklOCSEiZsZAiVf3y+vVBxXoORoVWcSZw1qy4m38jw
oAPtXDw3F3vDzcDNk/EY5ILWq5HoNXg77G5rG42GN2DzBc+6S8X+gt+iMkO9PO32
VOHwDQIZ4SQqDRY1nrw76YFEB7+wYetzleMJKjR8D3hcbr+X0T+H1LIE60/0E1F3
kxTicL5PTXYuM+UIBxxLNGLmUt98EbLy7abY3JbyFi4P5w/uAECQ6ybaaQSNHqXZ
d1C1B2kNcksmQ0d7hFW6fdcD7vbdn0lMx5l0+i0pEJ0XWljVd54gyJnpYFBltogT
gNQCcnNJl76ebgHXzlehSX9KYgulw0TQFDMnRXeDSvMgpnp3Hs9EvZOMLiM2R11c
lf6ZGIH+LXRdnBNkqIccJ8gN2oi/wObYgjEeUKdG9dF6Ta2ITtLLnT1+WMkUyEiG
toFSWRCKs0A4Omr4CaeI+syjegccq00b2hwZUuGyve2er2WorVUFjD4yRhoBnHqN
iTE4BzDRRiKcfGxBoleFkF/aJmwXpHh7Lqd2SlHyfBkIdNn0PW+Rx/0s4ICd3alh
A3QD0GG5ZwT7dz7pCHmBbF2rq7833WG3KYBUsILYQjcakGUke9wvu/pBKmMWMV63
dAJXO/nrf/cVpXnct5BoH44fALtileB7E4VHYa4IQV/ZNKPaF9K6KyvA59cm7Hp6
KuP+vRFWsdEGmMyiVJc5okCL3rz0UQzoC4LivBL220muhTlXL0JoMx/20bSd000i
7XDIu1gu1wwyfaAoTPDX8kp5pYgjvHXPMTKLztUaX/D4ovTntx8Y356Sw5CBny9z
XCEKe1A2EDgR9OubjnfOsG+JxkblOpAxj38e8COFmWF6TSVnA5K0AV+tM8tl1HgH
OS/Y0NfJDjsnbD0iPIZ8YCDaGP+BL33eyNU6BEH51FOtFdrUeCAF/bgfVSGX1qVd
jgb0MW5OZwQYbtOlhVbTVRn4a0dyZdEstEMhMmO4jKSFVuPcOZMXihCLYGyER6xc
zLDUFoJu7ixJbZ8pS+7/+j8l2VSzebzuhZSma/yPeU5ztmGXCRosxJH37ejzx4Fq
8vC0WPEy+D04c0w9LgRyDu96JV6RplMl/P/EXL0x0yfHEBWJukm1b0mYk9TXApi3
YaspObpyyajgaV+GuTQ6l+dAmFuz1QW/3Xep+1cBW58srJAHOBAqTIAVsm5K1XaH
G5bPWgDDEj99fzqb5fQ0KJN6WIQmMdYjgBve7ClLDWR76Z7BPaP16fMAVhq2FR0B
+hArbnpJNABOvY6oBmYVjbUZYW1eUXsE/cn4fkCO5x0k7lRwdEdenuEpWv23DXW7
rSC9u+9tQVcojWF6liRYFoAwdN6YNyLzSrI3bkdOLgcWd9CTJcJFGGYn7MqZat6Y
DiayDxtq3A40F5Qa6JGG9lVHaLoSR/bQDaHQmT1GmfIlG1JzBIivDBkFhJrCEWF6
I5+wU4VX736cJXqZKIIG5uxPaaBRZHRuER2NYes0xCDTqFhjMisuSBKBxdJjn1Rd
LythFrZu/b1dVClVZRqvB90/xZUGwRmmPZS2tCF/r/Q1gXo5dcl7bj3/YeX4FK+w
69J1YbnKgARKuECINCJCrYtf20Jen2wsmcHgOqlcasaqiiHNEqBumlJ94kE3KODI
HsYeTQ1lkuId3n4MVneEGwKmufHy2lsY9ZmcouEsJWEVyecTgcsnTL58cqHkCqax
JXQhnWRdusnp0jrt9O2Keusdkwdd9zKYIBO6MAmgW4vD6x4eHWdWR9ZBczknGVbo
Z1eTpfgQoSP7W6MRmVnPMx5enGU+hRPYuPGQw4PdMYLZ3y5CNU4OuF0rD1mHfweT
eBcM7lPoy4T2tloYKnIyaG5UHnS/1Exb5c4rCKpH0DTpexv6cekwblBRtuWf34gv
aqfT/taWAXsaE4PQ/ltbnl3kjMSnMZDmKYxHRvoRXDI2kZOji5wjmkc9Ub5QM4yZ
CFxBEFdwDA+KTOju1S0KiVyFwCVtI5E2JX5sISQOpDttUI9roqUQtWQCvZS3lu10
ojBJa7rNdBKKUf77oBmojUV739lGw6J9haJ73JSr4rtfZSiGmkrebTSEAkBSVq8N
ylR2zE5DaDJzmkRh0K+sJdBwhFrMLaYjnmPRpXcJUGs6JCh0tVP+24VEn1EN2yoF
pKTaBccfCoi+Q8OV2NEnD9rSrZ8VkvxbV88eXo56E5mXiDbC47JL/PbqpeIi7EGr
UU7l+b4SfTfzte1YC+AlxQuCCJ4kOQSp1Lv+1NhBjq397E864qxOAThm9TfciBis
5VnwIj3XwW7JvckSWlbReTSUSKN82wrdltVB5qUGIQG7gl5KGc7WfkLZK8cDk3oc
CtXNpUDiReMgynbJcQBq0zOsR03PIaklUjkgVej8VX5VF9cKqTlQPR97TO3wNGE5
lEPgzVLesTS+LFxFd6XH1TEoRxSzzMplE1NhaTh+/3YZKS9Pbr9SgTzpsyW5+4t2
3a45Eg7/foMXoFPAOT13eNtaG/usIgFArgUcU6oVK/nmAuw8LFQJA8nz83wrg7Uy
aT55AsS+kRJDVRwpW4U1fXSUwoH/hdS2Y8Cx8n66+N3Cysh6t5OPgyIkSf26zNo0
WP6wddwDiULujWxjcJ/cwlRYcFf5mWJI8lvDx7xbdeI0SoDiwL/acGxe0dQaV7hm
C+6uoJGRAaIJrI/BNvuj3sRzqwPAv6hP+TFTlOXeLIFK45G1xpCNmkzgXyB97ZBO
pbHgHTVFochrQcTaTalc/tJVuqt5SGBWjIoU9tIf8GTgzsr5IRGz6ixWgChIKW5L
frEjH+f2CdbhDiHNJo6do7xCNcND2wNqQuazi2j9RhNEtE5DECgEG5+JZtYZG342
ZAG8TiD75zAeAkXw5hxdwQ3hDXi4SOWVdGGdk/6UWut2HOY7NhpPnrZYzkRte8wX
/RWJlXqD7HMy2T3/9pSCun+YgD21bJ02byPt4/xuH6Hz9X5+xtN1xEPodaw5c5zU
SFuHOWm1pgIkMGFLBbwNIL+JQksJFCIQwL3FGFx1OcEJSFGAWnUhkE/4xjYisHoK
7vnP5PPgcKoM/XLl87Q41mCfMdIZcGZK2vk6tccd2awzDWV2MHnesy7fpPwqfxlm
cAvgq0bhu5afy6MmZ+fBehQP/os7petgd0K4ZhS+kaqROInhxIhP36oaVKS0V31o
QB23WwhjbH1OpEZjlHh8oX0M3IsVYMuC7AmIrKlaItwi7ZeXG6FOl8X1QJ8Nk/hy
AfJw94q2Wl8v8SrF4AqrOUxnUuqFfoS69x1agqLL2MoOseZgUlZJsCUHVdlkbvNE
uAnCX4mc8Fj6HUFgR9z5eEboD+lZktTILB35T5H11ESr9TZDcvjNQ/l2WWutwIfZ
FUlr1oBqJYnjFdZYcSBSpdnOuQnisubA5WtqGtVpnFo3UxyzhtTAe7tT/vo8mx8g
dK7/S4xKCmETqLP2VETjT0SQ0yC7+20Ipq/VPxc6eHsZ8w59iTco67I50hVdcH5B
VMkhNesf4gmC2Q4F/iQpVI3AZmTnj8UptFGCZtrY3LGpbVqqmLRzcCe5oCQqjv2G
H8e8ObCY0lqBdRtwIvPrO1LSkaaghwMOqv7WyJ5B9iPN+0yQ70X5AUnP/zY/Z+uT
WW7LzWsAakIpLofnA2IxXesSoK+hTPoa54lAjIozQUlFbO4xFwHGmt9f6zXvk/yB
yfHu9bbZN08LjY6Nqwq9CXXV39nvKeXaYf1v+E/Wvxs/qUx8ydnLewAKjySE6EED
KhB1hdi27+Gk003Xj7JRT8tGdbrC7tEYRyvLUzBhm7vbE16fF7q3/uBll32ywHub
CGrQIpL4vBChxh69IulVAs4xHikj4ytJUSJaICtRGHtiJ4nHZkiUv0LHnO2BUWTw
bIecWGqrq5lXnwSh8ulo9n4o5JM+8O/3cCgxZU0GTk+x8hjz0Hhpg7wDM6gypb0l
dSULq7x9LD51qpqKzujiSGSPNamu8EPl4gj/aamO48PcfbzHJDK3ySU9/4k7BmDi
CkAuRo4blwRFHpkF/wZ9PDxAkpZQhLN1Z+TZW05rYSBCuYb4VQp3GoABrgAmK3jJ
RDpwxOO160wCnTilPBHkK+CUG+9nFOj0ZnvdomjNsNVqTOpkKs/KZ3125iXulJdb
oDoBh4WVWfaIY0HXuVQN2nVjXvdnjjrTIWZLoUnVA+EqB5NkZFB29Lz7PWQjy/Vo
0nTQWm5oChnV779ljJ3wPzk3T17Qkuyvynu8/UkPqtSax9o+rGzi4mHTl4ZPuvui
gty3JF5ZbNKDnEdNHsXiUCvkcb6jMZEfp5cgvQAPTxY3APGJcKdNUGgnnsxNJgAu
FldZed3uQJX097UI9S2hoeJuFogJJF+Q27pbo/uwBmsernSV5mMqxcbh+QVziwcN
q1WMUNikgksKlWfG8jfib20SJwiT1pa0cI3sC2iyad1neK2wuvH9YWgfMxQ512GE
6OIipsRw29tUt0pwEwRy9U0FUPc+WGfmR3bHTtHjP/9OB918nH5OaKuMB/MpVrme
awkmOP1KdlJIR6513sLTxcxBpLV2eXcgfBPuVestTUTzoS4SHt+60tWP4ynoeRX9
W9SnjzdiTH1NHLF1tjMjJYywEAM4hnuXIvq+H8tm4RJm7FTauC3LnqZ5q0I1c3eZ
rG2qKm7JvY6Ez/W/BEZRbYa2Kk19db7Cpy7F4bC20k5UdtCRCc0w/YQ+AGjiu2Tj
Wu93gYfChAA4zs4VYlPUJjOt3r895N7JGr4kUaJCWd+JrFF6icnWbyIFnBvP/02/
lBaoGCdUI/mr2EipiMSYDZ0VLOAGKqp0EZvTciuz22LlSBbM6z/4xypUygE7fVQb
QMKPFyLrPzVMDVukQw2vm0nC0ZU7/xH17CMiQpZJfXJSdMiPpdutEzul3x0PqGNR
+Uh4hqHauVeBEthP95DEX41uTB7zBBLLaLfWPlv5Y+pXwPbltXhZygvCCqP7SzqJ
mxako0ts/YuxOStsFhCfIbY6HY/SavwGCz4PE7qCIjJfJS5jyxXv+BN/eTThBsqc
zc9QUrMnNNIt5KxShMjrgB4zRmUoe+jLWoWHYbkjt8bDAjHMoXFoeMyVWxG21N9e
/lTJSP1w9KMun1FF4EkqCQAZdp4dpOyelWGp7BLTwV/M9JWzeS2deHx9SZ9mVlJg
8B+nf6PtTZBtKNM0aOAv2i28R8LipnDdvQY8fa0uy+6UZKR5iVG/5RE9XtK8MhhA
2ehtzw3wKhhX+zj0JtUZlW+yllAvvvF4+XjC8Aucj/62poXHxmPexQVdX4YUuFQA
UKXatLhTeSlcRGMiZW5qJfnWwCYlIXs/u1EcIRpI4xOBTeWOCfDoIj3gHF7e2tRu
UBEkbtzXbFPIbi92CsiiSEnYytgKXd9iVebcPk6WP99mkhsOeEsDG1PeL/Evg6Sx
DaBeOtbU5n9PJ5eFHDktvGiu6hMjeGE+//y1w9FPLAsugNp62X32jVImmRLIJlAy
8O2fcMw0AvByC9cVAKrq40GeY/f67I36zxvSpasROgDl+MjegjNcGk6r0UIC7A/v
aGNIV1f0qkxaP9EXMBwmpFApatK6Ue+rUKiy0L9YSofUB2sq7Tde2auxacZ6/Z+j
TkBEGZLFoyVcHJ8rrsE+lfbvOwTRcQl6v+TDjFPMbB1dgSqqOlrMuIjrMpTIiMTf
eVh01aHQKBM65EiJDhamVRL3VjEi/L9bApIUDHKHgkTdtKoeKAaAd4xUO2+maPfI
DTviQ1LfOwdv/y3P9eS9Lk3HjOuKjLv2SvNVUOVDnMx2UKwvcQ4jFgLWvsgE/gHv
7XnFSJ13luMgTlxO5aiDm+64yKaTo0JMa6Eqb04g1Kxr9qSz9PFNEUcVO57NGlLp
eUCN57BiluhYWwSraoQK6XQwiePu+BcMjsjvaqv2kIxS9yIGAmQaS7vW/aMcvhPJ
UThJj5p0KSz5jrdSdO1FC6LsxzQoq66x+om0mkkm0BGo6uO/Oq4N04LC/0yNGYXp
uhnaSl8CgUfyIGhDpLS+g7aaP3M/MsQFocWhIbkLEZ3/4XGD8Us0eu3NZcwHDwZI
UjROqzetCJZaVVE1ZHGmGV0s1rZ9dbp+TfAsOJbp7l8oydhS8OzNcusLnbtSVMa2
v46dn7LBTMq6payq1XC/uHdG2vJNcYN/Q+mvo15WNuhDkPSvksEdSXj+7yf2q6uj
JuWvSqek9AVVQTRpH9jrqN1xrcA9WhYahSnZGlzJl1t09tmm7mdzTE8stH3n5LGy
4+XV6KsfkQphoXIolTbCtp6awXUs6AHYALTOW8OEVi7A+AYIvbdyDijgppFNVWsT
es/wTqGR54GWOqTTIyBwCd5hrmJRQF6y3eDmBtKd8fjx1sbqq3w2YnhG6hn3vCex
WDpkbkk1G8BteJuDwE3UY23CX6r/RrghAXyZ3q8bFDpuRjYnrsN85ivsjLx/Q+b9
NmUw2stgjnAzQ0YmgnMFOlbNetmOrSTrjSeIyEzz2oGpTAK1XCvCJf3Yjp+noHpF
U/BILH0vZTWmpnrjzBYDk8bwqNC27XzfdWtiCx9+MSKllfS8i2Ei3/En0n5fwwct
Cts0PE4SLDeyGZTS85gnKw6cQsfSHu1xXaZPdFB7TTlG0XQ6VYZM+HCKjnZx+/hp
dESH9Cx9rFvPJM0V1tq8y60PtGpoqPEQH7Bxyjk5jOpUohd0u3fRgkVrLIT7KBZF
fIP3OOzK99yzE662ftveMYoJtfGF7MXSyCegx1pa8BRvAKoEr8u2oW73X+eEiz25
Q/SFPk1OXSdJ4atdMDL5n7jqEu6c3NIiRZ45lBJ1eW98FWVYTp8X0WbywsO5RYtr
k3UWjaOj17FcG/jqVLAh9P0ZP9KO7cDZup924oI88xuxd4dI/M/ZcmHHfo3XmW0w
ul5GLZM5DiPfKjTNQFPPcnnA9E1Y5MBB0aJNEDWOcQuEHMMh4KHp93H0NXKJuWLf
8WJqQbeDvZjPzy++E1slI5UKwCBeNzy/bmtF3GTAN093f4F0WQGF5qOrFSDFv+y5
exku/DzeZbji2y9+1TgrAwTrpNXevJ4/wt2tE6Lydse1Q1D3C3G9Xpt7yJm/2UUD
4TY1mFFIWN4MQqQmqHeStizzOyoLHeGva7i3YIvPoH2tw+EVBQu2HHqKXyeYYZdO
MVdb4Ts7DWOga36elmjlPW4uBG4gWa1wWydlhMsk9Hwl0xJ/n6YRC1CclZSDSYcH
y5Knu7EpfOJj8JNlCtE7KzML1bbBC5woHWdk3V5yUIt30EYygIf1YeZTD5aqjCwy
ryFWd7JHG1Xkd7WReJF6jfYSVposN6/OFKWH31kH2bpeONzpLQNlb1Cl/BFQR21F
BK4B2idfkCk41dQUi7rZlDFqsATxmrr/EsLCTxHlVS7xEGBqwY54e30ru/W+qoLR
c7xmIGIQsLr5O7RMTa6RX8c++aZTH2qQhdKK9Od285V1Ueo7DEdtVNj3Q3xht5h/
fqifp8DWVoV8OkxJGRVpkkqxAwB5fJcAaFNLiaY9ppELApAluIQAylNnGa1/qc9y
rpvh8OUj+WhbxCfcvkStoL8BS/WWmtO715LgILhnGQxBEH+neE1ow7ek77wmlz7J
Z/ajtWv5obk4EJ1Aa0jZu9/9i5maJgtnFhCN7O8R1Spe4GwwkG9ibjs/68ZdObpl
2/XNGSwcfyKIYWahpkDx9JM9pQykAElbwut5EWDzEfuDrOiApk4Og6BurJjREON6
5co3nQABzSgpdr3S4wqslTXskm48GAAPRPC0SkPgVx1uJtCZ8M4TftCXAYhvrzz5
eU0xin14XRURghSIGWl3f5GUEpu04kMjvtltAZPOhrFFbGfupje0Esw1eYcPLq8/
qJNnr8YPcTQjQe+PQrUzIyDJ/KO1kx2ncQzprZo1Mv4FAgEwSpi9CChUZZu1oScW
7XYFhs1oGypiIT9ZIwGrS/QUoeXvXCo+W/fxMohorBAN4AdsgQMQx6r74HAZI4tV
5wcEwAuvqXlyrxl6U/C9ororDDn2ENGN4AxcV+ReCFyqmUhBWEiowECSrt+br8ta
CBM5SXMdpxYUJ4QTa09aqjAIjk8dzp6TJIlUAFZjku+xZNC9tpMAU6oGhSCyJZzq
MlaHIAKTwcpDnAH1VQAYlc1qmyslgdqunsDBpPiOreYHKTvGTvktonRXCZ6Zvet9
xLey1YMVA8JXmam85VB1voH0diymJLHH2+4OXYdNUqBXEy3noHeeTEDK3CRBG2J5
EaBGW8MpbHoDwJLuHOvE4sHOx3SbQo9bWJHIvqlSe5+NJPxMTnTjYwI86ZeU+gJk
wMmeuSYsRt/F7GHNTo6ILwGSaQNxsxyD6ZTWEACLDJFJt7kYoOELNZOEzFWS/Uns
kz9/G6F11+QEgNJcgB+I9LQbK8OzYEW8O50lZeWjbv5cB4VqXkd/txW3e8o4NfI+
mjoqEnHCuARCsNsssG0CanEL5T8RsHDHKtW2onIiYELMnkWWiM8KWW8D8E8pT7A8
/TZY3rc1OSjcKwy7Iz70De14gmhyHk60dAKFoM1iY94qyq+EZDqGINJbAekpDht6
zh9wQGPlcw7z7H3htijbNeSddUxXm+1a23Zr8kTT+rZCOxm4Kz0MJp2vJDsgYFNX
MgfrCpijynyou+TlL7BlkXqC3irzy7+OUZYfz3y0dUAxu8q0OH0Z7nf1SBCCWsPW
QqCY2ltM+Zc7SdmSMo7JJKn7E+pHUBMtuqPvTu5jK+P9SuyKR6FwlojhAmShJg7a
6FVeMF796jFJcbylIjAsysyPkcLVWLd/L3OHZZjZK4v/OA4Nj7Y3NBzzb4J8kOvX
J9eNs3nimG3Dp0xxz8IlLJKaGiAyXpoOMKySt5vVCPsLIukC3LeOWG/JTWdff+Xx
0xUuSKI3xDzz1YxORAss+L9QB7md8Z/g5JCOjjy20yJeTZ0M4LbMBLYnF6HIIS8o
VuMOZxI8V6JATKigXbMYVTueTgxMFxcSAs+2sPFz126a1VrfiFfDtv2aplVRWh4U
2CB6stQXDUuqVGMFhDrox986v6z+QZ3MVcf5EBKAyKobeo6uJU42pNNS9HtFRiWu
fN7hkC4gop3yIGp/mWp4uJygIftQkTd0g1oXkOcy2Se0vU1HGCjRNptD2Uy4UDys
ZNp49pyqzXM31RnUXUyzqfPunjd+gcPaHLpznLxPEGgSGMRsV3xf03sVCS+k+42O
7pfS+Sxi90C7QyP/JLr1a1oHV/fEwwtvYF6cUW968OcuTsMwhg/fJFVWDGjCjTBp
Uk1zwmdniSiVdGtjZ7cgMHikgTlaY5wteOa/CwFl9MY5hYFx64BZlVfeSS2xc4vg
6Nndy/R+9yV1MDMRaD6uFNylY9nKIu398GJu7UarvnOiI+mpWt6N9XB6s6c5yPen
0qwrIXhb3/YmLQIjFgMojNtYku9bEg8kG6EvjiLz2fzr7g/DbXax2Gm6AVQN84gA
oje7Vq+JN2SoTDZLFpk7cF5MG9R7E6UFJ37Wgn77JbfWLKIvR0XBBXzJ2i8y737d
zAnAji/OMxGSk/PxFdFLxz4mS6hSAOIhRUGq4SgNU3Bz6IhFh70VkTiZZ4rb1900
1zjP7vr+5LPfrdh/5ad90FMuCGB3xAXrVngWwnX2/C6QDPOGWtJ+7HDKVn5aOwAI
8ib62nPER1Od/NJjMzF38HS3DMZ8BhdzDtlukSbHJHV8YPkIp8iOXfHPRyJNk3Gv
J+Q5evJx/VoKJwJw3p4X8QYXeLFUzNitcjIPjGdcRYbrT+61XM3QgZG2qLkUWMEq
pV1CaTfJ+dY2Bdy7FiH9KjvfHEh2YwTqARyCNSDVub2fC6bayYi05lhsIiTZBaTU
3vPtsxTSiMQYIy8E7IvkEWHnRNR/UJbvjFJF1ySTte0cpH9n7dlsjEEmgkUYK3GV
7VXlgWTafFygD/24J5w7UFt8ZjXOQIT2Zh/dA2JD098oKEeeOR4fGCVWaL8Q7GOp
QULvZURqPpkLCcyRy4aVuNjMUzlyLeuCLdRxyTHvK2EZyN3euduBXuU698p91QPG
gKPmWBMfBWP6vJGmzn6yCi4oKqVS+hI9FgPspv9wMrzx8YUmK6GxsYD8kMIpQaJK
PA8vZDPQzSf1t2C2LKOGSvBJx8GGVghmNQxuNeKmNv1hyJTVG7RmxTPswuH70h88
J1VIy/8KVT7i31YxdHaLy9BDtxr7H8lSCU0HHy3Puh3WBGNa4iKkwkDC0bvSbs+G
qfmgq/aAMk4urWjAT1kXXVHY8dVE3JqqnsMtpBS/5TH68jiTp9xQ0oua0ALEefmx
PtvhPX4TrHYoKdVuATvu2nsSL58KKmfsiUnZXjb+RH/0Xw7C0iCbIMvUhWYGD9jP
+jAev8tCF7NZyOSN/lAPzpShHApH5YW77tSJrhliRtcX7MtA8RbYRxefkM0Zj8Ks
l8TFnjTGNPFPOUol7m6XLWUt8y3T6bOEhDHlL+S7J0m7j2YBIk+d+o4oztxxpmuh
Wbb89DNOlsaitOvApgV3S3FHv2M6NtXSKlhR2L2A0LeTkOPOd1OtJJjUO0q1P2WD
pqnn4pdmsctgabbKrvKwOpomu4JbxNU4IKHTTU8vAFTJ+4W3erubXvMB720XOoVO
cYPWB7tWYwXlSkSQ9+bR9gwjYMktYw/8y5iRh6FBzpxRCk1og1ugWefMMYeG0Rb+
tCfme3bvYuwtAaUg6+QwNjSgEqNIPx5h7ehJnBeUv8fmGwvaeJDT8TajtvbEt+t+
Ilo41AFbKU1zsI9ON+mY+XMZArisc+p1qOv7WtsoX5Fa9y3+sVNTXE3jqPqk+4u4
7bxJ+tQKlYnwCsr1hWeqI3GxKpwyTy0RsR24ZYsbmCN7TF+32CEQqlPzNdeeL6d1
WIJh3fquWu8V6Z7YLNiqdc38XYet3uOvudHaIBrnPqX3tdiW2Pnct0spEML8PCtw
DXiJJlxrtCStaqQpxgzzmakSFECAm83OaguxoOoKscYXZzilYQ2RrZitUS3WVPgk
LJIyMSyIFSCVtt9w9q33NMMzWo9RK0R1x2ofocbTJLrjc05jQSRybZx+NmKmdkf3
1oU6x+p4PBtf7M6BS27rPIwKv1X/F3rBrIWarMm6paFuyuednxFHldwQsQkdR2W3
arZoqhLDSI6fB/g2tmthiD43MVWD40wZT3fil7PSoncu1oaOFAiEUECJm1EIKYHk
iT7WxU5gU9QuHf3jBx/pu0J/YUcaOx6MFaOymWhEiRQMb/BiBGGx9FfHTxXI5YIk
ruTtnks89GHUDrRzhtSzrpRkH0CXVy1HLeGKpjZWD4vudqqOj3UzDG6z97K+biCu
DkCctpsrKCLihUAx9UQnMpRuLeWPoDn5iyRCZa3VKjOQzUXdUywqsXqzeElj8yeC
5OmdUEoXZP8D4NsQjOSy3+Es9DSWmwHXCqN07Fimmo8SOAvsMSg5OuuDDy8dxcxG
QreYjzpqwQJhbEzYx6MwOWbITvkY0JrcAQaauqWXNpqnuu5c3eLu4Z6axXcLUvX+
Bvagf7dSqi9a4p89NaedvHZEdFNJSDQ6hZOMZ9MbZkXaqwupKtVi4ILk3z2sjElL
AfUFZ+2kpkIWpF04XkNeLCBNn+Htw3kDeT418AHYfUmHldYh8236STS6Yqncss7k
U82v1yCqyPVt/97SO4xon6uLpLxR6/6ik33xqng3lrzVwyiRr31YhJ9RyhBrjR9G
LtlL9swKFB1Yon3wdjfqUXE396MpFSVJEVKadwrEx6Wdt8Xm96xa5K37UFAlOmle
CMbmVInyHwc7IxjGIX6dyN0HrIiMih644YwN7OhypZClNlN7U6bvwSZWcrQKX97X
7Pa+BOj9Li1aFVl01Q/tg9CHaHYrvl41P6wOogzd3feUh+WS7fxsrrkdeztU547D
lizLciFmaalUA4YrhlvV8ouyvo9bM9J62ynw+T3mVN6Ee6ZMhDx3CKutbd1YIO8s
PRfkdZPt6yPgfil1NQztvksQuI0r47NAMGqojUyGvjHKNcbu2TTU4jcCarsDr9F4
DYPk+IvMU0Mn/lsfj5lra7le2Xu2cCHYxtqcfGvXxqh7puB9Gstl+225V6Tz8xPc
0uSlWEm/llDyHc9bORVSz1ZDtZVENc7el1DIjlSAyq1lrucEPo6eGwC0Pohqe40v
cSbI1KhCTsxxA3T6UW2alIlV6rjKTtc0GlbRM79nJVmI/H9779QsFUDVDnZWHB9U
S4SeyC16VXsbaPRw5Pb1iIjFcMNQMHP+zUcsU5V86RfhPS9OVSDQFLE/4njEwnQH
H53dZegoJciau0ARnNKfQQ+d0EECPb9+VmrkppDAa9COqxEeTJU651oFTvrWZh5o
/YhQB862mjx6SS1Jd5beOq3vo6iaiJ5OHN2Sks4KecuS6ftn+JRJ8EXUWjLyCRnl
9YCsGOfkEPTnEi8AYeuFpYsm8+/vEmiaZWDuagIRbnK+RxAFYQGsI9naWuN0xG6L
TGrTGypCkvB+yDySyQNA/AbIq0wQNePI2Mt7c0Lvy2wYraznFjyeK8YgC2Hnk4S0
KIK47IpjY9WtUgFfeu8tw+BAgqgQkrFWcxMq8qpyKdFKKcDv1t9oY/oyLeq69IC8
ioHL0oAoXHymVD49/IU+kThm9SkJ1JCH4A7detT3NuUVFuxIW2V6XnrjN3QeZIm5
BIrgpx7worGj5WWo6C3+LyDiwl5BWGn3YGxuEm3UZ4DJq7J5iVwbm9QtRv2yO2LP
UgLSHKsQzj9nwef7OgGItuX3552SKCgROH9PmQOgAlmO+AwBZkLfSRcMKb4WaDPv
xFymhmMM7x7C62sv8YJNub/joGt+jhQ1jHw62yT1wRE9W6B3eYI2XuUc+2Uxqfn5
YEzdnlCR5cnA3xxdeyXvonXWD/Vdhh0e3z/reOYCvVquJE+Uj/HqhCYDIXBp1xrW
9UgwW2R1j1PZ9IuClS7ONoYTB21PxgKRizLMyBFtng4hfGvDT3IMoREZvSbAv+Hi
ootm5nv3tj3pInjIinPhm7wqJCLaFqXEjkKiemxvtg9jMGaev8cCP8V9tRgv0zkd
o+76MArb3Paka/KVsfKL095TGKjYSz3rD4vupeElyxDXMqnUvv3lfYiitBvI48s3
rx9eXk0/6fOof7bxi7Jae9tbKWIv9GLCSNW0qO9/XsNMlT4kCY9KqtgPEyFm2hgF
dcOhTB/wYte1opuVkyfVAOemFXfdXOzBJA23HIURVpxdsaIg7R+Ty5brt5+3kMP1
0UtIS3zS0j0NSZ60UOmioZGk46jnRdJPLsd4r3pVA2GrfezD8tl08gtp3CT4y9tJ
2BwJq4VB0DWEdL9CtAmt6dUuvjyUBrIGvVOW7x0iaX8+MrBeLIJ9NITrsfcBpmwN
HJkEniFcot7GpHPJPKOkUyq5DZjxMtwuCOOqQw77iT5eHv7NP/yWAuWQE42/ytSs
7fQILlVfaiEkE6M2xATkpUJoeBedw16FwLfLqWRrvytfN8dpCJoJg/oI/5DfRfqb
fgXsTyXtMiEiqFLS9rDi6PQutMeY+EW51mJVT7tGAfNxwUhQfgvGkv6TDRS5ZR23
TR9LWWdpHQXnzDoYuXGbjpTsv6xkxcqGwe8tZtPTqsRIGewDh/Ih15Vyu25qlEj9
MfAxnigpD40XvY8E7YJRKMIVDMWgmRvO6iaoSks/DnRHpTs4bRp0u9ookvkztbcV
NEnUa5ST48C74Qc4CrWDrufUJiu+BSLJqtPVUhSqvcFlQBwv1yDpK3ERqOI/fw7J
JxF6Spn9coCjLKlctTBRWEri/LHZ413+FyupwCAlTEzk7fcPDoxyZJSvHtnXBerP
R9mmEVq5/98Gy/1J0e+RAw1H28JQIPqSIciJV7YwTpI0otq4i3z8nsUEudf2jzBc
RFolsT0Hf0grKHM2Z9VlJsonkNkOMtzRmg8k+Z5N1d+U4OiCzjtZRIclqLhr0SZa
PrBk4SapSurPFaIn0TKcW/G5TQO+gDHWVNnKxxA+VqKcJJOSF8a3sgfL53TEgrX3
Yb7T12U0Q3Frz+QHUcIrITVQmhM0yDBD/lWnayW0qn+0B8k/tIuJpkVvlemmJjX1
Wek/pcQs/Pinuwt7LSHfO9up7tJBH6VYUJxJLvP+Q9amRTRuN9yUu4oxVfsO/Vyn
B3JBqzjpAMmIfV3ivKs2DTZ2rD3a7QvQN9yQMW8N1OfKJP0iQYRCUOtfGK28DTFq
WvykpareAx2HAXtMqFujKle0CFKDEQAlFtUD6V2WQzp8G20r6TIMMR2PK4Cc6xr8
cupwgvE72v7+4spS7wkGm4JHPlAZe45RF5WC8Rk6msmLpmhAq+qsNAVo85AsMhRR
Ntns1I8mYJIS4H6bShhcN17NUXzhQ1bGoXMn93KNaVzbY1Ged5tmOLFYWUxco+d5
1UrBB2DqTp6otrQ+2VGH4eRAINTJwS0VoY9OuDg/gm58ZS82EfDm/kjztaPAP9BC
Mhq8EEqM4/xBdOAMxLV0jH21VTbk1559rPYV5+K61mIuyOu5vc+Bs5ldXFE3Xe4O
5dj8+y3U5bG96XSYieyUHrdv7SXqoE9dngjkVjJrRSNA6fnyu5QrN19wIktM++T/
YgfXPSrlwyJqnDSvSZsXinlxOuMLajgxpRclE4b3kKj/WOf5UnDxa4JifM775Y58
vObG2RN7C3K9F7bh3Gqop3PS/l+oSF4GyGiEQQaak7vuif6log75TQG166uhNKG2
uvqR0l7RlJSUhd0RFMyVQxuIrw/ceAtf4Qk1lVc+2wNMmDJI7jqPgJ0yv+dcsn35
WZNoH4NFCC1gR8oKW28KmZccz7RU2+rE76b0gZD1lqmOaPvhWzTJYOH/E+FlMGdT
z+TZPXksqBBaWsfEJRl9XTgqnPJGxj/7VKifuk/0rji/94Y63jLkD2jBh3hdq4RY
sSos9SsqD1Vz/BbZgVjAZRoVOGx5GEKZ2MZHkK7jX9ho4uqo0K9StJvtzhdtQwhb
G5fP6HEWR49aGZe2v6kcUrhPyx8j6ZCjZ61adLTtrN6IlvtvX1DTl9hXnsVSAOGV
ec9/76SH+HgQL8estV2LO8UYXPTx3ecJCsulibJ2bftjbHgDBPDgGo7D6FnQK2S1
7B2JmiaZgLzzVsZDVZkq0KK+3DzSNws5nFtctWwyWxK2zFYm14XexcnFh8cfdSk7
s4LD3B4SQcult9umvcil7i0ylFAlopamK6Z59MTPVgbROvgvovxKr64YFz4L3geh
adoaDsagZjfn6sEurD+9gsaW8oZLgDcTKhVb7mJcBV4GjLCoy3Iag6AOS0SV3zl0
9CeFjfAr2mRdDS42T99Magp79/zrucoG44u8ocmys90hIndZldWaDakDtZL98KiH
DMVQaS4QXBKFb7ZOaj46JGxZax9aEKK5QYT8DmsPqqMCSXgACk1tjMoeCVfcNxfg
Z884IqEV3JP6axDVx1v4GtTs6OfaUPIagL7TXwnnGX6qb1+CbLqh3aqVJ4NHDYdG
B1wJjnnFlJZpcElmNZoOKz0EmNyehdiRD06oPFpuTXdilmsrZ9lrkTo8efbagI/D
cDthU7+bctlCV6I/jFf/FEXk+jDWB4DeQo2E3p2WZdWCcdrRIMvKrAAmO8xmur3k
vZwtkVzdZAXtOMZjsilbaq2b/KfaIjlIx6sqPZaJDq+raSeJyEECFY5f3lX86gIK
OLCp45R94E+cUKEtbP9ahJg1+U/A7P43gMJUXn1pBejklXrsxqcMQgY21rmoJr65
G/HMtsLjIk6fyegUOe3kT7v/L1mWHesIbmhp4afF2EZb4qNd00EnQFcTh0O0jjPe
s60U9eLKGFH1Lw45CXvdzsw/uNgzITv9gNeQ3Zw2CrOF9MH562dC108ObcX2To2+
Fw1wry/fEU/sSD443CfbULQPssczsPmh73XPzWKiQAWoHf4RWneXRTilEMRlINwB
k/DJcEXi0lTOB5L+oHUA9aRIyv+cThTj5Rw2+8+YO9C/075VKxx0mlh6cEpIZ0oX
O1wGRCPjJ1oxjScgLSIuvrgq/N9iEKYzaRtuZIYHqsVogp3xVAAO+tKat4VG6tST
hnBbDMtFZL+pt14p5MRCi84gXgO/PkdzReOaem82IBtOefQKSztgs5LwAUOawUMy
C++RnTcAlhEzMaf3iP/qfgmG1Zw1OGoydBzbhgyjbQk+JaFN/hWqTKOiA8JPu8CQ
nUQ635gc8yQe9J8c7PKH3ziAZZXkwZHfIgwi6mTC/Gd+3mSGJUiufvDPU8W1yPKJ
FoPY1XfCkXAYVC7zQ12uGwYFW/mDjYi3U7+mQRWTTxjvObKbhE4jmt8KO2SCOe8L
xgiQ2fH4KBoOUIQUj5J2mKef/D/UshYej6ExI51U2PK3DNmgrxO3hexUFI1SqGty
Sm++RsCT6R5G8AIN6yez7OCvAiv0T8n64bf+BlrWatzt/tRq3hs9tKtal8TX67y4
sxfaG3wYhDpRGJGEKY1Ap2+UmUAHERC2rUyo7btjkjWQbE5CeRzW04t6+SBTctJX
lu3ODmXnZd0Lezqb2nuj5pWAtoJQRdgiaWkPy2XzFMD2hZlDgZGgNGKfuEAoRCna
gnr6IAKmKvnUEX1UzbJ+YzfTCDocvO32XPAd93G4LUICU43Hhkq5jxqcq4prVCb3
9PUWutcydkCXVTRbTj3k9TLX5vy5fZ34uuIiMv3jvMrvreoqokxpjGL8haKpCnfD
McQoEz8XREeRZzP92kJcjcd3lFJ9VZDwCCNiCboWlXpOWdvEV/KK/mBwuvdk3swn
r9hNcvL/CaWMq8EDWw/dFFWTcLm9TMg1BOKGQSlGDeV9PLLurm1zeDPm7eowTxpk
KD9Qe6EhBV57E32FF/MPMg+Y8thZM43z7Q6JA5dCbhdSJreRxZcH2WstTrdPmmmC
N08KIHSoarxd6jDeMTr+plX8AePE1TjT7uXPqNp2KpzljbAmoMv5zrxH/qvp04Xq
Mr+Rq1SwcwNlTiGHfJLzYI6IlVMS9tc+NX7+ATplzW6YCsGJ2jA95GV1IU0Z/TEi
zZCrKD3WDVSDIFrHX2jUz4C1B1/1gvNE8+jZc7xPtJ69DbeQwMUzRwMaQjOrSl+t
+GQ0F9DJPC3jcmKpudvGQVbTobV2cUZ0sd7XYdLQTsu5xLwpOfx5ddxXK6a7S8kR
F0E3cvhCQhTQBwWAWwU4lYVv7oPMsAGc+FAwGRlbY3Y0FD5PLazh1jVoOX/8wUxR
lJlmol6kYlK7bsatNsFflBKUZK2MPHeeTJNg8zLYR4doaRmm/xjzoVCtGJHhCk7m
XCZa/JxtvXzCwGg9bJgY2zE3Zlyt1CzgzVkNKjIRAuX19Kp71hv9x3rv68aWcKxo
l42jTgRCVAFECK9FRnI0lWBljgYr8wcGZjtbQkmqpCbSBsahqgKkIaM6FB1HDKyp
61MgFlUlCmP7QDR8RM+Jz9IYvm3FIoqkLyxfVD3YfcfoYX92jJg/dVLluypFK+cw
8Q52FkYkdXm9UEXVArQa/GJ7Z2LHYSVyMSDxIsVo6IuzrKqOBz+I/dX31dgQJ42Y
5jLJYqpyEX6YeHVmQOt2R+8LKdRVcX5ZGbSN3uDi0HVgaNPM6iuh0Myp2Q7JL0UP
JnMIHxswvAyDbAcDatKKADTm2tQ6kbtNPHj61rppxgyfGbPIB9dDAiq8xy8YMhef
jv4W21/IUjZ1/6znZ9/k39TjaIYZYacasKYkb9OKBtKZxc4jH4VNPtTFhKu4s/YZ
srSjI/9E4YGxr1N8VO7FutFAuJZsfen9kuoxRShn61/gCJ6MwbkBB800K7P2bowU
TkvB0JAMsmHQG1uVHYQoqigeW/Q6sRgNCQCjfRgqMxX6r/cm9VDqwK+vXunTha1J
ma4IFxidn79fSim7aNEPtodfcYScKtw2B9w9dAsU9dv+ONBvZgr7sfag3sczN5FL
Qe8LEVGGHWSCkZyQELETbxhOc7609YBoePUkjGTD9dEwTND0zI0UqfxSDrM7DSqM
zc05orTA3f+a/pLclLsdSIFOZjrk55heRqO5H48I+Tj43ZhOscIP3TtcSuRcRg3V
bnVwgc/DyR33SoU1xYI8jbBs6sdsmHJKG7DdeSCQ6IpoYOye9UQo9LLlQlCWPSL8
VdVrzdaUBEgd7655fTzGCVjTool89hUugJpp7pcrGrUcG2tvZox/Oyda0ugrGNug
sJR0S9pRSeqZX834JXVS9+6hYpj5EnlHnPnJpjiTDZk8TaHs3dBc4PFoAhq/wz5C
ApjInB8hnnTCEhLUdTtcIoA3Vv+EDUxbpTgUBarPeA3SQGZRM6I1cXCNBq/kaGCK
xbjmvG8N+OjJYJT1qYQKaHUPClOXed+y8dkIc0IwAB2sD0AA4nJOuvB7vwhqQGDc
Wf8bHZD8XezYDpWxa4WEZ2gbQO6b7klCOPX62GI2ws4seI5UJvilE5WgGBGB1pgw
lOZbR9xmz35NIvmu/2wMFj1aIohihWFDPpQ0VQeCRhWr5z6JxaRA6oepqyyZH2Sq
mrCLDwCZF0v7I9gFvo5lj62Wo0y90c1smLoiVrn26aI3lRcIxQxGyExT2hZn2/AU
12+Nn53XsiqFj9nZWjciWfyJjl4vhfhd5i0lnUA4M3gKvEPLit4zlWjtJlnSAZAU
+Elo/+rn2DHIQ95+P41aOogks6Xgr0hDSPUG0xC0TRoQFJyOrFJaWIYKyPS/cGhf
rfUIVK7CXfzQGOwfaAp3DZycycWZ0Z5m+XnIAWaYWL5Kk45OLefeBIsRGxpJifjd
hmBnG1hoM71tB/XfSCqZspjBe8H4y4cMmS4Kq3Ih5Dzjka29lNkAVhkzbglri809
7BvoxmK+CUqe9qvl0qpoSGH1Qm9LMNUV/NYFLzh8WHCxeZkW2D8YpXGIMeYEX9Bt
r6DrSctqkL+HZwnMbuaFNKgFDxXPqcm0rzUizJA91zSGrYSGC+WmsvXrsjzLY4qG
VxUeHQQGUziyne4MymBbOUV4rUfSTW9Loo3RqWELX/OOUSG3ICpz5hqRgmg+oaRr
Ta8mfvUz5/Sj9fOD9wbGCqXvDtoXYSvW9Gfw2wAeC/C7qy8SOU56f21LAZbNUcal
lrYEWK1uAbGcogQ/gybuKAX/NuuHy3+Wmkhra3EJKNmBTm6erUdyC+aqLsYMme+Y
CxSab086HFvYa2AtCL946Wfcv5AgzNe8Mv9wGRgfZ6BSA9a5kUbKFeMTVtlJozox
y7CQu2YnY5cLI6jlfv1aBMW0QrNLevWJcZ7slZtfTeY4sH8Jj91BiyLXaklPzrEy
Npf4ZKsQ8h3bpkZG4u/BpaoNRqCIaYfskUrMUU7l+vabdKekSpsbuZ3KZejBtCyL
7vxrGDEpPhPDl2yMEOLc9jtzEpgo+T/8FHwOx5HJZMAD2O5ScgXbnZ9VPKnWERa2
JvO2rpz9eWTEMH7go+y/tMgLB8YTzXIRqe1fs+mUH1nd6xTSkl1AcCCHGGsVSBck
tmowpRIX9ep56pSYI0JG4nWOtH1hj0hfSLZi/LJO0leQkKo11WwW/9B2oPicSDJR
6QVxJyFQSL8oH3DgK1WEEFokIfon7O2IS7t20AhbpmQfKcQ2OKOPY5H8Uj4qs377
1puxC/r52PAYjN7GPZC1sXvzc0mrw0LlpJfwjBP249oyoTtVl1s92BzxjwYE7Pr8
4Nwfz0lKrSoJL09n2Bthnxgs8jkt1mn84bJTQzHpSNSV6Dx10scKzlfs3obrKUMj
I50rdQ72TorEZrKCGmlVOw7/6bbbEGCfaj9UgIneuxZ5KTVFEy4XI2RujCuaNn7T
+UXTwxzOmtz+nmtjrK/JEGVXbU/bUdoPNmvthZ/VP9Sq5CRf8y0xPpDOkKAGiacl
IwhBhyr3ZPUWT6OU5mzHcE0Q9pAH4GZ+Fn1pSoJGkdc58tjABHovt1GEdSwmo8SZ
rGTf+MrJDTYZMWJM+/z1KFZCBFmWXE7pdErQMk/64uT02lo4dlA6e8s7w4GKEtOF
42jTQzMIoMblv/1G4fOAngOSgWeBG+W+B1Q5iuhQMGd+TcY84HfrKVLd2Glm7SSz
xoQpAkq0mmujAJSS+wfc0MKDntb+nUXRevwAdJG1R8zbkC+14oYmy41CKieWFuEt
jdgUnIOhgGTUtBEoykyGmKtHCLQjxkw63DskysZtGP/1wjk5JvcrjAN/jjNTHs+w
YLNXE5SkaBPcLq/XzwaOJkuyKT9glah+25EqkmhRk9Ufrifu8mpxy7zxkT1wBizv
ewclZjgjTY2qtNMLgnPfShJB/bhxyiXLVcWUif48yK4e/rgExireQsP7ZErqcyC/
afcajLf/Q+kyyJPYZUGFPxxPt3F8FAXhmV16q2vctul5k0wxyq9SuYby70WvD6bM
OamAwpXcTDSgdpGt8Q2qTeBpqXiG3/ALbReenZq4jHZVs/3xJvdKL8KT8vf2EBdv
JPKUcG8UY+HOIIz2NliWhIY1EA8XdoFEpCyDlcNSMn3SUVAlbrgnDcgNA+QomH4a
/o/yeStxslRWJyaDvsjytNjVXT2BMaAhrmcKEyOJFzhuC1OIaMbSqFAV970Sjm+t
iGe1SYT5rK19IT14IA44uz83yVN9R0uwPD420APJ1XLq+BvVigXe4UXT+9IoFML5
UQ6doRAUlP8ACaKM7f3lTwezRqa7PVG2UPsxVNQ4ZcNYOASFA0uQg4khM63KscDm
byaRXTHdHc2hY4MsbIimNVoYdwv+xM1G0pQZL0IaA/R4hpD/eki5q4B2Qw5QDdPX
85qyiVmfWbEf/HKwKwyFOLzlkhCx5i/by8B+6d0EC654TSSia5fRq2Tg7qaGqhDm
uahk35GG+j8Mh+eU9w0WG+e/ZvzfOu8lQLs/qzNI8Ah2s7uUr6JsmvL6cuy3HSiw
LhSmW0qADzbFG/pkKK/OFDZFkEUeRM3f2MmuJvD9CQWRz4OUGvfoQBg6Pfu0z7Vk
PXaP/HcMwLDb1xyDv1crpm9UcOK+WCgF+CkWcmvgxp0lHjY4GNj1Jxj+odWqlv2K
wFLAC/JfDX6Icl/ekFPxaz+PFDXWcKqwCME88wcFxVEpF4kTuxrC+YtBnB05RnI+
SL4ZrClPSK7QaWT/Djc+AKiqwU1WY4HI0fm91NSvcuuPnDYIBcN2g/yWVU73SF6Z
XSdcheqrRuxmO/tFMqYLApwBOAuLTI2tcftDVO5TXfOOZkhr+4sO2yuSixC61dwY
cRcMQcdI3jNJ3eQrqA3ELUqVDkvk8fSZeRkOxQ7OTG/qc+X3MAZ2Ih8I+9tXbsjj
AUVN0DKKy/4GkFBMX/lm5OfHZc7dFneLG9OgL9QM0qMBj8AxGJqVJMERtg/mrvxa
LWBh0ES3+kbmdIm8+IrEjdwBoX6YcnFOzJoLDRh/RVVFxq7BfnS891VDV3y+ONvD
H4l1zDAU2wEepXRv8Ei2JUkJYFZdvucn/ndDSNtXAVjYCsjd/hwXST+M7Glo5oVv
oQIax4iBlMrIBu3W1t5D51BEFDcji+uHflc0zAyjnBIjBxUv3V6TufGixma7C/Fv
QS+VmaiGYFh1nruK3hZ6DrjaVQs84cZe/EXjShQuuQoTl5QS5lWjtmP3v3DN78k1
3SFiZ+797+J74F+SD0mSRS65O5Y7jpgxMn04XCTRhfWUd0ibCXsUP/5nD4wQACtK
EYljMlWoN3hVZMdi8pwx6ezFDP/IgZUnt50Wgoums5WWrp5icrBOiOlGq6YxXpBU
TJGX+TUnEGwzcTBkLK6FkkR3YStoxZ9HIeWoySqVz4lAV/qeu2EAxoZPr2mkgpSy
+zD/y8LyfI7GQNhgNvHpcaT3UeGlJObZLeOfgFsWvBdhNcmnY9Oxw+N/kzY3GeZa
rNt7/d2y/ol4iOthp+tLOhQ2oizURk4KE183avVzMlAyeDB7NuUlT+6Qm2X+lo1/
lD9XFYPuEwb5pOIqYn66o7hJJRn2A5VWJ/CrnhBtVCeBTHFzLpAiEG6QUAw3HC5t
qqlUXe3oPmHP+8LNLhro1cbe6H6t7h3ICwvIUtXiQ++MUMKUdF8E29P4SyLiMeCM
cqUobr+ev81TST/82KBxYuCr9pRYayLEcrc5xI5wGtYetqOjW0hNy6a2pxwElnn6
p1dwdAxq2u/bFd9EcBhHZJhk4/J2hFFIHFfVrJlDy0XWZ6Twh/soUmfotPHjwI9P
ln+pAcOqk2LlEWK2Hx6i0ulnDCGEkxu+ct1pb39CZ31IqCm8tM15xs25Up+XlhyX
TnrkXhGxHquLanVMAJlhWAm+ZBRWiJUSvHp5FANj9kqeYHqI/jdjDWb8YZcVjioi
JIP7VH+zVX1x7c6eSdDAEjwT+Qg8MCv8FFI3L2624rGMsttOlJiiw1zjwhQqIx1L
Mib9cs5jNvn+vy3bO9tWIfjklbhpbgiSo5ktRjaY8SbhWyCNapZv9o4r6B0VkGru
wyOROqMz7pui1N3+EoUg9p0WiSdFQHdcRRpd2GXagyBMo9mFXn54yKUTKB66A+r0
xTjfpVooSToHF6wDpcaFpLxq62KWFJG81eLl/utInBFiMx9yPouqrugoF16qECFF
8yKQwPbSYp9O66mNBO/znG0SP6sYmNeLRLWKbulybMz0mW1tgjVkbtTQojmrkste
3HwA+Y+Djf05d0Xe3EzFE6MP4CAZTzuBqjsjBF7xmwZHAIrsW0MYxdfPyugougQy
3dIslp9goikhglTuzbJ8lpGzyAuAgxHoaLceo7LuxoNe7s07o+LLSmgEjOZDZIKn
A3XtMAdTxY44Or8SZKFlaeoLyb71aGiQohX/9Ujf99rl9PuNuFWmgnO31KD2fFyK
PIEojjbO7QMsGoO8RqXNetMMNK8ZtivcKIRrgR+Y0SiuFudcOI835AQ/MgyzE7Zl
2CqUIB1GBBRuKvhRWP8v8cHchR+juJw9UxYKK/G3RTEXz2niLEuyCnxTRoF0OTBQ
kHmPUkWkj3bMflsXFC28/sTkRbDc4ULP4qi/pGfbA+KrvocdoIpa0HK9KI3iDIs5
kuE1xG7FX2fBdwseouJRm4hxwZcgrTOAf3l9uTgUn/eg3sz+4b9mdOfNisfj7rwa
kAAWicRu0JHyIg/9koIEuVoeiuFilTTZeVSqcn8f5VXahDCSRUdtPOnSMk28XQUh
z8Wue5xACkBjZOT60m1UCTyBTIT3Pz21oGaiCdvRft04aALAMMPYWgEhEgmv56CU
EJs/O5gbUAIlBKfb1wB7N8ofAIMxnY8sWpZTWxKSgwZyczoUL5phAOYEehQEM/1d
ektgVyfWil0AaP6OGYLhz586SgI34+sAygWkHbOqrEvUcEuLJbBJvsStNCODC3K/
ubg1V02DQb1X0MuMBkr1uODdARyCQVvh88fxyUh3wphGESldRhVoMfH7+BwA3nGa
GXN+MUsC/1Qo9dd5LRDnXvJJgc467zOCh/LHUFFmyCkU6a80pOnsHRmmgQMbpog9
N3ZagR6OZGqZTchByyYDdFARmBIJsiTj8eUC9anOVbU9uRKCVB7Y7vq0MNzikhxG
JOOfKkUtw9s2k/uoq+0qMN0kxpFn7hhJK3v1Z6hhjo4Zy81D08eC0ocU3Srpthjx
Jt0PDiAAHfkXJ+aPMPmF8bpj3ixuF8miEDFh4gcHPzLkB/7/5ljvDKHu3rB4vbph
wEwbuPsTBksKnZAZVlW5K/S0HjmPLsIFt8RtP9CFWqHSkEKbj3WKs6co9uIXW94K
naKjbPJ+UVSXWXKAS3bAtut8AXQS2YIwp+/X43Bxe6NkW3xtzWpY/HpYi1go3gSj
MkHlz6ZehcE6kPRbeq4enCqM5OrAZK3ocqmsrFIv0VE/yTSh8OU3MaYWNqKH0jwf
x4hTb0Dl4QKxXoFWjcp1NJHMmutJhJuWNcwI3mbwJcSDAPzxVPmv3QzMvz0axRRZ
oM/Fe7jb754IjrqsSqpTt/XqtSyiDvJm4yYmWJy6YxMm0rSegPGhwgVcQEJQYDme
zGLYh6Kjco3FDettH1b0jFGC7swqC6OpDWoupJ2rLhPUSmg57yLR6gZ1vikr71d3
uA7l/++wCZNuItSPlLSiTouGdTM6jaR2cuxAnSjlqOCt+7kpMiYj25vAw/J+Vap4
t9dqVKLOiDUsTnTa6rthqN70LbzWG2S4wUkO+Wfa4ihjoAGN6ZVllV+gza17g50S
17M8I3gzST6wp9rfO00sf+ItVViBj5nKUbw3jsKPLC6B50m6EmGqMkLRDk1N+5aK
Op7+Y/XijmIHfh3U7Shv9nNEpr87preBDBOKBRkJERCYxuRb0FCnukV4Tdayecv9
WBVkL/jimsDnlbphiKfCoPOr8Q2xcpU7ZSMaeRMo7eN9OUrEa1CTcgoQHJ5XaeE1
saLRZ3L1lTDcV/5+UqXAokCkgjcj+FSTOKJcqJMho4PXwwRz2T9YYv5NcdJWbLMl
7b+cDZ/C3KlnG2UNwG5GdhnDIySIUCmUZS9sidelUIGMCzWVYQRcLRbwi2eJSzVZ
GKHebTDfAIzVRgr9x1V82nI1xZBKosgzA97l6HhAxhlEQgUw2AFi4tbQpZ+FO73t
rtCtsp1Ll531lXWE5xD34GQGsVmDNelBxaMYjzbzYb96G12hgA+zhBN1a4bFT2v3
FOlKC53b2Vo5NSANe+22s5nKpP0R3Fz0naiSiqI6zdOCIXBVCgkSzHBlfRWLMjc4
ijByoUC8WEYDi5Q/Y9wZmt+lxbAIl9ZOmM7zkjBgUqzaJYmt1zCMoiE3/fTfsPjv
IRbv6hKu+4zpB4srn3MsMu0CGz9Gke6M7sjLhzSRhljWnY/RQYxrqwTsJ+F+VRMO
Z+j7kHKECvjkT+5vUIiXokCkzwIRbn/P0bo44Nfe9JJ0Q77SLW8iu21OugLTUhOP
nv6cTmbIz2bLqVNr1cMO0G1KkaSoK2mo4OnQoReggQcoYKK/763ktUFR/ViukfXp
DvtU9QUS0l82qCr4vVUhsBZ22N/YLckGYXtpr3aunq8gvMASxrvNcIkaDDMCAJs4
FkH9Fb7TjdtCnNxdTdTQc8RobactmSbF+C+w0PBhPCFHiWr3LXmWrHYs96MYFkLp
ndl/wJasyjKn0D0fITCFnXfYZIoBpIsfCEad4SXDkRbb8fDc5kwldu7vrGRCVFhB
ntSbOPL1ZwBAPynqDzOtrF0/z9uDeDvOQKE4Jpm5U04XMy+TxDIfvOidzoZ+rDXN
94AlpGUnzpZmh9RkWdKrZBzhabHe92b9uPcI9KaevNq4mUZxxYEK9bvcEG26oqZt
ECf8xOAOGyMlUKdhIsc2Rre8VOfPT96Mi31zfTdkmv3+AHsLuN6Sm3MCo577mYBH
HKZP7tUMI3nahItHg/Yk5DoPUD4aK6Zh80zw2+2jecrY7NuaeWTa+MPqzxWXMIoI
+8mcXzjCeClbKYF9BrkqgFf1M5hJpjjC+ocG1ESOVMUjo1mmrCe/xzJFDgRlkDv/
DJcP9zWmjGd1pTT9wBl/yirtRsqyTHyCXrVXXFEB2Aq2S2Aps/9bxjo+IskE3Qz6
vzs0uMp3O2ieICifKvsGok0Qcn2po5okN2NDosrvU+CiJ7x04eNKYuILTZKyj+3c
QJA7oPA4g6/2vdOw9EU0b8PKz1zmUqpZTQ2+yDDZetnj29zlUja0yKkLN9w2gsUO
DP/sqLSlFm5BBFKaO78DJmMxfa6KLIHHQ+4TinDjrVqsnxbiEe6R67o3K16PqRT4
NCtSiEkqLacX9RASMqIN3wGfQvuavmUT3DL5LH3JklmxzsTJxaKYQhhkcSFhnbfx
P3KHmmCsH1CZOFubw6+E/iSg57slo/RCGHNprWQrg8Zyf1KwORJrdBRiUYrRuRrY
zYFKitUNDhcSemCOJRAbKHfASpmLETtbgJU8j87OjfyDW+EjKByKV2ERHUMrleaT
bdl3rCCTo2igVRikw7kvsAtcwPNcDVa7GT/VQBBvSOV8mO+oIlOrRXPenz+hKR2I
zIXsZ4ZKIzuCObUIroBuhSnOXAMUTnDBO4NhYjSTH5DpLENkMntIWN6wl48OiPoc
zkpLgfeh/Ys51mYcQ4K/0MVuKOyOgK7z8DSD84lPraX17QRf0SgNXCkfEpFo5M8t
qGcV1QQ9nvJiaNvGB+s3TuHGFnZHZZJPm8ePl8LfK/8lbjO9Wbxnas561jS+lwiY
2L+71kMJoqwPRxUUxd73gJ07TJcHvYMjQvDTosmlOFmgQKjVHvzboiBDl5zuqjD9
+3SMLwo5zCEuMNRGH2CnKZjSMMvtIcaTR82Lh+OLd52ijU3k6RHiTrqK/uzkL4l1
t9iB1aEUuEVWiCNDutuCq6TZwGsZAneGrnpEMF/vjW8ilO1c2VWJlhq8bl4Y5W3Y
aARE15LXqOv5gFbeO9Vz7zMZyNZnHwd2/BA2Lca1ZpKcztC8lpkMhvkG3PEa4q9l
Rf5PxnCJNoU7FBoAm5rTIQWBBOO09rg7ybxH6RNkao+cIGNaP1Uroyd1K0aW9WUJ
ZggsGk9EeNq4nuZyw+doWf9yW2e7QnEjox7txpvHJORTvzrcmd3Ezt/jYTUvH78c
idpyTOSvxqkYSjSwo8TKbfqiNBPmH4u5GVeAg5sUi79JFKMwltVGL+hxqRrOqj8L
BPOug47EibxYaUXc7+4ceNz8w4qzjGBcmiCgUYx18xkuDfsFXk05N76VyKYQc4zD
ilD0FBt3PvM/wTmcwYNnBXnXbs5YDfpGrWdlWEf6W6Lw6bxhAqb9NIJvYB4krqFv
pE05km5zg3RTUN7AGNNn5BcLoW2snpJ7QFNsRBivCmErDXWCo7HSUaxo0zO+c4i7
jnw/ysXtNH5q9UafRzz9o9ICFWRH03a+LimzFlrFqNIYF8yZrmT4AEHwDBi0o1vG
KSedr9jPOrd8nNOH6UzaUTJViWNhJ+T+sx1m5PayqTChrRDaHrE1G8BW4xQHoWEv
ogvBgFVUO+1rhV32oHAtZe0gxeugKb+ck0eRVtW4+WkpbyicfTLb1pn2R9OThg7F
XVJcNStZ6um8zAf52OOCScAx1WUDOpo5HycwgVBztjZunKcwvm63Dx2PKlkQ1Y04
rYdC59Py729nVF7pemp9MuD84JlNlc1ovCg9funtYIx+KhNeGHjtRHi5dze0D4pB
wC+byna3BkcGvWf4eJYO5WAp8DEhgI/HBN7txl5AtTBLFdXKMMSHorPHwEj+nHDn
ypSg4M1GA0g6Wa7z4LzbcMt1bWrIFsjuVzEjHu5Y/OJHn0Ie2F2jog9pSHudGMrO
+bdvGXRh81EdPPkQLnz7t+4dDNt+F5jMeV1ZjY5tSz+2ZrtB8np4OtFI3OIVmtsP
qrKazcw+UfS/aNyNBifKBIfzOyAYC7Lf96qe9/t7itbn+Th5X/sZc4yFbSg/v2g9
Oc18maLXJKWsXXIU7qqTDN5Lvo3YKMehv9ecO1AUP/F3eYs4sKGcqOFN3Jpb9vzW
eGg/Nci0YvOJtkkcziXFlP9E66mTPs45KdZI5CzuBT1QFUeplEPhSd10Jl8ZCy4V
M5H8qFXS3EmBC83PBnXGf3WtZAfyX1YbyzwuSCeMAnU/f8ZRFf+WMJqlEslWV1ru
RT3JWeKSSYk07nyZv7aB81PcGa4LslAvo6X79qa2Jd6aXPPXocI0fe7Pkk8NLs9m
OJPuRAJ4P26WkJ51GuOKy8BbRhhaA6zP+4L0hcz3HPPoFE+ERQQDGpx0+na8A2to
y3QEd2vY1xFmqtS8BwOtBaZn5gOwhghplt6openuJw9toyOtaEEtzn62RQKDu9sQ
sGhebVJsBT7cwYF8Z0Fd3SX817DoOEyVeCQDDV5UXvKbBM63YfsqUvxZOR+mO8xu
fAAoBoe7Ia6Msec78J25QUBGdjbxWXJrrducNM/PyGY8tvJJAZWCWukliHSFC5sH
od5BxmcFtHvd2qvL2ueT+bHB/YnjTTDqhjtH6XH+VEZzL02E9gda8OQCpYgaqdxe
IXwYV2NtooeU1fsjJHNVGZt4jAzBWDW+/74nrvGGQkPAFTa/Jb5SRzL5uZ9bOHRy
F+uQyBXdktC5Ev9fOd/FSpTnqeLwadxRXIVSpzCYXntY/BS/mUhpZG6q8iVV7Pjd
eWQpqlR25da3cGhHck2tlTchAc1x+9Bl4jSxcqlTScIg1BOyIVy3vJJoJk6IHtFQ
tDh4lnrGtiOPc3s/rSQrPRTAwyWTlq961QVDy+tuB+PD+B5q+KRpiqSyruIdRtJ7
caOh4UDxGitgk4ZPHTaEIMB45Ic8K9ha1J6IIv3ci3wulg8F/C2awQu0w9ZrtpOz
YH7UUm9tuIj5qtjkSx1TYp79ilykI4yuFzbvQHptPDYmstexzemRXnIVIv7S9nLg
B8u7UFr8udKbjzusrNmnlR95QA2HYkrYT4oYFFnU2lmviAvtKDUkMk4LM56ivJx+
TwZPeBxGbkyyBYaLmgArtHtFRQkut6lCLU7glY3lgUToUolIcHK73QvlA+9PLTeU
svhnLmtYDgI4FGwK+vzqL7gZtWD3e5xHcPL97Z/sjLqarbb7JVBHuWDPOw7a7gEP
6kp1exIbGPavFvmHlvhZJmcpRRD9RfPjI9voXVyLGubAp72wjsFYp4Da+SEDFY5e
vcYTu/kL71SSlI/S3WjYV2y3udYDmmgMdR+/aqlbj/l6Hi2gEwNqrxOIUQ2H0OQp
bXmEgObJ0kKwotfEDVhOIkYb7P1Ehvqanpsy0Q3UQ70QPNpp+dYiYJxPJyi12g1n
bGhA9bYluSODS6ch+KL4fn1IzHaUyNGg1y4RZsuovmsk88ho5Zd4VXUZvVBl2p3z
KTf3lpKhby7Cu9p/8BnaqT4PGi8uIOrvs4OohgH74atZpINB1ZaDG5WJnFLzK1Uh
c9q8RLfZidDOCo1dnF6GUpQlUHUkNc0sQlJDwiQ+pyZODqWuRxnLnAZ3Gbn7xtVA
x6dl8SE4Eum+ef/CDquaFeiPKi38NoL9VpiDVWMUOdQTcfMwPIrLqO/iKB3TfqYZ
Puo6I3EG41yBp+GGaKgcMt2Atk4sL8irfu1kGXW1Pp1McvJDKuCUBzNVXHlEqB+/
snkDa5OPi2vx06u94uTNsrkTgP4UfAYbDrjOsaY4wWLvLm3Ep0uNg0nlZlPfRB82
sHQ6eii4eDvQ9xBcyfXKqNgm4Kw0REjEGQyJw17KVpCwqj+c/eloAz88s3PiBKcU
otoh9QABXgoGaw2Be3WyWcFnAffOB71Zj84ZaYCW2CNc5wrVJekkJjB7Qrc5pK3+
FdykaMTzjcZ796IKJ3mONBIZSQ5Zj8NraNGFyw6JJGqjoN5s09S//ANPmCdKhCBr
Io6WDtELSjmgmEX7UNpCPacTXCpvXvdgOPckxqrIhvWWM0jC6RCL1OVvkGLILDz5
8EPUZfbqn/nkx/+OvTtqrKiqwMrXam/zE/03NMvnskFoOL9toD+d6UrscbHbW7N7
QhkXQVYeuuAarLgL/+PJRFN8T5rBCW6Nzkz99S91+MWFHyVdjG4cJ8CSJwOkJWnq
tNNaF8jSGYqyKNT0IaxaX0f2u6AvC88Z3HJIdkdKoWLlzsaCwImmxo3JYW4llN/q
4nEBnJDLQHwBlazkXrM+362w45trJMMJMlI2Gp40M1qY8wDW3/5Zv27rg7jRdEHR
UZwqwWCJ8DqQ/Y4uWraPYXbWDnnVinGzcZneGVJZpJEsClMjCT/VeklkwQN2/z/+
qzTLR6TQKovPEC/BUMXrHjviPgzyEHwc+DP12RQPktbTcr7H8s7perGPda9tLAuT
V3VL01+pWShCyAqh/fRQXlpnw/vkH8Dns3vL8dWh4/SDnjkMeo3HO6f7UK8+9lE4
nj12EXexi0hJIymaPV5bk/g++/BB8O/7hwMG1HgOdF/Ln5M0V8+ngQVsMnbotoYU
nSUV/9SwJsaUB/RU3GMNfbMOWI60LqT6LL39oxwxyJGpgA1O7vcXNd0+TAN+s1g6
DO6g+CxIw18JyN2RsL7bMpk1hK3un0hbMjgKXXT+DnjYAtrKT0dtfMUS3XmuWZPD
eeLkVLIz3gS0Dec/EjjbN2tAqshosYIuWp9JCkmkt25kpPCcBOD2y3s2NaazfNlw
k6gzY3tEnqdM+xwgppDbZZUjxaEvLUQ4LuJb9YOjmxIJdYypaE4cjP7sj6pDUK+a
ALiUDEwEi/tWK/SGX+7Xwj6fwVGDmo4sM8+Qv2crXAz+VJlBFaqUtAeMnTsPveyD
ZEVgsC2OMia5xlFBo/nYBrHGp0KBpdOgw9DYNgd3ZTDsOm/Wu3WBiKi9Aa/VS52G
LdkBILKZoCCaT8E/bLWyYBefmlFu2rm49Yo48yaPnwZiY00Gr0cTvWYqyxE1oEUO
YCDaD9PuaFQv+VtJZVS1YKPOFHzodaO6OYRJVBqKXuyEpVa2TtEw0cEYJpMI4t22
3VjDcVskhbNswhywVWHaQW+WUiXc2BB+oiTsOJqcz075nWzNxQ5MVTN7DjAIT6Wx
6fEIj4Qmv+hqIehw6P8d6MgCuMgsytHX0ixFpKtZ69TDySxCZzLr0hG67wYWXY66
oc9QjhkXBILMjHYUK9TTkEjvekFerv3E8bU+mSjTCmozj7Drik4jm3s9uMOumUNQ
h2MdmHzYLVuxs9UFLLZdLGoNlHYmoKKiVKk84FuCTqNudJ/MpbyZ3NxVjyd3wWRj
YJ7EWtPZufHQBnotwXX/sS3vOpg0tdMs13uwvv/WAz+iFA35OV6DPn7GdJBQBNM5
fSAmcqBa1u2Lf/W+pkv+pJUxzVDATlcw7+lHXIgg4tMzZBFipVf/wWzbILkxWbtd
O2fpctXAFXdgDHK0Fwo0kNbSz5iJXJlGfpntRK4CaVNmhnDMRUp/muao8IOB283A
I9FwRe4n6U7EAKlsg976cggGRz96oqN8li41rAW0bGPNuyy0Ycn9D1dmZq0lNqR7
K7LIKHXhQLXOfD5Ukl+e68Q4hyauoORoU2G4PuAYPfn8kxXae9Zmw1oEc10Oh5wh
T9ftJj2fRfSrQ7kDmIrZxcTE5CH3u4MaG2RVHm1p6ScSiWlt1OmVmRxonGuecWvY
hAAvxw6DPS2WFguIXYiQXUtQXn8D63nVMitEkYGTL7tMXbEViEyI7bj5KwwhuaTb
buEI+NKyV823Q9uD6f31PXFyezhBZ7PsxuPiE6FQN/4Yx39nOYL2BsFmFBlj7XeF
hOtIDLeqsC/W0eQJNMK4NVEL4wZDddWWE4wisQFwFaNLCSu/AyaRY69iE41PmldV
VZorPTYsbctSVWGc71ADJW759P390HogNaMm4tJAAvAAJJHbiQaLYVrXN+eDW72c
K/BiNcH7eX6XHCs/2Jgu+OFnnHD1l0lcmxMdFTjuCAyH9/GR1vsiZFlQfFXyBQTV
LvA6fw/1+cPFbBMTtjC2gf7w9t2GDptJ07OtrN8a6QJZv4Mrbfkfmd96Ljb7L9LN
BAkB/3MBFyaIqV2ZaZGg72VNx6FP0AXGPB5DigJPw89YrXSdiWQHWNOJ6g95xPpc
++h9Ju0DVavM1wVkydW+K1IwUMI+oqOEYg47/MhBH1oh/oEYm6qImGVyCBerKUT+
/+yBxOk5JDKbi96xAHYHj3ptkDgkzf0+jb0ZxGhCwFFTdeIDIR/tD5MJJFPeH63g
MXV89fo9KaXls+nGmlLDj3+nXTbvvBnQpwb4rUUggONghbjGYqkMDh+WWOSvQHQc
nAb+i0Yd6Eo+YcU033yKdqCjV0NUPlQWuWi5Qd+F3BUdl1bEvCtUwH/8si28YJU8
dFn6l4ud1DJLgPfDaWV0ruRKGcFT38685mM5i1BbGop7t7Jvtnk5K2eQ6l43l5g1
rcHRFmLRt0jZWDWZC+nmDhQtvO3/y5rx+CSbFvNBvm83sQkwEKNmTTS0Usc/maKy
x4amii+SXccE35dpCOpcxa6y1rjFCDx4S3jKKUNBUvdbTG/T7CxyNT6pZFaKyDkc
9tHlDsYCB7H0I2vYje9eV4oiZEr8jFiNMjEykmPZKpVJ2s6UXWt6iB4PU4QOEXpg
Ib43/ybNck0dYrnWaOxAvJfCHzFX7z489cA/6wpJqFRqJn7BE6q7XL5Lc9VxNTQn
sqy8z+2qFH6FDoZfCcAm9wKPhsIQlCZ0mub9qVfIWZDIY+OXbQKy9yohyIot7UaK
RKWlS41ySIbh07Gdl3ER4Rdkk9yJ6gI1NwUONtCGChvX5Q2bZJbRq0ahyIYVQaQ9
0O55oxnSqJwSaax+TvuIa1Th4b+QW3k69h50ZMRpHjr0gEV9T0PHNEXFiRDjPkgw
kEhtQx0KN1WwxlzjjIgSMZjrdJ0Lf+hZdDZpqYPCn4dKFFCvNeIg/nSKfPo1sON8
/0/abbXqCESC2Qd7rLJ2P2CigP7oeFIR1S9EgKkveWKZELPt+rETH8yd2eTr7qHG
MN6t1qFUZbYgjIwgd1O2vfCAOXGB4emUSGQttvuAv6a10lg7pWKGlHn/Q/FlSm5O
TXx/V/zaTPtWr21AsSrqEeN+6thmvCzJ8gKgK9pZ0KFtK2ne9UBazMEAv4yWH+pZ
mRnwtgHZeYEoCCc9hYY964kp+cSHh8PQXuq45B7M7eRC4b5PubNxjXogGEgYhZXZ
7Ez8yuIKPMvpyfvgGjFCtZJx2339pehLYhnJfEtl34R35dPnRPVdqZI2TtBPvLXe
EkNpC3VlhS+p5sjQOuHjTE+5KmRKd2JREc51GQADsdQ0yF5cnMIjzhLkt6J5mDKA
vNme22dtg/QrYTZUG2kdHkJaUZ4CzXLHM3YPS0K0kJUjYz+jaTzUpiM7JpRlFWTI
aE2IsVJDHYY+MAOPhWcWWeNeNzlZ5g0JQC7nM6Waalkadk0meZBWeFOuvx6KHShh
KFS4b/MW/Vn6SFD1+hsIc62Ownb5q/V+BdnsCRs5Pb8FL9zzTPshrE9ljO1DZ9ME
vGRaA6Gan9QfPCQUkoz1dD5KFuoixpv+etXzlgEkGldLic58iBq80UeBwkxz+vBE
fGp3Z6c1XoAXYi9XGNKKMR7zZe0KMZy/BKmpw7+/SRQZNb54XUUAuzxqka361mzg
hUo5uBIgWfY91XjlbZP+PKb9gYmuB0g6iOok/e5DZbV27xOykzn4w6ZNVpPULltN
zCYfsoGp87lO2LWvKiTmauaKfI01s+IdjFbnf3abLxFQNpO77FseDDQ0z8MdE9Lk
taQlKqC9QzVFvBkGnizrvoDpNPmgGTp7hGZG4Aof9Uzct9j02dVPQw6Sje+InSvm
hxS2w4pbKwO6tvBbAmERYob38EjjviKYxR9EzF9ywapJk5QDanvcWXdFPjWN0etz
eOqgYctERlW9JCMxyiQlG4nL8kKptIbzxhIGtB6ej5hEm8wCIOkguZQNxxOnpMtc
Xz7AJhmPiPBy/1D9IGSYHcnmCJNRow9wDd95lNgZph8dYita8muDQuTY8XcLYejb
LIDl+aJ746ndyrKppeaSjlaiD1tTULSxi8qh2yCSVfmACIvARW5EBfxjHQSm3ATZ
dyJDzeNca9CRzoKU8z6sHcYbpChCIaxVzIHtDXizySBFNkCn/2mTXbQx3p2eEEpQ
gQhkYJbd3wYRTSvy8lhepnYQb6fDFaUPDWCT/a7N8OV6L4Q+ylnPPpYuhn50xHLr
BHHavwmny7cU15h7Us2hZo38EyDsC7hGnfSykw0//haEC1boWUm0Hl5696bhizoS
zedrBCfHOfsa81NDxuPMGD75Qvhd/COtGOicLNeFzHcFDhjH5jPQZz6Zka8tVpun
p/Jp4lPTGxx081gNDBUKhSyIhn/QpH8mulquStb2REmgrLS/KIp/5La9pItQdEd/
Ih55TWfQCPDLTUEs1v3qkXisgtHCS12pyThgFLZVa3axsN7IGxEBcS/ZdPjnG60z
K9KTQOEBwAMrsyyuxEsmjA4mUJBuYNt3pjTot5qkEtUZEWKft/Nvp/KHcmdgg6Hs
P8DBZMZUyRekeUENrT3Z42wbVflcvlxttpXMWjOHaREt4Hc+TA1mMflelq9uHgbF
IwEFVBvVJ1npuyEkWAMmFXqdJxhjid5A8NJbc+JvrFmzSInF3QhxDtrr88CSwU58
BL0FCXnvCMnSG++a396hhfZkLYwT4H9RO5vURDjg5WuGiOi7UzOvr4FwMrEyOwLx
BSjBfI6EnhMC8bW7yQOPFd4Cd/E+EKpAVekGJcBcGNdzDCghOkHvvSxoAO+L51qG
Of/puvqjzXFdxplCkQJ/UR7MjN/qsiHWGr2FZ2ke2Fpz0T1bEBurvd3yeDa47rGi
E3bOsEaedlVgOjS024eKl+7+PhgY4zD4/JTn8X5tomE2u1WHIOSFgp9A13C2qeVb
VoWfCe/N3LY6xbwI4NUdEN1a7zlhMJfVnEgsMJArnOqsNoxe3dfyT7oERXETDu/Z
e0iVn7BlkSqwNos7yWbQ+Dz2XwlGqn1PEF/Op25hEYfYd1eZj3mweUDobdaBvN50
X+0kNLq8j7+bE3a794kaP1lnRCkuq0nsdJgATHu2KEmeX+0SSkF5yhkkggZseFZl
7kfnWo+ersTz0ZeCu3J2hYDG0WtmMXIuOk4KKypQ62xne8zmxbgMQ3v6F8nC6yhV
vXh4ZLgmJ5YbYvuWPlZISey21PRZhYc4f1ucE0JWS1usknCqGKuEcGL3OdeL4xZ/
A/iDh1hDiUhAuHBtji7PgeIBV5g/jEzcVFT8n/6LibqoYyCKdSgMFG/xSjQtBgxg
o3mGx1fHFeysrAQZpqqdjS2BffZZmWwlj0O06SqbQFoGKCbRDjQpG2DtFxzUbQeO
PEDVDpQq3FInWcS6z5nFC8grEntON00dGaRSw87GxD+kFBEgRPwU6V65d80DxumU
pHAtUyHLLDfCoebtSsqjhG1GZhuON6OLhjqhvKbh4rmFPFcKM3PPMcYvkg8QQsWg
7anzM64HxLaZX+7cjnTVgfzq+Yx96BaDV8qdOkI/R3xoWEkL7zx6kOYjQlnwjdSB
OH7tVnZ1I9LIIVHxb3bH/RJ+pdtm9aRQK/jsmLTTad1he+HH2zMDAaGjZgqU/Rd9
`protect END_PROTECTED
