`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXJ6jolcUkUjoVQar6eXkv6kkSxxBqweKPT53sOvbIzJTgWEhZ+3z484jqhjuiMi
8E1u0cQ1VB0qKK3/jumC7fi2ZB6nu+LBq8tPy4XV8PZzbrc03nIOjsDbmpjfnXNN
nDgb8noTe48UhkAW83Shq8kdEKmtsCnyt+TlgmCBu7VBFguf+ED/E4NXrdFa99Lc
8ZevQmya+usW3NauwtqpvErLXnKcgDwW/i79YTmNa0IYIkewaVavFvuv/eCR/gt1
ewhsusUH09heKwfAgfnIuG9HHI4cBgGxbA65MiuXrAf77iL8jzIBqTKl0H/kkF6c
qcWm1xDZ16MbcaCK1TIAozT68gfT0pbNuWz6CE3ElobQAvahXJhyY8zApjk5XGh8
d6xGv0d/fh8FpaOtEQ2C+EiYqoAZro7ZTSdiTVFDkV6rJ3vSbx+0YxO2npofJKVd
XSRKIY9ZaZE4O5duGz3pLi+8lOo8G825+id+lYlHuNbCEqH/QbmggksjgkHLQKMw
vgXrASJokzYccYG3VbahONXaixG8CrHRmo0t5Q9MnQEXX7+fBJzMSXh35gTO7o1S
uSGp+9NMHS8grEayuuv/GYgF5IeWmhIWMsNNQnGGkTYwT6m93cCKK1d9OiDnOf1n
c6SWdle0i74cc5eLDHZgRz+TMKM9wy19cyzTXaT7o1Mbtle8OvcDuNJTA0wAenpI
D+br269yoexf3Cij8WsbP88V1+5hK/qMlzWqXmV1t6+hOVsXGxau2Gz6LDbUxJsA
I3yd/5HFxIOBT0/4L94O+qT4LtZJ5ol4nFbAB9krFPwBm83qGzcMKLY1RHBHhEj3
mDcJ0QZTTHSNEFxhBp+CVTL2Oe6K/8Jwt2xRwgS9DXcZM4sbqRTTPJElcdjzNKfc
sfBRiFrXNp/mXokk2dsMSMvyMFVJkWlgc9+raJwIi7A2tvSy+4U7eocJ46nXnKeD
LZ8N6sMmJ+knY2J70Qg8zLbATBASOxoporzyLYQnmXgnxMH1lixgVZRO3/UJeC4+
bm/fDQWfdnZLjVEyLSQd4qt6WYNgs4whoKaQ3siuf66C5dACmSeoLSTt7F4x/0ZQ
zj2IpJT5Nmb2p6OXzvrPO85HsBEc5q/yogqlv6mVXZQlQjKOfnKcItfpvhU4/XQe
Zvs1a6KduYDNAfpPhc6DYU/aDJU6xLW0wi0DCU4cVPD2l5KAEm4EIjzBSyFGjciG
pltDBuoBb1jeTDsenJ3ndxqq+WI86wO7kp+ttTYthAm3pEcwHvR49aOenAE0nGF9
HhUjxTpgTqPM1KuQogQDg4a7rhfKOTYJaBZYsT8PITXKbBXiVnwCgmavD6D7zL4c
EUOOiJe40fXL/K+nJyOQWdB0lBLNa6TQzCE07hIe2M2covMpia0+SwTH/oespG/j
yi+QccNMZZexW5VepGDdap/UcMpuqsC969wvnEqVYXuxx2yVnAbAuJjTnC2yQjxt
`protect END_PROTECTED
