`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YhdIK5bX5Td1neddx6wJfsCYAlUSq5PNcvANeBo6JT9nmNVU8wAS0M4kNjQ2QqRp
N1PyP0DOCFJsocWp6hjPMLjxp1t5MdgIJw3t0CqlB9yEmsTGO+5gzYn/JKNUN4O4
5A5uspeRZeAsrqxdAPXhoBpZK+8u1Eq/ddcHoPwsh0cAiWG/iT1COqVs0pWi19e5
20OIMj9uXF+KQEXLJRPT30PS353/zbeMYzzfp0a+CY+U80vNWYFlG+eJ2URijhm+
H/sgFc6frxPIRsLCRMWb06QLZXE+rot8DVKFiASpmB1mhQHyUH14nk5PqZ3UN2Yd
Xs7rD2NVj4pKA9pw2pQO7xDP1NRsE+Ebryl+o6kWPozam886NdDAMPJix6Nb9gdg
aiCxELj+MlTLxkmaovpuFJSkHqoPfeYIhpH6EtUKaxrH6ZIsBRUQ+pOYkFYpj8AW
+vjNeFanhG1AuPPVXJ3th9jqLoa4HkLe38ffcwGH64JUOcsWKlOLDbnzu2CLzD16
zLEeh3A4YPhzhnWYXkqU7WgukJEjUsq4UOFCc/hJFLYP5ujKAYa0miGt0TtYqBFV
ZFHV7owJC46dBVdzMpDWNJsyiWN7/zr1jDj4aA0kUcDDB5PASXbpQUokIpqWUXa+
84HhbaDZ3v8a9Y9yvgRwFIAb58dqqmgjVi6+d0GHdM5Vuyz0h3gQdPO9Nwq+wgAu
RwZ8hfIccooRDFIEIP1AbQRuMxtq0KNBnG2ZyJYMxlfHtjHO0vLI9d8ee92vWTcP
kZCprprJIbqN5ZE+A10hkA==
`protect END_PROTECTED
