`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mXAuREN5xq/vnuJNMobgHPCuYLRfDUATyvBoftawaRyPGEjknPbKkcqYW5it8xtt
GAIii4m3oGyieF1c4too1/irTP6igcfqI/452IrL6UW/eM+KBFQHTLUDqhgc6qlq
7CeZ1aCmUTEbYPwbCPfOk+UHiPlPk0JjMlnB+BvXFslGaPxzBDlWpTQE5NCFY05R
oA1S6KFv6PQ/oh0ywLhq42J41jGPJrrGm38letPv+1OwITXmx6HIgIWQ4iy4Cddh
+HTF+qXHCL85SGVLY3+bsqMXjmPs5JKYodLjB5AMJbbhGAHZjLh1QuixNu298mS0
d5skHDiLNsBgGXOl8ii1c3eO8ibqwIyCtx7ShyxfCVEnaS7oWmGitnMeAEDl3JGr
wfzRNenFQhJpNNzUADt01PgFqXtkj2PpKXHaaQeEpq9/+P9QgI6S7WUbwMszsK6b
lknPaEnyjqH90LnO2VvMbccZcfo7D6B1nuvGZbn1vX7EFt5Jwmsrm43009DOESPk
sh7nwta/Jnalx30tpk3JBPS1geMnNacbZC5IMuVTX45ZguMVauuXpvLm8/Ta3+KN
sRosghzP8YsbLPK806rdM1z7XbDyWX0pjEo3hPkeSTFbydWc//w1FiICXpCM/EJe
+8inC+8jWQEQunfAAFwHqnWreQEiITtbDYlB+ZXzFEjy4BWVq5AErhXny0HFUhBv
+CsEyVjb6VrEsmoHR035w5UmkfBXoIPNxPx3COc3TkoVgTkTp3vOEFWj0PQc7fAJ
VNxTF0doc5zjf1eCUhw2dMXFbxtLaKY8KrXb5JhZrHXQMIVzQAbkKgA6kUSYnxlQ
UcsUd4OSCH9KFfPvhVDi1W7OuFIiOYL7ieYIyeLD/z8H6zcLts3p7PYkhw1tA++2
4zZ00s8oSwcoA1J72YT9QH685lueFpw7X20dw9giLbqDeWot1EZ8vgG4GuFFOJHO
zIfQoKQrwJ42mNOFXifLManPN3bNmQDz1uUKpLOa5QglgeTKnY9OKGl8RV86SLcT
BINm5EXymBOaBLNSlgdaiecRYy10JZEcu8Bt/7DC7mksErJeuhBCCXT6RPxULeEd
Rg1aVrLKTGdSpRQKHXHeWxQuh7GH1ghpyAu/uqZ1c/nAw4CgeOpzwNmvpFpaPuSp
Z/XEAplMLzrqUnYrnXKNDBNjGHl+o9DWLPC6qOHNQGCGcSn1zvbvsn5K1dhe9648
NWlcAGglreh5JFZJoxxvq8ZwgHBF/I3sBUAX2cYq5a+wT8iFfzVRc7XjmxPIEcQe
ZOL7IbS/Z/mBXToPjt8KvgwIL+tvamH10XzYaHy0Qz6rLIWETwoxhKGxW2VWxL44
H+A7KGOkvGUZHakUZVQYwF6GK3J0mtIb//M0uwndGZIcTuF/wcGfQRpr7bIgCsRw
OVKlF10iT8m3fGdrMCVGEulnL4nzyPLKXKKMVcO4Duh2lTP4HkqNegyrMYCo7L7c
DHP1eyHWRhic18/+wq5Scv3+pHAs27H3xDedjM0EN8XixTsb9Q1qy93d8IpnogAc
85Fy2XyRIky7wk2rsAqLQ482LqIGym9jmcosZ6W3uY1pnX/2QPT/k8S98NnxK3jK
18dSTiUPXiSpX6h0W9Oqepvta8IRR5019BL5pz0ylMcZdZ9N9+u765WTX2vn+LjD
SR5WDSixBsYjbqVnWnBCshYQf0zK8WKEHeIQYbDqBPxn3zSNahI/2ExQQOu/IVAM
YiSVjCS8Oj+1KlBUBwG34KnwU/64+HXp7rvZDm9aF3hURnGdiEG+Aiu7XR+tdo9f
k65A1lJT0lRy3Rg6wUIpygPRayicP3M+fjyLZ6JnbrAgRWAwvY+phU1zWns9XwD/
oZui9BiFGN0U3NZf4FAtBEAf/Lhf7Eoe8mr2ynNRytA+C1Rt+B0mHH6iXPEAkWuM
wB5NHRwJTJ1S6lExCqVkyWwXcnlwUIK3tLUsEQt8qEHo3diEagMhsaSjB8WQ0px/
mk4OFI5nRLHLewKei9EVUncf1eCY2oeOvEaEgublifZUpRbTFTqFqDTD/OJrPSTl
oI26hAyHjaQz24dG2urqqT6YIizgf6h8mpsXxsLzf96qR6f0pKGNCOdHCt6CfdOX
0rfGjfqpnvm8M6Sd5hRvhjhqXZi80ooNfp0AsZSvQHkAoJfteJsfk6gOdTrUP4uT
/mS2inrilT3ptLgF773Mcs1FQpaw35Bbx0OmwHp53EVfzRYjN8HzxXKu87YD5XpR
nI4cudcaU9GwRMQC+tHvBzMbNtMi1zDV++XkK9JqyzpZ9gYisj2lpAqqD+Bl2oF5
+BaTC5qlANMgRwkmF51cWoNtoLaphNpW74A2Ec3g0yFlGQDKJnjkCou7ZUrDj8Np
Qg/Ew9rB4xyDkTY6wV0pGi9VmKNuOsZAa6c0nd8Rsrs2DwfEE+62GgAvpltkd47z
aVOF2ENPeTec513EfMEPVu3mG+GIBOcDahBCHZN7VpEzcz+XD2ueu8zbM4kt9d3c
zYOYmp4ex8iSqTWQk8ksWipls2n9migYluzjfQYljSv0Cg4/4wsJTFeRXaTAj2uV
9rKbn91oj6AfSFIOXBza/yclbqcGcDW8awqZlrECeEn7X7XnWv/HvC+ZF69UWNod
3Fl3KoeSW8IpjlyX3xvcYjlaYC5mxsGMidtZC/8HVcPoBw2US7ePgF32zDmBnlrQ
EcFqaEJO+1mwrczRE7SKfUSZ4te3vMGTa7X9FuUC+RLskESNt9y3tZGZANDQDADn
SMEOFhqIozFwMZFQhM1H9Q3JvU4XqXwadJbeqLDZ6JjEtlRO6J8prvIUyfxz46Ey
PqUr/hctv3tJMrn1QbSqHvZLRUjm9SNtiTXJh0JeSW8GvF8WVCry/lbXPWmezdGD
Fxs0ROAy/ADMsGPToKOG8CZ7IkfF47rd3NNPTO5DzS70w2KSPph80vCZoyMSDxb+
SvwyWaE8E4zon36x0eGGqi4/9s4LzDvV8sXVLFWmTEmOh4dwe3JTUAk7TTD5965E
gwdnUTJc+YRWZLFmvTo3ON7ew9OSFu3I2VGeKEDYQ7TcS4Ol8kku/HO4bHipHvJz
IjYi98nMjTRNe2LqUmFwHs1pCZobICjzIqatnlPhazKRh+sOkjsZsvVdnEzl57hK
E+14E5hGUW3aOulnPBJN7H0Lp4jHEtZYwhh8SYSgHNMAT8GzdP6b9K1FXtLcp4lZ
efcFvIYzSz+6o+sPKmbZbw4p+xK5qG+oYkfno2MrID0YBUBq3Lu5G/T5GJW8yb/1
oJvtAaVPa8m27MhlawvzYz/eaf4mGcwJ0ZuT1yZA4vMslqXyktcFWtXw38bLzLo0
6aCx8lqwpGcrSjugcLSZJYGE47+yT9gm3c1bXbRDFBSi3FcM40CqkQHl4fOnIj9X
HmjE2gjnCKlYCjj7qW5+eQxk3wDAxtDUFQPlyHyITM3/VDJnTxBrhbskGLB+zLrM
t6khCZQcUw8sF1L2Wbev0/vVpI+jPMdFMUw+wK4+RzRUhTYwYdwmzNtztnkdLGwj
`protect END_PROTECTED
