`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGS0Bnb7VvJBKTqKmOrlMB33VCkzVKGSopTcYhHJSH8Oc2PXjiCpjS+I7l8hwe+u
9Vn1iIiV0AQvp2sNYaLahVjUJTMYyhDcUX5J7JZtGC+33HjXacG86QwQBz9uBMTV
n5o/xBSDcH4k/TQIQwqsiBSbBXO7nugQoiAIKLw5Y03MA4FaZiOebdeIGCSRfQfA
VoLtF8j/EIN1RmGEGb/LFpYv6KD2P5I+V+sXFo2c0jVuFpHjf8Xza1C1+0+jXI8P
7u+xZdGOrYdvnOyrPZr+TtTAIJXbiHvFVu+KHKbTOT0KUV7hHz/jr4WvvqGMmgvW
HQqQ96DrXSDzZnB6yFyMlXhTps955pkywakQPZG3hAyyrrQE4/1nfrGnebRqo4qg
Y7U4fcPTFNCibJtDhzn1jDWnd1NmRg8Ik0wqgQOJyQ2weAeeznRKp/aK/VbCTwDK
idK3SWCeYcpEF7rpk2hZ2DOdQBaBCWz0ZoqA1Pd0naJTyFeOm1v+dvc+VxX95/xE
5azeockoMTc6R+MgZSfhxwdebywa33WcR1HYl70YH9HNdF/h+2O8gEI9Y62pS9uw
zjw874ZSFbToKVtYAGsIGOuiy+RCYBZ9B4Iz/q4XEN0JFaDvpRhVdRktceOZGrEP
qoAIRb+DkmzynSxwxiq7qsq1Ogh7mtQnY/0+JxuS/g0iBfxgTuB1OEMSIx0enUaB
1PP39jHdt4IhH/te9ZIpS1xxmxVdr8m12xxnYnaAlEYmdC9oBluv9t7zqaOT1/pO
KAstxcRMaYywpGfdW/Rm0egWdllbxtCaOxTvuDIEEvrmvhy6r6afFJF3R7AA7V26
2qSvyzb6SRwuPxxYP+k2EWNafdNGIULjjgcBTIt4Zl7yF21iem8EHGhQf+ptTug5
LYq4rLpUUrmPRCcc1k3Wf7WsIvlrbCNJE54yU0NurMTUBCLeOBkl0rjzJHoBEUT4
7NQrx15XaZ//FsaYvAyifCJo2piy6ZmXGZpGU62heNnG3/iHfOqaBqtTZQp1STnu
inYZEl/rDaENPpdhpQo8Lq1e0pjC5cN4CYx98NUmfdMJ1d1xrnT5tf9NfutCr1Z9
ztapw3+xEUNrjyD2KZvFSOvSD/6JV2C+B3JYvDhKF3PED0iUX3IasH4blwXj7/et
ShBc9yWk/MUzuMpC50N6xAL8YikMLtidr0e97FBViWbjQRofJygawu6IrpsAyo5N
ybBc2W9SRI06kjK1vkfDkrUyycbc0m+6tYoONm+Uqrr1sWo7WSmynf7UJWNKpFf+
CyTTnWrKyrNsh1f9J0EsbQ1QwFiD5ctglQMrZP1Lqh1pNlmk8W2Qy+ktGCkrodk3
9Tnd/UL19ujiSrfZrcU+YlbCfXtk1dcmlCyN5O31N4COAZvSS+WhlqeEUhsxya5X
wvrERKt29OdekwaD7NZXf+11jd/+YUuiSZ+03C9NXflU1Y/s6+Bu6LyiKPWu2GNl
uHZ+jQsiTrR0dBV1iM0QRk/Jbl4XEzUIDzH6KJRzvF6Ax8heGab4p5YOPfhMi+yT
7USV7F81yP8IefbDUYo/Jg2gv1B8qHiLlvKma/qsHS6aCKO8Q8OzcmFS+/xQImPx
Hp+8Bp9FLe8mOFtIdyP/NrJKdMQRQ7yKOU9vOBAVz8aBkmwxTDJvLE7VG3Z7/TKY
VU73K184rVM+JYb4r+UFXjL0RygD4QxLUtT84n8OddZElQJtxc6Th9ObJX5aK7jq
v3s4cfyOd8+Cvp0+KvfG5C650UDTlvzP93/K+wNjWqOU5duhieg4vBoz6pfVc1aG
hS0ks/I8LNERMqhKmdYhauMz4OLQ6zpdz957Na6T+wMZ0oMk2TTRfCKDARIdYRF5
ec0c8x8vg+8xBgJ+uiorVhLKpvmKLyjwdXA+CYaqoUmQq1PCmzi/KpBuFt/f69V9
U3h1vMpSkoEI4lbM5KgKVMQUpNr+ADoVVELdZP3lCZh8tUftd26aIZzl6QExqOL6
3yXUqQ2kwzxCY6zNS9wzz00Kc3ZjliBCAVhxketXArbuyiYS/+AA8XxDXFWa2AKe
MeMW0+cYcbGJ4QIRxWgqMTg5wTfeVttv5voE/VsA6v0JNp7jzV+LqMmfY/gEVZwj
vyNJ7k6TPk5+VFxMrN6D79MRFAQqZTRPsZ3ivtDd4fM+I3TopLjeu9uOw0xhHBU/
xy0DowzoGPmzxJTYrvI56bZWpu9BQQ49pE1KcDCrfrD9QUpIvQYNPW3XtcD+PKUm
zBPXl1jJHWLP13GNbijbibrQemRRo366lXBMDDWebELysAk+YnEVH2xqBrFbMSiH
8WdplAbYV7IlfLrEfNFG/OYD7F8S6rs4j29v1dfQHrQx6QmI74pzyQSM/YKQVFMK
uVw1of6aqNx+Jffr0o+0Exf9i0NNYPfe4PIBnviEJ3SF9igqCVwaqIgMfAV7oN05
qLnUeH+2mP3KmdR4qleFR2EOzCnIS/9uUJi/cEq7VqHQqgm3PWpi2gD2CU8fk6Fb
swtjBnNIpEwBKhGNx/FVHsUqOEJPektt+K8vhRQavKXPLuTy/KyjXNGSzt4+Swx7
xmhRo+H4wZz9VuUC9jVsaP46kvQn7pcie0KOAfDGLI39e2tihGmqpLFf5Ee0myBX
8wksL/VaK/hw65G2z5YkO03yT4efpLWMZD8um12H50Hyd1fEZy9Gt2Yn0NtSo+EQ
hyRsNu9y0gZJKt10NK6gRNmUYEXD3FYllwKz2BD1sWeOhZcgops1FLl1MFaDK/85
Kogob4oO1sNCbsl8PXNZxmVvAJ4dbGVS/rz0M23aCIm2gkglKMkCFnEBdAR+qHDX
IH5hQ1UyNVvtoUfPYC9yzTO35iv1yay5jwPlZ6KH7+16r1akCptb1HIRiHULZdnu
YUXBraUyVZkiXmjph2OtseF2jJyFL25kDcmUQ01ZHNRBEl4tYDuz04Iy5TnOLjr9
4tudFl1wc08rZEm2u8thZG6FNa0AE8pDn90XAxbzE68BzxdtsXb3W84/nhd3by2S
/S9qwW84TosfTRWh5g3jDLkIlkR2a06coNhb7TZIMTNCd059Ij91/qZAni3V+OmL
WV/4zNopEzx1PoDdv7/lK4qE+yxc6taLzGgm+WlIgzCYW/nKi5KbDtQH691N918Y
m4tZ86FLjfr9wUqkXB+mEQpCoNhxuxgYxTp7iM30VBAeQ3kf7XfWc3XPWhFv7ASU
M9UcOXB4J/GRHIKMHWhZWvq9X1UlEDmd/x810pQFyYERj68qgsjWwf96IUXA804i
rkknbWNyT+JiqO14ubsC2UnEmbY1h62ay0+/QeAESIUW4EVagsw/ll1IsH6Y4aMV
NfA+o/MsVUvguMi2HfbPFc7VM77l+oaKjoXhjgBWvjBJ6lGq63qDBkk3dpoQ7lG7
WSk8g60ihAzk4GuxbJ5Hma6sJpRQB+Fsy26dJ/NuBxhzdjQcryEwUXEDeMeTjweM
TvZUzopKHGive8OeAt1Ft98QRJ2cj5LxJUbdlZZk1xxmiedyG2fND+8b7GeEvyWC
CUoWQ28ShubxVZT/9qXkerWhF0WBlm6DC298s6XEOYmRXe37ccp/2rp48KchcHwP
dlIDFu5WBNP020hcRAbQri6VYBBd3kQP/yXwxWNZe/Y=
`protect END_PROTECTED
