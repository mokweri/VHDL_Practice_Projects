`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fNiBkr6+b4q0CAr6T0UX/JRX2yJ1t3ma+P5TJhSUwwvu0eJkyKDOS4p9GF+qY+w
bCO7LQ8rz46BEzTZEC/6o4/R8Pwu4bRlROOco14AuAEo78yIF3mYNpnJ7G97iPvt
nT1+yl9U4Ar2BJ0aQNYxjFY02mJQdKAUvhxidxJ5npsPgpuseEyyTR7XD3K5z+tx
86g0/nAWGTv/YS24tTdr8Feg7RX48Cuhpq2Qs99rx1kBn9vUW8DZnb7PemL2O8E2
LIkfuRdTUs0MFFnvgFiMvoj2UDZIlLisGUyXqP2Rr1qlxsn7z+/8CPkVW37e9FOa
msH8B51iEcqe9kdmn8fcG3WvuIfnYCqA8UozZfVZf2z32a0jN/LR1bNlEFBeptjM
r0zZK/8O4GjwFOaey6QMJb8PRxl6pp8A7hzy33Kcqyx2zUG6u/kvDF+Op1K9VLpt
l/WOVxm8ql7MfpfRx2ZUsAE4+CsWmLe7hdVf6pqdjniITp0Lc1iNEkMsNOFDLTOm
OviFfsv9A2Pl9/juQHzGaTZE37X1tNCQPrNe+8LKgPr41rC7w3ADm1CznCXFlz2+
4KAcFo0kL/07TJVXbbF1vpXGo5rCOEVxf6UAUmUFOduwJt2TdxASO2Wm/h1eg8zt
bpok1ZTOHEav5TzJRjdQRJ4w96yJqbe2fZYzXZtI/ieHM35HfdseK56n7lGSYAue
ylgRjSGHwG6s5QJC7LClryqZ0DzngGv+bxxlKJVJoaURh9sqh9L3pgv7GVG0R4kn
CIX18y1CJPR4QBijPgD5Yxi0b3C/+qrqkSfr1CcX5D1vleEUK3Igu2OOuzMtsKJu
KxvAZKEifsZBFwAUd6dLMpWOwNyLvSf6pVxiiENbZzgFwxuV5RoUhXycVWOQ09aY
u16RHbw/EZehgliDYRTx5enw/kiyu3mynqcrThL17rux2PsFPezeuw2z3WF68dXA
4W/gZl9iILFj/PaXTxMzTz9vJIwwlt0ifErGxy8JDfL46xTzkBBxPJuM5l2cnP5I
fD2E6fdLJuTpype/y6VmYIKU6wXUR71UJ++d8QwSllw8S8JOc7QEt+pH5sO3Dgcx
bsuUsYoYLO7bujMW2N1U1YHOWeOeT1XAZ97g9CDrZMOokldUYcpPyvtu+ala4SMC
JDCw8ar1TCevSGwUOrLXMVlpVigOOIg6/zQoH6mcLXmqqpb+XnZ0T19T06l4igGa
Mmq2+BESy3SaHQKzfb8Sk+U4FY7qqnPpvHKIkii3P/yYthfiBqiVgJFkJvYcMalt
VP1+fDbVik0DG9Cgwgc3o/jMSMshbR7hWeWSKve4o70gQKlpngrEmzhHbNQhZ5SE
QSqHbWVXoUmgIsnAh35gR72zROUARN/XYeig9hWxcQB9bizsjeZY8h6KjYSnpyWB
7qkJG0OU7YuA6QpC3KDTUTf+GS5HG7KtcTTOevIfkDp23BsxqrGoSqCQnamP9xS/
zpaucb7Ocf5i9L3/zo+z7c/7BPX6EWaiLd3E7MARMoq79I+ed/O4F9ktihvCSNPL
hIDq0V4DacSkbFEkTwiIF/o2RKD8ad9YBZJqOaZJmzE2dEAduenEgLmmgJG95WZi
TGMRDDDqmtv3FhknkSjREaq4KZvKfOgbj5kWzJhIKBmE/oA/xaEjhRaZLd3l2FJC
gOwTCtryVLgLz1OKwCK6EwWLGjDBS/uzv1wKVQSrrZkNL36Oyi3Z9bVgdeO1SANM
xaeIm+sBQLZx5q/WYD+KK15iQ8Mslow/ze2qomuJeIge0t9GHE59cRdY1PvRmNaU
vArkDeTO069XlYLfAz/Nbo6Ara21HLlDh9LaECCXhLWAJPDTBqOD2aYSC01SQAMk
HvgI5FlcIGrvT584nAkodWmaHHY4mfxibvda8PMJQgL6eWCxrc6m8X8zNlgKMj3k
dkntR3SpLZy2tptYj57lNZaPb14P4iNRmGmgmFp9UUs6yqAb3A3P7mbjWHN9UOPh
BNq/ExJwICFv3LekYSFdrTCjiTXqwnvCoZypTJvMMNh9Z+yG1VVKxZOgLHwN1cki
6aNOBCywTiaohCQiFpkd9sk21AbItZoMRJZOu+N9A3Nx5Qtw7Ze+77zcKjkXQalI
E2PLUXpeCUobvgEogjPvoiHoQ9xiUzGzodyPXt+gamXWdOI9cvH/qtLSirs0cROz
u0omQkryK/He719UFSg+Tj6ZX9YIAsfvG2POMu0Ewm3WvBDWW9ic1bBt6KbcSdB/
pZB65ftt13OK2LEb0sHEpGbl6UJx3nw8W3uoxAl8XRq7JoUXCiEw8woIxlhzHPJV
e2oXRFHrNhEbcmai5I4cHZlCZ/VLNK/9V3hQsL5Whegu2H72WiRS15m7QKzUMoc/
919AcFOqzgxfQ4LRt7t12EdRp3pKg1knx89JnNdTLRT8lLts7aSKzNc8SvnwaGOU
qGSshPOFiCIqUxRLcSG2FizLgT8G3kRKBQ/f9JOz1qvGH/IKp82UJOpG7t5eHpQR
mR3Yp8NBkev8kA8d+280MGuOiTbaIL+z+3goBBfJnzf80uQSRUQBXUm0P1Smam/L
2TTWImqhElDoVOEsxqFTipH8iCblR5woKFMnyIaEdeguMGZlCM+9CfzQSAfECEKh
N4fPHIZPdEqPFuGB0UgHKVIRaYh0iuckoenSDhfO92UDshj/vB8iFJHaoYmGfUur
WhHek/suRe5f8DN4AaxtH0JXi2D34WA7EFeotSmzguILq5hrtd1HWp7QoPut4Ecd
J4GBduAb1bdak/Ltz4pkxyWHVPEI92dA98jABbfw34r+NlUQ6kjPJbijRSZM1ZhE
hH7NRP4qfp9/XAqFevv0avKAV1oJjJh2Pex2wPx2JFt2hSAO4aZ2Ps6r7LMOP+w6
U13WSI8zQlNCROdn4N84OQchfoiJv5JDzjS166695E5iUau1MpE83GU8cQ8oSoEW
hUT/9hFdQD1drAFcOnCtKRMr0GyBL/LiEzTVrRffXAXCh8K/n13Ui1XiCe+4/TcN
hgnNua7MOZ59ej6Kyzpf1+FotCnEJ8XEkkJzZvyuHLWh96SRx3X1PsiA6bc8eeAA
rn95Rf3D0yTHB15jmG4P9aSsCeAD+b5niKdGxGveKTgDoZyfuYiZMcYW+jjXk1HJ
PozjyehCTECqUDrhs+C7CzMFL1f/ncDZxZlfaQaX6klFFR3xi7F1zBGdYin8Fuyl
FD/IxJ4gexryrm/Eg01D4u2xqc49oWAeTqlAnPOMAe5UFz3osA5ihaTsNwohzZXP
RSKvyG3d6QbzmH6By7Flml+tF3jhgIMkl46ycKDObN/oRzy0gjnhZr6JSknmFccJ
BQki1ir92yJ4KeELU5ybs3T5q3V0mzgw8Ma+oLLPqwGhanJ3z//L7ljy91goV5ld
QQhx0zrBeskhBljKOF2fxsPpLqgOFcRJbMzE84MSTN026HeY0S+vRX4d2OIFyjeQ
xg4Fe4cATuerkSn5KHqstnp2JM6gHCWk1YV17qZgikFKNaiUSIuDZO1hOBv76nr0
DdEdCmp4hrkSgOoXP+UVr6/GVQk+XH0QbA/jLKFJEBo8fWfAxrNM/eQ5IJZLKrvZ
P1WmZ1oRRFnJ6C0AeUBUmskNpl5vV2FBgYezRzdndLI=
`protect END_PROTECTED
