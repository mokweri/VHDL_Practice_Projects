`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R3SAmnPJlkzhXA3w2ReEEWz2jc0RlK+YFMuQap1WLAN4yH504bQGp/HzUw+ulNfa
RwF+2+75WaKdwZQKz2Y1i57vplt53bCMHSkeLhKq7esVLN5uh0UIJZtHVmz+c8An
8qlzsDfpy4IMKbP7h39+VEDmOJnzmIDpOmjNESWD6Iyp+a5dDJ917sDAljYZ79MG
03tUu6euJvdUJaxIFUEsOGtMtHYPuRl9Db0ln7Y9KYb4aHv0UD00zfSC0goscpsv
OI6SXUEY15mxtFjOKtw7mmcn988Pg3oa/OcoRN7+mYzNU40Gw3HBUIr3zOFhYbmq
rclfUYQIkUbX2acRF3HRrXHd6JdGSe5qeKtF85OOkumbZ16YNctftDUJ4xbRWxT/
gstWHvO9t9FunYRs7RJpYKux8p/zROOgCazWevVm+tDVeX2IvbnWkUYs4qsZbS3K
e27lcUh91fxGqiaPZdQXMJR2AxGrmpf2dIOHzNKW4/r2E1fLdhYc4swi8S+Jhpcv
kcdU6Fg2j9wSt3RYDbQT18jL1dmUma+PcCqmmo11YgDoaM6p3LYR5ATN2He1y1sd
3Jbge4Kw4t0eJvO/aSOoURYqoqrWwNLmsmeftz0pOC0p2C9QPM+zyAK5nAtbneis
XmdEXSQ/6/hC3/OWz2LY6XADEQeriPekzfy2gUObohnHXECE2Xrsgr8eSUgz6q5e
RH6OGS+g/RwaPVD6bPbIRQCvZ9jZRT7i/GxBZWDhYuw+ZNvMSGyWpqrAHamW3n2G
9IHIUkn94VljtAsC53/aRJ3tcfTiH8bsQ8P1HTQkDqZr5M7NkmylU8G+VoWqFgZ0
`protect END_PROTECTED
