`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dq344nbTuqX50C9cMr/fQqk8yZpIDOOXBcFD57gR6xYA48h7ipj/yxUnNLXonOgW
qB+IzsS865ppLavNytR1fOuNEuiX98DtQuyGxWnH/7OmBxtGtun8O0/sF5otbgZM
RznXLc6noqv40VeLlb/LwL1HJYdqkXgTgdZbb/kBTdx46GFybnC+TsdeoW3NxxUj
t4NrjAa+eIbIhRymrDx+UUpumP1m0apZUDJn1A8QfeADGumsCl4g86YBk9DdT+H7
I7ein4cTEE7u8Tq4wMTSiGLk8rYGE+AlAzcYefRZUkXXPqcVKNrs+tn696wKHEqI
vyi/S7fxQVfvmRBbQEf3wUaIuMWoCC9/FwYN6kX9I/Y3xMAgnYeiEooXE2vPTKoH
kloe1NYo9k6xDw+aFfy2BkJ4OSNS7F2FAKSaxSQtEqRf8PS37l+1BeoDEquU2uVl
0jeRlNa+MySTt90a+GDoGGU+6RcviQG/+6dm6vYNdWGMaSHwVCS2FnQN7aMy6ktt
oXCH2fdcZ/PEAsgf60s3XIIM+uRCS72DNyHRNK9myA5tWwroM2er2Ob5C9ZVSMHt
vcYz5wBoGOkl8wUfd4hhAmJS7QHG+KYthB+TdBLC2GRIJnkSMdkJAcH9uYBJzA5L
Jq64Qss94MP007nCrF6iTwwX7tEumw2fgoi7/vPlIIAicUzsPxkQGzpAOcb1ACfa
p3izId2GdGNqoQVNhupHSTkxMkQcjhMnQI95VfUjDW4FRDCdjjNQ5Jop4mYUxyvu
19/lVaSnqup+14NJCfeqQbrnHk8Wx1OPDGcSdYRNgorooKrGASDzvkQwvdDBupY9
bcxdFN0rDT0QIQKo+RIvmCkIvDPx33YC2jbsXCMiIKbQA0kFSoLo7sSGIxszIy6+
hxHq7suf3NvroP4DaHaLds5xAiHqkE14HM4qZ501jl9In/rBr+7HypwPWEBWcA0L
xg+J+sLQvWwOOedVQR0vC1FXxCM2RULp2WbIK3rH2bt4seZU46hwbKS3AL5oHLhx
Zld+r7VScCu8EF/uvbMsdtXTMdUhWQCpfcVviKkaewgpSkSno/rv1BEZBdunVKVK
56zPprexQ8qtfJutJ2RbB86KvDaf1r09UHLJC/lDISMBdEEhIY0U16XisWSpVa1f
uGGGH5AKAafa/UCPMcgwHnFl/W53EhNr9Y2V3v3rFXF0Hx4039glQnNhOzzScfoo
4TN8cHolFDQuEGlqW7sDPoXD3CL3nsG1jBWB1+kOc8i2+OKcWrF7P9W639zZSRqP
`protect END_PROTECTED
