`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/UbaDz3enevaCztACvI1QH3eL5N34Dgi4UN+lCZyEu8nQfJovCDVk1f67QBoL40r
DeC8znzIAL+Z99rbdKMVRFzRUdrwRZpn2eDoT9G/u/X7SBVkFmOeM8XYQBEOi/4X
Na3hZueVzcBtbKYNLdNMiOftM8f/adMeAyCvYaYyeyYfIdbU2c5++LQauxr2TZz6
WrCy+s1GZg1ScN6LyKp7qOfYG3Omac/CMupMovJLXvheyf9yfXHXt8D0gcL/kI59
CIYLPTzVnsXqvVqMGq6NK55xR+4ToWLmH7GbeCWa6gctHq4evao/RdKp1I4xgbqU
d0Ao22+feGgbeHzSMubvi+HK66hsXCXTG+qZhHLuyt+AAhvELO/FC5PUHnO2hgtG
NfaIALYIwr5BKRpdHmIWZ1mMODQwLJulSv4sR5II3/iZRvmnxTQ4z9WszygdpAYo
JcQi7iuRYhsX1AsSboYI6+EI1KNYzekCFSIuFOi0TpP3xCpUqJWrCug0hNdPP/HB
Nsm/RHKxcBh8arZEBsAWb87VzukAJmbfDXKJQ+q7vY6gqSItP05zkKt4cI++IdL6
nZOhXucqtwfvNocNtMCgtWq3j08vy7c7C+DCGuAiDncPhYHNszD5kxlAGc1T0aDi
d3f7uTUj3jiIzfYK9vGS+NInNfhl/mc6D5k7Q3gcLZUprIzVD1tgRTD9omchQTA+
/pmV+yxhlDGb02+Iwvcgw7gEldEwdArXNTw2kli1wXZNKwt1KC3jA/Qsl/okDeiV
SXo/K0rZytB/kW6VBRYN5mjyNK+er8nZsFLrVNxwkq+hV2kL52BrHtjZwMvO62DC
t8rFCeH6GrAdtm2v0ZijUxTz2/IRdI1osKbZ4M0lp6QTJQrZwOIIi2z0003Z8/jF
pzHtcz3FS0ps/BOd5tcvv/H7N7vxSyqjJgjNBD/VSkfm7TEoqC2OFymooY/IRqku
2oGxelgKmCLOHbVrgzQh9qkX9vLuFc+lrmkWZqRlCEyt1yj9ixMjxGmXohON1rX4
87zvYBtCxTjNXMnrfLUoeIe5uG8hIGH6McbhYzjPAlQnf1+DwxQwMM6BuDTM8QVe
pOBMeHD1xN4q988s92rUEGHC8kat2oL2ML1Z9pXLfEsrXYyLOLolYkL49vy1lyZV
Aw2s4jyDqwcEMDpEtRLmGjwdMoQOgrtVrjeoNTNp3JATrzCClELeRuA5Spcutt4E
F4hQLTVYIj3hw6C6Tt6BRI7tkq200CvMdwD2SDBeAH31GhKeQjYur+p/9jjyeyu0
MMOPkhY02QdHyllRdnKenjSgHKC+bgJHthfevu4kNP+Za9NHhXzfZMdqFc4w9cL/
dtk+QyE36yU4u/8LTQQ/a4fxS6YBzI2nfCsHcCL+qLhrpMHa1nP7K9wsBcnAP3OQ
gr9+aeRQxNpP3+BxV0GV8Cm47/zHUW+xyQwU/DSHs2Le4JZkdEFOTA38c4aOhYQT
ZwfPbUBNiddfMuGFFgPHr+EwZukG5R1051Fd9FTIuzWfauTR0wcqsddj1xoJOWqa
65/Dy6iYe8lLuZA/BI8V5TUmo5OQzQ8tFEIrgaU/2uXnkb1aRZlKyTcTk+HIH6wS
rXAGRybsrqBigIn0OAKZr6FeupitTmZ8yb6gub0+R1c=
`protect END_PROTECTED
