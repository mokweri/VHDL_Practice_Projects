`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lfvSyAuZtd80EMeWddNDCDfWmSNr7IVBmD0fQF/NrRN/OuWk8YAiFNcamKJQ5tnf
VfN5jYwD+306r2o2EZe6NMRX4BSa6nGxSgZ2KLISdwNSdwsjx+3vgMkpvpkOudhU
XrRoOMVeLwxcTD/FmYs6NGbWuAA8cec0O25eR2ffaZbCCfrmUHRywHq/vbGF0Ywi
lVb/Utf5V/YU+ag9ULWLT7ZlSqse3TD3Z2BxULa2r/j5fzv11wY8eDQV7O3gCLm4
cyWCh9wFR3FTJbFHVeq7lKE7CpSY/0T0DOID9pkFnTCshu1GhqQHpZeAmf3+6ces
hj7rsvLUp86z/9rLtMK6TypqogIG1b8+BK3hyjFitqioZzmIe7Jj8tfLnpsM+Jn/
x9y1O8sX+JfIdktuzbWnE5B46mM+X9TtIm/n9aaq2OgRKVp8ExUWhTWOpr144k9K
uNsoQgWrpWO6dGVCGRiI62yEoxg/JbfQnjRHF+duJV82qs8kuutMTLkA58X7Ozhy
uwyUOCBr1zpr9xX8T09MTiDH+cetJvFv1aO7BSQXxuqaswEwhQx8dauyS7S/aOkZ
+AMz3nvKnA4UGN7439koBoB32ibzm+ZJzgjU24OkR6ssbB3IFcTDE9uuvzU8Zdrz
sEMmvAlj46GhzdSHLtY/h8ZVWskmLMyqMuCIRMzDWlsQjBV6u5pgbhEIt22vBxoE
`protect END_PROTECTED
