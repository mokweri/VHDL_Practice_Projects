`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmLFV7fA/R5295rTfVTkqFR05VerwJSffOpGwdRUAIOBrHGKcBh1d4gQMONntgwl
MSBWYvqo1ft9A8C2PkdiY+Ma1l2XTDA+B67aH/hpU6lvStcrkPcfjqpxL4h1eBP/
KPnVcDSCVN7z8fJUrtSMtHxHIiRjHlcZfrTHU5JIogeDyQF01IsK9rVNvngXrEqM
GP/EDlJ6P7SdI5+kzAaqBjENmHQqYKtW8rLCx6slly91zhC2TAa4A8BT0w2XqsVW
/shEz3cFLkrbuoUfRKt9KtXvp7msTMKWXTWHzIcQB8yuyw89cMgPNJFb3xeIS3pv
JzCZswUiMYD756PrxZOYBeIdoeys0Rvwvky/WaaHTa7RPo79I0Z1DdWuraeV0E4c
JznPm9hFZwLIFOkL5x3Ozj2ahftUqCi6Dt69Ixd6OI9w2NdiriStj0X7hYOEQu3Q
htLlBbBwqxBv3DAfnnHcXCP11Zs1k2lKLOMsO6isGydre/TOrnaR1FQfS6Np3LSf
aJdCfrGRfVEqUFOL0IrdsAG3SxW0sHxhuVU1CqOiI8mn4qVfdweHl3Kn0Gsy5OtE
6UkhYEg28AD60weC1emktclKnn3y3LgJgfi7E/G2ekW3U9NywXJaCY/5BfZUqFBN
I64NH8s4eNuxh4xACYiPkWomaXJuUFYWFTEM6POPDGKfvLJVDXO7BzRj8Zhx/gZj
b21+nY6ZUTURXfzU2M0ZZUsfY27iVmrfz9i6aFDCtiQJiyaypHsUg6tJ17cmHkz6
9wrRTdEVkXze1kvK0MFSH3m05jdteemzLJvFQ+YjzyIfjphe3hClNxm1C1cHiX7T
riqAsHTqOoXtjUsctwyztu6r7dU1U+jdOUov5TqG/LtWiGJTFmNoODOgaJxa3Xze
b1dTv7+Z1EsJ1qFj+t4stVQZ9P+sjIDH3GrouKJKswfOs/0BYPR02S4nRzSvOck5
QB2SAXorw6tk0ylFN0pvk4ZTaI5HqQLKD6LRheVCySnVFaBctjZ7/q0cWY0ylZj3
mm4VgXS6HcNjrYABaIGXJuREsMLTRdRrEissThfrIvEcLqNCAu/yi23U7/odiJHm
OkYYUfIT2fcGsHgg+efi69iekH1es1GQ4pM5b7OjjHU/xsH5yhpctIcT8IcbsoTk
iqnZOn8UqUqimI7cmKwTmGm+pxs+HxPdZ7JIEfwL5QV8K1v2V7pLWCRwzELBFklp
u7JtUxSI0W3X4eL2oTYcDjbtinYwHjpGtpiCCIZNQ9R+0WXC0cSJ9QTvzUqICZ5U
txyk52278sPDRqahBJBD8/HvGsHft25iSEXJoQrT0MslzTtxVTGvUxhGLHamxtAV
tXqg2DkKpQP5lAprFn+QCH+z7oSAUdKRWqGD+WLz+fh5x4q+Oviz9kxA9cGtid3T
LMMpxvh+fFBjSaUdeRCGRV7TQJ/KfePpLj08fpfgsaRZSpOKng22QaT5cZcjAc82
B+AVLQgkZkPIZpgwfx8n0MBAhRnfZ2uLmqskmv6+344swz4QKbcY2CoM6j5oc8sh
z2pUR4totBEKcekE4R7N/8o5FRw+suN9EF7cRQlieqdTH2Hmxct1ZcOqzg/jn0+1
OVwRdCcKDVcbmpov4lbLY6p3uG1d01hAOoR8d+aFYJpRw85jT54o+J2LhvcjYQOv
BHCp0xAB1Ckc93Q9YSqE3OKI/qruwag0LVlKin+St7wrJVShlAJBCg9owb9RC1ue
tVEmqrJlmDRlN1bsSI+NNuak/Hw2Cpg+mfVRjQ29SPHJbLlRxwrwgl2BURAkPXau
jfTeKfUvp5WSHB24fEzBVLs8iE2FI8fcVWGEQZDfGgNA57fZv2exlwu1B8sYRTnO
LfZ45y6EynJZNegW436CBhTmxMcnv9s79oxwSTtf33laPolasLl/SqRfGyxtuTaZ
w1mWgMN9NIP+nt4834qah4nav3zvxPfyaG6tYGoUptBcBhA4ogWze55Fu3TlQhZx
/0YNDUu5Zial6kv59rT+SUmrpVc0mA89HdEUIAN+TErOdI9wZkn3OJ5stzBliSdE
py0zqhktRoHPNEtNz1FNLO3Fs4dreu0eSiPVa6juBzPLgRkumYGXh+IOlomZ8kPG
4wlatKqpKhG/4x208ppUCgzniKmL8osYcerfBMsKmcF4GynsKsAU6BWzC7v0FoEw
gA6jPeb/Z78GsdB3NHiphATIEHbV2U48HN23Ny8hgvOT5rx7BJHh8TSD1o/zEh/y
2XdO41jqA29u/hOwka5PRNny2levh1v6I8Y7qUr+90r6hal8Bnyv4JIW2BoVnOsb
+AjEZQMs1ng7fkOfwdA5zgZKaeuYHbdxjA/mEPw8AkvjzEOMQCE+kY2zToycfpmU
26HdZW+Oz6Z4H95qvENS8O00Ja/Ix5UidURM6sAIY63H6KRV9Kdex1tu+S0mAxBv
j8vnVDujv94G03US7JGy+uaC+GhECXI0z/IFXh3STZtnr5swX1HVzgYv8XgWfwoI
2kVTGVGnHE7cyLGNBeENDWkwFVpGuuhKzA2B9uMKndyFvqCt1uZEbApNh8D28vU5
/ZYejf167xjsDZW7cre++zYJXCzU7YiavmyjOl/95UWiZC1WXTifQXHTyzsxbX+i
mwuQUQLxy8ZYhakoeQFHGY51gOfVx5NrJjc/ndAmuUgiPjW0eClrho8w03LP0RMa
1GnT8PfRTZvDVv76wdqjSy/V1jq5cKaqJndd17uqKUzVwLxqIFixhAPDRYO8IDX0
CRGavdYOclCVZLI1xkOfbBAubrw6cooY2D69NziP19W0xWkCfWMMUNtXZPi+qSQk
/ifLzbUaXtsvAF22fdBELhJLP0FiGFaGP0p5H7vynyiz1Ga19x/ZUlfS9fl1+tz1
Vi8ouxjylvpZSSaNGUVcHqGGjvOJD0HWfwqwIwSl/jtWDpdi+pNm86ooGv5UsQVm
/cU9vMABYod4gNRCIystxdC3bfQY8lMnDXJUkAiXd0M2MHHgO4QaBoxAbeCKdaQy
ekloXNneeGZNwx29NV6k4UwyKZ1RfkpmCC4N/kVmapPuuiEGNsEBnRfjfA6U5xkG
9aC5pHcMpXzJuMSCCY91D5ADChOLY8Y6frk08QSEgrGyS/u2PMtajS2kbFkeS6sd
1rBn2dMyvUsAh14XbsJn3WchnADPlfym4fThs6Te6VoN2w1b44R/rj700eO5m5hk
P+sWH30oT/kLG2UUfbx7vMxhdeeqtW0rA5QjEjNf1JcBZwzbgoN+78njIxfJuHeR
5qu0HrNNVvgNhZ2bQpif8oxFTwihuWvut62JmUU+KbVzgtDJ9evx6eHD4rlpNM+N
17t1Vz8pqxnU8twl3bje0WdnmewmnSFMqBn56uYegH7FZAFH6A1M0f8WzO33GTsP
kzrV659raU9fKi960B51lA8xPaOtAE5KC5u282EBmLKAPQY7t2mEBjqOxY950Va7
SxtK8EaC4dFTSfOAVr50AIgoarMTxcMZJ+ORbqTmxbfmYkaEuWUHNhzMOgmuZaI1
gsOQAz+fONPeZRIz5RKc+bMCz6xz78OMVUHCRzqiKvAkAumoSirdcilG5+LXcVsA
K+vzIwsVDyf4494WWvk2TyrlD0IdCmKrUSwVKDITJANoYPIxeJw2u4I4tFj2w0Tp
KM5LCm/gL1aTt44Wx9XV1Y/X0Wpp1rof55OJLEFUTN5xHibaF87MjMrEhN5YteZf
xOQKHEuFZOqBQMZ0eOgfJRjXipROD79DB3vlnD+2Zfehz3Z+E3iwdJePeHjHUSZh
YyndEK0g7WIxdApxA5WXSvJnT1OiQukMGPNsXFO1QrDyGAFCOyD1jv4AHCLq5pXY
kcXPjNAymuiXpJqDq7fmKf6+aiaiBjgArquww1jbTyBwxKcGZW/+mW0XE0UuLJ6E
vbQgpLFb79efjvfGawKCJI8YO2YDuV3ZTCErBr/ug5raa0oFpwJIDXoAXFfJpuJv
hoMqSxMIcR0+Po16yxkHPEj9rO9yfUbAM0TWoBXruwtAwHzXnGqbUx70TggCx1y3
LPdwlKZr3RfVm04eMzmf/Dixucdisw+LiyQmXnqD6HBzu9VBy7XbPkDHFndk6O9g
DNewhPjYnUg67xbCrSG4Hw25EUDMSyQhi/wmE6LEg55/IRbugAfuczsLbPjIb9Zy
gXn8he3Bxx+Mj9XG69OL22z7pZUmPqEWKFMgUchGrCHE8JemNGQKucY5FBFkSdx0
dn1ErhwY8omaarWbXTDzaWWCrK/0w8l++OA5s03ZIxBO3r5z68rH0r1Q7eWIdb+x
xI3OgsQwjHelUi+ISwEkKR22mICHK26bZXcVZtiaiNscejnwdwQ+LhckwjWuA9A/
u4WNEIhqdmTRHtMI542N8tICPnAZ3CJGsSxdKynBlx/9vcZ/SVuDW2k4MR8/20AK
XGXUfZUmAAYkcM1pwY6u3XDPQyxC6p2UeWKwPIWP815PC/Lrsgg4Lj/L2+2TG/rY
V3XzeQykx5SJenNpOwoVTg+gnuil/Ua03fLbBFtNVuMId91VTSINZGGC1FzCgIT7
hT6L4VEur2KcZW0P2rYLi/enH0Oe8FAhLXYLJcA0HsdlFGbU2RXcgfPTNzKPx0rm
7aBKeoAUUDjDr9eda6JVeMjQTnFQwbXUrJSi2j9lMcoVmEbxoZnxSNl5MgcG4Fwe
8yw4v9vHiF/i2Fg41j7D+RCctV00p6hZIe2SxhgdvtNq3W/xnT79j5LIpNsWlzWh
7ZxbcMkiW32U0yrdUbwrPT5rde0pr1ux+u4FdGfhltrgajpI/2X/QQX299U0Jgzw
T1KJ8oxjA7OG5sFHjDU6c+10wRKGA6bWBVzvi4WW2eVSgVhEFK5Nh1uIqBv3x3tS
5ew84Enm31mC4LyHlInpsnxliKboi1jOf33Jml/a6A2lrnC6EQy1maow5LcTrTWr
AHXSPT9YfghKEcufjgOV8uz5s8mNgyk9N1babB/3rCC3Jg5QyDK6snhPYLzxH+UN
0/wxGtGAKfFF8BTjC2TRGOXamfYV5WEfEgv2DLkXnV0hs+R12zsqZ6CACJaL6Obt
nc18/XPjuoevvvpoUvFWBl6IIj+JmJrAMYRzgOfcDDq7SJ6J1UnGL8lfHLsz52rY
ctRHptZVkriL9vtAgVRWxqkDPy4X0Sv7Z7VCXx0ZRSixO3p1kk6T3msSu5FG7tKR
xI237HQWqjWA+GS4s9olng/fNBEhJUawxayzgemTj5HrllumypQj/D5BO9Wvwp/8
su1t37EleMY74gdc/q/e2NCrpy+3fppKyDLAcTOEtQYCmoLh8IJtGX/CGZJCh8PI
AdImtyMQ6UmgGmfAvXIbGk7Q0i7IjlDMsAOmu4rR123+PsIE0+o8HjD8uG8XEfxy
SUZox/Xak0bggVjXKYvUul4WfbVCYLVbUDYwQX+5GQxA2m0trcaSCRvMaVs/Q2+0
aYJK91nj0sWMEjjLZPoVkQKjNN7gHB+u4/DrAQ+mErub8BNj7Y1ahBYSkfS0VfyX
qGMTz7ASR0zcUUMAGIlyNBaR6HWVvMPMM995wC9Yao8Ae25ySPLbt4L7J/hyvEGo
n+CUmrKdKXYqLVMVxxHhaWqPcVVIIuuRsnCmstQDud//zZDfk81+BD0DOFG6QeYm
FON2w9swRySLGld83xZwdEdLBzvJ8Z1TKfHJKYqpHZ+6Uz2oEWcaBae9AdSGizak
CSCEdi+SUb0NpGU5YDZPt6oWh8ydAfaMqIvd9FMC+6XJUVjVfvAusmt32nUsFFFs
mTSCLxNDRiUsv+PkxRVK+tszeZf0lINHlE8CsARA1Q8J9oXknR/5z9frocEVp8AZ
agWovpfqxsb7eS3rU8JQe9Ug9/N0LeDWvO990aw2nJvG/xinF4jccFb9bB+sY+3U
0hdFXw0dRECguHT1QattejG/lqsITGrttfqgzJP47SAHJeAttLg3z4CB9ks1vgES
Ev9UNyQm+/g34AYiMqZQcxsmIcXlYneCR6bVvoKIxLetSBsUioD7BeUUaNmYU2tc
KEy8+Lqn5fRL0L2MhK+DZmLjNODU88wjn4gz+Q73hGXht9t5DgzJhmv91j5zmhR1
8JhbUruBz3itrxzw7NVQ0finEwgXafWyEWNqPCDo2tzJ3GvNCHMlv+U1p87ax67N
kXMXrOJEz8OS0ewiG3IE8NtGZjiwptNWwvTxJCISg7ONZDUi9vqL/JJcrgD+m9oU
mEJi6ndhPAJQCIMGdnXdYs4hPZqyBaXAjFDTzI8k4Fy8UtXb/elvIoZto9kMst8F
bMYVlJ6engeBiXFErX8UmnTVUkr6+h8L/emd7+2l1pdGGjJ0M/OwQVdvKSKf6o4a
NQsj/TX2wfg3ZgH/7VAjGturuHzL/5+ZafzXNOL9Cvz9JEhwaLJtZS7GMuFcQFEJ
add1qBhDxhUlpXUObVaOYHoUupua8pBIVhkz63LZ/9sJBwXHWC9PmqveDchUa+k9
zT/FrSOkM1Ki8kPOhyvTYDbfLJ7oa8fW3V/YYGRvveGQR6yBmfa/IHCs0PGKW3bh
9ghBqAckXE0sxVP7s5XV0hI3M6i6RRJ7Y2zWke1cnNwl9eL8p9b2zw5TlyvYL7V4
AmfWy6lTWu1OaFn2ry27+c2NqK5WYewt1K2mgNrt222/1I1860YtnM0ben+1Oaow
/n1cBMjo9eegk5T0HhGZkaARU3ccuzNwax9WIUxtwjNN7ILS9iN2KnzHxr/oH/m5
bUr+DEW1kuEUMVwc7e00GKgi3XMsLOxvHqazkHcxiugqC7FRXCnYxzWRu9ElCZzY
nqOlCA/3pezvEzgqLBeiTPTLP+0ZGuJmVdEOJ99Bm4I7P6ETz7P2LyiVDhDQLuN5
L5Y8C/NuQhVYG/WPNuH5Isu41VCfCJMDStIKFyYlJiZRE6ItdG1UxRSWSvIOyylc
m7lrr9RzmWctLavtdGu27rJHYX4D2tpsCNV5GebJWOLosO1PK9+fK+RUu+Eq4YY9
Djay7Yazp5e+1fHsaZUAXP78jtW1r1FEYGpj8uFYlOM+7168YidFzX5KJ6ig8VEd
IpsYc7m0TXkUxQ22IIibMo8O2G57efzobUdkcpjfv1xFdaib+A27qaGr5yfzxbKb
BH3yLXXJ6WbbYQDLQaNj+eAviVc3WQecBfHdQzvoot0Upp6B9YbXAGsubP/ACB+a
wsVsHofFAW6abVV65NcFwQARBx3YfaJfCMiD2oMkSptxreAes++IGuiZaHl1gOPH
B4e2Kgcz0RNVre7xYy6oNxjR904n96eGQEeSixEFgzRkqj61zM23dI8VPWG8LUlc
eJCpexoJ3P9it39yut4PZcMQwx+h6DTQvoVeqgfYz/bIbZJ48ku9cS2QyAHRri4p
haZhaYsusTPWXtmpXRMKu6IhEWrIisFZeqpflIPdJn3bAkKY3403GW2szZTcP1at
t50lp3lj3D04fumi23woKg6CpkNu1UQ2ccApEaZZYZ1fNZr059EhnWsB+2wgCvbz
SIRwrkW+OsKNpIgMQnf0JBphGN8vHYtrM3Lbdmc7pxGdyVrJSBCvgf7u9LfHAyKu
aNFUiXka9dZYJeTPQJKr/j+O31OcKHf8+9WzSnehn0JJPgnTcvmyE1Lj2KtOjyK9
LQ+Zuo9yabeKgutrlNpgiOKDE7GUwIC8PZVNpT0DGL2Gm/84uLNyd8KWgsSPAhUY
lqfshc731pWlVsOqqbhhiyqITNL0Flk1MZGpd2U3Vhu43ZWXvN1TDss6jRzRVOxl
qEpkPe6j50Bz22i19EqyauHkoSUvcSHgyjaHrqsl7k/hbDYSEfU2UUp0boo/tdHT
PT0zcOZk1k/2a+8hWlmUmaggK1jI2XWyf3CQnh18CDNbJTM5zA+qg36nGJoerFvL
lFTaL53ZGhg/F6mcdw+ke28MfgdTLC1kPYrt0ULgTFWGL+fdqWgdBS3OsGUdgeYB
Ig8rX0zZQwoy7UyGcayOoPVRSCjOh0lEs5tt6XeDC5x4kaPcg9mjUeEGQ5eGIElE
Lkafr4h8qsOznHtCCQALLjOChcOOkadRMrd7OJtZ4nT7dx9vhwpJO51VA5l7XLwa
VBKoRX7KxN0lDeJULo02NiWEV8oaULZ5MZ/Kay7peSEovT4ePjxKms1JesudT77o
7m2OVNxDa24KY0ylJ+YzG5F0CIDKTmAWV/j5HLpbJE1EM8ppMFbLgpAHHXSN0Ni9
p7nKKa6N1Hoy3XcH+DfHsFopmO8OW11ldB4a1no5jXntTpGnTJ9fbAswi0biRxNm
zHLioP99xQwufwyk4CF7Ad5S2N1l88EJ8Pa1g6d9uA4fFOeoRcpMleqgx47zpJBd
DtQpelH6vPiavOxqPg3sPDt9oBUD+Lt9y96k4dYGcgoQzjMGYy9EYfMLFwo62jSD
dG2/rF/HR6+7hfxjt4PHujb5PWn3mdGSpnGDoa7VBy4xDj/HgUZC/VpPy1lXAFDh
kAHqroZHCvReGJfTJQER+Gj/jFxm0jiwl11hW/+jM3HnshMuQLn739NUXe/F0Zml
XUxown+5uMGpD7q1VUPKNa5LM7HFAiuoh1nQDwOTBQ3INo32+qNMp05jufyRLJiL
6SMeciVYZOFfRPApX+cJ7DcXaNKL1j2b0YJCUTFJG8YUqqpmGHqO2bk1M8TYXaPA
Z7xNjSp8CoYd+kar1Spd0i/Xf+SdXZ/oai2fbPCOcQXaBKZbUgvwQGYju4Nkx1h8
aaMt0bv03pZ3uFSYJzSloP3TtIdO95sb0PLZGxV15Sf5yrxFkbGYR0QLbDsYWUIx
Y5lJLFAquUpkg3zVYe6KF4AZpvtUJ3IcY7zSVgXkLbL724eO9QbeY2iq6PZnj03+
iPFxkWs7KuoId7C5VfodouUxWDCjFejOs0wUxlm6pokHo6p5iYnInQYe+/3dTxGK
MdOxoFKk055zTaoiVE1kI3WGgX/ycurRjIRrXfUJGRVeOi1tJ3zjmlDW0SphiVWR
nOKDDNVg8aCkZnZpQc8kz21FSrgrxWrA1FyPYg60T8Sa7zwwmTC/NzEJrEKr5oDC
oCXE98xY1lF2pT9zvFsl/dglw7sl7lkrH9YNdEtH6OQ1G8rhlnXd2xNu2rVQ2LqW
F8w/gzhbyZHy0gD/YGy0wIqJNituxz13QLC2+C6zFlAyzQ+RCYvLNaGkJHYPovTn
9AK8eqm346Qa8fhPyPyXVyOBWe4kdNlf2Ci7tH8gYtlLnC/rj5mWk+UyiJ57xAWO
nl/YLRzTQiu37a4wt/upH8i/R4A/R68nAU+bwtISJV+y7uX86wJdj0aoHbC/EnA1
j6Gh2D56k7SJMTNLsCd1ysdm2OzayUYR1YG8ijOHsmXakV8GkR5T8BjOsHLyS9VL
Xa8llR2ZMdoHZpK47yt4uKmVrtu7FHxrXngG7wrUUMaTOFzIOsG1y6PHkdzvC9V7
pXmGtV/in7KaPinGTgLj9mGcoIIAd56+4xq0wqDmO5bcPhoXJxG8yJmHB1pHDeAQ
JJsan4wkrsu7oztEWjdnoJwMd16R0Yd3sUfonkdjh1aV4plMbi1s7l2D21JSEoHg
9NIVmf0Shj0kphzFRHs+SvIa6h+j0wPykbt58UoZYVrl5OjfHjHUeaPCae6XuTkw
xp95RUu6Ts1Sm2wofriWIIV8KgzL5vSkCpiOYIE9ZhPP4v6so3VqNscC7tZ/ec/N
FFt8jAuI3lPSw3COOkNqActuAkjmRMx2sPi/jHq41rWfMeCaXess+JaDcxSYg1Pc
LCHAvfL9kruAxL3enf5UlD5OvEFcCBeTGT3Wq2FopVnOaI5Gn7GfOdPKC7Dg0gzv
eHvwfV/7NWwZcyZfkuvDyKCVwjXAsr8KVYMiNGgew7BzudVPZrT0qeFPe7dVxef/
8rqfFItYDo9ma8EeiykFhaxxbhEJA0riB+iv+ETYc0zJOqUqmCJgWH7wccyi835G
IcNac5PP0S0AmOczbFNAk7voy2IQSUkJW1ro0H1MkDXXHvnvplojlmlqZYPOPskQ
pOMk9Ub0IT2ZKrbrNjikjS/qhOReiNMJrHy5xZuRYcySjrlF4XLTEu0NKY+vRBEO
tQbQh0LPVy8H4z7dUkqWvotMk47YIezIdrW3g5G89/F6Qqa6ItvQ0r/eDBDomg+P
c0SCYnAA9yQraKLD2C8IYfodzJ8+3Sbjm4mkEx1agC07PHXnV6KXYux/HPHa7SfP
tZEIF8YXJmtAIqOxkhkWeDoZup2INJJNX+T6dO2xQss3P89IF1+93nS9SLVC4+qX
KYBoKJMTaOsnZrBYQPS71ktIVedMhKEozo4lDQbFCu6euaqXcg11UsSQhqe29jSl
Neoi8txOiJWQlbMki7eVWYJ2JknTYpQqC/C2XlkStd6ycuzO1Ygdt19QwVVDpBDJ
pDQuB0I5Pfnm+Bf4ZkL9ZAOvjrHAgDwa57I401bnY8QY9qSo7akPl9qwJrawULdH
RwlKqjcQPpSrBdNrkolx9ABufMbUivXktVFD84KlfKZ7J5v4MeEbq5I3TUphc1fO
pu2bD+iLUWm64SQkx6CV1rhAcD7xiMPFhpVsy5DZONePFMCaUOxbY9y1V25qibXo
7rSnqgnIw7tOzep7Z3J32NpKRIL9Va2T1UWRa1IRZ1HRlqJfalIotbcFl96V0orT
vIldQ4J580EYXohVzZslyHx+OYOPVtHmjn5p0d3tl52mZ7Pzz/9PD2g1C+yNBOr6
grNxCngEjvO6RtlSvV06zUl6+EsjKyTvDIZXaP0s4fxsZtn0XEiAPOwaJBY5gAbJ
SHWaNJcljcUltp4P/MCV0LUtELTksI2pw8lhglhpHGszi8z+o9R3gznXqzY1ZFzk
IDeDx4D5PWdzm5TspVnaMkap0kSA6Vhj6xAhWaVEu+jPWzzjiSi2rzhNRm821TLP
svZ75+F8FHhcV4kga32rnTDTiZuJ+pf4wtYC7awmGqL6u37lXNX2O0GYsDM+mJ+b
Juc2yHk9jUTHoVr5yUv4Spy+RiYBILwwOYai/Tf2ge1VmnRk7YkTh/S2jxbZkvvD
0wf3lBz1mQpFeOdoEqGNSqV7livNSr4o0YmdkFV7w3KTs7fqGGYO7ooFMix77DFn
biB/iDF2RshQK8Tt0K9I7STrHkvSp8UvjZmRzkdQvmdnkWp27aR9qhiftUofNWIa
lkMzU+zOmrjcwvOsJp6cyw3DwfZumhFgyPJGTJZuPDqlI9W7Di12AlhN0N1WLEiD
/NKxyjq6vik+SCg1qiHGaSjioQ10AI1E4k2aRK+NGdCJkOEZ8LNhF2x/bGnyGNoL
CMAX02mx8+kmQjIffwEV7aKqcoEBspYXXT93N7512X60uFl1p/JUX3dJgnHzEO3j
ZuoJ/o60qBiguqEi1izUhFoWIWkGrr5N+49VVzBbGtOxWRtydG49QUK3beJkAqIP
+HGo3uqcMqzcN5z+OeT1obEGnwN4JLGQOdaPN8/urFRim45WQQXB6g0rPxgH9Q3f
7hibWwn/GNzjICC5SYrOUwiC4H/T8X03Z3RHw0au7YM7tgCGreZsNUX8WE2fyWtj
q5K4Jwa8dzSIl/MWMH3fi0Jymw+BqyriOPSJparTNutpp8BgBHTxf3/tmecOTD+j
YOnst7fflWo8rQqz4bPZQlpTh5OC2RM2tRXvgmh25UFaRwBkvH24rOrjyzKL0Sle
cD7UpT9mwcxCGZiiRJzMH++VUUPsG2dPjCU/NYC1biByQwY5VjGUSVI4AxV9CmOv
BHDuopv8gxHo+1hI9rT1pJ1Z2xiD11w5xGwA1fyDEPf5iYmzUgrYIWrKROv9W4cP
u8Hw62HKKmY8E0KSL2B5sEejjdCAYDgg1jIPad6d/A5c1+YlnL0eS8B+PXyoWg0b
Ag9jNpgK2LywQPdM8SZiXrPVu2tDRQsHGpIMkYjbqSUi6D3r/ifx6QBrbOa4DGKw
RWKKei4V5/NlGqYhH3ByLTJxw5yAWYxnjL73EL8hUHkyz75W6XZoCXeakGcxeSJQ
Ual5gSgHFRt03nUEoxai+wg+Wjbk6nEyiMSPlZFbeHRkVzz5mkd12ZrLlbmK3huF
bPpeYDNxxevVvMGCvtN9sxUGJWectwt/JwPDvk32cdfq6DmotgaSOB+164cXpV8l
zZgnftd23narl5Lt0yU9THHcKOcbAJNlGApVRf4PIrsguh0qRsZmLGmv3+ZZMIaB
mT86Rt/s5+PHTE5XlVidwiM6V9Tv4+cdbiM/Net68UsuRh0EIEq4ORsNsz4eGiMv
ROLLT48eiyPp75irt/X6dC974Ov+C0tQW2BkJW83va9pHqZT4+wRkTlSnqq7zQEN
O3EjuRFQME23hh23Ij/kof4rtOq1hr9RpVZdz/b6yjFxrFUvXYlAGJfg8YMezyBJ
1ev6GbgbkmEHHKwp63LrlKAQCK39HpEO54jIvT9TAUgnDxugRms1cxBdixueE7XN
G1HNaOweEtOiPyH3O572YvTxW3kkTeGw75nvLscggLj+wQHqAGpQYfYn2i04yKTm
uK8wNDazLyn3voMDMrTmTO10TEkRSEfcep6LjhWByznMAMf23iFFQnbzRcEzhwFz
aF15l/ZJAa8uFHGhiUlUPHvdDUMv/PFx/1zfkISJBBVNWr3d0D+1iJ4hqeUS0QtU
a8cGkBR6GGdSsK3vTdWAZFwFFxVlhoX8eaQ96OPNYyCUkGVUV6hmcA/m/QfJQkYy
SzMB9XRCBt5NdYyvZhP2LVMPil1U4HbAkpcZP5a6EY+rimcXqZPxdqTnN6RAdPgE
SHofb3QlJLSjk3gWA+DSKKeJYAlZW7xLH7eWXoBN2XM7CwZAHOn2/v0cems4JoiV
NIJXEkiXi9R1VRCy9xXiYd7zCwLdRFKjU0NatsROFY3HUfZmUG0hH7kVRSub0/70
oQn2VBKIqYzftEpaJPNTow1i2cRD3j9lI6n9zYbHUckQdiZjSdg9zBiBeFWdz/jS
Hn0F0hY2C6dvreDdFsu994OTvn2a/CbLmR+NXat9m0pTZ5tTMwq4NS6JN1lOkXWZ
w0h9oMNGXDVzecoPQZk+VZt2kkhsCiQbV7UpEMnlCSyblRzv2s6Ueq71jz4yhPIp
nmLkGVeSTkbswWy9EdE9EfUmht1iQlUPZBFBQldhFsYN87nyqPBQ1KJvm2OHPgJY
vw2+eMBw0SR2p9wf8AHQZBA7c47XwVIX4TvSxXleyU+6XsT+8dOdigGtJrhBSjS6
R/e52JHKzGRW+TGQOfyUJt5Dt70fOrwLujrNP/1FyyqckQs8dLb+3CRZCqbGkcXm
EVdKMqPDFsviyte8fOV1BZAmYcOB+ODgkE48SwrH9n6z51ZMOMmlT5VsIM04LUC1
69U3KUqcGXH4fPZoHlD/3ugjvz8ZWhtXPdOElM/UP8ZCqKBarGdC8T6uXjKDSMr1
520c2pv3h2RJA1T6QucKIylKk+mDqrTsYGHpRg53g8wjeZSTqZcYRme3xS8TaPbW
sjUQzvrH9WeuVbmmJHLGlhFtDUCFEG98LuHYQvTw/Mc4ewasMzhFnN7uhWZMVM14
8MQ/ecvoVmApaK3oGL5E1+R7Q9NDvI1MDn3A0f8oIvAJo2s/TdkuKB/9tmIfnj4u
E4uo7c5lYlfdzNwkv76wv9nDKC6iF4bOCaWzSxsqWS4oXVgYRzhVZiExMogbP1ib
2SKQ0x1l2blSdc9Y+gzW2WObTr5RbxsxcHET4LvbguoJ4TjkLvsd0C6tL09N+6Tp
rZnWWkJjS6zmTWwTJfsVfu5hXueiHm/d2S9iAw/v+cll0mDeeamwIr+t8xdv6vQv
zlilmongfkRuOvJy845BdhlScAo9XWzsA0UDoJsS2wmltCDBjhOLJvLW9Ok1qjuJ
k8ckhWZHtAx1Z1CHBYMsNbwugQi3lmjyedBew4LyML7gs9KCtSBTs2iifiKn9k4F
EgdPapXrl5xsCp6EDSuL/RlGv+OGqa/Ozk1j0s5zp8/Jl0tBTDkHSXVN/o+Vue86
7jue9HrDEp7uTkkNdgOteYT0ndjqmxXqLhsYpIF1/D9IxaU5QjdpPDHuxbcyPdV+
V8U70x9tVZETn10ZZH8TztxiC49VhUo4lZTV0liyg4kr02SkTMCG4+qAkL3eqzbz
F84Rn9XjufVzMi2oKAQFMiLuHBo8G5L1a1rEvJXel21mc6yN4W+fgM1SbanAFbDY
d+xZtS/bdZszpLaBrov0h6ZwuHBUHhIOM08QvxN5Hy5H1+5oA/CnIRrCareSw3L0
BXCQi7/1kaGJQs0dgMdZwBSCQ+ryU2zz5q7PUDD9xjL5cZeaMkf8FgieNihDOBiS
+c77k7wAPfZYfRF7iv8r8i/NUR4EnpAhBBnlI3hSZkqy1SaXOYQvHxEXULWr3bHl
KzeDCrkY9QrRqZTUIfgoP6ufCCQftBf0Kei7BoJKVeGOFTSw54S/8ppcmIr/87aW
KldZ8VkzdBTKTIb6KWtY8+2R/Pk25tcvP4NdVtYECrMg3Q0jk/rZmNx7ThcOZ2xm
KMCHMQ6mGpR90Wn93li1uppiL+rarcP6ZZyi0+V/Frpg5ZgKh2K9KDwy4Jk4Zxza
ZnpigdRvxWGqDft6d6vsivH4ZWKzB73qSySgJ7Rs63F7vU89BfCBwUn9I9BDNzZa
QVuHFPh8xQEvW6hY1i/vYJ3Q4Sf8KYXkVoJ4SXIV6atuDE933LzhKQ1/eSV+DJXD
9nCGcdrRShkp5nnUJLzuYZUPV3QkhZLIKkoDbIDL/mKVBSvJfyyGMBLJELOsyPKp
sPQYoAXo404oCa+8kM3R3PGkDO0KjeUeACS9ZbA48GX/hxQX82NCsdLUh6YF9eRT
L2k9K5kTmWnZArc0j7hsQrryC/320UkEfeEHC9U0Q+SOQIYUkMYazqZmkvFyEi77
VF4veGfj0DfbCyNckL+hf5OVbWjLm3hJPfRBpQVlvJiPgmv3LjJFAAPxWH4JuqNz
zmn58/1AyHPo81GlJszZoD+lWRcWgEZBGHiYctZga1vyta2NThb5lRfd8afUmmbg
I/F/EWq/FyFLI6zzCkj9IvgB/cd6r4PjiYNbbxFuMb+Yzz1a3JfQuzuI/BcIYvc0
OAT8RX+q9LHmkxmtsfH+CEieZLboqcanlKKFXL1dtYpZS5CM67wQnBrh6TW2jWp5
2bNxof5t/PyfKrSDDmSQkhWf9lxKY/fIMwdzS2331V/Z/RvEyFBQp/Et6QRzIneu
9h/yPPtvRdt52fYsLmP3/VqLAl4TKD/oLvxEqL018Cr+9Xw3VdTPfJ8UVqqTZTKr
Sn8Px0W/ymRLMmJ2jcdOl4SSmkobKSuRW/xMg12TnPbzagCpp9RNyKrksmApBU9n
4kD9dqtIzajhQrq/xAYC14RlLMbVfkKdqW5KNd0ehU1mqnLQL/E1qTbIOxvWRTme
azPZLOSHI50kLtYCs7ysX5gn90AWj1PUFBm5b9UCzZ2xCH8fa85pIqq/6TKlRfj8
y2i4Z+ZnbEM3hkTTF+L0trw9G3YsLmiteNiDY9G6kwtog1U4kyoHnl3GL2xQF9Gz
D9QvxhPHDKjfzFVLMkRt9SbFK7O3fXZ+xeYfyQQXs5mdUXt4mtfWH7KvuWh5EizB
Dt8G8mCnXXcFfOa7GeTUYOIA0rAtW3+k4FlhnI+Xw78VnBkmRHybj4QPG5FvVN6V
42MkqmsqJSuHLGXr7V43NS2lkdG+7BLrKAZA8yxfZIr5xankibWwcxMpUTZAiB7j
XQ9FQMoxxK8q875+zHm16aW6aW/4TGIBdaBT6Q1YG9488eccVCkZGnjYZVwOmv2M
ksQVkfSvmgr/XErbnPPNfC3pZx42GPfTwd4MKiUnhAhfaZQIFLgc1N9IsRwcrABl
EbppdZsrd1KrSOsWR4mY7a3SVnNFiYKoyED/DpfuwJ03HxlJbWkgQ4ADpynhLEwi
cq5uq5SAwTrXrRTC/N4501oZ/V+qNr8EXhzKBCOEzy0jmu4jdzF9aEr822GPoPM0
7G2W1nmWqcjJbq1PGx7BVT2YlSzM2RrDaSzv8U9Nl5GkDDY6oMO8gLKvLV+xSPOv
KsVr+OnU9hqyPteRIy49W1IngdKKGwF2g5L4mz7TtVDbLBXgHrQeBYMfwj83nxrQ
AeVXbvvlggSOxpoVSHoB37QpEXUl6Y3hwzcSCJTSnF8nNj8x6piGfTzifKoygqwc
/5+u3lWhRBzpzjKC3JEDi0DvzvsR5dyq0Hry2XjuQYSQhEIpgwYRHbnqR0xdNE3f
sQ9TmFqysBjC7Apf62O/ToD+CsSIkXU/Mh7tJJuce9HAeK7goZIEg43X05Shj/uc
sAirhKF/Ch143aMWoGN5NtS7Y6CjqY5fJuiTyliam2DrMDuUXdW4dycvhyLsw84A
Cw4vvenLNXnsvaiYkSo5LXozU88UCzgjG9kvy1XXTK4GBhcnzj3bVYpcWuHijWlq
JRpTe4kG1kOjp/aGpMer12rUXZCDZQLNb5punuHrZYKRDGRqR+4ZwYgxbzsixsxe
blEoQSFXNdHb20tYFcz0OBxb9lSMovU+lbx5hOECbHwAcUmGiZ1hAuIc+0g+c1Ee
vZdMjIEx/cWKWSJQUAvm+KUnqee0g74Es8DhGf6dNQR7L/bZdqtGLuPJphDzu4S/
v5aEQziznH/yUVnh4Cg2jA+RSJYHk0YkcnXKXkDtD+z25f+daFbKDUhPakS18MGb
7D+ZxZWvk5qg9M75efEfjb7P/A+L1a4tCC+uSAjmLlqsWUrpprfgId2x799+WnaC
qy2PJcrxkQYg6oHfviVdM6dm0DD2zvgIOWqD1S/70k5GHi59Hb/wwRq+Kq1sKz/m
Zx34oM9197paF+mcBP5l3/+eh9+36S7i54BuskFWTv4vnXJIzt5DT+AnpTz9Evj4
lulFEGJ41DW0zr0LAwEzngYUaR9k0ghk+ZPlGEQIMkiuziRc2MupVe8z2Q8QYgmJ
MPQzqMytb02WxcwJnug4D3OwhVQMGYvYbokCm/dISogM+OhnBruPxzmSNziYIagL
1NaF+Za5BJeA04egzMPcHmGOUN33DJMoMwQjJjZC2lJdzyWk3UzIF2NNbFf1cPaM
21ck9t3ZaavS+1SD0YvSt4/SQRb9gF8SGMkaLNM+S0ORaRw402MSUcCfxwcubvNA
UQROmXj0hYTLYjM1bh78Zo6JKkiU6s2q1ctLfGjhKgyu0oewFYepsaYZOduFNzvp
QDqsIGC0vhJjjsWEMP03qKp7WO4panko4nZFc121k9iSIU1BWVqEkJR9hiPgq6cL
eqvmOEcru5qrGl5n2Xbx9Pteu9ali539xY6nhyNfEKk17AAOzp1BGLR48Kj9h+tL
wmkgBoggWc+h9laeYbXBugTJWNCaqRudxi6g0NTKHp4QEpkpeWpqij2G1gDZbKK/
jKSzUKk8XeAxToDXL44fAsQNY13b7Hahpn/AEaSS3DFUIMMF9rQNN1Nr69/MgVWt
0lvNn9W5eV/32w/SSc7u/e259lp0PzdFkrPlBFcgfdr9DLHO46BWZj3be1IUa+vl
+YGp7TEJmftfidSrMh1k+a+8X/dzO429Ee1BNxWmNy0zi7oQ1RbRPs0c3oaF09wr
o9r7EkbaVH+mw0xUHQZgWG7FV51/wAYxmTqRnMZPdON+GXTArnp9MaYfUumfFC9w
V3nu+ONEGvAnob7gvM5068bD2LA4rCyyI/vHcrdE8hQoemtlEtentBZYUwjNvxn0
zcfnA1bGdvaUrGSn4VYqRFlYEf0baGOTCnW+aqRR816gaGY1UJIxL7Oypq+L083p
mkIY2B9xIewSdqFPMr7VXfNf3xYse/jssuY1kv6MFo94wN+eSsctsdZmkf2AsiVn
XP7mi+H+Q6MdFxyk9eT0NCBu5MfoIva2UoVDh5HkErMDRootUpKYiNJpxCVybyYr
K2SrghXVztAbfy+NmgulgWvKekVbQcWGh0xQ4eT1B+XFZBiDmqcA47+J7orQ9kTt
9wK1AlX/TNcAPi3tlRiCgFK+1kt5JP/aHTldoInks0j3ts59TRnnEbH7DWKji4cB
iepw6UdZ74hkgqtyXrmpvcXKae6ymHzaDlBfakuGLinUCeUuPQ65e2A9+t/QEUtQ
72IXc3VSQHygOqUfZ41kesl4Bqr1C3kLnuNBCr59fOefGJn5FYY5nM1WKSrDhrTz
BFj+L8iAgeF4/QpueFNQnY66+PWCA3nLXEj/62NXD365f/csCQ8eQknAKdWX5Hpl
vH+oCp5y9eqs0m+4ExvaFbv66GWwJfcWAW90Q8n4/iZFHMbE3z6MlZUl0AZe+tzM
jmoAho7NlUQf733kbul6oIAzhJR/8FhFzHy7pd4J7RpwA4BWMwRQJZ16PzS6w00S
7lnquqtSGzBy1OftYZ/90bL7jQYXZL5wKPWlZStjh0uBY+62qvrwMndC+jmIl2eD
g8dh11oZf9/24jojybBiKCwm1xwQue4ATWlof3pJBqmOw837/dgUliW/zaNPsWzx
MdDOtJxvYMG7YMnMS7DrkzVDAA38U7GhF7yunlpVzOlXiU/5AKQVsh8PMjkACRyM
9yrZqLhimxcUo5Tm0fmBEkswO/5f2Qj1+qubTjihtUXRAiq+9VWsOuSptF6OGLcz
MWp4xBmbw/BY19m8DyGFVch6MqDWeJKyzb1nUKLZdR0TYKA+ayjAsgBlSESEEnok
IxFTc4EnVisAZ3z11w6k9QIntCy7setOtvt+dmuZXyQkkpLFZQGYGW7KxSlKVFvL
6tLuHzPJIO/S4lQuicKSliaLtvTjB8xbPYSmCpjLrQO1rprjMEeAsJhGxIrf1gkM
IpYFUmcEJ2suu0Bak9w+bppnJlQHj3Q28YWsder4ZNEy1QYofZOcrZyWlrjuwRo+
uJQp3ZfQUmQTMNGz1K6NReZtwxc3IjtEAJYsaGop4YiZMiBZ5/4DODn6lKrr6C0I
uO55LRhWMpAHF3kVKPYYQu52NQbvtkIg7E+AYRBoQBdaVrsbJfh0IY07Nx3Vi73q
v44UfXurOdseeKBUcsFKeGffXcyAoC0kysMvKwAi8cZsU/UujDh1ozC0T6MxEiZI
SrBZGd635KLX8F8EsrP3+50+zvlRJgWlSmBQEF4ZHotWwkURzHydUpqiRKgkY/6t
BqCshNh2reA3l63yvdqVf4fP16vGWpcjcEy3yDuCVv+Hh/KXnTKOremjrufFovf4
+sP3rcD4ukeCmD9tr1VTMaTDxQ2ZQxfHmlOYhAP834ArwgyUWLCQutMco4Mtm90a
nGn2QoQ/fHtxjc7Z6rdKKhwC3J6w2mUscK0SmUxFAouK8P5XTjCEEPWYSDKKQ7tL
gKAYp67sMPY9IFXJ617+9NAwbWGTSis/y5n16Jc1wBj6eo+ZF4gxbKr3VuFziDtC
+JFaMrDTnACKK9x4nRxM61uGHm92cc+3rHuANplC8L3F/k5Hgs0wI2baYgxwjekW
hf+NIefA9B1z5niqkhy6bUQVnlgwcADCEm29Es5YzoFL8zcU1ObJHwgpgs7QVhPc
crZ+WyAWh9Pl8rUXgexVN6NJ0IvxzjfqaDVgECOiKecGRPKM5oZyh9ZopTNzT3O7
djZ2o6zElP14Ogtc2+G24NicDKeeBxcdLtc+yXg3kuz3B3wevJFVwdohxxNB/UtT
XKmvI2l48cZRe/UAHdbvHJYnbJc0nICtPoycU3cTOUe4aCHn7rGyf+m+gG0OzkPp
xYchBG0hs1PApo0kwgRNw96LfJQUtsdF3jny5OLcUDxrN2lUt0G/u/+wDYjRegc7
xF92oEzVP+jaBdd7abTpqPluXnOhUv4VduqV87VdXx0/yHCrnSmbqME/Ip7Ej2tp
IRifWcBYDXwG2ECQWRQXnpo1I5zTPEryKQm3ouh/k8mjP/z2VKTo1At+8mlFRimG
/0T7688XbKT6b7AR4TPb+TprYmVQ2jIVyUKBOdPWysX8hv3+nPgbsrOepKGCmnrP
4Gr+7Qm0t0HvWOIMqCEJ+6b2oECjHbZ8dskDqo3ZHKvVI2+P1cIuhySO7Sb6JNsL
lKjbcTV1kbloMTr2dlkWmPNthGsjFSugDjx5wObaipTXW5mShak25vx1/pErzgT/
HmKQYu9nWAr6RxozYbyqdbP2v70CCg+7xqRPvOpULLp0zGfjwyAZrVT9Ptph05MH
32oT3ipHgHSoE54+lag5Yz1LAs5sxaXLCwiXFA+iKdXv6BufR3dSkyNecJFidqCe
GANQTeD4egk8Y/+LaBwv10V6nmc9fA2h8CP9p+8v3fFuma6TphUSPeDfKvnpc07E
5wfOeEkmRUaOQYdtQUn7d8Jw7isV8iswQ8o6kYG6Yqcn7/HiGL7W5tHCWrkfkVdL
yxchHsCEsmuQ1nhIcxjyDsnRvLCxUSKGX0Rl+RLJbOqgPZ3z+SzExDQ5dSkj24ja
n9xhrBk8ZiQur+OJUXxPpcbD+R+fpSJim3SivjLBBD85sM8WSl5iUmijRFWkDrqm
040UCDey2BsZsqVnHKoEIC7Hda5HAcX0urPv2bXfO5OR38tfymhkPDIR3DZdEOFl
5THO+FSQYaUhQVAeUkvt2toV56xyOeCNHg4soTin2WLYJ9T0yB7F+NvIl7rpuV/4
nqRGjr0Ybuj/O7eBZ6pPN5Epj8jE06S6dhVUbWkAWtJG3wnE07s6ZpfljBelxsZk
kM6XTwV3BxQwhrpmubBrk6xS5uPVG8E+0xqAKd+Hn1Dvo0OdDHW8N160YosDXkZ/
7GvZqiJxASmEW18nbLbfuVjJ3hBqHwg1+DCBRZWNQZCXsW545QMx1KNcZU/q3K83
J2AgnLvteKXpCiK5XScUcjExxXtsT3c+k5KeqTQJhROeL7DsdoJMLuJx3sw+JO+8
DPcvve8hn94Z+2mq7gxkvQ5+Hz6avBr5dFJoDZXtvJWkV19WCmtTjwzcZD2mcTp5
hm9m/s5gf7ofPCAazZN1BEK4uzxQ9O5VN6Vtvdj5YQlSSizCqKmoaoGQ8UiUZVOq
VWmuw5+2nJKVRKeeaRpCEK5VXwwNQkESBISzo2KD7dkqGCXs4+OEw3hxYdQvU0vu
f8qUqS+CmEF4qx2N8JOO8IClS6Qo03wP3yOWiX0W0K9Qr9lLNHpf+IZX6iVJpNgP
+bwnqhbjwKOw3yl5VPOmxIU1uzsKZg3bk2YMalEDlvtaTIHEaJWyT4Nqey2X6qS2
P068OBgmX0xmtHtE9SB813dR12Kno8l6ppbgGYcc9nMeFmrxhoMiH/Neu6f18stf
dMx19Ux+3wAS7UZH710lxXqyaWBFerKwgOyYzJECxpjwECl6PoEnuv4LnLci1ID7
kgvZvm+pdU4d8WBqxh3+Henb0MVGf4xsd0H2RKMSERU3x5/cVCAJkfM+Tkjekh/Q
Fw9Xc/C3toXcwjVjX5ozOmkAxtkwIcJJgI9GCdNwrYFOVFnfzN9Z1i7ehxmym9lM
06AxqUjudkMGTqVlaR9vm491i4aWyDI4Pql6DyrwjHXsvWyoCxwxLxyFx77uuEFE
BWvASNgpa3TKSeujPX2w7AoSLQd94TOmIjuYvka/G6awK5jPpdomrOLTU5lEXWTt
LGMFkpM4cynxsX4BehfDkHhKHBx/Pae/RF8ho2ZynWnEnvUd6Hod+xfdEpNvFkoT
LiMaCSgpT3YAg/Mj2D4n0go9G4PdE/bnCBiXbwGWLX0Y7Z7/ppQ+0gse8JRy8tQV
yKjD0tAw55DsNe2USHZZr1TSvOx0fTmSPl/NQp3q6n6GMG6w6ulpgcmyfDI5F9YV
qfBffpjOZ23Af96hSuC03puHnctEa3LokIDce2OHdHsAM+eeRsXDPY4cj8FmiCuO
xZBDymYB0IDwBZDGaecULGDAbcO/+8ly/ZBmeGZz6goAZgfBQ22GD3/kX9otqYLN
Hm6UjMlzAfK9gJepLxTbBsQjZWRqNb9mHMB17r9irGDXmQyCwzc+d17V6yhGCQ8v
7PZYlz8bgQvWn+Kzt3kXBr/+uZhyQ1hq2t6pivBJFHjbm6NKKWzmmhXQodnfWNc+
eRp+xdyGQNp93NW5U6ilKYAjg6pFzHXEJ4JvH7bgAy8mK27sS5N81kc1fczBKq/q
zPY1nMVMbIqq7oZE3pnQvnfLnexopNTgFXnilXBiaF/qfELKHOnJWqo8YP5cbrTC
zmNH+fB4KmixWywI9i2L3eGREdv3HY9cLwFfImXXxdvXV6k8UT7qvTAEK9xFAQVT
GMSVwZgmbBiDdhDoCaW5r9USBc8hI3MS2ozJ0HE4510aIOUQDINoGqc4/mBYcbrv
zq/ycgYFhiJaT7dNitEmGnu8H8Fm0Ur8H/zx5tWxyfhRgqw+CPAwVqrvnBE5tjhP
/afKr3EjtgKhekzH4bXFD8Kb3HSAHZ9GlMp4eh6EB+nKjNyYPExaWXi+6RaqmfAC
SyYemctY5YDCK4R+jcTMion25nLqibwXKlLBANKcqxcV9y4DFpALo1li+A8+Lt38
drZd34EsUW3Potmon/FXFw/1UW/6xU1EBVx+YSiwgUhyeztHHXebJ5zbYpKJ/ZP1
Yb50TbN6QwNXjuS+36sgVay+UN6DdQfi/q1NXnZfUyaX5R7PntIwgAtJaLn8SKGG
vKeOL5460niUk0+rvztEl9xIAmH0qzgQzGcQa7TVxil94PCQC4n2TbpWEyplnzUo
YqeCMR+2KrBl7jVhnFub1+tCrkupw8cZvfGKYofsmC59Df0SFxaFhPFrN32nVZui
W4bZA2pYtB7FubkSFDVGMxmU/ir7qZWfUMByS+J1/YFwqj9LUfsSgsmG/eln7Dvl
RV0wzQrrzW6uxKompdSQgfqymgUJ55y7ophZFLFTspwX+zx44VnAjqS5EAR1yemB
gdbII+MwnGt5Ur+WaCseZ+cZYDWYti/fKJMf9tK0eKftRJg8ZgWBIFB8P5/BHccc
GrbDigPy9cqF5u80tVu742vWKdEqGfklYHdcJCbxGk7folV1WCIoXiJBXMq6JSaT
0ck/oruVI/nXnkmom9EeX/vecqGJ0HlkQQYL43aSP6bAN10ao82f2HWmMhvggmWm
7F8pIdLREDXBFZ96OzHMNhiMVAbbgJjw7TlEC3uY6hhpyVUHVdmmRqW2ogtm/MwB
sBWdJCKYGBGfAUU6RvrBhCeGSQ2Gmt14HFa9BHFpC2IuL+d4RptMK1UqItHptKLt
GK33vw1524sb/FMm4mfevS6aGIK/inek2cvusEbpqkthWNbTZKwaBbKtAiefWzq6
VBw43CvL5P6pmjSjPkfm/S1ZKDcUbqsBIm7oEPD+6qrrPLI9/8Ohc622CsQiDGNm
f8xHAAiPYa81UGIT9nnVSgBbw1HwV0926RjckFbWpnR2S3qxE93saTUbkmOCU4LB
/OhiMBxz4Tbmsrc817pDrA7ct7HoVW6N6PGOLnEQXXcPWdIGxlhVIa1+SYG0QmP7
XOTZmCVRjQUNYjcBr8QR6sW/kxrLtHT46MecV/HegGIXrKRQb29wn4KjdwmyAozK
hZwIG5fg24X1UEZZvQ7C3wPp2voX9o4898pHOajoK2lmS4tosCEOv/TdpEtz4Ktk
Wf7TMGErnTVuSlPf0leCwL/pk1VTSW7L7fOZRSA05OKyx/VMzH4BL8lKrgT1sIAq
dKYXKplrnLULD2Roh4t1QZekvgqtwEh2a7HwnLdoPTmaIwpnBF6f2/1Bl6St4mb3
tBL2jGi3EQgAsqOhn/zKi2J5OjVsgeseyVax5jrG9+dwH2Cr5AugCMKunH3shve1
4VbFKCvuVRRFDB9UdTTvyL9/3xbJULSst52LeagGMeySU8vYFp8XT0G+hZmUb6m6
8n4axUgCBF6ZLLiDgU2yrffS2Lnpw0sU/4RJdU1SAKVJo/tfEMG13iL1DoPCkXbZ
DdLR+Fpg76A1l17RC/FKU5wZAe3uANlcbF/gEd2zp7NTgvVerDQMforwvNEKMfPk
B+R0cdTSKab2IFJNcTegS4Au1Xpap8nGOaO+8BRGB9s1bYoO5Eq6pOfcUb2PdnP2
WQfyRUXWg8hJlFudXcNDSs+rOUHZf+xeKlASpawp/lCS5CvKEl0JocrfZxstB+2H
aflPdzDVPPKJdha3DVENWOljF7C/YkyWKkURjW4Reda1GyEwawvH4mZUYcF/Kw2F
ArNh0QNv5kYz48TxyPruDigQDavSS4Ekvw+dYclu8OLXUW8iYLb1vUotqcU9YO7h
/eL6pxTjLA+M/WfpXkoJrHv1mG22w51nkFwN509hGTallh2HENhv7+R43hntMzQV
fmf9y971hPlE/Y2i6emaTm2rZEYm1mXiwWg/bAQ21tcJiyToc06hgpfEUQZfYZg3
u+FtsSL5ygoaTU5IpzidnX+N0hRGQWXJhjUv8FhdUk1edVYj5zFzyNfH8pnRNpqu
jY1L+Ph91Z2psbWKA5QZukBfRdPPJ+6QhQOOLKuiXRfLmH6jIWxgfChEbagBFtgU
3mCPA+o43KiLYcFUMA/ZcEtrWudxzdOAyhyHLUNRMTyOZ8JcRUhL4Akzp8jQUvE0
FL8aamiUy68+QRpPdUByscdkY+CUPe85NNrW41qfb7IJ3A51k5zImJ9SMFcWJAXT
31MeAOzvlpuiDdVYUis9mgrmTdBjC5l+lDbY0/6b07toiWNUtdKwN8RGTALvXmep
mUPzp7EuKYBIixb11cE96Tw1ZeesR74T19JmkKpzVKaQ71Gpj9qkyIeUZ9EIDaTf
BKt0y5R8klYzceKBcKzhq98ZSSAFbQhgCiLD1gWPSPrlB8+Xn79Uv3Ezn+ybM6ma
pM0AS8OI40j1lhJH2uZ6PsJ10Za1ynnGUbQUHWBgijF9hd3kylI7GpKaXBSwNphh
6dNIFeg2TLjdhK7ph0S/Fl4GQpfmAXykbKxdlYZd3BD4M4GH/QeK0gpQno6vLRuY
8s0JgEmvwbgsb7k98SZo/THENxWhhPmJSwKHsnDbUBe7hTs125hS9q3GV6L3q15G
qdZORZexC2imx2Bd4zC3vssnSAkrTjsSEQUuJa8TzfZwZQJjjH3cekIC18WU1Xj9
JnCEGtDyiDb9oc0paiH/fOn8Ub07aMMC7pht++FGAPfKBfEZ6DCv8xVCBIhjZTMp
f0gfagR2IBv7A0sAhyievU/ZKN41WMK4z9MB1W7WAqrqd1ZAc6mrDkhhHWWHxBVD
FXZ25ZdMhrsie4Tp2oeXhyOXVGyYQt/gVsC75PCPPPCxTxIO2iiiSmFfI62SNt7i
xVdLjmd30uMwyuaV16800pqPHYtfFX8LhaGqtBdqyx1GTvPoiMi/HmOjSFwSOlEC
tZbNEYm5xZX0ixjk7prhI+Nn4rutN1ugSUDD80t3f1OW0DOpqMSacIC5Nntfgmql
nvbOI5CqMk0VBsq91rBIeIaJkZDJ24mEaFIBXn8DseewJGPPGlNf2o3oron3jKrn
HVhGaCDMzTrdqjroIPf6RtKXDvmKyYNVDBhtdTSi8iBDX5DbWpsxENjG+0EIo2Gc
btw7vI5LynLvaXhkPRx2SntHH9jQpR9namdQ8Q06y8/3dydvMicWi+B4KVGUGZCS
XTedk5xYajns9PaDyGFWSL+eX3kAIxV9vNTsRMkPrp0XDHp3XTB8PGuM1njVJg+w
Y61NTSlYj2eD07hLuvkhzJUkhjFwf5BtfpSSuXYxpnIjwKwO1NcKMAXbD1WkBEK4
8rZt+nRrraz02EjhkGVv7qo8+hddakLOvO1M4KqobcTuzKLcYX+AR8KJo9sWLuzP
GR7a1aZ6ri9TCCtDA5BgOjMNodGl2d8+wvznek9sUhBs8JXonJ1QzImigJ/8GHib
sQfr5JGZK/8BxYys5VuCqUMvbsA2ZkA1NkOAIlqk0rgoJ7spxrkxKL5P5cyI04ma
L4Sl0PXhj4H0lAsly8t9Dcza8tN8ECugr9jeUQUItSkkV3wuYndHvXAvRhlR74Wb
K+rsUTCmJD4XhDZKNLxi2MwAD6wtyqS3ntILJv+8ypFCooavT6btDKEFkISXDS6D
Ke0j/ZKwIuIvbjK57OE36g48rAtZ3brb2xV33xJqlsuQ6gQz+ujzoAb9+honoKNo
/VeHepZVfeS68iMJtlIURru7an9D0jJKMSr29WF/kSGgFMRa1gaSNDDTipkAIjj3
IuJcClNrImPJhN1+/9lZtp4RQMA8O5eWu1+Ys03Dx6Q28yKfoSTX/SIfu07axlI/
jc2M0HtiB/VVXIkIC3pksBOfNPs1r+BQMEo9Ih8Wu1cMI8SiL99g1rG573WYIMdF
3LnGfLLjPFytjpUn8UqF6acOWkEyJSUOVezj/HNw0TvSkcG3hk5cFahz1TEa8ssV
g0AQ0pr3BtsQJUZvlir2V6VSgInlpXNJa5Y8HPviT2rLXYuSN7PUnOrm7wmjq36L
O7bnWjquXfTO3HIBucPF4oEo4U+duhffOEDtffwtuAl8s7GtlOzbzNqbFvyKZQVh
soef5Hm0G+PvJTafR9mhoJcNlpmcW03WqvIrlta2pFD+k249mizYNONx+IEbyMqe
dspd5LJUMrceWNiNins5oxWLj2j1Kzsrk0UwWssfSYl5ysP4P6Qhpc65OM1f12FC
pEOYBrAWM/hYW9O3EXMNq/7PQr6f8my8ybWfmFkeWexM1Jb2Z11ElqX/+m3R2wIM
wNGOx0xlDefgwyFtyBkGG8q6yEn/Gmx5UXQ2/aKgRB6mMqDCv/T9rb2Hxkdjx+F6
4FyklAdLtvn3+ZntAYA6smcSfGYXey5YBV9EIHh3Vqeitr1f8H6ttaCFYfX0EcKC
t1ABa8AGY5Ssihb2sNTJVwoVzhlZEAmvzTDpx1VTkf13Eg83tX8qp8YmPhiSPQEL
zXL64GeQvVzgtyRIYWB9i9zFoHmSFtcPpP01Hbhco54HvbK4TekJJoWV59WG4tG/
cVI6+zcj78ht1jthd0hNuX879nSnuafuBVd/JpQj9xnyy0OzDnRukhVhuCZa4qCv
JsdngTXQHk0DsaSwmiFoCTKdMDb90gM+wTNjm/bCS89XDoOB30iako6imydOumM6
ZTX7bus1JSFMudYnZ0gxtTmtLj/2vygPj1Q22d1vW3dsfkmQ0RbLJZgTODvvv3Lb
Q4q5BoadxpNH5FUV65PtIwQ+kckITiVs2AYhQWN3sLfbXQ2M1gJ2WXryWGp69a8h
c4biO1bABiL4NIRWjQcHCylbpKzV4yJLZ1Rxq16bHOvtd+S1hlz3JJWv6brG/4tu
/VUeaABTi7XB+Gzz/11bvRf3UTvjc5Yrvb+DMf4AmNJqRnlEy8Bu75UjE/4+rMEE
qNolc6cm9PTBJDndEM45DxSPMGvUQMg7lqnJag+76XzoTE4CqvSs4/HPwJpD1RWW
rvT6z4KtLoPOinhxHH+f1xHNUwm24umXkeSE8+uXJeqrMWfOnA3+CePghWKeIfjL
5P/KlPsgcTit85zwMT717O01ef5zNOSYLyw3H9HQ/v/TH7wvdOpoT+xQEo4FucR2
pLbkbq8FkBpPnypY8FgVZGvv5xDBrcDV0zozc3wtekOFw6LDLoWmBKAup7In8kq7
YLSFdjF71W1SEkkoe29F1hTt6DpsUrLkQNqlpmtnxWcIZ4fw33YGFcaVUu8IB80a
9Qj9EDuY0fCoBqbA0fM1owM7kDfbvHKzfZpv9LTd+EcigvY0bssUCPcR03748JE3
RFWdxMPPmTwjQ5z+k40Ce+QlDjrv1aolORVTKpgM5x01xWuy3DtpZ+5yzIfgrDJJ
k/JNnTt0JmhdFkIvNjFdk4v33limYDmnhSG9xGYjrhvvHEbjhbliMmCKNFMeglrM
8F5a0HDtdkUD0E7Alvazs0Jfcy5q03nDFHSlsnv2lB86ljQLQvYlNtrYbWGW35nT
2Jxk7h/ORc2G3G9js/pe1r2ma/sFbPal58aYtwOymR0fy2b0zBcg6Pk/GTSdEhW/
FViHyypR2jjWYqnfz9uGDy9voA+rs9TMF9alpzrbkOJLWB/jboNN3Yh4FxG5Uj4R
G/Ar89QkUkKibNZvjMhawHZ2OD4HPqDeIq7TTv0CNftPba7xqCzy8QMAb/SDc2NU
CK25QNzWzvPV1OqMfh15lEpCv5iLEFXww/A1DdIjFCfcztJLdcOmh5OYEeScQCQ8
nUom10iIRhtsIRmkKZa5p1m2soSKRMofmS93shbXtRPGJbj1apweEL+9IbKaN/Z+
PJBDoMA6AhHazKUM/J1SKbazrmu5zLAK8ARGJ0ETgyengEBKJadXbZlB69RJorMQ
+Zn4YjC33af6ABygRvGdUtF9JYg6trd3Hsb59ydUCfxpNLTlb+x6DitDQG6cGYMU
dZWk2FAzEe7XF4mmuT26QIBTUNPlhQlvGaQZ+6aywuk+vUW01I1T8eJ5vGbvdpQY
XaLRvd84YU8xkCGuMl4QYOJF6UYayCSWLyyV7NvXWsLTlcD8Vtw6kUkWDrrFDi0s
4h+J2N2nOo19JFApSyMGhoMbYh9F99RBAfDd+e4fOk10SYnDSR45ZmbVP6KmL6yO
V/jpxr7nQCXB5Lpne2AW+mDAqd+yOfbfLR8sN3emnmrUbSnhgM/0fb0vasFScqmh
7h7mosCh8wBB65bT8cI04QzT4yCptJXLhwfXQ+KtmcoU6B6KQLuISWZR2pSqzdTb
NEbOkTaYwEqr/XjAHS52J3QUZVbK7BIMtpml7t8LRWGGS0fFrTmqkqhMApF19Bdj
1Gr43QO6xyz0Jyw1KuE3LeyKBw7AtfZp9xfnpGObvY4Bk2h3cyHvCuIp4YlSsbm7
7Ezv7s+PbyOB8gKTFRN2z9UwMGBLj8y4lPf621S7nyVQLRxQ8hgtECIYgwYh20zf
gQUO2HYE8qmcpU8C0vNzEyCZQlw4UyaVQBObDtff+hAeHQVq9whlmcbVvMxnb+6U
SQZocZyIGauQVbYIeD4wEUAoOhLokqYX9pXh8TjZrynFv/wKfCmf5AWhTm0Jgm5G
Kex3+Wc/A7dhryFyhvBdBwB9m8riUiXD7SBmUfawRcXpVzpLGl7tJwIzm/J3bsHI
5d6njPy/P2H8G3OMUvsLU89MpKNN1Hbr7SMqEVweYuTFQ9cViEpzILdpqpbO8bSH
WD4hoGCgcXDMIxlM7f1JzGkzEXGrZDIl0zc1u8t6oS7pRl741c1ZMfYKGXQkqM/Y
3rvTuOQxJN2aKMwal4hhfinydEKC0aaSarVkefx6JD2eN/kgV/duY9pUnAcSF1FX
paxa62V8I4p9NIxSfw31utoeEJklgIxoM3SPDRk6RKzVoEZmWhEk3v+W2nHR9HtW
rqOisis4RiLlmKHtj+DJ6wHcvAK0xDhlqxEsTqelTUGKxk+cNxdLw/J01kRdKB1O
dg3RyLvHdTlVj/m1VE7csOpbjyXnwonb93WG2RE0ljPcQXHZdWjC1Fa5qoplBQbk
gkJ3xITr8MpQW/ZwiPs9RCfhA5T2SJMPlUxKwC51t/87k0/B1qIs93yGteI+OTbh
lrCAyi+jztW0gXpHkjxqCCjJ/d0XxQWT/E9O2vCFgBUGQwpu1laWz8hmn4Z2ejwk
fL6ESw6fEx1y1nJ/Ytm4TY+4+JcvLD/YoXio4vlzduakvH7YOlgtlK6vl4dNAMPK
bAa4CF9PffIIjwk262MiaXN6w9mG1HSnq1Jz94mS+kXIviHG9tcR5x2RxyueJjD6
0mvFo2fzABs/mUXzGPTYGmlHlWt3QJ+/thRX854sFxwbmlrbds5crD9VFXzeMNxW
F9/teCb8Lv29GtLQYsA9iKWLz677DZ33cQzQ76o+OZmGPgHOsbIzlonj+MIx8ikT
jeHRttSX4AFmsNUg08pN+TAJLDSSZWECC/HIdRC60mCybdD0OISvumM8bFPUDZFA
U4/qn/b9stWG08sWh9o01HvIrshPR53smUBNNajbaiMvhgjJewl9N71nvKIZLskk
YewiVjo7neod65dJkvJZuTB6zmdHogP+J0IhYlLA2nuulzLD8jPJ3lqFjTnD6OzK
dMstVYte95AMp1K3DYvxlSHzHNMWt48M/rm2v5o6q/2rLfYLcnLtj1tn9JCniIhS
XXclYmnxVVVr6nX+HH8p1TUlhnw8J+UdCiYPsN5gI9ZDvCqaMds3+pO/tT5as5/J
aJPd/6d5VPwGZfTQ4ynlYhxhPwJqKxwdE2Ce/yB6CW51Bq49q8e/PE1ozc23m/Th
z/yHsFlM39F6RXkAQY0K2LupUJwWp/AkGhxG/j4Z7YWT/WW+hvOLx8DxRErwoibQ
qmh++u7//vwmZW1rfvZAHLez6K2Qtl2X3VUW08Ae8XRfvwTiTZX4rMwbcbUIxJRR
+KosXTsWnkJ5NlaJ3TuKFCF8FiOo7sIVoruiOdhzA1L33Jx/L1Jf9VICyciQieAo
YlJLRGf2dj4+5Uwrg2LiYOEpflToWpSJb2lmc/Piz5sJgW25xCkASgVLFn2HGeBG
mLQukgOBnBzCG2RXlTMDY8ZAzUtGZ4ctH2Xp5HymF+syGzTWszWou9Qqr/UBMIxH
NjQztFNigxcL1mshQNhvbIFQJR3Oa6goL36fyCtnz1eSv4oqu7ykUAgLHa5XwgvY
RZWgu6SARPxnHyrWC/BXqJngigkHd57jku6TsjIGFy3nde9/6rmk3ticMoG/LR+o
qOZ83o/kCcdkNpz0VIFrqMmYqxRjqzjhbo2Vy4rPGNl/1MqmZLk4R43Oyw191g9S
QLuZA892g2xPbNEY1v83CYhfdp3s9PTUlALO8NeE+ghvorEpqufCZDzLSg1/8RMK
Jf5TglJXHDQ+6eCRTH5xFUBS7M3bo2gtLXX1BQLGk0rPdov8PJj97dTzuC6CpuNZ
y99BcCJ6VZoOtC1eGr4uy3QNS7S87pzxdsgMwqsR0448AuoSpMQbvUuJjdE9YSq2
B6D4V2qT2/Ws6hh4I8+9uuMr8teY0Fra2u0tLoWdPWGoVxd5KA02gPVEtASM5fXo
jzRR2odx4ldEm04F3CFD8YuNmxLcUm3qCJbSWgBd6ehEzjqiW/u927f+J43r5LWx
wEd/kecvRp29X5nRpHx4MkS/NRR6l92AUuAkCTP0QzAriDGxuE0DWPYwuFhY4bqq
iGlNqySybOIBYJG4rC8WASG+gAx4D17Km6+Z2PpKicHP4yU7IX2+EhGjRndKfpgw
/GUO4cmgw6OpBHPziknuxLc/9Ve7qWcGbnASaJw5TBl1a+wLZn9i2COgMe/KmIJ5
mSt4ZT/vd3j0U42FZ796pe31FN4ZMeq4bR+cyS+FLkxRZu7d+ID+IZT14rOvr/Av
yqi0FIVEahr1l2gbo84H5k+1hx+bZhIjmRgjqVdlriYR5sjmvsjMSacGw2BWYmn8
owNPS1qlGgEhF5o59xWPuLpTZ26EVnLRPHzQH1JbIPIl2mLmKwMrk06ndakQ3NXk
n4RK+mgY/heQ+6FRSpaITL2id97y4Zeb0M+uxoyNf8PcmFFpc6jCUzOoYlc6vKH7
kWQjv1jhEFyhEfqJON6lmORsGi3AYj7W/f6gtKMQYQ4dUXzph2t8lCT/Ugu7Sp5Z
BrhCQAvWZNbrjM3QFBu7aHuXvdcqbTtJBPqm3YtcwhOH+0fPaW1ARtLNko5Q1Uvf
s7Q2UaPt61pRYD4E6OsYUAF/dqIcptI1YuYYT8LZD/APs49l6ao63qG4j+be8VcC
S/QjPTeevY0I5RENjoauDy3GYnIc0rmEHMAgzEj3HD+1xeWFVpsqL7EpQUS6pUZb
5xFkYkzzkGs10tch5XU/NOrW1vPQdYvTUYQ1//YHQUp9I/KXsg1dAh1KDITzcjGO
3yoMqJw/Gsr9yvxJs8k6rfMMjBcX1okarE4z5jhYH5rPUuDDpbQnBj0jk/bYs1gU
CWl2jXZLglxhkRQ0yNf8+YSEv+CZToCb8wnAecQP7J0EgfbVBnNdZee3ppSUdGTe
G3zJY5UzAWecFfhnaXx3iPosHmwqt+wUMnzUQZGwWiJ8Ga3d+qrBhUc4gQZyJOsg
bPt++useivm4nudGNab0cBqcqU/eu6LhGPdEXpnPIlM=
`protect END_PROTECTED
