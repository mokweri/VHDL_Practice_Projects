`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t07Jwtpnwwj97dr/ADDG+lvCRJ8Tcj5eXTA1+jI5zVkwafB6P/s2RNpm0IXui2qc
hZv93vPmA3Gd/LbFMM4u4OtvN0DcmYaN6ccJp2aQiAZmuSJeI53PE0XxbfBSeMev
vUKrfZbndVRKNax6oHLFdWgx2bwap8TAYbykCUVvE0tzhiH58quYZy3YfMQNQVn9
cr13IPjS3J1EpL0yu8uHQIM/UC1yICjJSkFd58ROxcoQwnPZlbZvfmS9KCoW+tKM
UaU+AiR61gn+VEMgQaI7xTJ6OGNW6eYRl9EBXff1fKY70V8X3HZDlszsKVxx8SHM
0WBRR/lDrKgp2dw4D25LhOD1fVnjun37R045gHBZa+PeYPewzGwJkdGnuC+MysFm
lqC30sYFXsc1+ZeGBn/b11B2lNJZnX7JL6DnLaJZyKc+5RGhWbxBdy6Nhk36jjVM
RYIff4u4wEuZbW+CsfyaiTZuxNXocio0HCUK7khK3baHPFvRcXx1IgAhISMHxYRj
GFM2ObR17xzvVrZ/3anReQ==
`protect END_PROTECTED
