`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DiXrzSdprbCN55MHqhRTI2aB9d/8+lYrRohflQG3lz0B8EJ7535SLxlB2Cdt6SS8
YLEvV6o+gfyRUBYtW2l5+3yg26kvTt4DWaFeeR8CeZ4m0fTP//cHewBQh5Q/pdAb
nXEBHqQIhPL/cItAAOKuSoJSM1wtaS0mRNN24CPCSSfnGm0dYQB3h3Four7NPMD3
8pMJ1CXGeWfaCKl5N9mP7e7YOLHd6x6/8Tocd++YyoSCq+I5cZxvGZUkCvaXHvGc
IBD0WwrPh7z3OpEIeg13p79go6OkCY9e/sVX181S3ABVg/if9tZIEwnbIbds8aDr
/Xy6NWstfZxpJIG/ADyLvUMqbXWQ6LeTDKLVFLC4vWB4d9aJbudptVTb45ASFou4
63unwFL/U7AKk+0fgu2vw9orBP5w7lusSoumVIhzE+BHMomEwJhrtxh+w23Z9nvt
nduhRgZXqIFRdIWoyALsCmP+gvr8v06DyLPc80lEGAcXsBiFZBlx+XV8MG1T+ANb
2feUJV3IAAkE59budzZhsMtNJa1EV75c7tYZI/DE+T96ywGQzlxNN2O7kGocLc4u
niaJf80Za6DN1CuGXlnsFVUDt/E6leWgPYklvjI+OqGwiL3OGtUqgXuhXfF41byJ
PIAi7qJhhdik2fcQIyrvj3iPI6/RKrFU9PG9NGoWbxCOBgAllLPXYH416VKhfdwd
STZMr6BcmpZoI3dSIHlLTto/4yZwJUhLxiUFPP3znSTCbTNtjIlhhlNTW6kvrPq1
lYQFKkGYwv9akgzhT/fBcK+g1Cvd8yjHjUb6omrs1tPVIpS2uWmniMnmtpP8VfrX
ASmOtMEvCveAHBv3wPeByAmlYWDAYRuXVN6ZHILHJ4WHBUAPDhHu+cEgUYZnAW3k
UliksPpGQQ1K6iOR04JPIC72wsnxH7hSNEtoTxdmj5Qy50VDvHFAyarrX94gaNyS
AZDcl9G29N0mOC60lWUqxOlrQ5Phy/1SYu4lDrc/J9DKWFFqYmKTdUsf464L6EVI
vmYlhnsACQsMIzv3guY38nJR1T8RyQQvp1eZsWLd1gvzqD9Ayy3Sk0BVeoO/o4jJ
715u/SulONw1Q4ahXZlzCKYCAyCjqF0HOvn5+j2Oy6mFtXxESuaYjQx3UY4KSkHK
9FM4W6RGLoWpGsMC40Dzmz8vIwxUKRR3y0tU+4ztabtAy5rPTYFog1o/zQDZAjnV
suMgBZACnAvOij2RcIwHfXiq+HWYCOkc4XeyaA7TQrreREPKphH6rBtdotSDRk9v
eKbPBWn9V1PTglJu8hhN7cdsulZmvCYlLH9WlwM8UrYnvmTKoEuGo9gv2oWb1ORS
zrONNuhi96z4SjBolv9YAn588wgDF7X59aAQ6ZfsXQvCdJHTE6vmEDjsvwAbHLBq
6cRu7oa2dWRW+A5SvkfE+gk+g2c5hXWiFHjR/XnmWKh6QM+4FmmFW+4EGg4xxlOx
9k/8h0+XlcT3KvX0JLm2xyV9jibdvP1wHDP2shrEYcOfgPfoCvEexLSCGk7XkRUS
VY5Zah436H5XGHEDjBzVBegPMzZgPUMRptRVfPTmNalR/bdPOYqLPfpRuLZMAbYm
miVUThFA2rmZ5985SSQF7nmg/Voy2jlj7nY0aOLHYxpnx7GEPsAIdsEuIbnt/yYx
3NkaxP++XXcWiRxlxRvF52I1nc/pA2xsOEuqocJSwDTOhUAyfOX3l/EfiPYWXQO9
0IAJDR/tsGIBerhov/irrOSCG1SRNJYuR0eY8BQDZy0CKyZfB5GO/F1ZrB80FTUC
+c2+oT1TjnxUWapKcdiP9F03kt6LUuzMKkF8SxH9HX8xpc6xwPAeyOepxiHmPk6x
m0ZljGNKHFXAF9/8wGOYT6dGw7kB80bJl1r9bJYbS0ZwiTkZYb6QluyLA+0Dvzr2
7YXg8ije8aWFukZy7AJo6bb3vT4RRUOktQSuKTmCNDLpQstmt6WrIUPvJu7x8GBk
V1Cen6xcsnwmv1mIuK3DAytbFYH6b56gmbPMwvMPnLGM5Uj8XlC4exxItQfX1BVt
TSz8Ci8bQs7BbxGbD/1KcN9QgSgxJthPDtQnItjLvdohDJmfwvNHL5+ndbZJvhzK
5QFvgzib1m5ce34Q9Fa73YDD+bTuvLMeIOncm6eP6Xh24ieGQN0SoVU1crXp1/Gr
F49tC3GYAA3Hq9MtklJSWqHgYhJLc3pgb9y/wm5YjkIxVaoUf11CxcHOi4fAnVi7
uEPbJxQsu3s7Sf2O1ET5FTXP+BllBABWCPpE6QpuW82WatMw2xn31wc1o+xBD7wo
21g/hJC9wQICS5RnbRLzN/VNFNC1eNdrWDgPZPsYbXyzql7gio/bJEiQMrtaIDVX
LbLT0faIkGNiJ2GxpuMUUGDfH99w5NP7E7cAGFTLWbDcnzHAEmzB/VhOfynvwOTf
sljvasKw+RXCUDZ7ZmxJEJw8yuIk6N4XMHFKDreYl2dIC2xmRhRW3PIn5nbl2BNl
iddl/ZfUC0jAssLTYox2ZO/+6ASrz7ApRm3yC+wlFi8KcuGhwYaMImNyggxd0MK/
S0UjpOAN00SJykP2gMS7D2I1UjiXK3Zkht3fHjZCnGH/yFILvbDke71E6+x07fqL
/Nx/8N+nY0a3mROurDsjDa+rlP3Djqlb1wozRnJjxx3zXY5QQZaHCqBCQIGkr8Ha
MKEUjH12rRAmmXG0aq2ohgycre3Ye020qT0kIuISOB1NdYIKzA+i/+qu+Lyj86Di
jWgaKQ/lfcoOPXYK55TNfvpgo1h+AdbRisiV3ukokhpfSU3gPZbYMjxqQ4o601r8
G343DPE+0dKf/rvU6Xq06xyMtX4a0230cDsSejSZrWs=
`protect END_PROTECTED
