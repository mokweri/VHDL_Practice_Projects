`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9MvZCwwR4oEDPyLeKputf3UHkSsEPXcoFP6/OxCSNFM/76NDTfxkYvfRVJtFcd3
V7lKsBcfqWHQzv3eu2Och4u8zK47427VPWfBLVZkETP2jm6YlJKrV1omyp9sLkhX
Vfcy9wX8X2Xh33hKhNkL8+z5TN4UA4y/djeVxEycRHe+fEBY/SPJSjGfBLJaxT1a
v8LMUWGwoF9jSBfRbgpJeERMoa8fFOfyyvflcLCKYTs+VK2TfdG+zHkH/7JOAP5S
1LGKVX/NjEdGXn6DrldUyyrvtXqa3hXXColV06/HarHXBRsvMJ0Vp2dHGUfikaEo
15qOsg4EuJ8GLDmAH8xrap9S+QavD2L3etyND3ePA3+HpY1DLekbDlky+wBKb1R5
uf5rnxXM0g6rcCYNZPLcXCy9YAq6L20y6Uj1XZs6lDaIZ62YLhw6EzNCzMDdgR8k
vG7IlxrIJXyFRqbYeClpgVdxghENTAGD2+U/xFvbcujjC8uharakRC+LUougkjii
jcU6acafHQcNwNr/CP5IgIWupHmbXINc/j/Id48Fb/nz7J009jAED43F7jT/La4E
j4KJAb6bfjP2plfKgUCE9KIXBC+WvEgEyT9B0DZdiJixYi5bVJnTYwZNAZE+Vx5P
WKxEjJCBKSi3dQWEpFWMEGrFJyDzFie7y6JcTjgbmC1MtVvCxrs9kfDEmyEcMHOR
5kreQArvdGum67ZUeVeZOULr7RT3/QZ9BLq+Y0WN/PwKJEo2YFY65dvGwPOfIbRS
Egfuy2TfaZwKwfQfVIu8pfEbIwI9k/2mC68mXi5lEkcWex3VQDxexbZy1Z8Ah+AR
l6NOZBZffT1lxHVC0/p2cphXako+q+hZvPtFbU68iuNWoGLd7g1fRkbvxlUXjFWc
6B3ZQaio0Xl5QrnLu3pjL0IT52KPrFfGv9RC+x+dH0ajij+gehTU+S8GDVxe4eSo
5sGVIJN4UAMcryJEuGdlBszN7Tx/0lZTiJrGJirKhfBkMqOTTAgT7xd4/nePXHll
JkosrjYfxFsfp0jv0cHfoui8eHg9srNMaptMCpCFe0pbftwvPSm2qwq8MMdX8ml+
SMGZcnZFUOgf8b/mdmFABxGBzpSUBdFaItu5fh+1GnqrLsmyFJ4m/6t/U5HWO9o6
8vT+9+aHvxWMHK1qpXs+bYJfAyE0e9m328ScNCfkU4p8COCR/Sb2kMeuYzEgyhV/
elckNBSN77hDdL5+CV3NiRJEOpgd5KNglacR6diFVELX+hEmGML2jjweZiUFf0A5
5R5Zbpfo4zKcNZx3fwooIvqB8ulKyT8HNOhrLxTMLWDNwKIWl33hAyjLjeaZAhas
Ak6D1DSfGWjnfad5XPzHbqRvusTW7LYj0rx9mxrzMzhh1mFPtX2ycvDW8wxH5ibK
yX61VRAbkJ9sC0cco5ywc7terUIg0cNHhv+ok9brbrmU0nOjxR33CQpA2QeK45Pw
SHDA9EUfVFm3s4QZ06cPaKnS0UjESK3Jo09x5hNM0KYnmvw0NMc9KKwH3BdUsHrs
D47XSNFYt7lHtb/aqBDHVPpolJrxHhK8PbtDREqNdsToFdEQpH9u7PRSi9W3klOC
1Pe/yBqmCmI3/mkEJMPQDK87a1GT3yTykJmORAGpNJBJlvnhqNY/E8STo9i/5v82
3pdqGbsbypCrvJIicUOuYkr23iySXK/GAMa15fZLHdlUYnP8z786TsqUibM/sU+t
Q9vwuizzxvHQg+hS+uqUB0ePHBMKxvmYj2Dz5JqYtk6cBOyx6i4NRFVkY0AxSKlO
aYd9RcF66zPsq8MMNfIch4nrb20fx69Ki0sWqq/8PDXsmshDRYt2mPzXrDfDkbQE
rECbahxRVk7pBykgiVWq5NIel5+T7gIhBLdA7WIp4CtcwAjwnaAYBPzSx/1U3jAx
WOSKDmkqJZleIPC0r7cX9lwcgnQE2A7bXw7mbeWQ82v3hVQbTWXowpWf/kQLFUL9
hcMZEQgiCUWTRDoV7vvxhH/TTznliWc1yX/mZh1tTk8BHiKFcaV7MfGUr7AZWtX4
rBSe6NNJFMu4yEg3C6f7qflOwE3O4FCwTDexVw+EbeV0ewiX/f3UdWou91EwYWyK
vjRAgCAzydey0+aw+wU/mLsBoz6XtZo7EoK8qM3yzOOTcrKiugYcTdncjlWVmER+
1cpwPZOxRjKzZ84BwOI1SUgh2nwishueyJzvirAzwk32PunNDXk2BeICmqPghlER
l0uvwKStC7CX+CaO4xY6OZB0fRATem4twz3+8ZgfXCNS+d7rzpoOmRKrKDlxDjFK
xOaqt3+7CHuBDReAGyKwDgI8XKyM0tI0F7W5p/EpkhsmNWWlTjUjpEIAvlR+xCpB
R/tnsKrH54uxfXd4dtF1LFxzY3r+L3fA10YTctx+QaRmh7DL5+h6YXgTt6U87Ry0
cfB5RE9jGtZhPo300KkoZQgjrijc3D3hmjGryuG17kueXyNqZdfpTbaxpx+w823J
o7Q95L/I4SGWE0EzD9R8XSn1Qxd1akK8CgP4CCC/Ge7xTpagRj2yzaWb0SMnmFGP
M69mJ2o65pPVPSVdccrbTEsMvcZpBz2ag771S8CPZ3ABMllM65w+cVv21+MKY/jB
tp81GwfR8bGYXTN9QovbTX6QSuvChHhx1wykplUnTyY88/1H8/ZofB+th9h4YvXa
3A/P9+v3Lg6xTIO0S/NfajJAzkKP3RKZNK1mU77cxw6IgHyg3IraMHWOG7zrW2L3
8PpTaWIE8OXVCWegRsbqMerJeI+gVINeLQ4XhN0Kv7LWtTF1ACdWkPIS77wv3/tx
+CO1dZ1qkmOFHBJx+nenxUiXQPUvD0/PDidMiQPBGr+Tx7FE2DK+YgpQbefbvokD
PK4fbsmaFRdmgoJoyzJ2nin72819idjmozTV9Xg5hODyRQZarx+DIUygasDyoslh
jV7JPlWzmr11cWPAmZna4rQjGlTK4VH7IhewqkCmLrlFV61StvHNYmvOmyNpKf0g
b8DWBG6+6zC80Mf6fbvJb/ssannORbNZ9PZpIpK7rVhsPXd2EOO1qyw5y6z0Uctc
nGrCe8ebibHKqlpt7mcTdH6niJ6AV822FHoQnScvtf9JeWPvntG1JTQQvGnvf5BE
4PltNUr4XKTEg8orFciheFVg8plsJAdDNTfWd+EVf6KLevLJ6Gyjp9UqfS1UiFSC
EG9CAL0r9/+LNfR2UvGyPS4qmd/CzkSCpRS1wBEg0v2CkWcTp8HyMUsUUqSsfqP1
DA+nAZ9+Z1QceA9MiQaO5v0PgUaoaoLhhDTKe7e7q2hDTm1Qlp0BFpsCVIITr9m3
KMt2n4iygnlTztnCdr9b6CdRD8/J9QlVBj13dqBvZPrZbqNYKP9wySK817KjUohD
ttBuEeg/s3AViGySQ3L8xzTW2yZtfKUxnxY8jDWDxNEBcjMa3C+GJi4qpFAucyEQ
senS+DeiPeOCr9a1FZ7digrsG7JMVdydo4ZM4Drx6GEnDT6LG3cuKWFqM7kw5ZLv
8ykgsxqqaAaeeW9eti85Uo8XJhf2u6kZkqJhuf4N0ojVa98VoUzpFBeYdy7BHtpR
dxOSExzbWHLUka4ok+mnKBPC7cepCCryd2RXfyu7RM3zh/N3WrIoIALu/3WOgX/1
Mr7p622/clyjbQJPXyrOeFn2liW1yqHMo/hYsIr37GqkGWSFReFXYRD0/7C8jHIl
KFnelq0IOeOIHyxzP1RvAFY4c7StWgwHsmMSH19xYFFAmvvAcu0QlgrURoTY3Iv9
fviwLPfjkB9LlySJIvln/V31gntCgi8LwxwKUqOfIGradcJMyS7vzItPQOU/xZJE
VKE4aP7C/IoaCGtHYvMcMD/eP0E3MxF9lz84WbusIJHwmHwxfz73g2qu8UEA3gXy
enNMy6budtwxQK1dw+V5psUODrO/9rYjCNLstWgm/rAWSGY9G/CiRP4PJ/OSG9N9
ANMd9n23Srv4vBKTJwb1EyMmoJHz9kYCeGCgHYTAcyYRITJUXwS76v5Rfjl4hJTL
ULI0trHF0pxmtMG5+rPfxFxhv4o250pfBSb1Ao5E6fblaoAZZ9MXWxKx/P3ii5/0
oi1Ns0P5etJjmudCNrhY8Pn3bUs5MharDu0DDbztr1RPYaJkxdrO0qmHQoHRFdeJ
/yKS+SRlH+Cu1FfVsMA282kRLgv/oULsQ6JTLTVf8e3fBKM3MC0PJrsNK8oByqkL
YJ0/Rs22T5CApisJS1iTS3iOuZevb/I26p7hOiA7SimrA1QRl6av8gix/ZXRE+pa
Rr23+RJtDh1rKocHSBMq/6S22jdP/Vt8jJU/HYqvOi8yrj896YowPbLt8YHW7jUz
CKSBdW0K3KwemPkk4LYT0Md31a91A69hm7YOq5hJZF/UpXKdZTLZxdAhleVOgcJy
GwGzUl1a7YcEHEWGZqU+mPi5N1HF7WNhDxjpeAz9GuDllKyTGn3k1aTIJZtibph8
+XAA0njNTVDx5HVSAwdwuVEqDa62Pq2I2Ka8gi8RoQcUc0ZiluqhO4Oz1tMudsh3
uy7azr/Uu/3ae1XN4AZgZbRtiE4nV4pKTd4DnrEesf+jy1GT2KWVqRD1oYPQnx7W
c3rxYtc1VPUQMZ0ontlp4BbE5dQVJNOvjlfcStNTgK7Ge6O/q2hIYkShbGb9cJQu
Z0eJemHxfC4snqbvDIOR/54c+NR/3DsWnB0v+I/kA5oj50joLgb5MQSBA5T2a7zN
rK6mh34ulTt77XB45EZhp8+U72m7kGZlFu5V95QynKltYS7FXw1yv+ybq2Fk5Jbd
Xa0gPGKuTFF+RL5g0nz17GFxJjfQDQhkYR8f+Hqm7pEO9ZZYFoHbNA878GkWjwyh
4N6sN/UKDSJ2RFnFx2FvevNRLuCJ6XuZYB9bzZRWPZtV5JnNM0u9nzD/vkb2RQno
r2D7Ypt9DkHRofYBiy3YNFLNVj7804n/BjH7pSlTmHGZ9zo5RRtzUFnfcZl1OVny
EoTEWRyVDgQPYycVpI+t0vlPty9s7MKYkOpc2bLaI3ODs5TG7AwCoOeBSdaPUCqR
Fz0tg83I4a5S11YoRvgzu8uKaA9H8nwJpfvKOmLRKIDN6KMYESTMP+c7vcE5+MgN
rTtxgk0huUrl4IcQSowhDU0n4N9iKTxwlvtF6tDpttmwTfEYDoLJ3patAh2rE7FL
8Xb2XqzDpFDp35kuqht+AHM+PMFFJNsUjg+M2t666hsUf8/9P0QR7tmEO8y0m103
5ksVxcUg80ik7zm641Jj8WH7c1PyNC4+B5dzLI7Hxui4xi+P92PL9049IUFmJGla
60QPwWehaBDyJYduIAU0h/cCf9gJ47olgnn6QSsBNPxEx42HjA4U92hGjWboqgHU
EM1+2X1dePsJAaW14EtwaRJCOHhsqK9TF9ZKe6eQSbAEq3RXwGq95M0v8xQiC0Dw
ba9UKRFtSzbfFWteQZbBqqFQKHc5nqA6QQpmBmJmRTu/Yq/zM6pGlzKrzcI8tSmK
yKET9MGfw7szbMDr3N9nAAICQjyKoaf41kyhlRZl9v9vYhJIgG+mBfPtnOCmdTv4
VplWXp4k1sD/4SCH8oeIjr0RmoHCuil8O6jk4kTgkp/P57LGh6GfIcfu6RPU5n0L
09xfwok83g5kn0Xi+MC9elz+VjFn06Dw9B6nMtlgnTwHV3Jc5xgfaESMIQFYuP8c
BMMfULUsaDOljhLX8zqKlnUDyqG/qjBgr+jPrtD+EHf3rVM2u/LHMd2gNCL558Tv
ii2y2IB+uTwXB6uWBbL+Q6oVTqfph/MxPBzSo3EGokeZBsXc8wE8vfB9gnMizPSS
1hm6lIe1w6SfGzmCKcVuazkUBRGvShaJFi/92Iuf7LAGUkZvf9vCaiLNf2E8Fe4v
SfpiawtJjCn848+o/1diRMfu1jxjRhxuqgdynDM3N301D2H+jIL002YTSgR3+Q73
sukn9fNSLn8JD79iA1lLUDSLTZXoOd1XNFmPWx1+MCS0Ip1+8vfx2JapDPpp56qD
CyxcuMiaCJ8wYdPFLBolFpV+Dsdehgm7rxqZL7JsVvCAm5dQYZxvtn4fyvLFS/pT
rxvEUxD0nFa7oXPsseEGdEkL/qpciirVpKgTv2XOhkw+DVrDe1BrgHuq2j9B7OOZ
DBFTnEQXXvs3+/lo/41ijDlPmeR6co1rQHucRSPp61hKjpRcEFMc4YD78r1obQgw
qNeEIncb7uON02PNORryDqU4gSUn74rLw5DnWfSyH8pU91Or/Awd4SXFFxt30Yam
b1ApGkgdrAOaOsucRLS5T31s1SDYWAqoSexE5Kljx9ZMKlP2WoWMgqWhhQfE98ty
u4LrHMipMtSKZOIgVStOiPoEt3Emo3GJSPGeDeS0SOJCovfFIi1XBww5GWmZt697
2ElvuqsBwZcgNkniMoNN5D3hKcf6wBmPYDF4RBTI5stbboVKssz3f5sk+mg5kO+8
pcJ66cQa3ykgEIY4JV7eRKQZOXyk0DWsYYd6E14rubstnho5of0lUmSL1tY9kJmJ
XbZAP0GR06XXl+6rePTk4mvG3YuAEIy4/ZqYneGphmzNWm/nLhrUdJn0DL+VGgL3
Wu4o6wRqv8XHfsbzpx2o6mZvkYbV2qDEEsNivjCb8Mk6WMmmKs2DES1OaF0xPJbZ
n1cYROjujsJDMgX3iZ5OtGSMd/f+X+tjO4sfMVfF1jv8UXHByWiawPL8GC4ssEA0
qi9yLdPujh5g6U4K3eAi/W4ATPpUC/2i++GT6Pf4bF5qlrBUZvWXJCyd4NBT64s2
397qgKkxI9vEKEN0E4Qgy3gy1nAGCOodFhwu2jbhOs0/LcHU52EnP+x1xjKKQBkj
+vJ+gk8f3sGWHQqhoRYa9AAwnHEwcnzCrmhiSLEDx11Ed2wnd88wLrxW1nduieqa
xdh0lbWaCu7AwDe31AwsxtUT8PKPTeqhFH2S5W0yaaKwVS8cTwwcEaKIE1K5gwTT
/Eiup3+OEUFv0KFR6ns5BaS34v4H87L4px8eXwlWbFhbzybeZ+bR7qX1hlQE34F4
QRPrDTDNaQbJWt1trNW1ePnEHxfbmZhot+zswU686cBfPKrncNEr6eMulmAx+bN/
qviIIuAxYH/sREn8mGFxpNaGmcq1kFn+02d71TwpNJiuGTMCGQQAgPLmngAQL+Lx
sYLV97mFyES0J83bHFA8CbpgIev6Rvz1wOdWM/3kwTwYRrYNpFjZT4b1en3c5FvJ
JC9+ScJNIDx6Obz6xpy2k+dsCDtrrRYk/6J8zVLXQASYRWB/EMcF5MtEi39Z27xt
/7N8FcrWG75K/RvqLTjUEWrnb1YaegbWFsWlkLjMlIuvy/fkgDG0WrJPTN0lz/X7
QY4NCJz7DTR31XS3bQyRadIpjkUvth54iQA0GVSlBTp8PsmumEBIjqbcQwF3FayP
bXlZ4k4smD8675vZ1lyctOuu4rOkr6zH2DdsHBPjqq88mmTL/6wVdBmwf4vq5U2Q
fGsTf/rxIc60lwvH+1xhsyKt3vRoWsurR5QDT/Gyj0+V46D1hoFbE78BduA7yv7W
W2JPynlTPjAD4rQ3XY26q6sDPGyHz5gptEV3IWKrBrHe6Q6vg1zM58HRzZcZXXKa
tDsmkTf+x4bVMYQtNK0Dl9SBigV8apcbKKbtqvHe5um4lPsTwTrRpB9NzNhXXNN0
pXAhab3wqSBoZGaiuHR5rqEqQUH/gglcH1uHmbD9kKnbO42RpTlHg/qrPTFLeJ2H
6QsLs+v3IqV0Nqw1PH/8yfgoNsn/XjvHvAlStUQhsW5mGK2SPQ6gpmn2pov3TZfU
ePXgxw3ePPF+ngr5Tm3mZ88RalILcZmC4kSQatMojQD4tBzvwxTS2TbHRdj8uRB2
NqAnqmgFQ0yvwC3kqoB+5x5r/ZlMM0H951jwRuZnn9r4nE04Mqo6a41fstvhFBoU
HnTps9QKFW+ZsJQwI7NmBqIF+yM0AG0g2cNf557rFzfZvt9ZyHbzH1zSN71X/PZh
B3Dd7QJJLxFvBiNTTK0+y6lyIyIzDZ/y0LjI/tOaFLkquoQy8gRVqlE4I9Mv/5NG
+AVexNZMnaXUFAGYLdlwjOHj8ntoVV11OWxS1Jb/3NWSJ/v4qahMvzy8KnzXgeci
4sdPGLjaj7keZ+oM8wqbCqzyt2lvSuMXrV0bO6NfA/YDXOPEI/M+/ZXMPENRmP8m
6vxzmJQaeARcuouQli84xt0DKACjp5AozmR7c/iqNLNHnsE+oUy7zqaNpmQUy8SF
xSxhJw9CJ7g9PdUo4CPNfL6KWJH13rSHCE06YzcKmxyfJYfAPqQiV+hSdcxezirC
b6gkLBsEbyJYce+1uXIqhYs14zcykGjILcFPibveSK/mxF50BxIdYI6Y1Bw3VS5z
4lT4ZdSkNpxtFItfM5HJr9GZD1ztIMrBVvutZcHotCoQkLJPrzI+cQT3oZj0NVh6
h/0cFLf9BeWSuhXsTcclHU+f2Xd0aPdK6P7RjzXSrS4BuVMFF85emviqO2Tu7AgD
OiqFA9SKjJ3QG1jLyvtA2neLayobQGwc/54xOugGftvHubXX2weAL319PtLA0+0T
RGTb1qJuPjf00BgjkSGS/NxfQq3r9LxzOX2JVVWf7aE1ULKSyp3x9WNUrwrLF/ZN
AHYoXdKgT6VHcJZHcR37QBetxNnBClgEi0SDiGUS1XKbpOpAYuOPWNGRPQ6YjiRg
/DwSLBFAKHnpAV7Iu1VF+F9DaTop9Qav1CEj70zxg2URs/r4I1loLyzymZYpfs1B
gc169jSfdeeAkJ4tvKomS862tVvI/X02tPX34avMn4rGaAOqpA0ewbxpNLQkZwoW
xZWHOt1RAmR8Ci6kwV+qdR+ix1lRV2r7Ootk6hOA/APQYvuZgfksGKEWOzzT00H8
mxR6H1ZzrvW6ju8ccKyMUIa+fbaCjkNXtNa0vGL8xBNatrv3lnW8k0y6wrxIyyad
A6c1kMCGOv8kYoqGIbKqTOECqrPVW7ybyrmqybXQTV62v/rCu1jKDnWDKqoNf5Wu
TE6X1+uVfJF8SqMp97XnhHy7hsgoa7Apzzq1j3vq+MKy5H2U5f0i6kPvTewAYTTB
MJtfEbR63YdUqqNrGxLN7RsdyJVzFHQQ27imEL03ey5CTxLpdqhKPL9oU96QbY46
rcwwmRtqiHzJKIw5xJFeGCY6bDir4IyHfBgO3bC+ncUbxyGAe96D0prs3Hfuy96B
VP9R9WLh6sEz98R6WRhLUXxmKQci5ew47fjgCNHhOF3phnU8rifCKnhSBev9mOKY
P0LvluYMFK7j3K+kfqr3gNL+jcbORhXNgf162RAM4LVZfG+NRF6J1DDu5Cl6TLsy
9TchR4y6r7Q/61NNnKEkKSwamGLvfIiz1NkEqgDI1D0SFrytVkopD3J8vAARLaDF
CR1tyhswL2xfgmhgIUpD0hQHZT5WwDw8ytnkbJkXBfU8m2PpB5WYyE53VOnXEbgM
pRZiRN8yz4v8eeGwayWsejPe0oVLgxI+E0V0DGCzLoYuJjug6PuVaE5RDfSXIpAw
JB9mZV2Q9HoTjXbpcKKLGHBEASSKqrKeU3cQzbami159vEasDAyAWHUVvRTVTj//
7Z1slG8nosu7LjkZYski9v6PbzIyPuncS6ElLI+bhK17URQfrOUaglAL3VZAGMrE
gXPjqLUiwBkCM4PVQGdZPcpphXSkS2S6j1mZht+vOT9/dP8v3pI+iGFdXSgPPs2X
L/Diidf6iOTzOIMfQ8qWg4d6o+Qh5ROOZ6L2ug3/UYJq2wBZ4nTTTklQrXApt6k0
EDZyw74B+1W6ZhqKO5D/yY2CBHAz+CF8MSus6BB7VYc=
`protect END_PROTECTED
