`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6UH1Eb4p+UTUg1Fwz8srtwZybkFizatNi00rhAk6Nz9w8J0qCP0prGP5vtc8L2x
D2UDsGDFlWYTen4duIe2rUZxR4Sznuhx86pug1YwL8Bilb2TTuT35jCRNFc7N871
OnMslxihY8K/Wq8jv8vJlpTjlMXjvqMErhqu46a0Kgg+ERXQKAMkRrwuwsg/lTm6
zmq31JbRcrMmmO4i0Mog4LDUdo1szKznZxtspSIV6vWRSYwHuI53FYKbfSQMruf/
xtwUSoeE7NGnqoqh/OSBNFn3TPB5CkSk+ux5yIED04whpSeVomQzdaKdGeUdkXd6
ZGh5y1seFamLScugKXfiOjMeWzXDlDO5TrDhAi75YOz80YhD2COJiFnaKywxM85z
YRm3d47O3GC44R7eiDpgT1PWp8H2J0gWjjTlsDfq1l+QxBBckF0IWC8cAhnVXu7f
Khh5ZkPCOTDXacIuFuGay6QOPkk0hF3NPw8LjE8AA0uWNF7R8BAjFR6qKxMo6l2P
Nh0o6YRevdz5FFIT8bA8nRXHkIsD6VbW1R0eA0iPRoRMTC9M+90+cPMEHLOPhGdY
8kmxNJeXIi7fmJquaNkCQipt4YHlChevmV/zYz5Y47GL5jaCmTHbiC/kTYD0l9T1
0E6xbwSgrc4h+kTologHdWzZe8kwgB0nqOm+aV3VJgK/giD55edoT6cSE3i922Ok
/3jXdCAhcSdBy9vlxO5v8kxiHy6NBchvgED5uhm7Tm7bX58+irG1fNgs4fkBhXiY
jrGb6aFdBBGsTvVfLr2ZmmBbUgSF2eJ1HZm0ogE5l8jVgI3govQ57OzdMQj2MBGk
SE/H8tW9/FcX2r9K0SZM2M4tbUHyIffuRlGSCrrGJnLjhh+0kk/YJ8SheYp6QKFF
ShR9Eb9kqPPGquaJqDKMlMfkCKLIVO/TQ2Rpx9K0bJayg2Gs4MjsBppL2MFSYQ8+
xdGlaPxGxTVmX2nDafCMF5eNz1HMscN9lU0ipX+ZbJvSPUj5JSbQwYws8JIqwAJC
V4lppHNLb5Ybbw+JsRMa+u9e3Z29XEpntGdv2irRO1pVNlQC/NaRf4AVzcqtJPnr
MdYQty4l2WSsrKwz4c80fw9XEN9NhUthtfM/Vv1ttm57WqeVOsjuiF2ZJ7J0Ny3e
z70gKP1kumgBDKJhhiSKN9bOEzPnr5RQu8fwHgL+W/hn56Kq31R6UDRPA8o+Ac5/
oDLlhrfyrOiAFW5Cgk1hGrlfa6EwP3yWlF/opdztbnFPBlZRTs6ZMtoNXWQOPClp
3HxFL1rPJFsQsOyEJzi0iQj3t7g9qGgsi2KkdIax5wzTRcd6k1qdp5tXNGIRpMB/
4b4CtHnSPyJyt/WMt7TPY1WH3VmP/OsdVSKh0RdCob+f1g74F165f52dGUvj9G3h
t6ejCdfX2/pl04YRGbKaJ5G208iYoJeJ7ukDrRawDy7xuCncGgqZcRgIf/tDhQ18
R/6z1svk/hGzU44BsRutI016JEPsTER6IW6LSTNdiF+eFVRcxvgAaBPTLuQKRWCC
gX8FG2IZSYk/3Tl3hDFSbStD2uybyIMmvcgWxqitMX8cBZxpVCdOEicToB6+CS//
kCwQ9CHBCSxtORHsW3KKnr6MKXNh0wrS14qgUSnafMNuz/aqEfEccP4f/er2cvv+
sHW2pztT1HkuaQbAC+r6nq+0za53qasu7ifXbnLoD4jyo8DXzGw4dpq3rif0lFBo
BwpqaHmDDx7fblzWV704hle5aZmEm+1lEoY094c+EY6JKHcZHqrFstEndfAG4cdH
povtS25Na6YzlUl5WOTIkzSBYb1UOwUk1yO9TMxLaJMjVYXN0b7o319g/BNUmI3H
JGee/2kbWGcRpnzONGJ/8j4dvN6D36X2aYcTAKlaDyADzchD2uImVl7H9XOkkNtj
iVY162DzUMskvIRAlTjeEOebT5CzmCay4IiQZI3v/hY3uqUAuN3OccyzsJPkSVTp
mz3qq1ynm1rs+IlBF0z53Weh9ODcW0JTLO7J8h+pK9wnLa+lKge5bRM+Md6hpsBg
lFWZY5ethVqoCMff3Ys44smyTICAjPd0iW7UjKso1fFq0wJGmbOpJ4RBWVM/iON7
M1fU3effvVaRaMdEH7k0TxUwxm9pgfah5iKGSgjGEBBRlDSsQUAhZPo9F+KougLx
BfdCc+m5Qktjq1rWQbe+HmApzpl/MJ/NBslF6YaA0VBJfAzywDq4S3sAfoKaNix0
o4jxAEbMK41m2OVd8MXc8zmGg8LQiEpnho5SX/knbNo3uFIiXqOMrUWbtT8tuPbk
noG0EWhUnG9EIKKm+IHRt43RJqPQ1dIGX8250x0c3jN5C9as3VCPW1le4fJniESk
wKugUBmcF1fwexVbByVeFackTK6Jvg5o397X+TUBkx8NAOCuojzcsafXDDZVq1hO
+gKcO2PwXBRBLBE4mkBFPQl7vC6kfKCmhTVZmJg/S8crue7xheRa8rD5t+GRybts
zPMx7upVWjuAu4SuvO9VfDI6/HNL2i5e4FgZjKBSiN7Ll4esJJyh8bBPnNwGwzAS
ASJEynxItO2QjEFubE9W2EctEA1EomJQylrnJxfPKBg98Q/hQMk1PYG0nCUl+Q/c
Cte7eL5P+xUX5ujKzI6ahj72fn8obwsZwspAZ9EKyVD0b2riCUcIuXUWfN4+W0RE
2GPMn20XhrKVFZJ2vZ0aQ8g+QMWsAvToN5O2lvw4jj0qomdxEKUhW9J1w8MyY39P
z5lt4lGwMR1FhBVKglXb1L1NHvgPedZ99B1ef41cKkfP6JqBXyroyu4CCcdwWVLd
0zd2Gog/zASAVHFP4ljOZtzRrwj9K6A5+G7xle0LpfczKEVWGwoexCQfp4EkL75h
dQNCx0EJQZYZpS7GHFcrcVSi2zSUUdDrd8BZtctJH3X205V3R7G4/mMptXAcuAk+
v3n7dwX4V6tIt1b94zjCrJ9y8VcMOvbiGZG5VG6ddknLp43eIEDV1NCzerUTdM4t
zM6QB5Q127N+sQo+XflIo2Yim1AtH9md7MIJ0DNkilDfGUIkFwMZEchrdA5fMsU7
sLx92vUE754HBx15RDmk6Sl087/7Ya6UgKL0DBl/tIIOF7g7jkcYZeP+7LIGZ3jD
IsXi1V23MzkJcbbw3hSy2d4M6v0vXCSdNHlN/ZeXJkAJ+KwY0ZbEfnlX24HbNjs3
ZaLAsd/RspeHUFMh8uxWJybslgJQobAF9sxl6C+vK1ENHWs5WNTWrNKHjp8hycor
WWUxVtsrRZj2DAJ6JthkjVxGjfJoRAHTZapZQ5fv3fp2UcUezsCyrFm4mWT3kuKS
mtdIL9MmKCpXURx+/ICKLfODALlHTpSjK9vNhDTAq6np9n1cpUwRp+aflaZEboP+
JVLHHvudcg9pD8QVoIiExmSep2ReIK45wsAA+REsRmVkE3dTOzJJ+qrgrFkvMtRq
ZIGQeltcIEu2JpMZO0/h0qZaFxEXdNE8glg21aIZip8STSjMxr2dRBJKv3vj7ujD
0vPMlBZRT0YgF/U5D9PEl+gg0vBnvEiXvQ9alF3KonxpkijFmUEmgknTGhX6gOYY
P8a6tAgwCwNeurrZSCeY0PYRiWsE5rOL02i42uZEGIjzoZsxWRWWv803RrleEQTm
vT9LyCa8wtubFX2qRLoWM3dsI1ti/C6ph/qSzON8swIW6fXXxoxE3mqA7hDQ+5/y
GvECz1M/iR2Rgtpiyp/GJ5PiZe7xFtsHmEwr03MZnyAQ8/sM5Uxu4WEByP3c6xKx
a34XD/t7T+3gS2diL0bYWqGlZkuzA8RTsE9xfxTu2+bkyJmk5a/LFZ7WRl38aT6e
NQ7NQROEON/FILxTudcuFOkl5Nie8B76DeQE1q2uXU3dNYyzgYxOzLUAH89kpig6
/5qqTXakzGz6I58xtim17KmYKZZjgngHY1VpcsE/n6+0yiePGx7LngxWMmdzxfwb
c7rVYDWtv8Wo+W8ixKEg8ptFfYq/+OqJ71GE18rbGoe0v/OEw9AGvInIpyOvi2Im
ZS/hrzRCIcNx2tfkSv3q8IWwyUq7r0CiGR+YatYXHu3fy/T07tiMBcr+kzGD6tuz
BYF87vtyLnlA9lqqFFxomiWSieI0yomsrRriiCClY0ZaGCyOG8ZLEej+dDRO8EJY
r5GVFhEqjdthX0mcOaXQZS1tsnDZmACFWnGBaK1f+U09LZZv8MkqRCAycJEBlza0
GHBAOuBfWwmMfCGAtHXv/CL73yhDldCDGFGuI8tjVD+waVNMvk9ptCaeLc6kz+xd
kHuJN3eY3pCfMO3s3UZc5wGFrP+UP7+kbHvbowh8go+bVOwxQDHBlYBY0bGcRoMO
/U9YEGmh08XlgQqhUjeswqVO+MVNoeVQF0R1qXAacnbHVyFlpq6417v2OD9BM2Uz
FkCSyVzVwm9mMUffhm0GE5vrWLA1r5ky0ov/VaY/12QxKtOXu/MvtSe9MsjwtwnI
BtOmkyG+YXvSe7pr1RRbrXuAYVIGBOSE8L8VT1t2TUK5e3jCQuSqfg0xlUmdzbg5
HqGVRERIfTlW5PAO75OQlZCvj2QUiZ6soxPzlKIVp2MIwMfpG2h3oY3jaIywCuqG
nsiN7QAFPAlkk+5i0KwFHsIxLGLmpNMKe77KVA0/jAwP6rocGy46G76cDfMABxZb
Kv4NYWvR5Xps/vZOlE4C9rjuBlmsMbx1D51e5iWpTOnEC8Zv/Hb3v48M6b/1huWU
u/6hWNRzsmfFdHxp/fP4hkHnHmG0vlJsMi7DF9KPbV9GvLIzDBD0pY7L8e8kNiyO
/GMO3JMDsxbjoeiZwXy7V4iwVSHF6KnpprwzZOB93zcJ8LJTTvclu4mxMPliNHvI
tYCblsZ966vQxrUfShP6n3clHZF854/d35pOHS9FVyr4IBeQC38MXCYwGYEqagMQ
7kzPioJc918kDW83tfwv1DOH4fLSWi0G1v/l4r1x00CTpk45GWxsn+NwLFgTV9Fp
SIKVx2VCD88RFsE9IogRde8kF9HUQQmOHX9hehNB+jjtiK6NRZVIUVUAMSZ0mrA+
TK/PiMl0J2XhFwjpq3vtGHg8ign5vv7SDG7DcKOl9uTEwkZv67KGWNDPFO3x/ShY
mhzpgWzx3dBbOe7zNAwtLZnyymTyXUYzTudifVhlMSOQjm2VQ3/Qgjs2KEPOy01I
bpL9sv/ChB5t1YBxtMrt7AIUE7BrbVmSNqzUnWlIux69FbobiD5zW1trxDHp0wgR
qHLMT9E/N6ubP8lCn4s6qIL0LNgdfs6OlhGDAIYvd+ti4IB82fpX64HPu8fE1YL5
4+zqgEpvCIsF/FWK+p3ClEIeOzebfdQhRTMB/rnBbn4ioGMcQn9fRkfrA8IX1/ta
Zv7Qjy0Jf9F85neSDZKCgySWN6PrnEcMun1aEdQw7fHeCWiA/oef+aaYirjnB3Hg
e122JLV6iDy4VR0l4xXstZFn6IiXSQsIljU4TxOLd8yQ/MeGw+tqsm0HAE6ljgTB
NIEUbtQOiocigv1PoJZj5zn3ryczkTggf4ZHdm9g/07fsJvIm3l3XnZVXPW2oPFU
olLZUrccEcELSgpYVjbs+A70gSBCCpS+7PjVxNTfd1ADL8nyShvE6QV1D2bV6UzG
Pja+52Z6xotZUwiZVbh/vycZOYRew/cTbbrg1qeX/WfwlYI777KJoxuf1mzsKvNL
khXCzoTiPUew1T6dBMMt2hLdkSSXSPLPVguJais3ZNrr9rRHmow/FcDOjVk4Zry8
aaTRh4GNMy3JeRt25zWXloAd0EC9VZ0P7Qbdrt7iQk0=
`protect END_PROTECTED
