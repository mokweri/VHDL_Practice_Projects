`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
17d8AIJepb742r3uh6kgH8PTQ4UtlgZw/c8L0vue7O0DgdQNlPZaTrUqzSFLijnX
ApwjsWP0LOIocwSp9bzxRfVKKC2zNNnsSSAi1MarL3XTzWIT8wZfZvy9sKBgKOhg
BvM7QkcPhJjPFhmV9pyiBbaGkeR3N0783tVJvAEx+sMRSEIXxHPp2gYBpU3/cgyi
3wIajvQkCCl+ZEAv4Od3luNIqNQNCrHTndEeUblO4m5oDlixSlUeHHAK9mxdVAnM
n+ZnmVb/7wufHSx4R9iss5MzOMDTSEuBgfa/SRvFwITh5BT7+I/tytcRQzPYrw1f
tfdC0T2VtNLbya89yDRTsVw0L3Inh3L0St+iqCJDkcd5GxO06sQIZGktyaoYKBon
TW7sse2KMjkaSirZ+9vL0aFO74DlfDN+RIoY7w4x08wP3XbxogTieCQmJ8k88xV/
kRHAponJeR9bD1B8OjWHSoMnoqFXPlvrw9GeOBlaDt7V0H0sqGt6RrO7/rDlDI3i
8xt0+eVpZ2MSTMsyYS6k5W2jEY1zk9IlF3pkNxrCFyYjYYkypw5hEHY5GE2gMP0F
fdi1LYf1fz2IiBwU7YHFAyK1luNQnm5ghHBTSCqQFdUhTWIbfyF7Lfo9C7Mtg5po
PvWN/jrQuTFkkGQSQPOG6Hly5Vgz44XFLeJVJoBlkBf0g4xLomsZVHOMxoX+rZiy
Jf1761zRUEWgSlyPFfK6fVLnFnF0g+7725vrxeD/1zkHlt1pHgqItM812BS1B277
l1vm2+cCoykJnF98EUjI4N9wm/kDdhrjST5CmLhDG40w1GCA8Kf40URlVKwbaYNf
qwHhp4kUbyemsg32jppdOBaTNl/8lw1qJoTWTEr1G7BZmPrDhnSR3pJojsuTf/md
f+4IJmq/cYRj7z4BVlyD8IkTiDgI40jFDIlqswSFRMFKrZhI2VUzuOv7Ezt8+VMV
O5JhJ0HqmlXos3A59LS0s8fOAG5+O5U4fVLMotEqxYo8TOgHxxWM9uDQGv5acYx/
4wD6QtrLyo8kGpkF47cfQT1Ae/uUvCROr5ZsxKaItWslrz1Ocvx2Rl+bPOofq0P2
FJRe6+aT0vvTRF10cuK3nDChXNiX9HPjVMHtYgJf/tLdBaA9yULZscG8BhOFMI/4
00gEioS4mQoJipOmjUM4XDIw0WjLpfkEUoBvCiovPDrHTNoVigfArjk4Z8MBL5Jy
Zrfxjah6bFbf2mv3O2znUQyafS+Dzwap8hYpP8fpWC9qUXbyqLsa8HvICD4wo8zh
xTBL2LoF/M7Gy5ogOVfyyWp0W88C+68RafDVjlYJW+skp4UAREJK8Mlw2yD0Ks0P
zEuHufHKBzMrQn6GfYozMEYFOveCAMN1xGe78Huu9LFoindGTZg2NHGt9Bes3QGa
197DX1mB2JJRYhZ5XXJHq48jvL2Jli5HyARArEiLPWQaDrZKKt2VAxwEbWnADj/c
UoIPb/FNvP3NFnTWBzkzbNhl2VobcnNTfbkbj3/NNNviLoZFLEiyRK/Bx0AepOhA
5ZZzWRkZotwfzNbOdlaYzGw5a4eNpUBuQ1DGMQ33SkNNwdbGBF0ctDDHERX0xNTC
jXBz8Hs0LXVpxs35QSacPnG5jVBoKzY6j7SwnqqJIGNM5tbcgaoh74Y6uE8EYzyy
cbLhi2fOJ3Ydt/TPlRb5CjCAfuxWvna/02IhKjnEzwxoFo2QyA+FMSsCTq8AQ83l
nc1SMdxfsKSWijvz1J5WVA+GCh47lh+z3L3N2UPU13Wk0RDIs36WeZcVCm91nVsq
Va1OK1JkA8IF6rtEA+NwlSqKXnWicIHQF0Qm3ObhPx/Kn2bEFC/J4rMYOsjdePG/
RR6qDDupyrOQcRQNzQAKsfk4qyYm36zUNB4DS4Xq08JNKakVKADry+FQbQbR4g+b
mO/xM9oP7jFrjWVQjvAUPvbah7jMEUeGVKWzI0ONNAufHAypmamx5BAjtNAQ51qP
zJiFUvWxcnqpR06YRmHwUwREgVg/KcxuIH2VXk77AK0aV36njAws84oDYx0MNSk2
0+sCLGWKxwBM8UhklZIRy+GX9XDFcykDJv8CleiCoWDRpQPpmmv+GmhKGYmYcNOn
iYJ45zyapbhBrrw3oKsBSM3p9UIUD1jnGqUxvzRGtccHL9fTlgAgokSoSbcjBA9d
2Jj0UwvwYxDoKvrknx5aAGfFReu1BzjqNk/jkyyOq4JQnOYiqHwsq9Tah1rqAzj6
wzDoynBl3rWIf9uXsh3Nceuw0+W//dUIHZxasAAcYw2YzE6lBJr36yceKaQSJ0g+
afc6iTH3dIEwOVz6dnP52zpd0FbPXqbu/7ehrwzjS9FTFON78BPdLMO/1Yy5KBt+
D34nhjQiwxNZCBRgU55JVjddU+IKoaP68RC2oHJAwZCpR0YRoUHBqnG0yB3Ga4Qw
iv/xJPoBRqwUnFdxoS8fRzqS9AXcAU6iy403Le0xVBngAOsgFSROB9b1vr0+oy8R
FKS6o2hKyTObuCHq3fBwCPms0pNBa16Y0scV+RNXGK6aLi/NC7HDM7KuzbMIkbaM
0w2MOi/lrhdmHWtcCyQqPfah8eIL7Y1xi1MwNfVXrf+E86wpOfrx04ZI+vQWU9BU
YCCXu/8Wmz7MELPXYE+LvDBlHWR/2mC5Fhq4pzWGIZ1WvQFXa0nXgo6znxIUzsLb
utLwOxnXJoSQmiA96uPoXhPkuISnnKF/4/D0RKNMF8MmTg6NcuchPWMGpBE1v9ao
NklUFy36E7TEncPusPR6GugHjpSfTumGbC5epI2SIaJnlfaTZPdkhnxG/Pkz8wSW
GVk1mezPtAutgHH05UM1YmaVLBHf+5+zl+vOPKzHdnmJb8GcPb7fG07fEQi9Qrqe
KfbNHEQTZmtRkuzjU3xx9hYZqtH2FZnATy67x/jvvxYJVCe9S3gkn8olLzBgZIiq
R+M0Uc5Fvlg8mHSbQIvp0/D4NNgAyfya7hcVHAsdttceO4rmBhBuUQL3nJGtacCS
jhnGVeg4IytcJ4zm/eZ/2RBV6LaxjpXS85Ktlwo1UNuW8JnVyLZ0MXfuntm50o9f
5yR/zIpDJ/s4AF+ugpb6znwawisvYgch/ZlUPDLBsgEFiglq0IjbXG2wlEcpypyK
YTJz1ETyfdMyazvHznUEx7Q/tWirrDwLQerL34AQRkjJf6WruoL8MtTFr9fh++yU
43kOBvE9z62kZlOF92raunIq8KnmG9r4IUUxs+rfgM9C2H5GX2uJ8GuN1PjXMyoC
gx3cKiYM0YaSG7ji3lwsajUf2+f0waxgYZyK762/rVW6ck8sX/S3bmgtPh6KdEXv
cqNREMljV78pnXulkMXcAOdpfdHS7tlDRcHDz8NiH7IXE7ptK5OZUGuDvRaCxpWj
uajmAUaF2jbZrJ9GedeCh2FYG8ZrnjGdtMXkm9T/eE+uZ3laXGgXfruy0tLAktTe
xf2fyXBC7sEMTpFUxsVTl+E02c8GjW/KZ8LP/amKNpSls8HD5+fW41174ftFBgSF
VZ9mxFuv18RoJFc14hqfR0CtZFqvkUB9qRdxmPV8XEo2JO4TLqohRF/4xX/NNvcN
uTgVkWdJ8t66fz9XrGP2kgp7U12g6VX/eNx3jVDfsWfU39q1xlh2gjI78uRJXjYE
y1gaWPIYuIdNsLrenhfkaUPaj+bDU4MFMen3aKkHz07ng86+nPcUd8Kq3LA/qF87
lcOarRrCtrSIIa0Tmkc/nBtKvRzEaPYMGZsj417T9vBGGY050/rRZkA2MJ86tKwn
b9O6OY1xMDN148SqTJ7Gh+2E7GCB8Hx8FPpDxuhcRVPEr2F9rheX/4fddn2YDw0M
jB/G0lv7RBSHKpzPkBOC9gA1mD75eh2ZI6US2hbFdFjii4Eg8Bh9tN/w1Y/CwlUf
j/LB7URYoXzhT3JUokY95xh+5Re7Wnkx8+7HPtuqmdodR7xeSKYJGmkPncGNDrQz
Mo+Hjlg79H5+Fhvw6+o4vD267p10XV04J4GsILQSIP3Z1boV50XDXuYdx/EZmVFt
Fi0SHcG7FJw/KQ5n1bHedvnPnFawgWcFr2id1jcmeavAqsqTvcMohYWGICwsVg5F
+iZW8/MLz1LcCsU/0WiomHlQVQ6KRbJFn+R46M3LxU0t0rceORvL1o3iWXkX6d01
lOPsnMft1j8Q/OAInIl0orQE7GtopLOW7AV0JaedibNJK5vMioSjDgCeXIRuyvhQ
bABtDrZXhjLsqCM8/D7ZoZEV6/GFMQnbdaHMctx+OLr2KwYeE6qk3gH7xVnETvRW
whfRojurUDbLqoX7zi73H6g6OrOVMxsp/bhK02ZbHtM0D90pqMbUvf92OHe/UW2j
VKHojYFCXPJub0ox+pXcev/7FEtzHzMiXajOeGlap2e+i79SuGhmDYpSDc0cBYp9
1xJGCC8RAPF6zjrHkp/t8GfnbArQ/PdtiBQnVGYW6lfUcydG1XxuxtfhNBltlZ8S
pleFgrGa/mRzpwl+UoDqXZaWMDcLPc1pAbZ7KVfgXabU5X35ClnvY5BeAZQcu6Ob
GPR3MSjGiQJXyhrRuXcM9NGkqohEfur4669BlZgtIdDPMsoSmmVpr0YW8PImeMJE
jI0F0c1T1r2xmTkTozKQZBGLLJWLud5kdu/SXQTf2nZe24WzYOpvrs0f+4bgxuPM
LAWtB9R3J6UFhiDgofgbPhO4kty5UUqJtsBeCeiUX0eU/LhpZVg8MoRAnFi15ghk
1+kK+TqVVOzGIP4kYQirrOxDnX8+Qx1/ZdYzJ5BABuq0LfyjwDFoxx8I2m3aGWOo
rz6W/qbmyZvwSe4UgmIoUbiBUAUr/RAiHVK1JhakFUGEZfksAcQ2nh4PBuDSQUL1
NjN5k1wDLxaHaYUtqdQJ8DYVRzHraMCvXzYLwMFDesSnO/d+O6rcdXDrEHTrLivB
5w02qLvjiC6aBduHarGaL5GT4vTgtGmXEu3ks3YEr25EQUT6K4m05IFgBRa7MIL7
6UX4teCfYGFX4R53LMwT05YDeLm+2/ap25dko5Or8YBaPWlJ78U4qT8HlqQQoCyT
bSAzYG7xoni1Mj2s1JoeP3ykpnaBgrjKxsWWMQyzY9jnqWfJVX5Gu7RpcP3QHlPy
HXmmCUGliDu3Z1V3Y4T4q5kjQVsimG50HNh1L4kDB3jKooas03jp2xlPb6W8uT+9
Zbd3+vi+PDcKDwChY7Ho6ITOcMIKRL1/mxZZYegB4Yflbln5tFqj4enSLzGUkKeA
FtBwA8g/wQR/BR6u4bF4FFaUskiOl77nejnPtj9Dmup1QCzYSrgRajcRW2yMPW9s
`protect END_PROTECTED
