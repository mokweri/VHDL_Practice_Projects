`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wli5tCa0ZA0Ecgp+hotnRKfCNBEEzSOPuppgcPlM8JGLC0ttLGlVjAsdqTMWI+9
Z1b841faWBZHQCFvjuv0RDpWS+uDPYgNhE9yldUVPsMp1QLt7SnCkwyAvwBBwuXz
STWcdNi3+6NLBK+SwGj5DNzXj05nO4ynvdqt3OM6TCjyO0f0tn5VpJVmgWWgjbUd
YXkKz4J56Y45KK/QE/HxIxxzObaQU0uxN5D7BqeCCS6BImwoLG6s2ASpS0tLCXjJ
ILg8L/2JTmbX9kTwsHYKuQY3puB/5r+F4bE4ei+b7AKfv9iI23IviVb45ImzG54y
E+tIXNuisvsfUE4OlVLPDrZKIiWa7xorOeg34SXHTgrJ7DzJrVkNy9IHPJHAIRnY
cGp/FINBFu7souvKuHmcCR5DndjXCOmLVCWSsTvwTnE5HKhvaKyu77QaRM5jbzkV
ijkmBob+xpwWGY5RW1NWALZn9/YjFyvodw/KSkjFI5OFFNj0B+oVPOy7Y9LLZaOK
3GlKe9dhWnSEBJEnKrnW8xI9Ro/kPm1w0Y83D04gvgAQkxUV8bNoIka8ezUs0Rmm
jsij2y6F7Ta6Vh7uCqaz/b7XYHgZ3auQwAkK8/Ze5wSPWIGrElHapn5ofOYeYlPT
ANzTh0Tw2ZsLZpkfiEc9BchY9TE/Ivn0UopwI7Pstk4mv53rP8y0eeU5ebkNuRfI
`protect END_PROTECTED
