`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4f4J9VWYZq3khIDmIpSYAf0b0xcjLqc9Wl9fV9gx/yv4io72I5nFDolrX6Ky1Lz5
aUO7n7j1c3/FQGDdQl/mryq9puOCdvIjOc40MHH5ycU1okVbpKyY1D+gXXGULtXQ
6BEP41VIFzvWnP/mTR/wJH6XiWvix5eOBb9CpIXTicZHGAw4Wuf3MBZmATdWtY/+
un0i9SLuLAybUAPKi/rCZ95ZFDfY+bcJCCGrIjpO+L38soIJpGt4DuK4ppDLbOLs
+Aa/IvmdhiaTnLj1wa6TWU+GEIjjnWFzHtndnCOK6WAsoO9pzqwYXibu5bpTd/DK
4xBDf7uu3qS5rZFVa9W/UlvMQyiwbu5HWCc6jDeNz/w5kXHJeoVVjLIIc6NlLpWw
2Q1pK/a38YypayOn/2lgt0lZWyvneBx28oML404Vlx0b0vdMAb5uXh3ql89eGlgQ
VB3sOU6SEZ9/hKluFjfTjv0QcGktt+CQDGnQmgfKbECf5U5GXJGFRHuggekAXNvx
0rkx/MNWrKgLL24nqMXN8iltmXdh7cuWd/9qKxgAPSqz0JzPeGjEQxNu311soPpz
XuCfk0oGrwn+5X9uN9OZXZg2KaeSg/JcVyvXy/skg78673AhFKTr1gHCYcGVWfEa
BmKCsfTF80nSTzsuWouZkmvCvp4fzAXMiE2mnVWq6pH97UG+ihJDzLe7icwcU4HV
+edTI7FU8yTWtgNnElWKiwMZhDFDzhW3c2AuY+3tVvJuQRZD6kT1s7tnHtKHPj0m
Ni3A8dvX+6vmzRs6+246U/VVjCRzsd4vu9EbRth8cgnftlE4iXzJ5aA14ZNSmZQ4
IZIv9G6V5NXWWB5rrD4cHHrkKFyHo8d8aJ7RVvG9j7pwzpNDQOaow1eX6igDLHiU
wj9g8fwgGkt3PgE3BMpkKHstX8MAq4IpHsTCBtweIgTd3EZBU1VJNxnTRQfOKIYT
L4i+6XvaTRMYNlm46bdzTsud6E4jLgFPl0nc4XGAbJ7t1YGByvtQikDiM/3NsQoO
MhKlBw5VRrwFwRFMFrgRmXVKMTEbXtzK7La2VNJ4M9pSbhdqN/XO5ZHDmsralszE
BqkSTWBl02RdlzIyK0aGgJaB7eI+LWk6NlZVRCJRatd4qFmwga3TFpgcEDKUfDYD
sjXwS3TWn+LC8cwY0CmgC653sHwxf76jDl/0G8AA5Rueg1D/cvXTBjqFK5GCX/Eb
ckz7gU8aWMrftzcN4tX7Dw==
`protect END_PROTECTED
