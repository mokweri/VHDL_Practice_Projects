`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D16QZTWqO9vmA0In+nTwhDduO7QcRCHZz+rpB1jWtNagTmMAHkOeFgCcVZEl4zB7
nHgRN/rRb0d7PQRF5CdchjrQRNRMdP+endBTb5PtU2dVEHAiANEJlxtZtMSFjxmb
r4oScY7LTQQCFQE9ev/iPmS9EySvTJmzT+cE2k2UTBza72qcy9zsF5r6KrHrhrDY
pU7PluvRIteBFxbrM00D/4C1pOgVVmFPxO7nzAH2ZQVsnPOknjghakydZ9NrDtj0
ySZPU9rKwNxkLeggL/EWXGN/nWDiN2EZVIVuqGjeFBcPWD3dxEbubrz5s9hwTUBl
OM/HIVddOJu8qTB5ckV3Szg9kiUvZesJmLVl31ctliQFIloCdDeCuVCYSCEGN5rx
TH6DMrKbQuPDpuC1L/zAlqToW3pyGv2bBk41zmbh5/Of+MY7MNMuKEXCBicrnpIK
i7eIrD8fwr0RB8k6pqvhWPV/77CkOIcGPl9o8ZNbR7nrHrt6MCXNZfr9DPO7lhYU
ae6HFZYqyzffkJq4VzsuBbpioOW308QepTdK13gIMOt+BgasI4O53ka4bOdid++r
l7kEEMUPpA79Q6E4YCo5R6LFaQMbQ7185O+1DK44VN8TtYGBIn+Op/xG67UFlJmB
YtbB4iDiU3pwIdyaHZi5OU3g0GGA3YZrPeIy7CdLJpPFwC+6TyT1/wvIY4RVjPbi
Ovk3jUbdI7xb41acg9UdkgV1kVkqyt1sHcdvy649TOTOFAGsCWzHLWAZB0RdqcT2
6XCEBMc6u+AgB4aNXvZHM9WdEeiS/3weEkBKvamcpa9ueJXjm7oRaVLcULLeDNO9
XT3hCOPGvjSuqBuqFNa6eI2XrHdKLQeb6RPMCUltx0wHPmcjHmDjo27yYSs6xH0Z
vVvGOd9oDlH8BH61TzJRhcC56oDL5NqF4FBFUStCbMkW+mQUWn1gsJC88P+LgPyd
yhpCXBBqXFOzMoImFj1NHYhYolw2b/kyr3uON6g3HnFilgsMkt4II2gsCa6DE0lV
b87IYJb13ile7gFVfw7d3CxcV3913yHk79hq0CLxS6EEpbGyZ/ZZv9BCQsv0QC2B
A+OVPWn6G393pDf1zqdA1fPYFn/5DySyQ7wpgIIq65v/4fCEDs6+9hC0keRyFC4Z
3RfR8NQFN2R2wGcaj7IByRlGwBgCFXMUZqtJ//lptTVvSC5YtSA4zWspUE0Zj7z8
2M4+pyiXDK7CTUkw7/rjUAEYU5xbV5FVEmXjI2ykdHRjsNjyBM8z1XOeMEg7h6f2
jp5ccS/hgfW4f8Xai1sFcOjrcdZcsqrahgSXSJKrlWn37KPQf0sa90voBz7OVRX+
jST3EsElioeg23NjTbBdSv7HC4CS9wFpUbLpAqyG7dEaImUoGDUI3mL1rCgOyRJV
IXbdgWx/7DeoW4mwznbLrA==
`protect END_PROTECTED
