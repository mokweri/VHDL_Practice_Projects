`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kv7JAzHWmLMjilLNNpVgnRdqP37So3RUcnse7TQtUxo8n2BXN7LhYJwxw0tImDzZ
08GOyV3koiVT2YnV1T84mpQWE6S4TSZcNcaPNquctuwyqllZ2ApbFKLzCZ6lg1oI
mO1sFV3iSxUKYMRcT57a4nfEXHNdAbFPm0cJ2Phcal5xn+GJ+eGVl4Kt9xGaluve
XGpOFn1RdrkKKF42P+co3nxHUuiO6tZIGAxcyX9dJMmM4Kv/xfJAU0NeDxanAsh/
pBekPQwL+L5sJLcuS/D3AqOyjtOC6gPUiCTv/UPsU6nosIwjvo9R2+buwNfCPTB7
fpNYJEYtVYGXtwar5hQWn7ZHt0YVKluA5Hg0GYIGPioePs1o7skReiJhtt4DEuKp
`protect END_PROTECTED
