`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FuRqyCzIlS4HMlMJaSEnfmmNT60n/wqwN9fNUSK9cClUt7y7yFLAeNrmaQ3I/fH9
E3pU/x7i6TXAKQPOduLbsz7Rh5VnCkhDnooGton5CIucYhJDyWKhg5Sx78Zt8E95
amiVxbGZnsdpQDSk+9PNJUSE+aPU5aYX/lfhf2jIHUfaLY5POHRxwyTH4eVbg+Kt
u0Zh95z4ku3/yd2bS30CJuIY7oi/qjob//qh87XNXzS1wjQaRQdvVyFz/GQN9G7b
ARSwFWS9ATmog8nGPfbD9GQoKL1lW33nSpwj5ekXQmfcCKtzrDXCTMEDlm9A6JJ6
d9J+MqXjxSzMlhfpjaZY0BeZZdWjS2uN3Wt3VAfOPn8Y8ioxK/Esrwsu33tPyVKu
P2pbYbUOZhIta5GROJafrcMbnBnrseQD6e948ZfSqfkW2BWhLMv/zAYGK2I7Uoe2
JpFvMfFXA+bfccoiZaxQFb6lkUDEdR2dlXRUqcRwLFvdySWfKQsSRrtzJZ1llQfk
zFCMIrCxwjof2J0Vij/DKpJfcgF2xHDdwa+2MYgkJoilNQ9GL3WdW4aJZTxEh6c/
xKF/URRG0qu9SdG/a8thg6re/ZjcHFX2ZOimRWn8Q0WZxWNWKVoycXylGygfYmJv
aCfKTcXhjpl8+yBggD6TQbG8O2CDgkhtEFmyC7gq/FdFV6p7MR/0p9LEHzRpx9UA
nD7psr61oOjENqirVuN10PjYsLCO6WcvKGyvM3P6TvNwDtUl17cC1MbEPq7d5whP
HJUkVGhDXc7LkSJSYjC9ifHauphayosGtNEO7Go1AjRkmiN2pUrovw0bbJ0nhGfW
E8FH2BTKId2w9dzrZxP5fMp/08eBQiNtwak6CmfFIb85NlIgS0XIq9sok401LAHr
4uW4luhKbDgQXFvEvbve9YYh+kdXGp41BzmgDc5WJmIkLrdEY6QG1EZ5iXDKH819
ILb2HMK7ld8qyOaA5drfCSMbsCaBriUQwEWaPOnYX6KmCGSRJbyLGbROyAhV9sYH
M5pGQSBOPcABKLebm8BM6QPJN329eU9UX7I30QumaACln466t3793RZ/a+NqczkA
x/roHozZFuCx6TB9jr5FnQpLen2H5fLdrk5FBjYdc17pazM89BmXxABwPCjZF1x8
SRYgNT+ARSPckycHTlKtrtApaxpljKOT9FYW+Aq3IH5eIraYgr3FPnRYqHW6qBMi
hUXTC7CSuIMJoAZipvCEY5eHghjPQIriD2ShrEIHAXL7FL72seCxK3SXW1G7+vEk
mKKEfzC4iORpCu0cobqTao3d+8fH50dEMG3EknzW57QTiHYC6q/2qQtKE3kHXwkL
mFamMIc+P35qOyltpHvB7xALyZdfcbRcdY0emum7fuai/FtJn5yDvevSndMsIbDp
jEFZCCjoqHgGvlzu95hQQZJqFRiOrQIcD2GBMswxnPuvU19geFSk7+upfO8rdg6p
whfNh6YpBeQvD5/N/yJXd2I9021fFlmgH9G/7/p9sENDS2K6IJravooPAvRoKBeC
wxaA91lAJg8850RiLgPmqprwyx29iL2UvdOp9xPNfbsUa4fkr8mtADX8Cq4bwlCO
pdzMFw/5mqbz5rklAJaURh+fSmeJYjDdcdn3Mnc8rcNUFDi7YyLFNekHw6y+KLon
sWjJahBY/4cCXIeCb1ByRksUH/1z3j0Rl6TPDfLNV12hATc33aBilZVGSrCpjI2Q
5c4lZiNKrXqFo6909pAket5B5WWHM+V9o3qIBKaHn5mE3WQO/YeyGTRNI1MXln6D
dMAhnCBI8+Obo4EQzZ8SoYEHOHFKq7/LS5mtCcsCcM2BHVc2Jz42XAWonpWq9AtL
RpaH1pYe5jeoj3++DNE2YPJs1DBhH3RO49u96+wZaVSeNTKlwe/r04q1KGYTott5
exi51Q+8X4yiQ2y7lYnV2kOvC75ADUx2FAnrLidNbuQYp73ueos4ZRMufDFcCq/M
9Fe8pH86/+0dieMK0F9/8BVt04ivpBVPKNGuWActJO3GaNOt+2Ss/KjrFgmWIGys
/Drk8+IJnnifBmR+d0sGiqjEScYPTztkrxPq85xqkmS3iEP7J8u5H/c9b/I8ma8V
o0OskahPmf9Eon2wcM6CRgA88/z8UJcB8LxDuKWdwAm+5w40cvj5HceNbg1dMphL
SZgyDPymqyvX6DQjtoyP2W/0N3+60mZKxXbvf1NkyHIyn08/GnSRFQtLzO/vZPTc
Mdmj8+5Kk0v5b6Bu3mVLw4lNDXTJL7DxfAFZpMQN/ZjlAvmHGAiUTT1OPFbBzbqF
forV6Xi8xa76pBIJCXOBNXs0xSmmo3SZ3P2healV1n6Nh2FiLtT5GDox7bTziuHZ
tck/V9/PZ18N8ADJGe+9SfG3Pj7FGOcx5ybEhRI5ht0eRKVzyd5HeyVjZ+9Omi8J
hGu76moYdNrWX3lBL1IPLrkZsJE1VZ6XtcmuWJBin4RkZqB/Oc79/2N3Aw7VJxnh
VbvSuTmpAzaHVgGjPAjVofVEEx4oTuUgttOypY/GBfMoxjUapmK9P6PtDOmaBuiP
pzo4IfHHU5jE75UVcPpZAgUlSkDx52yqnvuRkU13Elg/W+UG/KwzRnuGiSK2VozI
wSXKA6IbWMcXgpSW+dEkvQ7iJ9pe6qhYsmC17iBOOaOdMx/RrXxyJ0BFqV9F3WGp
OxfAyX/HWtiCOtN8dEOIL1tc7k2H5DoCU9eJXRpJFdQwuf0JEjjH4YoiM76d/ZlF
KzTjAswgqXf8ZSh8X+AF4du907u2c0UxmB0fzYV+COaBql6WsWY6C4e+E7rcPywA
q+KFkcAaFJi8RxBEG3hjjJrDb9nRf+NSg78bBkiAzhJK7zjz/TAztWj0QP7GoMSd
pOR/0JydKih1IuIJpNvG7+ERoMX33F32j5R2TVLCzHdazIw7AhcjHNXiMCd3PvTp
TJv2BO/viLpd1peZts69oZZiJRaSHrRLRjvI0ZHMTMIcRzlOaBLFOPaj9ZdQTRXw
MAc04cyhc1caawMCTMexJdxVrkAruu4jucohDcKPBb1QYzCfyZ83MOt/xi3pHboc
9Jhn7EQ0la+HPIFvkSulT41ID5XcjSFJXj6VXF7QcsNieZL01YD5hMsYOeLyE60+
6CmiYO8J4ykuO6vkkSSuLqBk2gIjdDgJJQqRWgsk+xI6s0My2Z1GL2PtcOuJiN2h
5EFIE9xadhCmRjcQPQDpKXXjHInUbdcRi4uk37t/swKHxN5DOIS7sSyLA/y2LN3K
zY5QHCNB/DzS+k+TT+4zIy0nVfePbEnMTnQm+TyPuqe0ZYvqV8Bj1ZgPwcGKJFa8
Jp1DnWC1roJraCJFf9kZn15Ed8duf1SLobg83zWXu3tLzRHp8xOK0C75Xy49uDiT
gIUgMewsuacuIRq4y0jjYsdVbfd5L7JidtUhUxYvcyf4REbDp0Qi3fyHSKbXSOZu
k29qmP94NpfVEEWFiUhbACaUoDQ2F3M+P+ptEtZ53IJxjoS9fX1bGKRmlfl2hvkX
43EN6JO72F4d3c8yUiPxl5RXVrwMvZJfCXxH0Ndnh7tqZyqTmJAnE9Uce6aE5BSA
iH2Pyb5Q+/7LZVwxwF5Br5cZHudzeQ9ZtJXyNg8R25NiyJ53IzbX8nAJFliU9tBU
fe6CRe6okKY4eNbJgZSG8NUA4/NwYouo0d52U/psE2PwuXlciKmTvqAyjqgkdHj+
iKr2b/TQMqPJzvAGBcIhv2vyywpaoWUwbO+K5Kz/1Co2rPmlW1vuywlzqgbLk17W
TK+YEBeMZ+pAZOs0pj3k11ZsRT3yvw879Ez1DHswldIXH3sa5bvWcA1iYUh5+JIN
NbZld/begH/CvG7oj5aFJPMAFbN+IOhGMbahmnGzPzqgtVGQfd8rk890r9V1z9Tq
syEoPgnSreeK60KRh4gsRTL9JmSGsbD76bauOUVyZ4ofwbqegNBXWR+SSm4dFG1O
p7Yvirxm/20aes+RdylCaDC5yWOABxfOQvjA3sruAODLgThEp7BkyJtX56/osP4y
hdqLiTMcog2AjZw58AX7ewZ4odeQZrNVN5KSWGAqoUbVg3HDEGsFqtAPnINmrFGJ
29iq431ojO54CLWPJMoMJuljydTClllBhsfFF5u++W6q9+L9n4kT1zftc0AmpUl8
tzdZP17B7dxCAUHbuLiB7aD7UlHcdPYjMBKMMt5StWOfF39lvb/bEVwJT054TVD5
Sa52NI3ER5dnvo+fDVAmhZnYwBj0EeWIEvLQtbOTD2701M1261jRyNU5A6E5gNPD
PN7NAiJMKL34iFNbx4CkbsQVJyeuTE0v93gcjHeiPL1KzqI+ashc5dbIebJ0b6AC
5OgwTFv5ApEs+ogQ+hAd1f3serBc95/KILV8axflGLJPHlbg2tLM73IjT0nxa4yM
ciFAxgfA+pcAhjhBUy+NloYdwV2xIGNmTj9ZOFbD4jFy/Itugbiy9zZU33aynx/8
hIBQLLU22hP21vePJBoBH0ZGjtKl89in2NmpFLJhcqS1j/BOQxkMoJmy6g/CoP+L
TxwNlu/D9ZBLzjA8zGZ9XZqXDWy45MvtpiTUZyHBBpUMC6ib5ecX/2/BL7QImvBV
kWVT3tWZxB4CSQcpEYzT7jn1u91VBzaKdIEpzzixj9WNw4V94YSnrTacRk79b8Dw
Ki7qQtq4/MNhATRq4sk+84fCP5QiwXkPWsF0x63kMdP+Q4vzw7VCJGT2RpFCh37x
vtAWyBp729mOyei2tvW0WCVJD0m0qO9xRx9GCSsTwlGL9GFor7Rg0miVqgTDDq0N
/WoCI1rEsKzd25T5HkIf3LwhtWa+jSLUHCIh53NDo1R5kd9D0J42KfMa8CSNLWm4
Rii+b2Ga40Q3exMgr9SJtYUs2x5rT+KEfTvl4gEwfQvuU++cQ9RuV6kX/dDbLIz5
2RycFW9KBvy/Lc6AfK0eQ3t99SEVXIYbGw2VHIaw/XcA+xxSHkA3Qgu2vCnMBpMI
Vd5Zd7NtO5TdUTCBZL7tc6tHUYkfnk8F+l3zkS8s8wZIqvgVm/mFwHCYuMLel4dn
J7P6c6iSkuqqSofdRV2mvW0pd+zzNFGMcRbwaadPl7T8KWsUUcJF5TCVKcA42dbI
4tomGqLcy8J6Q0RDyGo3G5uDcuy1Krmuz4o1cekEbhscie/89Y6Fm3x7Qhv3FthG
gwnH7WCj759hMz++GecAq9l+H/iG7vSg4HIpuewMsKJNbPwBLpKl2GiOrps9IyIY
HSzKkSRss0A70K6VyjX5QQergDhLrVDpBSwgOTdYkQBVeszdA9cBB5b+01yVwcEG
vqU+VZxmSFydexMe33g440g9vt0e9HraIcc02RnyyPl/OO0xVqflJc7L0rSNhrkf
PslgzkZKlVYn73bpd1X1+IHC3cD0Yefizh3La0ryGkV3ORKzQVXAAVbHHl904tUL
CPLFyr7o8OKLya2mb4AW6EbHtFnRhRePUGNfwfnyXewMcBKe2LOExw3FG1wIWk//
fvgbtXHR2jhkmE2N6/jB+dRDHmGNtFYZ+Cj2UXMVFMrTkIVdBt/HhYtFt87nqjcD
p9xUg8egLBCsL+dI8GN48AxrgStvWBeJoGLz6ZVptSFw7M5bK5y3czJuspyL5saw
+bk2Hibpp+sXuZunhSyUpI1B0/7IRS7yOcAyng2jy/4CbmJ/U3MMV9h6LizeN0Ss
kXxiH/qS9ge12sBWUe8vCoHju+BZpxu8Msygr+3joYk3z2cqAIOpAuPfxrCKoz4e
ShSYitpxH5ViIN272kk/gsy+tEIhC789AmhnCAFjhm8s0QzvpfKopz98ZZ/u52jl
Wz8xl75WCuhTZ8qJK240Vzj0oLvj3wjXBuCB7ax1GuZ1ZomVhhtbnagZxuSFf5/5
kTakHzvHtVI8ImDlkiF8lXYPtqeFu4zYO4SXSn/2SUGfBRpfwJZQ647hXovxuqR9
TyCmqBo4fvTmFTEws/QwrI5PfnmYnvbObYuAPikt4SOz/a7SZ3O2IV7YlY6ZR0dm
WRWlYt1ezGQZ/JyL5uKfzOMsdHxoZeCcOfMw/suugPhvChs+YkQ5nQ5pCjFst6k3
DY1iJ8BntwX5up0Myannp2xVWVMNjzY7bR44yZh7FHoHZ/TFhClFF17bRmJscIb5
RhgL4z3qJM2AvUMyG5BhG1Mymlkql19bYdvCt58q9XOL6zf0uVg5LvQ5RD8mijjl
4EMChmIGpmSWqrlJUvRuiYELfs/2ae6688i6tLsxvtfvrhPkpa4beewVAk8eg4Mu
VkUgHnX/7/5jJ415rmnhN0qtXN99C2tx3IRbtF+Ie2MhlcEKriRH7IEXQLznMzs3
HtocV6BAhu+kHvu4YuJDSm0jep2sq9tBF5Qi127THWcQk7K/xvycAtA9tiNBNm1Z
sIiJ25ZwZM7p2a8eCnXRzuwHkbRS+AS4hqhUUOdywuXMBzCJ6aO9+fcHM+zXF1L/
+YWCyf5Mzgs9u4Z60uf1lWDllomqhMzn/tF7vUqnwNtBAnxGx6e0cFEe29lZ9uJK
c1XNkfLYtP/iE+qoxEA6AeOSP7+6qMrdGqHuOK783PUoIeLVxQa87Fl1vFQjsdtl
aKfg28uePDNUsAgUr2EPb19cWUiwdI/kpYTQOc5/z+gG8nICcIb8we80Vjqv9ecB
ONvECWOnk35FbRV/Xi5gVFrD7Ayt/KPiMdtFsxudQp2FsbinyindosBJxbHguObl
vlwMXM+CLjWZYwRi95DTYSYK3BDqME8mkicxj0TYUx80sIU72gEBuokCg2PA5egB
dOKP/X85kJLQnOr1BNNeOop207sRBcjJz+yC8YlDTFfm5mdpPEmR8/UqGJcC/QaE
3V4Ym7o/zQiomrIU/qsmX40yy8nK8QHDFF2SRsgHm+GLxMn4xymQATSvFTF/6IRS
ahPuahsTr8N8hvh6T5pcMYcsXSnAxOjHX6BxPQDaoPMu2KGp110DLgvpw8lCK8Lf
Xfo/hnJ49d/JmPtM67IB7EDh1xKqwL8q0MeE1GqCX0oO6UO/B4OcyP4vRXJCJWCm
QPJmDWV5d7slacYNQZBj18SnW6E+spDnpX4cJmE1tPezT0N9fzngsmKVDzYq9dPC
AV2t/ikwlf0dG7nbV+Zniwmx/+mWA32zKcMHB2VpsBYaNNyZmFbO8rSx1okaz31P
KcOhEgP5ekQBpU2aKmxqdafsvnGsbVJTih3uNW7uQSZHOdGRhEbGxv0hJyHigXAf
pqTD0DNmFF3kILvBahllVgJuasaCsOncf39ndpsGZLASEK9FVi7Xs//JTQP2dIWq
1c2sClm4cfc4IXuLG+JZKPaL6MbHTGIMZbRzGzvNZqV4H7LHyUrESrcUIEGJRw/y
+auy+uOUrr8F/2UfVRVtIIYjGs9vbTYW8s8Jcpm3pH6s5ccMOoTH6ldDJrrUeNOT
vba0FbhEGf6V8gwrsAgGgL4LMqDND7F8cJWOgoXpehpD7KgL5lIuBCuSxAG9lncf
0iCMNR9JVeAodvuVYBYiOEzOQSK7xV2xFxRNl3+EJPvNeW59KLZqTXo801rh1NqK
kXMVgCHq6TlnjkFhUMilgLJv62EfHfKnLiZ17TaRIEW2G7g7p+/fLvRx9ckWddjj
1yYvVKTbyue/mT/OkuTAUd+4iBAPdaQi1GO1H+R5nsLcq+9R7ex1IqOTUUNKeLX7
ZLigJfXIBvVqV6Zt4+DaaeHfbbebeqA1gzy9BWybvXgZcG9jehOKqf0Bn6eHYybA
WLz1xPDxeUv6i++PALVWUqvESDKOMWANdRTpsSaXiZTthDBz45cQfEadMkRxNe8z
86oVOTbPT9Bi2bxypoZC/NG2yWtNDsbIFHr57y7SJ+BBVbocw7kSaanUPzDvjrBw
tnWJDYTxiFZF9kDQR+gCueM9Laduf1H8h11hXIKV5jl5nd3C1RnhvhCWMULNKnDR
5H2mrAfsXEDuymm65JKDP6NZVQEirhXnuFX0/7bLv2Uywpd8nt1Ev7b+Fil08ZQf
7Tx0yuOfCvDcJ9f4g1+QSZsp3lyDaQ1Uzg9Djz35wfERutO4+6oWGGD4HlNTlWe4
VKdlmngk1h8gl9XXwEG8ZzLLj5Nxk9ap6atV4DUK8gSACiRJ1nNxqFV5NO2jKCVf
jiCk0vB0gBbyjB453nqoTlzXzmOuSqeWaEbzDipEx/iItNhxQcBIlNDhfpNS/K/r
wbaR/7Brwtp4nQQ34OtwkwYNSiCV49Qiv+7zjSgADM7yhFrnJSrh8KsgaVXs3zp5
RE0IAWL/nhw/a6hlD8NBNEMN3KdS58lEtN+s58Vx7lJXuZqOm4TwU6akarX5LDb9
BtTfSUB9M59eOLVnxDmV/Wqel8w7cTmY63+YAzI+SPCG0Gt7mOtS0EzReU4pw8bZ
amZ1SrKaBFaEL4TbjkzLNXtFQCISgziAd83xmEW5Ce1Uqpx5iWyNMLuaWd9hS8K3
j6DNLlJA2c1LshcQPExvdP3rV4U2jIvdUvCR0JWGKjZCZ6ize5WjMuYfNg2VmXaR
ysaFVsQfs4ER/LEWPx9zJGBLsL4eMK3Mp2syuj3eayJcCJ42Nc3jUssbOVb5vXL7
bcpBYAZi2KgWVoBCAU4X3pquFPB/Zn/j6jwpH/mQa511lUEaAWpVr3ZC8RmGE0u2
dLmCD1gUUKOZt8T7tqcCQZkxjbJ6xcQB/F7HIE1mUMdeWvWxuIK08DTXwJtQcMbn
EmBmjiwpGHyer05XtP/zpIqG8B+jG983CJ1MIWlWsDZj3N6qhW3CYkKgIiSApIMi
VsnmzGDnunM/DcxJx0FzDpxPG+xkub1Q57RiT2Q0rkhzMRCNplmnXrGzHEujTN0i
nXcBI7BzYOWOXrAYzDRduy4Eq3szXfzfMFZYZbDrtCpODGIS0d38/cpumcfNHEYo
OXCLIFsYkKDCa0KgYISTJkOfBZqp5+Rgq9ojjwPPQRjHtybu2oK41BHrZZnNoKUk
APG13+VFWwSenTlOJ35h1hAoMqL7byyZxNsZOmBn/GW7ZYzqPxyDTuAZ6ZtPbkKq
Q+mT5udQm6rBPlHoxGsSD2YB2KkJmtGsPX2304VlzJwT4898SYPB8qyNrUHJ82Iw
KS1cGT2KzBbMi61rmHb1ZVrqd9bVFXPWickIRfLC4iwpaHVs4Z2/ISusw20Qe+fx
gMcpUzWHhAygH/nZsnSXnrR42QwtGGZzEBsl6wCCe6N3/Bog7BF4ecLiJARPdJdO
kHp7NX2SrmBcP7AxjWOennarmllN+X+Vc+I8li6GHDsbsaMruM90nCFHRh+cMIaf
QoTMIc9VeOwOIz07+DNx0aHtcuAqTd2iNSBDx65u1xZMR8LxpQpBcV8bnBff7VxC
Lbq2676eXTON4gNr4R5vcq/nC1TW6RVt7ijwpYFcXh2RKZQW/UBeUI518j6bbYIg
W5266pHWNndquTj0vsEBfjvMsvRMRMfcxWHaATsWybI+qr+46gtaf5U5vBCL0pZ0
2Ru1MJvT81iJ4Q6Y26osuQjvHRUKAcZu24keQCOHF0hBAcDDy35Ud2uOPGkqrTsD
qNiZQNX3NUHcGVLkXXQO7/49o41O2Iwyzomc3p4KEbppoBDFOwSu+YodLovhcE0P
Y3an7YShPs8XYzCaMiG34gV522bHO9WGtf/TgNABzLLeHZFZczJVxK/Fx95kfQJo
76g05/90sk/ftv0sftKMg99UYXWHDRYVBzBC7Sl6olKyMxasXaG+Ck+Z77NTdDpm
Ieqhgv/eCWwI6aKkupspe7ciMgdHICOMXYi+O+g5jQZe/u8Ljy9DmRKhV7BozvSN
gJVc851gSKLHXqKRsYkkiFgtEj8rzj7zlpY7vP7aTHHLWq6jnIWMjvt0ONqtZnrg
CZH+NVYInk9KVg6nxHFgX8hsYvDi/ShFrHBPTi5e8uPoUDz0ti05NOo7Qe/LJU/8
4UoRvsKR1skWVK8oWZe54ej5D8MEk4FVx0ecHPVcgrYVwOUbHp8CdtdPpbhtjZe0
Xv2n/FJ8THmvWyMakWceZ4sSAWvKshugcFyjCiOVCDxcJqC95kyk2FaXk7EOC9uE
fYbjJbY7Gnpkxp4uyGDKXe8K6uVU9g3E24tjXQzlnzcvg1xJ8YQrHfS8MCOOY8/h
Ef01zrCyP85Vjezx3PUl97pgel9zDzRdh4MvYoek8+26v1ASXSAdgqBOs3jdw444
7rX63WZMdP3Rk77NJOrUBKWBlAnbQMCnUjicaE+O6dNuZYmEiR5DpuWz8+9AuejC
2REgJ5P+FMcQS23QR5HYkGC9ypWGUyA+VGgF9G4f+5KW9R8s4whwRT5sGh9FcL5a
AWQJQe5s7Ytd2gEK+z6CVXqJWamijJmHC3QcIvCOqhUt6E8aiqc2L2yTkoil0KPc
8zcbeM7g6g/dghrKyQpjDZTOKQ6qC0E6ZEk5wo8vdRA16PwEeKTakCoNlKqpzAjj
t8P/CJg7CfUI2/PQZqm5dc+7dRpNddxL4OZSR7Zm0fibBnZjQ0U6EeOEoa9i7gzz
Gf9QUsAVuYQXlulz2do5fUIjTX63be4mUEso9uoxpKIifYSQxohqSsQIKzPIjMBY
BuYGrOO/mO6KJLdT+2CN6RLEqjjiPy+LKG9NHXdodq84bUOiREyCVwSwYGcsZskb
IWurYBf3f+Ha6sT56siXDVbEHHtCxOs+PQTwGNoO1joH5Z/3zeaW46PZD5SjC72s
M1Z0Xtzu5z2L5GyfgTAVIOXrNCgGEL6CZh2TvlSPk9Xas4XdjSqUkHPHrfCQgKq1
v234NdjuddIPfVsLS40ZmmclCUlJ/OqfCfyMRCH0mOaj1PJyfwYKAzM5scr1y2kX
aA/7VIACZviZz530GoeTAlAZRtA+tHFWLELtv7bQTxc=
`protect END_PROTECTED
