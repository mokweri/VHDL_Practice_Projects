`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39M9QKgU9i2PYfmvmcrOEjtCFeGwvXyJtPMj6iEEZE0ng2pntwNEbbzw1Ye+2e/5
yQy7Z+cC7FZSDdNdg3YSvCMJf9CEk875iCLMaWyRhhOWwBTsJckJTjP6Z8QRWhJC
LrnUT69OyspzGp3JVHtGZ1Yjks/wHzWM4i42iN/HdzGKKK/bxBsngZn3/erj5K4w
yboLG6cGQYQNsurjk6BBE9899r5uhTQROhqiGHXAfkXs7ecj6Y6SUwmNVNnSnyE1
gJxt0idGwtyZCmhQ50jh0rxtMISpWOGEQ/BI54wl1IhBpMIPnRtI71xPmVrEDgpO
AHnZ9JqbD1eyTHf35zs1RyVoYKQTH4PYoHKypbPUJzc9zEYxO9IbDbRoHiRWQEvS
HzSWqD9ShYPZBUfBFSPQtsXVjzWl/6ZYQylTMfIT0rSsDV+jrTxOMpKpn+J58wmE
nqkH2c6/Hp5F09sSbGb4+pgeVD2w5oVbtRVEir5o72zZChC0zR1rVUXZGm0pu+Ce
BkG797UM9ifHO9MU63CvAAODTCHfiDwGQvHM7gtDKn1miO36gP1sXT4I/KWmOwAq
xs3yVWP1HGLODIj6H18VfYxh9gJuB27p1LNinW0uiYr1RmgohpynXuXS7oJcDajq
5SpHjApfWvpMc71LXh/0IwhwGdtDjEJIUPndY7Upm+uWcmKzQg0yFVqwPO4qg+AO
hAChhO/pRSk5qjwlO4ijuPQilY24S8FdlxrX5GGvKFH54iLOSyuAVz1POK1cMVEM
iOsQJUyMAVCYsRSk41u6abJvtft49yRqZcQVVWLY1eOiBiKmrSHThxCggil25eLL
cTrK1G5sVlIOvS+0dk0RwmDlBU2mYsJwa/2Dg5enqPMzq2DUZcj7SHeXqhXdO6W8
GqWWjsqdPlh3mskjZUzc3d9yxodUCCLccAJ/eGE7GKxttBrulbrm78EsyZ2bA36y
g7PIUxFVxJN+O4olEExWmb5NVqu4lr/tyJajwYe4rLA9qJTksnrbibjxNzEUXKfD
D6hPl6fA4MqfcmyhHjsMaenkCNhGrjAVJrR5DK3gkXW8usZCeshCin8ZtCZBcR34
+Us+cwlQIdqy1RbbiNhSilRsy1s9Qz3TMHltm/SfKuAWHlBr0871W8UwMyudviyi
WSYAl3rRcrSbB2bdoyn/niUDAIVSxtLM9uWwJQpPOF8xtEonWPA4LCdKMEttFabK
bekOZhd+sB2Tt4AoZO6hxUdc7LgYJP1sqJ8adZypVBUdJ1Z+1o6h6+vzzGAiIltp
tIEQWmMycfJWUTct0oCKANOeHMK8ZUuU4uVnbNrIBm7xL0tChjym5xCkd2EeXvnu
1ESrLCQqd4fsA6wDABBV7rO95mRyrLRfT/YBVg6Yeiw8l574zMwaAMrOPtqb1Kjc
g2hEN5rmh2kvmM1E8A+bd5Qk5/1wJ2/dI1avUeWVsMi96NEwIKa/Ir+ofiqYsBT1
q+5sdzXdMHoiW+G5yiIY0kr6HPq2/gPLRQvwlvMf+t0vhQKmXE5lJM/j5AASeUVi
5q7H00FdZ7REbD0PlNDAGKqiB6qEPlRF+Z0zXX7ZWL5ibc2MZZZxFdKImRCRu/cL
sniEpS3wvvb8q1iWrfpi6AvkrHPszjWYtuIygn65T7C8Bdzo6LauJ3bjFW+6+BRQ
s6yJcssv+qBXzyE6pi+SE1CWXooBGiPhcr7RP+nbv60ERRhiwBeZGh3pkHPfxp3C
Cmt/Dr6b9BIarAdXrXTrvIucBehy9PO/pA1n65iFMBwqHD2n7XXB4zMmAgHnEYkV
Q95SJYBD556g9j/FxC+alnAWln0ysYd5umiKZrmqYlHYlOr0saI8AVQ1bECUZObI
SFwTmSbBXJTXw3sidtMfBQ9G7HUR9Hji5nmKSVka1p3E/8SVfVhyLXi0JhAaCtJv
iqfsXMRHoQdsIB0NttbzqKTKFKN/ce+thsoautfAUMxLfkGWVQxytlOR/msLjjpR
S/WceIPDnCcPppQPaT5HTtu8XSu147Bvj+aMSPQoaiKvaFANDNRa5eCZxSywiwcn
OTKYkCT17ol34Iw4ih/FncKFK1LoNnABu8KDiYJKqOyyer7Dc993UXTsBRMtJTUa
FQ6w60IXNftjeRMwHKcpM3rE3shOm8pjF1F0Y9+ubS5O6c2iFTcu9dyDL74h/dM4
n+EpJa5TDgcJk/NDompY/dBeTKkHCMusH2Tqf0G+eh7URWJ8jPZG+VdZzR43w5P9
1sNNEQou9u7cZBX1FneWBLiFl/ekJlvwbY5rdbz9nm5vbhKt5wQJrozKZ3/6UsPb
LSabmsmfehEqRsvpjSuPTR5KaP3KOmA+sJkBWSLly8IC3h/kYWrErcQZtbHwGmrK
J9z7c1eETs+rcGxaQ/9x+gNiQmSc56ycfMgdFhYkEGpOcOLV2iGEV1KiujDYkUfu
jWg5sixptN3R/o4qhP45g04o+w72ceULgLvpHvyzdlTqZ0mb5QHIKmJr+VUDvAfb
6fqNDrnAFQmbowxKLpoRIFeR2XTTL7hiWF7vVWhwWQT0WsephLsp6NIgC11AR844
9dNLq8FY0Rg/y2zXZ3+AliqhtwWyRyVwIa3o9scsXmUBqYIRD/99BBCAJS1U/gT4
Gcg9Un5SquxSDe6v1ygWqE5k9yyn6jWviPlexwlxDQ/D9ar1NflGv9SsDiPRruvx
qcmZ5w2uLiymCxrXgtQL+pkPEHB2gZQiCfe3Ya4iBdBX0xc35VMjTGJkS1Gz3UxD
N4dPQTupVCs8XYsIJ4lU5PXzy7OBZmlmcUTGEkL1IWrTuZhdW2HPdUY2PnxtjFs2
Fev+zsrtDIUlm2h6+HSbEqwpyAQKHtvgsczM/4xaLOGBLaAJNgDmQfmuS4hNnGlJ
ZiWnRQ9eRLsC0hxdzQ5h/q/Iv315lALpD5VIOY5PK8HK5bEMZiv9FADaZTvO88+K
jZwdlMMZGUQ80Iqgcqu/a2bcUwhFiYl/Ag668/f5yvvLhvMYNRtFrF/GdHxPD4Nw
Sz7c2swu1ONtDakpy0jYenk1yyaCl+TgmMDl6iB4qEaaqRmBGVesVwIMPhy8Nz5k
1R/HQ0KzY10UwlOjYSf31qxJQJcTAafGrRyDhPHQbaXa6uKLNBFXDKWighqs54xt
0O2NlHKiG+ztYsoopp7WWOX7qH8c1ykUJIInv6OraA/sGTYFEPSJwqhuLReFt+UI
lyAV9OFbQsc5GWm6baOWqdyAu7BVB5oaVBwveUwZZoc/kDlYFhKJl+Xiwv/qyPkW
JpJAGPD2C7W2Dix8XZX+wML/KFLMOX9qEC+1VQq0dkN9d/fdx4MOdXoY7X1diZ7o
zzKClS9xoyTQUTE/ORPiMXa/i3Koh9hx1sqpA9gfEK9SHDYc8afn2xFuw0shCZhU
c0+B01dE/sDOCA1t3y1rpWHv+1Cf7l++nkzrYSywcAZe4gxrKnwR7Sq68uocMu9W
9ztjCULsP8pity5tm1NHqIF2HjauWAFmbNCadrrWjmudz0YgHvES7ocALR+A0OMI
y1aUTa93qV0EgVLMF8TWD3laPcSmiDmSs8KlJIHLmkv+WUtNTVB93DHYmkePtY1w
jwrgDVYD05GpvjViW1UmnwYlvYCXbQTp9cEPRSdjxRuF0zHDgr6LYrvFaiLlhjYS
H35pT9+qlwfECMSGnMMBDb4qKHpHF8PrfhnAVVUwoHwc/o1SH4Lv3H2KutfMyPH+
c7wHlbUed1kiSH5pLbndXspDeftttoipqt0m9+pUMSSmUXm6xsi7NaDNuHHOfW0U
LuHubQqrPdCO4q3Vgxxpc8Q7eGY3jLKztageOniQxoOqO0bevoOPyO/PLPD1B/Oh
Shh/+7NgoUtJKGRwRGC7r2ZCTc6MXg2cLC8KONKc4CgHfQoEve7cCDMCw0oIhETM
F5PCDTsnOOa4Vfn9JDZVkJxcZGBwu0ySPcveSvbfet26NIOgrsd8F2xn3SeeOgiI
DpUhVfZRtmqzLRdOl4RV03ZoW6rVjH0jggbZAFDOm1LfPSSmJvBIRZzVvpTiIo/8
uSAewXtI6n6jlOcRjKVsr44145py+55ck8FWyNWiIXTUvCOPG1LQyByE7MzNXj+c
boOYERTmJpg1UTFihw/YoNXxodjT76g5qTnPkkcRgQS86c16wghfcmKXH4TwoBgN
GaZG/5SdXAkaYXUFOa6ZxEcAigMz7bYMmBya4tyre/2E9u5Pl8zOZR0MNXDz3W9k
nh9Zer9MyKHu2pGYGzhkeDnZxstc5qnvhpVVfs8qO+bc2YRbjQqQt8RyMDo9//Df
n8zCBvp5FV3uvfPreO4v0i6a2NxjrRNUNDxB/N9hRR/Wx5dqQLj80sgNQApEWPc8
8DEEGiQs2Ubm3J22gpc9F3Ipsfey8E4O0uIb8EcrnlrOXIvD4QHw8utVL/JRcDJT
ZsZgqMY6JVFl8dcolukoSFmT4NSrH1uSwPsFGxvZEE7a2uFpnvCm2sWGLwLRP6hq
z85XtDgdGDFrghrgNoIuTyNjlLL7+8HWRYhptna4Az//SSBWy4DcKZkUKszMioFv
aVzge0xsrMwti4S/PUzyZAFuC4XJz3+BnW2ik3/h8lj4LKhO/UXbfLQ9FmGf7ifA
8qeTfc8JVLp2QS6CmxEWBPiHiSDvndDkYAfuVRzSFeXY3AXfMXESjoASp9aqZRMJ
S7P84gAXkDN591VYqgdV/bjBSZXlmOal+ITLFGrvL0nt4Mw+ZomgPvYX7IhFSh9b
3wto9whiQqRoI3J5kLxqIumEuNej+bw64fIo2c2Yf3O6XGrE2D7Cs7S1ruue0Xq/
W9M0zZnEjusLM27t5YZ1w+y7dAbZg4t6guRj7rteEQG5mZM5x7abCXnCLg2ZPssV
PT2L8feO5d90zginyA6TIK7RU8AVTuLoe7pLkObrkVQfsa5u6VcPkaAfd4vzJ0ak
XU/lOJfJM41cCwpzCjTudCZ1lb3qQ9qVlfKdph0ROshgn4+/CiZdUzjM8fcigec9
nP0uH6FYFNuk+Hvl5BmFRdiDOJG76od1MfWGUNtoYIzMIi9bPV7SXzYzA4Pjbm7R
Y1XvzkO1rf0u2Lw68eSqa1aprA08FOKTjlpF424Oo7cK8+S+vD6NMHK60KQAzr8z
g7wTgkhp1J+S0nKCd02uHIVbd4RVQ/Eitv6LfqR3jampTBnD1Xl0sVTrCvV30kUT
4xm2r3NwfxJ/Vu+I8Aaee/6qTRaxpWfhn6cooxFgBWRoaGNcUderOu/BYWYi0Wm+
U2aaef3dnKQ529KSJDHgEjETiuDpBhbp4axI3Mr9+bmnAs6Az2zBT5noThmi7czC
aUpFuZqQ0EUbQuLJ4hWkGDnMadgBy/kCVtzpEGmm0RuGIwn3OCyvRli+umIInBMl
iCMaybTLrAezoykNknIitp2zE2At3WpNrD/hMl1Sp4b6DisN70SucqQd9SjOAh/z
BsfTwE66iOnu27AEFou+AN9sRRKMuU5UlyF6Apac83apAMds+koz4Xd9bexIQl63
NzmYVIDEMQ3/afZjcphKqQZaTwXo1Db4aejmDbSNH9LkTF3G4fbKTukz9nRIVRwP
BMNbnOi1l/7VVEpdBHWnv2izQZS4WJhlsqeSYVeLMpmOGWruJZWFT4ejqfB7qbd6
slfanwGdNdQJBLFAj7/De79A9eTlcI9aQ0wML0C7f0UwULokr/I0Pl+BBTwPOnHJ
WR+ROoTdnGt8np3gKbF2dFwJZNKe+QdbK+cerVDBhm6+9R+X2DQySuEVE8wXnVl2
UKSVzQI8uVBYU3OsYCqGYPZUUNCGqw94/9ttOx8WoxM3rwUlBmnR5irQ/dKogzr7
hdx2EZEKd6j7hwycpVF8jAMj/jVANm09kH/PtQyWPeX56S4fsOSY/rKKCesNIQK/
IHK9U0IaTGshdY1rRxJVOKSM5uBPoh8VxxZuD131z3Jgb+OQ0EdPCx2WuvmBc3Sa
cVd1TMyYIif8nFPMzihwXWbQBXYwwy2InP3e3AtqsXsAhzJb8hxhm2ZWdPtlUitV
gvnYx+GVeBC3ftWPGT45cQcMw5o61KtHWxKCnS8/dhgi2+gPbSlUG/HYgRVFbLy0
sTlZnzx8rz4PAIIZrIFr2HkV3QT2H9DFjt8ZiPvIxzIgWOwPE89qxR8mS6fvctme
p74CMl6JQVcH9kfCH3T0fpEnXCLjtucnG+FqkMCoOwJurWnJ74VkNJ9EafBl8t0u
v+f2aZ+Ifvs3vc7nV3q0tJUZZN323T+XhRQPDoU+XBKdaINLnIrnavSYPrwm5QzY
216pwbNcSzJzTX36QBHom/bSnIg0WPBN1o7XnWp8e4aQ5cf4di2wvx2D4tLnzwYs
wg4gCro2XP3CSTT86sz4JFUI2lZ6QeZo87YgbNIzBBG1hM5JobmJ6imXYYYxv27F
P6kvLiSRB00B1IQennczIP9OLPdxbFs4z94T81GUaKz0WHqfT9ja2aMUZNikkv/O
dMKGDF5F6d32Pg/FZq1r2b9VBC4DEov2ePpLFuUIb6oFahyFxy2lP7Sqa/aznHPL
NR+aa9XCeaEnJZJJdSMeSa4pZ6FJzILG7gWx2m5NUAtVLGVy7gEdsF8jT5b5boWV
sHv9AdixB3ZNbe3N31h7CpTnQdNnAo2NqUcC322h/ZnFqtRiJuJFLbv0EmV0x5CT
8Gh9yfQ2Lym6C0s6fSySeefDFusZz5LKCuuXKSd39kr158/59k+D/AOZrlxl6x8Y
qyYBgfkiX4dRqLLm3xXWKtal6auEpP+ixso5LulKcJofc0yYu9HWcEgebqDf9oac
jU0KWvc+ntN6rG/eEzlA26cbDRmB0d7XoqCC9EAUBBv1QHSlG+odigdgI2MDO8jF
TXFuQVJ+BpKihg0F60kYOGK+nldrjZEN+qYmMrRcJVSdrp3FnfUa3ouvUDQJiLA+
Tf9DKl6iFqixE+Ez6bQJgpjS6/C5FWfnFkuJ9dcAHf8A5L/AH4mfmnJP7v2ixEVL
BPgIMqCRXy8oI2lUzicnq90aIhVp8Xsps6perGvxcB8gGml3SFfLZZRiWEn+FUsv
FC7FC4k8BqucL1GichI62cNpUSCdWy47fKO3kF9wa3MaSA3USGegQOAomgB6n4cV
rWcxbGZ2JTltcw14YMK+n3qio8X5MhUwrt9HtpHMWXJgyBeQhAh4iDrRlCSFAOSe
hqszvzfu/EB0EQh0W0aEUFcWzf/KkfsWx+Uhlp1hae5q40ie5Hswo/jTMtIirSyV
B4hczXQcege3McrQqXizSyxMymx4WLI6jg4ef5Khp5IO5JGUgSkkG2X344636JRU
XzXMNPNpeIBUzrbeqUUTDfJv9g7fHkTaxJS4smWdjfKhFlBRnTBwDpgyIaeKWyOM
tyTHkFq5/FDkfSG2gHQhZYXMQlgUcxqEZvbpHOuBqLH0XrBQQ4gjNuQbo7oBIUWo
ia4oJYn6D/70l2wqnb2rgXUOFtzep1u2Ixgly2XEk4ESAo0aWhDb6bmHWFib6k44
QKVuggVO+mpvYTUdoJ1a2pb+MOiE8Rviesa3oj7032CD9ujYloUeZjV24XCpvtSa
4ZGvRAItAl9dwz7/s/1tTM4tNmHTNj5YZORTEgGhsqITzvfrbiRTb6AXN8YX9liK
lXQgYOsoYizfHfz2aKSFHW0DdsxgDSPOMZrO7D5jvSdinu88Ho0W9Hn6HaA+uXGx
8Cfm2+2XVcve9D3VNuHlOvyVY747aI4dZ1sy0S7FAp+FUroPdgR2bN0zfDSigrq9
ox9Ghw0fRbZ2ywZQqGS76wFo8xgjLHnRat5d+//Umlq32/PL1K2PPrMdg+qpI4bl
cikNKxrcmKoU3YeT39X6SRkFeDH5sYZUTa6VN/7DWu9AtMDWzHD+Eypx7b5iloBw
NPFjSx2zMP+3KD0ShcPskuzycmNwaiZ0pLdt4VkwnmaJX4OYrorxgJ49BkCcvGob
JuPDZbN94wYDiijHMA7iH40KtLz/LkYJMWJwKehNZ6usSnaze6Vo/ovvhQnclud9
mDYbH/uUFYsgJR5U5xZg7VMJ7ADmpT8SbzWst+VQkPRUwcbj8F28keHf1b0zKedR
7OE8CNP42b6rob448OfFMzznfWVTAwo4/5049hq89R44dwYs2c5isoPTAM+Y6kxf
bcQE3ah2KpI2IFrHOT6/orGKoOjHnRloovbaeY8agcLzaFxTUu6DATGTl5+k3W3A
yZEHeJlghStKcSzffp/0ek0V8ZqYLcf+fzK8CsRzIrS3fpmspdVwQ5GsEYWlO0F5
WTd4RpfwQgugDbYz73e2HseE0wmAPA2LUsBX4Enx3I7a0lmJQQbFDSYQHSk/N8NL
wVZuB0E8dEWUJtBzQBE9ENEaQxY+yXqGor+53FlThLtXPOy6/7s4Wx7AATSabxJr
ZicGz22AzhWxfZGcUtgujwvgpMwsOOOtZBOo369iO6Wqy/myC0o2OB9tJkodsExf
9DKPRL2KZ5a6TW87UkkF6kqUbfxS0j9o+7baJbbdw9jOIvh9+DkrmJ4oGlmiBq6r
G0h9WjrtgMZQu6M6cHDuRUZTc5TmoLDhvKrUmX4BIFeBe87kUvHBEc8j8p0vPRZO
5l6ZE9lOpVy4tYjyMgGc6bBeuQMSqsEMyKK7nmGQIMJDSUqg9uPID2RVz3nsSEqE
MKpfTYJpzkXp8B/2CKUcPCuxYFaPIh4PWhzXcab4RABMRHMo0WbFskHW86XGiCuF
n2wEkzQ2l+JzWbaEZXnMqlqpCTz0x5APh2f0LPgaN4dYZzWV/uDiCNQ90vLhCddI
fjBq/ni9QXp1oUbL+Fuqeo2ly5SwEO6/s3XeZoz3o/HUtoCbqGo6Yf/xeJ4p4JoO
gEXKN0WVrI0X01GCDe/2186ShPLAdFKdu/zAZjWkc6MKDJREhGGcdALLvxN5etOD
3ViHahYJ8ZdvzvCnhDYs60xug4jR0koOHJ6Eksg8XFrIryCKsKNI9TLG6p0IpKQl
LxBOaIxKifUR8DaXNfP604MLFtjRisha/NJIH+QF8AwJG7pPYgWoC1wwsI/HALFw
GRRjrml01AGulAXdfouW0g==
`protect END_PROTECTED
