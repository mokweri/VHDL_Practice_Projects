`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oj86f6qA33U1CsVapie5SNNeDPZA10HUOjI/A8YURSeJUD+fM32LuKyRxtftpf0X
5qjyTYt5f6ep+lqMNO3jsFWcJGhSaDUIwOxIdPJjaYmNZVrUWHm9Xgn23nglEdgI
dcF9yJ5oIWPBGwvb3fqfu1sqoushXLt+49aR1+ZxHDj22S4ke8P0V0N4/QOuaxjl
0YB8jMxWXkWt4WLZdlU9q+jXH3R/XcOk4r4UGUtUSmiFuV/K6Z3jbzCj69BqI6SD
nRTbqxtJtw2LIZo8badNran8dzFzsqXbauPPFrvRbxM4bnnrP0Pw4jjuDjUrDr7+
AHL/IETGnzH9C3gvUptQPeEzoYc8Xf7rQB6luV87T2GBUQ/xFruHvh9iqalbev3b
k8x5ChJ52TOfH319wfLa3SXQQcKRWlKwUWVDXSieevPRJmK1BbIo7mtzgKugrwnR
BdoV6UD5WmySXKHsHuXFM6ArLVPxIs8CEbrnS45tYexYXx8troRJp5RcsZMqVsOi
V56A9CMndqtRFCWaj/bpGBePc0qWd7kXL8HkTYoPSAlrGMzDVx18a9F9ZtOIObBC
P3HsRpahD8VvqwQdyG6eiAv65jnvc2LRlnxybVy8fXHQgahjDafhozz+D9+bnsEU
4LzSNQJGTbib1I0fhl2k/uj/XUFPJC+NlzidjB7eaDltJxHXxK+x+L7JXqTV6lZ0
i5yYHqpL3tibmEwd/KjzRXDlqaIPJU8vdY6FIdY2u2R6Hxb3e0Uvh+zAvTnoDrBI
PR9pEC9RXx0+NLWtxHNSTO9cgtFnmCbzvCS0ELPKxEvmh+OiegYqi8AwxIYAdqGa
vUkhPcmT05Bz8bF/eg02HeVY1Zk3xn2ikIkDWzQzHGq1iSsygtNudO7sufgjhb8c
N7qS+dnfqG3fFNhga5wFpUuc4W2XuJuAPGDVLKs2DzPiBB9Jv3RaLzORFTXoBB1f
gdU4nkrvBu0Pn6oR3+426ILOZ6i6Pl4ryBm1Mx64of0TlPwGRMIfe/9VQqU3V3h1
vrw5zlzY50wQDUJwLBarDWfjzv3Al51QfqdwBvU9pWrwvahom3DgUiQNU4j+y5YT
5NSNqYV4r4raZOakQ8RULqC8NL5T4Ca0IhKcRQgEKL8RElaLqKEfvdPyFeaZiPu2
uLt4+PU2md5YwYvNpI2CM2gYzfp8wpM7x12SsUezWq0lZLAZ9jT15RcVUNpyzr3k
JorTBV0ND4FEG7PKHh0FzUPQHlA2N5AfgfYsMqpUNtL6P3MmHqjf2cN1++9w0ndb
i9RqfZUHoTxmQ19sjaYKzoJtSDAQnVbqTao9kbcLEYbZ2Ov6yMlyZuqdxhqh1m0Q
3wfGqY/lVlbAZ9xsCwFVYo8+9gh44mxWhUajQdXgKqbUrtWHauhWmf+M4bJBaU00
qqWdJeY7bHthp+iss/L6dd/LwlQC9Cd6C3Pk7imWbyIitINkYGwPs7UergrjiYn/
uE8EPRYxqja/xQ7TXfQOvr0YA8pzMPmI7WU2ZHazeXKszz6WR1m7naeITah9rCe2
FbVGinZSjg7zRRWPZU4DO5Y7SSR+t3IzwmnVgf7KiyhfjCYiOkuTYS+bawD1+XEr
Wo/a+YYynAWyuFRoHZUGPjawl/7VPOD8z89BvlrRH60mfWkcuSIRG4WeVsMstRqW
6zG/6yUuMQlWct93R1DtebmQlx1tqhnc9p5gIkosTDljc1XwppzFLCmRrQY6busm
/h09o22toXUrg7g1sy++0mq01wDgASTyw8qCJiGuhlE8HiiWdZJsyDYyezANL72W
qIGar5/XF3w6P9gIJc0PYH7p+mlfioKvSPY67ZT2SP6XIVTsjGYAl7Ftx40PEhtr
Ri3W8shWlBVOrJd8uiJgFQRaQ331qH6afCIlcPDtINW0wJNhkkHp2UmaCAjphXST
gnsjty61070wLNO3IPOiErTRw/vc4K3gzaRxpzFVH5wgYXj9bs9tz/mBnvNcduWM
xIqcpR2pL8xJINxWm4yXkWmr2Rjl4bT5KiNV2K9UkdBz08DVzIp3pWBDx731lSVr
dKt70wNA0SakjrbwRkT1l0MWLeDMKGQByZLSDCaqsVk52Vnux3dvckJHp7hv+Ozg
6YiINUQiq+sHGHAYLPCWscZD5sDR+y+Yw3yP/L+cHcgh41/f/k7eN6RFEiLWO1iU
eOSSlrPd6CQGoNHDOUIP5C8L85AzlI2gPhjj7U0KJEgyaktrRPha8INkdn2awe6x
K3FG8ifCAbPMWAGgIMxD5kfpao5Y4iILdDL1spvAD6Bm48riTcS4OAbImY1Gm2IK
VVnDuTjHXX11knmlJb9HNwkOsUk+9QG4vX7LTdlyRZCAy3MWnHZBKoXyZF5qju+J
Id/hqT1KDlIA1Xews3yUfFikENExF69mfJzeKRVj/mw1/O6ws3tL1o4cyRaYzKDP
bGWrxfB81jG4VcfuTHHwUInQ1MAGmkrEGUFxlX2s4bPqJZWMSLKV8xg+90yI/P7b
5OvgU8hlYHHNmOZOH3mfD70Aqv2e6lEN09pm9ziPUnxnPPV29D/0aqV3YD9ek7qM
DS5URCnwx9S5I/t7AoYtzQZO3P5mfNBR2CLyqj57hpWAkWq2WyOBefTpbfXc1/Fh
HY2020tnms/e3IL2/RGUxlvuzQe5J3sbL4W02aOQ51rbogaeswxrC7xsR/HhMIvI
zuaozZnVxHjIEUwfeXjQAQ/GxDMsKsyAb13RcPe7qMDAPfEYdqiPLm7QIXrk5C0o
h/Od6rWGXHEzs+MrGfvI86ZoHb+cr+l86Rl77msN964JJsV2Hj09woT9sM3z4tAl
fZ3ZxV/WItMUwce59mKI2LB5e8504kBOYyPQT++fWdZmwyLY4WOZNEFwW9UcsFKO
zljJhGOIhlcEJasL7gEqTYTXrGyf9fHaFw3+AO//xEoPh2RevpRndAtvH6DLk5hl
KqJUhHjeVPieWg7NE0ghzkaeUiBW41ChN1RXUyFwSNlyvvDN5XNEemrB65KJXej6
VAAKbcMJ2Vg1tmxpOEhcWcp3fC1FolXrR4geeR8NXmBXQ0LOl+rUUnxg2PAxaXIX
AAykKq3moDj1lwGcvLxxhoH6dlVVPpuaVXJgawbabMcht7/H3ZtMtVIZAp+JGYsg
83hZPpPUKy8EcQKmIOMNk077v6RDq6aCpBYtLC2dlf/uIMR1Xb+VR7wpnYD449jC
RKo3ptqoXSGGiRwFCm2pE9NAEvb4ow+eaygxETvfJ/YPC1T9lNM1xbLCEzibFqX5
cc0lLx5GLAZ5EU6I5nVrqayvSjs7e9AqNjBzLhIoazqZ5ProyElbxpKWbgPNY9aB
OB5xFQlIweffrM97h2TV8AfchSMtc0/HO/fnjCW5DihQjiO5YHU74q4TkFyRrdrt
OIY2Z8fmt1TzKUMxSJKzLkesNjwN5mfmozeZ/G3SOEYJUT8/J6GZ8bmhrOViVRjU
96PlrEMG+pgX9MH0TNXE1FsfRit77lGCCI36q5BfbASGm1T/jB2Wmj+7WbnE4fT+
65xUz0JReL/UsbyZkhGh7uEBQ1VwqkmhooF4YbXcTWpKzgAm3nnXBhTgI7+jaGsi
irJsgqjrm6KmH4UiXPL/hNCaltDtf4w3/OxrDyG8S90o0h4/EOiUj48qcG5U74T7
u8qZiTi1KdKGS9msGYTN6zNCNBeY9l589PMVm98JB8MEUE5kqd99TCHQl9V0QpQG
7REeBJ1gxrRejxH3Oiur9QMRbny0RVhCxxQ52gWyqzAUD/nBxJ2xVGCR2ZLYu+SN
wIMAbbkFLrCszflXB+gAfPSRDlheHIYNHMi/NHpdo+nhw163B+DiGSQjQ+bbs2oe
ixQVshZO1qAjh3sxdsmfbOAQJiP2NiRW5VdCWFYVi7hwi/USg0nR8gcUNox+K04Y
PpLzFX34mgWXip2Qfa7BxLT4JirYZ5YJOHvGHqsMxVKcAinnJrPPW24FVXUWHc3E
PQs3u/Qu9iC5Lztv9N0yfLMRvoSga7JKK+YiNRkvmbvYKnKZGoC6y/fWMRDfa4ce
72LYU79sv41T9c16x+0TC9BPFtWKdtnZvmfuRN/io4h8pySR6zISmmwudz1uDSlr
sQ7+7IGcg+EnYBz+DD0PWZUpoAqT1l7wopjEWLUl2nlUuwOQWxzMI3Kh7j1AC/19
CbkBwE2DsKPKv/6RZYVlieSp20Kr/3P7XV7MFwrK4kpR+qZl7tJIfdyzFyuoXx2M
s+eP8yhOB6FW4hlD1y8ynyLDALYd2whob+c+ObQCk7EL6jXgbal9SbuoYOI1XbZP
PMmYtfXHDhDUStASKVH/8S0esJJlkOGubUsLUFRlff3jn/VkFo+Mp1Kp6OrXyiXQ
PAIFvprZ/rcNfYFYz2ebO+G5aGHeQNRSKdVQXYgqY7BmlAbMqOz9o9hR8oYRAIRI
er9/GoxkodCv4nazVILmUOu4DONkOSD9I14NppFptBN9FWH4qCEzdJgUusTroJmx
wrP7iXISlLY0OWuGHnpKU/Qad1YQ2JD7DxSuBM7Ey8WB27qmNMO7UPSnc5IPVw3I
Q6Sdl3NtpUwwPMjQtj0P9wV2b+Syq6q1omqRjO2mUJZKoV5sL+jI1z+tkbR7acbK
6ju14LQqOm99Utk0oV7Q+szoKdWlJDrYZEdcZlzKrn7wwLO74GeC+stsI5uQ2OQH
iBl5X7TSEx0SUvdU6aNKA4GfPiymi+xVflipd1wTVWA8SJcrlHsrfoJ6UqGNRgnX
5Q9wxRkKGa9PhXQe7IXaeYXgjAd1jxdH8QVJusAwW4W7LpAPhfCU8AIwY5cwq3CY
pTtnQ+af4laEEPeooGDJ1r+XijnJGcEFj+b5uqERkENAz/nqaqgDS0/YlMmbuS8y
+A8/Nr+uKY7LLYaJkZvtAfdLCRXgfLge+wwdky2UfydpZvypN817gv3qjiYsM8SG
RNoBx5u0vOkbNgpvghpINOjEWP6oy5JkdWruK6kVj/+KsNKITrci6DVMZVKCNNnO
AjyGyb8zdejhJ7vXeKto8IeqedpwXjf/lK9sr5bbC0SAW6t1XrWUAz4Oknt1pD11
oFbutDu/uGP9NVZPqs8ZKRyuPuDYxb/ZjwV3SAQ/N5JKhOfPZRTWHRV++kdt6Coi
ohyfLZoF8aZnhKDvmMtsq6qJsnmMNzpM0vNeiY79AMUyWlp9ZfnmGBTEjgbTQZSK
17ZKl3cBDR7+AkqhZr6p0Q90hDHosERmA5IQNoY5CIqQKd1xo6a45EumfzeThAKu
GpNakI6u9IjJMe0Zpc3q7DDVTZ7u2hDz79Bpp0xHVJktxXo6jhY5Rvs9BNF5zqzi
7t5UTfNsE8A65zr8NijEzNY/qnsdV4Zhn1RKt9zixjrYUxThuS57/JtCQ2ghksqb
3eC1T7IyjrkK62zZWg4EooM53KF00GZQOy5D8SMlSwfgc1Ps3wQTR844rKrWrZaR
Tz5hxggQibiBWZsysu6w2JpVcETZzGBwkVBwsAzcrhhzvS2zz48pPFKA6aXho6C1
plvrtEQBC9IwV/9/qpubeJbZjuSlid+89c17YWOHZ9E7XStkoEO3qrLqTWA6MZEJ
/bPYNpmUvborrNNgnVIWsbyg0Z5YGNSm51+wWQE4yE6aj2SHQ07QdAl8Vd2zaG2K
rLpYU7U9i4KlngUuOXdwJqXmZJzaYJhsSvt1ophMnN92XVOrPStW/jxTnHyFNbdJ
qw2XpezsU9fMss4tvEbs0NzSfakK0f1e2X/zHEsYoKYKFARrG4UyYWI9+D09LFHZ
4v71NshcSlC3qzGYn0x3x+iXyAwo2pj5UiWp5BDej8DhP+r/Bv9XfJFEc9ZEcMBP
qamjTy8OmyJ6RCrreWwSsOnLwXsj4P9Yh4k0XNDl/HXO+yTTDxYmSVs3hxYZSKSM
Nd5TQ+jCouy9H62xKGzpzv0522RvOJPLskCwfWw1yHg7CuBklh1+57Nbk+BGS1I0
B/ujRF72SJFPk1u9/FrtrNl26eKjwasBijOI35s9YbsSJYFLcK7opU4sieUC1gt4
TQUBJMznZpG4FaLhnfDpNi19wWzxA5Q56m4AQQWUGkpEZwQ+9XtiDT95qbSm0klw
y5qjrWCt9HMdKn9Tl18RYKMXX4N8gLFH3kxqUnfCUl4zeP49lIMRqiAbK3os8fP1
K4YWnwCi5H96GFMTC5KH20GrzS9SV0eVfmOk4JwiBpW82jC/bQfMD0WB+snnPUSS
fJ/z9ulaqVtcSoZpsKncuG51BPTxK24qycdIg/X6prI3w/HbThf6ZJ8DeXGYPmbO
PrEcN0DV6kclh8BDwXCcT4r+x3IYnpqdZOcEyt+vmO8g1kDxyuNvQB8ElYqYR0Hm
gLJWJ5iMZgcMv2SUSB4TbFN5FOlAFMe5H110Gg/z2JxxPv2I6np9kv/11D4JVm6x
oF6jLyVuL8R/opXjKpKdTkfYUhdNIj9mQJdKhsEx1pHUGYYJkvew385OMwIJFoCQ
My1P8dSL+/KC7odnpQWp8jmeMefuIBoSVpLrvC+7aFvyB0jNYXAxTTJ1oVD6laKK
RD94tMLWzdzOKNYNzET8ei890cFuxAHJzup1a5PqUQ912azMilIqLUApqA1SfRxq
5RAUmqYhoQoSzs7UKAcW6+pUdnx5Ir7So40pVbVqA9CX9E2ggUoeZ89PNpD9LIJf
oXX8d5idnUY13We8Kk4XXcWBw6KCIoAC+2phxY8qC0gwPlrPDCdpd9/g1kKy/S0S
gUGO5vw8Yr340d6PCOqHZg==
`protect END_PROTECTED
