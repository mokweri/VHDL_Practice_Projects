`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69tgDsraft/01U6OEoJZfazDJuMNyvQEy6KavSRYBbFnsYLmENOmgeuqxHu/85V9
hyJmEVZpqXKS5giBVjHDoLivVdjfc3lrVlnmXlXvMKH3nrHr9ZHCdmCh5Ug16Ork
8oQ/MGwvFGx5TEF15FQkMXUQ/IMAunr1jOhkbUSWwCHMMkswEAgOm3VkjBtHAKja
vYYtggLabVQ5PE8KmRn7hHdLpuAQea1EvYKnreUCUnND56TVyzjGsmMWaLH4Hs6a
dkIZQQ5dFmG5dDPNtOGRqIGv5bKkryeti9vkVmeV7jZ+tBWxrXMbNS6Nj/PDaOmu
9TihqsNTUXMQTBJEmFmPAp5I8N0zsmXIe7MdaGjnsVkavQeX6VxSgDpcmzymibus
PNGWEstLOLhvXDPvupJq04aAT1bactwHiQH8xiEHyX/idXddu6OZ/Jspl6lnB1kX
XHVfbJxygrrJvxE2HEdLiau9vMYB0e28aWMOsUUUNqcW6ValhCVgqRjlMQ9fFNJz
gFt6DZqPkqCjINIYdWe6hMyN3lWVOnX/IjLp/Pu5Pcb5E1kMWjLLfyVcnmIjmh2y
VD6a/Z58iQzcN0wmoiV8GcZgfjuRIKLinhYhq7OwMLYXOAkdJN/xnkhvXmTRZeYz
z1X4rUqwJA+ZXHoB7ndErDEpeYkf1n1dkwrfJOgVulfQXBkIAjivrwKVTfcrll3L
GtuyvONmEPdVXbZ1TVQZMrxnQs9V1ZPnOBSdXb1FMtnBIiW7JqkmlndmvazOdQmZ
lYMm+M6h3h59aL29OTSfgIPrL++JHNbWBcGGwLBlB7ZXPUwsQDeIfTlaLPmWRzNI
/GrH5WervEX1KE7xxm4onvSs0o58pHMzcyd09dg3Ftk5lfqB7MIMck+tTs6QUszm
2Mt7Hq4ahxBMAAhaw1zSkf6uZnz/dq8GjTyGK4HFI1DB1PVxmZF1PXjM0XN9Mt7Q
oEiLLQij541rQKHup55Y7EuIwUdz8oP+p5Vh0njgp2BA7BXWWoJ7uFI4HY8z8wrI
/B8D2MXK421xalvW3/GBm81nzKhd+bdenSVq5WdE15L49N3W3mAs9uR24I77xjkS
W2eV2M5nDir+LjhMEsmtPZJvCkHF79B5nuHw0zt/iS7JLikoBMRn3TTYmRgAknUC
TplvDEQ38KH+R4dbn7/db0HVAn3dJI9a91JVmIFK557Yjv+LnslMx0DXLTNFpvS/
ubwfWAjoh9TGwiC+jsG5Lxza7Qz1fuV/nlksvnUt0yqfErfqTowd9ArbJVfdai1y
3CULmHYL7TLsnziS40f7YF8wvNCIkSOhlPRrsb2Z7e/qCJRht52MOnS9YHf4mZQm
XawPxEAMZ5dSnoBjl33FkTzSZjajn2WD2G93U3t/KVp0y8Uq5n96chAJhVxptim3
Tb8NRBCmw01JpN92WY3TXQsPx3OfbQP3q5E8X7Tl8pFFwQB8gePRanYJIlelooGW
PHF4ttQPtWI6ZNOYcLUy3PFvhqk1YdW76NxE115DbsuIc0SkrXKmAUN6FekruvdY
HpH/icitBTkX+/qwVaevWB8jP0NoYt1vgHc1YMlZFhJKVkvQ8FvX/C9EQQHDeQFs
i/VvPhFcoipEj77qmWh+XS4R9jv1aG0CQo1NF8SzuiW1VRIV1sVN9t5SLtBoSN2W
MQxEzxBlcaTbu4hS5kRYAeiYn0gVwkvk/yxD/2fZNB4q+KDwEU0fkqconbZia1YP
s9DFNPUMHTUBp3bH/+a0m7eNquqxqlLb+N4iGGtNOS8x1F1G6xzBCx1C7Ng4WpAz
u9UyER/Lj1lV5Lb4k7wJAFH7vCQdc16az4TeCXFD5TxZAnF6y5Gtpyj6K9Tn1fSp
FlfdbJ3g2E1lygjn1xuFioi4dwaJJS8POgI9SJ/TXCczWLeX9IIm1XwZjq9rlySp
ruFgIJQVWWS3rYhTD9K+alehHON6xqnj3fw2rEOvirMpc1CtGPb4f2LLk0pqClHR
XfqhSTIGJsASmx1aOynJ6PYa5KicRObPTBfRpbBo1OprRMvzcaWx79F6MC6JcZBr
MKlq49UUfh6W69c+d3LmQ4Gnq49CqkDd3uAeDGiSNcaZFQJ2eQnDX6rxn3MHPefr
U1NPSJs2lX+AVBQj4w0g0Zh8Kj66WOokXXbHbkKFFzgxcDoP6DI9OET2zAdGd48Z
DtNqERZ/DiYpcKKNo6xs41+xDWwWzgbtB/VIon4gtugdgNC2RwvyErMuEhkp5ufP
FT8GPFKqp7Qjx3zRmAWX2ambjcdao6FchEz2jaetSwo2HlvCjpKxRlnREZu/dfd0
6Wj/EqKGBR5k2eLdvnRFLPKKqnWsaCvOJ+XUkaTMa7kHX1GqX1NFTKeD73b/qrSQ
x3YLlUtvNg31zRM5IlwsbI+fzXAlXRh+ivOU7v2aNlKAPBO4VOHauSafC7VXRaZf
BnFiC6LvORSoqSzh5sFSt51RbgvpXa4piCC6m7QILaDdUB5fv0k3C3OafcBRokyK
wxYZN4g5LIVCm+P+d0b2uhtFGzpBC9fBIY55cVRDouEIAyYl7imtJ+/gbVMJuIzv
YZlHL7Rda0HQj4UeFQooo1N6dwiZxx4d4IuPj2SxxUbua+5bWtUbyciLm1f1xSWs
cx7kbVtI2IDZYU+/ZQhNkJKnJDtyLUhSX/N03aF57nlJM3ACsYeT8PYj75Yvki9Y
0dj7QXdpfiVfspcTY/OwhvXcPmrfn7+wGhsiZulzgLduyaZA6PrbvnAvCBEkPsVa
x2UJQBxVB396gljMA3jwml5jANcdI5NX2bR0GXr67p8PrZd0K1O9FesWAooSj+2b
C36tfwD+hEi4x3Tzw0el5Mcy/sWKC0JU0ekL972CBOA4l9/mPKwPkUSbREkJu/K0
tBeZamVMFH+6kzInq0Gw1R6bvd75vJXicBYwhwtRgsMaic09gQA7MYvwhoFcOrmT
PCAw89XZh9ejbh5QEN66l2nCPfBgXDK/bjfbAcvq2tE7Pu0+EIYw9Q4qjRINEsO3
ZNi2q7Paf4+PCQo/faXYk48T8p3QlNFTaHISVI2lw/oAK6MWOuJq8pW/xd4Vptgs
+mxm/sYbSebBZHOON3T4zjK39VRwmYni80MfhCA6Y5hzRfZPYr4wgsTxaMWBcIYV
8Up0OcPqodgy8Z89kxw4v/w0AR9NqhctnZjKxNu8Qm/WZVQlQ3R4j/gQg3SF6ThM
I3GJRdxLPvyXdcNTdSGFoB2ucOk6lMMAp7YfxQChg5gY4O/mMAfnJWlQ2YXDuQaF
+EqfMEhVN66R8TPwhZ8zOoPC1boJ627tluiUKKoJkNg+KiZd8Kls5/7BVLF4PuIB
Juc4N2o3wLo+CWrrglwyTzNArTccVeaJt+rle7CEUfW3jMwSQofznRNOKKSuC0BH
qYSRD1Sz8EClpCX61Mo4Mqv/OGNt8GvIV6HXphyt+JGVGu89Ohcc9B7Ssff+x3FK
KDUMQRxuDh1Yi5PRmmSRJInGcmzvxx9VeJD/tnodaY6fLV85nJhqeZIubPWJjlfm
ZKyK+QSlcz8C6ccgcWQjS1y7eOWw6Q+YwBqUO6sv3dSix4F8Bkl8AhXUx0bfOpUw
iGSuyfRxOCXVHSuctq+ktdXf7k1us30OmPopd6uwOa6UWuSUFOuCn2d4tPrQfJDr
9EfhhOhyWg0zi51EZNqeZhSQvtWtD1UGWfF2gySQtZ0dC+GADkbvoq32BVSi0QUC
biCZ8+ekgnNzrch055/XaZX7tFPsbohFrYBSgPnlCJ0yprSXmaS1/1Ezy/h6BFiu
cclS1s8GCl5Ic5Oxtshc+j1ZPHVaWK+ObgduceCcKvaSGNU9fCMc4unx4I1EGzFy
pFJJ6gxC+IdjCMoVmY/KQTXWq7Eq0Ry4uejICb6460MnkF24jnJzFrdrAVL8s+ES
DWto4c9hFOtJ53rze8xHsHbg8LeQ6Kqu9nnMK+SY0NwSfVY7TUdsZcmdh9d6FnWW
XIbRmJIK1TWPv/O2w4FtLcXIVitIbdaKhj4HkhX1+8j8U3QMKAeMBWWPVX1Fx1PV
8aAYLvo+HrfQ2pv1c2+Ovlq1PpdEnQT+Y/GcIWw2P2pRMUzotEMAvmiOIvbKLHIX
YoFcUvYcYs2SA971YHw1/OUYC2X7l3HgZzdHSYakYPsvDZjjlPz2vAzaN3Zz7ZHB
hlgFcshJbEMUFiLtIMIUhFr38HHfqnJDeIPGW/Q6WBloms+XT099+HCnlcw/IvkL
RSOYuhNFCGfq19lSxxQZmOV2LLZTahW+ebf6533crN4ICwDAEOBeAFmw8ge/Shad
B7LKqG9R+r1TSe6yrUknQKzvPndcP3XpSdTBshKfSleRMPTT/1L99Le7cFlLuN05
3vgsiNIQ9SJek2iZQmYba6E2eSg7ykcwuqRZr0/sSwwTKR4JINuqxxWqzL51BFAX
l5NSlvfXS110jqJCurxD8plVAGI9G+ZmLng9vMict067AG6o//0UDHIDUz9DGtzL
5nEUUkkBF+Nxh5jLU31//L+85c9mB1Lm78zZeTSNqz3833jee67ZMVSNa2+UcJZ5
5J42jwMIfR+G6eIg2BHh75PWHBxL4+9PmStxetJaPkO6MoNb36zhSOS5rQgrohRU
DK8qc2uIhjZ1qCh8QywAHOQrra5sk+3QxaM51FzjNMYHHtFg3+08mXA3AxTAcVb5
7sPwh7z/ReG/MfxS9L2Pe7TDfeFRBfAtU9TZ5k7LIjjsUXzPX9JrVNZKDi7EdyIs
aNfbk30jFawaZSd2Rca7DKuEjBvrBd2suHKQ6+Nb3+BWxmESTPdhgd5C+/L0J8zn
1v1tBNwveWgnww+uNXRV+6SG93wn15wvfVZZm34WRMHumt7cEA5+MlqrKBnLoemT
jW+h8tFTeWDLl0JF7LA7H2JaTJnaoNGKNX08fF5Tgs03VaYJHDYiyyu0ikvi2dRX
Ev3Kj+BHe6gW5t2gXf+IQ27phH4f+8+c3+DliMAaLUL6FMxkhAk+P0vlA7mSKffJ
jweTXYWzKdQQVl4RLh41STwLeOVzOCE9pS/P22imCoSQ7cJgcFce0PstVjXfeicd
+hTQyOB1iObFqMrPQxhVVw==
`protect END_PROTECTED
