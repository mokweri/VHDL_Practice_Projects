`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWlfySaCefB6ZlwnqUN/iNdUMHMB9MoOUL+UefV95q3bLLlDcOz3gGVw2RFdYFwB
rPFnXX30FIZJsa389KalndNHDCgvxKDbhMWo0ag0V1hxildeH2XNHgrYVfRuXXJA
mWzpWs0bNoNz/xWVHAdGV9NKva7dNNEHUocgrL4/9jZNfY6vxKRrtV0I4293fcOM
1juOCu8tbEWdWDvbuQIWXqo05hM2WgTzI4LOWhBPRmHxmAMX6O/vIG6eEk7PY9ZN
5rP8iwfJD5EXmP0OipKb9Pf6/oES7MidGXnQGLnw+xBtq92MdLYzz9qXsiJjwY65
RD2Y5UGhTUwzkdXo0D6Vc7x77pytWrlZ+A5UANHaNDQuE3o1cW93MVXv8DdIkkWD
X4iVu0JuotAyLBslng/VTtzGdKQvNoHsAo7kDwOI8fqBOw3LxpU4oru3jez0v6lR
4ZMnIR9Eo/2hVIUvnQlFTOvKFZp/6GN/MVXVKvsIk4LByLACbW/t55A2nzYthOmd
DGXehoiKlhYLAAsH5puCDn8eANf0IZnDYe7seEfauFMTQhRffRH+xFUk18jnZ+QK
4AMQg9lHpQYtu0AEhOKaQIWjd51dSqQulXAIxTImTzX1lZm7M/IJOHbg/fhHkr/y
G2m2R92UKYsBrMhHLuF2aGSUue3BX2OQ7WdDNV2d3HPZlEMXF8mOn8+BjU/OJG7B
PCAezuOuJ8lP9ExojVS8iiN2Ye0BLhPFLil6bBCLz230Hsb1mkJNztML0+TEgshA
YZazRUsAgsdNluItQQCJ1Cd+/dAdR2fttKUWMavwIX+Z5+2QocVdTlAT0KkB+giG
2BNYWYp7yWyH91qYL9iVBahdESFqV4PCUp577u5WdK4=
`protect END_PROTECTED
