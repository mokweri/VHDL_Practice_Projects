`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afsWu8JoBHIXEG2QFm+6Rxj7VhAUAfzEe5I2aCe1TCVW9XEexcicEQX0dXT8SO9V
IONtq6BJRmWUHgni4p9XEkBOXUlyn3nBOx9qTD1K5hn5+tP00rj+mCX6d9ihg+ca
5PcfpEJwAcEpJlKY/h3nxO9OtEW2BDA9KwNP5QvHaRua/Mm9lKra/Gih8uOqgrY4
ocTTmGvERrOsRPLlIILiSxrWFpvrWJpPatk95VYBkeOVBL6vU6oP3HnDQDFcv5tP
ud4mSvEH8FJ78gtYH2vsqIHn2A00qOisA9dDIvluTe9v9fck9sk3lENt/QYMWv4p
W6pdiZZ61+SgribDgqI9oKFU/KfvUNstbf8mioQBRYL2Byj3qjsJaGHYjkdII679
3iUcARo9oB6Or0PwFPJ3HR4FE+keLaauW0G2ZA4J98fEqVCtyn90pPl91VjAZm02
W9bqqeUGdTxitztf23DYxhNgZ40DE3u4RmKHCTRMJ205962hT4EpPJAwFtv2Op12
uY9Wq2h7NMRoKTdTD6/y0pqqO4Y6C3+D6dDAthOun6Xk+HhhPoKERv99slWYAzEc
qH9LJoMbuKIdCN4QPQlRqRcOtgoEFugra7QEXRg1AcKdFhJ/zh0wmHQi0tzPATn4
iaRMyDBuv8Az7zqAU2YxFfx7y2e9Fh/ineC0UoTpIDgw0JKCpKOvGyPzaHRJtELE
ctQM4HLIuVMyQP/6moMNO8qs74mjWdIxcBLWtQml8tfY4Dc6Frlq3Anmnsdg+g9a
yeaK9QZSzk53vLtnOjKTryIgs89UOYg1I+eIyKvrxjsmIEF3LY2Ij1ByO+9Se9Fz
rmauN2nnS0HEdWtk+WoCToclALS/UKtIuhRl0FsF6kavF+Yu1PM6IzcgGS2f+Hdj
hWeaMNIdymojXNdvp5KNsbrygqp4j8/sT6RZoBTKVtzocWkgRuzZ7ae3JgaClq2+
TS1dDMhwc0GhmkeYa/CplAOB0oee8u7yr8o/9gSN85vsyDfWhw/5QEy0bVUDlfpQ
pf1nDknXZ/oPo33Ai/EPxKraT+w6zDvaLSxVtRWClS1fkXkI7OxWJQCugmAxV9wV
Dpf9WGFkgsCAQDARpEA8hyqKxC7JspjSLnkT2lBoWm8=
`protect END_PROTECTED
