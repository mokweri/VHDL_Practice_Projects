`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8FKlc62DP+qJNOzxBdA0kLfyBl3eQ6tqam9DcFLhMFy5RBSrzhCDDtBglaHo9lm
WtGW+ojf6c5gHkwfqXeQcQfi7P+O8eFcmLZvKZz7fbovlPG4VR7VnPuo4MPrVqEc
V9tY7sCqg3xrG4/Lv9lic+bvl65/P2euoa4QkwA3471o1WySU7q5vPr+dMDz8QVS
jLus1eQu2lJtETx/y/8Wrtrn1xR59eWYok4D1tET8wbLyPWQawsf2kbJw3Sm0rNv
ILQ2x5Ux7OZcQi1mdSSEUZ9RNz6NSwrc1iSUZ7dQJXh6wF1gte5aT89YbtHzsZ0Y
3N+hkXBfKJnBWJ13OMGOL/n9kVEn+CJ8ax8m659n1tX8BZLux3Q8No/a2XbV4VOm
qh84u5VKLv/iuc5coVy0ra9Fx+reeR7XB3MU5H6r/A7dLvxg6CN3PLirlnbfUqX6
1nRbGVtiG0ZisawHWuAM5CrV7ALKrawpH+TePLMmeS92kho0aso4qyjWgl7EKgei
6ytN91F/xchVGOWBV6/kCttHjSZfL4D1qBVcn++9UOU0TY/j6ZqB/210qBI41Am7
M2Kumua2tEmatYp3aonuw8H/3d7//2KG0ymRRx3J3E1QZtUvoKi2mP6VereVLm+D
hP4d8VtpMJOyBYfvLmROlOVCJXK/mq32Md/qNkdgw/eT38QdD8c6dtXjosqbfi8E
`protect END_PROTECTED
