`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YlhyValCr1/H1imvvvTHhmJJW8NG72beb2rTqY344tK99ae2GYAu1dOjvZLsrnEK
r5+y2gcNQ97RiTUfn47o6tAY2LYcMwG6waXtcGmhAIWotdwkq+cetkyiUl+MdVLc
zBfIfJqZWhA9YSL+8LhlEvWqCNuNU6f1dPCTmTm+5T/EkDRqtJgvQr2wolraL/mv
4qSM4s6h992vDUSrgx+cPMVM25qpEv589WkwaqWwMFc50clO2WE4QENi9onOxhJA
1veh1Cc5VdwikBqrttgYuJ8yNztbq7Rj3CT7+B8T3DPm44QZt+alJnpENoTh3t3N
h13iNXtJWrxu3/WMxSW8rl87MzVNvQd9IElwsUtWJNo3Ci7J/9T03q4utg5VaPRB
dXqZX7wEr3c96Olwx+HNtA2LjuY8Sl1zTrJZzFW6b8ODWRh8Ph84Y2oWBZvP1ADs
fejDcbKeRTDWPh6cpnCop6BGjebMu5J4PR8MUAty9AYm8rnV2sSU15qQ7PFyLc2v
cBpn9wi6uAmUd2AxO2NUebCZY3+hsZ52VjrCEzD0DoXFSAZIm/z9/O3sv4RZkT9g
UAEDQOoq0emNJpmPMMqFsLSv4ZpUswWGes+Lu7hx2fCGFisXDhXd9sQE+QOabvXH
bJsqgnz9+8iHgsP/m73WfpjjpnZl9b9kQZdy8wlrr5LZrkz6RlmUdR3IwKVb3Djo
/42iCM+pW0Qwc6hIBO12UexCaquJB77LwySxHdBhg0G9u8PsiHhlJReeibZzyYFM
57T4CuoAMN9njzovj7SXk8CXHRkb5UcN7DLCxUAY79suv7oTLgABOm5o/2yXdSDK
a7PrSuRUGXip9ihNNj/dgBr3/Rgy8cV/jlfOHTnHLLhkX1j/c5kUQei+uiPBBuZi
CMvW+xL5fSqexj6wztN9cBUsM5l48wDgfdwC9vd+ioZqcotCT9tBfuYVGiolG+SX
BJ4Zap/JT516B/eBAIdDg9BiUmzXwwEo7mR5v0LpPtOgjP/nCDkiG5M3W7hY9X4J
x9YnaZ0qyd4tL4kxnwsrebnKlvdhqIw/+/fzgeFeC8NH55Pb7h9l4QWqgocAvTbS
`protect END_PROTECTED
