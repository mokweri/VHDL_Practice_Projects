`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vStWLi9p3JlMP1oPnZNDOcYw/fFP+qrUPMb+C1VcHZgrkyNp82GbcGJqcjCr5b8
8uwMX9BCb1Gj8Rh/1CBlVkWtQo/soxQcokpqCndhwTddIiq3KUKIYlZv1gdEW+j0
jumTu/wL/WQCwMhYef7hpHAGTMYW+2/mwOJCtxK1EIvz3Pcjibed2fNJ+VfWIwRk
nrfLhrxbC17xWh712NWxo1k4Lkvj4SeIFmua2Yn79c28n2A1kk8l8sOu2Q6fKsXP
v2r4nD/cPsTM+8GkEb4JAtfn6ASO9NZfU9wTuHcEg0UURAyP5GBk1afidM1/08j8
ZALX2rV8RhZrSmzBR786GNN7VBCoYCASb6L7unDxBJt8Rf2+KdSshGkD7a2dNF4S
wCeOaMNVT6xbjk7lYtYRfcscGK4f/fijUykyiHFAvcIE95re4oYUx3aOYgWDT1sQ
1eAKYdkb54C+8em2u8ncFKgJ/P5w82xoDAwoi9wNpwvHLFtcdYr7hLlZaan0tWNw
sdH0iZGI8R4r5DzHLtbrExwsVSHf1AYxeOvJFx9cj0xC4MA2Sn8zdd7O8+5IF6Nv
XxR8ZBoBbztOgHU1NyfSmbD45CHsUJb3yp+fdIUagmzh5hTyYuHy/jG7fF1/MM/d
TNAmnIQb2DbRbE+GCTu8JNQOL9h4ZFCNSFc0q1U1+xmbQwVrlb4Q5uS+nbY+cHb7
6pFnvciEwMKSWq/hMMdQc0sEIhio0sEl17AyTBJsGiRayAQZ5P/7ok7kwTMK5QGd
wViUKcj9+oHP6qVxAjbV+6ZVsacXKQNRgb5eB3BulyllYRZS59khRTnzQZPEJi5f
LeKdwn7S39DUkVXZVaNSj1hwjE4NvtXNm4n3pfH+4iQ8i23l7svwM/TKVtZHt6l1
JeP0XlfJ5irej3lwsmu6EBDEswoFu4Gno1bL59nzpfoYJeoVVyP3Da88SgW3v0DE
e+nq6eqMPDSHiyovYNA5Nh0DpT948jC8d1/veY+0ylFyxkSGShwRml03yd4SASqX
ETN6TVMNFl6VBq/+CDF3kwdopyuLw0k1GDT23LKwjxdLv9Zl7JRx31LkJEvQ0MT5
B8viLUEJpNyYE8HJaKqujEfM06EoATVItSxx7Z9flGBGrAj8zmMJ1TQqHUMbeSmR
6x2WHr06W8wKRPdjIKq/UNVORgexkuVKCIF46HJk1Lm59yr2gXiqXivWvyJYsmw4
SGsp6h1VA0swOhtt6I5gmiWPBtRDVF2N3P49RueaaGs=
`protect END_PROTECTED
