`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAZlQ9lF2x0awOIWkiwM+dzlSe0JM1Fx5BqLiV4MNQrQOTt2svqiYTTvt02X+gF6
W/LtRf9MKGpetKf5C5mac/TP3m43DxrCEPvxW9VqFHl6b+FWCS03NiHyxe7R2e4Q
EpPYfvCO+sWw/abA92UOlNv7s6PWWKvRmAjuhUrc74iiL+ztjRpwgXoIyVcQzCG5
usQSdt1pseAjTwLDVqcTCAK69vNYlnwWxN60pUa3iwsW81jOBohgg6c1gztO0+ai
zeI/XpkWtEhpfPaMTohC86kysZevwHEWLD8v/HaBqpsenjvyvHYypMVz8uKJ/FZo
se2d/7Mo51+qmp74UbyPA3UrJiI9GOD/jwffjmBM9rzYRCdpV4+B6uBvXEuW8L6K
Fzd0yjOwoIyUL1/k8yNLqr3DtlVsyNkUTcgie4gk717cp5EwbnRZKw/EbwKWIXvM
yvwtm9X+IAelgQujcckklZpizC7zc9FtEWcpMeSbhrSSOxrPmrmVjV6aYKMvabbP
futBBbaOdp+0B0KhAZVeaNcJwC1dhU7Qvri0/4Ned/n3TkyPXDACEbPmlkp0WVa3
CGxTFpyqrrH3O5LmCrINjJdAOlelbq36TgiWU5Djy3ZTU3wQBbF+g3rKAiw0WfAA
hr0Rjs584Mlv30B9I8ehWcTOQeZSVunbYoHttKapPaUSz+lpHOOprS/RyVquV3wR
RrO1n5BePKmZ386j+PNhZV2MGjY3kF9etd4xO6tcfFZSvUStAK9yobOMloPcN4gm
iloMQI3W/t4onnnDslELmpZ/sJu/oro81MclOz+lGmnCzjmcb0xauyCxldT9DOy2
ZlnV7Tb3s/sOOwrze7rTHg==
`protect END_PROTECTED
