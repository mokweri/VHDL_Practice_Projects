`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ZO38yOacWUh5I+Px9rE76yRxPRj8ZlZxMoAt3euduM/LSSd4S2tB2OQf68a+wf/
kytkT8ABoP2cdgAdmx8WcraOlheurPcFj8nMi/fGQ8qa7bhW3pPwMq0qDZTImQcq
6FkRWhPsTmmnPDWrde1c+MFi5H57+yRmtG/wir6MxsGVfSc79VlbK0qpRkvdevzo
nIrWptWLCU7CgcNVelz2q+6t2VCjy6/PKql9IFibff1RA8tUGvmRYMFPGhoAbqzH
TXtWiViEVjpJ88QgQEJfKls7zzYuh5clZhz4QKh/92rdCvUX6JAGEd7KDoz5W4uk
TvPbUbpcW/PDTVXLZsuHB7iIPiia+U91An8Yy4gns01xHMxiu9J+ZX3MB4TJxZgB
ePGyexOAsyWpjYrdfCc4Mnje4Y/GJYAO0h+FQHAaNRny4ljZWd/biIhPMOEeIeFh
ZdPzFK5z4pg8bNkzWy/xcKyp3h+ff4+FPBAFZvrXKoxpgod+YozuO/1NdH87sPGv
I4Mv9w5NB3hjQ3P6grARnCfw0+A+d1vvFxqy0Q/jgZf6sxzW1f0MRoTMpkleXpVd
qdNBn8rr/au8OMup3Fm9rJmQUMh8l3mTRUJidfvJogEO46yxKnuhHtnQc+Ir6Mwr
dnr9WnnYLYWM9OU0dblPtoJStsT5pH5o/ScLviMOIY6u54C4MU6NIm8c4BatN9PS
HYkTOeWeU91aTXFMX4nDjX3nTTPnrjtssnRiIonicCqWwCdn9VUzauUxSwNnSsmW
mcEyqwHRo7rof8yiTKQTsn5woq5CezgLN5ayWBaYOjgJjTO1PV810dMnFqauQy4Y
SUv7ecwM9TtI3KgD6teBKdyRuctrtv03AVGIf7+J8U92TBYVxzlRWQp42e9wVkzp
gJpnC4LqMGZI60natgZIFdKiIIOujs/jKpHVqdax1M0+OmeFsuDcEpB92MycL0yx
oSYk4DjU7AWSJFSdW9xQSQAmVhKhW3CE19HawcjUK93GWxKwI3JSQW26Ir/KPtKM
uU4KGTZvhepMJ8H/Ok0jBs9m8QA2jx2IlN3GoKKHxkzGQcY1EIjsGOfJ90lO0b7N
Ez4ylHVPXcY9hjxylp6KOf1h9yzFMvqfOsTeP0r6vRM=
`protect END_PROTECTED
