`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8R/z3Yr5Ixxh5upw4F8Uqh7I8+/hdsdYubz6lS5mu1+KFx9rETq5CqIdTNTW9ux
/VF7N1KS/JZqsWT358mqVJVxT3DVkej9TVwXMdkRNA/Lvv+CDAOeqgCmKUiXi4qe
qeSapOMzugbvz+os+UlMdRkQMed25hm31Y/ca15OhZMCYnnrjm+gyGp0xCHRBPAL
pEs5kQGNtjwtiusy5w9FFw1c+LiAvOv/wE7xoerRFDpYuqqnlnpYbjbph7fnFQ2e
WkozBX3FQODLHQvmhzvUp7bMML4TajrhdIvJwPaKd/GHCl4Sm/9+BlFXAeRTqYHF
7uOzBceLEfECEk/i7ZFoZpsHT4KL/uRMjCZK+GXXT8YCh8C61Uw/MDlJ7b/O+sB5
9DSa2ms67wMQoo2CngXMknxaRykfJazHh9gOnPiInJZZhBWLzLPgfMdr8iW2YUIJ
3qJLEeeqIKsd9dIHUEgbiKlObVUsWP6XtoH/eN+5MRvg43NC4HwflvxfAWLJJgPp
HFvGomCbJ1M6e/q15JjsVMYQd7DgQYprg8LxUywy6wFRvKv6jSqXvuLP1EhCenAQ
qaMQzp+/9yoC3CwcfHn3a0OVLbw2kIxhpybCsM/mBvthyms7rk9jMmCrpDCb+d0p
SAS35aEl5qR48uq9qiXv4t1YDneiYhK+bbZ8FfeTtJvPtWXNOjFAY8xlRKZwfW4s
16WhrEQUR0/MgN4hj+I9m029KbXgsXCs0GfOXXDbxjrS7IBWrPPHzEG+1Jn7SZ70
`protect END_PROTECTED
