`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eyIkE9xKwk2xfrhvDVgEdd2NfZwj1laZq2e2yGgnjdYoqsLPbp9fvi1cZp/rkdju
sR2dGIhpoGfVxUwF2qw0vgqCcmE7sp16UlKREInSQU+zo8Xtt6rtEukF5frMZXQN
DDbjSoOwKqrIpti6TtW+DYVZE1tDf8ENoQicz0MMqVmdIzp3MFHq1loGpeWGTMQP
lf7wIzxdG5ya5EzthwvF83aAbSmCR41X/BOc5RYUxiALzOD8Pw1tMCXvEKUnMGka
74kMgQsJNBDLRIC5vdJ8YKIlE42vR4R1Rwq7Pcy6FbuK0Ze3B1TEcEa0gwqkaHax
fkrqY0r/aXzb6lepb2yygfAfSpq99SZmYgXl1pIHxPn5oW4aQPC34majqXYfMdKq
mOw+S+q1ecyiQTY1N21s/d/1CNAXBoDFOepHr83hKGNFjHnWcIB0hDWV1KtQi8/d
YhN5FgGSFFUA1FmjQQtxz+A7aGNur0mXh6IyCtxW0EsEsl4xitvEby6b4/yW/GbN
MA8UNoJf1s/vrNGUwlUX10pgd9g8P5ZvbiJ7rh51GLXsKUELh4vfHpQMhZaZ2FeU
5FyXFuWTTd8A0r1Fgs7Z6JIsaGp0RmkWXP26qGWvBGlpHRtY2TWFCsF/RbKoqfd7
qyWKvrpyX6LIv0O8r/7QhCxVstDluRUiJ/qsBE7QXIdh3VngiJW3L+nZ2Iizcor3
tLSRGAwHyX+t9fTjzB/z3xX3q/5t51d4Z7zg0dtAaPYZJ1YfN1fFbr6Ne9p/XOCC
wFsM0DyODVGt43rP9L1eySN91vkBOjt6Bw7hI1q+h1ykxDsuCFB/g0cvyYvEkbpu
8Qb9HSWaZERd1AupuYoVbjTGLIxpUHLm/PMtKlNUzL/YUAjEV0b5fC+zhsPI3i6T
gtfdsqRD1cG+7K1S8AQNvz/iqhdRyvky8qkUhVMSjLgooNe2Tb5NP8ckTss+V2oT
p0a7RDt3QhwWmA+n8nHav4yZudGnKcoJgDuftJcGmE02bapK03ExLMcWvLpqFwIg
VR87jv91KnmazfID86ETKA2/7b6VSjjtKb7G7dsVd8Mt3GPZ205T2+2+b6YkLYqq
P+iPbK2ctWeNX9qgit9fl3oH7SRIu0oNsk9C+ro0Mb/2d+ekjOznwvecAH2vuomD
76m7V8r5e0djAmFj5/knKlyxQwesG/SArcQ5YWQEvGZGqxATMI7Frm4mvGfrLAZz
qzTTjYRhI+1tqn4Oi0bhwxkQ0YzfEwNvrp5++UNHFTRFXrYGHXQEObHg8QuxrC+x
bF/iKL5Z6/vLWBWGYbCbce0Jb+0tFqN2shcD5MoLjqncwFtrmAQ6PBUHAJy5gAlC
3+nJC3UKVv07DvQYdP88jQMzjtx1TliHgZ/V4tMOx6oUa5W4nD+dOrbzFye2GlGx
vGuqgFgDH8/Z+DvCcbYx6CPrrvu1r1A7Ia7fiHt0iq2t1v+ZmdBLiiTeQ5xVsDOZ
hJFZngBHI1UJ0QoY+3s/rRt7J69YYAKSTljiT8Lh0zLFVRVrBepuXW00FlgFNgSQ
VikEynrr3IcR5uCCwENSVmoi9GDC5uNKXvU2G80jUWPrbqzCp80apZtgvLsb82HW
ESz0TgboJfGYx8jxgDmJdE2QTm61v6CppOL4xQ3/hi3iNs0sCnvY/kybddpuGpP4
XwYGIi7QGUJ/4gwEfLwV4YfTcBbkbdBFgvs5gc3W4IhXY96Sgp2i9YRPLHQfew79
mV5hpzio3X4pXtu86LSQOFK0JlShFqlm9HSlLArLcKKmiyxkJeb+TnHYK+8dp4FF
UF4qv88WYDZ2yJzpi/3yJinKUl5BTwiVa0rEp2N2mj/zliuy85oYUkF152OD8KgH
fOI+nb/lashu+zx7d5tHUDTRvQYB9InudoZa9aqb3Qq7KjhY9hW0fDSHuUEe7ti4
8qehof+Jh5fHHhB2KRt0IxoFqR6QqTpGqeDj002eyqUBgL8ktTMtzKYGa4IsfZqW
pqumBA/h2N6VPO+0vQFKvfB8MWqS7PszKorVwwd1nYHCogebkE8jkKuD9gjifxaq
PeOZ079EUv82QajsfqQBUjcxdhPvgdQ68bW/zPa3cOIXw88mQtjUO9mgm6ij1yh3
2218SrcNvlGrcNkgm8CSXTFbXcupzC83JRs1WuMXGv/tphnN1WsUF57eCTSAfl/7
adtNpnctWHMLdAvTVZUBSgzllhBBwmWGeYg6jc/mLlH9Lkj5YmNWKx+KG5QnItez
yBmwFOT9RPbl2jvABbCchiPSJ16y+UYQK/4BL6hyUdAhQMxYJOpAWUUqY7aOOehm
Em4Tbo6lJPbnJsiac3B2W3+E4EBN7O/LCUmISGvorJr2JwVXpW8tbXVpBhaJbrGt
VkLdkbxzrxRYXpwciZYi2rqKMeDpQSV7XUZm+//3IAR8Fm9ePz3EodGK41pxfOrl
HB2yayJuu5IFxlhTgBYM+foND9aQrysigsQ8tf0iTVGtZAsWG0dASB7g9OLiHAcp
Ea/mvYyJ6D1fsPXwYv/4CTFFrwhhY/g9OlfjjYvmVlpOy5UNS2WijHGm1x8vjVMA
78Kza81I8jCF+pdGhrwaQFQvjoNmPbhHSNWmmhI8eBe3cbG3H9hp/LAMj/O9njpO
4QlL2kDLOnKoBFg6+mGXl+/I4KUlWvS3OZzKJ3hBR+llH0IMTc0rHCnGeiR1krvl
LG8f7LNIecpFuAw1CKuv4fdHVt3h0GD+cEZyr6lSajWdjUINOPtpeZVIu4rUakBo
7qsgUP0WrTGxlIOyElm7zI47g45TaIlndNSpVhReaPJ5ODrgjUqmNrSzxdDfjpRA
ajfOwNLjsztrb49eQddHyxTNjNvKirBE23x/0cc/2N+YM2YrMJBlb/i9GYuGdZuX
kGyAXXbx76DbD4aPJMvLz0au6vOwQAk5ebdiH/qYJ3+tUzd43ZcDk11zXDqtKWG4
gsR5HWEaiIPk8T2Rc3a5N8VW2jteSnVqN9wh1JZzi5VHcSe2L/dB1ArfdB2AuPNG
opPqPzNAyZo0dsMVomiQB7mGntYQUkEzQKsEmUajZqWxHPmxyHmI6l6OMHjFNLRH
E+u8XPrBjymn9ni5nJwsVUZRGMEElS3DQoA6AK+0LnS2z5OOXc6k+r0H2ln0w2QX
ymKnCrZVzucIBA8Q0AtvYOhrZxYkOtYBByR7fJ2Ju0cLDuGiTrFG/RkQWlH2j64t
ehzvMH5kDZiFULxLYfMwACtTQD5enU1VOiX+8XUF4XFCl7LYSE4uZWmfLbtjYezB
E/CC3RJGUQmE3d4NIbAoRecu7SkzDaG+RErKV+pPA/BrFfM3cdPFK6cu9D3sYxco
YRabCl8xhl8rrXwmgRtaUtw1lch/jELE4mayZmaAIy5pTGlF9rRr/wa8139iEHDW
YS2TBvBo2gPRYnprA21eA4mZe1iaj7Pr9YK4EE7ksJkjoQz3tntGt7QhfN1uUCXc
bnAGGNAd6TaE2ag8XoT0GfSdr/IanwppzX13Jv4OMdzI5zt7nGwyoga22n+ZWkHD
w6VcrhwAjp3RPeaR9XLAOPfXEaD7mgcFzxsGH5U1MnbHuMFCWf7lvOP7Zy/twJ4J
1Oe3r9byNKjW21oxKPE79FwmeVvodUYmSL0Zqc73jMIcQO4FBngYrSn1Zetwrm4A
SMdqguzidePB6FwURUj7qWrEIlo67eLZinc+VtaHYLXh/VMaebXYX/XZlPO6NN10
ajFqAAQ30Q4v5aw1bT2/Uz4x2oki5nM9YNNKKtLwotTf5f7Bif++ZwqGarnxD9K1
FmrD8o5STFeTZaH6xgXUw+EcWeUKGuQKa1t+N7iMnQpyzmLkOwSdpmautOIuAeD1
W+PvHIhs9s8EvDBfNAd5s9RDvfJyzXEppQPuBpUaELcpp7Bho4gVX9jvK3XtXDn1
JTwUZrH6Bq4Pacfs20S1dfvw+lncBpNTEIIjVeRzvp+0S0GRAKUZ+B/q8+exQdZq
cv+vdd+a+Aaxt2RJQFCEAEA7V4VY0pVRy7nOcgftq/oGu1JNfIK8Ng7Pm8kY+ArO
nGYHsCanQbOYjYXECqwePr5FRBFvTV8/QVkN3uj1QVs7ehGeZ46hol2RrcosO4Vm
EkqpzfgA1oPX53AMuRUQRiCEcI5v6ktdlt5kz4QLzZG9uiSsRpz28HJa6GVdes0y
9YywiNF24uar7W19qFtqLxObWOx94rdExpNmzEs/3texVVsricFJ4vfAS4J49RMf
0S9bpXoQPGIZQgTlm04gEVOv6LAF3T+gGhmveo/O8vMI5tIqQDk0XzbFSeZrKxvR
YaMYs/r+sBxMq8PteYU7vvo16ZHq0K4ZSd0WcP4tZJkeTEtvhYZmRbG4LXprRUBs
XxJkve9vBHAS900D7a4m0yBUOzGaTEwl/+Qs4TyPhbjiQR0zJdI/74FNZ2qi9JXw
qNXnDbDls7p/7VLvGA9QQ0yu46Po9Ce70Qt9EOnoCqs6qqUW+eSV7eByFRtDUv8i
kDL2PmXMwX+Rz0nXqmCGfviqfZBe8nluyqvPPPEjnJp1qYBCM6PJZYUhnaU7+8k0
7fDTFk8A6SfigQCgvwwgf9rei8hOnWW8NnfH3ot6mlv0Qu/bk4SuRcMWAlKIfqHf
s5Y+EkUMd8/4PVkdAOhrRPF2IPq8GsunRCYiTUcGKyRMUyOc6VvfGevB9PtUVIcB
cLlV0Ax1lDo0P6cy1gnc6ZbUjODDWxLAMrNz8gm9Fbnj/VyRhA9K7bgJajcIai+S
B8yUQouyXfZX62VHY9X1u3gtJBmjeT7z61XNU6HJN+W1d7QxrPGIJx7XTedAh9DN
I/kX7tOWLtuzPGSogPjG1c3hGAPp+QkYTHDZylNQcCch0ogfq6jSO1XsbHzrQ8dt
lE3Sryd4Sw3T7HC/m4K/psBLk8o53DsLvJlHtxN2ERzkJN/LbqUcdWs2YK8rO2yG
ypaqedRbZRHOgWwTWkRCtbKiN3/6/2Mejrp6U1wQdSGMLDgtJIXvLNn1Fx4bbl9n
kiXuQhMCJrv2+/RMOIqM6TktXfcCVaxcCFc/MUdhrajnvmrp7ToJNCSFaw8NQuby
CR4GGsgecyabdmmi2R9uoKZ2kjZ9OeHXTTNKURdx7VWkNmR6Saj1Dx9ssdjWXCs1
0sAsTqAYzCbxA7iqdcclgFhoO3ssionfoBVa8qyY6wGs7Iv1YTIkxOn3dwLBcVML
enJBMm9v9DSFYixpSMfKUKspvyZIxbnDLEMNNR5YVUhzWWZ4HVrvOkn/VyoYZJOA
ynrtnI2z1X99k/Vh7eFqWRwndZyeOSwhQ2i9cjRmmsDTRwSxfBVYWdqnTnF8tbmM
XY2vZMhLqlRmBiuidJ09xP6uiQFx1D/LV+RD1MfbjlKrLC3KlMo5PW8qDyoJVv6Z
+In0zJm/F2Dkr4F1xVqI61qZygnMoJRbCPuZa1aUuCoBUGXYZik2icEU4/50w7OP
b7qAhKxNl6qPVIyHbDV3VPqTMnMR3Yo9oMpNukYgk9aIlTtE5CUBHaktEcas0ucW
kVP2tj2Q7dbPhiZZ4EPArOpQCSDY1GcOD35v9g1VlftYw+iujawCU7wvGLKtXZdj
laDfgq3wa8CKNyWmkaMoXbWblne/1JgLzzZEttMwrTs9rwgDJQUXn5zeVYoEHKP9
FYC4nSGwkDjCEmmBF8qdtun7MmUK+vpQ7T7BjjaBwMMu7g0Jqw1/WTilT0LBh2k8
mgVynV7tJpGP4vygSK/KLZnMs1bnzoVe6/FePHlzH7DqGhqCNY982xrIYzBvH6NP
wh8xl1+JDkLY0GBfSY9EhOikDOMcv9Zd/bQqju4wF59/PHWlFLSERXZckdobgTqc
s4MYWIE+fBX0CJT7BcKaTGxFjsjcLJYyADY6is4Y7lMRmJubu0HIciMW2nHF6Qt/
u7Hv8texOTibMSGeLnNd16NOgHaClVJtSNoVlpMXjzbC8ChzvFbkUyRL2bR7qQUm
4dNr9hI52h1iJt7zPbiAZd/LKKJCvlawKoqXJc+PRJquYAGzJSAL7Kn9tr4LZtMM
7VLaQcy3UZ4dJAzpkM1QdQsvLWZ2oA7TfwziZqwD0089GJfkkUAT3W4Ktjzj/L5Y
rfQmr4t4AnpLpEnUrnOej3iM+WqEqn03YJFOo2H+o9dY5km6PH8cqXR4NO7YdVk+
td//2CD0Uq1JcBrp7BYZBes+YJUOQUtPJUpvZcAJoj0uA30cks8sOUG8Hew1dpkP
5xHJ+7n+7EJj4yZMakcwj8pHKyF1toKQRUMN2LjO0vBWcWXKugWJ3O8em03CiP5o
O/YRwqgg6Av758nSUDqBKV2RpyBLhZdt4oADU53GdFe4VpWv0FAmSsl47xr2xAai
VqvxTjMGqa6tCe8T5w247hKqnZfrvnudc5jqLEyUSAIWrf3UStG0mfyxkJdpxByb
kmb3afbbJwvFDSd6/taplKfq7EnyF6nOYrFB7diFqcTip/rDvWIFMQUAIsWBqrd+
4efPjvCe8JiZ0vXhfW9fn9aYWptLlSST4K3GOVOcNFFwCrU6e/3yqxIhXrFCF1ib
c0ohlYZrKZJ8Eqg1dg22CsV3PI33i442Fo3hA58niaufTRUEenq/cE/JuphL8nPT
9wAUxyRMcottUGe/hRexqU5OoNRFQXQLaW9sjBuU+BVSWO3qAnXVoLAcspY7QnuS
ekxR+dNszJIUD/Z+xbK1mpKeGgA+Uz2uRxeA2nqsGk+tGSjrtCqqjizNVzjK6bkn
9oNLJEk1NmwE5XNlKSCpwEy5G3eB7i3EV9OgKXJCRUsI4k/wCRBWjV8UyggnxVxK
LJKidbFqGZNg8EiEypQ909PkBB8wLa+I2+liLUar2x3/YUbeD5Q9sKdrglrhmxKf
x8JPV8Ir4XUVKdjvoPuVo2HdcDsOaNgi1YFBywaGyqsM1FPmqDXQHFfxQRswXY5v
8wa4glZ734fS410OTZ0xg0yTbp+kh5Q7lJB1LH90KmQdoJd/oucmn4VSpmMwUQQd
4SvcIxL3SwwKwCQQJq7X4uT6DVX6r8r0PVZemN8K5xNkAl3IHetLmnBFd+x7Zaqd
oyjWVVw0nlEFJcMUm9IdUx9Wp0gVbtTa0vn9cXrhYAsIq9WAQfBwlcbeiqFQcSMI
pUH+An6hcbhFaKn2QkcX3Izwg3WqqfT5OKmwzoQxBQedfcM6zad6/7Y8O1p8BXqV
jn+BfMZzgvkeFy21QneaY62r2RKFe7l/CGDKSQvcHYdw3vovkbSOyW08tNyRTaJr
jhzP1NVO9cfPxl7Vovc61cyZQ0r7Ehs2VvdFL8Nl7Y7EzYJxFcqmdXHb1e2IPpSJ
07IG3qomZIfPr1t+uJTxezSKHnjgwckIzsahF41oJ7gypSzSkzeyMnEJP6DLmb0c
XEpTygNehwyfrxL+5aUwNKDS22vrf1iDjrKLRnc3MXFiaf7Xt/hm81ruHRod4VoI
fsLmFopeafwvFXFdG/Xei3eJV9ww1JfE0eQNdy5rYGUSx7yz8gFCoZmjmob/p6xf
V8i1Wu1VxrpRzuBylS11cEpLmQquYmXT933+/0VTv1W0b8tzCI4SJJ+8FByrYLme
VJ9TD3CAdvMAGR5/mKl2HtJaSvqYNy4HE7ZSMJiyepm2tZX7724cYfANfi5qNj0l
QHcimgpBLDhPD8T534rdkpWmJE/K+O8xG9Rs0xxo/pyWq4E244gnYUvrCj50HG2N
1LMSLG3uCt4abooSkGlfLeH+1MMB7fzN8J81AL6uokh+monCKG+pFPBLCuyWkD6/
GIoi1aA9E6FMjP8WIsKg6ucMaQ4z8ZlwHm0mQVuLNLEpy+n4khqYHwbuMxUr98BW
sT4a5px9v69fV9OlhNDJCjr7QGo4WWCkxPqmo0gG8Hmo1HNO6mZ6IyLcnMMSzpKQ
dwa3slqAFb1OIrXU93K7hbX+5CGzDh7uirLDez0NH8auo3vBX5wyOsTq0yFY3ORy
tTXbCLhfjWEdujWko4ZAo65QB8wLpkAj+5yqyChZgbFevpNk+zVlGl63Bw4AWE9Y
Jm4ZDFDSY2EuKxBWcqbPxTwB4F90eJHI41PSicFuTfkoLAiAWmiYBUd5MN1P13G8
vMiXolXSNzQ/qwFTbZ8bKEyMaa5polrQaceBkyElXYwjeqDkt+SVTHTQ7lHBcDRv
NLwZwR+egiYH9CVXRuBWsI2M+1JCFOASHV5nHyX+DeP9oNzCWoKYeKYSZ7XRibe3
VYM1I7Cn/iscn2OQukwnRsGfn4QoVXTSv9aH8IzUSpRxp0S1OyDbwvx6hhymZFao
V/pWacKwNngeFelUKklsyjXM2cdqNfmZUmAOQBKj9x+faPcEbV1DJ3eV96Ip0h0G
dNlqYm6+WsnM7dcxR4hVpUM8aMau0pUkz9a25qv6oaDUW6gih2Bh+nyPtq2VpGXz
yg7Q88VD6rKlZpTcZBFo+77rri7lPfq3jNd58vfRtkS/xDgNAOrPRPXxD6asY3GJ
PloGGzDwelKsfAGeuQnSjenNDhuc2KshUF4VVj7cP71wc4nLCEB5Hs/bVTgU4We1
uMM7/QbmlBDHspVz+X58MF+kp/gaE4qoKMo859Fjcbo1ngrMRV97CjE802qrSbHc
oigL9932AWQR7GGRFGemaPL72YzrRP/f3RlL1K0gFW+d3EX54yrPzvMcQgZJiiKd
C9rkWk6rTUp1j2/VxqM0G6Zs6WjRilYKZfPjSkVha0GTqLqzSGtOdCdBofUH0GYk
ycNCgkpuFClL8xl3iu+v4Kif0lXOu1V26BL5DLhdwaW/RutxathkpvONPeeVmFYY
HkZTpoaNocZ58yYQ/uiaczZlWmNETO1lotLMHsnsOY7gWQy9CB0ENthpWvN8tWF0
Wbpujhpvwg6M17/aRLMBV0lfXCjwR+xjPo5tCP5NIKnhMMpd51unNDCywvEzNy7U
UuI9EE9ebDaL3m93NJXNcROhpWiAcnKG/DJENzgE4T7qEQR087wSRfveJavI+dSj
m9vOjBvFQnS6t0C3EsylJ0j4N4wweSyx7daVl4iI4lmcSnfyC/1Sic9VPeGAdRyH
G5I7bqpJhD9dcxTx1j3HL2l9xhGCLP+ISvFYbG7l51UHV4RNEsRemBAnJBMp1Phq
ekpCCDRgYriiHPiKQloH/1PZk99gxUbBuWytCdBjkd5awnIfHAOFpeZfAvrBvIDY
S6YQcCt2CK9SRJNynButO29jS9FvioriZUqF8sxQ/BXYNsuy5vqdKuMwHmLO+Qhz
Ts86P/aljR98yDQYWs5FpCj9iWNr7/QAtIdFG0KwzE77liSKQ2VZWtVF2/FRngSf
oLwzN2NAxJKhvx2L+FsBSKn/D0/Zo4c6QZPfoU6MsbQWjl46qKRB8nfPisJ12f1D
SVj3+1ppym0OthywanLEQsBwbWhqJbca5HtkYh9wXAeSWVFrnYO6rNGzbmSk36E6
sTvwqFJOS+RHgZfVXFSNW2P915ay4HWkLVQjS2LTJbYVQZWw6/inO3ZVGlfY1t94
3tY4JncuKLDDLbZEXlFJc0Z91zaY0QO1P5Dsxlo43w6wNRjo70ua2H9hUhYKs7j7
E4HZmSLHsWU79TUXaqhqj6Wl2x4wLd1D907b0iFlzXNIpS8HdcsWB9puIisccoBK
AULBAJUEwp6tsQ67CmfhDl0JfFCeuGyjEceXwoXzR27C1Fb52JntAUJ2WWA4NcoP
5iJSzjXdmYqId1ZbYCkzC750PaLnrwxZ1cerTwkgV0xIMczzjSlIvAnY7G5X+zP1
kWHgejMpW4oyyTOmjEUKixc95kNLR1G0PxP5DK0j8nrNwmY7SWcuLt9ey/LL4Vuu
wCd1H2zSuH5NafgloEhUnta5sOL0rJSPqHIX88p7KL5ADENHdpryGEQ7UesluWHr
zJpXBpAmCrdyAMhBg/SYutO70mGC4VHOrfoaHpvFTcti5dzqASxGOBkFYSUPXXlX
saf3s3O6oGjgLlVuukEqMK/MUT0vsMC9MZzP81193FHZI0bmVVdHhNGl/6s5qJDo
unAgn+hqHq9U9jhorgx/teBRgSM3HybwlAKYdsyXpjoByLcvI82jeoUzkibDp8nC
IlzZ9CAlp/33e7snymu4TSvPElqIz/yOL8lgVce3hJkiNpt+HiT1moQW/1Lw9oLS
xLzOzKedgsYWkVud5LGpaDnYY7OxPm/e4tg+SBEEM6FizShH6ebMfrFEkp6qEATb
LL8QHXL2ifb/Co5tnKTJj0KKGfbE1XfpTWhu2VgBNfK87dzrIxDnSEoO3QVKzpLC
JTRK8Nl1nynfcqoZhetOnQnfYKfm8vn4/bacgS2aolNfVgXS4+lSJeVMxipYzPL8
hElJOC6Hwl13UC0FnIuGXntk7rHiHQXOLJUzm0Xzsy3hzXZVlYhw0yP6zPb72Rr0
YQDAdIVU73Eg/xjWCeuL8T5jVy5S76zd9h9QXEfjevxPlRTYc1M9LLg1DeZViClK
/h+fKJGZMafjlHT3n/8U0YVzOnTdPzVfavawridU5taKZi5jI43q96aSqQ0vVqrK
Zds91dc8QzVPlW1jflXuBPloq7aPHfWsfXwzbzcN2+DXPPU0vOV+4gsOykWcvoR8
TweIEiLVZKsbLK/lpzzNoP7tcAWFza9PpcTCGmZvKstYcbtqi73nP/ezLfy6geVS
fllr6F24OQfQCSO1o4BkA1APudBKFund4yncUK2BKhFMdt80D6nLL5KS/ZImnI7W
WvvwI5or3BdUQvUr20ZwdUD8TZZ9FgsnDxfhCzPyiGqiBSZu46fEOFola3qgIvdY
1a8xlx1gElrraFJnnQ1JifxCGpAoZyX1y6zqpALyErUxit7II42cZRI+j9jwpPur
TlsI1B7cbNWp4KxzL2GoZFYHbz8gxJqU3xDnEHptXuUIAeM0vcjVxvHtHeb1ZFGc
noxdNgAJlXVNVJA5Zt5A9sM34XbZLeLtUQaIwhLjcw/ApR6zUv7GrTezqWQTBJxQ
BI1C3ZNVNmaadDIFFkIgt229IMLrGLPP6Dt5scPhK0ZWyCf1Lg4pHKie4jIlOEpq
aRm07eA2EXpX7XM7+N9VGKgbcDO/sCDwpf0VuYGvM6gnXVbs11jtd+t8cg8XKQMh
LjoP00z6dvfbMKgpOReM4w1I1vXnhvI4hspN8nWpK5T6jfL1VZeiiVG71RyTWwqU
2sBvxwyZoAOo0YzXuJqpKl5dBhEI7FIUkdEYKLHDyXOazY1UD76RK4W20SRU6Ypw
rFFLn9zwN9lEBA8YVcDjDGjRZwnLTjZSgb2ARSyEB3gayxp3wLoZtgjlP1WEo1Av
5sofNqD9bF8YYGGD+Uq5uqwhfg4FRsx/Ib6y+QDsu7bo7YyQrBP9HafWmKyI4pzt
p7i8C21PS5Cd8ACiFCt1kwm5GPcBEnmtc+sGJfBVGntcamTQJsFevB2yrod17VB0
6L0DZdbNWdpGu+Sm8tOaGRDrwoIBC6rvx9lR57B4wsqUBZKdRcgZcRjDLj9AD71T
zICVHhnd1MiRSaI/x9ZVREPX2bDVeErrVd5p0Ri9aqxD2nvEuTi7sEDcP6o4F9Wt
MWvlVIZmyrm39hnVVSg3YkE43Ym+fu8tfBAc/IzJI7E+b7g02wcXmocV2ActHKKZ
l/DlhbjW++OLoeuWyeoLMM9uMqqP6sMFEByRA8/2a+3/fVOhFtiQMrcaz3FAKvuv
h5mDGlsnOp86DtHB2vqFqyQwiocZSVdYQyKaptErtDIcZAcwJy0LeQZwspSuWm23
Mg0qkH62BrYY4oJIkC3bXFrJE4gNPv9EMx/ZUXbSkBkNbnZEmXTkwZF7sc3NVIdg
bwjjGBbXjpuCIh+qjuv5BlIdimCIpyIU41HWoWAr5HYcjqPyMjdwOO0duFGERpvV
PrhZVKEmnF1KiMZNU0x6Ht5Hu2SBn0RyupjI2IY8QTaghgyoldB8YrQSPjoUaBy3
AW+V7GxwJF02n2qdAAWHg0KfMqCet+TDv8FZbgPfVqN/bPuxSWdghIYbrv0HXNBx
zEEIWSRPepzTKmFc57808xB5DxxUgrnaVoxe3nTSFGZWDl36Cu7NEtNpoNAhdNXz
PyZIQp8fnMdLl992qDtEHwwitDYOzyCmMLvny/EpHxcZ7+XQQvhGmqgmI+V2wRw3
oF0HhWRlhKM4dE/gqkrogbYjH3nDYuBqy/9Z5RQal5kfedpZNgcAZYFVJzUFoONS
3wAjCmBU+dmkW95KoAuMsOaO/0pRp1mNCKAE9s7MEQtXBAoHbFuNfe8ZpGh5EdTF
N9WKpnaeBV256XMkxBYyjfPrDdaZI2dcoIgJzWTCRTjuq5YUxSUgB5F+Ugb8r2Ea
aUN0oU5nhDSh/VjNtvUAu6kATo2x3yfiNp5kjV0/P7ImhxjcJm2LDlOCDj2Cevx9
KceSFJfRlcSyd8juMptUVhZhoo9xZhvJM2154Z2Nyffn85Ss41no9B5u2sApdbc9
A6vzRAqP/GdtfnMSjFkId511L3bBlzy03WNSVbmpcEuiuYd0fa0kCDcJiswGA3PC
0hhB372i75Euc/G8lCgrfTVYdOswT4z5+xpDd8Ki72w=
`protect END_PROTECTED
