`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSAG3Bp7mIFIcz0ym5rSHkUuchB5QB8uI/wxdHcx4OXQHzrrsoJN4s4Fl4Dh1JsU
5xBORU9vaRCEIPR0xqaBTd83ohpxvtaRO++9pGD9YN8vQhTr7+/2UKY3kO2mG1AI
TSdgAQxS9bZ5vwuuFFXt0tfBzd3F2ybcSdsR6Wj/FDKjhMCLSWQvpYg6jz6Hiw7l
uvGKjJUbosrte69wmOaQ1gLhgAnhK+UHIUhaath2izz4g9I/9dn+o0tpG8lxA/nK
Sd9dDZgx7MBoyRLKMjbGR/4upE9PUVCOqMYvt0twStQ4XQTJR2XxXCcKbLTxisZD
Nk9iysnRpnU1kwsZ9Q/QFadRtgBzJIfvSgXDMuvnD4TfwIFBn3s9IiUmD4dL6Cy2
ADP95NJ/GRhsoFL6AbyjZ36siSa/gaLosIqmsWjVXvVjstIGiSYB1MKquHWyGwMc
AtSYDlgl2x+o3g8o0RSvFR6eapamNMWMJXytGacggkH0CmjQmrbeG+6TABHSGX4N
Nbls3Vr9X8DVzBEjOEcWCzrvntJP1xyFx1OoTz3WRMgm09U+Z5Vo1qCI48ECbA5I
Xzvj1rtgewNnnO3G3wJEUKI/0IV2la2OpI4g4xH/CD5RlSLR/DHwHxJhkPaokfqO
hA4IZl7qI0iwATKypGxCgtZXqTJlCTIbtbgfOPojxaZBCqjvEi6+h/x5mHPRoWB7
TOuQicolsLoFNWgvRYxbMD291QdW7pBjwG1M0H7KYuSDO2nsJ1jC6BegVcWI5SQa
qBX/z5cnARCHXlx53cBXpRd6LnAfAObvuMKn0vH8lEIJ/Ui0bNFeZDQgxFPS8pmD
5vNI8PsYj2pOzufXTHhKDZi5AM1VIS11yxyJOKqSQQlnmpjlTn12mXbGpWx8HvoO
6OviyA3sV8kEzgnYE49yiu4+wM7bcxtjgTC9j7yxa6GIvUvP7ZXtqLifO8zkp3Wo
uZwQJ8u7aQxlZkI/+sZFcpLGNbD/3A5MRcOSOQ+EnyzlGbaiBHkzG4vHq3hnEdQZ
EDriaCMTTnv7SuKjtg3eQ0HqB4BXBzBoX1ZdSedUl9ebPgSNbxkFOuwMPXcaIjsK
d0YoFfFuqNss7AOAzQtmNnFJvLTQ/+WdsONgfbbCf4iM+1Ok7mg0ik6jTrC3p4p4
ZAC36Gkws0HaXtiAaTXcIdKP0eb7RvqNrv9t7o50xcvq5drjRtB5iTqzH6deKluO
CvK0dYtRlKuI5uVCmLpIm1UBHkcAm7xNrK8Cfmq5JvFSYoamHwZXqbpeLcPFZwpg
o8ee7iOKAame6QkoI3x/x4Ts1XjWkTTKau5dieTeX9nxMiEZveb5FndA5tPfujbn
kukhLFSSgQkc+UOmfx+ubAwMrruCleLXW9bRFH9jMwDVEJU3VVqoN7AUvceOWa1R
BtcgnwkXmvEA/i3USNzvTuAeH6Y0Sz/UfSm7jjgLQmsImYxxlp2X2SBH8LGDVpl6
ORmN06jx9MOocuEc/yHxl6UTp6U3yM+ReZG3lOEnx9zGz1VbmHCKL4jlqBmcaH0d
c+Beja4bEh4J2674WNFSydgcmV3ThA+c+I2oPzkfsCEWvmyvuZtOvlnb6PH6qBcG
+jDDQ8GynljnV5jK6A74WU3xMFmfE+xIrT3WUr7NhqA=
`protect END_PROTECTED
