`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cKiJTbVVjkz6+NmEI1951LvUBVYEQf/qmiozlozSENYJK3hwAPX3faJ7OBSity/d
5Glc+WilS/4CPIk5AlW+XyChTZnUtLcG8cPWElZu4CURllcJuL5lDb6L1npHgquS
JfPokjL/7EgUs9a68x2O/MYOp3d/WM8my16/uS5s4a7dGCOqKUmolMSqgfYPEKMc
fn93TFLiTfVKKmhVwuCUkPaVTefL/H7/0j4WiG/Osx+hQ/8bPEQ6fdLmviEOJ0JM
B3BAlFJto7L+P5PkovjWjOKy+zTwbsgxW5enWs10v8DQYml7MW9BuJZ8YTeFDXy1
4Ra8ZuJfOblkFC+6pvGDiY8uJHrNDuv3i0yyhlVSE7d8TgPKkQBX1uZDQp4LQTow
c8VdPGx4JJkVQSYoHlmCuJqTVdmiktLmWPAmtpk9CSZj2iZQqnjrzJSN+ujdmkVO
8DhX7naaJj3CNOQFuz9kdAPbB3vg7x4MncHL2kMAUwHEQy6GJ+DdZp1lgQh8oVIY
bAVR34VYrLhbNFm3HyBI/2PVBCWC+xk7GVz08BQ9xK4bx0+zTKoQ2d1A0WxFH3XU
N2VvtphgiYT4wSxaUy10vPPuANGhkz+y89DSrGwJmqdTCKdvQI3lxKMqwo4fmJpH
8xNO0dBCHHRcPOGUVIRJWngXHhHFhllQWfi8SrqFoloZimQAqWfxC6mgsm8luU4U
DvOMOTqqMgeKSlOuc7WQdau6xV5WBkOMNvM+Wvu4ZSkdD2Aoy08yGcZ7evbyZCb9
CBzboSxI4xZmorsiQpzSLTF5wcjHq+X9QKHLrHBhs6LdaBG7iz79PoriCL/isQ+V
IElEAfSfjvnE+R5/FJ+lTNr4vO+asqDnhorulTKKK2OzQkDLXwgZti6J++ptRl31
7w0KAxHUvrx4Il1vi3dS15vQWDB6pXVkDV1BqNZh79JivnGCASvhkemvqPMuWIdI
3r2brv51ejDAiRv4qasZFjfD+Nzse1Xb3WkP+HlOEgHybAIhryFJr0e/kxzDNxhb
IT+OwcMPnP3kmeXtfE58rZ4+qtNze0EuJLWhqt2if5YZ9Zk3V9m67lUV3vggyIFC
/RMrI8lB251DzGE5Iau76PkxntHZSFZQQutU/vedhRSsEh5RXotVmsgldb+jVESM
gQqTF86cyqQ9Y4HTapqhMAyQDPhHNtX6bQ5pzNy6ltHvrQNUqfOG94n8CC4X72xE
0eqE1x0Ai5ItZbO7QSDMnYOd3F8yhB+4MWFawm5krhIBlolfl3EzzY9DgRB7AvDP
frj6Gz2Y4QiPdZ/ATRH6w8CVs2VKlIvlx6BVEouGPZbrCPOL06R08/ZqzpnyWa7n
36IW9sLJOHNv/3WVVWZyjOR+riOwFh/MJtouPVxlvU/GC2XEk9l4gY0GIfJ0xlbH
ygkiShSd/SbFwc1wrYAxhZOssFKACtFP/9fszjVUuJmunOyfng7BoRS1CFlbIojl
3XF+vIQmMOsJXZqhE5aDOTWMz1YyaIMThKrpWphygMN5+eJDxz7FL/DE98Qc+8xt
RJLbOhNTthRg98zOvBADK2vU6OD1ErweE/Fvb9q6i8/hkbW/05QunZu0iAB1to5c
ucXgNbPahLs0DRN/1e25lDf0qoSCgn1TiEN8jZygEnY8S0AePeTam6dGjryikrI0
pX4F61Vc/pWdVZ3T8mdJuCbQHF6GSyGxdKKrvz3lLH4GaBgvbZcrNIzqxsK49Nkz
z431QY0kMnwhj9nF0G/y9q1+i/dSgPT5h3Fk48DWmgsiSRuWwjsJhmmyPgMkmmrX
n9sjWghX/wYIYqwj3zDgat4eHDK198yWEC0NEM4Ocy+yzP+2gbGhR9obr3hjglb1
/Ft15dkIZJrLXJEY0qjRLqmsIF/NDe0oCpR43oyLITaCT1BMrZzRqjMLq3tSUt2N
LBalL86cVAtA2UPjFaf+8IO6yWNQZZyJtP0oe5YXE5Hds8jQIFyN60/TSOp5ZBpo
4h3tgklZMb67jne4A81jv1MjlcPjW83qIYGlnXOg9qOG1Uhi2SPfUrZIGMNZEbzO
opdtf4UOIHUBfkHuBRJ5X8VwwkATMDTnhsJB1sQucZJ2LFCIQJcrVxWHP6ul6xF3
mAGEqdllHhgiqEdRDrun+4I3uzBc902kLf8F2+KFOrv5OAJ3fMV8n4w5nCOAbEUw
tpfrTF/Aso2rDKgxCQk8rimXBJQtO5tIJtUGRH+AtCiQLgZe1Ty1xC4ZJ0+CnGz0
4nhk/un35ilaE9nmWSUnP1LQidApkxXOgnMwCyKFEfrkNLZKVKL0XN2jDYUWxZA/
LwvBqWIgJC7peW87CM6sLy85Gkz4Zf5fARNcTzSY3XJ5BMKjSxkj9OLHKCIn2nXu
CvBvCQDkMiHO/NDNGoQTx5C7VVCqmMOBM8Z+BjW9o10Rc7Y3V1oqVFxLjDtu2xGh
VyylponLaJxv5BdfQLfSSSezxbPpaoEXwcCa2NfrkUSMwodWR3nN2yDR2CbUod/t
PHHkgNKwbko3sokH9hipaYahFYp78dJHBmcZmslHmH0biReoI5CHJLLBN6ggniAm
Al6yxZ55KQxk5mIpB8D+LKnFqlDeQ0wvvLa/0LUrj2b4OjZwpaXExZf21b3BTwi7
yp2OAvFaQ8J23rJPgs68n4YBHKYZeIgZ9inMwUrVUookktlE/qgPylp5wKuQ8eyZ
5559ENEv1j2ffIRAXBafxaR+BJCvk8ZnuPuw/EXclujA2K/8ugvU34ykw3e0bpwd
rfeUCRyYaDwRFdSk/fIxd3hJZ8IXEJVIkEswDU9wchDVi4XYsrkg1MNlipQsjZxZ
OMlDoUTkiOFFHdpW1b2VTd64chxkc5ICzIrzq0ZU70YEc/FhB6bG+xym87zXBFlI
/v6hU1W51fEACZgJCfdxpw==
`protect END_PROTECTED
