`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rH7HIiZt9rlzL2SWIEcNV3qwomT6mRuJbHQanuz1CkV8iGwyXkSgUdiEGVobv1Nj
TX5OhaP8l4CrqQDJPy1YmRaGuipboGVX96NnE7Pq8WWRpTWMDbwdF9WGFYwEUgAm
+vuqnNID5fcEjBGnXKhfnXVosmLWftiR03jUXRCxFYiIshKeXNo+beOqI8urZfO/
scY/8+SYNbTOiAWend4nTllniE75uB8Oplq6pDeojkLiIeup41mUkPHE9vNSMNX4
H9bPGjfL6kzkibHZCrXdKruZ1k7Mqf3ycXgxhOBevKHLFVkGqou/t/aM9BUoM0ER
kzEnSbzKaGLzXMHtyAppSlbf4XAIXBQUAan9tvq5giRZ4xJ/PJ1eTYocFxd+wk3z
FCxqwwWXc+sJaZoQOpWztUHDP/oVnt8StbN0EdZA4bkiIBzKvkZjPBFMrmviutEO
9XcM9PgJnZ3y4dvehEGIGmb1LIJDalEYQGt1j5saXfUgaQM72CMYe0y723GqYW9t
6kSwur6WmfcUUxR09piNqHa37NTfZmQXy7xu+hwTjAHpj6VZG4ez77/DLzv7oGXO
utYJoK5lQZxcE5W559AzSKFdYIrS0T25SFIlIM6/DjJcUIg2AWhaYKOwA2WdntHq
O3lAvpBpRe8W/NV0+wxhdNO0FKjuWjKuHNVYRBCnk7UgC4qMzNVHGDckzkHMcBdE
JEz86Bs41ODzE4tYd6nMDHztzD5Eob3cv9BHOLVn4gw707Ovb643yS4MaaGYmM5v
SrXPkVr3V9EO7UMz85YaOkTDwRWRLka3jNHxH6+Ze/P7kJl5m20ws6VoK3Jm5Xqj
piAxT0Kp2M0+t9EHAuJoD6MqHHxguHfSCbeoKonaNdyW237rBRVcqVMpcVLaAXMZ
kJUKh4Ly/FE28yDCeso0EyRp2uk4HlyJgtyR8hEwvwOR5AkBXE/H6a5PKymMAoRg
bhEo+ENnrvg/ingPphZTQiQMYHZAaRSUvtVvA/knMx5oi6kAzIMvI8hoQ40N9VfF
fxhBkgLmuyyHej+CplCe30bOt5My+19UQBaDaWzgxHdSR69Zb0NfckpXUNGwxFpk
m+rlPvACvcmD8LLZ5IeWd4bdo9VJ+++uZZNGjGjc+rbMMlGfSu0Dn8yjFiAwfoKP
xPrZrbB/+8kXJLLh188OZYLHbkM45xY4abn0OtzElTEU4AiG3s6BvOkUa7LgVtPL
qWiZa3SOO78UMU5c3qUMT2EPXvYIVE4QMODWUgtnGIjwVQg1zHGkkBY008te3AVZ
/thK2J6ah+IqffvXeL2rGG7/ROX05FsrnupikQMr2Los936JepblHeAplHQuE687
jMPXWIakELEacTvRo+RB/fe4R4dqKkeXQvknBDJBWMREPnSDpWOq0kQ9zxMFf9vn
B8JIqKgFirqUZa9iDTN58JVjX2+n6oezOdqdd0bVOQAyWL/X2f9MDBogSX+QsTUt
+TmmdnfjtbKDaGIXNx3RYU+bK9GJNq6XiCVsmUBfBIjvXmadvAfYTs9E9Rs36F/v
EBpSvB2s0mCYYS8AIYb+ckGOwFTXUbzcXCKO3JpURQz13X2ZTn2thba7hsalKW48
0wNY1VW1keD2WSIZY1DdnG4Eh5mL+UTeGGThrALVcWXr4rmTQ8VgxVavf3YFxd6m
ucWpnqv2FcEg49cgzuYwzS37n4hNrqPzvYl6QcptZQjHe6PAA7bspGkRrbsyB5zq
XLCnEUjJW/a3q6t06El/x2Zz9CcmyVNj2GjAH5XUnCpsHXwICj7WlggCfkZ+BTe7
t9V3jtnBXdBko1FgKCGWlWx2HEbEMg/KhLbf7Ehw1TpEFaU7XBf98PMCiPxTjRaj
GTPau46k+zlyls2RzrOjZDxrvI448NWAF/C88IQU9elBJdccEhSDrCCERQW2tD6p
dg/SctWsm4Ph7XDd19Kp4bN95aDNPX7WbWtdOkAVck7tNjkW6GgDE0FyrCPifKY3
vCZ40c6omkX5fP3e3ZnpqkcIrT68Qqk8bFpwLBVmSbecPZnN8vAwjn0kOAgUGVxC
F/99brPxGo/4qweEPOCpzVLsrtG1VHCa9DUdBwemx5ePUrqtYuSJf8/c2I+He5oU
CVSAkNBwI1X3Mw6M2By6LQlx8unxVhxob/i7JREor3Wwn3H6lrMq0thaUM7kfx6+
977XR4yLnh//nbZ4lnqcl2czqul7U8YGaW1kr+Kfe59Vdy/u25ZxWQFVoSU+fK5H
+j/ZYlqeL7dM38xb4SZesdOj3JiurJYTKLlxmiQZK486mU7hoDsOSGvxKDI5HF1K
Cbnt37EOuJlJJnsSSrR1IKPBvFbEiG48UrMweKcQxHRoqanwSJkpI/YKrfle+x5V
2zw2lFBpOpw2NB3LdMUUmd1MuP8hx1cccoY3efoygZdhzgS5jb8aURqA3nNveT3s
7tmNMwxDZ5lJbvfQSEjEnWp9DLDTXef9PQr1QYweuTuWOOXO7gph5wZpsaymhR4Y
vY6KWczp2XvAZqUteXJ4dmEMApMhH0X72cxJ3HlKS5v2wPPCxP9OQcw2YBvIe6wA
IFelxd3drzgDchnXppRVMUyoSfGQ0w5pLVWdNLfQOFzvBnt80yPFkVlSrtWOsVK0
H5VixqbBJbFKFH+9Zl9iYRDV5L4vhdRLXHhlPwfMuyzw9HcbMbQoKemQg647zuU0
Wire1err9wtAu6YSTkLUQOiVpZcVNecYLpbWavQNiMwIHhwvHQec/Mk25F/p/lvw
tq53iYdTI7OyWHfKOfV3Zx57o7ManUjOXrKIHRX/JIysA4rSU4QTQB1/3wMmOJ0R
258mMPIdO8o7SNry+nvMhMg/6FjUNal8bC0xcosI2jh6Mj0puzLP3cm28z2VUiBH
hjetY9Tk+5vdrQabJCEmt0QTZZ3i8fZjiYujRhZvgIgtcPT5coe+c8QIs+YKuM1Q
kLHXihOHm4GIVoSpO4qD9fGzGpuEJwJVGAqKljoNjZmyr+sCaPhVb3EBn6F5tmHh
jJVB1zIKzMsOk6yQ9esNapnp3jGOnH7lTJ71ZnSM6uS4zJkj7ixPBOOW5KoLVCu3
ZlwcaQ80/9PyDYaCrfCSxclVFWtL+iYCclPITR6cuhp2B3knOfhZjpB2Nza6cDXy
TO1aL1sf5rK4plwwVutFKN0iJ4U5o9OjHLLqng8MxpHMfZqaNhjCeiR8yGOHRfOo
ESz+1yIvb5dp21XXI3qDAy7MBVozjIf2UIxgC5poRNndcm2oQ+T9uHRIZU5MDgcb
fmWyE7aVRaC3TzjYCYLnEjjoRhQG9M8dtarkphrx8HVprmtOtuOEeS+smYvhAR89
wIzRsX+dk1RJFNnCWrCd8LHJ+bXOK4T9fmO01tf8VuQU+k1RapA6Q6YZlg2gm/1D
w+rCvVopKh17lukRch+HOvrmVm3NfY49/swhxQYW5rgcEbh8XQCYgpbZItVR6B2O
w/DBleG5jQRiifv4EGyS1JLFIGOJ1RzkUG9t9JFSkdfFVEi5W2xYooR1nXBfhQ9N
/iiZwqC+nk9Qs/VB9UrbsA45r74AWDhDO/ydWFl3IUOPExjeE5pS1vOtiAHQdFMb
aItO9BpFBxhWkUC45EYjtxobxRmKCZs7BdvCR3OPnUjlGUn+mxea6Dhtzij42Tty
kgEByQshr4f/2DTCbvlqC1wP60JL//UarfV0zAdwxHCp79gmGc6Jpgzv7n4g4BOY
cAF/ZFT/KUVgQn3/ktLEwApA5+JKIlurlaCQSosYnP1TgrHLcG727mj1tBUI2j1u
vMUHIgpypffUtSYepOZhVlW9Xx4G6PepL9sLERfpNFdBgdGohi92EdcT39fYJx4w
SpbvtmoH6gtxJoy8yMwckQq0OhHSYEqfBNzuc8pX0Huz6CY6d9kJ6/SAMud6CpI5
p3wSxTwVnriByc9ntglFrJkkKrPbPaYIZ3V4WQ2sAMDqIgUw/P4PZ0VDCop4CpA0
+FZSbdLn1QrKoudTWn3dXNDh3tJi0N+bb9J1g52h/Lo8rhF5eE7hpkaezyUaDSN7
w10Wi9qBhiGdZgSNljugn44QXjRv9TEYu3mD6ynMt/lSBWFW+Em+gvb94vMomJ72
SWN+Xi0Juektc4/Ya7PL279rLmqSpALFQc1D6lWeX6eajKnTFICPig4E91eX3tou
Oe5gmTbBANkx2Gy5xWD5ofzNYzUNYXKNEEoX380S6Qc5xu7zkXckxuGfm50mBhuR
30jCXmt0p53pTBTBYN5yEIps3LZCmvn10grBkGDNpTWmf2QH04XWENVawhF3KfzN
PeCDi0Uukya4vs8wODcb5WuS9zE0uz5lOg3PPOCLEsMbld0J0V5gE1u7ocu7+Vj4
m2i6pxUbNJ03Kr770bp5UpmTYM7yJQkxTRbi9LH3kC3ap64BP0jtioHnVTTmk6A+
Qig0oy8BrHmHlkG39FWbPrra6LafvnkIQCayZjxI6Wol2eXEDdzkVCt6UIGr6Fo0
FuiHZxZEBjA0UfEQR95Gym6CnQOaKEkn9KjVnQGsCVZgm0mm3Gr8HTgxwWBM4ESw
BwatjSjIRLwSLS56fz9u9mY7V8xrREn+9YSI+EdqXqj7t3jV1E1xGAdPg4Hz0Gdo
tDNtJ2NcA0jgTStgmyO29sqpZEHnLsSFgpEUuQzJ2Af2FY4DQ7FkkR4LlIRqEzpo
RY501TGtV7b9FmmZ/VhbEaTbXqklgvK2qtexQBGwn85UY6Nvfu4K+vCtYdv1bczh
AOc4sff9bhcVdPgJyWQoLbZ39Rgkx4id5ccvgmLHs/Ka73vrVTResFdQ356y/DPr
hW3EpaZ3EgwQXTaRFds+NQOxal40DixOq4yV2XLQ/1UuI/X8zJsZG0apr+nmo55Q
NH6VS0wv/Y47k0skL8hDtO8Lbdtwr0eP3OGfxz7rnpCQPWXdD3kJaAFs2AzPjW2j
gNPryrmYI3Kywi4UK9ZHdxHOfnrpRuSiIFzTRO2Rc0lGQhEAFyMEFQU6L5ZftCv9
COqgp0E8aziiGZ1NMiJnLhoDKpUNC4FYTww+TF2UOO7c3USB7Pfdb+qVQlJGbUFd
qYJJX/UOl7e7TnH9qWCZzHhFACoX51PcB4BHb7omcMR2R28jcTSdjqemSJf+yV0x
qWIshZ/BLbyZtxI0+JIpMvlZhCWkIqs68Ni5Pq3A1UxX5AMeNoI2DcVeKmT474th
NrLmhbkN48i4x+xIXJLBlCAtTNur4DWzQjxygRduf/I0dqhM4g1b/R2Gvvm/jV6H
isCe5nNEz6HDjKInRkjqY5mcYMGpJiPA70oZz6DVBCR/631gmanKwrAxAc8TG/XS
Yn3cbF8mS849QuRCODifp3MSMj8wY8CJVSHi2nNXxItUOxeBljzL2GM7Skyz9P/c
qLv6SZ5HdHRokABVwJgZp9GqIFiOxbHVWdp3dLVjv2Dis7sS9FnxGxYsAT8N1Izl
4t3wbVw4oqlWHDcYR0yW3OS2g3qFNNR1iY+dAx0a6mu3yRHN/GoISb0uLOPSgCvP
myYtzWsvvcbLXkLJNdxKJC9frAwEDTYahIbl1TKJ5hb9cX7x4apTSPTaHyIMkKck
4IWenU83pAFNSu1Fv3XXqpqvAQUzcEwoxTMSu2MlIa8i+KCkqzKRu5xadeH6YrX6
oe0k/p6AdFsmajq7hmCr8pYS2oJc5ALU+t0upw72kYICUmW7zqBmYRdWnqNCMYS/
MNi+QDbGj02kd9uZMqwdtxibBmwa1ufeG0whyyqbpiHfdqU8imiZ7bz00fWYByhI
nAZv6zIb5ZQkYQ94cs9MHM6pqHq7IYRLyMty3K5oOzUSfKUcoYoA1pJaSFtXzeey
HcFSuRe/oTfhdwBNnmvKFBN33yr10OgeyZFdEWS652qzdwWH3NF2k1tpdLRgGsJT
8BhQD6V+X5EVz1uBE4wn+lRj7TB6GS0ubj4/vPWKxKHsiOOgdBGDdxsqnvWlfu3c
DaOp+rTmvqUeWPkIdyy6sV6RFF7KTHLGNxXbLyAjQGl+LFvJlz7IaF7D0vsWrXu7
7hJtofYNy8Z9vsusS6KP/F0Cka39ZhICxvk0P15E9Sxep8W9gVVP8GBti79QhHEg
tN+7F+jM0r0tlFj6yJi1kNvAnyuGGJYkDcEV6ubG/25YqUcChxs+vj18Iz/HFESG
4IW7A987VWKdGfhdX5eqU8FFg9qUnSjidS9yVJr7PiqzVqvVilJ+IDZXBHxWrUVZ
jhSi9KWTfiXTw2lTNoUbDF1ULGoH4qaYjg5I/F3PW44VwF69p/qDNp4BK+rwAkvc
V007ZuHio9o+vyb5Ooyf0FXXoskj/61z6FValo9KRMGc1kuo73a/T3TrGoa1U+y7
woEd780Y8lvbHL7MGSdvrp2Og16gfknLpTgfitkFn/N3QyzCvKzUQxxKe51fDVDc
QGd+nRGBdCfjEll8ajvXrQ1DvoABgRkZWCu4b8oM9WoTiil1XGfc8t1UONhXo9De
tD65fNRCquirIT48WTOFMKDVvMC9scERcESIirKc6WuTj9SWS/tY2lRH0hCYFkiR
q/iIJvIsssT1nb7J0UWDTNFJ/dP4xe8NH9h5Rg5mPP4fAt2QtPwfXx+YiKxo2vLb
jtK3EM6SS2g34Qzp6xIxXCKdAea2Krws3KnZlNuve7GEB/Wo/M2NgXp1g5m6NMP5
IEJWdctbZvONHn0szc4V+9nSedQKqKdWY88pBvj8yaXItM7RCYTHJ0CH7WIte19p
shP5se0Tq9LxMKxMxemORRjNvul5lV1hmfurHWObgvMSW3VyPHYaypgk1Qo/+nEK
Zc9uRYTq0ZJAL2E9Gdbxd9xkaXKcryjOhOXF8VP0GPNQPmZ4nam59bGoMz8OZb3z
f8V72z7ChG4JZEzXR5LZh6ykvdxC3QdXyFJhxql1K6Zl5ngJYTOHgn1sGXNwfI3a
Ll3NO3jApyHe7V1xlIeJRB13/aRtJJpIuCEiJfRwQ9Xj/SU9QXinvL0VAmzMktXp
Sqgl3DQi6QqNvEjhGnxywuKNtJg5zCeRrwK4Hw4JY9n9KKY+sGKE7TrGNR/D23Av
S8jseqmEO5x0FuP+o5xpnNOG5TIcUGfph02jsRIcff3lUPcHX62wcGlMDXM4poa2
z8Lzz4sE4Z/hVDz+VJZYO1gJ/9l7/ks+f9UbptCm7hd7q8UpH0OqWx4YbyXfuW0C
brv0uQdnuuhJNKdt030M1BFyrTA5w+sRfCbUU1tMhixKXx2xxU8RWFpM7c5Y0p+o
wUa57NrpkNunLi3fU0S1wUtnlz9Zbb5QBq4T7eZH5gLMzYlUDq6HMerTAj5E61Uk
0KV6avsNgtgHpZPh30FB8SityhgLUGRtEsXfLaK4TC/qWhKb6I6OpSQBzc2gl4TT
+TpAZSkUe8MtqBItZfuV9194LR3ApQTfxPLdprZItu4OpkldTSqGFYOHyzmQhaM+
57HCPV81pZthSnoOEUq5iq10J7zoq+9cgkypHKLlpEq50RlHhGZh0GKwlbuKLep3
xek9TbexG02WZfx7DVOL4YHmmxGzvg01bgJNYwcpe2nrGhGBZc70HJoN2uVqqDgl
CLoxLqh8BiQbMC5oJhnDdNOWXQ6TbrJNnuQ3YE0F6Ub+zPQOtoKELQf+sRmgMF3Q
5UPV6zbS3z8kn+QXjtNEV2qhJsrC9ItthUXwM7iiCjCXlsH7dS8z1Bla8cnQ7+OD
hNyg4cLuLBSJe69WbJD4h7dc1pZEgRjfvu53/F6kJH0dqA9xs4VeIq05yrxWahu1
kYaK7wdNv0Lwa7rXWVrv/FlFOXsf4MIBvIWraRX6sHF5keDgo908z5dfnD2ZmZAM
y+DpXpqY53+6LMFSE6Qr4odPapIIYCkpwe7zTNbmdukyZKxLu1qt5mptgQQRvlXw
2v/cl8EzhyJpTQ6uvpyQUzkgvHtRuCLB4rZ+X8x2Dv3Fv8XMcQU1GjRz3UlgZUXc
jH6/z35V6UCB7Jj9rxz0l3YwGmbSJTNbGTy38oa04KmfEpcX4GMCtTnbFS+d4p9C
RSEhO2cwWGXabmeOD1hHSsWMyXWIWQlLmaeWiHSM/lQLw5BXg5CbeUq1dSmmQa9g
9iYIe4SW8VZWnLZvzNwkkcXPSBZwJhzpJedKV08UbCSLr0Ve8McF5k5jDcxgOJZD
+QTkX3GBhzoFT1Mz3Cv1s2YQfmhEvAtTjk8tRVWjzOTLipJBQMY5QkpM68vtY/s8
p+rNjDynV5MbbVmfLUERywo1yPMqoNtc3GdHoziHkpHdDjXmABT20xLeKXKdPB6T
iKebbiIzpwfy4Wq+bk9WWM0GE20AEDmFW09W8PFX8QpWMgRaK1bjWsfP8F3Xn2oG
Kook1fgdFB9J7FD7OdboudZeTWww/bEOdOAibiVWICl1E2jxVzVdjl+os8D5DF/8
OlVvF/f42xkafYRl5lvnYCiQtdIjF8tFbH3OrvxPgUyNtwMqK0KL4R7KGTR7pUxA
daGEI+hZtnCTVhc8nanIvEg5eh4nV81O7IyWAlTiodpqeFVvgfcBnzTIw2srZ3Uu
JUcs3bBeQr5WL/yT7AbM7FiArTvVxrTN8xAIkA6dHxD8/g6/LLIevj8d1EKGoEBl
Rm9Y6TqwGhztEvTa7skZ4ki/6vuq9bjqA+xGriFEXHvHo21UsReuKCnyHZc6ydbo
MPW8+A/AK1HrkyT/uXJhJ56c2jZXnVBE1CA8ZLWtSTVhXohXiYFopaQdNf7WYjiK
UslxhtDqxadX0QaZEikqOJkBLVtrdu2qcy+OAeFIXvNvr4sEnmDFo19JnnLmhScA
ActDvWmJ8Ozda4yD/S9PvuwqvrVODGfS56BbY2XhT0pH4Fm0dfw1vUPMjDZsofTt
OgqfJMdlqoSWWcmRcy7weMbs2ia6I5FIuFFY4sKIhkvPjNHrhBGx2XigTkqYb+KH
db9kv++LlUr38fWTn/CEUDYUAjvBlQ64nS7FeAyKM0hCcWdPEjvtY+gb6CkrhnfL
SMqeaMjm90+v1SHgf+NNlnlws9nmFIrZJ668jZvQ15M6/SL3QJ1csLRPhjvVWXaX
VRCxsQVGGuzeIhwk7W1Wz8tFrUM8saMLX2q3pRrnlbGT5iC3ajUO0TlyJrdyhk3X
4cBm/zCL7RVqcMflReOS9oXMsLp2eK2ty7J4/7K9JOHOeQf/0qcyNlhx1YYtlgQd
CxT51j7IfD1SamYJ4664DgnrF6KuOSG/cSs/96WBHEuoeAa2H2ryJe2TbfwUGApd
15NoSTAphzgzmgeYzJvlUVmG4LbCJ4Wi5r+GeQ47eG+h3PiUqxE97yRKhfbtxmKa
6pSHc5SHoPQd9JruuA3+0Gd8rbhkj5tshU7F/sOA3d723ufchXUbYTGGK2dA+5k7
7RKsohTdCoiSnDuHdC7ttneaOzykgJcsNbDhF2YJ9282Rxq66aZRudNtlf1cSGEy
nIkvd9ctHnl9WE2ASS+h8V1OPOfMCRBvqKuEkhfzUnoWzAblt32lyNsIr0m80UzD
ikxNWOsu3KDBiWhJlvYHXKN1dEnXU570gxkLJbvLMwAQ6T/iMNDL6clOk+mDXPpd
ev2mQOcm4fs2CyY9WWNBvlSRsSFN2PAhKY6vDrwoegxMg0+WpV5tyobbXGhegR8o
vxGTfURqZm/t/O2mK4+gnkpRDJQYreVueoujbP+J8q15NoXXHCOiHLEQqeKkprYp
n5ZyYtQkwpSjeQfx6CTAs2C3OpLpGThNVyDLEsp1RLpRavm+5e/sC86RzfuWN+hV
zSlGDXFV6o1pEQOqAX+rexpDaQErs3ji1F9Vf4lW5iaopikYgDydqgWj7jMrWEmY
n7dhf9eoml21jIVsRtLSbJtxaXJeouc3M75rkWiZcJCJiH8Qk7uiDYrbMuaoGDNL
qtLdp2gD4XMdlJaHWK4C8EBRUQ/GYRDQodpcFW4C6F5hlnumQrEit8sNY4gGn8y+
2B5dJfXiKu+av3idy4o8btGARLURf0LIRcS8NKttVFp6CFixPKCc09xcWH4LC6mA
BqWTcjUIRX6Ww/yV0sxs4Ap/GCdqVUWjM6/9cj32CEbsCZRXvKXn53MItHSu19A8
BVmIYwoJ1+XQNOJqNYH6UoCKJ3gezu7b8PutRh3o02rl52c2WPsxk2WdXlVmoJyT
8jX0/PI0Iujp76pgp+JF1fZ7sippmsPIUqZXHNs4xDbClIjHtBbUzSzgOZfUD7kg
vgih/0fIFFmZ0d+I+y8oaO+Mp8mlij2lxRibgfKQ5XT1gmF4GDgm1wN43pqVlC/0
pnikhZIqpH9nK61uyikod3ickHUaaC17wTKXQgIW+cQLO/d4E7m/YvDTAn2nL1AN
0K6hbq4TVqQj1IlCkE/yxNDVCj9AEt6xthjHCx0Xbr7NlyIZTg5ws5jqqvhbHR5u
ph6sY8scTA3UeByVv54ZkXcDufXxse80yLM/nEZo/pFkeZwb8Q+8+x6WEbs7OedM
wkmWt2eDmlz/PGT1rcSX7ASE//jSfC6Sc1nBPdFWuo3hpQLQlosvo0/DBx1tlnNM
MDLgsqUsQt3Nt0ai2dOUYCYQm5KqGt1fZKC5X4M9pnoxGaKq/umadu1CjJxNtY5X
AHRektJMZl3uurZ+pmWc4ixq57VHOriViHmSSEFe0dcbwDD/k9IlmFKFI4+RNT6y
hZxTCbkXnddgy2PJdp1xtDcrzlOuMTYXIZvdBoPWkrTdHKf0KfTIKZ9Vt9fgGL3g
VGcA5xcy3N9/6kL5jJ/rtqNfS7kXqFAMEdKzn1hik/tYTKn9b4xxOOL3bOiX04K2
2VivNa8ROLU3XwPt9Fuwgp3SVetEvQtYcsQmvez8apil1OM8F0YYz6bwxWIKLYT2
mR3fpVfPM3oRzMWBYJMnuqSBXiRRN4G/BBg0IOfNelTMsSpfuJoo6trzqQZJx1a7
hcb+gWR4WG0EymJFGNUDyMiPU+izRj6A6J94R3ftXZOnBO1QRSqXG/ScWLT9vlX4
b32xqom5OIsOCbq9I8AL72/5+rOa/hjeWbnU/SFq6vMG8ct3kRCM2Mx7dUYv19/3
f0WNU17ku6A7sSzu/d+OuAR0fUOZXkrGITUD/6dxGS7bXG1loc4Tsgf4GEv4HcDk
EP3wa5ovPkSKfZniB69CHSRCcInhQxp+D4L5uQH1jUEh5diEO9GZgHWR21pYVxLK
311XH0ykFlIKLf75Sqx7Bi+7o72+Dye8zAes1B+qb3QrqDuT9nfu26Uss435z4wZ
xLKejmfn1WxwEEBmtcRFOERaERtTN//+eblmgbsHNPQy1iaGAq3mggf/kKZYMGYz
VCt8JghP+pFl5tBQjFCQzhxsNUM0/q5tQE6CARC/HqcYaJAVjtcq4iVbWT2LXUv2
gYDRThbICwAVYooQ/FtHWnYHuAsY5HGw1X+3uPSmha8nnUf0wVRCFlYtJQHXbzRg
qgIyqb/Ey+ZuEBRgCFIWRkMj6ellJ9hnqwCwRO8NAB/eNBxdD9V8x5GAAGNHYBCj
o5gH0sd+L77puAnNO85Wb972OV8mCdu+o2SnpdZIAIKaog9dCkZI7tv6mpPElyEd
0bCn9/nwd8E7BBEnaoFojKloDxALQRVvJxSLf4UCiYa8rz0YTe/IDXkgzXHmmbGE
tKso+rKSbWTO6cWHfdTkLPqx5mKWl96nBJMqQpZPsL8b16jrqkNs24gFJZikoJn5
h+qQ7LaHxFknNWoY5k3fYYJZHUESz2AnTrK/ewLkqJceoGFUuZLijEHZ1+rGKqKR
d0nDwR7Ybw4WZXDr9zNN2se46ajrTfWHBiH5dx/oQV+Ol+Njmsp4L8FHrZLlnLkB
SmW6qFF35PQhuliopDn+hPMow3uOiRC4KfBvXTPGUkIFVKHLe+g9Wmqm0dnlmhVf
QkkmY1LevLZXzQTE+c7eg5+cRJphCvQxKEvdogWnJS5wnoKLeiSZVvuKY0D4vZ7z
HjM3HzRGHfn0c3DoLMv6E9IJ0SNNx9SMrl0v9xE3H53ncc78xtDdrqyEce8UVNj6
KWeRTHoTuMhymjaFiFdWcEYGkyr2udnHx1Gn4XpB55bapjIxSBNkJ98nGaMR/Lgm
GNv9x39SDpZWzHX4eUSGw8MQ/GVj6+m3RulwUJPfq1cj2800+hd/iURXwJyew7d7
4OFGB+iDzzqs6t7JtJJBQTZUpu5NRpb3opzR1LJY+W/14JMQgPMr501n0OmOckCz
fKUSLmP2gtjGRz4gW1LyK6eywUL//TQXg7S+KL9gqK+tAC7t4KpnMXIWuZt2T6GE
MPVmhCdzBqSoG+BpY7lEzloZ5FMWHBXTOvspIGd35pcBF0y7T2EnacFS0nSd2TNa
HH17K0DltDkotLpxYZz9mzYdRQVDmKvCwQfSwb8XCFBGXKnBtJofXLYQlGiwZ3B5
+luLuATOYeUx3zPTZMQ7bP4j+NXl2SuWmkk9m8mpDgEMszompMgK9TcmwYdGDPYr
WvutqoiJB8Rhxo9JbKH8kNpb7ncOMP9npkRdTbu1TvxKWrcc8yEs+EspvP8NdubE
0HMxfXuWz0S0/klTtle8GqWDTAco/HBbhLkqiuciA4LPBmR9JTn6jVERVkeIfZeb
YE/w/aF2owetC6xZRWTA7cwS9ysxbC381FV4IHQBW5tgyoB3VS8nV3lHPKRJRPXg
4vk2O5X3JO6Gu2VwqrfxrIJbfnw1qfDH9KKMLC+yRq9GMZYAg4iyWfux9MXy2mTX
tOrxeh0YCdsRYC8Clv4F7DzAaYvgTrpIgOSOySiL23elv82FQL5LfiKppZEJG0PR
9V5xC4FRqYXzaTsqVJWoIM+6F88MjWfRteRd4vo6SICEURl/ULsztDMAznBtmPQu
L4CmPdYzjKGCiL/P6CIDcZ+WROEJn59YFfdm43EXIyiEW6sH30jrB0A0A5qi1Jb6
v/IgWckx0zd3K6Cxfq6DMRZnVzYvIU3aFH4YOXqY9gfZFyHy02bRKhkjwNe5GLR8
JXiPjdoHtYlig6+Nq1mI3YfmHO/uC0z+/JiAMRcRWPLUCyvyZj63TZ0ConsEqFQN
pxd2aU31rU3Pij1Or6sOvbb5xa6aEfmqC9D2Ffxo3rvKvMIBet43Z4ge79sD9CHq
mRAxYGBIgLI6v0CSHFfi6Yu/9rQoNPq/N+LUfr//nM5p78tJItdgukNbmrtnVjQ1
z//gR5cMcQugnQT7RBxx+Z+jNMMmu3m4EfvBk5t/P6nTX3j8xKGTBuQ0WHdMED4n
TMIMwFH2jCXG55eEz4kO2Vfbz1IlkzGtUhOEvUR5q5XxJ6ZVylYM5AW6dyxvFFFM
x62qrnkcE6nkP4DFXMqrDtOumCkqln5xnBLZ45B1a9F/F72Llpt2HkUrrmvuoDJi
F3cWUC+C6r8mmgUY32GBN+8ra67rmohPmKaqBQsQCSqTN3wZwYMcOIRjk2339hyP
gH6er5SzUw/XE4eJtdcS3l2ErPs4IPYGabe7BbVwhk1u3NB1BelCxdyybqUpU0pI
uHNT+RjHR/wKi6BJk4dLq+OuSYIvDmmuP2AcqEXvgol1SHP5aH4Vx1NKJEIgHowQ
aTN6SJ4sLaSWZEyAM7u+b3kRCd+TK9GNV4a2SS7pTDg6pdqqnDMfzDeSo5Z69fk7
W/SByej2GKLGzGJ0sp4FMDqvkrasfGpDwEzC4TDMp6ugGYZe3wUZDg5g2jTZnUGl
adjBSzqIW3MqIn/x48PO8GP1j9IRcVDFGSxoZkXyCS95tvink+QIT9cBW5Jel5oH
j8QT2WqRE9D5PyaT2cgI73mMWY6gZcC0ZDa5Nke1pUNklJwwjvmT8CG/222eX5gp
UP+cvzJDIEXST/P0QgVELlz/Kap1z7ee5AFVuHhruInFCbe3/iW4cDDcLtdH7aN+
h/NSTwSt3fyl4THxpMfJmDtdD51us6ocMZcdsd9iPF3dVxjGQXcfJ9fF0EU1hPRO
Krul8nrZ2+JmGOZwyoqUTDRLYL327ZtOh2Pf3DwKNMoQW0G09yGB1HmSkQV7+DpV
3EjfU7N034KtdBZhkZHTLa/ekRHSsPW1qFXogaQQ0EC+KdYas7j7JcdGU7DcMeLu
OEFFrepkBMrQv6tZBE3s9DcqeHFVpfMTBViiTQ+xDRaa5s2bdgIcY6LMPHlTNXdF
6exAJ63l1LZpj8bcSeStxMlB5mXZg2pEcXnBhyzxoSOV9cNiSYCcor3vXnj/lJAK
i9UY7JuPhOQUxVr3U4YXe1zoDaVXje/hE2DO7QNX+jjGvQsAPURGMKWf05gC1nkk
00xYv5azQ4XZ/Vnlqrt5DWN3ip6O9cHsrUpCgiIV+DwxOlSyqTgbRCl54TQhGvaD
LoJXCemWhraoel3Y5VyczigFEkO3buwKIlm7gUilSCpbVt9Apy3Lth5TwBXH67jX
rn01FenHjeL7aGrmZIuA7rYRoH1aY+0rNMiag9eeB5HliT3CkBDlgnSaImFOoUz8
8bneHhine1OMKGnpJs2tue+gR+k00QCv575zuPUSlhSlayAgElFhjyO/m8T4YiU5
+Y16vNMFBjB/pvqEG3BPZHnFKxSczaEFBuGjshq+TT7xx7IBOPN/S/ZccQ96bFjQ
JmEAy4F/zUv19p8QOgrEh7IjQ1vpz4ZiplqYAFOEbQhwjMyQJ7IgH9t1Jdh5CWk7
YTcWXpcQ93jCJYGjj447bpKgMitIigUvaeiOf/lo9l3ive9YsQTNdvDQTCPdWWQO
44NZa58qG8VZNh5XVT5HcoUyJv12IC46F5SJI/k5ss7YlI7hbvtQ4Mx6JLRdzAKS
+5GEjaP1xmY2i3JcO949wvZMVVwAe4Idc3PKdhkluzPj3jICrw9R962xtAmCJpCP
HDHi+XsB3Z5YusgfYVPVrzo7KCKuGjpIu0twu2+P65S8u1PfWptbvqb+3ojEneNI
245j28z+U9GPsJYyZzC3GaCo3t56cHa0cJlhjeJcMhH9wu/dItH1gl8W/k6rZukZ
LqCFaFcg/4z0xJJ8VYJq6KMmIFuvoCECK2rlFvcYPFeWp1oVzOoohaAnrHsb55/u
PTmsEQ0rf05U4wO38vw6m+5FoNG5Vjhb2kGZZ9ZnI6OL7BvwdNcPYNrUuumCoWPD
BvmV8Cl6N6LbRSyHo1kAA9sAizna871oeg1xrqEa6WXnpQKg9yVKvDVe6pc+YKTI
mC/uOcJuqVpy56puJxhMCghL4oh/fqRAXmP12U7FsdAouTlnzyErocwPqDlpZcmt
875CnqTw5lAzw/pyKkXmmCUDxHPfm1JrZ+tLtVJro0FGSUdgpZ+qPXSSvic+FOKJ
qlCAnleBnw/fvyFNZVwf5i+Hw8QNkZfxdhOO2y1tUt0aDDtwpxsYKAjTBdrHdYiZ
l8gmOlMEJYtoaapTWe1k9T+4HgJ4qcVG1CG3h45XX3ikOKUKmDmUVeShlQ7gbrBW
W0uVt64pQMvEopCmCwm3ZZ2qEK5h9y8PLudcl9esGGQl6e3+V2sTkx5F/ByRk5WP
cThpyL7YtcTyIb2sjyJ5b0JFLYl6gqVfUOARn6Nuh9U7gyW5XNsaNkug2ZRZZBki
JtfpPpt5zrwHDWZ8Opm6dXiCP8wTGlFkOOBHPXy/ZS5MzHsKhbvSz8kNZQCcItxo
YNkIziwjmoBW3VIkkWnhP1z2mrFLWza3G5piCvphgczMIFcK2pVh51sdj+yWHLYF
yQPmxwbJY6oExdUpUUP0j+oGZIl0hU4jmj3XtndsAz9VMfDk8z6FzY9sXdXAW3Av
qXQeA0+/R0dX7tFSgCziHK9sHrxjdoS49IufhdFGK2eM7gn/oHEBPYhTW9dXthvJ
EyaMUshRHFWduy+nDatnxpPsM7UNffVzff6wqMcNi0Y/pf0NNDC/+IBnrOF/QZYr
l+YmWA7p9UUZ7mi8mM5pqjf7+Fk/r7oAIBBRmHaemFrQ9usjoJ6A/jsLiI6a+okc
g2Earxt1NKlbpLd+1b6rcIGijD0AslAEuG+1Jyhi4xBmCwpv/5wHOyCWh8WyCMy9
0ay+hPlExY64+3D1PIY/3c8GZQ/svFQYgDqh/lU6zpVaI+vGVt3GV1MQTL3FrnCt
Zbdv8ZARrIwGm2vigrZZiofozJsr8g2zgXeLO5VWFiOEuN602uSjS/dCM+jPVI+g
UgoI+88uInTUtz6z3qzLpqsr9zrLWMnWWCWMw3QGxwVrIB5CdfAWPcrIh4AmSYla
bTIM5TnHV9I5jC6ljDXS1zcP5Pntqphb7ssqvx54F7/VzgVzR2gJIeUEQMGmdpaw
dhVHlSEIeegtRbYfMBPHZXOBgwI5Hg5xGazi4saPkmKo7ETceHzUQyqYEDsuSZSS
681yl+ErW35O3EDi8lbfZH2NP0wzMb93PIm87aXLYsgK0zkvtf9AC2DBXKl6TnFB
nvaS3UpyVU+51X+AEt3S2CPoTG4M+sLT65oiFMmK4BUI7UWVjgTEZ+h/mwMueze1
jO2tU2vogaEcI4YNFQ/ukQL8LizbEitTKWNtX/Bw++/H6bxQzcURoPg03pBb9anK
/zkKMAh4GAkq81IfwYEGrtq0va3xxQlzH3WnZyPdclX8oaZIU3bEnr+lkW497bSk
uyQepW+mlyelieUU0nJ2xwKGDCIqZDNhLnBh++2M5JlIAFEbh2NxuWJ+AKL376TZ
ZYU5YVZ0oDOAMq3yp0jV32PgoI7YPSdvGizZZwQ7FZNBquGRz2lUI8UaV1/iMjFX
5xG1sRA3bv6r152ZWcrCR3zROMON3zVN9DCAdHdYEgND/JDgmnSzvi8eXMOfuXir
JFzhsdKuEONPznXRexO6/rILl+qvSpMsqdKMB1GZIDTN1eBLSpBHBqbRXyGy9dD8
USoOxf+55xNUVAQ6w+1Fvu4qK8SJzdrSZ6M+eErQIPK3EPCVntDh1rZM7y7lSHoa
2aD92mC0Co5Ac8HwHppZYJBbeYfeD2WBWiA/6/b1yH+jRs470AubCpe8RHpLDRxn
91CjhnLlv+/57TG2VfqWISohVHYz916oG/e5YmrnyW7i8mfytN5vvyvPzWv5+Yag
D04fgeH9FihhpkzmeDC0bVmzo1X5vZkEAqPBURMQhRAam41evFvn3854gedSWxK0
kAs/QCWIfeorrE1rcqSkq36pugkdN8/W5OLzahYbS70mRmsisAcdxQl7x+rdL48+
3LR+jzY9RxtfCvSwcA6vzgIa4gULYitGTTm/9Co+U5fsWheBtClpb26qc07HIrVS
mYyuHiPaCHhI44lNAmpUewqxyymvUO2McWTCYo2ZvrO6h4WRwb+LkxmevXku27oy
ofqZlQY9GjBUXm5aQnmjVG/UFox79BRqDKTCkH7fvizhjpYKhxNDM1Zxv5b21Msy
HrIjFQ5ppx97iUDHcGclNtWEdKZhyoB9KSmqwYjrv3LM4j4FUKACSxovM/sE6Kr6
n5BUtBOqlxOSq+uJ8LPImKhNy9KrJBKY9pHdTqCxXTr/UPjQ3qqEaRJuNQ8CahqJ
2ceXJEMuJe9HAoUhXcgRLdaG55SRfcNd8iHRQVRmM3y/h5w1NvJ3bVoFZ7Mn4Nbg
m72w38EYgLKq2SZRps3v6FljTNx4LHhL5y8YfqXb8rtyN4K8DYYCTCuGhOP9Kpo4
RVOKWc8bmW9Wldyk8QcKcg4EY/HyXT2nOis1yJBuPyWSYwaKGNRe+s7yJg27VIdf
8QXBut0a7b2BXBzO21CSel7NCYmR3gKTb10Kf6QTlPoWK9593JCBUjZyMkItt/A2
ZI4zUg7assOXo0Y+e/4BnRFLeW/Q7A2rjXh7y/g1FFoGEsYZoHSzYmUq5Rq/Slhq
mt4ISQneC2ILhK8pCCiku+JbeQ8W4l3DcFd9lzItEYIq8jkSrCJW2Kgic0uJzlQw
RD6mTn0ufrkQNMHYGIJLxX4qgn8Qmg5F9eGrRK7sd0qkLeBGvLPZ/zhozVB8luQ+
rj/hDGP6TMJKmSiz+leFay+qFp8WXbHymj9N95BgG0Xfgv+572/XBc9bRvK+tn6V
IBD5IuLmfQLoHHN/GWH9NXVFqtggST+p2i320Uv8ipdx3DvBB4S7QoXvPLePU1tX
blmSGFWQ61zrGbboJA9x6KBr+cW1iBvDauosLiNdscrNQVS9bYH5aGW/0kuKCsMb
EN20szn5pvKcTRni1biEBbTkC6/Gs/0P4idu5y+Q9dBNc2KyrRufIhPjEdnGmn/9
IToMZBFxdKMcCTYMx6A52HyXOSdG8qYcfLueisQo/WNusugHFWBgZFWHZUJ13rYm
NDsDBhhr+26NcNb8BtWIKZiZakcto7I0Q3Z0z3sOXv5cQ0Vsl029R12QQ8V8lKzQ
BccPeFuSTKfW7Ktk/Sa+o+npS9vKX6+eN7LLIoLPmcVenpJLhI+28Q5QNP/G35m4
E0kinYOa2f9A1Gr9BDsSLL0WvT2Cmrwtvg2kUhg+/CZ5I8a1CiliSZnE74mTv/S2
q2O52QaKZULRToqlmaIsRPJb7zmjVtcUAkLP5JBwPhKpJ63jf0Ixsmt1M7hspNgp
ptkbW+cKQL+F5SsvRGqaS+rYzexy3sXYluS6JV54OinbeAiE4yDj8MKPCNwhNz1I
5lr8OgVqr9ztMm84ViEOUQcxcWECP2nS+2xR+ajnm16LKhI8kz3jahKjN/2yfxTp
NyWgXoTBXf2nCzKmAk0jm52Vtz0oQle+vWtLzLNDb4VFJThluLVEtExgcOrTvZ2q
tlCttoQeVoIJlA6OS3eRlWv/Qu+4qh1xj8SJZj5ye32EMfOWkvjB0KLtbv0McpAG
H6Hq1KsOpFHp29LL2tijbEQ2tsEXgTrtfRq0jhpLFsngexoh2rB7Foy/B9p3/dxM
FnUAISZFy8/2pkkz4XZWfoH6egcHYM82Jwt079pJ0bRc+yfoMrvsZcKRJ0FCOodS
7mx3ipoN+5bloGGRNQbTDdOVYLg5hIO3gDGoZc6qen33RfJBfntKxa4Gk5wQWacM
VQuLI4NCK8hGrdwvwB9Tq4dF6Z8EwhvUVeHTW3D6nH8o9PSX5hafiNTxQqfgK0eL
uU2Gepcl7CFC9Ne2kNhgack4qo7eLL9qODneAY7o60IFSns2cokyvIuNwM+gWFwJ
r8s53/1ZRtm7YmEm1PfEmCkK7AvTytsmujYyz/kLStPxiDgqL8b/XvBP0kjWBsgh
gi+LOsYHVyp2jP6ulSXtxt5IjbGlyMtFskoiob7CjLCIzXTbDoXbbXOnZhwmB99n
Vregfp7dmPgUT1I1wAxzocwzoI/catUCQYky+2YEiVPFflbo9/zs0bKUw47h3AJl
J31r0rCTdbnDacfEiINUhKbLzIuWMP0qefhabeyReTJJ2fQ2PLz+hHkG0HnyuRw6
sT6uviF7PQ/TXwNEgUMFt0/oIsWWqKKCtpdOOo0X3emT3Sz+Bg5EL9mKazoF/zAN
vPTGR/7MbmOeDdKUEYd1/1gohQwvmYGswIZ/OHTEP2fClUWSXP1FBhksiWRKNvWk
Lnl+xoXItTjKOhdYupFDsM5SI9ARK3Z4HLngmqVmuMN0W10BisDw3+lwhBfKbv6b
97XcdYt1v3cFSlHyimoxHIJMpaK40D5lnh0m1dw0xUOvn0fU9p42d7ex5hkAY2Bc
8E43Mzs67Pa0L1SEZlUkFRGiJ0xwGplUhkOdErjsrHNtNFADBlMYCSOf4WWGjOEM
3F91CbGdgJmfGftKoYqChfOpZoVxQofSlYk6RgyG1hbgF2tN3jzMPgsKVi3TRMbL
cigmfYmiDzFSLB/CzVL0cqnlvZDidSOKZpVepb6LwJDqnwySLSoNkSBpQPLp07En
YPrX+piMwpUNiOBW9FJ7W6ZgRIEIc8ug0/LlRhO+JFD1R09mOitvWjJiTwlbY1Cr
ZtyrhKSyEb59Oyj/DMTZZxwbnxOS+Ggw8ReYOsZvBIaeTW4m2p7/kXqTNLglGUBF
u5cgP2PjADqW/wWXoRMHFXK6zrjOn6fQLPc5hRBz6/vJj9eDwkBYP7uW7wsHMeO8
j2i7NaCljetCCqyVuGReG3Q+hYF9q2xBcWI5NpwImW8+8tRejHfCLcCaOzqekHW/
W45jknjGTnaBHmfkkXlhPJVQ1KgZiKBuAxM7GjzQ7Z4lygZC8FJf6fM5kgAH/eUj
oYvhSRkRiEV4+aI0ynbMQLmmdkMtjJBsG9/TTzPcnbkddbgKhte10XbcfeWasjcU
7M8t0yQI06N8ZU17m5Pf/48VU4yoztDrCD1wEOhlzv6wBkJNj1aqGKNbVZGt4TXr
Z0SWeU86hH+3+V9c3gBZEvAqIpdCcP8xhadLA2GUjAlGPZNzhyLhQrUTdFb9AAcV
NhhhK38iELfCy//OQNDRSPmmTG9JMKLKfvwDr62A/26uH2Qk4wVFl1ywWZt0PluP
MvGiUPfHCj4HwzOPhkWds27/CdXSD9SZCBBKdH+MQLgCgnU1qtRsNUTqJyqW/QjX
h+p9D6ocNHUepuPMqW0wAJUfRPNT0hgtt3LtMCxiXHTUv5XdswiDgryRveENSiLQ
PD9Tm4LztSlPZgx161SfEDYsIg3Tmm6u567R2MvWgdQemI59qxOjeoDShhvL35Le
rOSee2N0nUoUyrw5VV8B01CcwPYaWOt0wuuqhs03+KgwjoEFvEI9OrObSvDPbxP/
sGDNkuPMqau1jgPfbdqYoiJYbOdXEglQeVihpg8+UW9Sq+ZgCseW/HRrCyoXL6dC
CrIQ6ECoPohwYh6rgaBT6XMGIMxILbdqfsoxFE3Fc337O3LndskEJYs3jaLXCg2r
J9Jam1yJOdmQgPpdfATpZQGzLxunHL5tTf/KycLAPcCwf148AaM2SpB1M/Fj7XML
PJZleIXEUca7KsU+cjcIRBMgpsUTSFf/YYFmlouIahn9fUcph4z+P04Y7szyB2WD
SVt3eu3qXIkiF74Jt3/eG3Ed6xa7cKMt7RXvC+tB/z+/VDSD9JGq6GkTgWSFcNlU
tDRjNOvOq3X9JZJfUoRsW/h3rAONGy3ejTX2bTtWU8RMQWsof9DuGfR8Gq/w4wKA
VEdTTqUuGy+9G64uZ3KSb6870yjUg3peG+vidPKhUKUJoxArSxJspWax3k8qRTQW
Nz+c/nvwLH/P46UIIQHlmHlQE7eyMa9YCBoKSVYnRx7n31EgWtOfFEQ95zGr1Qi+
QsFs+v6t+wUMBxd1ZfmgHgmCifnfmCbT8ngzFrQsUrtbF4Qbtiq+FDmM8sX5rw6t
mLzwpmfm4hu5vQPKyUQfQLv6LcAqVmHO8PmXd+m0o563Fxr1ltYMzBmqeT2AZX7x
Jp8A5sVF3/Kx9roIPpquGPeeZCgXb5joGxRGH8Ek8udZk/kXdkHYP1y5pmbnRfwr
ae5wWKdSpFW9J3Ukc+8Kc2JOvVY8kJb4A9zY7bpPLk7QJwgKhXbDyPYBv5XAw8R/
oA1lVWEUgDyqdDSIUqQ3aZvZ0KI2e/OA471pF+nxjc3hrWmBkTXLnqMqc832HBcq
qC+F9MmARHACOgzl2EHL+6NCnGSLjOXIKpcu6RAo7UmLej7a9EQHiBRgYyenjUgX
Cl+2Zf5sXHOa7HUxD7xH0Y3N7dahhjpA3//jdyLeSybXEeMScuybXMBRWovfM9g4
S2Bmgbk+Zpxfeo67yUAcGTewDiGtIwsVGBjgFnyMK7eXk7y8sDU0Ish/0/IRd3oX
asgADprsGvJATAMXdKkBzm8g2XHuTA4ZtlXiQC+1hDgbsmjga+mxadk8EHA8kapk
EHQ9HMTPdj+2IEvD3J9hHwbhbggdAG0IF8c5l3tkc9lLpIvJNWYKes4mNPYUB+14
7Eb8Kb6iaJ/tBZ8kyWj4jF7ajE9NRNQRW7yBTb9ej/IdloH2XEBmnQyDVVWj3Rr+
7uhHmULm4gBGcg01mRXQsgVJlrR0xz6Qj3xkQ5lg5/68J5t9euAnsmPS2fVZ/phQ
6TTG+z6LrDKVoLVbMXOjQeuhjUwuxlRz30LxwlERdmUbHnrQdnsjtO10VVKIJOS5
To51g2dFry9rmh0H2APtL7DHHdFJDDXoCvZgfkAYuAju54TUwb+C9URYt4qCoyPF
Vnoeb3hx7disN4KlpfRcyVweIKMCBs9SI3m6gCIifAjL7vIbax3qEAd++Zyj/tYO
Vz2x9poOF/NRN1hRzp8zGdoPZaif/TiUPR4olXwNJ/XVI2bgHCjVl04cbpI1Dv4F
tiLzmr+MtLOHU1DZpw/po4K0Mx5VYctoYCXMv1mF1ZzIB7uVuH8LyVHKRt3k+id4
ROB3Y8Byi81Yl6DyQ1NZMIPzENFM0hFw8RnIyeCrKQEfLh/1YW7koDWi1uKdeogv
6JVy8rz9OlfhNdahMs6JYXy2YqjDKHcikROOH0mearx5fel8jqhwm+9BEWw2GXoG
5iW2cfWLn/wZLgvoA/Wi+DLonjXozHCYdOD0oplXKlQ8j9A5M2SugWYKH11qmCzk
dulZYwbN3MnV7J2dhZgClPXbxWNR5GqwebJCd5VLsi+1+bmGzv75iOyIk/eq57vE
WWzfafjEZmfS593WTG2MwH/9iC/H8Py9mNgtgmJ503CKsm5YrdPwytoC85ARwoG8
N1Nj3n7EZJNgt2EM5i1dsuN1b6hlyx881KM/eaYp+sxLnfasdjdWf9kSsMk3gD2X
3ubPcwkReFKks9SE+fRKLX7BKDOugZ/R/cscSFz12kbZZhKRWXJM0A70rrkzfBk9
C1CItKTdAeEwZG1N0UkzRaK6FUlWyHvdQoRqRrmDuMQBaeT+9JtiWKRzFxkfgR+Z
e2232fCx/fkTgoxPsiuS7R8OU2PPX9ex2IrfKdWe4Nybk2CVRDzdjGaYWbNKBWR+
HuxaG91csle9aO3j5WaGov7cceBkV8lmoCDID4XCdJAd6CIYgrZE2OiZSLhSD8Y5
sU57+zXYUozU/JGjCr6A7s/kiPnFvUlX7TnC+8WgiJlNOHPdVQsQeg6GvtGxyUvo
bl+WBg1ElXKhkyIuP8Ug3KctoEhjTTEeWOSZW0LDscPBfXXUgkUDwfZG1qFT29q9
zn8/EQnjzyCtiZmibHmUaMx4UNDCyQ14V3Q5zRRXXCoWXCP3wKg9zQ451N3+oWuH
HFVvki01dzecvDsxSTjvNH0kDjZpNtff7hOHYJKaCBLh97JhhHWlcRUwy+FtUxs0
uyFtgpaqLf8941A6Qv9kD67/44rGlbqG0Mx1zzefukfdG8CUIp3iSnBO9Wds4gWZ
mvu/MuFDlRIADoe38Q2Q9skFewUX1c4tl0qlN2nsW5lXRGxzv1rYenJAImGS6PiK
K+6ac+n3/6QQXBdz1NqS7yHxGiO5QDOmziRA9Fifag5zOOE4GivkUwrJw/FKBcX2
ves5NKVL4HEhFWcUgrPaf3cjxFJpesRhFFG0mjBzKcObKNTlfwbCXbJ74nlx5hyd
1SSQDYl2FzRSLcter4jvehST2YDUYAH0eB0VFGSOnzVAFh02qiLB8lkXxcBFg8lG
gBEnNJRFsbcUBLk6EdOaBMTrK1Z10B4hBDBVZSSbTeAEnmy1qGXzD3jLqeoGwhRW
UH/rfNOeV/5UNhom1Vkk8QGaRaTF8sRTzo8WRVPKxvH8Yb4MxJMmqR8ZdLzeJ3iM
0RIGKy5eHYhnTaJWMaaELRA4wLyfEz5S974CWwaABOyRXVLcbZE44VaOqXxtGT/p
Ys8ko2fYUT6pVwOK4zR4TYlCFQxFGAVlaPpihulG8ENJ2iWbQLCKF0Zu9hSwJMJc
x2oOJx5I4Rey12xQNDEJmCGeVw+ZcgB8p4Pt0GMALDJ6eid/wdxsRkuFR/tVz/f5
CnevzYzl3A0nCNKjMgnNI139SK2toUBHLXNPaOxjwY2mD5b1I2S64OH7d3XJ3hJz
TvdkXqOUUAC4bR1YQ9odyOTYTvJXwZPWwCBqq0fRh6F5Ow6OhP4SK3O48UN2wz0C
n12Z7O+muudE2dSVYaUHGpyKcgT0BT3ZrTuGwq2U7VW70I0syUi61XgrO2A9A6IF
1rcYOwiAbOh59U5tppKyF4BuJwMGfXFnwuxjmFQlJcBYEyHO1CLLxjyxaq+NMmtY
FCn280cFUuiKX/SUBg8JxiywkBNkd78GnqoiVfHvsO6DCkeFs7eaQuNJpb/iiNvM
RTKm3iSBG9jgbiNrUbeHTAmOQKqVc9g102vi9Kg7O5bFlBh/cx/KMM/rtR9GZzNm
bc5xBhqQU90rNI+yNKlh8MHP3pOJu+RQbfOntebcWv2jtav23GWZnDOLFAV3xB5B
HTiFLyA9qzoQ2MDHcIblWbuNq5g592TX5viP3O81+EtGSK2EFK4UjPZDxohtzQsN
H5tLrYBenIiKr0FobhKbo/Z9WZ3t+swug22HDh+PqIi9l5uFZJqbXASeG7grm5BO
5FzhQmX6CSiKc3W4alKOVEPGf7mPS8VUAjobFNJjOmRmwAWn3d8OramgU6pbyAId
7iK8oNzkjeNAHMIcGjurW4i1e0yLzlojkWwx2eRiunI/fKWUSB7LSeJdIqZBC132
hP6v5M0E1EhB03jg9QT6NarsqXDQthU+SGLgwaiOPo5TdkJiDMvGOq6bwIo6scOk
ZJRtWi468GzK6w+oOuWuZ418aUK2XFGzxKTAD3yrR1VlWTKWY6CBdVn/efTMzrGh
FRbcTIWmd62cLFqB3ui27zt81HG9OCfMIW35m13wp7mLEIZfqxyWbGZwDOpj3QOx
VwmI/96jwV86/WW3UUs4T6tiKuBNjXnaOtuoH+i1W+zLofarqrL5ikebmxRECGHf
iyC+BvCsRUqOBVdbb3I+NryW55Xsa/mdzsB4VPkTtqSCiPpvXBEyfX95yyjsAXwb
jx6IaP5Qg731L2knr1YCVql3/H1hgXSJWRTKz0LzwkvPpcZcPiQWLs4WQtoMGL/2
wrI7yQArM6CN+7rrzYfkkyGjC7ePM1yq5e8H+0P6NJ7iAJuWWx2XABMPhRO2naKq
I76pmNd2VxVIYSEP5H+AmCql9lxCSWC2td/dSk8p7lfaDZtzOaesUk2cUBC8HMZ2
lU+cp+jDeKg5JBYFISWQEeQFgWKsfWxN9inl6hqFMrDzXhwHMfmIkwfUABe+juQF
jV1RjcDXo5255Xo2u/53ah13zZzF0/13kBclFnfwbTZbnc5GM1EEbsiqjPUiqbq9
evAriQjJaFw4fgGCiowuUhEL5QDVKZum2QjRBt9i77xZE0nhS1AhSEoztg9JdBFI
MtaIljBFpVPUzAxBAYjLqtzmU2z4DQon0KHS2Z8SAi/nSlHxmPEebGjze9mw9XZp
7jUmgh54jihH4g7PypJJuioTKScLj0zXSVKaUckdGlsY/NSEHe1hkQhZpOBAWcS1
fPRAsclYBZHh74FFUrZdYohf/1nlb64dbN9Ir2sP6Dm2/k1XhXq4SlAQ/ouvfsCu
dXd+3lhyiMR4ZSdPLUysYdytD7546BpKJ9UIMhtB3tCBzNV9bWD8GtsUftxENMqE
DzE9LG9FREJ3nMMyqX3dD87dqnBzs7bPkWWy69sHdT+cD2617Av+pjvIor10tWZ6
XAR+Sz7gH5WjUt6zjqYu6APVdR90Sd4zaOSdNp9w/Swetx1ZOvRRL55IjlHdbxuC
C8f5eLy5JVvMFlWY5FuPi6s4Pf0aDynvcJ+M5RtAua1gb+YMsD8eFjForcky48NV
2x4ixrF+F9Mh2Rn3PTesA6ZtKygqMaC9dqDXRO6tixTMhq/j93ZCwN3P8mqMNEMK
ef74e2ClMm8wij6FdwUuvJxdF21lUyQzMqlUlRrFKG4auZ9EQOumMKJniLlhG6pr
Ku3AEFreXRgQu3FRTVOkWJoTHbxOKRl+0IByFp95Yi5q1/8J6dfm2wLvVhgSteOh
+DSXCHS2/ycLa5FH7fPa95fMfflinUdc1hGPZ5iydtFqN0E60Uz+iq1cY5QzFB7t
eVxalmCkF8D+vt++MdA8kVR90MNXEN0oBznYwDxPlCMfvRsGlKyzkZlOokyYK+Hu
V4Mbmy5OcMmOWSrSAiXI8x69s963TAfUBJuYYnI6Zd4dKpO3stRrvnyds6neenV6
j4g0KkP1UF7bzI5mjl8A5GXUIbEp3PBmiJil8IQmDKVUKE2+eIm97rdONRdH/lV8
UAz/96tS11LTTZOJD5igkOYJQjg3e2SgKyAMYpnYiJReaQqLCsNLeuMFs9MWehXq
03B+Ksm+36fSVuXzH4ZP6O0vGhqKDqdr5ifbQHhcH4LhiiaM5h9GP7Dy5kwc7vaO
Ef4j4aXKPUf1MJVYw1UziOALRlnfebzZvMnkFKvqZbxqIB3nNya1jlA+cUUApnl2
kVvpDyNJjyGOE2yFKR503EKJocyOVdh/I/p67tta5uwgx+omQoXh+LSiq/Yb4Nkw
AGxbIKRYhsG9tMJUnz1bvMD3VkqzOrphnNhWN2ThLF1/Mp7x+kG/YWPPlyV+EQuX
9UzhZVVKhYuosrk8gz4W8hZSFp3T80wEDf8lVNalt9wnDhIxe7dApnhNsQD2p5dn
Gt2Bgw9C5X685IFrhZ81NRYshVREyz4Qx4t1lKXaWenb21gqRV58wNraXmoMuUr8
EqXd8habl0BOrZ4DagnkcllZRiQhhr3r2BfbHUsq3j9USTai1PmQCEYFUQ5yYpab
dFVPhaVrOSV1oI0KOXW8bc0YFHxKOzUd8UBw57yNr35JH4rGtnrC6m2NVzVl9LKO
E/e5dR9S43OeJ1wsPRrYL+9lmiwVq/Ib5bd5kNmqszgmDCQ+0O3V+Gs07Df6vpND
xFgjRIStMR1aJk/8U9kEXAwaPcyO+wpFDW1XXfT1gn8V96oUEf+PFDApzQzlNZZm
YmdTlX+8x7NempQtwqwMW6hsM2fpsWNGA31S8z84b5nDSGhFHBwt261nCNjQyWa2
nACRxtmsLwhpmwi6L9fE/0tMRvAgKhhaeGIdc4NJ8kXyCJ0u1TaVG7t3rR0qie9s
GVG9RFapJTNHKiki8zr55OtGX8ISBzCXKcJBS2wASHf9n+JgA7z6A9ZTfuccRlDA
ABtTopnmzAeQ3189/imoQdaGLDA8v/5CUdHvAAiZbDG7qXqsKqGxW2SJfK/USL1y
AY9e+GwvA/jdWoyUdoeW9hKBieE02ZrBxnv3K5ohVq2tMYHmmRq/gvMp4UROAw2K
ShuILJpM//a7R+OHfCYhrD+oIlDTHtx21cY7Snu3yqNIea3oV2uRlSYIpuv3tNJm
K9elDFYqayFePlUw6AgkAGZHKe9PsmDNJ58+3C4R1FY/zwTOKaD3IqwcvjMWI++3
M2D1ryWazGYFrO6FaFYTnrO9z43ob1rXBXjRystNeoIyhv6zOuDgDzx+79qtXXsh
gUHLn8zVyns3QMzcf+AIjCFoZ4nJYxZ/4b+/snXsaGhyudASt9XwVI2Z1dii7UVM
a4WGpIMaSJG2hT09ldE8nICLd75p9BzuP96PvWR8JWaEdJXfe2oLWs4RWYXJvwz/
xxDoMl9CbZ0MvTc64Wt8kooXlir4B0G6H7Zc6u40DIVb4xNxtYkNSYTpKwzPq5M5
aDw7Gh/BQ1MuWv0xoeeRtgA0/OrvFN8rLQYcmv+RPqYgY0ZxYmdcVE67cLJDeLl2
kRn2gcbUhCshVTjpUdkGBlJFJ0pMEOuMStGz6wB2lSjFMIiV9SUY35yQggGgczoY
uZG0bMdmzRchBmZxrEzrjQCbBxCp1WdCwsHi/Zd4noCHXBtwLX2PfehYVd7M43gv
QTNtiE9QlcmtRiyR4oeDa9FB1uNACgCvzEPJhgSCA54Q4ofvAZzKLXAtJ7VJSmAO
lbptllLdvkC3hXlg44/s6Nv9xRCAUVdLfU5L/+I6eVf6DxwVKCpFYsIM995stjF9
eqqq27iWoKgm1iaD7P4eRhAwsMIcGqVs7yjq8MxphCLLxvKkaqRkwD5P//NavsTf
9J+Ttpp+jL1f3M4yEpd7HieAtqAS2PdiAySiUVXWQWjpVNzRYktndYHuRd1s1F+U
t3stsbD55kRl5EhG/qW6FkOOox+xWns0qPSchbu2XutIdsRttgC4xOYPEl6P/UrU
kGW7EBXKtfe/6aR3U0tsKezzIxACh1QuR7j15mQaO60P+yCGmuobmMUgT8xkaJQP
8LvdY57+jnNvGi2MR9h65WZyU4ozixdXQwxmE5yb7vBKaERI1RSruKFGwr81j7EA
LAPGY2VvnAkVmoNIvfCIPSsoVy6UZSc3E4vcW73mtoXRl5qDHlYmryKac8BYd+X1
RKATqKWcFFfIc6wbplcj6SYUK4nPr4TCnkD//teL0R/fGggweCHU69w4gWo0TF1a
7ZkvJHVyIsc4T0bV3UPLrsDB3p1eDlEjd1RQvlqR1pmMkB9GVFjTsh38TiO5yxi8
n2uKGufrEHmnvzm9BMBt/u2js29g8LqCU17ZGK3Ia8sBoqXsm+0lGnrYsTvb+AD1
B1K1m/Y9ZjJnG2pDNZ/CULHWszkbHIM23qU0Sm+oviYMX8UW3+M750/zcnhTWkk6
DfKw27gpIY/bqkfq3+W3PQsPZCqRumC2dpF0747zcezd5zuUjebKmJjorrUEshR1
NgmtwRK6JNaoPHws+IROW6pfwd5GzWj9UwgK4ZRFDVS2V3su6m/7RiEWF4AgvEbq
I9UUQvWwibtXjNMwuw3kOoZEZ3Cvwx+I1IYNiYH4AeCUq4SL4KxaUVv3MTtNuS6K
cwvyx+HbEnCbFAkcOK0khKTAF7xOODecFOIezCxvwPp1qyICyH+Y4DqPrY16CVCV
/HTpfpJua2y7Wr/eICjFDwjnenC30pWaoSYXQ6/Oq93QfAOk3dzAZiCjmXun0H1+
WmRgyo/ccOijbwy3k6jsx01Uy5Pm5H7CrFlW6DIjlbXYPhiFBcriNEo5X24pLfqA
SgFG9Mu8qpt3ulf4HCM7uFOMvPBEBA/3zF38yJHjqEQ905NewUH2iuoHOb3aoxEu
Z2fL8AaU8mbLA1o4zYVltTgvT1K8iTZgjnZ8AXezRp0bmSAZavezVJiL/0wlep8l
AVPFHVh4fVr8WjPOBwnyx6Ox3x1qzMk6gH5sSR6Fo3wirGUBiImgnOqOnwem61fP
PTsyVyOFav7h6DvEwzHw369/QbBGg/ppw22ArC0DMvoVSZV26ugB7nSRecsXDgy/
K4RIPWzDC2XDb1wfwj4BJ8yTVvtnBins3eeQSeZ7Mvet1uSP2Ai6oDN4TLBDs1GM
HyoPrcKFi3qzW0tsoj17ghwiN3M53czeEyCaf6zwnMRllIWC3zd68Cm3PqcLwHLa
5Hzu3eUe43HwP5k6T9xq5uvIblGnopKJkh9zeyufA6+AIRzGTZd/pJemxdMvcAmb
Azi88JboHZOijSw1UWGU49D85ZdjP9yjA40qY+wkFXOnq8YLnTk79RxqcfMzD+mm
TDddfk4MVVbKtUyzmb3wz+4h1lsAfwSKf3dnZrX5Al/YSEo9Jt+NBY+h2VDjgBS3
5SU0HWf39IuM+Btlpy1tH31P8WEHm83Si2YO9ZjhIu/z4ybyhqcQ9+0UGEDB0r7/
MbHEZDFPNbPXqnjEKlVw5uC+jbXfePJiYlFuY3yU9E77n4C7WgL4JakyFIs53dA0
w7MNpCXdgAFSfelOVH17/k5OPqa/k5H4qHmjB8atkcuGlS7Sjg0ofXoYRY7irS5O
FP/mHOy23R8e1D4dz+TY3grRVc9nVVjjw0yMhq+jmvAGN8yqw9G9NHcDWfdTqc6B
TMH4NNNHzwN7CxC6ko9LSRRi/s1lx27vEc41poY68sobvO1o4n8gtUWkTwigkErj
sT5NCdUi99B26a3mQrQFQjrRzutyjH5K20xtt+ZNuoV3wZNsQ/tcCx38hE9Zq8n3
CW3169Wuvw55cBrsU4gi9DCyDCHoGnSoz/B0m5MIDrPH7mZtRv0VCB0rI6Z6lc5G
qdNNVZ7oSDcPgeMDZXa5tLRobsqshvz/9Cw+adRVVUwoBai/m3naa/e7auc1I2BI
JqYPZbY5x93uWx9TZSx6Fz0EruYi1Uked9Pw0yk7dtMilyqqSsUGvbU5XanqUYjz
3XSuuITabSTDf78+ALsxIPtn23yVQMn16a0LVlI/e8+n5Tbd0gvSpnwuhjufRl42
rON0WU7SN0KNUyXSkWrHyQfHxATH3lWtDJ1WcM211/4z1dzYvjEmFjg667T2+Sch
W1otZgqSW3SCSe/ETTNrn9DUapGSbA1L0PPRctven6En4uc7fgZwGqFz84HWm5WP
GxkZoYWXWrxahs8oN32jbXbZ8RprqJ1j/nB6OboIX1oubtCCoCMXcw73IFmFVePL
EQGflZ2si0VBAmIPdnsjc90U9W7yqFerq2olrzS0YEcIZC/XqKiTnaDNwodF2WjZ
wKWAomX4KqcNhAspR2mX7Kf9QWBBOCgZk19bh3Tk5TZZ5OluNIn7QQbRZHe3O69e
MU8qBb2vHunjho6FI14El8pkweAN6G9oYeqpQUYpstmWAubPAoaAxguVQMykHlvu
M8et4fIl2RzghmEfplQNbxngOHbh4FZAQL8AmEkvnKCHKt23eMTl3aWO5Gg2jvf6
CEbBQfA4NJ+hALfV5zAD7CvTddygPiWPcAsPxdxzdt8R54V3lBeSXl4h/edEECzv
W4uq3/MMnxh6kLQQWkJwqgMbUGry6JluiQtoAD+XL2kI6PlNid32kXBDKATyOgsO
eGNPILjRY5gZ6OIXJStv61QhVNpiZgCD6232Lwy4xLUsq03mEuz0ChThEKT57ZHQ
Fyzb8K2BJ4IgBg3PRw84as43gefPOeTHi555dQSephuIko5dM//9inQl5/bSn5ry
71BBfU2v11wnxpZZlwiZ0qlgrcreuzx++eksvddRmHMR0gEsdH1rzusmWQHKyT0v
OCgn5+xkUvi4rr4Ks05dV86CFnp4m81wiZe+op4zGCnBHKwlJz04j6zZII9TDwsQ
ABDzNqqMthMwp4WEgkWmToS7c6jsRF9u+NuVgb147imKylNB8T7KbNoVwjPeAznu
TMDNmPYI9jAHjYifd/4dAg9xG8vDUHus84VpGwlrevcIISJdaG1VQ/rBtRMwYbC/
BXdjMQQJODRnRfyWqMQnNGb+W16Nt3iPP3OZ5dQcdhXkArlfDn/HMh3K6J1qlZun
3hoLl9F02lwvZ5mORfAyr8igE0wN4tJaOWlFJjwGLAzLpcgTfQGjqhmCSlspeIOa
4PEKREFLeeq5ndEA4jYkv/qQIuTbsdnuLJ7HcwAZXBIbOl6ricQYjfMeccOoPRy1
Jjc43gpGMxsIVWAK8nn7Jsw01WaRn4QqSnez4z6wKfE82MVtl8plNs4Gugt0l6yA
MwUq31cRlbl6yXmFYI6UmArBGqlzjR9njC+KoKi/2C570Ebu781B3LmExoe0eSJe
ufyWBkWim3JRxadlWVq9opU35Ak0YKu6HXnQUh3IYTO9BTigyKpVnHMm94qJmcFD
xAlY4OOjzuLvcMFYde1WP7ppPELoleBhFJ5bXy8F06orHirtICplPJbzuCxSG4id
HEJ+BFistvVd6VILbdow1hacbbpOaETrkJYISFZTbuGWREbcKcSG8RZtOLYiP4pj
G+KnZc0wEyMXteeI8Khe+kb/7PdF6MhkYx4dmGEiQBI7VtExmtFTSqYMurGqDYgN
kTsvlTH4GXRSG+g67RC3JletkUyGARQgnpLs8aj700oiqdPy/tTLusgt154L624P
LD5arufo7UrIzvlALq9ARdQTRkK35BkS2CQTV1i3Uum4dbkvRpoLiLe5Y6rLpLFk
BYZHJK7qUuCh8siMNI/nGF/jXxuB3AbkDQsEMs4B6mshIWzdhE6pdH3Ef3iCGK3C
PtXX8cGaITjHVULrmdIvFEBloRJ42R92kw+lVhBrFrkX7zJKh8Yp/W9BIFXIckKu
5/Mz/WpkLsM7rQgkM64VKpZ7d0Nbj9Vfuhr29lVaSIFNUTQ3nYakQ2EC2xQvvgMv
2CsaAt1/fXYmR2cGMk07LJmfsc6a8qR96ugh5z8TsvxVALi89yrP77oPBWzoKYGK
ui3IEDyhXM+jWcp3ohW3LlbojMRl+H/VtOwGe+os3ael7BSucKpWpOXvLAhkBZxj
3KP7cJqiR9g2WX3jgH6uQAwY2HDtEf0yyPXDKhKV8+VFB1EDVMzGjPrDJW1VJrv6
tuIBZ++eH5wi0iN3B4W2GFDPGslVFUNuQAQo34bUdPE0L5aiD00VdOs3OE+9DfuB
ebN0JQmL61J3IeeXeLEaiIaCPBq1PvfRfk8FvqMqGWUdEsjLDMZFOqI4dpvjy8Et
5T8rl7KOh4M1a2Dr48zPUAgTMusaZ07voEfgJtv+7v3Ub53gr//pxRoyQmQu6svP
pRFkBebg1MHXT1C4cE7dH7v8zp+HilVUT40GQnkc7yu4cHfVF/sLl8LXi/STWLln
XfR5+5YvTU9xMch2a1BljdCx5Bby04HHEkcpasU7itWNq0qH78M1DkvAlk69GpSM
Ro/1X60iteSr45SmBsx9/rpF3sA+TIGy6CDTrdb/vyRUp0Qc0USEnhtSMiBPGoz4
2+ik6++OHF8Q71O3J/+iI8UXGjKbx2CYQu97mcrdwwAgNSH/XQrPG+Ep49+OE6Ls
wTOaX4J4xxKre0GlnB0GCK715lOaFzM2E2W3tcIfqb+qTkpQnALqcuquLd1jH1Gf
5GSteFBWTquHm77o3Ya50LFogmzsrjPdcCnv0x/9I87pctwJRxCwWqFxHLTYKNTt
mnc20Kzw4PbnxWoNm4wIpQ+SHriG7axPGjKntMMCmrtH0W+rhyFYbER98cD9QHDj
GfWqyRsbwWEPXowWht1mUjNbdC0m5oAqKb2d+QWFeY7ETR1GA1VYsp0e0Ia8dw9h
huhMnBP9+DmOBK/x9OvL/RUfGrOapVqO699Vk2UT/bNq7QhSNMYgw4ukpToEVBZF
JVUupGn+SfysirW4EUT9DaAsMcOO+47PF4E63IDZ079LVHbgqB4ES9pbiO4nuBaB
Now1gOAEKrAEoaU5aCJbAXAgHlvVhDnzzJicGaVZ5MeNru3GJ0m5bC718jyk+bIR
Z0ssn0X9GMV2dayahk0AjUXHF3Rbtm987OaaNLap/nMPiJQ4CJ+Xg805ov22SS0q
urKhq3j1kEONmPrnBV6tVFGtsdszwSgTFn0jGrHDJYhdwADZj94VJsipm1o3p4xG
hFD/8myey6ZXFLUWUyCyY8a7II4jwgtxYKB2ynA61wBdbi7RjwHO/JQ2fVOhjBaP
ZxD/7pnoVRI4KMIYLKxJ4WpurDdBGPa/Nl1ryhUjuNFKOv9TeP660mdwEgZL7Hd8
sosxe+/gTscBlp5AmBa9r573PW3G5Qv8ZDpcxTLYjja9teqJJwBM9jRnatuTYdOq
eGSYjNi1yW5KAJt6/d2eitvhky3q4RCemexlj8/OAzd+hK45Sg4TfFQdL+6UJJNF
yoWk7gJMjV0xpF7u+41JyPip9qWZJ0Ib3wDnJzN3QBHHfTu3FbJCeYLeNXLokgV4
zlAd27xCXHgaCYVTU/sGXHtC/TkpdkvwoSG17T62wnyIhuGRjocCUy7X6V4FAu2G
Mj/9BUwiNcsEne0TG/w/5wyoBjZY4Bj74LrtNu9zZIZmTX3xCwZ1RIDTgzB/EeZn
gFDf4AjFsmG1aVGPjtMZ3bTWsWockqLUsYbKoZUlm6xQHpSmEAg/VMOWQK+ZSrwJ
BFDuiWTw3B4rTEbZTSkyaV2NWQ0v40pq7SqC+5gNG24LLmEfgT3pV7i6dFY5caog
PR/H7RIECj5q/Z0ejGOCQvefqxB7oPlpcC+cqPUkO26OmFtSe/GO1+FYqlx6y6Rq
8j6w6Sz3KVtXT+NUqkg8F+m17bpvC6NQ7OjK/Me/NgzLtzX4D4EjCG8uh57bMY50
5I5jguJ5UrHHv5PU2L0GBn6JY3OZc8KwmO8MnuPN6tjvPcCSf41s5QxZQrTlMK24
4oFKTNuqJ9mpqPCmJw6Y/MMqJ/+448hqmcYXwZrc2+cIs90uAdUf9y3DEfrno0KQ
Suxu2TLkkL//qo0k9xbL8vQwv4DRf63kZoJh6+C/2zUziP90Z9tysKUtb5H8xAJW
idWqip5acHu4l04s1/4WZcFH2LiLISEa2n+k7nlTFK00oqR+W3K8r6/Uk8K3sDl+
WUjZ244Renw9VYYKhH6pL61p4Z5GRF4EVcaOdubd91apMsR1bjVBsOchzYy1J049
9dzUu7WY3DwwaT9oZ4nh0Lli5fwiG0/m0IbhVaXu65B4zsZGDKf+1BPyqGW1bpqY
V3d9pTYOS7RloecTTDoF6Fix5Hzkn2mfk/9l50dILmMyaM1wnz0fJMI95Exu9EFc
pWQOggu2mfIiX1Qj0nPELRoft2MZqcK3PLvTLPXfE2n2Bjq71etJFqSBMlnXbMoB
QLdI89Yg8fZHEBq6mM7R5jW2aBAZ1N+iIPnJGjMt6C0263tSnPYpY8wE5FNlkE0w
ndtuPKneejioJaM0gMH8bqbYIXPw97hcMLsv3cUGF6Xop+frajLeY1IsY//urq/B
+5H6+JfYLCn3XBIAGotzOcI4LQkGrNeiiw71tMWiIfJDCBm/P6WgOObenX3B8nPZ
+BP/1bEMTqp2ZQWSTOUaghy6FSZfbMg731G66AM0O1zXsPrFLs8cNZqf2lnQnh0L
RNTUD9Jw4nFIIAU3+4EMtoi+XPYJYFHRw4yjcrkecrFNDv7QecVan+AlrKj10OQj
PbfhPttX/TjJ2EPnfG8Bbuova9N6Ubzjg3tbSRcLPjuAHTDRz4h4Vs2mEonIwMT/
vUmt6ogMc4dFiysUmht+CLL67sUTRKjq3QuhBCvAD/T47YmuwSX158abOp4wM0Up
FROp/4JJEI/WU+aXIZm9HeYKwt3SlSQfqixUxJ8xD1DswCrO8l/bUsyBbSooKuYQ
6yPE/tUj7X3RtW/2uY5I6bIHXzgBXT6k6xKlBEVMs9PX4Xnmnz6Kz7oUzfcgGcQJ
vloPkyI4bnnkDPkuFCSo1xO08wYP/qPntfvZQTc2EX44zH8I+lJThuKF+IbpduCY
lhT1IRYiIsgEBfpJQ2TkiPfG1I6s77lOUNOIm3rhIy6z8KQAe41oUqdJMNdSqksz
048tPu1j3yfjAyH+ugBdcV6Zpfu7kuvy9fP/xc1s5eVXDeuj/+gczUD5J4dMfq9f
5iEMsHgW87txcyz5NLMVTuNfLCKSzYLnwrogBVJ39pTpawJaa8tJkmB/V1Jo4zdA
NVoHu5F5J6awNfdOjcet4vaFOzQNRtGaGSP/b+EJsJM/IhkI9A5vzKyWKDLd/cym
1DlxUt09W4VrjA88XWyJ9LsLsA/iOEEA8K2v7l3O/9hQxbNcQx3GB8IZJtAm9oMX
cEsCE15VKEQehFtJyNlPi9AatHg1TPiXJU/Z0vGKO2UPcsLtGqWnQicbEIgdoUhk
x50yYh7eMKedgQzSKvt9Cl/4GXDPsHpar3KKUHEqIs/NyPd1OpsvluymB5sAEk2j
SfthpLhEcqhAdtjVJDZZxh8QBKvbv3NVe3/2qTc+pGTPlIurcs/z96ucBbMOS3E+
JsuNCUZ8qL7Ev/ucdzfGOF9M3rnDagnl5YDAn+eurhelN2Wga84UgQX835xWepCf
Qs7XvfUgA5y8JqkkuPDsnM/WxlBrKRmMzKi4dAwBgNZDV6/LZpUaWcsYRFcgQ4wu
Meg6FI/fQ3qDLy2aCVkjh0MtG8eqVzKPRMJQobFHAE6VH/RaRKWaXTMiMwX9fCPm
VlOXi6lcV1OfwYIT1ndqT4hpPduIZwUZIA2FKEeE0ibYUFfT3YDEomXh0F4GAv0X
gxMLUFUkGDwwrmvC5nS2tOoGYdzgELYFAVHG5J1AwSxq7zcBJTJwxzKuMIOspJW0
HD1/fK3jPRC9epRlUwEgi5WC78Yu8hZUJidCwzRL7a2WJI42/fwxnNoAzfuosFpj
z2O1Mhldd/hjcZhar5Ehzw7jd+KRDh4XozeZcgATl+PENcNorR/dCFP7ssikbeAB
LztKCv5/0bvHWQjsR78nli/M5gWqV9fxUqUFmoKU87VcqqNQW7m0uljMSj+39h31
gAgfrJAY3xRX6yJYS1Ek56cUokui2fRWAoa+PpIANvg4ECaZ7snX3wOLQQSbn8w3
ofccyUF8W5iXizp+PGsFyE+V7tm02KVScQH0MjL/D8icRn4VOwda0KyLn4kbb6Xl
Ui5PLRPK85F0neA/USgYJ7LWBsIu11Tpd+HXuCV485W10ynTe8mnEEUGUBwbnu+o
atLwoe121lLDOZ4DjDRPFb6wdAOuyG7TpMPZPpeQR41xAMoGBuL1Crm9Z7MHuwKK
qBDnsApDyjHALW2PwKyS1Lbg09LE38ON7YN2lPpIabMFytqGR9QxxlfvOhXMaKgS
nozvGJ5G13Doj+xuXl8YuXlijtJ/LUedtyi/kwSVzp2QltMNZH2xIt2QPpmBTE7O
U7Wp4sKgxoe7boXDbwEeaAr2NMplzfc/7gpuUa0ppJVaaV7Ol3MtM4pbFzaU/eXE
XqaOo0h4DdhaNqRFOGT2/5i7OIk6QMG/3eg7bIUzebzhx8xTEgJqDcFcE8cEK1pK
ZQNfzA4Be+2qTXUYBdGNA6u4E82Dq4gjAPdFS2z3KKI3px0nQGFzcJFPPtPW715q
MFcZ3WXCvrlu992NaWTQVBRBtoW/TbUkohgm8La/a3kjzQ8/3IvvScfER3WjTYHB
nXw89zMKOQkSTSM3hZJJz5WQhSziL3tleXhqMRDcdps3RrfkKmK5cTlO+/AQYy9s
RgVOkD8QPYlc++dEY+cAFzXdpRJqsQcNjpxTlG0mabOQ9/RFQSlfsPnAMg3yY9HU
3qgh9VigxpUanO0qVkzkTukbC36luDhoapBuq3ivMFFkSad3nnD+w5C85XUXCfbt
mAVWfYVRXNvscy7TmHbi4Ubof/4zNJz0DLABchg9FISLPm/KvF+WsaJghWJQ5xjP
jBFISlRFIB8GUOfxQHyCCkbjzPpIhXQiPIz7EKcnFu0ZtRhQ3Y7LCB0CEcWMyJUi
bKfI+OtUy4IzpZF9BJ6kivFKDFPs9MsUJQ20/u5duZEchBvx7mlLjIMvwsZLA3VB
xj7XSmO/xJ61kuR2Q0bdMY0UtdHEo9GTXAxsoaT04Tnj0Pk+I8jNsBgMNMseNpL9
AG4cN9kAD15ftEUUHo9zjbnBLqa+yAoUVuoievVvjuTOFk7BhZGx7lExoZf4yc2J
R5qVESNGy8YhaX5UhTa3j3BjIvEPIM9h1ONGDiK/qOoA6RZcq5Vnhryzpa8gNPoi
jE/8fwUHKWzgPxqY3Ofqt2oKJwx0hfwlnSWO6fm3LNnAjV3kRF3qaMUuXIHwdXaL
iPcuJzMQvxHX3t6XZD2SJ6IajP1u2p+qDVDKjE1rbUc/SEFSS/R8KdkfRRVPBI2g
c7Z8g+Vm5+YqZJrDEasp6Z5zgG6TvySurbbQ2NQ9HUkjyS9HTFWBbV7SWnk9EHZT
v5qnu10rxfmvbkf7aPRD5guFZfKyEB2jvosnfovBI4GqvWnnAl37XnL+aq8Pccs0
7Tz5/FmcOllnou4JbIXmRZ6GY1RUHkx+BJN3FL9biYjUhsYL6Ywxx3557bkYDbez
VmRPQxPYqfAItc4lRkL8bPgsDnaco1E9ALLkyTYJt5mjUuzY5jZUkhPTUkXy151i
mJurEh+tmTKpSwmsCiIf+yRBdpSxQ5fmA21KuN5PxJbHaJuxd/FbwSSb16l5o8nK
/4vfYgbvlUTCLkgNM40xACo6IM3iqrY3O8oEgIplfrY7A5LWQgGvt1+AXIMDB2VC
k92l/hDt8VG97uXI3CsIzaujbfM37NA6P2W81U2MtOvfLFnzyliVjjzeGmWTKH+k
ESPzzAQExEuf2kR0UOwVE76FJo6LaQxMjSCcUP8gdv1AWwFAzni86b5foKu6mK3z
jBxr2GRNv0V2+ieMW7lRQecKowzwELaAWx7n4H+h0acDDg3Lr7CpXWGmtmPLCBw1
k0gmUYCauYqd4kE370cWgdqW9NP4We6HILVfbdS9JWEbz6qb0N0Zx1tHQn0IXeQE
EoiHF40UJywPIN2UBZ0eWQr7lKrusfrDSetsPprUYU2zXZxhTTXs//fRCGYuWIF1
9luJQuGK4vWgYYhJn2iRPB8fuJSUYXQbIrNWYO6q8o5VRK6EO+Ufw/xxrDpf5ouM
WdaCOj9hpToTFYdT1rWkWcTThT3+DXlh2D6wlUxRqVJ6pstBpzOxJdl+0k3Firsz
nq9p5Ud6Q3rWeIaMknLNT3yjZX+M9QbO2slbD+JY5E+uHbBThowkW+TtnWeXLnFg
h3CFAg4Ad7QgkSAqU3Whj20rWCBczi5jpWLPQkRj9GJGxZUIAKT6rrF0qaOxiiFo
fg/WphcmYmV7k0dMmgBKbqN3tBgDsJR/hI26ROqA79bVjArTPc8CNoEBLgWpRejK
QcYU6vGzJ/ECfftYn5TOrNv3UwLN3BR6z2B1SSBkvApdLV5IomZ/7rA07/GazSXB
VwmEkCenjCpO0AUWlD74KoFNcDCxg2zvW5hQ6/DeQzVyFhQhcl6d4T3Iyr+rOMw+
YqJ1Xmnv8M1ug5XLUz+m6D6yb5i0a4Mvskxfjnoht2qRAFX7S3Ju0Kh0gOXplhYe
ISfdsD+hHm7fDj1RaBuV7MYpNFigpTiA9FbSPRF/eSCmOTL8fOw1aGfiaoyYxCzC
gV2RQedmSfH0IuDubgcbjroxZ4S6Hqram/Yrx+tUrA2q+W3+dcFHRQwqoIaTxoHU
7VuH5ojosIiiWegqXJWI1DB6XvV1QfSB/HBw1d44ix97e4UuG7KcWZnHZQ4i9BPL
1jVX+Xe02OnmSNt7nhYVLNVRhWPWav5AwaCbaBYAdJhi/CLtTwzo5P10lDYeh6mK
4gUsJEz52MUUSOPKiFKPyKjMYGdFJlglctUJ8225wmKJ4YzulyhqoX9x1/m/KnFC
rTXB3YxSwJ5PA3qCJwGwF+RZq5qUrDdmh+Wu56784w2ufnbwp5kqnuj2jBy0kilu
GFP9jTetm/YrvnxoTIzlvAYYcBdp4tvye8+WPRSPsz1ov9d/ULsChU/IPdLZ5KlI
UL+PSf9COkKRJuncPdJqZ9zcgFwbO12lUn3Bw39yzyn6A0GKMcMhKL787FQds8rE
IWRopL0oJUZt7HxLFhs0u961dEfMHg+JLCspOHytEjwyffyGgBbI50DrlWz9fAAf
naaBaDmhSG8mSTKWMyY+wE/Np0EKBj2l1b3GYpSvUri+OCk+HjCwjSR531NFHcWx
bAe7rIY1Jo1ga/DU+BQmjV6GQw4566/C9dUlLHuHciUY6AgLbTwa5joOTdyWpOhR
2zXpZuwW687KVMfqpJdNL2Rs9NSsiJ7+2UDjNjWJOLxRlmCrnWtu595TtUM8kNMc
yZZIhnd2cZKR2n6Xjd7ukHhn90Gk82LZ4WZuIqogv5J1vCsgBR5KyZe5RjloaTdb
r3015sQq5C7NrS3SbDEMKUae0QHy/A+oqelj04FdRaZcTUTakpVin/0K7ccKUdg2
PWFz07CrjQoKmocSf6gszdCAuPPtIT87WSMKRDk4PpSqclE/AcJn8LEPpunymhC2
dv+AObyFSBY7prGLY4gbCSHZkpVRePZr0cA3zwJBuzZdM2xF/6pMXv8vxatjrQhk
e05Zv6T+rtYGgaMG5eKmE0GaODpnuzAbwPuTZAT2Iaz9mKiAYkOHX3DWVnYkm0dE
tGz9EVBldtj4WZh+v54pQLH4UAjVIV61SYtomxIl8dfFevJctSNVdSMDjPuG0VYa
9+Xnjb29TJ82JKa+sbLKKOOWqgDeqqK3t5D6kYTr8kWiGGjGaT5FUNaJhIfx/mcf
LJT7wbJvXA0eOjQu8lcRTogF4MUJtZW2txwRKYtXl+K9V4nmfgzAk94TZwri1qqc
dkm5syc1maVb27f1G2nZdCZkFSNmRAhoLSmiFOLrbUWJDBvmBawKEkxehAFIQXYH
jLf5ljrbrFQ2lbE3priZl7pIAzCnMbNP1Hiz6d167NB8Rz1rtVRNlDQN78RYn0xj
b6AueJU+Q1dJjbqqR9CGotiMdPD003HXMEbqrq7buddSoYWn4VVfjq6fA77/EUIf
ydreEtkTfv+xCNa36/TcunUHmYPyua/SbMJRzCw1GR6yUb7uFc2k/+HEkv2hDD0W
+X3NVE3lRSkH78lZiv609xbBwNp6gVEnwe3Bfx+lSPmZV4Z3mOp26jtp9IhCwttj
yfdT4RJkqGCBs/ACFEwmQON8op6hWn4qvEfp2HZjDnXg93Z9GKz76iMrmAZb5ze7
hCNcqLdwOq0wyWwareytpbzk+cBSXqTnTMlo1gWFFiOy1mOglAN5N4MCnyqWmvgN
EWA9Wx47rTWCNQU9sM7PnKtbRKi933uOpEQ0cr0lSIFED/EK87r1w9hk9B60hqPd
rumGCMmYi2bqmftV7bSaAT5mSpU3Noa/ZVMgYac8DqM3FxYBsLEwBFZTXT5FL7Od
n+Vv5/EYU35iLYhs0D+FU61oUU0OA4ehRBvnmO8KnBuZlO8COnF+uhnN9edtBSkT
abr7BhvRgf4pGbWJO0fYlMQbs+5axJhKsf6O3rqoGxncXxmaiPSoLMZwAHOyVOge
EdyXGsUBg6J0yPV3kCWewUEvDLgp+cKymgw2+LNJucWtoTooEv2UcdO6CE7yShbz
tJUnS7CEWvMVKrHUgCkyoubqVns/4rNWQVjIeW6c8wAvgqbvfGowHP0xPYVYg86i
Pbhv+alDUAgKiDaANBD3sY1yenJagPtcU1xIbtxOOSISpLkFuEchns/XKsC0oiYx
aMbzVOj7+z4qmb+GHuRsKYLoBiNBVqznVKe0p2nLcKT7yKIq5JIYZfMfe6XX0iAG
Lt/lOkIZAiutDgeV7mrLqfix0SbwLp8HQjnSsxp99JUI+0nShLXbfSZ8hKLq7WtE
aNjw3/kEwWPn71mJjenZYoEUtUPNAG6XU1FsYZ+EHOUre7GQvcnbBH7OcDnok087
ZEBg9EBy7Vf/5vHk8vLmXwyRzFLJFNvkBZPJ6rUVHoIdTIAzcRuLvlj/CQIc+Fvy
kehAmE/WWc6M4L0WcuXOllk2vUqPQzgMAlDE3fTfnhQAHclOmODeifa0cejeTYdr
cZbR8+UYZomqCvm7s698lPLv+9tq0E0M6GX5LNFVVeeUr8AwSRA/0NMTCE4GO/uy
EtO7+cc3TSvc3YG+L8dKUv+ixrcDAiJk2vxvj4UbFmMkvhB47eE/z16f0C6zDHbN
5b/kG92pQZEQke2IKJaF/SLyI5E0PIjHXICH46Hn8v3ByaJbpxXV8ms9x0Vx8zL7
2h26UuzBM2wDwMqowoyt4Bk8VM2z+i/NqXzB2e3jFJwhrBrFPSjUlqQh3YUuKwtr
ehbfzFQA8Dcwh5hryU098f1Hdk6gvxvP7qWhEH9yt2Z4ELCvi7ID8/dehGdnno6p
rLiolemR26eRxIh+/HVNPeYtNZcqCbP7rRuQ9v7D2iVX5BEr/MeTX4WDruNhbBaw
ZvoOsZZ24xMuYYDXlMDNiKe644PIMDsYGslIrchG9HEuSXCvmM/CI1b1Ri2y0/3n
jAjWWEnqs1i3R17rOz8kQCILoDUuXIhdtJWiwJOZ10BHhWnkBwAPRv1y0u0j3s67
TEcmyZOJAZujXkasTIBBKnzX7IReClJe3UlhUjLbSrGW6/9+05q/D+PVoEGySMGt
eFPvR+fAUuN+Sry3RSt3zCUPr7hf4KwnYFl+MPpC6GrTpBYMDSBL4lTTGThTQ510
A616l8/l2YBjxmX2hKmr4Dvhvk9gMe2zq/+nqOBChpoGP9RsS/TRjl9PvIQsKwoj
5KKC3T7gTvZVV3r48eFfsJZ4RE3kO+mV2/K9X9Yh4pDXVSdTWwKfzJ9FJ42dsswf
HkqtIDYYHa7mbvZ7w8WeIF9QWgz89EohlxjuHtCAUJZTwYIPpW8BKOKnwi+460KB
SQWczNRSo7aRi+bMGwsQ6O84cu9sTvuqDgMF3hZIXZpI4/z/xcah6ZUQnoi1pnE2
u3oaGzJDcIlsOFlEE3Grh+2yKxPq00D8uVMDmMJvgsKN2UcCdWcs6eaHq+0UYEMe
BCmxSuzwIYefcBe6w+L1IcAU6uTMbjd6FJ4D/omSIKpt0JB6Zv7g8osSJoCmqDk4
6kAhlneHTUrBKzmUI174dpMIpE+FPW2MZVw5bGrBq+dFAVnzXgPuE6metQ5ZbbNt
qb1mVO0Lfr4sR8iX8dHLQb6+frQCgdj987IchEcoaYDWs4mCmKAAe9/ning5shqM
5xP6H9/ty9TpsL2xI0nADZ+QKQvDjvwf49yFsGIn5w/V7IvnGwey+T+E5VxbXqzU
eUKYzVMSjVu4+RYMQbg2a35hqAJouXrFlh5Zndqw5mBYxF+yKD91FD+LNd1L0uPi
tS2RS07JbLUZa1ntY+Oth9elXAvGZOctOctAyKFwSSBMZOOSWKdQKHXSFD7Yk1Oq
E6GagmEbDXGbml5S6c2kuaRMbX8+bkRJo6vVSumF9usGDY3M6NV0Tkf/7utLD3rB
kKY4FVc9JBTAYgwDMAZmqEwy1H1ByuppMcPq0BfJeTK1hPM7MDxV3uJJT5SuIqwl
lZvqndzHJHzBPrI0Rv9yPWYyzK7aXpFkKHwcjij9mJpciDA+R4ALnF7VsQCHekA2
RBHuY6iR0909Qen50p6RQmebYtxPzlEB34GxF87fd08Liw+q/QSM8sEL4HPPgSP9
1LEr6gmX+TswP8ImvzrGgLqmT9tt3Gf1GpI5JiP6MgzUsWNWHxxB9H6OdQ9+S5RM
KvzcjD+rbotjamtrAW/vOh0Oh5QovomOv4LZOqSzVSQMkSaaSpBFvZXg6Yxw3z1C
LuhWTtKgRT0GPibBR0X2LsNfE1zCQF7Q3V3JxIo4AkEr/OjdJYvtLhpEQUpDVBXD
thvhmrJlRcKSt6jyrHPSZUhy9XftFMbLFeLjGsvnrxyp20qAfzofaTT3Lmm75POk
qe6umj+oJ6k6h1O6T0InI2PPVpdfas9rzfxf3md8yz+Zd3BKM8OF+74AXCPnPTOs
jQzcLqFfIxRuNEKiL7ht5TxDIzm2GIwJqRRzaBaiUyGARZ9ZS3VtjlXdrYT6yll/
V/7kVCD/dhq8n7d/w0HGcO8vXQv1fFZ5XqgqdLxxrMSY/0bqLSies2GHptMFx0jz
XUY/ER1kJV/z0bquakMc6RXpvawaN6bfWfC8sMV9VcmBgqC+e+Dt6VBLOztmzqPp
2Mb5iyRWhIhDqsyKX2bwkfDgEeX/lMu7ckoPWJEkcy0BYtYVwNuQEyOZWtD6OHCu
PdhvJZ58dnfDIy25pdRORQwz0wpZE4ddAPg7dSzeq5+OGvzfKtlDduT6M72qzkem
hW6N60YuvP4seRxXzfFajYxIXmzDMKgOgdg+dJ8RALi7l99ftTnRmxmmPIWUi673
oJ5MNNIc23mlz2/rrSWAA55otQJvc77hzLup5es71hd32VtWPmDXu46L7WVOk2+Q
PMnOPqcccxMbLe3JktNzxpG5kbqVPG1u4dJFesWGfTeXNkIahmN3mmV4mqRlHmkP
KX/OYYM1ggpDPktdW221w8pnyPHYIb72mFNKD6rucZdCgzlhYmNjBHZtm5dZiWsb
uOC+U6u/3knY2NHqGJCgRplkgWzaQglr6BlhpTIGjv/KducJ1NMOIV9T84jAsZU3
XzaUoImPmqTKyd5/ZwwfZsWj7GEERKou+mM+3zkm/JmvFOSmdTsXQES5ws271/gW
xIBNFyNvjVMKC2BpBSksbIXOPdCiuZBj5T8SmQAfYWuyhJgalgR8InSSGVSKel5X
skZU9wH96PBxaf+mZfme3FgjY+6ZCb4KTtI4ZKVyI8T7smQnvvTPFa9j3mZvv10t
/FNnPLjaiaCff6XEa4k6HhNTH0vyRyEMQHvMsjW37BdPfz+odktyF4QESqyKMfwx
W1+06oRKxWVX5oyTwZEGi2XMno4/h4ho2IPDcvdg756yK9Bw8o7XeOMDLmr/a6RI
NFKg6ywy3TpTKLxn9kEL9B8rerF3clrZ7Ndeyt/H/S7hfeqQmi5eFnxG/uiGQql+
9ZvzQCELffbRA7mEaFkQtUX/G/5rLpaLR5BTS347bA060AA5lgKX6cvRkt9LKzsr
lznAJE08on9FYKrWXbe27YP196dkpEfyY0WlEjMUtW8HHi1S1L4KtLbkuE3QWYtT
4HfPzb+6uEO+X776FevyGKncJEgx2P0F0KyHpNhzJJi4FQWUtfLAmTTkVNuKBwwN
vlSghdxzqzYYs/ufaFpFLIKjcexplcMQSwQYcQ68Hn2wbi9Lpqc8fxJHXuX+ynRF
qnnnetPAUd3U1heB0OE7aQ==
`protect END_PROTECTED
