`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idB461FtzYm3cLavid/l70TuMf7Fe8EPBKTWuxjljA0SWBA+O6FfiTO6E30IrOP7
WYNVjL1kp/GtlyfTeScZWfwvwrkf3Nqs0IluO/5uERK7FFHtaEI2XCOdDEQmMBu0
3Z1xrhg6eYJ8qmjauE0RmYdxjIPJns9o4Itf01cFrqxIwhRq1JOIKBRdW8tn8F+K
qED+O2n+aoCpaUV67QZ7rEsNabt9pp3ABDDouk/kdVKFhM+5x4Dw+6rqskn1dqvs
s4FYex4p+dlInTQ8/Q4D6ujycZZvkqBzpV10JPD+qBz7agyooMrKmYhEqjqqwjW6
2wSjIyjZwAVqH1OFyaqAmQvUutqYxo0rMtmMYo0uHV/6SwaO6PTFaJlVxmfBefLQ
IYtR4E4MJ/hT3QRYZNkn5OUhSV1zS/vRnlERMpciVj/ZBQABVs/9etfo3aF6DIkB
OLqfFNb6aZVqu0U6gq7YIRhIJhkYXCOVfBqYAEs96R8t/EjiHCLNg/3ZNjiMHUjy
yRCbB50N/xEPUc05sDwh9d1WhEfvGeB6GRSTsFDwQZcPLuZveHUcSGapiWYF1/dj
G21HuBAYelCS9CYUEngemP6cSezfhoL9CzyTv9ClGJ9/VrhljXbPSCQ95z6YN/Pr
77UkI3TDtXNO0Yet0Zu1YMuk2L+G6cMhNlhGw2Ci3IJ0EFIO1oLvR3KhrLXD9oc0
jP0Nb0v5GXvB6RFuLTEJZZRPQIwggpSYRBH3ei5iUJYCMoXE7LEbnooyJJ9TAkNZ
naiooVT05c+6yRzk6lzds6let5A2nk0voA2/Ijvc35I9o7xJ6p0gzw2fgilIERrL
E09Yt9nlWAahmM5nWtDCI9pxElIWcxO6k0APiloCLFUzMo+bLOSTy5WvBR1+1aow
CaTNJpqG3Jn73AxWei2iqaI2YfaaHqHGwroFXwEa0YrDjIZJEU+Z4h3xXwj4v5ba
0DJsRsxol+spwUzFr0UFSKHjyw3zi4qd+MemkmaOpukeYjou23n6xFujB9KAF2xm
ODP36CfskLMprLNXKIYlpFEOFkv/HjuudPTOAIdMCglAaq8AFBzmK8rekXEY1usA
MVCwHcVBbkMXUjsDo/u9LU3zZAmjmwbczLFWiHhWxVq4/JHoMw6a7Wat3OEYxOZX
mnjbcZm9Y40rkVaohHjRRfoZzQcIF3LAsZBprrr7aqxQaAEtd4SSXB7bBa6J/nak
aaavtr5uTysI02s2IDdRyySM7OtJt1CTGTH/UzLytk8yjxN1zd/4OvNxhLJlzJ5h
MlAsRliB5EPBDzv1IEbo603WYWmB5T4p4fFLVuSa5yC2e5m9omrQrZH/l2CgABR1
VG1FRnOGl16JVSLk1xHOJDmo3TFIz4H24ZLiGxu4Ws28upWIv/nHiymjZvc3WfLm
NGbZVZ/0/9x90gbaMcWzoxMVjmh7DtdO4YNj0G9DaBVJ746eCldec0jSysP+L8jW
SYNGs4QkdBvsz+xaafMKFI++6t/Av/0LX7oLkWLTo/Pb1slIMzA18+4WNehjk/Lv
igpVIDJyNiybJQz+qvsYPYu97DLdDXmtMZQ9tY6D2WLAet6mICg8jjSJtEDi5N9D
gF6OxbCs2qxioybw+F+Tt8PiDzaKE/b84WG8PM0qxQsD4oyjnNq5HiGWxdzPBJEx
s7f76vp20ww8MZ5WCO5UyobH6GA4VJ3oPcMG0BeT5xLmwAwfeEYLnHUWLSoKdaBW
zDL+T/OPXRpY9q0crWxPq4kKs+hiTjnydrDE83bGoHyhORf/4Wk+v3alUlwLszZ2
XG5Hs+qSCDgBvnMw6O53s74RfwM2eNv9tSAFpejo1DHQuE+TedPcIbU7Twk2x1Da
SaHPDec4JrOkt8SBESllFDcexty9YFxBlybWk4wsFoOTxwDYkpYidoBqEL0j4OO2
SLbApvxHCje4W94FgicujqSVhXBuSDjpNb7cyJ0QDf/Y8S0QKT3bPKAqPhwWpA1/
6Syx/G9+IFucuVIktFC/L8BK9yFvYu9YXCoKiCPeo7IzYoXaFmPwPjEoWbBM2syN
t74RYy/DqM5HXrylvh1qnD+zKTfcU0mlM8S/NZWdN1wRfGWb7f/YGFj+mp2fKMJG
JcfMBEyjfDU5CzfFDw0F8U/Tp2BgF0rYpjqwvaGauvyXMHePu8yf3/z7gzezdKoS
1mLLU0rUj+FE2yRHMZoZ0UmOphSa+ZFEJ4QX/byo8RnSTnB/pk+EGpgZL4LCtpeV
jKuoLn6GXO+9gatHCl82dxiW+KXgFnfGBe6MESDpwZJpiBQYvg2x4Z0R7VTT5AwC
7AQgxoHBswH4bTpE8oXoIQ8VDo7HUq0kV7anNu9W03dcv+7fT2HmlnTgoVbVTcDX
WavkpE8XAdyhsYE1IO0swZIXtAMtQjJhP4+VkoSmQbUFbnyRvPMmUBI50hhK+Joc
vvVD4CWA0Dg33NJp1d0msDuB/sLH1qXUEd4UbJXjVNCLrWL6u/Uv8RxO1dEZIu1p
AdkiPYxpUBm45PExsl7dO4mLK+SReqIkPRMMRwaDOTaSDHbxRuji8XH6yA9EGpHt
emqF7FJx2PBb1IRzMk0Ellh4uLNVHz2gAsrrBmFNji2n2N9Isn4LpREopwgZIN9r
2Z+dPijA/RldLlEA04J+lkL1OMKFx7Py3toGweFsN+MlF6XgOgrAS0Z2nAKJ4TwW
0S3+5aD4AnxT7UwZLD9JMkRTxZ9UDmWF5cUflGI3sWDd32bpyqcR1LnsR2AeKn47
pl/K/2e2vHlSptrq0hhEVrVD92hff6QzRZ/peptxcHuRk+KfhyDb9Vp+e4L4oM2s
V4pazw5bjbrCLHkOj1Fmhg81q8ap+weroiBGqUv6D9qbLWSGFemN98e/9epXl7hr
bXZA2FZHKSsaYSb/vl2WMZZ3C5uewS3BSMVQ/VlDLIlT/oApMnGgFbin4dY0unYg
B4tSUdS1BVzBcYW3ED1Rlu09Xd+vUWdbMvNIiBLU3sWEVFHCXfwpwDmSR6DkOpo8
+f5m20tPlx7VzhObDew5ci3AZ6eRfa9i6B8GHeoX7asJiDw1HhtIeDJCwfmOLxOb
zWAhM3dpFjSpX4LhuRnGlEbCwb7TBWoQ0rw1KW9lBOWaNF9t6ngCZD9zc1T6yQuo
UQ32rTXjusYc++9+jpwgEpx4UqIhHTnOTr4L6QErSyloI5FwuxEpPY4JJT4HjzdP
OX/0lROI8cnHUILrh3W5v5OvuXcR98wJHsddUIeFlxZ+RFfMcIzlldA/tRpaofOT
FdAsrDlPJIk6VXdbp8q1A222t9A9OP8UUCmFzN5Uz8qqhkz/WghYX412ENttkz9v
+LOclTkBOmKbG9JobodYufgGdh3gsOqPHqmR5sX84ghp5nBaymK4SVIh08X+qzp+
U0/1vB3+0OWxfk6h8fsj+0oCI117Ku6SuEicschRD3bfFh+4LrcPhMzYAMXf1Jmh
C6lX9bdGvIdZiE7eAyj+1vt2NUAJ264T+s/0XK7SIj8YR5oXYSNBckb9ATSJzffr
iLX4spMWKnZUXqwff4y9bdSyjIyez72Pgg79Uz7T3ea2D7Ved3XV5iwNRH0ZIOhX
MOXP/0LeKrDy53HhahfaXnoo9PDSRqV6vKNgSb4Q2PZ8+2IENd6XrtNIPQNGgAX7
fZh244oE5qlhm8jGNtfB19GjN3yaJqzhDsAye0TZE6q6Ehw/s1rSiOxddf2PkNxu
jUTn6WsMdU5zY/akjjl2vonPD/3QPKEolDvd6yCkXeixCwKAfPG5bTBuUytuq2SL
wfjVRrxYpMbGlDB966i+A/g8kFkPz2H8wu18qRwx36LfWR+FW2kx9aHNY4idyQax
idflErNgX7MACc99LPZoDhYZrwhwd5ch/tDoYA6g+g3ILEANkaXs7uKxIdCfb6xQ
6BtRwd+7WrXIunxyZZ6a77z4PS29vCUUe0+e8vpaFr+aEwvnUgoky+6QxDeTrpzN
g2SiX9I0xYJEQ5xjXxrCrPlT4vrcRKykg9omFOJoqiwOzHo5+xUEzeGRSay59af6
nfj8x43jRLMxlOQy/z7JP0g5o4FqkSVfk/ygkL5yJxs2E6ipWcOi5AqxBVT8bUda
NPvnB0b6uQDhE7nWIiTa4fg150LSsQXkAmmiCafQQldi2SH0zhy2VelOmC7DRLuS
8n5MZOH/Kxp9km/EY7Y95PUPNbHERx8+UdZsEsrZkg6l/bFL3d/z7uJymbJpBOxg
zT7iVKJmOBMKHuAfnHDJjAM0qyieXJxKvPW4jrSGVbWgNftZ7Zq1dDTQ3ew8sjHm
5ryPTTYNq3NVCDfqLC7NFUnWXDlBXATO+XWoEQ0dd1nRSIU8jvS1IlCLv5+0llAC
dWK4FF/P48I30BL4qdwKhZ84bOWrcB66tAf/+E1EwOzZGTTEB0O+GbA6gvfebNB/
/CTQIObPZEwo5eTDBC/7vvbVxRORWfpheVUgdxB2m5g2gdVNlakObES5ryzrp5Z1
4IV/EQhPmkS2IjHyCIN80cGtC6OJS4vQzIoV0U+w3EOWccFsm/5bKEYq3aYFkOSS
PKXsQIYItWQ7zYU0iR6mJUO0Xa/3ASjWjulpY4DFZajACnYibB9oMQHgv12nBk1o
t3AuzcazlJ5a5wkTuGTTq8BafuCfZshOMukAsQslX5T90QvnehoRi9/aF6HDEAcr
qdOwYYyfUl5ikYTUFHmqZgz7bDS0PS+RZ3pG6bS6L8dDp9hO+fdq/5dh6wcLSdTs
/7wxJ5I8HjDEAsDVlTDu9NCoem5OdmAl2tRXY8VdteNfNN8OFGy8ypkcprIjbY6v
2kdPiQaZ8ndH0s0ndU/Qyiupb0OhHCNi7tIKCcZiuaWfYxTvoW7ODRnyRibxF+dp
L5F0hxQv1+NsuSpxA530OESdMzxJnOTiFwxBn26zWn20scfiKCVZ2F6jQS2zCRWY
WFQaKCu4lvR7gINDGIK4KxHC5juNjaEuLqFbQGHRZeLBGG7d6dAW1QABKp+YlhAC
DvPeu0BetriKjhUBbWgHOFnMko1Qdt1RMAE9Zf/RAtPG5W8Vo/FY+tBLzW7Ihwa/
XUaZOqVtSdum7HvqEXTomByBm8md454NvNGRpZF9nvWRyws6gjXAjWzDFGxXbgvD
4rvISetW7k7KcgKVBUaTw8PQJFeAwZESvV/t6CA4QPRbuFYuhzdCvW35Js9RcKWB
/24hyZQrDLtmE6vrhTQGo22OjKeXWsvtKF0fya3F66jL6OwC6J4x5ujfZW8H8lFX
s8ibGQHErh2nabPw5req4quAt6B7/HZGs59tlU8bZ7uwNYh5jw1mqHCGm6tMGjrg
/j06xSrCy+lO+iWOMzkHQI3ecjCdkbgoptpsXHoBlbdyWdhXbNW0y2+jrjJMPAp6
jIWBTovjAf8cJEIrxxA4Dlz3GxoGpKWBhY1+7LFwpEkajVtYCZLhb0EtxStF6hPJ
o/wOouMTJYRAYAI1nYiZnwh8PNqYt6cU+FFrHlx+w6xktFdJqpKiIYI4JS6QNolk
2bBM5Gf4K+BhD1TiWCYNqhXgIugRyaY7mzG+RiQ94cdUXt6IIxERHC9RCSZ84U7O
G3ntNu2UaSQ2pWyMSRLq8YwD+OkHYxD5E9gVsR6TklvkSzHFCUU0lQ62TzdU594e
xTb5Ew+PH1g6LjpSB5pnaPYMVvZ8dXFk2HrTkxb6qu5DYorgvD/4XvplRSk3927b
O6Awbu6a09evznUI2qdgZM6ALlyhMprtvUX9l4q49ZJC4ASP1kUsSsqxZK0CD5vO
g4H2GLEtIc23W6BP6mCGeDllUkxdS+m4KaWUPBxZCSr/kPd55CWTKRDg2UZmWa7s
6ahTSsz9EubzDd/NRwhioYo5TDzFjJe8xl0LZrhcGmSSlW/98r55ovut7KesGnPF
9Jz5m52ISx4R3i59xOa2nnljNuoovSuv2Ar4xBjDZPzru2YTfxnTLlPvVjivolbK
O8r0JS8e4gi0HdBQtyarnSX0YAi/06uICn8aPplgCG4XSMGUBvSE4WEOOb2tJ3KY
7IzQvoZ022dyst3fKReHjV6yHwRmWeAVpuKdawjVSFB9NZJqQmK61ma7CJ37yjBt
OyJnLZ0Ufcl7V0fqtTHEGqNpVxuCn+CTwrBDP5QjYD7Lbd1Kjk+bjZACySZEQ/Q3
/U0iYAn96U3XaQ94Hi3JYxXIarjFAnnUX3s1msO8jyH9apE5a2kchT4ul7CRPc9/
zUlukfrk8cYoe8ePQBy0zPdcCZrcUmZ6wpDCORsh9s5i+7IY28WNnc1855yrzZWP
5DtmrxmAKIzc04OrO3KK1Aof4xA4VTZn7qqMkKk7GzhND4DAmjl0x14FD5OCoHMo
9u1i46w/Ep+MkWQgXycmP8kfLwUUAZ7kpkGSoRKsfRO/6VhUv77QrmxIiZRsYo9A
W/2FTTdGWkUUXltdfAiqtnrpMJi7P0XRL+LsvYqgrZVi5HGYCKWd1cJkpg5YWWS6
izXGk1N43Q5YhAreUMHxSHVARPmmIxlf0isR224OHnYXSu4bQ2rhBlIg/tQ+eqeD
ZsiLjTDd9SYOVTSDzXTPf8rXzIDw6Pg5I294XEX7kpE6mg4kI9f8HJsctjLQLywG
mCRp8B7ZhdRJffY6wzVjn+N75FwD3VKxLtIqcRwF7r1hl2I8u0EsTgtAK7JgOqF7
zCXL+N5W7BX6wjSpoW3i08udWCivcOOZPFRjjva+SGUNZBQFophRRweFZ0gRcpiJ
G4aS/aOboCcTMvu5ylrZyNvDrDcYty5Vrh3SJXeoSSd7fgLNzhSaCaX8pDF/S/Xj
bESCQlntAebImCQ6n/lktGnSKY6WSVQ5v1XOlP6V9vxb/hTVfH4gRmOhBcrZhhLM
Z7KeSH3GyKPNPG6zbG2LiCrEkYKNLddXNvCjLW+x4xeEsE6W485mkgTzaDEl5/gA
uPfm/dDV5IQOKXeXNHnCIEKlueLI/4fh/M4P9gaWA10O8ORfkjP23d+xBUYZPp2v
/kqQ+5/2cYfMsMd7aQ0700dv6I95etDZc4mstuvs8Rx58iXrz/RFuv5H6mAqBsH0
muaZ6YNRHpFuUk8Jriw4tlW3BhT+iSEiES/KOGLKi2nKSCdb5QVFRV54aX9s3AEf
1fZzMsKV0mskbJM/9mMFcNiWHgPCAmilh5qeaH6dQx2TcsLSPwFmDx3I5wiu9g/+
3QIvWE+JcFNNTULgCi8iGuAawiVvh+ApoAw1Ojw6VMG7pYoDU26k2SdLphk1rOHi
+KgEORXVJLLXHqWOPR9IWOUu93n6J3zcS3H5ebpMk5jDhiF06DW3xPLIlbIZXRgL
et4QTnN01AxFV01dbvGHGMBwzUp2mxWbBz6TqRIWGG7Kr0m99c8LoqHfQHvlh/ZT
hLEDU1f/dB4OFaaCFW0rENQYtd9OEhFeaPafuUvUG4fOTbq2a10qt4mV73IMJXQF
fFtAtM/z+VaC51C6j/Q6i7IrjijTvOjiNwgToaXmaI/envXujWRquNZaSq9hWEvy
KhXU6Ad0J0CG6eNY10WgFgGb62tytjHrW2GABJj7L1qiUm2Z8Dj2a0QsGpWkNXtL
t7fHwD2ikeU4LIvP3CYjH4v5kGSElmD5h0G9DLTvNzIRdVikLnCzc2hnd5GYjBej
YXAH8/p3nCdNezQ9dAsGM/DSO2Zn+bVasNlFjF2mGoIryBNo79KO4s9S2JGHPsYW
wntuYV4sW8zerEOowj0Y3PYQcANUMmwzeEW8MVx2DYoh20Z909rGi/vNovRPB71t
m7PIzffgqiVpC1XdiQuSIMEYtKZlyTgfOY3nFd/V6yVZVK6EIe5Ej6rSiIwQPWi/
fIMTauUG3WTAN89H+/MAfUgcROgYYV1yZLpl15toGp96Ks8HYgTbmE6TxinNfupI
k3jeHQENcQkA9KmNwAn5ZPfS37MZ+8nLv1QGee9+yLus5xuBiz1qRv2WcZ9fyaT+
9GAYC6rO7LhZI1sTwfbyASmle+uf8R+dnb1FQdppMiE5o2jlrNxuZKxvIw8fMrBq
98HdBRgCt6nnr3wqMp71yoO2p7zyZjnPz9kDOOdCwfk=
`protect END_PROTECTED
