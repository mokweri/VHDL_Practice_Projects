`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AIoErgFj1slqNwIj7qJDm/EuYmMYUbrxHjLfHybS/mxZLo1DVlYQOadabuggn8Zw
SmGitFFhQvNncf7ADaMqXUfMJscCmRVAr5LAdXZ5Dd6sdfz9tWWjdg6Fbr/sPwhD
k/4pqXD4+q9uvNbvTO9z3KJsicjYgmt1Z61ytnALTNszX43tl2OeofxugoSGLTd0
/CZ+541Uj1CjX3T5FfqM4EGhyHoJiibk84Ci1iRkRiYlM7JaI8hEiwzjHc30USg0
il9i5ggthYxnIU6z7OJkzgoJgWjKVPrt39Ri1pKuLBkvambd+OtRBlVNVjuNMPlI
ujWoy76GqoKOxAefW9ioGZVC/W5heESP2xUuOr/bCHERc/Ka2hu++oHFi861h4iT
WIamD5vDXME6zvxN7Q8b2Ew/t8mzswxwaohmHTeK/fFf5HQgtmC7lHx/HgnzWWFT
iJBcqxWV7UU1o12vSiX0JIxdSwCeSFfDGsVP0X0jPSWdyBxvqqBEcQcU0bpnKc1T
Gt7pjvqyBEl3XGoNIXIZ+KV20+SUiQ+h5NZhI4lOhMxu/mdPzb6U/c4puXk2R5LT
0FKvI3A3AGftUOZ/kPV57vk6qd/bX93PlAhnd/IZZiuyfsV5OGivKUEU899ZZP0p
4chBPbYrH73klC50nYDS7P5y92sNG+cbjT2tiviz75S3OyI2++u8XC3t9x7nPVXM
0b/fA7qxSaVZU7EpEQ07WVlkWXl6fIkLrVUJ67h21fPLZpm9Svp6Clw0L6ADAJlw
Ju0HI8Fe24CYrfzRek6wA1ZoP85JSEbA+5jGrJQXfgZILrG+md+HsAB2OmxRO+1I
4UDV6x5l9rLYezn+7cqII0pZUTY+aUVV+bHx7T2Qo3M6IoK6xMGE8BnqfQ9uNGgk
CwAiIleOwxALuMjVa3Myjor0SyQ9vjMJR8hyQ5Q0FXE=
`protect END_PROTECTED
