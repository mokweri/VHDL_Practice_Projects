`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z2XexfBjcTIroWbdLYCRXujbXTo48Qcn50c/dbxxLFkfaQF/29jwOnLm0/bkY/oA
vWNSWJ+O46SRZ5UzYJaPiEhXOAa2edxci9uPvzFT1OVaupghcK3TdvsxUGJvbLY7
0LqUNZfCMdBxuW27PyDf+EY+Z5U5Nc7ZT8W9HZJe9itc75ga7H8EzWydFj2aHwp7
mImx3wo+LQt38mEj+peZcNqwtzbJQAvHsWl9vylx/Z/lJFZmTLVDU7JU6b3pRSCA
K+9WAnN+dyTebraVMIczh4QoB68rwUZD22nvMbCYBIn1SFLk5gUu2/PQ/jDcPNbw
QqTALvemRYe1nZe+JwwoaTvbZl2yY647Vdo9cCoLENgz390RILUJCTU5Iw5UR0j0
/rx48pHmmtwSgiKfI7trLS4izeHZ42a/BGlPAP9YF0UjwQ343SVu/dHvRzgZxeuZ
twAB59TAQ7rdODVRudO2HOBW/DgBK1eHKSmplVapHk1d5pX7td+LDToBZ4QBqLh+
b3+gR6N7NGOnK0Df33FcOr7t/BE/zeRPriO0BM5QFdmjXdmZ7hKNs72jV53Co6rj
k3ySDFugNOjJbgT8HFGIh4Fp97PtCYPo77vMDio5jzT4NJnEkwcTv4+QTjK/FUq1
Xy1jE2AhEZXiUcoQc90xzVTUywj+wOnQXrmLE6GO+ujZYisp32iczasmdP5CUzGM
eMlNHnKVTQ3ytLEto81ywwUHzJOiSyfh/0T8+26ItfCgyyGYbyDoWN/J0NTArwOB
nMckDvzLFgdDdraAqbDdMfURJnvvd4JYN0q+6xpE+ATa2SAdRnTFx+COUjpUgSRC
n1KYbBOyELkQhU7apE93Xt8Acne831oUrtQ9xUgbpkS0jn/K46BlZA3XMxSYtW3v
l6mwBsH0W8HQO4Z1/bHoTktbtfyd/RXVF6glBWa/uSwy5JXdYx3Va0Z167z9FUIA
r/3X9TkfyYmbNbGzj1tKVq+qzFjANlL1NlvoXNMNeSJc2q+magQOwUXtVzT2bmkb
2X7pkESI2erSd9IBfFG81c/Ao1rdZO5WDZnEABHeB8KtbWLNDDOTQHfwjeKFb7Yf
tUkx6LBGXTTfVfcvMB3MYUWAfuliCOPc+/Zl97sY0B1l5ivWceusNOBSaICGXYY4
9o/kDOsnZ6jECDPQODJndEcd0qSDC96QZEZmRzQp9/MlY+24ORcSxZjP1C84vbE6
5Wnhq2fE0TJJnjIEw2XqTaheNw5T9SvIroyGi294ErBrvTd2Oo/vDWFVJ/VlciBD
dsCl+itaSbmLmTxlOHMSrWOeLwSp6z5Vj/vEbf7tUtDXHhqFZBMq59D3vub5/HKJ
AksjpXpFMZZu0v9KDznMYHrxx5yBgrez4YrDHtWL1gbzWC9BkKclPIE+AxSZjR6d
Mut/v196L4J7VWpRNMVQFi3cKWDwNndvTXvf+5HIlqGkxqzdKe1+lludkuT0x1UR
2Bguizdv1zYNrZH9gwFAVf8BQhD6bvOrX0ndfQVhk6B6m3yBetnI91ohYh0H9PxQ
E07q0lF5SCX1iVWEK53OEOAO09xzPJEs5OdkHSCE6/ir+6j6IKLfVN2QOgR6a62S
dcgCosusObYNlV4BtZ/0nREZFIra53OaKHox6bBe0v09luIA/+0dTBJx/B6XW3nS
ufwJay+Gzs4YzxeFUsDhm1i3eg7bLHjhnCgMfpQSXMb266Oi/skOV17Ok2lvyr2A
un0uIRkRv1aul6jBw0h/5X/cIF+znTR/0h9vs9A5uizCIbmc/8cbz6muH6kn68Ck
fHb18GSfDYm0JK1ny9rmDB1EcPtUSV4R5YJYS3j29bE+CRF39P603nfhi7xKTZI6
sgrtdKVJrphM5ZN4Fh232JLMzbbsIaFuNOPqxurdS0HthA+ORtdwcrl8a8f7DIfF
p3E+FvD6oQG7RiBB6OvjmtNxSk/OOpDfFpz3hUCPFR4oRmOkj5IdRAxaaKl6LET9
DqTOZ1OdckcSrRtoQyYEfn9aikPxUY/Oi9mIve8UYH53JinzMeLJtLPjoTswy1aL
2cT/a8gYQOxhayn9H83dfSkU3BZe/VQ0uvMCDwbrwbA86FOJDGwES5QqLQdQodMg
tK8RYjq/dkoNK1TwexxWzersMokxjKWRva6c4CPR+ne1PBJj8fejTPMiVb52VAsU
z7ARuoZPh7n0XRO0MxeU/1VmEmto5xD1t9DmPh1fj2a9woIeQMMiqq5cxdtCNdsk
qKF5UgjVQt2j05visHKK67/4rKPsI0XMsyX3l7CvLStf5Q4GZmfo1Hm3L4kx4DtT
abWE5WsydKImlwNlwbYwjrcqGlUXFOj09WtcP3AvBQCn+SSzwwF03CAlwoXHOXZV
c+H8IN09tF4GnSgrlblO+cRQOU4natxJf4GYr/YNR7BEwDRWKLWJ3za3XwOsQCc7
VN37XOHoWz+b/iIohUm3xyRU8K5vPHcvytbvKlaDp9IzLUrAeFfUBUkmryCD19AM
c74E4cB3GPXNDHxfFqxAaO+/gFLz4oIoOgRffDWJTqKFKyolv0Lkm5pamuZv5R/x
lzYsfp/gT9XxPR2PQWXO1z91L6PreAIaO+svL6AapGfZ3zxLO+pYp2IVyoDxBmsM
S3V9aolO5g6ps3MqHaq9qfK2T8UB6xeOE1YMHiTnFGKFHT89QdNGixu98L4P6nlW
aavpUADdVhZ+Ba1whXUEBQ9L+bvtbeKo5ZieL0dnPX0ZlDysXzn6rh8z10aF7SwC
pWFLBAMPtqKL7er+s5K9o8JzYnyNduL3okzdgqq7GbdzBydzB42W3glmYS34qaMH
BWGi/nYPKaJngWigvS87ngHs30CW3oJaph3/+izG6MA8uJv/Q4BQf1tjTGOQuMaA
Sk8MdtfQONeKkFhpf6id6NNyEEpVQAZeud0fKotQ1+yT4uWVDmLlJSZIQKBFhYc0
ew/0Rg6g1Zai/ImnoZAuuNyjJeL1bL4jCBEDuxVP1hJ6WwV02CTDbZ2iAYmjsVtx
CaSEhBoWRqQLUdghGSIV5ZKXhm5TAqXJYFjWTU0ZAlcucD4PN1nEYu7b7vrwByoi
rl0cebjAAhf1FIqH52P9PIgmRwsuUJJzdrzzYDZ0h9e7Ay3xmQEiGJglhA6gNDGK
PS0igKtdB+T9BULU35+fhB351hAXojAVXB4fVxe5009aFcsXnmnlEnoap5K3nDqb
AaNvNOBz9+DqAX+2LGaEbgjEGqurM3cmLiv0S9Heo6LjSDBIcU1rQrE7NIAe6CjQ
jT2odRtpnPhovX1vDu4E92j+koEXch9jo+xmAqv2e77kmcxYWMPySprHznNAD38d
XPSqm1wVvyewfcgSjNlwU6f96SnrpGd9WKy/TF7jfLXpQWTubccejuiwFkbp5vsu
t/7o/FlgAkW3SLOnjLLwnIe3vCklcK3ZohoWdyHNdB/nHn53alGq4NDDAxCPxT02
mcTp3001hte3IW1261nH/lfyipRhCKWfyqKm1WxetWSmqh15VgIaTdYdgCTtpxZN
XVmr/bl0jNEzDGqOlyGd8dGBYdG4PsAVO+Trosu8XZyp68N/qPJzqv5VbYbXtA0q
jtbKZ6Q7EM9zMZeZW4ysjWxejHU/7wjAZMfEbMi7jKPxXoRc4iajQj9oZEnaBiNA
LD1Kr30I/qF9npPn90l5D1CnP9YHSjpptIOwfpWf9bFvK1SVLtylZ3H/Y89vv6KM
A+3RiiY7A2wuFUP6cVTpbyDBbm9EdqFX+7eO8M8a0nZ8Bu+U7W0kBk4brvYgRbZb
9iATW0H6eNEQzRlPWdWayZtDGCMnbOdm6kvMhAdU49tmCKFbht+nsT1cj52HUi89
DgxGFcEVmMNiaPzW8QtRAgT0Df40ct6UZlBZuJ+UPskCfijoCtJ1D54cmjmCiU8a
WZlon9Lo84MtPSiIXi3EUTKGSFBHxua+z3H7SSbXwNTrBawxgQV/brOebDE1rhvs
yaSlUp6zNm3y3Yf83l5XWPaa/sxTeQ1An7hafpM+t9twJ5W/xxuRYe13IIcKd4WT
hCfuwshCtupT5q/jB375tK0t5o9kx8zVZsuI9ABtZOIsKXWP2g+H83bi/qDdBi6P
j7DLWkn8gH146O7NgnLzhXAFfzXTMscWDsBWpfvXIg7wzAO2pQz6H6wsdhenuXEY
tjXwZOvtnbngiSahdXydAkUFx+7yQ64BPOtiB5HwHfLwqG3bQCjnUUHF7klqDUAS
Iazz4daWIP/JcKoHvnb5O6B0/+nS0gBI8ruuSsfXG0nC51oCqv15xt6SJe0ThiQb
wCTCNQ4ct5b9yJFGnpWL0A3at5s3GZBuGwUP1gQtch7F1MJuOtDlxhIYJm7HDuJJ
5d60BjF0QHLOvuwSWUQKlG5BRw0OAZDBkrPa9PbRbXuQzlulrGQOj3dy85dNS3NL
RziDF/qO+TkPsMgF7OwR5Ldjzm9XtCmGoEvKtmRBIl9Ts+k68Jx4k1sCp0pY0swW
CaWenvCedoI575OwqbHlqcRfPeKiSCYQSz3ZDMgso49uQmjvdXHWHZt6Y7mHufFX
EjDKsGPNv/Hs/ZPj4ZWnI8rnMllXPUJnhaEvpGNS9rfPP/7AtP+XnfRsZjAA4aEw
W3xz/c08AwttQaz8MSVdwyF+/6Oizaf4tTmbfZYLBW8olM1Vh+F0n4MRNfGnu+HK
UWzHRZOD0ZaTaWyBsQTozmEmaWRVcsrsIu+gHHH/Uka9t3h8xVUcgWMJ6rGYhZZe
jt6qBfwCp14Av50lZApllVevoxzRWG/CiIHNyFlktCHPZ8TM6a3UAgaQyLTYCHYZ
yZ0Tb/6j+R2/LfOMfK+0TSww+K5iIydR9KqX291qH7Gp8NITvlWttqcb8GbX65F4
1K/POSIpxyVfgdS1L793zkLxv/6tVMfvPEPGDKFc1guQqFZZ/l1/zjBIhH3QK5rT
bOmkO5SgK5ltdCED4injWUkGEd47G0cVHt1Fyj9J0WGIrxBYvGp+APuUADNcQr01
3XjMV8D5AOB7CgyuFdOHgw5IRRsr6qfmB5Y7UQ2YHLMW9twjWkyFu+Avpt9M1HKw
pZMWNkBXMBW4qmilpSJMSTWiC0aayPU6B68Gr2rnudwQBvhCpKfNvrj+nlaMCFhj
zW0XPS76PbNveErk6HYO8HbNyXdRPsqvE/p716tldagYYU9vvTz10QcR0vt3KhZl
7cz4/zMPTxwI+4Ix7aEty/vvqI7u3Oe9o4U54pYqOwWHKEchFnmu0uI73peUNt++
GgWDlVUZp5G6mqBbSTYFUVIjUvJMHXquRlkSm/Wf03jXxEBC5mgOvpne171nNr4G
n68qU8OwYJ3TLL+R1syrKHULPyCKWpmyCaf+4rtvAlnECJ9tY2WDeLYLVneM2kHh
AnshAgWYEEEKJzKeFLOrJw0qG6aIOQnGk1kHqwvn7xzprTdygPctm01/KDP0D6DJ
ttshPwFSSzbyrxt7Fyuf0NqyBKlnPZ2RWvB4CVLKxkWdlaVhgtG5UHdTSj3OipxM
/ok+0mZDVaFbzytO+3msNwIg7ro2LbAX1nNmoYmlRt9AS5dNSahQc/WyPjwQvy1v
YQ9ne20CdgHc750tHlWDkHyBJf/gutSPVQV409zJDvgE0qRVfYF+fSz13qsDncT0
U/8kTEOey7yYAE0r1CT7IIoEcTCCUZ92Dl4GWbXvDlMwIN6NWG2Hb3fIJS6KmADH
OVkhuznumZveTri3/bzizsx4CNWyk7LGBDrvtxHRU/4ASPiFPxNOqrD/dGuByaRc
gvZrS/FVM5FcNyeDfC7qmB/cBjRJcgSqydKFW7Nb8HMMTrzvrY+i+XOVEli8CRp7
EBLQ3a9DCPfDmw4t9eLUE+Bzf2yBW2aya7kIDG6DqGQyHyyM8pY4zfRqIxKvEEE9
jdWO3Rs5cRdINwANFpKjuwBk8LRDWo+gziseCoahiR3tWWPMR5zzLn3o1olcyYTX
YtYhV8U0z29F8ss7TjYKdIIsdvoguGR+8RVgMxF/dCgDPSTqKRm1BYo6jy/jPQ47
w8DWQFaMp/jF7priap9/YImtwLvYHGMNgGFvpyW285GR249ya8ZItrH4Q3BEhNTR
nj3yjNHmJ7KXUGGBFopnhdmJBtsuoynH/Ca2llduCgsbMOWxQ9oH+JOxMYdwFGNn
DnFOZknpC2zDlqnLDpLhpCxL7k9Abez7MgO74AjBnVX/OxFc89px+tWlLrpRk+9b
m7sPeOjD4i3ov4qfLxTD80xIN9DJdiPD++7JmhBqa6X43TXxr3ZYLepbyL2cTCCi
jcJ6/Xrax6tlRpvogiNw6bMXh4wSqBhHGxT9WJIl+PWMok8Pf6a5XRJSS/AOknsA
z4FX7RZPRON5SRq0xMmpu04M/dzIGDE2YJTlLEfG4SPIjAPVZwFxUjRDsNkClbK7
YpUGkgYkLr0zvB3NWVjd7C9tN3TzICrRaSrw3JJr8AE6eddbkPNcR4GwVAcKsDAp
AgBNoyl0UnPrAjllnU72+JOZFay6OOTFw+5ldyWagsYeYDs+T5yCSmXUXi/8A4qy
HzMSbCedhWtWWYoja1t2Zo5KU/wDcwlAew9Y50iAT06houhFj5w+lHINfYLuvy+z
qyFGQRVnM+XI8jASu9yonUaR1rSNLdmUmaK0eV3GSdda9sgiURA4IabjF7o/T9WJ
cv2vFMyTy6a7L1N9McPTeznmduxSbGIuXtaB+VVsEprpJFm5Hblhn5io+dAhtHxt
ATgGzGHrViNN+Q+4l16etfSv3l4pMfAAff1oKo2s8GknLzgZOd8eMOR2dh+0Yxqy
1LXo57MrT4BqDFhv3s7sXYweCxvVOHNQeiE1xkL0bUKyJ5vJZM3o3wolgIqb+IN+
fErG8j3nVSV0Z9NZlLR7iN5c4RJa3W+pwCCMkY5+lLAda8LDY69Xs15/w/qTIct/
+ye7j7qnAtWxM5nOvVfd8OrxPBPcPNsOmapsGLqbPfqvifif/PPHg2zVf02y6V7v
SDSKvZANRAKECEjdU8V3yMCD/a4Kk4h0BhAvJcs3zlosL7lCjnf4caV+41HTWtPp
j5mcQAjE4mvGHIOMIIXXzaI1qcSxUtr5PdjaXOozHAqPNV0X1p3ozz2inqKWbAbz
u9iGKMmUqAij84+TK3aApvK8/jaNXgMqPA4RGAnmD9f+hi7raQwBk6NCtLFz7faN
pUU4ukzmGVTnKkI16/vaGOU7MPIvc6xQP8r0D2p3pXbtSSUl29f5n/eppqR07gSd
6JYZ9P4+uOS2fARhrbbNNqK2syF9J2vQMtAHNRqU1ujVgRFojLexMSp2Ftb4Fhe3
xYsvFTuDmHJ+/JrqSsdb8v5JyBQf2pYprJ5YFJvqYwSK4QYMO6jSQr0CvTGW2l1Z
BiWLJFPiNao035dMcJBnboG37IxyG+OIiIwdvf7b8JCWorfedQRqtqBUCw4Pynwn
XvSdzlsXFl5cE0yWewOzE8gtrQEOiXGjHWHB+zRXiEi/eTpXRnZ4MWX8dcW/Ytq2
HMYyR1wvKL55Nn1/M5DMNnTWltTTIuv43C6phPvhLaGqN35cc8WgvBMXMZ5s4lVb
+S0IM+qD2wtiQG6CebgF8JfVDWcQHq6RHV1m2YC2w7608vyEbexM1pjnUEu+eiHS
lBok8aqbST+adqzx3P2h4MlSJMoqCPzC8tVb1q0FjAnJuFoQ/0y6R3ZAB5tT+u3y
LlbNXcZZg12BmFIiy1qCmMdB0+vMdbLFxTgQQXwa63Twk2UoyNHLqmDKryeIsEsJ
XIyWTcqp2PATpYCQoE1VVY4tb5vhx/9QRK6T6+oT4Iuf7R4BlCT+x5QE6TZWgJCF
jiQWdTUeDGH38WNWuQkfvEqHlb90rmohDfF+2/2QMUQKZmbNLbQoi1TXMh64tdJ6
eDE/V1mikJuVUUrWMv1Ae0yTSg68y3hnomGfQNtVh5BJ3+9m7QdmH00Rx2H3vCF2
pKF2yovlw1l5hBbNf2mN6A59VRQmEKNSKSvYYoKuUe9WFO2wfN9uJ4aADzHRB+Iu
MbeUE/DwZbcWRkqMkm24L2h7pdwrooTsMrL6sUM7i7Xpi9AddbwfNTl6OPrvvvuD
3fp+pfSoH3du9G2U1LvUOkqKk0b7xm0vk9csDxm30FNyqzqqIPm+kgL5BAbfehKJ
TRNAq9GKc0I0LaQ9rGynD+uHYUNv5flr6F+vaIKMAUcmeVeWesIJ+HUl+ARmxnxX
tE2eJ6DtZ4o1nKp3Lh7cUesgRiFhNhoEqrUtQ4dukOw1VITaojKQAA2oESIqTWZh
fESNUCnoOIQ+ErjftX/EK9xBdOO/qr25rphSjv5F0XksoeYBT851o80+9FIWs9D2
/2lxYtb5YyMHVUcHwnqEONFYTI04eH+BXXGA5Vf1jMMNgwn5SlO5MGILp01gCEc5
VFfJr9NXBsGjM1qqzrImQD4ESqEG01A4ktUHOLlugpf5LG2NgW4q4KBvAc76HOqq
yPBJlv05v08c5j9N4hMRKsOCLDDXVApjQuYRVgnpU3cwbZUjyWym9jR3U1tAtu2P
bTbeot8SVdTrsb29U9fFj2DRdIuWX/1kIW2fsg3AlRdWHQFu2eTOZ5TEfCF8qFM4
d5IwB9MsxFRPRU9GbaA1GHJeH8e7rlDOljN4F1HDmkpGYNNzpJ+7IUTnPEqiDmby
AtGdvTo+/8RvPuX4w1ZiAfW5/f8fDSLwsnzMH0JA6GDXyczlPXu8YZTdUfVCJE+k
EOlzziuaUFRofHOOtS4tInMonb2mDNS7bhvXOLCinTWdtW5FVuceBytARmO0Ylh5
ROoVDfiElcEmydJG9puCHvez5J5LAm63A79iT7XwWSfc9Y+owhVaIVfWfjrC7l1o
ypGw3JUWgSf1dbz7TZpqq3RULMnCnRxa6ZqHAUblAkzqpC17ZyHzGCLN37SAs5OS
qI35yTcr4thl/RaaMPejsakwXjviSP13gvn3czfALW75DsfNQNeQC60BPbL5/MTe
Is6y7cJEtcmAsUn6cGUhOsZALfFzuFD5HVVJOjrbfdWs/gqHupjJH71IBqOANdzb
JNSuSviW280hL+eYNm7pU088KO+4ZEnjbYb+t9L/f615F7CzkA2q2kUBGsfnRjFF
YyGhEwPEvMYA6cjxXA0hF1IexH9Pbc5+aiyTqhP1HOmLhy1PSKHfnPedxFZ9zd2Q
4AWplx0r9YjtKeCJaAScnV+z8NZaH9jfU9w61Ut3yoGeiYZj/hWCba2frSvuzEuW
vcB62oD/1GYuH9XewbxN87bMEjTKk8ur6p8Dtis2LYEBzKzBD8hhVyuLFJUcSpJJ
QBANUosoBHmRvG0rYjE1h8mbo/0yaPhsQjNBbe5qwHgOquz4x4iQkyYFacSu7E6P
3MqJP1peUQi6GVi00yXtHHm7rND66sXJnhLo3moWbS0yJ1xj3HTXxyttQyewKMpr
e7yDiMVKkBj/pjmhaz5xZKkmVZvQXfPhdEU6P6E/r16518ph5//cHsrpyirViqMg
jAzq/RdMWN1dIgh5nhCBEQ==
`protect END_PROTECTED
