`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDYrMvTImztK+2TRXADyhtk4kC231BGQaAwgbnKWV9zzQW/KvixVpX/BH0iQd0j+
nKau/fK2QgmEJzdIX01XxwPU8v0QS+huNIxNMwXJWHGSTfzuyUskNlguEUmTv3Cn
qy2KejeQoqGOWcmZtkibi1vb/j0fKk6Z++KLoq/5KK4fDcZQC3BwgDeivxBtcDBB
pb/WvrKgLQ1JUN4AZofmRc31hj+6TBVvsuiKcYO0WbtbWvSpYAFr5oAXz/cmjaHx
gXJaEljaVOBV/zx0EzwyLwBV+QSoeobvNZSBroIlw/HYLzV++Ez9dnkm8DWATt/O
3rqaCSUCIeX9so1GEgRoWj3r9B6tEXFIfT//Kn4FsOMrD0bFkb9l2A2puols1Tqc
JeesOZ6CMl+lB9J67ga8NkCD/bibTtF/PEo+JLB1O/7dxpA4c9FvernUjhJ2EtA6
WzULoGGIRjNBx/rlSHbzDhzihgxs6MZ8B63WVXx0l6WsnJAtxrgZz7f8HTCK4QwP
qpOK5t7b4kFPa2v+YRNV5IhXLj7JQpd0jaaeGi/Eqk+OmuidRPVkMecn1JPEyIvS
B8/hry4tVlDlQBQECmR4I6eft95YbK0ooK6X+LbGWzS+3JflxbDp930KzCNBcmEd
Pry6b0YiLofwERoVQ27g0mwKqwJEvciWGM6kqE+uuElj2+25C6bHOUrBV2qgcHIt
q6UuffEYVFlEgWPWhJ+ug7sJvGu9TrsY05849p1u+lNXiOVfGrXDGsGWQgO00iml
CkzXZGSzNGIZKEqEeb1XEbe8q0SraEIb7uXGDPCIVr1WV/K6ip8Z1FfguV1FRr9Q
evzIopBqo/KfWypnvpgTjrB8x5tx+UnCl72KYBrhNWajR9r6vjDD6lHLTTuTuKWI
92oOWt6jAF1+p+HGg2nsdK/izDCXkTFrfuFpP4NgnRyRHIjJfVgPwXIDo27rKeHg
yWUTBbJusq5m4B88ySrdpuTSbyBv8kmlcKsyxY+CtUPLqBDzN+cpUR54f01XUYex
QJ8rXcvVZtVRxzZ7Ie2l2v2gJuYuZkhE1HBY8/PVpv6Vl1E+qKdOoAhvLrjVVtbN
FZw86TRnlX+CL0/x1V0cit2j9qVpi0Y0FWvvgaydracO0fxXUJKRmlakq7Blhnw3
vdZUDn5vVVMTldudrkrY7Hh9RBT6iZZ9qQFoKnEKcpwtCXvfw91j2xkrCMZ9tFmu
FgW/ZvfNo8mFpksobNwpOr7Srj2+UiqgeOdKwZHWyuBRppy1GqyZzFhkqzBGBDAR
6hvQ5ygfLgfzUGe4G2fOOLeWgB8CGN4R9EC4DVlVtJ2wLNf2wFkSULK7+uV4R8lZ
1AvKlLQja1us/xnqxMqpbUPb6lljKnmLk99VzAFFCjMC8DLttH6R2fF1IjHOA8QM
x8PWsNfTK2fd+qmO7w+Vttew55O9oHiEChJv7+PWPIavL5bpa/G/azyaycZ/gGUX
LJgjuMeUIt+DNN6rbGDIMDcN5VmVsQmn2QKtzKE69pwZkDy2jRc8bHPGHxnwJo0e
eEcO0gBkdNBSVSt/qyQ4ZTaNU9O9C3wxL2nJfp5OQkSyEKNzik0sN6sdRzg4XEAv
BOtwvn3iiGNiqr20lIBcamLRSSdI5IAvbl2HCYgtfaU3bq/CSKTat5UzKxUSDJCK
unB68jlV/V8+TN66vq+GuOHKYhj+BBbBLj21LpuXHizzwcjXUOB3dAeBDx6sRTHJ
HkbT8eqqbf9D94+7AQwmWmfPQDq1vXyrL5OixKtE25k0VDO//Xy7DG+pf8/XuKm5
JYB9HLjcGye6sQSYXiRoZEbvTRMqHMWEMF/44EjcbWTyrytHiZoaRfr8Mm/MwtRm
zo6DUX7Acw6B8wKadVsG+D42mpxQaz/k/4m38W5jlOm90867aht4/796niQd/KRI
uJ1uQzrlGs9HucJ59NdLW+eFtv4bpRanzJcEDk4UPfM+9mRWsFsH49wpKyprI9/s
4DfId6dHmN14cS6muBz/bLRUiivKnb5+IPFGffunbkFJmcx/f4l9RgcqwMcTCyIl
IQeHCrHinih9vekQqx2mTREStnfb79unLfDPtYkEvPUqf+XJ+zlORpiOw7INI5Nj
Tz9+6LXemoR4dlqdMI8KacyyX8Lw5KfsIQ1cilE+JxI=
`protect END_PROTECTED
