`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8finiWVFobq/1MNXARvIdFxqAIdBxZRuVOypX5jurRLRoiLHC2J+ND4VCh8fFzT
FLh5c7n6ch/JWuUVGqMigUB25zL8SFZPF5TDstVrpLRbEc8XTzOA7lRQa6fh9SfT
nvwgQr/Bnlev974fsOc+VC+g2khhXaTEdPDW5/fxZBFkCipkigOXV5URReeHdbC8
jOK6ofVoKKuxtE5Rv9isXVd061u+QJwrctJqUT//wXi/Z/Xs5RpFAKWhVyGhU2qC
gr41R/uFQDfdYIgiD0Tj72E758EmEYJyx/6eLZNhlATaEwL+Ni9UIKA3N+3L2uoC
gLJpefT+4KjqdZhwrObacAaGGEHEwMMmUuWAqIx5MS48Vfv9S3GotpOj0fOjp8Cc
StbIr8REd7wttZCk23GK28ulrNdY4foQyDFdIYXIi/ggroQkEfjxyOrEQNJ44Ku8
ceRv8g1Uyun/5WRl2+zG1n09l9Ux6IQy5GreRf03VgZCsFRtelWo9fAgeqYQ0xni
HdaOgmIU1+Ws6gZZInlpjSjrmsaCBTG+HBgBBORt+Gxl9vE2XH6vclbJsymC6dK0
C+E+WTm+oQUQf1huoecAP7RjFsF8YHjHNZMjGAzISS0Vv5dJnyk5W0fFnSdi/3/0
z1lRMrtuo6+El6w8c/G7yPfpbSjG1j0Y9/EipSMvgc89Vg+MVDsYuUjEaLFHI2tY
H7hE+FfATQg2V2BHk3RU862h9tHMGdt5xXUSTEWG1ujH6OTXS57rRf74FCNmd13B
zAVg1jw8PRh24ntoZX+ZHvoeA10QyxsCtBBiznr2MkjQ36zA7s2ltE0CqeBDwrgg
tbd+NEyH5c8JuqkV4q2THq5ZmLBaMcEIJoq9cciwZmIN1Nu4hy9gKfnKKHB4Axop
QirG3DNDlqsP7VO+Cn8Yfp5BT7eRUsH+NQGvGFqQE/WImecyZm1r/Zqc33N9FJin
Vz+xXEZEqLabZlCXkFkqJR/kPoSECje+JXvQTez84qPJDRiCRSDdtjMxgj3fFmeG
tya5687iWZgCB3GyJBYXb21HkLaYEkG1qRCcycj+6PsfQ+YbTP5gM1WkP64MraLx
Rb3i0HxTgWl2KrQ2tH9fa4GkC6ML62ELe/QccqxAEZGWaOgN5qsVyh1d265PuIEb
WEBBQiVj4V3AlDqUXdO/kFIPhc+NHShZe1Nlif7uiUmlKLuVC5/b9A9kNAyelBVi
Gv+/SVytdWiFHOCqJLRbTjr75zQg63rLQjYejzjjTkfRRqS9gKJDmJWuZfat0waJ
fkdD5rDRjfSv9rOWTGqYE9EPRLSpYlrUgai45jIjtE1pxUV9UmAIOUQ6jwpKkZdz
sZ8Z9s166qpre5ipwvs08hIBgAckSBPkjLCCzTmGYNysyDKbmRfuj7xsjmhJPEk3
YxctRTZJAuFfvEg+mG4gUOLoXWn9ghZiv5q4VqCnI9TJOYGQtR4Yg6kND5QsjUti
UpKCrTIW2qsRJcKDWB6aYf+6OqCPVl67bKLmN2QClZAteSlYMc4JmyUmWwFirGRN
gw65+T26X/pz5QntYXIILPT/HbqXEkYgKYZxiw/hC/zL78YpNoXdG+P/43eixkTr
/N55/UO1erHrQgy13uwFHvGGhGBOweThsSKBwhJ3ITuSZ7rd3tmNzs3AXinMyQMe
JBZ4G0BqFSX7JowlZLONMsrmFr/Rkr1i0uk9TF/kRhIOGoOLLNiq+2YPOcD9kB5s
EDmJWdey9IbK+0p3lTU6ox2N1B0+tVX+bzEV2FiBqxE3hJOE7x3P7oZ3sBUg7/LG
WS4pksIs9tObEVl9ER4dBSEgvC2oo0olXZQ9fVE0NdIywsJbOnzFhPDwTrILO5Xx
dsre95RcWkPrY5ZT3SKyPd8fEh36Gyjp+5xIAvLpJf2glv/Ft/I+sGGlyLUbOhna
3WjFbaqxEg6NanZ8Vu22oTMgy/eiTr0mk6T37uULdMkZ6Nl8LqP4pmvqfYHibQA4
J6/ri+NQeFYAH8SLxQ0j2yCxrvWrZaCIbwVglofzJqGcdTJEHeHVL2RlSDAjm75T
6gzL5U1UQPwmawspDd80BfLF6xXwK6XDa2BfgLiyuLY6hSzrXLSwS6W1FU+iOYaj
otPdr3LwFdhICLi9JGoJ3ViUJ7ZhjeDWu7QK8qzpUmwGH53HhD6UBYhcQ2Z6W4zf
CyomibmYTCzICSntYCH9eEps1fn2y5RasaqV54/Dj5PDmRkzQAzKjgktbgl1WZG1
uYZtDPcUyG7MqY4EJ4+pBu9ajtxjUYtwxnHVuTxHg58cX9N5WZYQUzfuU3lI9xVE
0p8k0oueV6w7D1jmL/bKqqfhmUzDZ5E46HT7FRWViT4anpVNEMfPM/UEwPg0vAOT
VG5r2I/3sFilNgtTLNLQNID88Gnye7puKYDPgCRSMGWE2ZlqprIUAezVJ+4KtGSK
vMERLpYRU7k5SqeM4a8pEF/H1lWG0lX5bXybxuDnsbFqVW+saVdWRnnL2nMrSMGm
oObhjkKrhDfX3gli1xrPJi1/spKbVPWCRtntOhT8mxccEPb4k3ABxSW/r7cj6qZw
QwmEj5xaiOxhZaoAYo/eX8QYALebM296fdO9o849rMvqHlTT74OUtWCBPIi3Vf/q
AMfZ2DmMzgMslSo1RFlcxMB/BYVuOqYIY3kRssKMv/OTwAJlwwEoLgrdtA3SYWik
j4oH9rMcfx3orG9FJtzqN+6EihYVK06rBk+qUNLNgzAJoVC3VLlTYXxvZHyGy6qt
tmhPugun90w++I43j+YcTJwub/C37iDJuFqZdyr1PfwlwjBVSuQkevhpifvIgntg
TGMXen9YQUP7yuCuL43KKd/r2HYjdxO1TTHzsKX1xdWPmkF3cMTD1T/WAz0WqjSj
yAGZ0k5oWBMmBkwNjhrACkx6ujEFZZR5QGAQ3K8gUM1UuWl97Yg6qLQLxDc0e++h
93HgLTYRvStY3EI2nhOFVkqG7c1kE2Skb6/n8tLmymLNCmt3UHyYXkTBL6dZC0B/
64F/HxfZVIWOfNuxxtFz4/M/plk49jnLsBbflChLM4FwDP/23UvDTUBm+zqMatXl
iwDdosM8NYvAfCcOlR++MHXnFrCIaWVBXhDwXad9Tw5SQDevY+NzhMJCJq24eu+5
ygDLjvFwkNrbqueHkKPObXZsrwKh1EY/LcrmKR6k3+IuG/u+Ci37ujGYBBUwo+AS
IKhxFHFvvl/Fa/OdceWzkl2eYyrqgXSoJT0hIqYwdhHRmFDTrH8eGew71Bws5bUP
PKIawlfhsE6ubFIgjXoFHxX8lqXnAdjdyBjsZwd2k3PAGuj2cm2aoFDSBg9j4GaJ
LwihYmKFNIWBR1+jhfL3H9Zd+WsC3Vx7hJM/GwIeNNeHqR2rS3FfKHMNnICfynVE
fAeOyJ/lyzMkQEOj6QJuOshlSiO+fq9bTb+Lf7zD5seAh+7s0ad66tD2w9N7L0oo
B4Fp8vyPqqeq4j44sVP/OLSULNE7JWhVHq64FBKeoA4q5nFrMIWUY+J3uJjfImYp
zBAwwHtZpQxpJvwgSOv049Ee7yZMsx/cJJD5wdYfp8BN/z11SI01DSWD0LCwBxou
Li+tEKE1hPOn9eDmzIHgKvvEVe7hFKDHQiYO0gj2qjIaeYGwLUIemb578X5XVFKk
2dfLdfmh9JJPfyZB+WEfhZmaCwjeDMjLLQOFScLtqp34h6oRrTxUBONwg+IKhgtY
5/24nTVeYSYstnhtArTKODWqZBhZ+np5JMxlsu7vQWnZsOsOynxBGUSrlvfdTpOp
1t1P5TVbWMGSl/iaVYV53O3VUKdeZI89AfGe0E+aX+Lig3LeC6dqSm/BnHCDhqiu
fb7yh8HeZnX7q79yPB5FfLj/vzpD9FWXlhxODzJX57P6MhDnaDgxc6SIAaDFufRy
ymTKEztDLbSd2djwLRBz+gVVqN9r9Ak1WDLH7AyZIlcXcK3zAHgXSELlsC87CjST
g1JBnvzW7xh89V8WMsgnFpogI7itVDOxSg2nA71zfjHd6H51BeCddUTfBeu6TOOF
QvVqFHEaLxAH/ktTN4Wz3r9duqJkX+GXHYTXFRMmUpmuqyIeIWLOnkwKeXmXqDsC
`protect END_PROTECTED
