`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZ7f63PFetVYsA0XpSnUpudIaa3Wk5te+r6XrE3fZXTWJCUM46AYuf9F73Ak81O7
7T1IGP0W37Dj0/w7XVufF3loSNwi0cRU607nd/5ICrlFFuxM7OLsR1MV3rlmBnQg
43zLhSgVt2aEPUP91ExilwnNcKbU3ik+2nVgqPk//gIBMpb2KiBA7yHPdhoSSmF7
/CILBbC78Im3QEp28r1Ppt9kizPXzEplDi2nEvUVCjdiFnM8XBoqWbkAg0Vt08S6
8jQY2af0A0wNLTGZAXHqzqGoQ/SPfOQ486lxElVwKha6S0OZCF8o4aknYgiXqkMr
UygqigOGDDzCoO6ChZfaOWZZbBF934XI88thrTk5M+VdhkU7jFCIjfYav50wTDYN
7LXWUXUv7NAwJi0mG6K1UWy7QesQ6cXwN1mKfzNzrJtM6Hu7aJfv97EYMPpH9xTA
1LoP1gOspnER50dODe3c3xiPkDCv0JRPtz2DviNiEw5tqVZIWJKbcG2mJiJpMr5L
FrIHt3Wfsw0w69uD8Y5IBLEUeViY0CLIoNVFCG1Tzd2JOHUiAD7T+zWJuB6iqv+I
b1+CsJfl5P7PfveSZeJIH/DhmhgFPXbELeFCyKOMyFQbReemH1jE7dTTFU+oZWxi
zefg8T08DgCD+VFM1OiYTAGDAH6iRgTc3/N5Sv31JfehYUnZyo0Xp96JVUKSVQ0a
53yN1YtHgob6TSwP68hj94obp3iOL5rtsGRKOC4ICIWbres/9NQRtCDh3i5jpJVM
TyUcWROnSBeY1vOAyOtcwdFVGKUaOmNB4o2ACGXDBDWw9ZeyqldCZcnlZuwVMgab
s15Tv4sowDbbrOxW+Ge5lBwarVUlNX5IS7qUnFBoahrn59ubWnkoi4LK9PQTSayi
dNnrL3Gr5nhRE92MZX6Oak8cXRa0m27ijlqQYZ8ltX34ysc3xcn8TM/WWCyCr3R3
RWXwfcVuc3EsT1BPt5Jwvys3Alwe6y9qQg9HysUb9hfLcdjziHCCNvNHbABh0yqR
wfUPbUlu1R0d2HzcQkhqXj1IYN3iijTUCZm0HTKhOMFQ6i6Lh+t1zWcabofzPgV/
nScofXq2FOhxHXcy2oUJEVEdapSnqhw5EWgJJX7/o0s2R82uj4U8YjmjXWFJSwZT
/hri/tAryN76m3FhlNhn9hxtHfWQWgjkP0V0BYLZaDbnNrT5Ea/dbJ3PNThaxB2l
xSh2fUf0R4k6Qj9ahowj/RRAn5LKlHULppHXXcQEWltOx4ZHu2LMa7mqA1y+4z75
oi/iO2u5t4uydmMjdpM+ihffHPuTYNkXaWi2y2PsEJfwPx/l0iRMVAL7sFYDPyOR
fEwdTUhQQ0RZxSaSLowcxTuQ/HMhm/VGQjhxyCCy1csDx5WBYkTF9P9mJJVGQDt8
OGSNbPMK1/VKK6lwhNGkgsdHlX9Bke/eqTK0ZDLkDUmMTrOLvgW7EBLmLqO8vicD
gEIRWouDMjaZzwNZxDTZN3zVRjfJhWvVGuQIbe5QP/UGDnDBeGiE2IJM6CjqrOLa
3g/hnRA+6X/FfU8FxSlkcwBZBg5sVFz30Zrw43/0ujd+L63WQtUZKjGu6aAU+c9/
xOoNAoBwnba7k9jWMfdkZ1hhs3nNJSa3PayvdGZobJLs04EIXFDOGcNttLy2SxPR
jAxhALIPfqec6l4h+E85Tg6Je1h+pX+5GY4ZBQjfMkjEIVqur+Z0Gp/oY5cplksD
Y+mCz8/3AmDxLuv6oitXobmo/F60CJAiAo2MThNwWqb3Ut9YBh4ISpFjgHtcNgBr
gkDGGL9xEfhr0oxHSI0e0hn4VbW/zCslbluFjzX1y/ZF+U3+Q75lPZXOqvYTlvDi
lbBbsFDr24jY3FvEE/cZ7bOyrAxPgGaoTi6uEK2Q8Rk0m0VEtwV1gtP+71NZgYNh
qp6+y780aT/yPrjcCNdGe59G5Ib08h3SDGpEZzyQCSm0Yw6i0HCEDTAc0c0OInwv
HhGNUN96ysIBrwokg+zFuGiqbEkXxPIAtxyPgGgeHwsubgTK5FaCoMvvKi6w/sag
FFySGoT7KxuW+ObEIyicWZNbEvwnyhrEoNSP6VYQ5lQkiaIhvm+HSSX/aIhEQxM5
Oj7KIsnxP+9L/mPPl3AoSnWuMnol44tsqK6yugDRFMWgeWnvelNzMaiAxHQ1M7cG
S/OjQj/CjnsHiAEd78kXAwPbVYZVs0RoHtwxXZrsaUK2PVJ4y6a1AZZBC851WKqI
8h3AiCs4yT4+m3N6ILA0ojEElv+S82xRlcXhvfxS2fcTtIJi3cZnUE3U1O4DPGpA
M+LxZRbO2ZYDOzjoehuNNX5Z+E1WxoTysoIT4CMN4wSLhvHTionqQjdevqiHeFpc
sdFA8dCsO7G8+5NoVllE3L8HnE1nl0UcsKAJwRSf9WJnI9vRCtVH0Bmr336t9uUH
3wdj1WRuSO37S24j51jSRV3qItzw2A0qjOL6nmCWOKdJz1lDl2+9ccM6LreaRDjE
Lab0Aeak0+pD0W3FSzNpqVLtZk2qjfO3Loz5a0P/VFbsUjFHMHlEDS0rLPHAGvJb
jBozlPoP0/UElrzBGC+lT38xVQAjjw5MahMeEzK4cXMoAmtijloklLfkAfF7c0gU
yABaRs0Vu/NQrjn6b0Ty3xMyHjxUe/bJbJW8HSETDsXiXI7kZ01HMefoeH3szJH4
PfPunt6ykzkMe9ZTIac+7dXALjXzDFjH9By1nC8fMur9w+TbxrX2rCu9w22OhP38
+ckIHkSqswHyNPqBoPgLB9WTJzdQxQEU0X+1IDYkcV1lQzA+ppJdlXV7HXPKFpdv
7wK0BuSsC2yswvKYC2W872u3XHURLbbT3Wxo0soRmmI0RrtNkM8bXgAOdxlQjZZR
Wi6+MRS8uRLm1ngeFfeYji1l7FCfRL3SyBGV7lt+j28qu1KKhE16TnSLggmToLId
mPEUL1gavXTd8igghDlkFWGzGR6fFgOhv/HMiR3c3JY1Rq0Jg8aGGXDrRt7Pm0rR
3Z3eMv012q9V2EfMUkkfWa7Pu2psx4TOLWtkx8qR05l7IOaJ5QzXB5hkvDeH+Mm9
VxkAeGNmaFJabj4QURTz1Hyk6dU/3m9FP2+HDcnyjvFgqdJvWcNoyohGCy6jhnrZ
9z6jLvotOaDQzPOryO4f/NsjJ4Hv11Htyn4LQb9L7mA41w+tFIXSKD5jumzQbyM2
3Q0r291cDFyWXg8ARRMIUL8PZR2h6OEFduqOQ2B+aMOxkOGDpIYDOZQIWkyOtXe5
pQk3oTNceCEVosbKx+37ySBZabFFfZPh3Vzz20KubaGmqy4bSh/nWwNVvEkbT9vG
zQyU58XhR7LWAZ/5nlzkFTpcpMbfeAA21s9nT/wQHu+9hQF0XCq/FknRxpogEdQ3
mhZZsPv2mpro4nWi7qoe+RYgil3/xjXePUWdfDxpfYlDhyWhXIw5C/LZ1RJyNMBU
YwzJxJnZnXt8T5IhOvZy03xQYISJfPTfz1HXnWNKsHwanwK7yGI8gvHjjOAg6p9b
KCveAE3Qx+iEScCvo49DTpcZ4ExBKzcHPJV6fBTgQ1B+gxW7CvJLMfY9cSnyCbHD
r0ZPwF31p0QTIH2jAtDj59pynshUlfEGFm3v7hz+6/L/Y/GReeQH3dpehojuJ7SS
1TTN5+I3M9rXUsq0K7bSegPDniy3zcBrKmkrLRXTd2wC545Av0gv6XkS2Sp2Zoka
8oL8X5geSPLePsHzTgGjWn3+4zE+dM355rN6d0pSlHrNLrtEIOp3M18qUSz+15H1
VlTEBg0VivsYQ2Yzgtf/N0nO4hO2t195USLC/qVHKwmDuyk7UNuNH4hKHUQbPFdo
MFdCqBBXTW5ZKcIEyiTa4A3N8FpSNALaX7svuORHhEem7xMyf1Ss9YQEsR1oFxQE
+adbwRwg3aVtr3R9ZeT7mcQYk7sUtLRcMdCXXeWdrkAs69WlwkiM1idAY07b0Su2
NlJlDkF9QXzCwQb0Lj4rODmbC9iWjzkp+Xb28gy+WCrxl8Oyw5m1HLMCuqjwW6xj
wu1SmeaNNPFnPAzoo3xadR0mvin0CPT6sKk9ahfggvrpqG2lwaehEFQiGbxXbRTI
`protect END_PROTECTED
