`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHyY8WP4LDlxj2Mmb20GPy0D2GtFd5GH3MHmOXpe5M9WXgzotOfDyQmbUriY7j62
I/gJj1W++zdVDV2gJDkGmSkVjVwIMPIGLzfjYNdud7yIjeFTCoqGPhJTlD9BYN5R
Xel6bs12QqAJ8p2mkrteIesDLY8w+z4hIBloWntWhiatOZx7Jv/yX6sTh5gRIVYH
rA2ny6a90HByw4CuvEHE1GeHM1r1QbiisKRQ5y6cVLPDo9RKlLogYkBLq98Edfw+
0JbM0557aeBDSiOKwJ9gB0bw2n9t0p2VrUuxWXAVrWYHks0H+sQNL59dWUtmxx40
ctx+QckNITXTaSoKr2lgpz/znESA8GIkq8pJ8yeW++OaJqFJ06K0tRuYh/GNSpUk
v0S0cds++AH5OnbJh8W9MN9zyQ+gtbTjCbRb7Lvf90iR6/glVp008C4OTBocVEB8
Bffl/d2/TGeFBPLswVcX/mTq7ArBt8/t+06Wnb0sfEqoYdnhpFvIhqD9+f62V6h6
shObkMsx7FMkoxqzS3Um2bvMLkij605lYwMjlgurUL7hVAFRap65UQJZGTgHs+Az
O7J7iYdXfDZcbKSSyn2t3ALGeJb7s5IihidXiN3HeBmJ7gYyK72AWcWwjuvzvOAF
NHnWo/JT72adPmjjiVzy1bL+Kr2cMsh5YMn4gau9i0VID/PvcqC01m2oDdDmWsvm
gdyVJONUY8fdDfSG3BWoNUvulYSBdPxmcBPtJI1Uv6B79I6gQ+2cFvjTcMIJ/ziG
mRM2tjgHZuu3fOjjPAVQwSIaaf/11Ww31BHOW0U2BiDregUtFy5Y37w/ZDV8gGD4
fUq1DF8VTqWNK4e35eWWP+WU9nglZO7rm3xghx83rn0fV2+Szi9dFQSV2pOTxVl4
a9YqiYYBzRelEsachRl31GwKSRI9xpqKOFpBS9xb09wY6Ty89LCdITpYF1yADa27
0jTeBP+a4i/KwYxGsinluZcXKt6W7Sg7B7PUSPDnFGHICppk4CMzlVAyS4Zma04M
+Wf8fYkc/MkyhQxreWX3Ow==
`protect END_PROTECTED
