`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yrirb5vNcsASV3eLmDFhQFsfz532mZ5Opx6mKeEsG/oNWYZgDwysyPbOI25yw4IP
j6WUwKp7dHr3vg8m2jA8dJQzIC+PCQTQcdnW57bRhWCWG+PVGasfLoEoZ/Kojhdd
Gd8IyXrPmLJAcEyz6sUjGJg2AbtzH1sIk2AwEI/sTegfnPKtD/GzHN+BeEZBTSWm
chJGIPU6D45Ht/EXyDrinVnu3C4S+Ov9I5UK2/xOC7n9BvwGeKvnsF1hGPI8jVWm
Oi/DNbn+3P9+weCYZq8xYUiqh7u6GQai4sdy5DgvSEa38bvOLj+VEtUw1DjJda+o
+kPcEvlL9B/kYyliiFUSwlT3ouSshdHYvVPt84tRqWK4CYv4aABUGVxrMkF8IjT0
PU7wo1OtwW0YM1vnl7j57eUqAv+irTrrSScT+OC38sDcmqLNQb9jNo9gRTide0rf
8EKNREkvdmiKzQlY5cK832/Gyk/FxdENLkJNhKixNgBzQvt3ZaLGCa4PTrEQ/oZ0
GDO5BXOyJ2syYGyqjf9TgeXMOtQhdPNghXev2cU9vm1GoXMuXKDyUprDzzaAzKz3
I9+n2jIIGK0a2dWiSjVdQYp7DLRKHtRnlPfIEv0lBwwxgTr5QKp5hY4WmIXPbMLg
tBsEa9jgMTwcoYM2Nx97RuCIDcKmuPJ/TQevVaAQFTstFzYG4rMZF/K+biQAjKMe
GhUrww2A7SnRhAIrejXbJ//tkaKySGsoJfVyl/5bXtx+N9f4CLlVhAytfkDDaLoD
woZV1oi24U1A1m5Eh14L17HASEPQKP93KCeM+qO6/2R91ODsr4Aj3BOJJE2TGrg/
HaEZXxhSUmkb1oz0eIFtKA==
`protect END_PROTECTED
