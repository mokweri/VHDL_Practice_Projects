`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2FTg0n6njB1IGs/fftWmIB13UgUssC8JVn03/Y4q6a95RrMNi5LZMTwzf8gmli/Y
4qiKP9GkAnwDjZ4ztDIrfcgCwzaZlBp+k/jQOlivIYWtU92G9RDrzCykk5fZ9vVt
OrRyNm6RaiEK9LVnyMDvhMnqs65FgXyC8EU8mHmXAuE=
`protect END_PROTECTED
