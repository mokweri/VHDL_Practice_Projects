`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uXaHlOkCTDjP45KTvZr2lJu4jHloAFkv42RwDvmoM+TiUC9fxhDTppk8QgaGe2IV
Q8ILQWHAlMHXoq0T72wgmamMzqrmcd7/103Vp8yYd9ZF3oC0jFcoqFTeqEdZLJZk
aKNq7PEyUKNnwSml9VtfhR33NTojYj6FaGpsVW2nal9PP9lbJCtiiHUOxvtFLWuF
KUI8x8l/YcvYNYjhmBURmNo6v4N+CpEUCbJEpAS90j8tldKPYUDpk+R/JFpWYA94
8lan5NxX2LJ879/L4R6MI0HWN9rEwmotDRcTkYM7ti/YA7IqAW28zxmF3GjK2ej4
t3aPmXpPWWZ2zLp7wC3tGpMsQU633WjBtlloiF2IJGGYxqs49LoYTOGew4ZMgREN
MGeGRe1lI597ZCz0vw4fOcExe1knszcJjBp7PKMiqT8NWog4DOebLV06o/Pfivo7
2NiN6SomdztbYJoHU2VVByr7VvOahBSsZNW+IVvoHcEmdFNbhc5ox9GUddw/an1q
kT2H1upNmJRw43zeV31nV2681yfcGlpwXwOsMrJQP1AzJ12myZmqadC/toBWwALG
mk8J2sY2n6BbneMd88G90O60RZ3Y4k2+Hcbhj9FR2jWmT1Huafd+ZeACBYX/VnwK
RBXe+TSvuznztec6ML5RMdhvoilg3MA48mHfujMMxsF4hNE41iVd6JZqod4DVTx9
rRDf7EYN48WJ8bX3Itklst51FJyGYvluw/SPnT6sm8JD3eReje8K1F4p1ta2uxtd
EtlGKncL1Pnq3Es2OoWa/eAVUV37iWV/wD8SDAWFm76cEe2yu57BiBlem6jdTLab
PCuSa2gXXEqSBqJu2eGDgFfG8T75uKJwfk3LT0jbE0Nh9fLR8/0NZ7ViXgVT00EJ
UHn/cDkBQYh5HtPdkA+Ek9d8U3xMhal+qWXREKkofDoroyJQvzwNmB8rJkhB8wc0
Ryhs6RHeLZJoTX7AlefhZOLejU4Gyt+mWq8whhsG7nCfXTtI+Zlkcy144ukAuwvV
nwha3qPuPMTEr7rB3ibocTsDO2sid/yhHLN/vqZq0mXYF6vSvyBUh4We3mytj9gV
Ci4VY5tUaeTyZGOQadOHt2sV6gEzxo4aWJGQW+MHGvCK1WNOC2otK9lCAiB9YPnl
kOeAJSJk2pVuoAD8KcAhWwRnQsv2upgnqS3+Tfpx85r/dysUtZUsD2mfhqP7i8dU
z0ANT/EWafuaTHWj/ynRJ5L9l30GZDvS7k+1PJ6kO04NnBGLgo3p+EC3X2klD2N2
bFYQHomAVyHn+nihdALinUYbymwlDiNcHHs1sUXaM1JMAJwLwAk98VLr4UqMf8im
lkct9bjFeueIU8ikEj5pKoDIj4mh0PGKPN6igWjuqF9WWS3enK/w30Rc7Md9hKic
DQWUoSnv51MU7EU98wvmFsZ91Cggnd080QeDwPSIcoST7Qtek1p9wO5L1lznUZz7
q6e9tyiT7pcP+tVnsg2EaaBbGbD+tpZSp8klWcNJ2Huam/+uYjpiZc/jj1xUPcNc
65hDEUn/WbGCdlckpAKFBIV254PK6UkfLBi5o/4hH/SW/tCDEESngg4HT3qY4uf0
Qm6Bl1XHDwT0YvcxfTC2fCyqB5T3SJXRJWQcs4eBLM2lCTMo5OMBbGkhppViGBgB
czrPrtgq+z4TWmPNJNnfjE3zjKCtR2vkXtTDNHGVodsbKnLt3W0SGX9CSPL3zaOy
F39Ha4h2wdJJ+aXyhG7H6Ssu3P/lTLZvcaiO8CGGGbWEYk0ktqAG9VKaIOJ6z/sl
AUVYnI9WKdh1qpejkuJWgacW4mnjv1KXYQeOdrP8DOWgx5NEcQ8GN2KjwrjUqi7e
Y+Ky84hmWw69sJiXeBATjVRaJ6g4XXI/i06nXV0IlZwK4QaAQAbyoST17k6uVjLw
Q33zbC9bgBLag5cxgRFQWCfY/Q/667u1gDDKFVCsUUktCokuEvC8GqkzIsXdRijh
6nH2KDVZLVIPTkod+3efPj4id8LfpLlDJPe3rfk5JD+CjqZT6dSnd1qW05cqJayL
CSAeQJ7r4FLsV8bf0dHbfRVSelZYdLgiQhZCTprT0p76MzBdJwe1A8DY+3XW3XM+
rnoUZzezm8RGNv58VTR4Dk7MRuW6adzEDT4R20y+BHUmT5x/287OMDvfupfUgV6U
7lNuI4GT54DgqR2RtRaJuDshmONlv8OYZkyHA/9u6WrP2bPv9wHyRO5krt16ALfA
+We/FAecLZcLwtaUyKBCTQHe7b4bqZ4uRlSnUIc4OVyC/dnH5FihiVMYqNZZQxhG
AV0CeYL6g/G/LkCzJRLRvzgQa3r6RgvkBLb+1OcZL9MVLcN91I/1KuWk7zxbwRsl
YdQvIgDacdct1BL7wJiKbjke3zmNKDjyhYceHHSQUdtEtJLx0MPounzVEu5b1Q1j
cDYNpWJ2YnFIKzW9KdIBaJvqNznLQPZ+TaWMdH/g/rRPJWYjq7UhZ59fUTKlGkDo
rAsWnpGhuMqBh9p4+nzSzOKQtYQ552cUjHCQzmyNA6tZ9n4Lm7uW7a56Qy/ea8/E
nvyqQNBBbgB9AxiXvsQYp9ejbDDajxogayafgwtNHMxHkJH+IElGnApIbluCt7Vv
AKg9LVjmleAv2tSMw1hhsJhZ63eDltA7yCVV81cFO0edU+2OXk0mhOtBwY9/a2fx
+75eiILgqfzjo+VcSaxTuir/MOMO4JjMbOEIi6rkx0HAGAnEkHkjKhY/BitW1xpn
qrW8nFKM/pHm+afCmdhSgUJNMbGCwuktgHxoLJg4VNDPX2uEWG8HjQ0fytkWHCs5
pFu4mIHsaL5INO+2tFfMJ8bMJfcb2VASaeEMh3LcCEekuRrDsAv2/rVp5zCtnKZD
Guph8ESwZOYSDj/IQinZmBQfyJmA1S++uLf0PwknIT8dDOrgWdlVh3Wfp4K64/j9
OVBacRfQRet0N/Myd9+p84ZuINAn4Mi+20847fImCvs+ZKiDPkdbTD1m2kr9WEIE
0wkCUR2SkK+f+Q/xd3sZEcNVHK5vSiVsSd84W/8Sn1w72RuvkeECIy8Joull5t9C
0oXBV7o+xFsa/tp8+X7wkM34G8IhEBIGyNm8t9W7V2AncdpiMUy2clSmrVQaZl01
mWlueb8/G+M6dg1d6I+rMgTew7zRTJp1nIkdq9fucNtkl4vhSPxXQ6NAmTmcupT7
Cbtc3jAbOR2Br5bcNwO2uP4tc1Ilg6RxqH9URQhAe5gqvbF4PruUc/Jp0bxR1VJU
EwE7S0RN3KXOricj5fimSAMj7Hn4/KC1CKIimqMyIdhg6gS1iFlvmnLi2EcEZ0kI
crGygqGjD/3Z2M0My7s8IT0utMWuXC5Sd07t+kB0dAzaKOcEWnu26/+XgimJYOEa
Y0U4ghQCZIYPmL2vvqrGVJzElgzXAY59kOtb3YxZqZpFWEw+7jWr8nTzPZlw/INB
VNWQdCWGyOtYjCVdFV37xGFNyvFO1XZ+YZmglR7/9ZzwYVZWaUuzYel9i/8gnloc
KPzUmy7W13b14WWSXMRS4cFcyEWlEMb42HgnsmaQo9e5YA4qrPU5SGvoLKvZZ5C6
buwLvTWHoIvI8xq+Ehp/QwFb+6YnB1wbFzUk6GleWOtAqNq1LKMMqRKBjMS/n0Y/
5YSIM5FT7q0WFSYWjdA9z60siTze/5EF8TSCTfWwnpcAoJJbaD9JF28IcVtnIqfe
vZYcbbRhAyfVIirwzMsytSoqA0dzxCvU+qVkzPCK3uDayLJvkrnKK0Pc5XJoT1F0
55cSkn7Q8keOwYwgdsabHh+hqYGvb3z7bQlbuh71LOdDAGdK0Y0FaaWZBb3ihcId
APOvEDgO7V/hewvez9qshRV69TmDvxFCfHhJ4dv2rqDmw2qLac/F4pXrvaQbWIwy
wI/GoZNM+6T1fCR4BwcNcQokXBED+gXUf8qjzr+06ZU92g5g0TO4nfqo8RdPL2/B
1SF/86WCL4eeR+s0WhGX/g8bT8VNfrjiVRdyrNKCN4/qrNQLY80xgUo6Tvjfn+5v
7Q5seRFJ1YCioXZUxPdDQtV6X+Yav6Vc6+hDheGziGNwjFjl4MPwhO9nzHoEIoII
HeiVe8xQPi2o3waGCPP2uoNdusaptxG691FbVeJJubBPt7FIIUStzBHYHKqVP05W
dXpdK3NF0YVWfth8/7c+u67HrZC5qMdhYfYW4ydEynteJbp61iN+VFSkHxRgFuWE
1vjVEjkYnYXJPzg6wOcJcwGDMMduPZ+8R0kRE5xu2FOC6fbq2Y3XEAsbnrYXVPHp
J59lNbcUB9PWwbuXzU8K/wbWqGjaKL41MTxQ5Sb8Gf4smEVVWmLeMMNE5cCPvNEN
IX6Qu4XAUh6DpUPVkr1+dZyYiXT3Goqk407P/qHQtH8Gh9L4TmoUFENPtTayrR+q
PTkE49gME5dl/CMM55dpVxuyhzBLp6QFryc5B6gBLLRQgcttllq/VmV7f8QwaFkw
sYbAO/KaA/86jgEtIuwZzgvkz8eL3BkTeCrn4IWDldRZE0bhQDRQAWOnvpwYJRWJ
6pfY6/QD4NiI6QATzIVIcRM2Q7B+WWiIqx7wNKXB5N+awVNtRN6x7AQoucp+KiXN
QIXMBIeVYDc6VMuqawCAAQge++4h8wG4Xt16LKMoSiEcH1xTdbF6eRhuDJBpIWj3
nSHSwCGDZw6RwERql3qHlig1z0+6HW7TrFv1StJZ4JRKYVTui2/YwsAU/KzhVjW0
a9fNQ/4OiWExDyX+nz9rHQMUNmqCIuGSn72xZD6xSjblzBRFEDhP0fuLTL+/RL+C
7QcsVPeM8SjcXTU0xOokusiC/x511OgDwwZ58fz5Oj/CraUPiEllXHbxuPSBfXcp
Git5iVzWzF0B5uHW4bzls7Rc29D/Q08/WFP9I7jV3MRxo2JnknleGHhawY4fOauG
/+noMHStIDy7Iv7jLRqocJbn94U6tcJe9RgsadMD19xqA1mIfaB6M59ScrUvvlbM
bpKiNBdvbUBCKhyjt2zPH45mCgLzgV98rFKMroqEVOwgNASPVLywSqcIhsfBtFzo
PuXSxccG68AzRwC4bdPdACI1e+D+XKFAasWFsWM4r29S7+Q8154B95T881aK7ah7
u5LC1BBIpkFNTatSVEkewcv9w+G3Onlg2eB3fPw7UJqHP+1p9/OZDa0qlone+9KS
vczAKyks29fyKPLZVoe+wvgCjJJndVodHjbDkO0zxlZzO5Nwt0+7d86jez7nzTO9
0DKYxubx//p1U+FQmiCDLOig5Pgjn4kdbQf2uAIt3VGAqyXIEJF8Mc3hk8FRr3Jd
gC9fkrtPMAYVLTOsRqVh5xvbbReej7ykwcoLvOqwZEk264h188uUNU0VGUOCwirO
y4mbfnI7wsU4SLpt3FKnMyKTr7uzTb50iKvZErsRkAWJ8H2KkjTTeXgDiDKqk3ZO
tZiNfBGHEdmn4Iaydvdyn0iT7pPxfFY3u51RZfSu67lQ1Sn/r4N390xFk3V+S5tm
2CiDUbhWOGylgrQh3xCV7/NP5r/mBuGO20KkuG1jTmehu8VgiK1/QuXjVEpnQOm9
2xRAz/YgMZ7wkkX4hfKCHKUe8MbMtBwifN7ETCZokWLiYjPm835s6o4S9ucJi4wk
s+yk8UI1PnOlOAgQ1gbXFY1gqQVvZQ1clufKW57ZRocjjqTsNe2ejOXnH1cBqI4I
Lm7y+WzCOZzuruVQ0zq+0XXjCHdvPAGF1qRcQUsj/+fa8fb5LhoNltDIkSxaZNtj
yFnjGZdGiUdG8TFYH/c97KHEPSiDV2skRer4JTLRt01DElxN2yYRuFw0hwYjAjbt
W0F4/8DOabuICzzAGTnvZSQPAKdhFTITFMeTUNq1X8K6cqLbu4ekNsQs36dxgOpP
DNs5r7V7ZslxG1wS85KtR0NUZktyHVNED/IIoFykw5l2qxzyGShwyP66Km4QZlLW
DGuaJsKa00SrRZ2SBI9AYWzjvAj3ia+RA/sM9ID6WhUxlQ+tsqzXP1BKEkWazSAr
0ZvwlCz1raESkSqwuA63wO3OiSkdmYZ62Wc+6UQsjda2ak6VDw6a9VEo+PHbXNfg
yaMYFKFG+30DVSRp4YU3vO0tyv89E3x1LRtslZc3DmhuxGFONnv/M4qZ7HnqvX20
xIHkpmBHQ+BYbe8nAU5A9sU96UP0GV6Xu2CNFqjYU2U9sN0XfWehNHTzNhCD4wNt
HH8i9KqctzmWjAPEaV/WJhVM3+qD0jK4a37NZQAVgcydlIf5iwL/m2AJxiXPLt5+
BdoaY9oy570ORaOKLGTP2+CNZPnXkZMnTeQNu5BLCciRU2LZvxfUzOnZW5Hutcu6
t1+A8SzYdMloRdYomCFSwlrcljXQcpLzoCk43K3kyhRfOLhYl3NtkG/1xuI3q9qQ
HMJ2URLR2+CP1dtf8VP1dqOg17r891GQU18uA1Wej77VdyJU/cHnnzQDe5IA6DOl
UE3kCyITZ4QcQ8+MpTWgVFNlPUUXji/SVPvueTS8Aja0TLfRwGGHOodj64LWSbrQ
vJhPu8+7h9RjSlfMKGdYjIRy1ULujwX2uuJAQqHuC9OZppy1dmHeZoUpxD97dMMz
ry0Zg4LSMo9CJk/K72pxxyXywNxekqOQdhQErQT5nzbocCXnxJcnN+X93kupq++9
zSOBX2bMwaZSFSWXU0gc52tdrIdgQ1AAtnJnmZ2cLQceMBKYxKN7rbZJY0veziZ9
COjdMTjvH5UxIac6i7jKehMjo3ioaaSKx8n8FN5h5EUtBgY20pe3UPRcuM4C6LYE
rdYogzF/oRg1sFVwlr9HCYRj4BKqjBkgGgdp1lIbnWTrNdTkqTxx+SaEIkSqlSfD
V3QJazWBp52ktm54EdqInN7aOBANb4NPGAK/t8YxxgrF5zdh8DxRWX/+Jc8krcxd
81OyujtjgF4MWbf9VdBX70J5R64Nwm0WPfL+pdEUvHjonrCAkbE7Bg9Wkbjvpdi8
aVBh+29gRgRr3pZVMvC/86ccAiDYvpKBpoSw5f85ML5ewz4gbhFgBnu5NOr+8sHk
Xe6UeLVPhPebcwAdPmrc+rZo+Z6MXPTdULSnHCVTjH/F8dCauU6SfxKrP38NQonI
1nVaBi69tzEh9GtwRK0BFhcQFFIxVnLdxS0i6T+4H59dya6O4U4VngG7y8iaNM6r
8y1q7T0mQgYBzJrHAlAzohu6ZjvDQdQOtSCd53DhhXQ11YHy31cSeQzmf3DvCXBQ
eIvzcezFOKh4+js6ehn8qnFrTp4Fogz9MYnkP472yYfUMVSv2gc5e1llEUP7OX5t
1eOKu9tRdOoc+6iFLNm8fPGEKa6zPQ0NdmClCfft2zUUTX1zkHlboaDlUyASM5B1
kfwFzpOjyQEvZgs6sqPv15/bJDGV6UXtZxCJWoylTl66acKsVEdUh5+eyHXz4qJH
F6Bub2vFE6Uidj5Zn2B95qxJm3LH8e2+CA7LJLpvnlsGt022+IM8bd8m9y4XiEQp
cwTBdXkhMR9vlzhD10kkujvmZSgiOOaCoPrg+mlyF5bVhkN2EOZLypCgUPcVmdDf
CT/kenDFZAnA4RGIRDaggngzLel4H/FEupwCedPOEeFC2/D+yOZs4rHMupfjL58R
kyJ/kz1PUekHkxjFy1dJhxkPeX2kdT7hxdsU5kiWv9KjWHTCSOI10jF4lfUqNhXO
65SEUpvU5CegwIVseBTkERv2slnbSd70slmkJEYOUUoMp1C82L/mMDAuKt+6O0Rz
lNKUqDMjvfnkX/xeLnMn6qiY38fTW2fp2Yey2QRQtff9YHik8QTIMXYlnwMLyOHw
g/xR2StvfmfeQvt5pcDERLxcvmK57aRg28sKSkkqn+K+rv0UfqmBddgnrQHche7Z
8C9MaCbdNrepzY9PUzcI8CA++5DCW+Kp427mckYUv4uVimLcoIk25Zf52rFry5FM
UojOxdJrq0NCS1bm64xWZX2VfWb1K9OkqjT5U51Y36rSS/ef35WhFax7CTJpImQw
kwoxzzB1u9/92E7Uz0ACXKDKDj81eIlel4A+bEYiKyKBSXzzLiPMzTjdn3GPrLMM
b3bK1EI6ShUIOEY7OjYhstGjE17fb7bJjNdnKNoTCY7ZEQp2/2fG7PA7bqTQSbk4
+o94UHyifMJeqxTOF6cafW9MLrVatYlwUCsbkdYI9G5EBs64WeaeRHGsMVBBjRHL
jl2QXOEwPZTQStP4hwTj1hTKTcd0elMmtO1DZ7Y4F18J412HpxkptQD4n0hdIkYW
f/iKOFqPyuKxndasMcASd30J2d5KDvk+7I9fgqGVaVlsEQXakMqxb4m9Q9XlLLa2
KB80WOuqh7h0wO7rtNPDyFxI4asyxGz69vqzl1C+6pLHJQjt9mXWl5JH+wvFzv9J
b8bp9ErU96pvQf9uj1JiX7IdKX9bnyH/ijNlH8bdtuEmSAzWWePgzMKvCyR75gcz
KOZZosxOilJ5TTpZWnpMXVGHDGsbw4ge1yiD5X3lNj79Iovd528GMD3QG0vwyNrB
p41ULyqAD0l4JPsruscpgOHNpq0B5QGS6qPfiWbmut6yXRLfv+Vwwf2EgiE5qoxb
jYA3fnzXJIpCJ8Gwp8XoaXfcLmn7Li8Z5ME+gt2e10IZ+6/g1Rwx81R37cYTUFPx
89n94h0OuuAKKRhTiTRsaHYaCkOToAYec+gNB83T4TX4ii0INcdDCFmLzRMYQhdy
aDhsQ5HzOhuhGOZxuGUi8HVIpBw5HpeW/9h+cVw/o1az1q1yQB0F4wUxOIexGt0w
76a3m0RtiqPToSlIjW72RvbLjs0JG9iA1Njq6tNHPd0lUW4gf/JNymd0D6I/+QY/
i2vw7mWqZArxoVLVzdkZgx84v5g43L6enBizi8fMR+nVfaMcaF2aMQQSmBHc3UGf
+tJZEPP6uz1Wt+Tb2Syb1QHjGjLngNEe5ynkccQbI2fj7VHZHTN5qq8vlo3Cgm/2
f8nY0uDqMeGqHqFlevSrcsQFikFkpr7p8LvXs4LFRaNzh3R+zoe9aTzWBZLSEj4I
HO5F4mIiLn1OziNlF9hzNNN3KPcSzjXEA6uomC0Vr2ht4JphcVjHSKXhCxoToR+E
y22OEWPTu7dof51UMtTZ3f+yaQuqnd7/Pf6ZCVyTTf1o89R1HepDLgJjz2lwsX0j
vhB6pu1wJ5Ttl/8Wsd8EoCYz04gu9MRwI7rY/mL5WuG3ed5jG67/1DIewHIujttm
qhKXPnnScHb2IfIKYf0qedUx3YhbcV0bi3UWIpB7NBK2WY7fUjHPePaPdQS1zhjV
42BMRBUdhB9oIyHiMH+KrGtplFrs4pYAho1q1JWajqTC4nboyWDs8mG6u2FBTgys
+nEUxk/UNvo2BTg929lamvc0KfSCwgdwj1ee7IfmzPDjov/rD8VWAefjSj7gLyZK
sDEq8Z8NuVXkpEar0hy3w9TesqvET3o+ZT0YkHfjJM913yECG/TBoN9Y19P94mN2
yP8Ntqiacvmhx080EKjx8p9NNRlJxlj4pMep7qOynE2KR66v93CDrEtNU+vduN9X
z4MFHjsuZ5H/f1lRhCK12YVUDzK4JyXifPq5sgVMv6iZV8O5G2FqTbgXue5bahoK
Ha2OSAVjpub9/RkVD7xn2IHVr62ifwLdifqkyG9mCihsWWM8bf56qmK12SxhTcaR
nU6bxSlXfUPradAWzTKppAQGo0gqaskPXwqX8dKUF/PikyMzQOoDyh9Nz7f04KZO
9A/8r2TyiEd/M414AoKnfZZSKXv12Wah9Ar3tFWTltnwmXDzT3hkVJjppYWOe2Ry
pn/lY91DQoCvA+hVIujZHigoE470b8+qngq6n6HnUP8mzJCg2NXZ0oIBVD70IZdA
t4xRlS+v49iu7AchGzUDm2vWr3SSg7ekwlEUYYwy43ED/CfNgyvRJiU2XI5J4lga
a+uQJLlRIrvWAMoNBV9XB4xCPgvllqMGfFzVqD0i6nnT3ZS41EV8yvl/Ir6iFwb+
WBO2iam7gWg7SsA+uqUDfpD+VdzNJeQhzI2u02QL5S0Cq+Mvs1j1ERj6GKtQ/HZZ
SsgOsCtJZ64ICvcN8J6/vNAIYOEzc2FhKVTwXOC9QcG+mNZMcOwDjuqUIKPcfMHh
j+6NGIdUSfJjxqNLduU/q8/+LBtYxG/h8QLcl6jf8a/xKzA8C16fNd5eXy61pJDt
4rPU+Ku5fYAV8iABNFq5JXoMoUFwvtJF6HqwGdvny5WNRw1QP9PaC2VRiQPq6PPP
kUbOScRArU5S8UIZgfYMTq89IBwH3vaMvihp8fGU62pngXLLTNIQ0OuDAjjEXE3R
nIfv09RPf+HXiaHx7Cl+s4XD9eBHGmNtN1S+aZcZJi54yD8m1wsax/K+1vAbjkj0
HZIhbZUTV7j8bXzwrv3AQP9OpvUmyLjnYMduVVBiJoXY48qS0pdA2ucfTJLzwSbR
hYbOKAOulFONAnwWA0c+y0MKUuIpJlJKcSe4VWfr0A3j6YNFbPfZ43qRhyguQHM3
cfEi1uzK80cCp1jX1kjIAQxHKqF+yldTFBL3bsDOXjm6EaC1eZCIL3Zwrxmb82RH
kbLnQKnETXAnIyHXhBdR3fcWDX6qIRL3O7sVIO+4h8HKHYSvWp2iM+jhkh1LL8HK
zNHT+xn++AuSB/6i+wrc9dnFnEYYwZiCxIcf8iSVKEYQesyGkfLFnckrchpSAnPs
8DzZ7TAAJcbi2eYhwlSrPlxh3VimhiECJUJTWg0nNDPG7WSTh/6hbZhooLEoFTEP
bp8NxM+e9CWoi4nmje0pU3Wh+ImKvS/gyatYCVsb8QqH7gHlOAGELOWrESPWN+bK
FwtVSyVxo7eyFZqF0yV2Z4hYZ0WmIKG059ZO7LB4hLeyjFUNU4DOwga0wkvrCCCe
wnVYqJ99qhR7+RM0/r1i2iC6hstpEdYafikCtgKZgqSLTDRQUJFX+50Nd//KFPev
mlmSWNLQl+QO0TW5U++w+vi7vPsVTcHOOIzQiT2xYw9ANgrY5pBazSn+ko2fiZUx
tiRJqE6PsQgP4uK2ZyMVTMLLympxTeB+lHn2J68YgbTJSqtwiyzruSrAzEC206lZ
juHU9r1updVdslVeaQvgVmedre2Z4tqydiKHyUVMIkrnevEraIGO1aFiVuDGXzAm
pp9q+d10MUxAeyvd1+YHaMZRaM9vzSrHImh0MBy3YkuRePJ8d1Xdw7Ns2P6lQBX6
rOrdBuni/wiAci01ol9SA6QoPgCA9AjM39EpbOE3FkRruIZV3rmBX8VgSaj5OQR1
oVMZFaBP1PFriiSBYpxxjT1gA5mth3p0cidoLTSFXw7Ol9j7UNSttti/PZHeEFHO
+gNbxLzgQTeREC/bL6NYIMFcJuSB4euTCyNWZpvUrMpLE8ySsnvRp2VZK6mMFAAZ
yn5QFbV+SSWPEvoY3I+4PoX6L+8BFp/5an/blOaauC8EVQWty5HkHgePmeg0Iw2Y
WtFnQW5doAwHF7UQwFm0teX/+Os7E+XiwcBSVKkGo2/M5bwtcGSVam7HYQ4cjpHo
MXCD5V18F7VLni2ZUAnTbl7+VObXPsB0hR4CEhrGWHfBwM3K6zl64LGNnHJDtZgi
ewvFio0H/mJ9fycQkZeWfU4zYdJQzOMnDuPXssN0SmwAUZXkCCEGc5z+S0cW5fmL
NTKIcAZIOZI2xy/513DIgOaI2hyMwNOTVdEW0Vdjj8R9xvRqPSMV52ZkEisOGKT0
2sySt/yUbS3Y6g0nURzJcnk+ae3Nb1bmlJsnACViAnJCRLMz69qepo0oI7PoBn4d
hk6cOS2mhuK6n21Bm7n1Bv8PdPXLTCepQ0bwNbDULLNMHTTWXcpk//tYezNwfl4G
j3BnE01LoDxq0/dgGumCUD8vmM5Vv7f4fD5Zj8lJ2wlC2L0RBnvnNLy/+bhuT3EF
XclDvwQPqeTmgEEXvVdgoLr1nz02ol2nG52nCU53yILG9+FdthyY4mRDSHfGr6Ww
A+s+GU0ugwhVTPYYaZhT4ACfr3/PkkcZ+aH+C6B4vhB4sdo68X8t+Qo1dQkJXiIT
IhTi5USZGQZS4KwBKN56tEav9pNVxk0FZIjZUlcxyIwEx4pvpuq8kyRrF/Ayb4pP
fN4BptQMhAXx31w+sKzFqZAJZKHlQQ4Xz23C5h9zXyz+kx7wZYKiB3vE+V/LUwBT
6cjo+10Y/VSKOwXULBNCvP5N1g0R6dzWRmbWfdCQpfbJ5L2Ic66QxYsEpALD/BZa
h2ejZft9WnCLW6+hLb0E1VAF5cWlrGLN6bGcyl/R52UNGrPLMLtcs4/klkz8AbAc
x6gxM9ABerBVqt3vEyoHP+ATR7Shj6JpLkxF14fVd/KPj5cflXDDmZNLx/k0tJXk
2QlOKZdY8MS/1mwf18DIFvvhtpG/gm5y2/eHuaTRYh4l3pF2GQAxj9p74g5n12zm
C5FZ/4lRxSGv68ZTGDnfeb95fhJwONtytqeK5QAVmXHa78jM5bd4ejUEtZJa9AM5
J3OQAEufH82MAvtwd2vTJv8mc/bzRuqXZ7KlGgKakugbtJCm5fLjMmKw5DuHr5yG
udhK29gzfWwcHLqQOdJlg1YAZfWAzHUAuqht5sPQzlDGKelAVzv+fyKI19e9ry9h
rINGGi2OnGEYNH2egaT2g0Vu9y8s8E3CD/f4UEDecI9RXELXB21sMu7zx5Sousb8
6xI0FnW2ULweNx8FgWNdiuLQ665RNZWik98EiZPduv4BamRioX+FCpPO3gBc6s1h
GNgNO/+t1HAQ44xD2PzPIftcIJfh6AdYfshS3/MEyWgyIHDlvVfFYK2RH4HH9lZu
acvBQLsq0NKgTuwnK3tv7UWqXNNcoaRWEzXpbBgFhxUAHpCAeGxxMB34RyPEfewx
X64nqXK9gzsCyDYpQdgvbM/OJmqEtXH0JJGFiOS6JSkQtHWqr0QnBh/JRtT1He57
pwEShOdvqpf1sZS7VN4iGwEhl7DHD/RUKh3TEMWxSMDnm9L1yzot3SHtBGTYmDj7
PtCgrRMEONlnkaPTBO0fqHPAKRw2lwpreI1yq0TGfS5jn5Dz9l9PeDhcLaTpbuCC
MuP5M9TnrXZ1CcjzuSDsxRpx1jgJ1xTsEMKw0lLzse0OOwiNJ/cAHvkwodDzHbSv
b1Z0oUPsNDSaFS0HhfHghGypZc3vSpoCBe7OPixozfKFSj+BGchNxULHsmfdCE9O
OsXnG0RfdgvQTPEU4pm7YiXXHydkVy9BsTptCPYaB4aZaeQB2ibecXEipG5SaVvx
18bIuFJC46mu7g6/DFVJS+Altty0eN1YSF7dA4e4e7K1gO60wRISTFGG5dFIZeqK
Gv5h5fLvdBlGgjMqTDrU3otD5BqNrv/R2nkrPDGiGj4akWvzJgJxHT61IpKA9iEj
Gt6kyxPZLfYUU3BsLMd/3V+uXsLP0TZWIacqfUCHY3jkx7ShUYKwY8a5ffI+WHCv
NCmuWxM3fYNzByg4U7zDRUFoIY4O1wtWr5YudEr6oAq0nDw6h9/wISb2TolkwPpJ
b7XTCQvNM0RXjmpsDgDP+TQ0xDFT/6ty4WDUONrbEBznUbCrw4Xt/3GSVLusN18X
z+RizZjQnCf7rnMWpS3oyts4Sdp57us+p7l5K3lcy+XR+0cTMj9A/GcpdhDdbAlZ
Eij4VM7OJtbaxu5nlgownCqBxeGGpn/E8eTNsgIm38zf+XJk8FsnCGoiYgO7CP5K
/r0t7yaWv1K0HV1fYC6ay0KKZ4vnSegy/H5TpxgFCVkqmajkaQqHOdY1PO0AKlJ9
sCjXrXyZd6TtWACZom0AJj17N8Z/y30ft9Sj1SPrFJUcFbaf7mqGfrL4kxoc6M1B
znP3C2gS350GekcQ+21EuXwRQYcigaGXtmbgeXlEirBLD3Rc+cNbpIqy/wsdVW4z
paxcJEcSvgwYKoZOEdnTyLZDz23w4sRAKhsGn7skA/ZIDJumao9fPhBqWGcyqKVn
uoTdSoHc5RxSM8Lack+91pN4+6qvipJMPKZlYv61ck+ySS043Yv3ku6cJ9RhSVUM
oXZyTSNGtyx55Q/JYZG6W+YadeSXIrcpMhoc6Zif1tXI7dhPiZrgl1p22HOYxCMC
viXEKfYmwrhCKPpHwIZIzt8ztcDL3u7dEzmiFsht6k9sZfVJi63wiW0FHa6dv2v5
ttcHPWX+Yoz/b5Ie6yxe32/2YIHJtEiv38PeN4vuy+uWtw5pDWTZff9yXxS1a3Y6
/tA5Z/9U8O18t7ElTWjRsiT4KzeJezDnVDPYKXydvRshyat56522CeftaU8JgKPT
Lli6hwELE66Oy9Ehubtv97rjEOttvHu1lPORtX7cCr7NrzO/S5q9+u0W/l0pRlb1
ypxO2xGeJa1YJSu5C/uw1TIogmarejb6+hA+M/I/2InSG/DQOGyGV9m2ILD45h9N
SqPp568HYPMYLSiNBfs55GP+pFYWpk39LNvJ+eWo2elKkMEPUf7nS17RdcosHkTJ
sNxCL6X9K7y4kpUkM4mzkEjSUos6l6E48dxqXTh2Rrt0ocvU+VsEH92HKAmJozq2
ErIH+zy31Pi1QB96oJ98PVVkuJy/MSEC+HKboNoNoVQP81RDHhibUlK9Y/ni+v2Z
RLtjOkAhpBPYGg3Y/0wnmhbLJ4hlUarMGh34WbVmsQJno3BpAWZKVipIvO5RrBMC
by4PdHnbZKbfcIulxwiCNjsE9WZCDDhow+n2t0+GzX9mJ62DPCFYkTE14JyjODhd
x/ZqsGGGlAezfzL5EaNabl/DZNdDPXfluoYEHOjfaepJ+nuXsv7W8E+p/xQWtk/W
ujX3IiJmCqpQm8yZnUajMOq5qPyAtGs6akwGYCLXQfD51TRg505R3p1qiQb/EiKN
oOBmNmWF8FjiWiqTNlDXQ5Jz7f+hOxMnXeegUoMmAj3T1meLtwXdPQUHARrbkqId
CmZNvoFWTDX1RuwmgDXJBuxsFMTCaw0AbSXmgQqswFrnQOYZy6vvmQI1BTvdwXTP
MsNXBwLRd+BSw6EBE+numo1soFAwOXoporULSDdJKK+6iymSihmU1kmaaUb/6eYF
DnhHClKQzHeBoGj5z3dWAYAvmu3JLsGyRv0p64QBi1UrdftkWm+Gyl6B1Ep6/I+S
J/wChtJE7lWNAKKHTKa4vGPx//GGwWyMkin718PGwUdoKN2pQjqbjTXEWr1IVak6
yLUtE7Vgsr8teRi2exsC7p6AitgRjvYNTDxbsSm1jTnED2IsgC6evnUneN2FiviU
asOf16BYmNYJQGP733kEpTdEOAsWN4HR3TPeIO3ziHYW6zCB1IzTBW3ZbDJFj+px
q3SJCu0YcniZGdDDTwtRdIPGK//hNX+Cc8U/ESH4MVexgrxGwjH2emoOG3kABwsT
TjtTK1jG9Jbta3AMo4EnMF9Jofa5V68Q3e+P/OXCu4XuexkeCTsArA/CWRsk534l
zPNf0ZjOa4y8HQAIagUGEGp6NXh0tbEQFblTL5F/KqfRCdw4ReYrNRXfdPZ2A0iF
qB4lnWMdJa8w0GcjJvJC9eOhiRe9CEJ451hkL5c7nc6rxctnTXHVX3aiWAo05UWs
/42+ejfp6KOkUKg+2/3wJwcN00agX4h3ryLGgqpVPx3fZS2CTzDFT+X92mPCVhWV
nZhwhrvpKucDlKWSOXtn0hAR7lBzOWLvCKxaI6W1TrPwm4l4ETR8B5BCf1Juq9IN
59Frer7PHpk7bwiqsl2Q15UwC7btMTF5KcWKdngY5f9nQOMYK2+TFtQOF6jpX1hT
aOWCcxxQ+5gYPsOku7KpGelJjcxGCVQ/S9u31vY6LLP8LrWhOa5PDDWSgL2KY0LD
xnedT3vhWBfSj7hO2e4J+KZzCiO5LllxgSRYTTy/vliqx3nyTQNTOX6bGGIdIfAY
op27nLIcD/ilrYqFo2QZJxCqWGYcthFywgbXdGZVNWYrFlvBwPkX2oDu1QSkP3+W
U21iZ3O+N3oFF07MeV10Sk2G3DOBpfuyKRxiDULsLkYlEKJRsjfC9USsLhoz6Bkg
lI/8rOgNQsxCC0WRw5BWd1gTZ+5vt2o56cGi5+8aZkIJ7naxn7ve8XF4SXnRgmlv
ypX2sncgijrmJyE4jVufBR0uGX6KSL/YiaiQnD94JFiAk7RRum19qbOoaZfw8I/a
J6narkYB4oAIa0mgd+EVXnuSF5VtuOzBJR1fusSQGxdIavrgHknoVkU7QPdFRroC
8b907RaorS9VpOMAp+A0zku+aKfuFQow36dm9eVNaCuHkrozqNRmIDHKxVNbuI28
0e3amE9Rdm5arhL5/Z17Tuhl1ufcNZY5ZYR9AvEpTqu26PL2N0eDN7alJhUVm9ts
xNGLRWGfQq3wcSXJglonDLP/bk51RzrOmF9+c55ABG9BMGzOOueLtenVsltGk1Cm
U4T+CjzAWsf8mSGDGCjtBiPM592Bd/+a0iQj5ZekonT3LKIEDh5687eKJnGR6iuC
yUX0QscQb17VsD7BEUYKsW6Utu5JZMLcqFOjn8Mhh8HbtXlLxniNlShJfPklyb+I
HPFn++xu4gXkYPi4dgoCLKVQhIYlfpFRKQxoSKjXdjYUZWRPfvTrmrxL5R4SPHip
nPzzEQ7l4W31qhxVFp09oQmm5bFdjwC5HgHg0QUyDZafdecWnKlPW+fZG1Sz3tfi
K1YIMRwO0PleKAGWNnN59N5xkUOOqWKAbSrJaXY9Q2Y/9fKlVe+7iJIL1bMXpHN3
G5HgEt0av1334vOpjNaFMps5bmU6FDasZBb0wV0oxkwZdPJ5s/tapwBEdViQB6E1
jhphWOGIvaBkEJeWefUZUa6M+uFRrc+ET0ikNakrOiBq2UOtgAWvWgoKTTSnYNUL
jhZuUKhdwxbCnqtzsV7b1muxoV0EJsNqfWWsihUXD1B4d+X9Mhe7MP+SWF7OxHwc
teDCME1wA1aNRXxad09eU0QaPYiiT2e+EaqRxTB15NbeLjooeXZuQOGGNLyDejw7
RAv7/gDSpFIWcdFE+pcQGq5tls2T5ghO0FnOM2S9MV28N+IDYA2uq/kuBQKk27Lt
Jo2vUDtARy35NsYS69IxKJkAts8JEsyLnpuUVZPNxpuSpd3qrALbLjaYbLgf5MWH
Du6oqjweETw8JIIBNfGqblcPklEaUK3M54H9rNqyX41TKqtFDUxxu/6TUVl+80Te
VhYTHcV2StZmWsxTHKPJ5no/hJ6DvVEXxMTRvY+R35HP0Eeje4OHMknk+SXPWtNK
g7IBFpsY7HqIIo4GWeI/M2acj99RHIH5wK/QnOBdyJZ21kTADKhjyN7rXpYODK4U
xUp0riqGk3SGolubJELOBolBZ5LI3l0HkTLobJC2lrbxeFFsnKWjTtubSexK7ly2
PtDhpBFdMaMTj+mcT7STryXOvMPxaCT0J4GjScz7RHhe0YtBdHtb1yeXqa/PnxvS
k/eHNZI18JJpgbxsKiG9/ujaLNzV9kYnZHSQg/7aRK7CrrFkOuJ94Vr446zJK2GQ
5EuJk0xPfl+ompWn3aBDf4sNYooKG7QrSI3KKZR1ykQkbnPqJyLRTTz1XrVOSNWV
KrR3bkDMM1++Sh8nwOTOtRO3HtvCEbyaPyTfhBBp0mi5cFu13oBGktzPF8HPQKKF
hA7oB7DLQafKmuMxsD3q7TBRf0FpXWdpSSNh9/uqg5B22N8MLYeQiPF2btmS8kUy
P7J3/tzsESj1k96z2/0Ep8uzKEofj52fb7NT6NZFzgHhhkWNVFMo16TQKhR+CYfM
gz4X+1XaUx/dqvrhNq8ILSd84cIPoBGKfzUwEwblGuSpqevyiM9dIR9YSvMVNvjA
F7k0k2FZqTOV6rxniu1URpauS89tHNDdBErU95uPTvUm0OcUxO7lqVbA/bRwbsq+
1ROJ6X9v2JN8DFyT+3jXSr7ZweyT18/XM589G5tPa3m5iNpcpGsWSSU4ft3YPVen
UEv6nomQ1vhCL4rl9XjPOFCGhiqO5oXtu9La0cPHndSkhq+s7Qi2Zq2PJ+pFBky3
3uExq5JwG4UrXRNFF2mBo8TFlqACcpE8aohBqCuQ+ZW1AmAug9dzAQmwnx6UGPKi
ad+QwxDxW5e4X7YUEuYucg9un80kDcq5zkxLyNpOaaVh9+KW7wmA0x8S6mUlxy67
aqcjVV1VAT62CvbTtj8RWTopOgTY9wYDasKfM5hw4bcA2XTVWGQmtYAZRKxMQFFg
dDYtw4byGMA5Tpyu0OUkHTY0u/i7nIyj7JpzA7D4t56J0xfkkFZh3JHPxEiIkzf0
JJPXIyI/RwaZvm5fEONMaDyquHMJguUR7K5lhEHJfZcjakak/M4JcMQZRlh2cnlN
/OVBWh13Z93lpBCGIx2zba9quD/GYDqpMDgMxf7hSPMMGxMlRUZJcRV3oYQeyIZH
xrNQdvdB0GdtwxnGjXsxe2Y/qeUbJYkMNFSJnBgoObANUf3Yx2k/PoJ8G/nZ9t8S
sv1hYE+azauXBSgVchB/ZUAUdGJlX2X769kv9bfCNe7fhZD/Gz48JOjTrbNCDm4X
Y/t03BQ1Nq2ttcDv6m8Shjb0P5ol/sHd31GSo6bJUMDD8x8bimooO9sNS0/C0C5J
kOyfvJjjKLC+YP8r0OU8Pz2yNdm5nXdPZSezqSIzZnQNH5buPkkH6Tps4nJzj5ix
XGCeVk3j+z7N43eLgPiZ7W3sBgYHWgEL6BiApIxsWjSjlP0fr9ty3VWeS0bdqytO
VcB2C+kBy+OfDHCrOWhqHv0FkBh0aVJWhL2w8kiVv0ByfsjoQy8BhlQyZFXWvSYD
TK47CFvqWAAEIerdJJvZVj+dN6q487ftXZktHSt4jGIWuQLsB1y5ZqPayXvIlWRJ
1CNP6bj+5j7Kr6e0JQh8OvEUi47y+K2EzdpkkIQlzUXJ6ngiM1xpCDYm/okCLli0
Hd8SKOJzI4Fznzr4Osl8RUjVCjThtrmT5VEY4XEK4VWNL0rNl4kORUo7xAcERBmS
jF707ODC7jqRkjy9UEsp5nA2svh3Jd6f+rvkDdyMvCn9tF8caAtP3OjnbV53EnS9
yDytDmwgf0NWdlxfGLVGxHr78m6yxSZvJrhJt/mPrOgXppvpv73ddwqCLsjhJ5qS
pm1/vmaNWcIfL6qHyzIaZXbfaA+/YeD0neIWKrBMHfT6ki86V8rTA0Smrwpq4m/p
Edof8tykEFkFCoRaLhdnn/fY+QftJuUWD2X0ro1aWD4RnlyUkxqdbJfF2XdBQiqX
LrRV5/4KScod+rtq+ihifImEvv7Rfa3BdgfxtRHJ9gf8zMKGLZzWrC8wjw4d9kGq
IBiBRdYihVAdsOJAs3AboawrZoa2PGmbH4c9VZyZ6epEy+JdCYQNmADeeyJDz0RC
h6X7KG0uWbwJuQZLa2MwE8Ls9wQ8hZQocPkI3CX+QJ00p+rRgrTXNXadON1wEZzn
0qbrdE3+k3HO9KEA04/j9q/IeAw+BINEeDdBsKaHrVrvQEn32ciOizQuqMBWXc/u
EbmDXc7M4aR5uqtCVjc4s/aTAfitVh77oPz6r+zaTBdLJB9UWxf9uxipAyV8nNIR
JZ3oNx/Q0BX5G88G5wh3rdvRxXWDfoRX10n4nnxxuLL5wjfb0GFDrM3NQSjt9lKK
FK0O+23QRDc5mPHgornK46upzLkw/iwmA0h6PKTpT7OfKydoNyzKrKojYEZs/1ba
NgIUTwDo0frjmd9Bc5gk5ktxyiSyWkN96qu6So+ndJ2k6HqOqcnJe1fC9msckTwV
V77a0wHLuriPnCFbnk740Y+iDemD4pRbgGQfAHMkKbq7N+2YC4hfxxxTD7BbSjol
ST1yZuBacX51hhj+rn1y8L51DwJOxwpaBb/wqJH++lRdRO6uD+IiKw6rc/lE9IzA
BSArbXWPL3G7VFHrPXvIrsB9WpIzIIzCNhnMYZOdknc8JTINjh4eRfmGIGs36TVp
pkomfBPaZIN8H5ObbSSmcNOY7hdEz8OhNmPzUJmR3lYZUrMbUPJWmAmvTSBfPLJf
9b57jnKQmehNSsnbVevjUHAi44+NSHV0bl87Hzc2hgONsTSssHCgDhxbIHfvtvPr
fpo7KXA2zgPBXUkZ8r637yWvwjrgYYz0NyPyr8QlVbJ2DxmjTYzZH8wNP7Q7Cwro
pUCvuHLjm68Osb55LXYP5ah+nYOhIAmqyXF7cnZAx32fGhUFQN5qXQpOz45r11OI
49cvoTRlcFplRO+aQiaWVrPsyuP8Ds5vBqgFWR2kaedtwCtu3DPDpgRmWIbVJkyg
/UklZ/o+0CeldJWn7uC8k+eOZgVB8Aux5QypcOezNWR3V/gxo/qCCSh7P8XVZRtL
vo21zHxTSd7kcLRKGicNQrsefRlGj/AvN7tU5PkQ41UZre4m18CDlfRpwHXySIN9
BqLO5qDrHTOOtLLVgnWcrlVu1PImNiaBGo0XrN3XOiC+/vipQUXkA4zstodw3RTw
3YjJnkA3/udRc8dszEtb5y7NngkZftL5814+6LyJxljUfFXQkxC8Y8L7WXaa5NeY
wc0GCRIKnXtLCGjv60OZGZzQlyx5rjedM9zlVQJwRHwmWfxvNmu3n0xP67Q7jM+/
Axw0oBKrl1/pUkybGDag5uEFKjupqR3jk60eIfSwOGaPXzy6v6qb/rKESbtUuXdi
L+oB/6qLoDC9GAWGyoFuJLYUdDMWMGU65E6nHePOhWo60MkkvmnNV7KhTqGvsA6+
ayRuaxqeTQ0D4bStiK0nPHucNvzNSZGfi2hsf2IHLvCRqPZk5vumVxkQ4z87SdJu
+Orkx+ZNg3qRBXiOd1soTVpq8sNE0JzwPtMyXYD7C3y1w6ohNE/wIbAp9kBP8NAb
Z819P3RznfZWlWDOfnhqVHAf8NfQ/HPSwYYQ4c4EUkNLxj+wmvHR2lte0W862rf7
i2hxGv5t6dq3be+BvwozTT5KDH1P1u336gJhqHGictOS9yGBzuLt0tl+3RsQZkH1
5lDCltLGDsIBjBQoFUb8D7/QcpQl5YckSAX/MjOoWl05FJHyr7MTJ83usrIUobzx
FCKVW++RjXZhj+Tq6e8bVxphL8LVuj2+S07uit+38/YeECejLc5f8Y12WLT6RlgR
mNb5hm8/Rr5mZPL/ULQ2lkbniiBhWoF0qJhgPU9HEoRumWHOKp4hqZ6A5G0ksf3c
YflB81pVpebwXYeEZSXIHp6eO5ZKy4a/Uc055/1xzqspDN8xmcKUykg2IgzO1Jb0
BfeDQQOoqi7fwsijf20lW0AOIfCKzy0BZ0C90fojhjMboIdIJc1tq7qDxc/r5fYe
x1Cq59C1OzV2FGevmkOCAucvplkehThDJZzy1cCM2T/Kcamv/ftoAjNqTcPxTCpA
vtas65wxXGJYucyvOFtY84ms/S4vYYx1xmmbT+LmA4/Y0hPHbRQoUV5fJom9Inqi
AWaKE2oKZQ8JKdv3dSu71FAiIUpbeW9Wc1189yk+hGZf0r2wI5kmQXLv0Bfgvz+M
+FQI6L88hBKSrm9uiDgbszHAKKTXLHJ8cYd+9h9pgeojx3T451CtsEDaXtHkO9I0
WFqbtD6NFMxlbS8Bps9dgffc/RX/CNRm7ZPqq/+9NvS5iSB/YEMmzIGHLl6R4kiH
JtowRWClLu7A7rsWaxIGjKdDBCZ+nyGUaI9QJtoNRUy24qjOIKMZUjOoVL7oXFY2
E08CPWu0nUpSz2xyW/FEN0mhJ2dc8Ts7wSVpnQ0PEzSljypvQOI2ZV6q3NwXhrbZ
DlCk6r/ZLsgUIh3+6AxVaYRPDUL/0IOwIB7XXQfGs5EwKbeNitos6S0SkCctdFL7
e+usm0IdxMp5zb1faMtGC+nVaSMU/9qTKp25Y68Sjxn0mK3kjCIfg2JCzdP8tAtP
frmNhIxYiKqZUmSvWd8Kjg2CEDFoMM9wQZoY5G6m06p/gtntqjQVqB251o9xgnGB
7kUmvW0D+S3f6nLUiUtlcK59wSpRXfiX2ev04OgtpVA67OpfZa274A74NmH7OwkU
i49q9PlyyZRcTC9CHBzceK65k6SzThHrGXW6NZf3UmzZfVbmXplVpg2Wzm3MwVnn
b9qVXQkq6FWbR3NvzF9EHa3UCYU+jEJQrOIWW9k72DvgM69CPgwjWjCl4f4tBL2q
2qRJQFi60gBWGoTUS9z6UHM6QgVapUugk3ZdjagY/MXzwWZVqHnA9qWXMd+hUKqk
KlKFe/Dq4D9SLti8xRvZxTtk5Os6vHvtzekknKOb9sXXU/nnAk/4/ItvH5eYVwNK
Vs8j9mHGREBYEJSGRISvMM3nHT60KCAhKsRiQQ0dVvqUNlmpUi+oflBoe4vYhe0/
iZRhVMXwPVg1iu5Mb+AwPvIBzjq5uEs54d+rpCfRzH0nUH/z4X4cBESTsdYBGw1s
bo0CaeLoSaOVeUUudM6Ni2kU1cOen7zGSD0xq71x5hrkx8ZXxArKggBiVcYbMKSp
W5ERw/4HUyA8XLQdUditRRYjiQQl6w6u1sbJ45NObb6oEAmwBdwgES+DwNmk6FE8
9FO4bhH8tUMlmFKpnKSVLCKtg/8oRYUMjTXvHOklyjRi0kycVuuj2PDid/I4CDGk
aL2n4csr2R/y2EcNyzgKIxNb2q0m+d2wYrp2Dl1AVDDVBi3IbN8QE7bntHLAF0b+
GD7bs+ssSiC5PrwgpyetbABbe1SXLGIb31zXnIW4ngkI37Dbkdfv3mhovMn2VY/2
vrsEpWn2IsYID9SEZ6YSsdOg8rqQlB77veSPWfYdvtOp7mVB5I+ro9arXONjIHia
EMHMBpX0CfzmrJRRtUs1doogXxD/TMLhL6GpnydjqadC/ZxDHAHtsbcazZLaAM5o
0as/fdIcXq6BvM7ceNMVlhhlCyDHhp5ogTZtZJ0XiiysUmFkUbKU+ZWddC9PopBZ
eD12kpopmcGvn5iO76ScXDWMyE1mw9/NNoVOrGwH777TP9JJHgvttN2CTG/3jNeV
1gY/OHXS8um8MHn17grqW/Jju4l1sM9XChW1hCstbjvp8O9s3WN0FyGgel/tJOU4
JYdIst18+PFWYTih/GwmhXTJGHO28ZF3vCBUMk11HmzE0YLfnfg+3BQYfbrfPJ/a
Yrqs97ys6BO6ffJbcfg/TnKHYW/7EWYhd5zhYvD1VwmedpY8QZRAEuuCnswZD0kF
DJkgG6gCI/abGCQmZLgCdJs9ynw4jdvuUsfCcLQdRiwu8Czg8yR8fZW/30CXCQXw
ST89om2wMMUjvG3v9U8It6i4iz+NTdoFMvfDancwXgOUBuq/5cpY3AWHnJTNmShI
Lx63y5BKQ6zRBqYqdkhqDRSv1uKPWIiwV0vUl8cE96CnAxXO+x+tj5kIpP3E/I7W
9bWPgNTPW/5yc0gsTcKdCD4pss5wzzcADCd7mwdvD7izSw+i+VmbufOC489OIKfR
LHoLbEPLLQ0xxZZ361R6nLWzxER+mp5f7id2/kcmE1NqHD4ZOzjpmAjOPjUBY4LI
p3a9aiBi6oHcp1VdxplT1biWKUjxzObDVSEI152naqExSoRjuB4zwp7Ug3ViCkir
mn/PWHrGbLgx8nand3nQ1cN31BV9ZoOS1Sw8mh7j4i4l3bhL9L22h8QRnvfYZ9Ry
499BmxXRXBzVUcoSfr2tdXSKM4XzO9oLip/U2f6RL1ofTsMYUWnxxS9s6o+rjAmB
Zc/SIrCjWwJmpH4fl7rVCqQHEZTAEFijZqcx6QLZTKacbObTBsDO0Rb3nUdz250q
652yf/1XpxGhugnfimA1ncMoBiIWyGRSGbqXoymaPf30DAEfIh0TzR8kP3eoWv6T
YjksQzxTuBuh3Q7CJXvoCl6BLF1c3sdXxN/IT9i8lPTHlnYisUuQLYcgFxtnt0YO
53dLkmCxCAQwMSA238i696ODnlfVR5i9+3LlHPxEF6K5SuNW5spjsBsO4dluIlLa
wlsYXDCQUjGiPFMRg63zqBFvJF52JQ5QEGOEpc+o3PCHSGyMXzrq8eH+Y9AIM443
G/hANQax0LGva573q3XCLn3GiZUqVKA4wwEBq7rUfbLbGXMvceQvxXV+YLZv+Sin
HDuLzOxH2TnPpRa/RimbAmX6U0xqxCqKtYY/KnEIA1NdCUzfWpIm148k+5D7/sp9
cBLQoQVQv2qxfanFgj/CSFAsrXrvnHKj5cxscX2awUeZtu4ZRzeKaZVKIQIuNGSA
F5H6JUXLt9I30MTfSOgx/DEn1QTREa1ta4alaovt26v8HWuuh6q0T9V71EPjyvbm
25hDspJT1BFVJHe4pWNoKul3BmEOcQZR7aWNC/dmG4kO0dnBgdsUGb6JXu7FUzH/
PyC58gDyWxoxkD++sP87CCfEFr569J8X6o6vIrwkPtB1nO+mgdg8pD8RPLGVFTOl
QgJOeB7haLUcgxv1vxdujdb8Z064sP0qNj/3sH33Rv+0DhY0mTUdw9LL4JYnWnR/
B6uTU7sOqMO0eCQzHqdpE1nAFoW4PhXpXRMif6Oou2V1ms0FgTTP37BbVtb4oOuU
+KfrXAA3SAtPvrIxq1wZpAXzJ1mfO12Q9An3ywIzwLtJ3G0i32ASyrRbDnBf8oiw
A738eCcO9wDzas2gFIls9S5H3D/1/zOcyHhP+qbkjSDMrpcxL0nFfImje4QBIRZU
SEsPbfy4YWuDpuJXJiX5/tqNLnbLTFHLWi9JBcW/I4XJi5qoC0PtAdedDFjnBJqE
Un9sP+Xh6KXWBu6bq16EkPKc+K2bvrWSb6MJy8rdrdP4nYX0PRfJgDfqHQfGvFof
mvbzZifDrgvDQowl34MR5Z/IHWBTQy0SWN+pixMgtpcL1pvKeTZRa2pyB+BG+w8G
N010kjDrRsQlAXctxdJZGt7bKyT8+zOw2YzeklcwphqRwHROZHkEqEUyfYCL/PaF
KXwaffRpfUkoA0fWutgbWCE75MhJHlCdsieeSxkuakqnLgyHjMCUP6/JlS87ygv6
PuJHB4idsqDk7XaP1iMAFc5QceOjpqvd2ASgEdRIs33HAW37Wd8/ij6Rj8vV/8zW
i2bi75JycQXulZBEudT9dVrFPoyKmQSKKiyrTKZO6oci7bfUTVf16k4q+aFT19sb
/RZYg5uU810sFqLJNRfo6Gb2nNrgIvlVed6HvFvPruXB8cHzylM36bQYuWV9i8Cx
OFcgb3IroEzP5YGkYxn3MGBW5DO24T6289S9wInOjEm03RKJeAuQSKfoBi9npoQg
TAWk6v8hqMX/SqmOSfbOiJRK4pUnoN7MR5nLr1vj24XyauMOPekDIb2b0e2ANEt1
2gqRETS30kx+G4t/fVH/DcGQK5BUpzZO4k7MabSz1zhoODvvMotFJPX55e56z/4k
qSkvwIF0S34iZXx62X5ZIprNzZDg3FxO9s2BHzANODi9vtYNY1TsoZAwqi3kCRna
VaEjGjubHifajbWWimkBj6GoP5U3Ez+955/qbVj38ujPuyIWcxeCoZb37uqdTtxJ
+Alvn1BBomp1nxp5sxsuvX7a3y+rx7Irf8VmPPQ99lmTcP0ars0+iaERFFwscYpA
491cD2K5NPzVgIsSNtcIcNT5KTk1qM2/digDM/wrWLH7u5QUSkyGwgnSEo9AWzhs
YOcfRM2n1DWMhrAIxHH9HNrV+zxKd/s4Qz6GGswYGGMKiqjnu72vmIo48G/psadv
9aiobGRMubKxhXeU9tk+StBUD689+NKctzsa/VUfYoqnTRa+r9MhB6j/oZuwxGGR
DwTQksphsCLWJSA84oJJdB5qkYMptA9OgTKhqCYdNvA5kjGbiuvcZF0vGquBGO7C
Klm65aT8940T28wjXf5VTKvXJE4RfQVwJReJL5F9G4DAZPN0R0uHVo2/ILXdSVGA
Dbm51bNvL2L+MI45EEGbB0+blF0ERIDGOt8l9Q6NQa6C1mizUM65sSMbHpNFq3oe
dvv2oBPC18pqW/ccA/nX3A2NiTViAuhI27TQGP81X/LVvWonV9GEjhm7ZP/3r8ak
IKsFbXaBai7htc2j5MEYmc+27nX8wplDQ/1gpiJYWAvyPy0WTTupN2yxgZWO/Xvk
tLnCZDJKtcXQP2ZxcDT1ely3t0Het5bCjZtALfJcDFeJzU910VPMNe0X1iwq8v0e
SSIxtKdNElLdLo5qvLVhIWRCTHXpsdwSV8vVK6R5wqF+zu6p3z+WC1A7mxdcGbgk
bkFSH+IWdvfAEoq8V3+vmTfCtSJH3F3AZmu7pkodxBZaGSKlLQcVb4rbg3CWy0f5
L//kUg6vZu7N3BwBKUj/y6FnhiznlVqjkKkOAkUhn18qzgbJgfG8nH8f1OtGRKE7
ZPgaiRb0NFUZePc8hZV9r2dqTsdpKSsayZSDFjPMl6MNeG3gSTVgizauYo0A2vTt
+gPscegrMnAZwLe2oh1cmoNKiV0VdlYeEVy6Ed4wc6wsHEdouWfyAZcF3AkON6/U
xm1in+ke1t64/M8R95XtlB6ZlZsoKZzCl5rw9oOtECJfZuRRwdppxTXg/+ICd03w
dxXIWmkHtU7S2i+1YJInMx9R7hYy/IHntupRVJU3fa25sqz1aEqHG3Yr6KDhgUyl
q9to3WQP98yr53UY/abYCCallDr4n9IFHZlQ4rE3ZQQcwRpyfQfrJ+JkUCRvyQmT
UaFHLz0Dq7UfbsvWLJYeJW1I4sf4vsNTuQttggGn8/1tYSXg6/+oNr+mJ38hPOos
NpZd48/kJKOOjd2fF1OxBHRxl0aPau5DttQIb3wnw0lle/mJ3vQPTcyhq3rE7s/5
WHcvA66v768lxfP3OGYKgbuofkaqaJgH8GHBg/hEnfBQHLt2EcGqgekB3zTk3P9u
Gf6+08KW4JVY7NSYVtf+7TEPyXJEF1nkzaYiSchEBgrqp3sNtf1V4NxDVpGlSVFe
g9pXPBQIWWwA/uP5905JE0xy7FY78IGJTcQ3stOX1wGg586wGuPFWkEeBhvnpUco
dJ1n4nFwaSrKlAlBGaRjEVYkkkmtliXnP1bKQQjdMacItdL7AwJYzv94Ks3L9I/A
rj3OZS0Ht/2R598Vvet/lPRijTf9VaV+Lxs730OcmFrhMVN5Ztvw/7uAGTsRD66R
70TpsuczW06vIdxj/yoJNz2GLVBqGSSQzrJSya7IgC0eFblKjTqPJUETYSjvhitY
PMp1cdHhxh+HbCCkmLIdtgktN+obSOi39qMvTv4tNPjh/+id2VWjhRjFeJcRkEPb
7XikJfpk2gxIzf2VhAx/lJA3uCLhH3tjBaRHa2jjVzqOLB8axWkfVauMmjuudsrO
Rnn1CdR9zlgCxNKb1ZRarHoQuDuUr9rfitfuI9yqpL4+5rdIChTJBx3ghbM6j4xi
KekdZUMZnCjJrN1h56NIJcDattJdRZ6oo6z8HAqwzSEkj1+YvOKV35V3XnZXhamX
PkLsII9J8E1WX8gAmGcha0HoA1fR+l2T7vqJ6RiAoT19dxYK3b9WZ/0hwzCD7M3I
o/ENwbu7iGxqosLKE408phPFMLcwMbfMa3vNvsZod8y82y2pp4q94W51cdAwYw90
YyyG7qGrnDKhjARBknqn3hPlwTdyPPEK0Ha0NHxCDMiGP6Fw7ENjKDzEQeIull2v
DCXSwoXMTEwhUSy7OjAtHfwAYW4nP68OqprfZmGymRPkDAEWRr0NMMjN2Sacdye5
mBTR1XEOzZPIDt7L+XBY1Zrk5ulYxN/5jOtwjIDDLVqiq1H1rz9c/Ii5RJ+2Zh4i
JavPhPCxTxbQs0a20GgFM6RLuCNEIRkMxLtkQpLWC1ghq1pwZfMAgmdR1pi36oRi
ekV8yV9mUFLm757GEsgy2JVbwQHTRlucptabxTfKLEPqucMLEhGBBozMaafKQN1D
1GYVP11/yV+78sXojhUiUQJGwwkACRQoUoZHYuuv/uXMeHyEwfB/5TFr5GKQoIu2
CplWQeXbBK6NqgV/ibaUkiMxJ9RkCHbSn8f3WN5Kn3otfdJ6vJegjHMWJOoDwKdt
R431CTlAQDyJyIefrVw5MaJzSV+32EB8HLo7iH0OfDZ0LcKDwCSm0HsGRVV4laa4
3hARDdHDn+QmKLlEmRQLsS671l29h1dV+5aAHlMMMi25FwF8+0vu0qrtj87GBSkZ
mqG8LY46lHfHOcxADsAVM3lVH9M/cAc8XkFF6dxk6gWHJGDKY3QRCfeSQ9juRrmi
i26QgSNXkVKrhsEy5hjun8b9w2cBzU1Ka4k5Z3aS6mdANjh0OHcCZR2zEqpXLVRl
HGU2HcuxO5YYB7fYHTDUs5rKwvVDbOhmXoRRTflDNmWTL+VL2fX05RDHrsIE/VAW
o/kZ0aY9LDV3D9l81rrjA+VezVNtiBp58SfyL6gyv3MwhRwTa8ymkFJIrtDjJcmX
2bXkcvjt7zLPxBEkm92eDLNvRlQO+5Z98sMtQof3bbU/+1UZZ3sOEQa5afNHm5Wn
bO/MnL2z92u/ERHhr+DHJ/N1rfPOOUNMZccZK1V8kycTB6vlbAkHYfL5g1VlRdq4
WLWg2jKBMUwmT5oQ3GoG+ULqUwz3M5KnOeEZeKDLlhJNCY4bkiw2AbgUs3sBNYpl
2+9zfC/F3vFemVvmmt9XzZ4AKuBUnYD6j8IPeXxdFQOVE3OWjz3kOF00/XvAnXnd
OrGl+IAde/o33C0JYhRbE6lEZc0H8AZmShfbCertjH2QUyuSzPUP8M1dqMO94Zcw
If2JXf23wV48Fkf+mtoxN9ZreioOpLWUTAAYGhHO8cm79GnZciZPIAM0nrVrn4cC
kv+YBiOQ98im/N3UkOtrFS9KH/77ZzGt0XakKSFJe+8Q4bptPbf+wKXzeXeDN9lO
GAmX1I0D0gFWcIq669VfYViwlSzzHbeJre5VOdJZ3WM8VCkId+9AAvBfstzMx6W6
1ONJHDoyXzlgdUMpRNMVuVDPFgNjc/1SbeHEMKIWnmow5uuNRmAJEh+Q8RPra/A9
JS3oWEMzXcWf5zAGQPFofQbkhC9XcMgFrrdXa1EjRnkEJlDMIUqD5mpIXHNb6HY2
In0kwzLfgp99XCzLF5A3So2ogxluA0ZhLYf5T+JNbSgt/pWUB9WLqU3CIcvPgcpJ
JjdRmpQY1iYfr+7rwg6CnIYjfRadDIvD9umb0E/+SPfsLA88AteabXfT78bDa4DO
zBGct9pueRA+KDlFaQL+Gw+0n0+Sshl5UmWXWE0Cf6SHv1Mg6AsrBYnfMBhhiMtq
DtOzmhqaHChvt5ZMY3k+XU07LCjaMo10SXv3m5y/PK6OsUSaUPU4vREX14s/aPA5
8lkP2//CzQ6MtSZN4VZFU6qgybW46xk99Txz5HBRST267W42mSqvJu+BpE6u3bGV
SikZGC2aGWehEFfJYliuvEiJaTnyAnUIQd9wfUAKLVRkCy9v9BHtlugdFiyvSXW9
+H9cdQ9zS++Ke4Y8JZkM0/aVCgokWzzhmH3RN2nWi/DspBKnmSlgOcMdgfrrI42z
r5bkrYKdbieGPna0AyBpeHFFyyrIwKmUhANoe0GxpA5X2hhyZEX5OwY7JiV09Swe
SNQfyrv/auhhgH880I5fVoc5t0pGuz178fypBEaQelkCA6ylwm0fCpJep5Bi47yn
2qIIsirAepr0RggWo0O+QpYw5rZs22Fd+gdByLXNEJSyX1Kf2jErtFr1aPX9WWym
ulz0NRN3bCt9Wg2YwHpalLnabgoFs0uWMJV6RjfLzZrO1WfUbGKOAHMQeYBDYtH7
dgBC1gaWv6QErPh4ygXQTisMiB3U6k9z4FlXtwqvR/Qo9q1tOawcPlQlNsvi9l+3
6urIJ6TrcSQJOOD3l4gRUSCcoO+8NtRG+kPd97FX568DVGv1qx4XBV7iwCmMpbtx
KPy5a73NC5+br1MOh9JY74AJR/A5DJjJ6QwVwFgPVgd0X9OB/4f41MdoKv2uRVLt
Dy3L6SOEmhIfZurMFbvX816VfJmB5cWBzBM/Sp84EJrxn71GQO1x9NRWrxiJLst0
BkDKvYxHVSTyYH4++TfkoXwg32ohgZk043yMnEmqJR4DF071rCiwIpcAjyVrU9mx
Y3l3BFgDuzhCnwi4bbmdevAqQdL0GdzRAFSP59dbTbXOvG6cixkg55+glMM00gn3
su3k1GQX5H6jOMxzNhPtm5GHu3TIA2xJ25qs9Ujl6zJIY2ouqo01IJJrQPr1kE2T
4JiCYp+PE9LCdGCH1uRStlmRcBTtE7prWE442pEcQpnyqkJRKsyf1TT2zL9pC8cS
HBQsa9/1mwzJZuU046X4S5g3n/RRtvsV5AAuXrp2QVNkLee7sbR1kO+8vmZhzFO5
ponyFpPF7gdg8jMLqOtkHKWX2WEAvtR7U7boGrXFzxD7wLJR98a5N8mhzLTGUnka
PnnySufldG7criABsFbIqt6a5elRMkYtGUgqst0uymPUM61kZz0Rzgin3c+9t2oQ
xFcF+tdZ7Euk08BnYvag+CBL07lvWCSy65VLOXGrSDY3vpb92c1stxfyARTL3Req
A232x8O/YK8CAIHfFoHRkuFU/YJQhhJpW1JG72pesg+QGzvfECuruxvXnDPcQ3OA
Bxo+KNuNckAeQytt95mIcQgDZy9GhgmxRv7y7NHa2K5dzNTFkDG+KPWHkzQmFWCF
HS9myBWkKfS9OQLr6f1xRyju/0Qe1SQAIWy7dNFjRAnfVggPOQ0JnBJs5+KFTxfq
ZvJV/dL9PDcnAegctUfNpyTMhsdmiGBWJOEu6wxRqPuj2RL1Hx2RzYHVrclWg8wk
UlfcVV+Rbfn2ZRBq1DziY+Xm8d5/OVQoMvprqwtchunLT47KVydSQL34lbt/iqSF
Oz+scErRbd4aLXMWCH3iCdQ7vpwixXLuE1SXgE7l2S/gUhcCo/VSFzAaqCxDX/+s
Iq+eV9zy5o9k6mQhpUDqRd9SBWCmejmArCtTgzdWIqWB7APbNGNmNBK72YJd5uP0
rPiW2zReZnKPnemeGYZk1iZh0MPBUE3+9WJtO8L1zS9liRLLlVeMVtjgUqdymSJW
9EBOyZaVeJNXvwe6El0N8C+zFwRL0K5YsHALw7aNvHw+12HXNrzsL5Cl0nNXUC4q
gnyDMXUWaQVwCz5/DKaPt3ZSvxOfIaYVB9DSXmnFN6MHERA64NvngGL/iw6BF07/
x6TPQaNx+rhjV7bQ1zifD3iXjQrpX60fBqaDx04OpFqrDtN75DRIlmmW8OIA0Jyz
bCiOmOxOcSQFeEpUbAICZHDezUrBDkbldvMjCK8XNSKgjnMgeB4AFN/rb0+g/W63
J42d2Y5ibBFp4owzro9FQSBkHVNr78IZc5p1kRB4XVWJ0RPr/PcihZAUqiLcN6Yw
S8GtAZVdKZbwLlfEWxVMb5yZa/oPx7//x2ywZ2/fMIB3rG7b7nnoXXRpNHfNaFkl
URYqNS5kfaw4/vAtMJd4BwSxcFOG+T1nO1w5OWYu0xCoheC+YEQ6o9La1NCJAn5O
xqjaCAGUu+2CAPw+NegL+6Fd7mDL4ZXMKKORPWdmvAtxtTA5J2msvYVg9iJU5PvX
bUHiR+GXjIIOGtJgZ0Jkwwcea6+bRHmdqnqfcv8URpOj055l6mX9ktZGze6eJS1G
dKhfU6uKHfW4YfEMi3cBhE0ChHX+nfnEIgN/Z8SVw5PCp1ve80IXbt06gCpzUcXy
pukpJJw9WV9jY73aL1FZW36nK1+Wa5MbPzIeJ4yBRTfOMQdQC/OWAl2KERvZEzSb
hqliHkkOGVKihYc7OBedArwB7q6Z7fH4eaDQO/YfpDROJswk6p/UsxX57iGZwz55
Os8XKikdIyU2OTAIvni7sarMIo6/XICjmV3pKfu7vF+WF8CYdP7S3d+to2MZI6WP
ndB8bREKUGvLymROI3G/QBveoxHSwKEirfU0HSxBQ/pyMKKcMZ65ADCI7kExJ4Bz
Va8es3b2Kb8+XbtQb+KBIQX4xJxnJCqe5R/2NNa6FrwQPE9tpeXiomVuezTNAGLu
hEyJjRCovVG1DebfYv7POd1jzrKIyGV4tYY5P+a8bti2O1BRo0dJph2jFMD2S2os
NNwfasZQhmUpmUnS38oxim3bpbDXQD1HS92SRmQle/GE/XMSKXyPB36NO1NsSRRh
XU2ikeEcO+VFjh21fAoBXE+pwhb5MNx4TrXVBE604KCESDqPH5zXlEXjiGDMUEOG
7WKsBR16YP6tM4K7dz9hGHLa/GveYrx6v36NF1UMDWEwP3vO9Y8gUb/+xjq8yoiN
9TW5cd1LBglWd2Xf5c+Yvt0UJ/pSMGpoZSlUkiWr5ApETzuo3lf9qLZ6dm39LP5g
WuwQGgBDr7Tq/cfWxxS4IXb2pDCuCH7mCx/dEfuhHSgUr2zSI8sGt1KyspWrCUWw
svr0bQxPszcSJaH2vwN7/5jNgbPQck8YFlBlgG5Y2ugDl9CoMe9x+ilGiHH9Pw8w
oOQz9vBhLwj/3qKWrIiOG3bWBrj0LuyYpXBaXBMB5RVmPsX9a40+wp17O4ak/KME
6esJbJWDYa/JssLol8f2CavUkbdxNK6z+t5JiHkft6nEhNVkK/280YAmRxK5foKE
Pb0N1Tx187lwOf/uzzgOaUQRvzTufyCvhmpWau77S2THdHJJRePYOGSTMyp8G1He
NcTLPclu5ZnUpgEXZ+MHPYVQL3lpb3VyCarDPahAZGl80n3LttiI2jtPDF6zKeGp
ThUW/Rf++6E8Mdd0ZbY3txO/7V3h6jr1VkTZZIOIL+sW97AaX0HkvvlnRFzBYPbs
KU9KpTXIDL9O2XP6OfMlE1e3JSjMYkPz6wwAG28IWy6FB6c6FcGAdm9I4PZb/75F
GTUw0u8fHMuJ5QKNK8NRbNqJIAAAwiecUEs5LtDlbiLw98Wgpp/zLef6YHXKxwbD
K+ZIW6vpafkMqAWDaF0EMG3kMpGih9EsUWOaCqEhooWkelpz87NDhanSLeprKbA7
kSFcUp7UAdrIhyplkMxq/9h7poE/3+gJ9ZDQf5y7z1OjoF0284aunrVqQVQTo+8J
pP8bvk4IBKI4lp+QdNaVxlFtzxovo1CI6yDZ4IENx4Ba59ZNFgOiCU9ARkspgrkR
V+ldTtp6YJsTouHeYjM/CLeC5vRZmWzu1FKpQK0d8CH+xS8JllCt9sX1WLMZRtpq
A9IwzqDrXzIbXMFrWMOv3vGI2hdMY8v7pw++9dcc2qnzoGSnT16hfxE5lyTMjsnq
fGniHn9vZLqn+TQfLxyNhzmkcbPHKkZAMmKEYHyuiEkz86ypF5KvN/Pr1H306mBK
NvLID7dxLlUKdJhj62dN5K4D94BT2DahRm6VCRipInW73xYSTCI8hlVc+BBGt5yj
9/kVkY2Mbe1KuEDvfd1plHskB78KFONReckmSiShSZfMoyDFMO+W8BVsfMJNhtLc
cTeZsO1GfYd0A4JRcosbvRK29qxE5hSFzCDr3cHsMWuIYqJ+py5lLYy+uxq/MQqW
Iu1fb8nVa2cWsRsZZal0mD7AkdB3WzsytrtkoU7aTwKOIEKbnpQo8+LP2YNnF9Yv
IUO2WYy6tCtK/WqhhNZp6E8UUGkWGpy3SEc0oJgxKm7z2jLLiHTZeuCtB6iGfW7a
+ZcpehWuwVN1gFJQdDW/p967MPnt0Ilzpw+ceA4S2h04uD3GCv5OKcJEDBhTxroj
lfsbs7d6xBiQqO15oBhoXeN+Fftidzl6PO+Rj/oBdHmT6ldx18c64oMHTVILJTY3
PPBig9S+FupoONGEFbyzJ2h2r0qLQ+MWgiTOO0k2SMmexGl7SFoowwX/iHRKC3nM
dVvDsOkofHgL7d7y7zPBkf/sM3ozYov7QaAHoiHNPV3FkXoITXT+IZqiZvICQHW6
CZJUeNFEeLj2sWKzSFCzIPrvKyRVR9rVYRinZNgVXuELJvkAlhi1oGxi3HmHRyRu
j11ktsRl/iKRXtpR41kI+gpZFBTLCukvtXtEaLJDPFIFTr+cA5uSNMYbEnIShuG2
XtHGSwkRy8tCKtnTYK4Eg/yuf9bdwefqUPmn6XrRHd44GJrx6pohrmIA25+XxFYG
AxHpg7G4OHJUWX1uEUvsWwd3+hRMlNbB/PGC44NGSnKI4Y2lUk65Q+JTv1gfPuWT
6EPQ2EFbqzeARJ+hQrGw4U/ZXmDe1x6+9FcqxixIUoYPG7hkM9LdZu5hUeLscPcn
5HZvbfyIXu0BKHsVz0cVaOAIhs0077/NldYkrIHNR63j1Hb5Hm5sffMd1EZK/m/J
RIq8LzG2hAuqqbuXrBi0GWYTPd85eoeEIDK/G+iyNyrwfKuLevKdyQkxoRwQCGMg
MTxp261BvVY3aIf3Rd+4Xj6QERHDW7ohHM1JZllAWyeLnb448riyiyO7Xz8kHWuR
CK1+OgBAar8zNof5OVvU6zVgTPtD+maP5Edrhb1mImSfYcWV7d2icJGazsfEw9KS
lmoXhPLyrWUGFAxY46R0x4t+cET0d9pBka50filgJ1PhJngCec+TY3NQaI3TmN9w
6myUdlEb8LvDpV4vZlo61LfDliKh436BJ2X2d44rZB9KXh7kuXCNTR9bL7cILcqI
5HrfdTQylI8LJ38SZ8WW8cqQn00jEXkmRNi7biEcnfzADJmAGH55tIHpEzYZkkf1
jFoZfuDqjPmKCdaxvQn7ca9D3fsXVNxaySx8NdhNW1zbSgkjRY4J3LCA3q/yQIvJ
LUmq6p6tl8+GXyWbJaAJWcBArbX8U8bzEiSY+wmySwe3Vv/fbZFt+CfzBhaEK7Dy
2NFbYGNNE45RHtEPKs3sjmP5Omt64HM4MnRGSMlYfG4SC+fwY7ajIF7zpXsBtpOM
dgyAu7lbhvge2WEqv0cOO72AljYGW4SvdeSfZpZZegt6rmdSW7zdEyxyjHE1yJip
ekn8K9TlP8WzbLlW+Z1WetMsyLt6PMXiBqRdyx+1JvfgES1uoHu1INtmfunuAB69
zhKxORfXbGUrBjqilsifIRnphMaXKJP3+M+qs8LVGm1fRDcZXt1Q+tjcgGJ1NdoW
vtGEYrJAIVtLHH7fZoVy63eLw0niXgUcQnuXuzG5yePdkYfIzVHYg0v07obngsuD
UtmMh8ykVSkLy/P/2v6RZc0dSRUHswBH9WC5qQFrszD43yW1MWYbsRVOy4cqdM+X
kVIEf+3ywl0big5auKsasW5C/1G/RcjEsKP4WChAtKeTyqmTt8abnWdve/NE830q
L8GPEKwOLYvvAp5e4eLzlN2oZ+1zPqDR8MqaWmavwEVncXPpO784tmmWY2JNdZ/q
d7SjB3IQbwIUmLc3Wm6VkkARjOP6Q0vHEX2X2OYhum4ukjiZjGe5r02VW6unj/fu
wUBzZAXQcr4xYwhqX45YnAaODdA2o8sas+xb5lFY3ZR7rXEgay1tn252cYI8Ruch
LEhkZ1+74tfGBM5PPqARqgyN8xeOZdA0Y5+NfhMaJeOoN6ciJGvUFSwho8FTl637
GiGUxjU0nCxU+t3IBgHSOiVOVrIaY4I+FqI6CDRzJSLBMvbiwWroB/a6n82hDtBM
o3wWiVGnx80Opv7bk08+UpHslDZGJGX3CRf5B/kuWOZboFDy615dJ1cNJw91T/e1
CCZQ+br6ZmaJ5Gaz8U3sy2OGdwllqlqGo/i2SHAGP4m9vZBn6eaOmhPbZPL8Vsq+
954hw+/vT6yIf3KoiEvPRxu1EDdtHDfMH49JnXOECeHGFwqo6+5mgJVKvZ7nO/ga
klgRHgld7BirITvmoFEGvi4sGztWf/IFjAAdNJ/GMmvXV54qa3sxXkQN2MpMV9k5
xX5CLilvfvauufzo9JMt/cgONrEFe71ZlJKah7rNV58Dx4BMduDfDMIYPBoF0hsJ
3UcOhIhrHgL//icxhGt1RM6cTjzr9ymAC2nh9ZklZoltLaRZbWccf3vwARFmPlV2
pz9w9P/UiRWjQzUcjCzMh34shFOe6iMVV/N/m2Pqj0nR+ILINkL78IkOj1bX75eG
EaERHKfKJdexH4o/6ROdMd66hUKNe043YZI2OCU+OXUzhSyFYVcJ/aBSq7c5enKL
rGauePZNx1P4nc2fVdlAG4ZGvT3EzFYuK4UU9bxHccaAwE3zwVNg9lpB2IBT+Avk
gMEgawiy8vPMKAYIoXnWMsQeu147LHHko6SaH6fzKpdGgLY5dV8HVJf+C+DEt03t
n1r1GDRWZwWzOdeQB371MWbnm01XCmDvn1PyvS797Y/uJjghnDRA4m4Ib+EiXAgi
y0qjdpL1pG+G8Dsj7iqNRVAWi13t0yguKya8nUpXn3QpNGhQt8kbGhFUCVi9T1ey
bOSBwjY2Nd+srOOXspMIoAzX3hx6nPcl9CYm97lu6DTkUYZdtKbYIemFpnY3XJfr
zMmkJxbRjeQ1LQeCcI1dKdD0nVulFAyUlPQU6bW4yaqsRjPB+SL5jMPi/16paPX9
wo9xX/Ol80Jhk8wQ1cSkZ2wUQPQZkL0cvX6zbFlRm/SXHAycB1gNqfKBualaQBly
o9q6WZKQtpZI3S6bUVO3ZBPpWHSVYpRr4351AquJNbPDskWKRIjBOp1b+a548tfz
ondVOKTERzyl1xygIzBnpiMsJUvAQDBM++gsCKHobuaS0DscXyBhIkz88hChpNEh
pSGsS/IpVd5xURK8dYE++MXXoyByDbUcjBsSVJzRtPYx3+Z64TLOWOtY7fXyHY+O
e1ANfIpnhVYnEntRmB3i0iUVtR8gW87ISPnAFxZRAPZKMt+T9ts9i9admzQchv7Q
lzn8hyt1v0hiNdRTUVj0TfVERrFX7cadS3ltVrqO6LJ35M3vlew+XDJBcot3n63T
13q3XOssLRgICIr0334YfXhH/KQ//wlaIVHwxOcz5ybl4xYfTDVLPhszsMmofgAd
zV4Z1GN8wzVbsj8a9atrP2yIS3jesNN6tGUBUZtfI///fofeftBIoLTt+2zecNk0
BRsoUjtuQc3qxOKwY6Hd9P9ZemFLaSXZLSc6LU3+x60xGPIcnosxx4dC24ERWAe8
X4P4s2vAe+fHxybUI+o8vyWm024BD8nl8U1J6ICzn8dsRIHoS9zShHVnf7kCiMMM
eSQ2OHqfo34jIMiJVAoZfcw5TfWaOxtQiK/utcR4mYzR0UfhSBpquFVkff7LNzhA
3+N+EZ0T0MoQPiXa9mxFWzaaIvh2w3ASp1S33BbMxpNqw3v/Jj2zvrr+/55cl4Ki
+tpM9nGZODeY6VitiZ/WU1QJAEwNr+JBBLFl2q/TZxKE7ruDVF4V99CqFsBpIN6v
ZTXyvr4CcqfF7HSF6q+iGg+ang8WlZXcQtYaA95xSIyZv2xhge7blV9mW0a60NDS
9BkXh0B/T9luKA8GNvYvntjXAW0Dbp7KaBwSVy0ra/yo9W9M+EHxj36n88AOEOYO
hmRVrua+parmznrdM4tvUnYFvrpN56SEUJcHtR+aYDVNsM8lJFHszGDjJGK1O5Co
H8uREmsu2EyatVx9Ws7Von/B1qDlfUZSLiyAsqXcYDx+bfgilZ0aGy1TcnGpGZm5
3BcHvSzQV5Lj9PwX1Jqs0Jv9CLKkZRvqNa25GpUBePYAPzSQHC12z7kBlewZxNoK
qwMYzFJonbHTYSX/A9V3LhnWhCs6H659DvnN4GL35DRxC78x+1LNym932Kgqp3V/
NMKGff3wXGd383ULkiJpzzhFy7Zw11Rdw/btFB2vuz35ZdmnPMVrepC/C/kLApOg
0Ey1aWUvjM2zbmays6mdTPOxSaa6uSqYMNN2p1wdzH/G/wU68q+70ZDtqMpZdVRV
m7vyA7YI1r8SxPw7GnUbo7grv7HjbE9wSUHEXXe4NDRlRmEZ5BP/9sKcAPI/gjGa
bpYMH8XdOM69hRSJog8AAoGme2hSeBnHyJVuSuZLbHO0/nKxom5m0Ay3n1ZoxOwN
O8CHkuR0BiTLrdK4+2SilVTlaHPz6qgzOv5Fslgw/C68tKlFe4SgK2pgViCv3OiV
qdJW1raNCG8Wm92DvnyUrt78mtraYBL1hfLmNSYrQJhSdHHK2IhLAiItDYIcfWmL
qI9fHle0yURB1k5WeBbIawakuecxLE9YuUY1+GaOjby+M45Blaw/Dmkanrr2f4Er
xaOY1EOW7m7vwdYPzNH5rbAoSNLB92BAy3DyoIKA0t/B7oggtZRhLf9Hmto+PtCz
FHgX6wiTydS00PuiFDIMhFGaZiLT9rEbunPOjpmsG43KGRVEdiGdK5KloYaksP3O
eBLy3rqGTdRMjT4pZAqkj3/B+Nu5xoqjBrgyVRgkhLjvi2/ObcxsV368Ec+aOTe0
+a9FmGty02Arb5hHWcSO580JsuWJdjiCR3UpWogUVk1dkjXNgNI1L1Fy9aCZXpzT
kfv9zMwIuN7GgniS+6aLnY38M8YFqCEVE/OXT8r4xodUVVcj5CSCtSrT2DTxcoM6
GKfIy9LvPIDQ5NCjcMP2AUcXjrCXjpx5CqG+ErBb816G7R1KBPVNzpYmAgPGTVCd
XmwGMgFAoZF6HfuYdO9fUkio48A4G3g3zTQxy+bWGZ2fX9vWQAT4ozPyq9wyBqui
XibYPITWOgMdwHaq434majIaGNrRt/vqs2CiRsjzhvLLgqUAMuxPjUlLFyaMHBoC
zi8ck25xd14xPtO0khcAjiYjsVy0tK3buYc1JyJ/nn8nE62VXN9vdpkRV3CMR3OS
IdAb6RCzYQiiF4qzmBJwNE2AJyHjf4QgvQr3GSm4Preib/YgG6nhC7JF1YifI8wC
t5RvU5CKxdQLO92Y6bHfE2aBhxYTTNLyW5tft5vskEmTmKWRrOt9fN3kPkHvSBm3
InVDqdgwy7fQGJhlgpgYM2L78KG0etal9R1dlreA1HdW9c3VoHhDsKfAWp7+DBHu
x+deWOQJZ3kdZydNTAsiWCT5H2ffoDIT3kx+RSkRXhCpLppjNoJRAIv07CU2PnAS
ryIlpRuDsnpty0+nJhfWz2TMX4tiIZjeKZJKPVa5XlWAVxuGXpsKmYW/1Em03GbD
osLA1ehN4IpQ6rRpIPxsWYdtjTbQrzq/eyzfvXer58Z91GOJWA5ToGTsOD0kkfRJ
NYQhVptWjmY+rhStql3G2eGV8QtImKLc4I92MMe0LW+Caf8uUvgg23kVgfFw1Fvs
JVc3Mu8wxlJLjeyuJZi+LZuoF+PK+dcNQqpC21gMK6hZ66CTdCCVIVakZ340ujnX
/Hkbyrm91pFzpbdVikybSsp6oRL/qGhx1oQXpyX+nO3eBCuT0f1i8QIHO3iDlx0Q
zW8WmFS3KOtpDE/BOppGL/Okil7zwf/gs6KunhT+owh72EB0x40XtnIOUXRp6tK2
oLxYNY9B1m9rruJujaOcKSzwL+tO4P4HzZ1fEMqKQFdJY9908idwOxKGgMvuBXg1
SaiYXYJ2ihBuJ0EocIN0MlZ40RkgYym+1gdTzVy2KYJ0X5vgmiBVK+3+peTgnQrc
Gr23pKrvyszouJU5ZwSupHwGOnfnwt2kPLaCmq9vxv/7omNr8EGBVfmkuL8A9skk
PNW/AJl0K0CCOy34fC4s4hqE86Bcrj/nR/nEygO9LbeqLhGeM8aMSqzGugCpuMiY
TuPXMr/oGyRx0VVmpStnTGJgCaVBgXi+6U3lLNlDfNJn8n9E0Lc39v/lhKSktWV+
pRLqpLZCDJiJqthUOHwVXrSXrPoe7lyvsapFwRsmrPQZkcxrOO95Q/F7ZTLbiXhl
mS+S8krrEg+jC8AyGe8J8mf0pqpGUESXLtRt5exWw7EQ3f32w0S1jssxkOhAyeWm
UimKvJExgiVLq72WwQqV88LXOapAZzhY45EqIwnfPyGzmAOmO5v37HqA7U/UwLLG
5DEq1Lh84TXOLXZzPLTTTgE/a6V11SI8dQUnY83eEs6OjAGjhj7FLEBa8zwwOmMk
n2uhaBK0ZyApqNl6DJFuV4jGnvyMB1UfcfCDjcrgp7GJ4HwJPtjweW/gtHIlq7rm
mCtyzgH1Wziq1TJMdOHfrYSeSe9yt7fQX6o/1f7jW6x8ML5mx4M9cszlDuE471R4
KiFPQ2Bb31UZn21Jm9QzEoc1csK6JPKaBeT+FTDZHRcCYKhfMpoJ008dN6LvPCHM
n8SOAbfs2tO7PTBj0YWnMXJPjW3ritELBcxrKyKWAVNcQqvzf3b36tr4OhL0xAoh
qFqfa6xCy6zSfwSXKWsZ5EYHey8C11eEKQFvJz9/SzSFR1W3y9xDRZizSwesOLul
0dnIRXmL8XeIPhReozC/hbhKPvAQndOiI4Lnmj09Sl/20Z+0Gs9DtBG63GB+26Gj
7yJDoEfD1A7dA9wysstp80HKoqlS/cAu14vpuydP3bEwRGgaUE0bQYVKBwjzMmQ+
1rAfNEb406CuupRYjrmkYl/xL94WUCP6i2Uzy/aL/Mrcjs/AuhDHcLSRsrBYZajG
JmJFETBbHbsYryA7UlEumR6f93XthsjDTGABAFxWZIuTjdcPXindoPMvOnOQR839
Z5u3jwmkFN3V4zn4mkGPdw9Oicfd2QhGlnI4abKPz+SGZBdarwe82SSYU8VCcfEP
iOf96xrUf2D/HjIquJ+6F4H52G0FJxEBLU9HuD0SJ63zzRW2JTIdD4T9eDXa4lSN
W8lwrF4iWLYFs5I2ITkeicHTd8R00DeZZjsJcWyDyb+8NCfLI8I8GEUHcFpnHG5J
1CmsxFSf2DwSfLm7CA5fJ18dWXezs/os6bjW6uZYiU1Q0wLH93kZYh3fFqbtCAJk
fU0dO9xw3TUjMBdw6oCb+dt0CG3E9/CeLrwwUtR98oIBqFVZbDaAYRwvX38bDnz8
i5FUHzP2m7OgjAryf8gLqRfS1dMoLoKx5A0RcsRz8+hssKFuKylNSjVDFRQ/KOiD
6fR+fdSv75t4k4kvPHEpKNLZ73DBBT3J/frtZ80CnKKjcIu7Z4UqDDPMg+BcuglG
c3/FOrzfE3QIeop2rqREp2M7fF7gdrjWHbzt8rfT9/6qPBGtJ5gHDwpBqFkOE8yq
CrB7vNxcFo1mFDMcHktagm44jDj30zcC0eAK1e9oZxnI+jcyNLjZPSHVlRYX42+S
X36TZnvtSI7GPNvtYR1lsNg223cyBsR8nPpkCrZ8UvivDTgEBzDk4vhz9lKMjd/g
5Iu7Ilx0xMj8XOnLrIqy4F0zeDZ9hW0UYmrm4zkf9rvG90N/tMYWa7PH6DeeJCuo
H7yvCVpvEbQ2I6XNCWaxEGftfB+Y9b9xP3DHLzNFU6UAC/c8sfoRhqnpfTDHumwn
XYJvVFBZk624zlg3xqN1M8gu2cxDOiKNsn2ixbFDhekXP6IIoOBkDbIQUYlYyNDs
OY4xtIo9vtZrOYR7N98Fyy9ZafAbSxsS5Zi55UN/TXGyqGshkN6XC5HtCvoZPJbY
VBYybpNQdo3MCL3yUi5oGPwx660mYxdN9wl7zSYSXKQs/8iSIRhkw+nFQlMced90
vE2yFxhvhoNWoVFXBwcrXkqcFrlCabFcMnMPxECYRhqUFH2Kku0qDRSWVlufYiVp
EEOVTsA8nNgonyK9+Xith0aAkdBvpqP7pyJP2ALHBmZpfJ6V3+7Gij5K0Ih9cBiK
oJsySR8k2StA7pxWsc8/lyB/tlur/bobmB6IyqgMZ1GYxuGeyNcjMFaFFB3whef5
AqMkcCM1J85LVmZ7ocOFeqFOi4NmwZrNK7omTQfPmhidkxMAe1G4BStpcwbkGNMY
iKwQzIfPexB6lS6Qc65k1YPKzdbldQSu+kW0QtQJOREXjymYuRRGlFhAN4sLjoQN
EbNDiRK0jy7sU/VZZngz/ZmhnjepoJO7ghRuObz3NbEw48LBfFp7bvEBCxXTQi5d
VC2VFOBV+qTF5jmSdJjzRcKbEIOnLGJ55m4/9J/GWyt4BpnuTvGwJyiFLCBMnTWA
G02jLZtLuffKZ98B8eXLQDp0g8b9GlypHrnsNleeFrdxgyEBRoDQaw51PCHqrEE7
1StbGlBfauY87NfKWc/cf6xN41z7UpVk0LR93QiHo9GhOCRmLFGT9h4EQ/Wmqepd
IWKE5xvdi2uZV4DPtA9eOs3J92pfCkCw+JkVub3OvAumENuoFz3JIroc3YioNikZ
093cVf3esCEmnob/UhLy2btEbh+CQoKxhP3FoknEw8gLDCUlByMR1+CLm8cnlywa
dDHOjLAPNui4lOwDK0GGMMQuhOWN3Zws3Pb6ld+vEi2mMoEJp7o6ma5N4k7m1rYf
wl/Z19JOGwtJxVD7mr9hxjYLWVEeEzO+4xeoyFNuZOHRb5+cB+oI8sHpRHEY7F+G
/vguCFxn/PklZDNWHZTf8XeSpvsoK8NSgoLFSII6/0m5U34THJoyhuvmhYHsfzQX
qrIBQGMnElfy2vcLdRo4F+ownt8s5hEPlN6Ay1FMbaJbPneOOegmbbogxg1Wj2qL
aPrr6hBjt/YvmAgLcT2bBqELcRXbHiytkemihJwm0QuShQ9D/j83r7gWSd3m0ssd
WSct3WRpDVgsfiKYvnnGLNC4NIj99AULUFt+F78l5EcmzhCEfxassRKbIbqV44GI
4fto03Yw6X4hkVK3u1d3DmftiHblXa8gNHyKAiNGsQZkGbQeBeqcc2C6hwh09KSL
HZ42i/uL10SYv+JWcM35MrqWUAx+X6c0r8RWDFJGSNtWl+6/dYLvhMVP7SjuMQ7e
aBegyoqCPcFAiltvGUYyG2V4K7RGL++nbACg5O73ORSXcsYnO56CrzzSf7iAhnxF
mQS73Mm+2F73eQv+Zu7Tf0XpScBaRV0emdS4u2pY7jCjk+aK/wcBEBTcFbCVycsm
2zK2wuvH3nxnnd0AXVJiE20UHZkUUDd4xng2GuOxcVcAdvtUOEZfIM6RDCGSZMnG
Sssg7Kaspztu2fSSgF8seGwQ2+5TP3NMPdr6O0fOinyHUcxDSpFA56KgpG31NdVZ
ycDmB2BKB6oPzUoXLQ7ajV6DVXqtEyEpdjysTqggwN/IeJdzdSz2vrf3XrNJOQVz
C+VVQ6GSa0vm3+Pwv2EF2gopSYaxKNUTuQsXrwTd0U0fmNBGN1c/6lgLpTZI3kBe
f53+ajmEuR5CAEFsPnylOxwa37weHkmg2ocBNS+MNJN/WsWAMvvUQk0nXwa8zER2
Y924KlkXhzy8pFTB9lHzK53/YwtN7teohwWs9z3Srq+tuu/3lTeci5ECnWA+4QnY
aztXFEZ971B5qwQI93ZgvHB0WtF7fUaUljbme7EZmIAdY3mWIXUhTECOD/f0HssE
zLXI3AfwY3rlpBYY74aizf4w6z9GHk3Mf4lxpcKSpddmol86un9464GkYR0QcE4v
MKLDsEd47C7jwbYC/4FTx6j2ocVbylRRL4nzY/vMTB197aY4BCdwYtwZZ8I/rICC
UDsOvNhoq5Z7mQNfnhjM9AzA6OQo9tbsgWYMMRmxvPXh4THrESQ50RbYKDjze2hh
a6FodfqSssSoWzrCIZ0jAPeIQWN2cva9VvSL4h2OId+pXnAKQP3cjEogjOLayl/W
LlKugezupzoXyDPkU9vaHv5figYjh3s+yeRQllOD2urqrWQLUcF6FuMkVp9OYQOR
rbyxr+KHAVkyO9SIW0qEVGgbDmnxVwidco0NYAXYYgV5GSvW+DwXWiP7QI+UNSKL
J7xO6bMNHmIDxrnHb84CpIT/fXWHlTbuWI/kNleV9/st5x78KOdUsdx2oBxqnNUU
50++GGGAdVmDgaeLgMASgaDrg5FXdg16IBx+gevREMSiUspz6iXrPn3I5yhOQtp5
45kGcbk23Z81bZ+uUxLgs0fiCQW37DBVDXtWFKtbmXyji6VxwaSi8+FUZKebderV
MBYbLq1PCko2V3qCebHKAKZm5AvMkhve7kPWJTw4ftnnz6KFFgvS87QMqNfvUIy/
ZBYQlXl8RvR/xgzK3TTCCWDPP0OehXuJbZXJLHwFWM77jmJ7ev7g1IfXx1iWs7R0
txrMGhQ/YPu6YPHX84zN7uREcw8OLpAMupJ+bmmxi2iV74fpD2/nDxQh+6M5Onpw
hgwMCreZVkleoePCYCxnDBbn7+JCu2UxIXAvoA0YZ+RU3FpvFPTg/dV7IXF+MbGE
7HghA6Ny+E9Laou8iSkjF1E5IRI8H8ddyvwZRjMnukAsO/nIK3kSUnN13qsenRhT
KotbkjPOg5yrh80ttbmwiwrwXXuhMjgrbWMpeIdNAZYAeDRNvUGCLqwPtNPzA8mG
Dr+z+ctZivvovVz8XNNRiayHyzouODgUmRS/Pqe72raeUWvVTf6+PtsRw8HCqHmy
sB+kVdiKYk1aQeu51jyDRodb+aPQ5BSr11yiRBuTFbN0TP8TxMNp27D1YwP6mgPD
7OeltBcE34yaFZ5Ncs4fPtNiY0Q/K95UGI/xVabnvVI+CRauoJkJ//N7ifdif17j
WJZ4fSZKwM8JywBF6MmTPaLMxh+oj7i4Y4ggPkBP7CNvzc+wtOqAh1dEPJPSr3KF
6Btlhs0BF3WHPPmCZYnGLP/+5/MlROg/83o/kb3Nicbtr6FaOdWruXEhaYOlI0lD
V4G0jCp8iI4DnVhJy3WHhXRGVakqqDcSohbGOH08WX6IR5pp75eBDZdbDiezSV/t
IKuDuR8VOJgvojjRMhbKH4uUpuww6M32dQ5sBzhpd8C1Ov9OWVxyuMw/vt3RShBw
h7AMz2feR9FckIPZjdcwwSZ3dQ+JRFZruYgsMMIA08F1/1ywa6wHSIb9WLoc+FlK
3lmuhPW2S7D41naCji7aEtQUdEsof0byAoFTzTV+WY7/T/LqG0fn8UclDQ5Bm6Hc
YzANYll/umg14pReVtBRMA/DLIDnFiDEqOuRgrDyaWT1arUwSFEhP0BQT98ghcd+
R0tYvbh20w34LxsLar3rFP5KtOB4KFaZ3frjDD9e+/px/VcEayf/Zy7w8Th357Q4
evzMYDXSet2OIfmNaVlG1i12qPhodFezYYg9fOyVIGBlLBlrOgPqc43kXOMejwpF
FDVJPENmZXTx82WkLp+SZ37jyYD44E3yuCbaZEJoSzm0Sko0WG81sZJ6XyUKGl7l
6Zld88LMPQIAmLWaJ6WB2kOGBB5WFW7kLLKP7N/l58dmgeqMHLzPQJsy+6SJ4+lR
++9rr9sSd+OBN+FMpho0oHwNJC0oljB6gJshZ+33TQHvQguqb84Qi8Da30NY9JT/
1EWBz3GwcKu74wyybAuToqhk6JOe1zQHF29MpVIwJkgJfBBcktFd0B3bhW2hhOEI
4IrmqzpmRdAxugYK/G9BxTOOkTEWRsS/SNPrEREHWUjkzfyniXIw6CnJwPdYyMCB
wfK2WzaPTgbSuC0BRzWQ7WND6mtaEKeEOi5lfVrdM2aKbI4GFODaW05yQZcZ0ii9
LvO3IJ8mMyeKASsm6UxkFwzM+/4SO8dyjCdCtAWOIp+uWbNNMA6dDKBRp/q+TrUw
wNDIVpo5LT5YizGRR2cxsoufHtfW2gj8b3Fa99LpwLcKNIlK9CGXO1a91nvepTcI
GZ4O75eUo5wpNezU3BaKuMKmJsIKC/O1DbXvadCE14SoCoAQVvYbSJWpXGTpGioh
v/tGTSc5m7HyFVxvpTsf1U7vpbBCHfI1HbAtTQene6b+zlF1Dx1iO16mDbDtrHG8
TRxBzag4fbxDaCfk8NIhtTdQ1LAepxPJGq8kb/+rIgpmJ0IjmreVXse5+BNhdhPi
Gzum0CRvhgWM0FktuOywg75icAcH5LpZganwSJBTAOl/n027UjiSCtTZ7RsnT1UR
STAD4Bltm3B5eiN7gpiWbmh5AWr9tj4xjQGnBZoyUroiHMoubtT53iJ+McJpNpw6
48tqZkcf7LzPsVcBB6G6Lh0LsUUvNbwh4cCYsWLdN6mZTvMsn1NJb0BMbHJrNy8G
anHIaSDd1xikICbVrovN2Mg/0oqaagnrHwgx0AklGpLxCll5rCjFCFxioYG3cG/+
20HT1xXaBli4S6+6a204AvQZ09Xo7U1PsdHSyy22ap/6cq+sD7jdMCDZFtlpiz5r
tz51yyzcSEC5l5PFi/qZMsxaZCGckbg7zB+rhrlE9CH4NMvYY7Ln3KUtyYZLGJJo
jCVo7AytJlWGXIgHJtpa+CuEbRwJ7ust8SIIPRZP7SB09M9Iddx5ObO6v7sXo66J
R//pmOSVkCIDCEvGbXC4P0rfEBGIoIlUu0DHQZpefRvNL0mWFWJXN2/OKZr3y4HZ
B5XzOfP1mpm/0vy5j+HOMeI1dcvodaX2UfmtMqG3o24sCiruhsFiIRrK3+KwJBRw
dSdCkaM234ot7fuk2xhC/niWmAzMJV/DHhGTu4Epab0Kv2KO6lxCILbnyeaaQDSq
5/TErJ5npNX8+tfl4Q/Z3GIoq5hnCLKsd+Ib1QUQoj7+MuLKg+hRReCrj3/Otomc
/uwR04fiDiQx0wOPj5i9T+owRhqa/17DYFocgSakt7KJet9BNsq3EmPcC6LaIBoG
sXqHuhgk0a9y4iICo22v/VyyrODynT08sEIw/yACHO1GtSSN1+3tZyoqqn5J6y3V
X/tSXX+wVUxBCb6lEjY96tyRAqp2s4XGGJ/PYwL/b5dpVQFsfmhRjCtWdkzbV/sL
tWUNH3dAGQhwZdwEpIkhWmNnKNssthNqwH7faQ2H3oP9/E9/njZnvqdUoFz8xCdl
NmuKrpW+dp9fB/0JLoKQwuwmRIong+IOErJzf2KtbB3y9pE+H1vSc7ewbNQs7Q7X
7vruIGoumSN7NGTmj2dvYzLbglc4YgpNAgm13KHuLDrpkPQXSb/07zBNjUpitBbF
JmuetsnfPwmJaPcw8ye7V+7KNwgHupLMrmAccZiGXIO6IQAVoYjxoaFdMNE+qjkH
mWyQJwV0kpPC6DvzCuMO4U6NG+heby9n9jX0UeLCDwIrKdUNs7Xz7zHyeIX2fk1q
NXpMkWlgPqE9GnB8PHTG734ljcossQ9JNpYUFvpTY7QrKNpXWQnHVjWxjC3ETEXL
LYtnh3dZWUN6oju+LZ9oILamx0w5BpiNmMruCnmX2zzXbAfMzON4TfPlPbJ/dt6h
YLHZoLrUYRZyWp0tPH9MXh6/EH9ZTUnml0rXKZ2IQa2smPyxdX/lts5Fn+ROyj2G
TCDWArh/pRg5bVgL0xPeyFpy8R7fMc0ve6WplgBv8X+JwgiEJ7JhX8ZYnFLwc3pL
MD9UwRqd5NZjBeNCYt2/jEuhQFIBD+OVTSeb8jQPFmQsedLnBjrtUHIjM5KlH7Vd
d2yCn7WkJEkwAxyJJbcZR6bsadX+j3DrLeNV8VXBZDg3vMP8/zY8t7MiU+DEDaWI
lr4SO+GOt+sMfzMGAHG157vceZdTXnV8Y5aRFdIzYM64NNp+869yrubA+g2IPuEy
XytpoLw5YrjP/52Wdzh352DRWD86D36AMfqFYyE2o/++rfcX9/TEMZdIugwljR3/
vtIeaKc/SNoR++FHWrdXHdv6f0NE7kIjL4lbqE+5QeGNgcrpvEP9NlXc0+gjsSi0
3VFVeJnLm6Df6q9q+EAqz6jSPeFZE50s/WpiCqxhEqDxDbjfT/vtRtd8VrxLWXhl
pCf75OTpXgjzoh1rZzokOE5c1Ej0uaFkl6aYc+8ZxHEmF7GTjcFOD2oKRK20TU1G
HjRyhGvq1l7dd12z39Cc6BfUvo5slYcfXUmVYy74hOv2e8/wtIWWdly+DVPZZqKZ
kERLmgmBNgr3VatDygmSDSCIFuHXKGSlzEkFG/50BuBWKu/pgkZt7W21vjvHpEpp
Wmr/Vz8LCchWyah+LGQEsWCosMAOaofJ2JunmRMmkN3Q1HGv1FG78NIi0/VgqNJS
OFM72hVTnT92iVpD7swXzU3p63owXRwkgNhapaa4V4sRfY4NDyWqoO29Lz4jRuRR
ONbFM0MP6HYkfLAmR7ARPdbh17t7FJkOy/X/UKe6TA3fKhTpj13RXn/flk79XgA5
9vpy7rKwRm/SNXeG4MSfJGqU2DCPu/ilpkJVnc+PE8PJSz5U0LZZDGRcN10r06+1
KDO699Y5vZ+oxvQSNvmcQrC9TD6LJa3fH0sbweq49/0CAlKTCX34lFnQwLKoCNwz
eSiwuQC/u8AYBZdlgirOMerPrH5YVZoF1H1f3G43Xfv3TDj8YP/sLnUnxg/v4kCj
CZuACi1UJGvorW5oLvVY1bvX+Pgtdu2QJh0huCvIQ/BSGTvSttJvUMYV0/wD7ong
2hlmbBnRrci51UrDFGIAR9quqKPpXdA58AR7+PjkHeZ8mbkf6+csB10ONAdBGLLX
6Mk+Tf1gVPeRrA60MXn2OtzSGHV0F4ew6Mb5vPER/ReX1d1shx4CtuhaEAmy87fs
BRL23/4tl5wdOgJnI93qVMLMGi777LWe5I9LeNfHc7rRqps4YL97tsUbIHEgg8ch
wfS9tzhdO3jPKSNeqNjXWktLb7Kr8peN7OnqvUGVsKj3LQiUWk8yPYzR++iq+KyN
7L1RcRJJB7JHoAJzo+nJ6pn1Kk41SDrUhWlqzC343kpI9s8M5jUy5u308INSSfHU
hrl0Gplu60ssJobc3RV4MHHlMRS9i5SY1A5L8R/wIlW404i4rodw2pDsoK7AGgmJ
z/jEa/zgwf/4278e3lZhjNv7LhsZB7CW/REA6LMCWxBQw8pM+3GFVP862H2o9+8z
/7hfmLEWdiK3ripVwfuqgnO4Tgkqze+oC0xALYjTqg5u3l0hWn8UXdjwXGA68wQV
3G29lhcIobsVDGzyDzZJemvuI3xASjWu0x+lYPtiIEblLjS3sAJ3wgj/dRsKdFvJ
MwZZrrMOHQPtz3jeae0RhwZ8FXeCGOsNuqzqsZry8ezIyYpp/dt8vTfkKWp1mdUm
4k5mQI6lYseJp64VDm1qQi9pIP24GanMyWI41fKX5MuZw3tYgotSUBvY2QpULgoS
r66uznSP8qjh1LGBUmHTjnXTjWG6vV1eC8H6UW9PaKjR5a66q6zBcPidOCfzdqUY
0y7dFXtgXGEZfLPgHnqJhCkUg9xFb7/grH7D6qDE6zydafWlfSq+efereH0e5xJ2
zzOPykoBPlPxMQeGWWLSawwIEElptFsF4nfZZP84JHBvpc4dBfmqLDU7tSv2JKWz
t3woojTthQTGJ9msJ8/5eGf42X2OhOvWfuos+fL3DtwD/CWqiSNAb2xY7rPoVYeW
28SEC26F7y9g+Cc0DJgP8qUI0FF2Ycp3bIqO7W1Ks3QNRAWReeBusfLfICf1ey0y
IsWBH2p+q9/arrAXpn6lTj5n8UeifXzEF9fUBXrKLJvK1WU54l2k+6anYSeSY7dr
6cQYhY06Y3G/XPkocHva8ODbkMUBlbpd4q+hAB3M8oZ3XEvq3UwTbl3G5RZTpIoa
UvZaDJXkG9gQxTZXv7gYBfhU5FgroHB6AjC3CbgyNMXnTtdEocgFvPAaOGK7pCpG
PR87CPi/4CEFSzgeAQF3c8SXPXrHjGIiTTDh1c88bBGDdZqod/WAi+Fncc4mr7h4
vb4f7LHKScw29iFl3L3M3X0XRxkW8C67uUjU8p13ikvRqIA/X6a7DFBNAzcH2njt
calEV+70nlKEG2yGsty7P3f900tdEsH2GL8LibBFzcXbgGHipadurRu+LfRH5cAu
eeTQuW8q4QhEg2KpIA+dX8Vsyy8P9XLYziY9O/LrRmrhocXWXyvqQ2LqEJVOxXBE
sOEzQLjcTp4ff0SsnNqrbNec7xOYaM8TJD/7bB+Y/vh7ChszuA1fd+FUGkZawe4H
UBw+RHo/NBz+yaH9OiqU3woKGSRuEqG3pXOWWcwZsNCJ+lIlrPv/QxdrfDGMuTNo
QxDsXMkOXFo1bg9MWYO6CO6KnULxwRCd1CX4fc1ReNpMjkTosvFmIwNaVmjKjNbq
EBqtST2gPx3Mb/0Jqxo7HHj5jnq7MjH+gi3PQ6GTofRsBDCzNTuRTAAnifTfNQjL
BxPq06rXC3iKlVA2vRZ9aPZxDSFAueTx1Araro/9Fd1C7UQDKYtEqEcoutOVJxGv
RMHiC0D7EDE7FI7C6E0PogV0nvTEre/ijEeQUQD0VjjeLRjDC4CkITckKCl32VQr
gjnTNMmCKmMUFazCqPxD2HJehmYdkwUtVvdmlG/aSCXL1GW5E1VzlA/EJynIgD/N
fzgzUUAACt/L25SRQeB99yKeMK30BdDWmCScSK8JVjK+RLN5jVPAndzocjBk+/nn
kQCgg7WgFK8cu/DVlaG9s8EAVl1zVqMw6dJolz6Zg+P5qJQoPXOyZuTdYj0RnNSk
ROseopZ83Y6JgzxXv6ujlCRxMbTCptWGNReGrN/HwuBcwv74Un/EM822jDR/tLEa
xLb8w9fOHcgrtFc9e272ylmICQFkgWv4YvP0Go2mYMkntvRAY/KH1HQlgE9Ba0zG
66WPlQ1UoK/4rsFmiCzDKjifLSEyqxDizJ7SuboEqyIdF2gfd8ip4iJnKaoMAuyb
PD54fxE5nhK1BRlICBTPkENNXGy0qtMqDtaikYOottio0Aa6lFz7m2G89JSwACo/
ABL6cg+bAWsf6ZG6SNe96QnSPkAdt+uxJ/zLY+HrFC+XrNfkCBlbMwK14RFJ+iA4
+JKrbTPxst5xwk0hW9tKsuNftUtSBIpeaiHdYDDGh8SksqXrG6T0Yu0y+BJ/Tdgp
PYo7MHK2oX7w1VQRpu4qLzamtWximMbbIUCKcs3zxO/KepiI20yhMC2vzS+ivoIb
bvntpeRVaTPIvNWdwHx+hCY2JsANaR2QdfHinD3185spqlS5VE3/TKKpmeMiOorY
rJe7b0IfP35QQ+WZuVZmn/jk2R9JlON3bVQEe7R6lLe5+nZCheyCXQcgIoBpCGRt
FfAZHRDISstwrvZdBqoXhMqkisDNyaUt0Mx0y6MqeZbPK3lk3fpnY7Cx808Hji1k
a0/u20JRr/3iY86U0gE8Q5nY8b4v4Lul7ZZt2IdNKTufOlZY842p4Z88vaee/ySf
72BtRZHgc6l9IgGzDI8QrMtTpRy6UMnJzQmNnG+kc9Bn6Armk8EO7vNP8wRV0bPn
Ck802ZLt34qdV4apHjVTBvzAN3mwCz7Xy5o3z+zhUU+d987497EJTa1A04OElutM
fRgASXSq1VsDUdfNzfvMMyuMDvldke4tPSI8rO3p/OINM1WatkrHr1rbqswasPwy
4vGc/E60cekY4EUGBJPRNQ+P5punKgxlfzSafok3CZSoZ+VyVq5z/o/zyis+F2PR
m+CTXc2fgTk9IMtqdKO/NlKbYc5DpduyQyzZBtpKguGqtxvkGfFd+CsPQ++X4QNy
UG2xX+rz9+SXs0p6U0AaAiSi9N3fNejiDX0U3KhpQ/5AGCqxvAr4KCwz6gjAZt7l
d2rVaSD8XUshFmWsdgwECwBQa5V11+nZaQik+lK6oJEbaEesgA6bRGqXzzOFly53
fofnsubSrbAJwz/AVk0NPRcYOd2HsHJKk60mLshUXkQiJt/JoFmUXY2V8ZwItMEg
uH2LV6JYhhGpRK/b15ka2m+VuzabXWp5rcUcW6Wkjfh7Exw7XD9hmenRKnP9yAEf
3LDf6H4KR3SMWKHYK4tM41jg5AFcy2yYEpWDVTIa4+sEVtONYCAqa60dUBtY+Yia
Fw5xulzj97LkABJSQEe6i+pjZoXmvtKi2vXm55tRyipcdA8YnxqUVGml+L7RBneo
mzJsai5AoFXlWUoeyl7aasgASGVZHJs5qDcqVy5aleOo6ee9loo7S0Zh1menWVww
tcHKvwsOLPCf1Egb1dS5PbkDd5u+aX1/sispBmf6MMG5o7uLKnXUHfRu8KopEC9f
SO8qLEHMz6LD8GsYbbrjKLRxFNmOlvWuIcTq2Bz2baW7Un/kSzXRb1G3xz+Iteh5
pCmN3P59FqkktVf/zGcLT2xAl1yB1DyWgMKo/Ex+cwhdOKIae/5BPTFykrrUQUCB
V7c6O19errPGxOMP85TzhBP1uHvw7CUFopjDrx6y6HuvhhAxygM5iwctWUEa6uZp
RbOMPiwWc0QVEBDNxpE8Z/en5j3vUmrLOqXYURC16+RwXhXC67GQyrIhjaqEG+xo
eSNWbM0KAY3+yBlpJQ2bo6XA/A3DxHACGMD9ng723yZ4LiIxmP0WXvpFFZmuSpXk
TuAaCLpw+Q7erbrgKb7D1y3GTYmGmkWetuz2AMXalfFOSJ0qi1YY2agUAV7/iUgM
En2gkcpTGEx8DviyuSZ9kSJaWQ/Q2VBOGSWZjgbUY8wlj0TxzbgGurbEuWisbcA2
2MHG42aCHZRDo5YYdI9db+Nt9m+pWaIZwedIj0eW2Z9DSfpTuafsGnewJ7SWMnON
AO8oggZ30gRdF+O86TvXX6iO6qkbJKCThzqi/f9sfVqukUiW8pD/gxRw8pbE7p/1
f2n8bkVEvhL7YjHn6ThfNVTNKclOJ+LkKw2DRiF/x01ouvgN7bquNEvomXNrSWb3
ipnuAhpWpxTr2oCNuxt4ve91OA1FNvVORAlOjqQJd1YGXr58/d8PD6OVDRKmjvXw
Z2dnw+JMgZqxyekHnIRMpd67BHUS4DaJYzjKusv6cayMnhfRlbGQy4/BhZixwqs7
SdmDfjvhOMymdVz53cv8fO4u9zPFiyjOtOYuNrnUgHUTaqPhBrohXTsJAl/+rXWI
gw1NWXYicgHYr6WlmvjMbF5XHSoWqBUdZgmWt0gqh4qN4sk7rdG8luWHD/5anbIX
iVgGsZA+/MQReSp5Uy8rl9PQZdo7VQkP/gCfUusBfg0gW6Naxh+ZMK2wKuVNtqDB
GZbQ0oSzFPX6tVEBJhXPXHLK2Wdh+bVy4NQdFgXoOoisjpE+o8Meq1G6HOkZAbUV
Vc7Sd14QBjV4ofCmDaMfqkbbCUlez0ocK7fXFOAu64/cTzkhOibF8KTbsLY2DW4/
YMBmxAS4/4xlf0/MTvi0O7Ma3GP9ZFBkG9GjJRnm9rUm4K5FKOkw6IdB6EmXiDxS
1o81QDjUowrU+1IOlcdxhwT9fQzALNSLAbxbAfk16qwBFaYtcZW+T4eOo30/kusi
qPpyOUtalx66gcqDhjKKgbPz/TtG/2RxF98AHXJO0KQtW57Ofb5HUtDSR4drpHir
rD62famVNxN191ON4pWaj6dPOsIje/1wJ/LBPh9MUTmT6RfmGBGft+6KLqFNLZYq
zvFWn0z3gpNW//MPrEQ7k6PmHsX5JDoafXmZLumsINY7N+A2ffdDT0o2M+6OQbH4
lmAHMxntUx+zSyZ/uAv9PqiBoE6PxYW5lLga2glIBdy/SfeiFCSv1wdeCklIh7ds
BOcl5nUG6NkuL09dB623iUYxCBkPHGEW3MTfTMQxcWIGm5+MVZGsDlq8kGXeOTnW
oAPng25wK9L2cPuiKByWlYn8VhjggyS0Nhpw6yjA5iWO6rLq+quqjXtGLKCsY7zS
N3LHEeEsbkB0FwSuVpyEsZjL/SPAhg4mw9G8Eq6aKBZOZfg0h60WTeI/ITHH9LVI
kOIkRIIcehkK/4H+YO5WB7d1dhdqFJDJ7+CFFoul1tdJHbrbIUxxLKtZ5GNDSHcP
Hf/syzMId7UHGani4qczfQw+sEW6co4zduHT/m77+b/DQ87HpRRvnqSgcaxWzKJ1
avfMmtosoFChF+BLstBhrEuVYPuxD5zoM32DH5bBgOaty9a/OC1QBTcKlT/T7Clx
EirW05UM0JlYTC4QyT2pxdrEGJJQ0gEwMOH+Toq/JmTtlPRZIEuaJldqeAMPZcZX
8BKG7znAWoZumwlnRiOKa3ezxSFiLoHWeN6wyLJ3kdUtHRVGueErKEmFWzpiP8xK
++aoURZpyCWN5ihaj150qgA2ulG7QPyQLXlY9/rl3yRkZipwyrcdEeYz1JuMTJAc
XQJ3/yLjEL3WOz7enTvh7VRa2ucHJI5TogbUTRFAsnEcQH6VhR/cvXHxozfVQpxy
2g/Fj1LB/VIkw1NZwUD2CUp8kQQIYdlxlpkd3FZR73BFbhdFqjERbFtpYAyEb7Z9
zhBYk9TghKuGLWlmhn2VfD/vi1W+99lSt4d1JQyYDg8/SLa8QB2/vcwbNOO5cA8F
ylOI9Zetga+wzmxdaplNW1fuAtN2VIn+nj17/j69yiBqyFCOZshLrR87JlQCuoNH
D6cZPf0wmfXSv6VcpqBLUtCWXfd0TrXLqtr5flFhb+trR3BPBST14+iNlrhf8qOg
9D0O6kbZxN6M9/An4zHFKz/UzjXPr++QsaUMr+tLdB2LHKlsD1KyMTNCanQxH+B+
56dClQ31zLfpGlChLmB4Q75SgVKrk9zUq+GFIdO4PpXrpi2+vuoJoVVhHpgvk1ZI
/aOEtNIURDRlHdAY+7eZr1fx8fy3mVUd1947dk9nVyxlLmUn1tx92zP2m10e7Ibb
sknC9B0rrE8XMzOpRw9MuXghoX1tb8jIgMGWIxkeysFgbuRd0buAQOaoOn3QfrJk
/kUJI15gML4bua+n9SWdiq3Ig90cO4TNbY9j5dfXpJMhD0Xc47jAYNgzDcFZsubL
bZucdfGKi38w9nWW2wRtOO4MqEIhEHJooreif16MKjEoAK66uioWc+lUCz+JC8Uc
MoHbQaoIPz2Wmu5uKigPycTqesI762zHzZ/L84gcKqWiSQkAmDvFakipJdBPSlEs
66Xi3ny3n4Q2ggHgormmHfUlg4KxQKhbsWMAvGqhvzGi+nY1eIOEbY+h47LOBt1e
FrkJzlN+vlot2Fpnj5Gr0H1zmTedl5eozGmYnxFvIUrhrpk0LWlOeFcXRliAmKwo
k3HufuwlAGVvo05+ei+fZx4trE/XM7yKdf4NHtxa071NU04Ejj2HEj140EMgh6RP
Oj9DCma6HlwURUBsrd2mbX37VADB0pnpmRKIh3Pdlyds3wV6lEzv4PnPEiHZ8Kko
bMQ1DkKrOhqWo97Vl11BH04vIJVnJ1Mfh0hbw48xMEnDHW4J4YkmfttSy23vm7ok
Uw4jZdvbZr6HUWyX3sgej7o8Xoh+7ZIRC087Ubf4xDbKeWAFvbtjcFNRpFhFGems
KlUYdw6J8fuXSOH5pXuxMw9CryZbqInrKAuOqtrCnFCTvFrMkfWH72Yk1QKK5aN5
lHcRuJzsomD4yDnNCzixEw1BwVpjamIQs7Ith+f3Uju8woYwFnHNDzDK19mphfrw
GyUQ4tSy80fcnZPNvHPcNFwXsuVxy0Yq7xNadpUrhdYQSfXX5cSLpr3uRbUp5Vl9
zPL0DeUACWPl0Ge+xG1IZwu+l51ET0H/16lPdiuZA750SbYIXnYbRmeTAnxOJld6
OTre6ceaIRaprEGylCGpD8tO4PMmbZrPisPel76K8kbs+UepajE4sshE23oZGfkj
yQVAYpRGdEZ78rpoWbo2S/QQNd3QPFDfl11+jlo1/wSXrJ46IXYyIfQQiPk2Hhwh
AeWi/S0YJmMQ76LPi04vQZp2H98W7e7/XjFXWBdbPhFZAf/nzaOMucj4gjgAOMQC
Ogs/4mmjZFQkHs+HRKYggoeNylND+v9FYXadZ03HcQa0oX8eDOj5YVj8UmrFIsL7
egO81BcSg2iMjVsdpFOAeKDLjOjM4NcjNclk76qDWoPn9rjMvzgSntgqg+XszHv+
K94borY6ZZdv/4cLIPQI3uVRhi3wmQG749vU1OB6Kpo6R7cnV4v9s3aHZXsB4Ez1
JyEQpXt8IuYmTQG/1LI7/SMeoR5hdTsiH8wGM53uZ5L60H7GZ1589MlqGMp2sifh
KHugp9LN20OuPDEnHtPhGMbh99zjpCUJkaA+ypZ6nl4WRTn75mkETcQVfF6a2UFt
NBI/2cMta3OjiY0bXMPkY7ShAIbMUcKhkSGiZXF+UXeyIV7SZF0tL8eeGNB7LAgW
gae5KXXqDj9Ia/cpddGK9vMD4wlKOTNSqoEpanRASAe+5MM96NFD/IVCCcchBpvm
CqXjX887V3IKuq1fOP36K2gPnrta+TOMvht+T5w+c+KWzNc/ZpomU06Zrj+lbZOp
2EYbu0mKH7nNzIQF15/slD6vXfV/ydw0cY3r/04JE7ZyN5Fas3wJnXY5agljDNKk
0Lue5Cy6WfVGU7kmysGwTXIW+QYgPeRDjVnGtAIxfshxMhEpYqDz4ad8rWmc5JPR
rQb2h6csYGik5V4hTzKX2SdJz696AMPBlIa9Ca3fPVOfses+75mYN7CxdjcJDEQ+
7Dhfvw+/LtVJdmTHY1fla57O+EGDz4riqUxph5oJX91Qso3exqE6zcgaVEMPWVX9
mGkJV3MUvdxn+LJy0FcPg3iuFFiQ25/TeTJ/peUW7ngGBeq9DT9lAya/jLeCIPNM
BgDOMDPxzXtT8iBw6ZUFc3BxQGADBoJWqLJPKwL5nAlYyZ54RWP0f+u0HJn6irej
c/yOxIeN9rzLxtptXVym2hvx0O4HhGh5W4lJ1tWGZCwnNttvDFMztq45Pc3r6yTB
qX6FClKkz7rVnI0YSfH7LXwFGJbrelpCiirXC3xdL+2M8kDrp5FpYmMyb3AfWRlY
qeGJPc8idKKQtzUtk6NSV+o7VF+iAyQ9laHd/LD4FOtzpUV9khz0aYH5cJJLNBUY
bwjy+zCyVoPRwOWUzB3xshNw21JVAJcoU24Bb44eKa124Dnrtf1wYqB4raUFuGas
EoXCgA//HAUr9EjmFi0tlc+AmBASsKVyWTjfz011E4oMDlz/ANozPW0nGtLjmWN1
Gh2/BwDP7hxIoy+20XnfJOeGqL701Ua5L/VjvoE4Ozdm/2ROTE7mDOb7leBSBtHP
MDPDNq26a4bBTzg5I5V+wF3jPAjy67RZSTNBbeGKSB7zoZGHTvgxV9NqdiLZKOpQ
jNxPdFklM4qDjohg9GShQOavmsT8AUTgh+sA+lI3TOQBN1fx3WcmrpeAGVmM4CHd
TLp6ZPHD9//wRcp/JaTmfW0bI8g/HcP2OZborCCEzgAo1BsWEbOU0HGTOzR9hcau
R0CFfORd18zU1Vun3AU452gU68tk8zJvre5p/+Ewz5qHAoo7F763tTiFd9wYW8uA
bFkT5LbTXbelvCaXNE6mGI2zcpYxkiAu5gmxhIfn1OsHSTpw2S+/zjExwyWxqqj3
96OrRlUNbHIfm6Xz0/4Ear8/cO/LWys+KG7WrhK+AddtRTVp1/w8e5DbPTKBJuUA
wKV/NS3GSAQE+hw8DK8YcHicqsL3VOa1aILvNKJTlwEI86dymDkQzgSkqrjt5I/3
Ataw5oCJLrEUbbRMiQnOuzE4tqSC6UfHrKDYtKsK9xCt4oCOveMpWZ2aL8H3q+pp
L/POW4Npo3pyfl0pk6vm5skizKBJHp4XuEj1f6uSqKLdC/Qpdi5mX5L7pTtq0TnA
kMMCalSaOrVufgtePkP+ERpebbMM0P/qWvxfMsQvoAPQYQk1cGnmC6NKF2mdALvZ
utbcUtmaHIO+DJ+DUjTBoOyqf8zqg2ukfpKxHvA99qKD5J8YkF4hoCsAh0ruvKpy
dwkPchz8Zcr7hEyrkUxVurth4aETp/rva97lfrp8/PtNvmlPeGzGp2aEhAEHG8Ln
ok2g2k8+AQKwtI1G085gjoD4I/b+0Z62zdZAUkve4wYgQlazDvNLh5Cxpb7hw8cT
peH39IYpIvCXgG6Wgh9G1kRQW0YUbQju/BbR98JqbcqTWpFE5w5NnDskAnnbuHxQ
J0u1HyVjGSlB1fGOxoF2ipIHwLMXl6A1uISNU79F/TED5ncG3CDSNEX511C0Ag9d
VG4FXy/e0PpjcDL9gaJBpedqnFIN+rCyBgj6oWmNw76VVI4LEm3/u63ZpatnqeOR
1BapdFQ8TjXr5vTn9X1mvZZAAom0PQug0dCDWomgzZxM04HIc0D8P6vqWX9VfipB
K4kNKanEI0iE4l9Fq9P6ei2kAn3kjiSDt3994eDuKfUnXWkpnFx4teLCXpWNfpqM
ETsNjc1w28NkRMDJcckbxcUs5z+9JZm0L0uS2FPO0EELVtnlTdJM6QOigFqe6dfJ
FsOkKMhSStv59puocDccilB4qeUWroAjlR6C3CH2VFk10JqnwbEB/VfV4aFlwHjV
jAGi8ruYrEH3g8Y1PZzdEPiRDasC0eNUcnRF0b/Ql+uh2yx6KrOU0Wlg8BKXV/Oo
+1qOpEDrOV4FlYeHdtK0whz5rwCCRy5ZI8ol5DV4X1rjzOTWbpFIMov4Nofjoy2A
etERrLDnLeq+HLThEje2xeMc2odLowiyYLLeltauWJ8xwuxoES1NIy6i/c5jO/Y/
0UXj8SvkoMg7S6hhqv0Dj5IqdfHj2REjfXR1XqI6tRZSaawbxUopaLrcUoA6I+3u
+WTaeKo+R7YCkScTBdKQyunD+SC2/cZ7DWnoS5OuxM8CCxKq5PIQpCgtEXKOYXZW
SQ6v2uvH0i/8rEwvkCAwn5ilh5Ql6Ym+VwWpQ7ZQAPWDWlCbntsaE1ki8JG4ihnt
a6//0Y7mcdqySgAqTJr//NF6dcq7T0oeRrHIfxaIQC4ZfRjXvuSfNSUhP4LpFkJa
UD65XjUtUdBFuuccfUaQBCK9ajyL7d/EC2Ic8mFiuD7UMLYlI+bknBftGEoa0j9r
hS097LH2UsNcjQVF2O4obMbJRXcNIf3YrfPQEucE7Gj1dYRDEUvmuEx2uHD2YftB
KA+AqDCqRHDPTYTdpN3j7NAROfRnFz1HxO0qS1SHwfikTaBV9elC0qrPAZrs9g7I
ZTra6VtA1dLEFUVnyDn95N5QkcwZNNb0RDuSSU+WNL7T4oT7BUenhdyjFQwPac1r
zpb0Rf67/V/RYslvRPWVf9MQt5UDGYse3Djo/Bq1ePfVIdQTkRC6n9r4twQP0E5t
jkARox35EUdNSXmazj7/qy+5k9i7Of6986p5HsI6Dnf+BKf3TmSxNGs3SHM1ICl5
0EZnhYD/HrpUyAg3uBF/PNa/mONdTuZXfmiWlV3dTTCQDy45HXFxYJcxEGSV4THF
yc1Ak/QkgJ6pqne/h9HcC1vqppD4P1ZixGBMKBBmw8ru0jQdhfIbpEfBaTdwBf+e
GIxAoQ4OCBUxEvu3ZyhPAAvynEEcCvqiGtajrohT9p0qAS9sMb9ck/ohG918RhIo
2XyN0IVHP4UJq+mCDZRZusq8gYAy5CT4BLF76ClfV+7S+F1oRZhszESLPPks6m/q
cQ+u4kx1fy4l0gAcZ/1n+cVRo0hwgmTeOR+pkzMxMdfS2ywJkdscrLVLjL7DQtZZ
I1HM0MuvIi+e/rhQvK5dlcv5gDK0xyg356nPexlOMthBqgxIxoRQU4sCgOUgU/JM
/ml8Zw9x6hhvqKgh9VkupSWZC1aWf2lQkNpRHD3C7WyDOWOQxD1Iv2YiuQFcUBOe
KZWein/ccVnaCfDpjI8auWTGQUcJDWUmdzfg0zq7s0hQbzQT+eHItGOu/BRG6Isx
e8E4t8/5q4a+HTjofZZNO1lDRDohREW8R1fMGz4QBcxUC2HBwkf2JmI3BS9Oepc7
45SiHeD/NUkRWGl/9ux/99O+wXZ8YCUXkZtkEMDoWw3TyOKjH6Lv9NX7wrptTaEb
WD4xWy7iqxZ+OumBPnc5++kPgLAdwG/V2TDdeBUwTM9j/A19cd4soI5KTT5PXwfv
97BSKLjTstPtyEkQpJIOrESkoRTiGQ7NdhLXwF4YmdvrL0N2LJ2XEdjhZzUgFdsN
zX1h+R06Y51uH7KFdlvxnbnbITMzh7usBcgXPxUm5cMgUJb5Vuijrox19fJH9cDl
Wr3Xh+EZFewFQ5WUp3jjMNuR6eeIuxRSSVn99qOp2nwBChF/K+3kusLgQtVw04v+
zfNuVI/4fpKPuXFtT1oJKyD4iA+VHX4CMRRHUGxwWZ/yvb72LJVAepCdo4VofV2U
XYWOX7cADCj7jmr7iXSnDiZzBiaPar1cS8JJONMHdAxNY6jGRPNxuA0ILTfUoqwt
3++pYxDeLLIB7Haz7eIGkE9l8jFFynA1brqnUav5AEyvqGK0G0NsoICtgjG6MB5s
ai024n8kiIvDvAS1bl6goZERjJEsjhup62kYSq+9WpoZE9QxaUJaNp0DJZ3mgbAX
FQeKlihbp9XFW29OATKz14beogsnn9lZJWJMKkDa2QAUi4iZnq7I345nqz0TSdNN
Zro7aZZkw2k4cjMgBwk1LWkvfAuNn0L/RLzs9cjFygi1t4gUUcF0yHWSVh3+rnXW
L8RJLBTQe+yy7+vhoMLPBq1SGfwpMX1P9UuffygW6x0G2xCYxYZnPfhNPyFn/Npe
b/Lk8yUPha5j+4NB2VaSYTgM3U8ni4HRxfADr9p04fIr+gDRe72xWXNNLd+WJWNd
nU4B3hSS6/XdlkP0IkY14wMumNYhj0ROwCw92Bzo4yvBhgL5U0VrnhDt2G1bDdcM
xu/qtkxKYWepFzmPRJcwRL5uoT1HB0oI/xUO2+YAIPzyUWo6VpQjV/ScmN98/xzK
v9rRladkwpgEEgXXd8ZWSqi3DZ8cKCBF0NBomZMblo5e50OOliYRV0gRFbTCxB09
PJlTHwpXQuNdEuOiMrsrzGPplmB75BX/d3PB2ZStSlEVjMeMtnio4qEx2tc7iySx
LL7HW4u5I0pVA6xhDxz1l3lqU5KxShKo4oVNtRfwFol6fLsridQlp5KUOHRc09P4
a0q2zlWpF+faMr/A6hOD2ssr53qMwBwXe9g7Cwg85s7yAd0cbT08PaXwXtq/lh5t
kdl2y+95N3aOOuiyGvkS8L9xp2XP0Y6S2W/esO0dGJTeAHleF8QIt3WZSQJYt5Ww
zC6N1EA7pp0PhHx2HBKUeKrpopDTiR/+OyvZrdHp1VMOgtXtHUnu3qdzLYf8LWCc
aAXzQwGfAEWhteb94Jr3S8tWF7hudmxlBGKGKfFXi14mNY2iATfOh+QOZIPIX7wP
sOhj1Fqdn/5bSTC2cl209auvHn4Lf0qkxogemcq8gGpQhtIZeTInR4pZvaa03n4b
2s2CP0MILDiUDzjp13FIBVc4t9U04L1620HzAH0/q4HmuPJ7lnTnDe4Rs6RZPYVr
JvekTu+sGjoPs1A351OzLC+2IRdQxyX5ZpTY1SQriL2obh79NdzHjByOvD0rOMW7
Sy53DPu6p2dOGHi4Tqx4Q+k5hHUodW562ymlxESQL3C9ap9gcdbhKJv7254+IP/b
ELWgLYLxoMqkW9j3lfWMMY8lOWKgQFbd0CsSVvRYYL5gLZkrRIPZhAUwCL7Ztbjp
cdggkiHE18uXkYEMDv3KDBvHwoQJbiPKzoKDK9nHCdSEsKCp1XKZgKKpNVJo9ir4
Amdfa8CvFc3tHdVHor5bJg0c5rLwutXq7otwCIoBJUzGl35C1WRIvggaklY2uGPF
MtfLPRUtoKleMbG0VltfZeFDp4fOXZXe+1g4ONwgiGWNIPVT23ym12yaNC0hoVYC
Lqp/4dQlfiR2EfGaPDfXbzeCocpWYnttrrcZKAgaO9EOVYO/eVM6AiTnhMrDvVpH
3LmJFYmV3HqtBLpgDMR7aZx5rK4wVas0lo9qV7u7UApnYC3SsKL3VCcEwgk5feDP
PEd0gGOQLfgeEcJno0uMy9I5SjvvQx2s3RO/7E0JFCiZqBljkcocrsQDsEjo63lz
XciLRslAsBXGstuOZK8+YBT/CXQly3+d0MLlg3QOL2K3kCEp4a8RES66WIHFCJ6A
tUdCBrOogxc4X4GFdaX797eMMx5VNFGXPl1ntmuQl5OfjPolCBVGCKmnrvj2bPIp
nFrBEgCi0LL7SG9ZAN3O2CUb6XjvYPu4/+9O3+xyYHxO3BZ7E4itOyXy3yqHe5Ds
5EOao1s3r6GBaoqcV91iqmuIgzsI/m8LyBXvpJnd6kfe+01lFmKIXIrswsdHlkGA
aGhjEfKry4CXb8WIj8VXap5ywMBGngeWk3tk83lDt6blJ0oosF7UO9uM1dSyAeuP
LVXjSzUfPY/ThsHd0ELhpNc3eBdbwHK6Bpo4MJpmVqxrBs0h9c1Q9Eg+rRI8PD0L
jK3bvwhTJwRn4hcql7HljW3EqDXT1Ki90utY7WCOQ0/Lu6jNZ5HjD8z4vjmph8oZ
Nvs0CI9W4V741R9PjzBgqLlRc56XpezujrO5Pb4fPPdcdbrY/Cl+YYiGsgZk/fof
QWyuqaz/hS512RVJ0Uatu1d2VkIHTAd64Th+lS6PcNBlq0Ctz1L90byY8iHh3Ifa
sizAkPIzMYm95EbHkmjX6bacy2VkDm36358Gyn6ZyG5Ba8AUjw+EJGJ8MJ1n6+7G
UFqrg1DUD9E+BVd1dXbI5HXA297l73xCYcTjvH/+dVCj3wMnAWzaQVNEvqXRWLhb
o8YSPJjXNIO55x+2SpSsJf2ZgynR150WXAqRJSvP8eFXhKUstmHuaIi/TtvJrTBr
pvgF6CEvYqa/DNyEbk0fqv4pzEZUVEXc94CWNo1q76XXeOKSM886o0AoHL/u4NYs
Qvgp8ZlsOPu4niL1ZLBDZ6SMvN1dNehmFxHApyw9o9EmHhT6n6ako8GEa9nTc6oa
f2YpFkFL1fHekNIN05X1wE5JtbqFijO8PZrPCOKTPjW592BeR09cThwk+e9GEa64
g2xd8lzlVNZ+5rclnU72x0G6PcRqwcXu/KXYefiiZgYj78nzaR9wTn4lgRv3Uavp
X8+KiYAyeKHCJvzc5KcBOOYzL/TqwfdbSma1r+5O6mvogXd832mBe1F0ruT74BIj
cSdYwc0CfRMy79H8o8HQoBiKYMkfk/sEPYcG6Jdyu1WFOgYTmcldxFez94bfDJCR
ng4Q1Qz04CJrUbw1se4Mj94jeJX0B3hR/isYae6njqf/yBrE9ZTd1d8kOqiZmMMe
/mktTtmGwEQuoxdpfV/Rw+jjjTibn5UW95xC1nDSokbG46ivmrOlqBnom/sbaCPC
r+I0N86y9hRs2T2pWO7BR2kfqlI35cLIjfQ1jBq7ZUlqC3bhJMWEgH8YUk4Ple9D
KvlGzFWQGDkFfbxv7QB/aEgXtZfq6AtNIxSld8uOj7a5aA2gC5s/GeG4sFHboyoK
icGuCC5d769A1YnRjjtvBcj8WOJZHn0xMPlZBjeGa2h0G3LBS4ObP7PpUXZ0nf1b
5NbSfb0jJzbuzUcwnQTlesEZCzfpT/ktt8fbR3nyc0M6h8NunBWo7ydtr5Ne7p2p
ytsNCTSZ74hI6DJyMaw3YlPr4fPiQLB62lL8cZcIYMm5xRqpYEReNnCMBPIQ1/PX
Ep/hDigiP/DH188XI1gV3wdYrcmjIkhe/fjyMCXgxY4n+JRkobAs0oFJNG24c+wM
7AM0MpuiXXYr8+YV9cvKARUXMNSz4bxrRlP1hHpJgusGVcSOgDhy16JdnTesmrbA
l7GC2XPc0DPzbExuIXfCsXoi5qlFX4IHJuBQL0/nsTuOSgFRKDd6bG4eiNxv0ZlT
q6KoWgLOgSc9n0CBV2vWLpNpaQdVjY2/fGSvcgIrpGo93/4yuXYOlgev0XZzNBl3
BIJarB2R+4rJqJ9Y7BCkCOY8TXFUcGPpBOHE9swURJh04Fb2v3zYBYEhA30s+/EX
znDRbP2KtDDwalOEfJ7367/HHpSKpLZ7dIkjOUTexgoBSCStWO3TtdhilCOUxRJk
Ww0Wc/9GgVPlDgAuuaeeZv+aycYrxpcEFtSfw/dPCEVDDC8xM/7WEh0DrAthTR7a
HkVwbR881WjpW7AEZLrF93D7gkZ7Plj6ruNOvkYjNsyLUmQWscA+5sRKPJtScd7o
dqMUYl5IMiJIOVf9kxUi6qJOnXFokuPNAdIdwz2OXXpZskbLkhkoX6AHc+ZPYf5g
E3d+9sqw6+1WnF0LS3axB63Wv2/Tfr7AvmBxc/NoScm9XVwRPU3YqXZJ5jN3Q6BL
Me2w0FXoM/6Xw6KHCSm9ZI9iryQz+PcxsYGzdNc2ORgKqYu5dXDAKB63qbkGniOf
3MbSV3jkLlrcdSwD0JsYvuE9v5ZY6oG8RBnFXbIoB22IHesGd3e3X4esEyF6ZoNF
QlKqkvjHiQVjgka0sZMnTD91Zp/wLhL06gF29fkevV2YjsE+asPml/ZUcOZckhBX
I7I9SnJOI+Gdu2fojBvcxygvTs6/18SWhJuzePyarbVDc4GIqARo5EGHle+qKnt+
w/re4kvm0Zdzv055aRN4H8itiRxEUkZb39+oLqnAB1StiqPo5dHQyBneiCU6EAXQ
sxUqdROz2dUUOOFUa5osGghwMhnSo6SPkjLWfxrxckHAfCqNDA57p2BTMlDH5MZt
42RmdNxVVlg5MlYQpjmBGRU3LdtxEi5iGIuTMtAT5JCbj4VHJFPhWJ/bDI32HI4z
LVy1+mVhEIUfMM4ONlQa0S2m58HoIZTqgG8e2ZFzujUVNUuzZEr7eU6Np3gb+slC
Jv20dkrqKYgIIsWrctXUtVEiHAocl0lc8Oo7K8KDTQrOlaPyxN7n4Sk+nNfie0Ih
SEDmyirwMjaAJntYNkhOMD6fujP7r8Gl/ImhS0bv/itTsa4uLewXQcy+eh1TN6rZ
rQ/BIDMcj4XI7+UU23yyxX8CVMn4+YslLLy2LqH6lY8x7fkaEkLdHidF3rR1ll+A
zHKKCI8xl/2UFlqV542miCwSJzNVqXiVTcNEWEmVFUgNCHLMQk969B0gmIOjXPcJ
87LVirjF8D4oqwlDwiFuSSLRhslVQs1OZBsZjQLs8FKx1IiRgOwALDSG/o0aOD1l
/McOD1duK2/N02VVvLmx5KC78/kgDG9palhCupl3W9LC7DZ7ch7DBNq70sQoSAYq
Yn7hQBZhTiVbQad52TCpdOLysC/zMEZAUlHO+X2IrvdI4tmk0FEEAH0WL98UduHZ
EXtSZpz1mdqOra5KEwYZQTH7EhjburmEV0bWYRZjhl1NQ37eojgu/+cvi+/JBns9
iM/zA2kfYLkZ0qiwGUPF8HvdGg7QroZmZKdSaQkqWmuWKCHhK3MseTlvDd8fzDOp
Q+SBcYSFIfh5L4syBHRmT0Xm2PtGLTJ5jclefVUwgk2qngANIdZaa/LeNjGIMtQr
xjL12zmJPtK+NGivHDWJ8DPNRMhhWc+gmCwuOPalI/LgTOVpW7V4HhtbxEtSiOVw
/AO/TIFaDBOTgVBTF8/Yc6PrL61LXDIlBV+tNHuKJlCMnBZ7Y+ys5/+16KFqkvtf
UNZNg8D0LNg2tUHtVXK0SD78Pous0weuefcAfnXKX+tTFT4tpa+G/db0oujj6MCj
LGnYg17l8PZIRDEgIZ/saYnCzbbPco9T/ugOJA67Xv3/x8fqcL0EncuSM5bsbiBa
WicDlyNn+U4nRRvvylFwBJFiHDfMoO3FivqyC5QcGD9Wr5mfkb9qfdZLg83KtcHN
XByg39ZaqWQNeTsiZQYXtxk3D2BgTePCt25cGrJRXGj0zQQhxkhn2xJ6zpYcY1Nj
dWsMUY46fUL6IgNFmTYd/QXTfCHXBubnnXru7Gb4yX8EaQWeeKf2pZ9rbHpEeuqF
rRCzy1YtZgAwqNoQpQurcfjyFep+G3d0JW5Au4YMZ9n19lco3pX8dowLhB/uD8WE
jYv9ihnmI4BIz8s27/0P1j0XJsBYaQNoNmI00iVso3EKjw6DunYaDZJVcFNv+E6R
VFI5LI22B+v8Fwz9pu+o8s5aI8ybK/j/WIg+JNsTChqO7L1rPZWsGjA4EXuOGv2R
C6kFunUrQZhgGH7EftYaPKNulH1cVYy6OVHsJLcZrjVdmBDEhzp28L66SUAs0j5b
qek3T+oljJaNY6yd/UtDQbpVdLat6TSFQt8fD6Pn+sW9oy9H6xUTEpzbnqJqcfoI
yzaDWT0xswV8z9qCuitJj0ePupZNaSnaLp+K1zPOFco5iFQvT1hCW3Q4cHhZrXw/
gi4fNwOKHRmWCZBMhrhUzDLIcSibGlq3L1PR/MMiDebagn7OLCLDNTRNE5Me1W+s
pP0UR0bAkKPICfldMmCG+TWGoAaM3vZuszSbZHLmnS1oJ+1wbqC6saWFyMXdKOo2
kzpL679/6IiyjWaE6c6f2L6rhly7HPayuPlWRKTv69YrSF5GXRtld7YBuEZEKq3M
UBBBKIN7IH7+DypeEmNp2AnL0z8kDD/zkYyY3RCei042HVf1TUiQ1caiaWwjAhat
BtMbzcj7iLs6fpyy5+q641+vLGsPt1p3Yvtum6FCDV9bzkUWgCrzOLyr5zzFOI6O
G3Uk8DzHiT/hqpIOFC93fdU41IjVe68PXsyxfr/b3AMJu1kZqfCzAu00Zrgsox0a
Pb1nZ+yQMhe+WVsF5AH3mBowKi5ThVOzoI1SOfOGMxx/nCCTIdYL/t2RWktt3ykC
+Bk6G5dNGtoCLEQmxcdmEdWpcuvpjRygt1Jk/0I61tYtOKO11rzOdcb1JX+1PJCm
/rQ82JD7UwtqaZQ9XRf2GQF+ETZQcxEHoWvL4Li8lU5Kpw4ISrGlnBK5JfHJLoXC
ri/1JhrADn7/E+1IAeCsnak9Memvt65xEEfjGnfX+jS9JGmy4UxhVIeqQArnWr9h
IYDElKlB4bpMBbQ3X+CYeCoy9H2Wc3oXz4XOnEm2JhVAZYGlKz0jdNSBpbFzSMqO
wS2GnOzx8za61vH27GGqNkvSvbllXc7iSMjJ3Z6BbfVp9rUnpvc5FFV79Q2SQUsb
GWqZKg3bfXSuyoiRMRLZQEyg6pTgXFRKT0gzPATFWK+gf9D87BBawliV5OY+5+eE
+LV/gCU+MLdl30tRPxwxaSs9e7oriGpKGTOpIfkQizybaWHexCYKDIefN/q4umJR
swLiM3OtjyefT+5KQfr8DmL7fVx0aPjTVYbHIerPM60w4wxZr3aNXUcmjW3+PFg7
BY9c1G6HvuB4TDQEtN02HAcNFjGTadc81UoqAu+S5Q0mdAogRzAOTbUTUxphSney
K3d2QPxl3HAMrjmne2mWtvmkL2mnUabE447HFo/a1gGtClQ0Pri5nSeq7A6jV1P/
BaHr2DRYqo5ABhirtSpzMEbt40RpM6IRODtkY3+99bPVw4kq0OgW9rdeK+tkJ3F3
soYpD/2jzLQenB/D/WTAnBKVdAAYhnIBByF6om5WvBfeaylVRU4KiNFDYDgVPxi3
NqV5FFTGuRlsiSt1WpCmHqpwuKaaBo8+l3Q9JEqU6SFkyhPjpHDGjQyp1Djp75HI
HMvuu9mW3oxNiIPZareDxfo2vNiwPj8OCaX5jKNgViJ34l4jveu+tGbvpWy/Zo63
yGEpirGTGH7FBdPvmVGOVIm/w6AuZXOPvAlbaq0nfIgOkw7oR/il7nV9CVXAyuBY
hLMg7bK0BmPxXrUI2iJpwuDZYD+eb/AUjrUONu5Qow8jLoN4FfTdXsDF97LK7XVp
xnVKrTJsA8WMYed8kgx19bPxxuNgjoj5jFwqRCAJiqIy4nA6ZZQevAv2vqMRPLTF
CNjzRVhm2hSYmYFBswNgd+bIbwcKfA2CB2lyn9FMJtkS1TpUUDHpk6MG4wEYWcok
1YACcBjtnYTxc2mWNHtcmZ4kD0mAZXZhN2XFyI27STQVC9vR3I1UlSc5R1naJXFj
FEMGKhl626sNTS4SWw8FMGkzZU+psx3HasQEWo+3FGRux7BJwcLjAryGnWXOkRmJ
HswAEStKA6UC7oU4dJshqw9BcQHlGjqXKfm0dhgv866I/S0WjDZzlxtC5WvQAXv9
Gt/dkXy711Mnmr/Egvtb4AAXYCgvungK6CNH2K713534D31ZJERcXZHm7C9zDLYF
e4OV6txd9cIvrPsD2laKzzEGdmsI80xAbAvrJi8UVozUoU+ho5u2runHsivvmnek
2r1T+MsUDu9ZM0rwxivFv0zbfFGL96OkS4iXAWgGJikJNmCoQzv3nQwkqrmQ3Q9e
aR6w9hB5SNCIOs3XNB7XtmxKRDB330CNGGJdsBMqAXnlSL5n3ftFUFr3nUfMZf30
tdBudWC+IEur5681023nXKRv9luXMwHCWCbUk4ObwRDL/Q34r2qE93bfyFtkGUJj
cjTKAFArvF2BwM0jbeHD62wsKVNEsUTyaWYzK/I+z5ehZ63PNmYW5Ut/tXbRXkGS
VVnQlAqQCzRKzKSuSVfgvcnx/etevi8FyOobvQv7uVcPAsUa4BBFTW4GyJexxayW
CXg1fmdLYjJ90d84S84zxhMPB9ZQ0zDRQQ1Z7irUz59v5asZaozNbO6eQdVz00O9
j9XbySXSkzRlGHE7AD8p+oggKfbTf4bKCJqsFF8hNhOdJMwtzK9fFeWFWDXu8XPX
olOpL6Tg4hVWaZAKttBrNgGFyTdkR640xsEL+w7ksoDYexVHe+BcNMH8zABY0WcV
pLex9yN+2MmEtqZukPf5CCbphn3UktqI1AJCUJqrp5xeanwTyQtItwcsrANT/0Gz
cOyJpODeVbolnIYOfVDX1mdx6HGa3l+B+kfHg3Qkx/y8a8c2OBaYt97RKeehckkf
JIW5E4IR/iEEQm2ABoFd1azEpT+SmmzKZ5z6+vlm2yeABrts05wLwXnIaBG73cdT
3UytPByU9DC1pf9PFBc22xjuyhy06NVhfG7WKs+doI6KS7y5lNe8LzhsEEC9HRJV
/uXmsPkIZmqlJ4WrokY6MfKiC3EpxJ8fBmGZvjoCm8p4pK1GqAYyGiAV/mVvaFyM
qKmkk8JBAqDjOd/7vF5W+QkaowjgxacRoP8E4CqcEIHLW39GQAB3QcdohvC9Swzg
Z7eCmiwxwct3X/k0dO42U4axbgFiyOVBtgI0drpMpUq5xC9hPn7zoRDSf8zLwXN9
MyAMbyBYV42Wv8U1LatptdcjIEa2UQsYvLSytuuwFJlTIbjhfPTF4C77DHrj6BG0
vjNyMa+9KalvyZ9WrLH/PNHgY11lza19wD614IjsaG2wfSA0e+nVcSPHTVL6bm7q
Q4I5YTP1ecSS5X/9X3lUjkxF+2ujJ+A49kSv5jqWiQPQp65D2a/2WByWKRUbu6IR
arWBkndqvFhZZw14lYEiOyEZrWAAooBhsdlhEgsOray0rfKgrzYR/HGh3lQ9H4Pz
yymRIQGz4IM2Dq730Wsz2Q0Iq2/MbuRwU5ReIbLI5fU6+UatgeShkXI/QFZ0bjpi
OggueE3tShQ3Y8PJeKWpAz4tz36X92ZYtq8zvdwAwTEyDXuu/z5C9k1f4ixJKXoe
wVn3aNHZdhq5X141vwGjgoHc7uo172KbrQ4gX8TXsOU7ZI6M4P7KloaOpBG6wg1F
XS9zABueD6u5U1MqAKAvuuQAoJCnrSgt1FeTuaIOkIzrE0MBNUl5vcs2IgZCR92p
oRcUwv5ik8URYSGHIqzHYVvgwfsX0BVpaSrojeuTcyHJABlmZoobLS9K29EHDd6K
Dv7kVyLjZ9aXUcLyxWj+Vi7Ne2SNc/mu/fitKNVWZ6xDGXQ81o2ZXTmdnbWIlLww
tuGqv0NfijkBd1qkAD65iq1GsXHQdzBFCZdyJpLTpnKZA2+pEzzxT6h1dHsb4EWS
DMYtOUZNdqeCENB12QJpyhaaAyHrYW2fAqUMGpdyTsFphC0o9fz94KQ3v741Joas
ZaQomzmj9m18kzM/PfycKrJMSQaRN9E8D8IYgZmGKSkMfH0vBvoUNXwOVl4O/TeO
8s7tgrN+TEy8K1diqWgZDW4nCsvCDjmwNkCyTfKv3/38tWtIMWLqfrwOSA/Auzyh
J6ERf5r3zRIxuhwIqxZ6Iv9w+SVxZkPZQUQcA9HQbzomTKSCa19vDRyHa42tH2/L
DyXksYHy1Y4cig44CQMqGntnWPmOwLsC+ngLxvhFunlq1ISKvIFD0v2zR/ey0Ypd
0MWN+CcbbqDYE0rpD4YGsBZLNZxR7eHz9RA44TkobZmOSeWDJKHfn/HidTl4iXvg
1DUbHeys2Kw9FdVt+GgL411eBiFPtdff4ngbMDrNBHgIthG59sWn+S4JMbFzRazt
jIwq6cuFgRnfX2tiInG4kHvrK0+68mCXY8YHUalfN9izjS+MhM14wU5ibPtqMSPk
kIqUCviJZkbTpLSFtU853i1j0Jn2eKs9iZMcoCfVtkDFhJIigAVYSW5tZxwB4MdQ
c8ZZHjUtZ4iPXTva/uFdExbxHvWfMoy/hGxQr7G465DyXBYno8Y6h+aOtD62YKbv
k5SIQaXQE50towvBUDTFTLStElqnMX/Vnway0FLykWCMkbR1JkiqyaZ8BKhrF7WU
Ww1ioJPB1XiU6g6NJlmBRxOtSl11jPQ7ckJwRHwZuqLBYu4WJWUPsHfzyGay7E+3
2cHaaWJp3hOpRPjRi+8vuJ0VzSgIByThe3AoPWQwGeZ9C2Hc0j0C0+5ni5oEBF5B
ALeY7HB5HYSAxfpK0VpvwNgH2IUW67ZdMwsPlO1K4r1rYzqLnwksbcf+np+6vndN
Qti9M+n3xZ/v3mqMIliAtBXYEyjIlrTKAW/dZApcj2FLtuwixlCqteYJVepe6fKv
5CPqDIpf20V0RuZYjFvQIO5O0+bp2qsSLsUO8KzARweqeIh0850MYtTTukY/voEg
LrqSVhDNBLCnMzVPEtnDskqv2LN9wpvvmXBewdfF03ocrP1FCPoR4hRlAJBQaot7
DgzBHQXmN/Eq/q19SOMJe1KKgqzvNApQ5C6rdWL3daK24nNSNwa/vw3vJth0igaE
6qqKZgpHfI9F7BTc2IlZdmli+2tydbv3fnPZXdb+06S5ulO9yz5wLuWlAyTNVzAe
N0yG7Z7p6PLO5W0YOzW94gisrNGkOq6WJpCp+epROkKMdXRC2ywHPosFfKL7n1B3
DrE7EGst/HdoecrrgFAlFBgtrjZAC21aducZpvQ8cki0WC9Pq75K4AlxwVGfDjT0
tl3oqmmnKy1rRRwBPb7HkBI4tuZyjx3QHfa3F4PERCGQNYl90Qb/UGmeg3fh5iLn
skflOYKEI7vkgpmT+0KgzjB4XYGmcxpaq6BuT1KO8f60MswqHUUsu8DFcH4W7vjv
FersOk6F1eD6qZkAtFsXRtpXzgbaOomvH/U/cGaB83j/sMNgqrzDLaQYA9YGj4pW
U8Kwpfhlf5ZEDohTN7gLTtNvr+SIqju0dUWn56kYeiI6OSdWmmtlWQHLQYRsVD0r
4awLfJxlJ+f2ivNaJrbyD5cie2zwrK5ozfz4kFGOHoxVvihzIRp2hZUAfuO1ZXWa
dgdQnUL1lENUFgrtjTtbM4CW74TSp+/HguWvUIMabdHMI76GIkP0swYnxPsbX0DA
VI1sG5G+E/jADSuMAG3kpvuMJouvV3TsVG2GKGOLcffqDe1dtvaq1wOIVPZ4Z7ng
56TjN0awtkS/TQIBxe+bnUIk7Pgx0Y+G3n/FT+m8aHoaVxbHrHJKDrTBMTC3dlCc
TuQJg4k8DDay6HBgdZZzWHtwBW2qGUuhGAl1dscepepLB7VsraGqQlQ1YojgToMD
LGMTQFS8cAiPrnqJT6Cz5H1/qtZT9l/qnsU3YpD+9Z3nH93CW8l85BC2rfU/mq10
d+6e/hz9B1nKVIqxzM1DP0EXqk9VfhsJl3wkMrriaOW+BAPGTahlDsxnQat/llDR
/5m+ryL/4brbfWksWJRhNb0vxe3TJH+fXQmVf/gYK5OTeJlhvrytLCMg4/rzvPur
t3raQl43TcWz/QfsB6F/YxuM+hsznFOoOtnGHCO+wJ30YKZQly6J6YIqdY3bPOwk
mL2Q3a0TGqbfY/gh4cdk2d6rLXsF9sCiHBQG2phgYAI6KVyHtx7UWm5tPJQHozG9
JntANVTSZ8c3h3gfSpqoXA+2fqpPWgm35IkswNX0Lt9H7Xzm79d/tyo4P7b1IUy9
YgmUHGwC0nvYjDt2045csiIeGojXThrV9gqiWuk8dDTIO1LK60Q3hTbBtPdRM8GS
mdTsL5n6eG7xOvQuo1v5HjvCgjjbvus6IFXHxHNXer/KVKHKP019MgdCjBIEXnsn
HK6K+A09xoTThi8KSf11HcRHpwiQsFa/9kqWezlVFBRhLKYZdFLPl6AlAd6Ua/Z3
qaL8ojV7qviOrJ2dCFYVTQUSuQ2KVevzesIJdrUDVvVd7YjEpOxy8PHqubayTlzo
7wYLX7hV9JOEE0TRxrwzSD3A8Kkya842qo11gpNftXj2eSJunSM0MC1DIayHoujk
cYFbvbiA8WI1glWQRXLqkYgVfK+E5fspqfxBF5lJWH+IRD1Aj2w1Xu2Mr0Dxxhj6
vd5SvqKVS+I2ABDri8MKS98Hquv61onzO0t6MfZHn9Pa2YcCOF7iR8wzJ/k+QpWm
qvAL3FvMo8GJd4fQY8hNESDTg0f8++PmCbMrE7//sanu1cUBpMCX7WyY8Z4Qq/6L
SwNFeV+aCxjf7LdkoBI/aDDpD5tzZgVU9ILSfAJvqPM1gqADgXQe4snK1N1ccCxz
arPW+13HuI7bpzmT7ETslVN5PXwJvGtpFkUTCgBIuLQYGIaNQo9kUHM66L2adR6I
TIhDeduWwXdQfPr+P8tG47yNIE7KsrJb3xA2hbpsiFdNyCcTRlarzCIsI7sXFKbQ
QtIEW79onUFw+JW4nN6XYLvkIUjIr4Su3+bBPaLfLhF3x2ADYaILHrQyf32O9has
UlX/Uht9E+F47GDKJHv0YLoUtzV5aJomXHzmlkavnM74JVo77dyciIj8M0gJYCh5
Rs8kj7i3GS4uh0nxXO35/VdprX4WlwSWVUfIbuGDKtoVV/6LFkYmvDeunmDUSTun
seA//FwFmFptlXcMlaJrzguR8g+qdFM619Jfjx3WaK31YwCj5n+kuFL2TwRpvhbK
72E+3061e2D8wu79xBugECl1JQWRD6kpW7Qm78VMwm8IoR0EXNbtcTDhHSC6XTN7
fj77VljbeSm55pJK2JvVjmL7m0hpesUQJpi3EHvi3aohk9Zqmx6lrv9eOjSSZ5zU
AIy41cw3NSVCqEXHAzemA8KetdrOgsXbMYTycmZQaGt4Xrp0Opelcf9ZDE/qRY39
dZ1CTGBFyH6XlR4/qR1wXGMInWpKAh6d62NTooNY4SXmSTugKCmk72NR3yX+ZU1E
aUBxy5HHoZbN1imRYw9WVaG5qDofZo3V7fjMXFnacVb6GSRRyKG0omvbMo+O40Pp
FeS/ouNeclweiHJ1ZB2Nzw516zxV1jhZpH8WCHQ6gQaj74mF42CRvtDzGo2TQXHD
ike7SeIy7wzSlV+9amvu3/5V1jl/rl3yuEXBeUiE8QilSfTwOtoAK0WBAa/4IH7a
nrJPfORu4T1/YoncBLK97/9oKSV1lxw44G1kHfb7YRl8uONCqIGnArlHJqsUQZyU
YhwIQ5rTRuhxgBvPWM/Ul6gqPo1ZN0j4pl81W2A8OKHrk/ziCTy0RQDkGaP/1Z+h
3ZZXGSeMUVvocuPcO1a9fbqeNOrmb9/MyLhv5GtckYk2Amt6a+B6KVpvdhCl4h8D
nauL1VUTKRpju89O56OKODuvy42gO9Zu80ht3WKX7sCHrZZwGxrVI1Bq4OybrNe7
f6X3X4eiQEefx6ju6Q+6sGSY/Xf8Sv5z5q3IBjNltlG+P+NRnNO+b8e7xaHsXeLg
rHDMJ9kXv5EQOHcW/094T2evxw7hvcrovPMz+/hHKsHmMl62K9uNeau396s4gFb7
3P2AzNuDysxmHYDrU61QwX/e3whYha8SasnyyowuzA1rrxbnoqC2uQKRJoH+54wO
KZZlnGpz4gLzqgHbh0nFaI6f5t2tbXx9MiP+3EBTtVJ5QxMCpicJlrYISmRuKhC5
V/m43WKry7FqrbNjiZyOu/2KgyaAuhZzN+zUVcXp2hQZ0RghOGijOoXEE+kHz4mN
paRqu6fi1oYVGzzE/Vbi1hoMIInLO+l860LurVLTdJC6ZazWYgzjGTdF8zwajuAr
I+sUdy1enW4Pbs/LZi57YSN4INZXoEIvaitXgmtLj16OiXHmwyqaDmQwZ8GSl6lH
nLeJnKLPnkZt0/FL59Ac0G16zDkDStysMsPhSn43Ow5UAJFtzhw7Msubku2iaFRc
HBhhq9DnApzcEoB3I8ZIz3nUv8vp2mnopNhSEe0o0UUC5LZcrC3KigmNBDN2WI06
lu5AUP78hIeekLyoHKxxV4bHenTKtNlGVJlmWpIFv+QTv9N/AKTRUHi+ckI3EixX
3AL685OR/3DlwNi3vJ6aUod/tlhWfwXJNUBP7di8DN6jnjaF3oE5H7NRwoNdJ0cp
YRIyuVvVO3Tge5LeVTDdDetjdsVQKAIdH1xJSwh5tyA6Uas4THXyuCuRMnqgkkc7
v52o3Of9YmOh/Zz1s+ODvXshsM22WmSSW/b4U0Nf5vKJm73bTSpUIICOfv59DVEL
L3FLfjI1rT8Mjm8edo6ebhANmc90Y80Q/eVdzr3RDGYfdf+iNLzztBA1mrHi9zSH
YWKE/4vc6UD+tgf1tikUtrB4IXDkq74UrtKTQLGC0VuyxpOpf1jYl0t0EjYZqDnw
aWIe97bJY/VvZjrDuPOx2ATJXca57I3Vs21wFbQNqhNcVYXm3wRtb38fAguRyDf1
eI7p4aDTY+LMe/kiAm2Iw8TYHV+V7zafp7HciD6kcwdnVr0hZxe4QOY88aoigzHw
YsiiuS0SIYu8mvMt7QkzfBPatBz6amY1LU0NfSZKWAch2TWPh7nE+F5aBN0gbCyz
fdLV94XaXFwvdDqQmlDXB4Ct/D9cZB52N60Esan5A6/C+cH9jcnXV6BG81jtW33M
0WCcRjOIJB1zoRbHtwtfsJDuvcdl5YTAOwZej9kz64c8B+ZARVVRfvYJ0nafEdN4
mdVc1gzntHYyaWc3rwQDnMQb7F1RRIXcheg/2/2mhhN/enPrbZHbInRLF7zNPz5h
9xSPc2iMA3LlXmzK1L8Y1qAcNgdu/Qw/KucIeNPifX5Di2nlRauiy0n6QRCDdtwn
2B3ybM8+mqx4ezW+e+Qonggxzj81r3z9VhpCB9gVAxA8aTtute2UDXsmd/R9pGO+
dsjF8WfjvPZlPu3K+IQVPp1u57TMqCK4KJcr35vXVyipN/alW5PjfDc7jozhvgkj
cDZGrtkHRw7SBfE4n8w0hMyjgBS83bcaVCQtY1ZLb9ZR73Kco9vH7GVKnxHzJP2e
2LankL6xXDk7f3mAbf0NjckRblXBuEBJ78OLgcdlugRX984j9OkkcdPoQRq1JTKR
UPh/qn+WXEHgePBYgYfymYCLmB9yQX9KJsHCLyfqDPrUcmqa/MpxvtVSjOcIk0hO
n2X1jeERD6Q+33m8fu7WC3wVI1f0ZUf50EWz8MEc4MZA4Jh6yG4rr1kr415MEIId
gmfhTbsEsdSNpG0ARv8qWybn9um4ME6hex5kIZB2RIbL1a9H1LeU3AnX0+tTkG1v
WCRMwPs8B1buDi3dTTC7XKLe5ec69XxTKlDcTI9gnuXAl94tn6PPshy9DwZlLeVr
dz4m2Y7raOokSr+aMzHLiKnMtqbKH4iEJ8kuKp0QDbDZsAZkilAE0Q7tlCzKqlv4
eioyp1Mib5OuU3xcXzw+eOOMEBdkZs3OAh4e9ykRbeL/rsxSATTz/91Y3zManQFk
cJWOa38g1xw3MGux99JSQtdfdc8J6osKa2d3IPAfcT0kCeXGd9u8EPXuNhCNwrIx
uRDPdPDVCKWkLzPpnJ45LnxPOtGfLpe6qVNj4KWZm/qTXw898N2WzPmPIdm73h6Y
RmPMzpc2VReiv4nGYERTfJYi423icNCEsSkhZyzHWrl8671b36ijBJ+ZGHbY3XCL
1auCugG5X4w3m0UZ/LW2XXikzdNF0oW71Q/DKn6gcMkYrN6fwn6JzS4jKM+w3hnX
FI5ws7BvZtKNlQuB6RzsEcZVC4H4+3RVKzA2zok8KV1g/y/O7uO3ulU7qvN+DWnR
FvSVeQvPmmfo2P2ijxxR/tcjYCtbLiHRcbcdPEy0tLAZyoN5b2cTW+eay7G8x5pt
iP34p+U0FyCFBlGnDHmbE86mfvnYGziBgTjZWv3aTP8Zk0ZT6atVGPakAP2voBFw
Cp/16MqyK64eGTbHyA4E80gJmVenKhJ/BYFk7Q9gUMs7TK34MQc2Y4jsTdxhUB4V
g4sUSJ91/z9lrQRIJ9KzVRk5a8YTiPKz1kVDA/s/ctjLrmKkUN54ZtJ3r5ANtFYy
s9xn16MCDce2SMt0+1SGJLHXVQdAGfPkjxHAK/xLQH+epQ+/aUDjTraSoH8SEaDs
dS7tAynfgQouU408phDFXujBECsJZm/9NLexAEI63AivlscgOOrJRn76k1DG1Fa3
M7ll15YOitZEE9PRxiBQmQZVDMtoYP6zEDiyVm9wompm3iPwohY1hH2y4g8/rPYR
NDIDTcWn210Z84MQn+mB1j2cljIjBc87kzMth16FZUk6XL1UL5iMEC4caovzoHFF
g/Sq420vGP5TiP1qB9xk5dY6x82pBs18aVDe8EmwAWAeYGYe23t0ymZoIMHSs0mb
QlZYJRIXSHNVHP84SmoXY9Q3H/RvsNTdDFtdnCHDmqv13mkINQ+zG/7PCEFfxEE/
uabaons7vZF64SK2wwMcZsQURXRnWly1TLgr4ol4YbQ5koQ5LLJq7bdUi4fw5vuy
cnLz6rOTMoFw6Hezt0p3HGMpig/bg9glGilAfWMnTHXQceXg+Y3U16KxgFd7PoJb
F3v/ufh7A0JHU33iTwvUvKFl+iy2xJ/SeMvDSfIGjnKDwYJ6QrnHC1a28pWYgsc1
HIRp6KM/M8VxB5Kg7df4443WZMk8bLDxYcPWSthdgfhlOuai/dZitZtfpCN6uM66
PdkN4kS4luv41bxh3DZ203jweYoVd/l0RCHv9jIsEfj0Xpwqmy9lNStT3aF3H1Ps
ACNQQV34xaLWKRjOHC2hytmC+nYrJii51Lj6m/NUcb2lSVLTSSBrgFiG4JHrDb79
6b1Hl7L1qCSinFkOszMqfCs1y8VI+eUT9PZnZf77Pzxdqo88FakVbPpl9+0PsF9G
whQ++takC3LUGRYXENsdVTHJEw9cbScoYVUfJgJ/yVzG1pZl0LLd/2XZ8Sfo4sKe
Qlkfv3kO3NxlPHFMfPDePpH7IwrhsSnj16fWf9QnyPWt54b9J3LZIutmj55r1bMy
zDkP8apHBvmV5glbdHMGqD9XD2l2Fl524Za65PHvCU06D/tWCqTKIDnihzqqjvCQ
C7D9JiIpq6fQuAtwTyjeHgwcBHFyFOfPIxKZXuyDIZLp7vMSmUoix3H6yrxGxpOm
pLyMBb6FXqOPmQXbewkoMlqggE3bnw5wFa0CGtszNmshRqWCSN/zHwGv1Y1wCqsw
7/fxAN7cjaVzkNH4+HKp+2LqggitNjLMzDcLOavLWO5LysLosg/ghqRU5QUmeS/+
Y1o2tL9enK/VCwtOTsupiMqzClt45SNB/Kpg27xTODhFPakIC2Aczz0u8BpPzFbn
6jtXWCNdC/CWnVk4iCStlqW8f8AfzVZmDX8qdLNOoQOCNxE0G9gEIsRZsuBxio31
fBRLk8uLyPSVg6l28F75chuU6i605/LchWOYwiChu+eNHG+EivNkKgpx8w3P/zp1
XiTQwFfDYF+bWKOG0sCwsSY1ZSo7iUTNBMSbNY2WnGDNDY6kzif6iy2n2QX4g4XM
KqnKK5sGkbr1dCfDMvBKzKtBMW9SetqlPA1PY9swF9txy4dZkZXSTIW94o34NGNS
xo6ccpyWaSFuOXBgXd7LteJSxefujMD7sVpeMuRbRehtDrWc89D6I3BjrHosA4ev
V0/T9HhOySs+SxQ9bmBWp67dzMg2Vl60vNNwd40tGYEZDllVJfQIUJJ3xNtRtTeP
5A53ZGzTLjFTIQ7BiWhOwBHZKe9L6gC9xC6Hj/M6y3IRN0xDElC5HNCa1w2K2rGc
fjCh1ymv8BrxBMyYUQTKnGEWngW1kY3OThePzZWCEwJPre3dP48roIT5+2vHE8JF
hpZlh1UN/iHbOQx1aRJlfoxLUMz1lDNby4HTEUolVjKI2OjuBztAHk+Awg5YhmJM
20nwmkcMYtUV80txv1/oXNhLbkd1vKAjujIw8UWxtav0ZGwZZ5zO1K1VZQ6JXBOC
pCmXpoDCpo9UdSf3ErJcUnUFYJdYMBpQpcV5c303K/MeBZlW+mJBFb8YmIFne+Os
AA7BnJvDmWbjLHb25rbxOtn4u6Zdy8C41xwF0Dtv2/o69/D6i9mOKIo4XjwWP/bw
bf4u8Cd292TXAPVhI1GfWzQhfyrBQDOyj9Q5JneJh7/SiumHmL6NbX0q7rMWNK8l
hl4Xi35gG/hP2H0Q8e5LCnBkr++pAaFI3DuW8LSblytZmvpNZmqzqxeOCVAfYhc1
F1xYVs6ohFFD82Yr/P9UqZoJ1SPsE1HW8+SS9McYcP/JNeVD5y7uPtpsvLKyzv/w
5EorgKRRs3T7y1+HZPBJQxYcFRicN/ukBKbE3IcO+tic3VhZ5rCIKeMaBEq5whXQ
lBvUJvgp/rNBKHO+aXZb1/Hp9iOWPJEf8eN+NLeC129fg7PY/Fob5PA8hQ1MNue5
x711kCggBKUD+W88yYYgv7D/zGpxA6b2P8/09FoENdpoiWZFe24F2HbMkjJJB053
hXTzSvS1G+gkQIrRIaxHoxt0xN2p8MyI+NANtGkNDcYGCw82KhHLx9/TDvKHo6ht
u1Ygz1ZxyZHnCC0hZyM+wED5rym6j4fcTfg0e3j6+DmaejEwMAmpxDh7OVQ77GlX
jqIudMplDaE0ov+tHcnGDRL01/Hk+2W0uwuVBOhhAOp46+FScYlw2+tiVMCQYAvW
LyRFMAcg43ivd44C7US2aOdoBjlAZ4EzecW+D2Fz/VWXR7AYfhmNixMaeLhtEOGp
PPRrSHQdd06dyrbpb2qGpH6H3vZbkXWa7IOnYKSnivupX3V92903T1Kwo4F/Da9o
+1kgUJfw7M7ofPvyqHoIe5Yv/JU5bCQi8WInq1OzZ/TD+l3BJ0kSTlDokD+mw4L3
dF8+fGcThc0etfv1ECx26HlkCCs8dv58DHfl9CtLWXbxsb91p3Q+4KYtthZsVa5+
En7Ry8Amx7+a4r1LO9E7ypGH0TVK+FJ7w4H7pk76djUQu+fINhT/jmxXxhRo+m+y
/r6hx4tRQfs/lgexURFxx0g2rML0NX8du8AC7h/0FQzcr7pBbqygVxj4r4XCvlWK
qLHawLcb/wrkRM+kFgUrJkhUvDG6EVg4OpNqttAXKw131Vgmd5rvXU3piEmENA7j
3j3H8mdykOoXJdIzq02Wf0+Lv93ipIZl6aL8ceoKFl0dt5V2kG4cVuSMwry9vZhO
KnYKJImJMKolnwOiB04KqAf7dEn4aUbda1l0DdxhrddlgaWTv02emUvmLVNMuWkj
O/5qo06ksIm2NhVDRIb8+JDRa9fbzyh7fQWkuDNaxU8Td85MGyeNa6/XFOCtJDVk
432H0OgtLYxSWJWkisaIMFR6Ga+P5+gu+hDuuSijYHTq2+4qqiqsPzaV0/348Qts
r1ED8MfsoC8O7fphedR8jdtaz9j9R/9OxUPBBbD7sQlbv4/8Q6S+yAheFtJb6dPX
ZywzGu8uCVghMUT3m5uAzZhrndXgdjQzqcMNsqFrf9SXRXLMjUJArQQDkpagTRcn
EJY/TRrsxhmewfJQLfJD0MFVtqPhQQB4XErXK6jVdXgz87RNk2eWfnOOI9DK56Q9
njl/VfHTAbhDVQnmYCjb63J4QGjt/M89e9TQjn0LAmSz9oQYKWiWMwdLxzCjdQ5k
i7s1WTYr1fOOzvb8mM1h1VZ9z1dVoyPIbljWkxtGrz/aKuMv4AqQoQ1P/WUBQqAz
xcsIImEgPSIAGuD46cMpOP8aSy4ECTWgg/IePI/ZR8RylNTv0Q1/Ar5YO3rXKyGi
Y8hSBdRMQ90FNbTwFaatX8vbj2B96Upp6xfbY4pI1fNX+Uk3xAmci4ry+veFOtk+
aTN8Ac2dQN05pXV6cJeor3cG7gVU7Dxg2sK0vonTYavfRajq+WoCLDkQ0r5RJ5RH
ra0LuJxxcORVma0m2hM3TZ0A4N4Eph3KaQUQcpFVB5XEk4qmP+KMJMjY47sOfflA
g1FEfe2C6wc11iLy11Qo46gilgvtj8lAgLuXbIpfHJO9kArOVhwrWtcRT/IcRNQO
4epx0k7wc3dD+YeIsb1AGgjgnOwptbhPUdM/OOvBLpZqh3pforght4TOHmdm3prc
uCQafuFTwqS2Nct6aZjXjsnibXx8s+2Pw1bliKsukA1QY5FlV4nkUm/BIR64THBl
jEdp55iZ5PpEk+TpPNpYdnsetsLIE7Gw+lrOI3ZLtyzSQaTRCUjfHMEAtuPrEXRv
rnVkXlreCnEx+W7YLiANsoFHW9oIdvgft3Zs3qGthohGy891OPQkwaPPw4NEEHif
QJ7LgSuEFzy4zt6E+Fv32FBakTX3qFA/q+onzQXHg7N8+gAgKhOh6SJO7uyiqOj5
B9vw7leuvqfzwWSAodN+eQl2tsbk7pcqZlNqBxqql6mku1yM3q3RQcNwLWtrHwdY
zcWgVWLxoYI4gy1H+fpB5Hu33MHGJdwGMWsLocd6b0pJrL/uECpMuLEy/Ke6dkcl
LstEswn0RGGIwF9F8D/IUUApFOx/VgOGS9TSmk0WlP5Ht0wbbU/4SgFcZvlnHRQV
LQdJ/QkUOvhOj7/ovoTDE20E+f4Voqoa1XBChccoIQr5RCxs8C2vaH0gbT8ik+ic
HTPzJnU9J7JwQ/HEXe+2bTkJ+SVNxISgLN3JR9calwwgAUcJvIFHL2pZsQtxrr9c
g+heqv67HnIIujmcc4Ni1YCUOAZc5cKOx8OH8zAT86GhTPoWdp/Y1vSFZFFAk9NC
kLHNf1tOsgrWlA0FP3CkPkuvC32zOT78q5VUArgUq65uMRBLMuH+RqKx/V+fhcQR
Oags68dQEGwdemuzYw6A8DbBWMbjv6+dR0ARqF60PF5LvJk+3xR+6Wd1U1OIH01b
mtjOwkGyV1KWiPTnXRgMcdD+6pWX3S7NXPpjyBWkm/avAzhJgAR/prLp4PcnoZf6
Rh/1wRmKC9Q1ZI3BfDskXGnUE2hr93MuGfZ7Q/qExw7fRhv/QlsTEXUZUEMCQpj6
jNlMUYMLnZOJBdnmo+77xLQ1DljSkpCgXW5kiD/S2ufIaDm+zZv13hurRr2KhS9U
GPPN6nWIxMq5f+BE+MwI5nZo3kEfwGO4Db9neA1/hxtqMoovdeRDN6fRgbtbV1zG
6mUrbz2w9ZoXuDkjitS6s0xo7shVhjdxzZP3gxWCsBTR2HCiGIdyzd0Mqiay1JdS
dI32UiHk5DHeAkRAluWzD8VKxrL2MriSsvFeKKTphS9+ouMPq7iX+vMBw4LBp0v9
0HrY54DVOrB2w3mon76pzmOduOAgIySpGDbxdaVt3LD/nJvAAL24t7YLzG7dCEw5
gJge7dvn7iildVDrOZb8Vr5Yx0v4RDqZAyRPWR11UqDjhlTGcTUicvH/3h0h2wIM
pYlVdLIXQohzvPu9wpbUaZEYGrSuBISPK9cd5zzCxhzh0wKpRZMARaU+blL6ZcHm
VrLHO3dH5WN8aItp27wmYaKyF6mDPnjmlXVWcoTK6OSipzZyyzNjNnK0ibl5MujC
dvDHrU/7bWMfO6wnF502i20YHpF5wXZ6s3zSMBHZyubXow5JDOROVtqu8NVzRvYX
qJPqpRVbMlvKZUK+8NlXemQL0E4sqRV9KfI9GssMXSjI6Ga64ZXKTGKAN4+ofVqb
FECXTgp6kDsreu6FHc5uet5Phft7MNhgnCW01Vhk8ANZfjQoYM8MvDHMFc3TP38P
y48LLPsbC9hwWQtuguP7rXoqG4/xzCHo5xVr8yBHm6h5CszajOTUL9ceGjdzP6ns
RVCPiv+H7ieR4OCrK6cJLgGFxll3sfS837CcCo03Z8OSSORYjt/+svap3LHRZLMI
kBGOz1e5+ldQgeHV4C2JSURIV3cS8PHhiIYI7Nj6fMsnZgLdLhzc/DUzEDZWUA5w
bU80gzWVaUdAvhJ4FZeiVfm/1TmSQ59bEhX1x3cXKdaRPGrSRWfnNVCFC2j6nnYQ
a8upcIY61C+JINoKhQ1x0ThEitf0cexz2Da3a8y1FKqcywEAtPG+gJHxVSHKThah
oIs2hFMVTs+a1P0dcJUuHToh6A42lgL8fYVsCiWNvSh6bdoV64D5czCxshzUg1ru
CeM+FwpYdlGA77HrCbCd3KQ1arfEsj3x6IKXppAYLj1CLwu+ThdWF6GtX3VCmsvV
TTRfL+Eny74WMV0hXzEqmASSyE+OuEJaw8DATyWQVG3olJmgsgrCEuBr6CPS57bg
0p4yq/F79U+BVoYlzIfWPKxM7TmbbCAwSNUDjH6kHje3MiKnBXEhems14IomfAwB
EvLhDjsUIkYw5gbQOcvncylvfuVK33uN394YRs32QSg1v7OjDWaMk5oOXyLrv/JN
LtuW5La+9X55YkXyIB7L4c/Uw9mioph2TI9YckRNs4VRS+gV0G92TQZUaEMD2AMn
ifwnIcC8vU5jI875v7Cq32C4eBl6LfLMZP+7vb0dTyA6zgXUEl44qt+MOE/BBvsm
cXAWwRqx/sNbFYFXW1jZWuWpDvS9pRgph11tHWBJ61ussYBChu/5vgiWIcn130mx
qm+HwUKLD+JehiOZZgsexTaZ7KcroXo5EcBgzTgkrN2oZVrMZz2kr/AOH06hVGw9
2nwg2UV5gQo+xAROO1KOCxOd0bpulSmC2oZXD0rq1K/9obBkuWQCbcUnnipeczjQ
ZIzaOkUMom18JOEAQQ6ZxvDdHShCqqT25nSIFc7v9r/VXJVhA2b2uJAUqViZMai9
zS/TFh8/F47k3frhwgj8H62y2iFFcrNxG8xXze9GMeWHTQeiN4muEilV+q+r2/c/
DvfrhuNf3MzI6Fc1IA8Q4oqq/FcRBHY1Dx0R01LNIW5iiLy+H+ykxubliUGiRCWi
xUZk1zezaMVBIP0bMjjD9b24aPHXT6nsKwxhHHsWNNNeCQ9wJ5QQxMEe7e3YppyT
rLflWAYBRWagV4DcOIY5DAZeLhGLp2m3Nr2iPd/ZZkNRpiDBq1bg4ThWdmG/cpAc
NDFHjHxgTIhHbKdJrgNr4o9CXtWzr89odPZ6uN3xjtZ9ciqr0U6+maJjZ3xsGYy7
BDgTq8yZAchFmoCklxRSs1dlhRt5n2NQI/+SInibvcf/Urzd9AHjp9lPiEYaAU5Y
7+kISlX1QNPo+2EM5HpGRYLnI/Yv0zd/s1LX4py0bCmd7w8eidNoP/DIeX7izag2
vOQrMP5wfefSLImiNIWLc1KQ7LctSS+2qI+GBhTB/eJ3K8CmdmWsV/lGArAJfE9/
S93JIpZZUtTsteQ/HTrM1U1DUL+4mnTjYgt/KbA1cQlcd4Nm99EDiwNdHeSQRxze
NN6m2bGAs8Jf8zqTuJxfPrNEMeqbdZ2znoveOiKneZnkEJIyiT6BVSdLM9+j50VY
2qffvmc5tA3NNKEXD5VfBM6ldawDC7vHWumQBvPDDif5KDZs4GSiy3ILXecT14lN
xPtCppbnRy1BGCWiVIkWV7YPMf1ieP5641FLQDqbY1mPOOoF/cDe3X1xk4oE1o0S
NDOPJckRyFUaDbtY38y7c48WxTGRg3R6Q/8fzBBAm0mM4Bp77WrB5yLc6h7S4dhj
xh2yyAscuWVrWIfMBYm++lNncEML/Kctmx/UzOY08RhWnqML0H+Mb6uI9an3ukTg
tEPRtUb2fsTvBnYlph3eV4i+o+7KIQMhGF2SwjrILAmqTn09ePWxshD2ZuTjkLwX
Pd31CUxkVXZazWJFImHjLCEsxClqxBaDpaj3aSAVYlPd0SnbDo0lGZvFFFYH8gQK
YpcsWW33moJQa3GyWGf6ZqQQUFNRbTKhedZiF0t6ZJMLG7FoXf9FAQlYdtsIPnqP
JrnC1sLpRlV5Irr4qPTzP2WkIV2IKbR0/jTWufkuu9KKfkKWzLSLQjj0Jh/SXXPR
2VgJ/7hmOrm/gRtMCDUO81BSaImR+1xqc4aEOG7GjbzppRc9H4Mx5rVKYygfJI7Y
tZ94JD/KNMK353L3M/um07EMFZ56RwzfQGI069/L3CIL2xJTa49APtAwGilaDL/J
OcOsieUSuwtuF8bxNxv5pQ9Epp5riSUn067c9zvSZNIqHNdUy5DRQaYFM2MDQlyP
VEtUQGJ77eWJPna/a6/JAqpub1z63ci11MyAunsNHiqGXVabigl60zt7SbKUi7ZT
AQGmmIWjmABaUdIe/6jOt3guW4PhG75ynNNb+zhhrbSfdAoT605KZifg5ESp+3c1
Zmbw8jjB/uvMA8WkzdEmc5VkXNqLIXqgao6sOnsDGOdSMaoj125l0z4aF8ruSLTn
j8IFQE7+8SEjhbqLThtCWcTlq53+enMw5TmBicQBmWDtV9fahaBXckKiPGrwEDLK
/gwo4uvHH+ohi/ybrMfFwkDzlT+wdSGRKJNc1a0Er3qjCXJwMD0VrQ/GCi9ykpb+
kHz682BAmrJuERR2s7b3BzUU5z5DXpkvG3/6tpPI9X0/7fm3/g3EMbHwLRVHOsOP
iRQ75r4leSXluproXh/HgLyOlJjOzy6rpLuJd5yvwq6jTz/AieET7sCg4yawJsnl
mdB9NsmlbwSUo8qOJNnNzFUJnaKOdwoEZs2zwFo5SKtShuwH8iQPiXdeFsxfL1l0
fUTdkpvd1r3Mz+bxrOBG36+1cDb+XLrbG9MzYm/fo6gYG+sF5qzNwTvg5j9faprk
8O08FtZX3H/j2KGyyYt/9YcGPAzCFhW+ZpzU+QmAYklTHiJhaGBR4mLIMPJTX1kp
fiFRnreOTR9rb4BJHueQcjOLrr/4zaeFofkI5+tb37BjBmTvjAZIPaNG0DoijvQO
UcpCgEEVyD8NNdBgyE7nBuOEpyYiqcVhYOZwKJZBmn2GDdEhEmrkglR7nigUKWDz
JwB/q4aOTqS5DwQel5azXJFadnX2L62GkpcMcX0RTRE9cbgO/HLmtkj1ZNkkSbZb
DttH68QwTG8v17HnBDtWySOZ+BVI3jmA3OiIoNcdAguPSQ/sZjY4AoFBTg/YM0pM
6q1ZMhDEUreL4Sxz3k3JTaXpCwutaoYy/t/i6IColr8awpE5QT/74YNYwDvzagL+
RO/nQ1+qFOTPHKmkz4giXLK6XI4oDxPPYQzFzmf8zkCgqizH8yLDAgKTKij0eeC8
+LDuxAvgWp920vZWAGOJwXXvgOSA17Qepvw+FJDR7+nMuDZ5ZeNZuvSvMXaoWpd5
QR8V+n1WEQGvhA3oRYR/UVN2X2nWLDJOd6dOMAv3Zl/W57CE42H+9mlCwzUBcSbp
A1hdALq3wINtWZXHa3qNzsVvaqfE03RfecnULdbcLPMOB9N8Ew/tcFfxkrHbR3BM
SXWnWgfLwcW5bW8Xch4N/4LwEDX8lzs1fwLYC5JVC9TYIMlOHdXEAgjYIfKzT54g
Yv7+emeXkNwmpQgSUV0R/vy/Fe/KblJQv+ZCumc9xXJ7OEYA3WPO0lOjmMzjQqgx
lmVsmw0imaB34uhmiuhg4PDgGzlhxvks6US2AL4wrCyLTLihZQaez3XEP5giO0pR
He5ANBgAYNWrQzHqI1QN0EltYTSCnn30c8Ch37qA+WsBjyVIQsyENz6j//b4r0gZ
3/XYY/XCEEeP7hPnIJ/yWMk2kW+1u9UfkTteZdl83HUs3+hz6UGPkeXjYBtNaD9s
Cha2Bn6BIxPhOesUgNU1m9FG+vzQ/+yH7CaoW8mgChIi8J9fpgGWCe+ZLW7PGX+8
+ye39/P2hKptnzgK971OV+j7IUluTlf/hC/Jr/CKx27KOSApJO5PXDCN0SXGvJIN
nZcw/7XCH+H26sh2P1ZHturE+bXRxyTtBo0OtBSxg7rU2P8MciIJowLM+wtt2ov5
tDVyrcvxrzRaSniIkb5+HZTfwwqbCTR+phDUecQrguV+Wvf+Zb/wq7nvKH2vGhkT
wOP4rZk3yfVjqH2sPvsuoFrfr7a6mKAYrePs1E+7LN+pJX/Rn7TplKJ4ydTv8xYW
iGb13D7nbv9JJM1mILKDXz2tc6gicZOqCIOW+Z5KL66PgpdMjqrUwZC/Rp3DYAj2
fdof9jsa1jDYa8io1VsAC+aQ/Mdoi2lyZCgXuDwM8lwREp5A1ykM5Sha7rmLYRRb
/QdoAhAWdCrJpkaDDsUzNIfV2n0SaM3RgTVbmq9GQ42TE6hLpNOlorxh+ZMSRcO0
nWCH1QgDxOrUFagwqfPKBa7v8PAn6Iq/9CIJgtRVuWavgZhC5x8A4KlI5KczCK0r
jn6qrwVZBbLUxDbh4ooWw4wqipBF0G++USK2EPbdRSSayDYGEdV1Yqcf0+LBTiyU
Mt7Uln2tyas1qsTadOlhVshy5iVnnyeZI5SFH4BiT/t1BE+hqwrRYtoLMB+q7hAB
pU1dnCQ1ruSFX3QJu+cb0o3LxTFBxHBRj8phQwSXm0B6mQ2F4ck++28DV53qVLgr
VJk9YPRHIjkuwO1AUTpQvNyVXEk93+o5vxcIg1eHyB+PPsliNqpTLAtNWPzO+I4b
EptLyPZbvubGVMobIk2/1WVgOvJLc168fuXr/gaIvkUTCxCehxkvrr1xNN7DHgcd
R7gHLhdk+Lpqa9IVC8GHOaYnkSSlAxRG3Mci8bOzf96BDohXU+qi6f0r6fcQmIsQ
sJqL2FzY7B87ZxoLEf3ORGObmztNEOz04h7Js0YP5Su5xnyf5iM7wvDz8tbBbJLs
qDyBsGs33Xh5r7R3zGEzcmBbcCh3G1MTor34lpUsRJMXH4dCH1t0yjmDYIVBNk32
nY176XAQpC1DjnUOIv/h2bu4nRA7vRIx/Nz0dzd2T3Z76NE2K53wC+4vm9VPMJ0Z
Row3fWSe0vnIucslAFGQio/O1wTJbca1CU6RcjosP1MFNTzv2cwuTwxFBa4YRqNx
agJV7mE4kqj/GPpPBHIL7lFwrS8sLMvM0zSQK2dcEB083MHFR3qDsxbOo1NiY4ZG
uw/oy7MBtWmacVGWKT5XBTTxo6CeiFfaDmcmoCGD+uydSAIDyNJtxgswO/yCSndn
OLl6h9KlukJF4iW4Pd6i9mYVAtXD4ySyVRQFX2obGOVNIdbjHOUdkyiAjuURKWaG
t4RE2HZXaA45jrxjbc4rUh9JrTHtCG9K4sqeTUiSawWnrCl9rpg85tBJU0RiaLSP
K7askWX50Iy4xgh/80G9fYW6YZk5yyeFTNp91aFEWEOcnnnYh951xHQbExwlTOmZ
3Tij+gwjgWOUN7NBbKHpFGoZpPaI8zcapTWWNjKhfpnGcjFS619bBkZ0BGLt6/Wc
kMqE94GEk98LiLsKjcbMnzKgadpx9fvjcWX4LBhWSKTQLddOCjgDXiZyhcT7D9rv
UDwGrwctsDZ5JrJOh2Z1WhD3hnrrJo+b80E13wjo9ggNNrUdA/pX1eoTmT+zdG39
6q0uK+1NNiT79RxE/U+zrQ7YixjXEbBK8NsP0HZGy+ZcDGKBHNaCr0Coy7/DJkND
42r5e4ZLKc2+OkQhZnvGElJmsCKmMOdCxeGBaORZE+WasTjjpXWm+xRup322M9LY
91iCXB1ZDr3z/RTq+bFHn/whXbree5l8OQt2UlrW9EsJBC0WefamI/3zTZ/TdHfA
42tZTzvaMVHvDq+jC/trkmIDA6FIVTWOLplrahAvNyFfVFMSCjoi0OfgjYKPjopD
m/aQss7JyOoyL6KteGLJein6khBLQdki9bx5cKvY1thafuteza0/m87kMpuberrK
vX43iB70jzdr/2edu5VxWqSDcHw6KxsKb8GTq/OZrAaMn+Dt2CdGvWZ9PlYqA5p2
uHfqUwP2frgmkdXx4BbuOAsHGTVD6I4mR2r5skwot2W7+bx/VwIbluzQLghzEEjc
obaIHiFnwfQYNaiqwpEoTlYO2/4hRyg1WTx3odFspaIcqgdiPGHg2OxzyF3CDbIy
JrF4p0Ehm4rDje3TlImYiKa+1a7Bhn+fugVFG9R7bpmeF4r2v9SHFkY5n3NjTCxg
dJ9W2pro/8G4RMSFxKBuwDmkpqH5Fa81qRH0PeEjqWGDWOKuVkbwCBCnciboCeyL
F0zTiNyGrKVhP5krjpfRm4PPntwpl7lnsLoC8YDeEmwcQQNr6ozRynZACIvANfLo
O2keePqI2oDSyUkLWG7tlEog+AB6MCoBt/RkVyBhdndbNCN5jdSProQWfYI6ZrV5
GVgT9gmqfIIIwvl8KBrwIWaMBEDhliSdxX/gLdT5YR6il5yLXHqrgqjpTNjjPftI
TrNkAxWU9vCUWidih/CZ1EB8kGKvUzjcwH/s2gtJAM9S93RL7Kh5AK8JSby+5Fa5
rOdptBXMKx1xeYFFhIv1jjyhqe6MGGbs5Z8fTyCiNpF8RdpNIOVYL/2PqoG5e3E8
nIPST4IXsJf4PBwvPX1DMI+01fFIxMDMy4u7Y1PwxGNWQ7YCuEoYFbdW+sdSFCBf
5PbA9LbUKQbuJNVQ/TObEX+jMypTRkVbVqjqyYOXa2xFusRD652cyPpXhDzgiYDU
ZlzgWGk9qPjth1inxOex+n2yzmlQTRI++e6YykP9L6oq+FZyL1RrhAc7pCaHY9Hw
LI9V94wjqQEfKthL+uE7L/dCehOAPXed9GPAwKn66T4p4MakKBqZmqMPcdjBbYIB
ZGMsRu9JALE1x2PRAwtL3NT5SWy0Y+aG+RsLwgv9zkAYoMtsqThL1aWtBzMuj7js
hg8r+6F726TVclYDaGhbpU/kaCrWDlh8N+14TTdJBt9G1/NVK9RIdL7MihJVNBkh
kPlBfqYSMO4gnyH+sXCO4sx7u9BPFgAFAfk3TqRLQsixxFPb1L4S77mGpkXY9lm0
TsBRBU8meMXw2eW8kg2d85ALV8BTQmrfiGEdLD9cn+q7HVKze5n60LPxbuUNwCai
vWACCEl1femWlEUKrdAJmdj4esldsJQxUEMLMHFPX1kHigNW7mUPdNrBo0zsrXIN
u43UVT+/0vH3TuwN2JchrOnrvaUzsJaB8RezBtL7enqFzOEdHkVQIulDLOWizhsx
mqRrSjVXRsF2yGBLCrB9q8u3PksYm0EZk+5K1/mc5PO/ojBqvH4ggBhi9xApjCsY
UqqXiRN+klPT+wTgjzAtB4DxfDx1LBo7fZn5Yhu420QaSawbqsTfjvlOvolHKWjZ
geyJN6gXAOqXXnAYVlDQEA4MdBY6jDK8l8PvA5mFe6m6StKxow4dB4hs32BeaPGH
bdOAhAGHyuWIDHpO0HtsyVQSYf7RuvO13uMdg1E03IrSlG0yFQhYHwR8q9qjw6B8
L6qbYBwNZ0yUbby9yPeFPTrjklJu4qvDHGtxiwmIqlOGGZ2ivEHiH1PxnZECqkFM
clm0fxpZ384LWGBSKfb4nDRR/7KwITjuxw94DFHUuQZpeYHqFm4yg6akPal6+she
1/W2CV6UVwQClXjIlIh6KAHLQ1fkD2EME3hXN3xpryXzkCIfbAahk/4dKl5oyJCK
FX+pVBEtP4jTSL5kiHM8OCp6t6GmVOpzZ7f7YLeK7i1sDonS89N1GDBpmjLVdpHN
o2xHHZ5lCMfhr9BHeg9x25QE4yeeSGLuWtMdKOrQLbVx4/tW5WwwbaK8x4dKPRnx
C514c8u7Ce6yB8YxhcZLUIqMm1xHFHBGn0bCwmbzrF1JKw2TPjiRoOk4Lh1+rYKz
na+vlG3j2m4iDOC2n5kVa+ad3HatieuwNeJElmEBs7xkaWausjLlU7a42Y4CPzNG
w0FHd/5L1w8vl2OmHl/c31Z5mu6Kk6eLQ03ZKlYLZSC/3pE9ovAs9Wgkb3QAJlw9
9InzbufLKmh49Lcyp8PxB+tdmFdfFyNeteXK9JH3JvDqOvb1PT6uxPaU2H0nk5US
e4xCD1lnhWIOs9a+H2eu8hPKaghPMOi8Phoq0dVfshuCZMjFVQOI3d3xvoaWzz53
crcbf8iZeQi0Qg2RsZWiSATHrBMi/9B9jX8LH4qhiVGwx4ruKiXVaTYwKsrUXWsb
6IhGwNXtaQMgskBnFjq+VkhXo+K/efWq74U47iT63rJ+jR+majGmCmOY040ZiEV3
vpLBcZvOxe1xRgW0oSjZkne1SerlGrkNLBd4s+kOtZEs+0PXH1NzEDITQXsixG4t
2INpudVEDmIl02YJzE+dFJlwErsKKsSbQCZRs4M6c8hhgT2wg0W4ecOUkHbI7wZl
M1nAsH0gTklAnv3QKQZqNtZ0qfwd6OZ3V2oHBTMQk1l0lJL0hv5SLFT9fmQUglVn
yOtfLD2UlPAINdTjD9YSVqeKtOpYHBumKT327f0oGPtcEyc+78DJaGU5XW+bF52w
NQfSphHeTSwqU1gIAsG6GMJTrhlAzTE7WtNpdaYXQj/RiXnww7nCzCpjtZZM0Xgm
zvW8mBAgb7CnTWyD/JIju4E2nJlnQlxPaSWJo8xoYeffFAq/1ctCNT0apbYprUqI
lfAsSZq6boB87+ZCj9P3Yf1OHOhxC9STZWaZQNumy2345ZUTwiBzyw9ewH2cQtbk
CY5ftxuLmqXRnmGYweoiNeG4AmEH9ZmVw2MMWa2auf29RC2/PxdgotTYCGDllMbO
YQfBK3imxGcnAF/VYLhdGAw3MYdnBv99vgRy1+pRGduUTN1JGv3eGjBwYsLUplUb
RLwlpTlNbz9VxXe8ERlVRorC39Fp8d87kRMgNO3LrruV4GgYCYSSi/cy9mdQYDKH
nYuIaEcgpF4nL2hm4TRht/TcG0dLGxYHxqVbx5pv+PrnGi7nn+WQbVMixcgXf+Km
qfRPtKkHPV3E3JxztdnGNagjZ1yxuAi5eJw/4n9euBL7u44Z2nDtXMc41C39hb2u
jXtPpTZfCuu1v9+w1I5lhrjnBW0Jvw9lCFYpbFZ8eD43NQiDBaCNNGDd8gTpfBU5
Ha8HicMyfjTc4+uHpXUA0cnyk8VlcZoWjo8r1xS0bZCc/W9o5EYl8eG+fdHYtpWG
TQX0bakM4MS/JtoAe2dvEwKT4iAL5KucOfltgyHaOgWSe6W4mnW5tNxPNPLu8S42
vExTDfSg5YcmZaViB7MXUxdGVmcxEh7v4Dq5WN3KM+C/QstDmTi7FPfE5uj+hvqf
3VsTgJrdi3bh1qZA/w4qhnFUP35jRYZlIpGJFOxAfGHMYvUbjTVX7I0WBDOTpxrr
b0RDkSgd60kXyu86MKE4aC0cblI7NxccCboyyA9ZlCldaY/eaT5oGcNJS7C77h6/
NwF1Udk+qCQT1ybuYL6punpmd+YajLY/ho8UvNijP73IEGdQfBZgsUnVaVh/uWz2
saY+5Le1/shuJvRNHXfNaXuH0y89ICm8Jv2Rb1KkNuETb8JR3Uea6h3RHyG4npDq
BMgI42gNsoETlbu5KN46EeYjfrr0hnW8qcXKz9phDRmFp5ae60WhGDnTmY/F49VY
BSAweUYxXCUBEXoVYntcH8H5gj1qgoAGZrdwEmRMyozjc6uvGQBAiQosT6BBYrZh
t+ysVswtGEg2yIQ5DXfhqE7XBdwHK+dmrepeEeznphz9Yyep1v/EIwD31+xPA6XA
ksZ3joBnMMaEYMi/f7brpmGaEUQ7UHd3qneGKSnfsoUAJhlOaX2t1egI02jPaKQg
jrVn5CqiO1BfCv0Btk0FvjWjjzo5aLeTiHHsvmcbduSWnfyMkBe54pJRTD73SMoA
ZgiO2ejgqIcPRQksyrVV2dqallnct7X+HrZWm2/Yojy4FybkoEQmv7Ayb786fpvd
8FthBe0A3QU1MdIpPDm36jB9BaIPhD9gIwYDwIfkHVfMbRwM0b7F/+kQQ1S+uJGm
wuQRDEQrKEGOJtrGFsqjr9j5jdmCp0EoxqLpduR6NmMeRFVuPArB5A0zXsKJ1MWp
ftvyZGWbCyoM52uB/iNfWANTvWUN/PW3JbsCb8gDzV1WHFCw7zTD6XS7HmlWHOLG
d7peHy7gLdJ/b0eNzB2kdNBG0PbvIp0aidOv4oQY4S8OXq25mDWZ7ME/xmu7M4B+
F1ONx2F++g+lesMH2PF9E2N+nNr1kUv2l7DNZpozoIPGr3bJ3URYloZRpuz8hgxy
0sU944Gjo3I1QoVBWVfGL7Sr/x/pLYIPhvpmz4xb2yGaQPN6GP9i5cS8iBAhyXOY
dfnYdvn9mJ/UdARjiIEs9cBNZgE9Jza7G5d7dN0oOzVHulclqLgQgKoeztXNTePz
dYE//96a7sceG4oNpVxCnixh2wlvgncK/1gNVK4NFJkpHOYZZku2LJ8QNTNgnndu
yTjWCKtqswyO9j/lLEzFhxJxYOt9HYhn+wQsrRGq8PGokvXdgolU5gCL/2MuZ+zE
kbNIBW+EtUDoCrNJmUaA5fa2HfoDqtDEwVxLF6zwMtlO8vTXD9dxumn4URPoR8Ut
I4xclFBYkN/+OOII2r7K8b+yLZsRNzSNbv6ymxMyKVNeglbye0FZad1c79+djE41
6zM2h5BcTmVfPYiC4783QOrqwEGewhTvPsZLNQMrJK60Q2w74Fpw9fnL/Ewgh2m0
HwQ/9MdtxwyB5okAoGCMvOGxkt1qBkxJpHax6MC58JCKXDWV9us+JG175K/Mwkpx
qJi+3fceFcUDdEBLorwx5UyJntTwKAIqm6AiHYnfP+iQZ+qEYEdFQ5fauOXgscH3
s8ZV73v9uQyFu5xhkGOt5u9zxg0NBQttFAyjqKXxkPFeLf4c+kT0djT1c13oCvjk
b2ZseIw/40uTir0pFCSgMcQFiXXhAripq7YBv3y8w6/k90hHQJMyux4100a1+pB8
tHubHDcZ0jZ86DD1AgeftRGrAt4iNQoH1bAQ37CCTlhiXrZYGkAh/FGLUehMyOv6
9e1NaKN+PHwfM0QnWc9r4qlT5lAVKtuQIwKuKkfOxHITw4ctZ75YCFxj1bqHpCOO
+uf9bHJXDOCiCDcO9rE/19yiVRKa2nqc+bUqhaDJoi8No6G9VIvHqSjBIGTvvB1B
5r9hexsYgBpq7HA4L56BamzrY5m43Z+G9XXypwfiml4xXfhub+C6z+h9TVi1qxvK
mCVD6Jhp4HoAUFJJGdZydISvMdXISiFOjLerZeLIjTOYwHmrUvOwiCOe4NtNN/AS
u+ZhFdFkrVhARL06bXuReQFEyu/jd0RJ+R+BMq1G1nH9lXPngb45TpMioaVBo6dw
x0LgcQlv/Kizq9i616b+ZS2au+L3aA0QNTU43y/wAH+2LvvhDvMLyKPywZOtIzsD
PFW7gstYaBvFUiuAOBOWJ0F+WEOJSvDedhVxTog+3orlRhW/HyFdObygzfIvnIcJ
qIEzE49a5iGiMrg/IpG9Ml3e5SeNH6q1ZBPmWgNM/iTrGkEOWaJQ8f256urboMQB
xIfx8VttcGSvmyl04uTl8FJFNkBRWnv01qmron1E4zAvgn54t7Bl8qy1e+KySC+S
WUJP/1bTIusWdP1S0Z+9QGtzToTvNYVbTykFC4W90lDv9sQ19F+OgP6AvEe/vVo8
zMexaqDxsNeZkGGk9Goeyso/SJFo9eW3aXGLWRIXoQKlv3YNyel9kjBgNuDilaxO
ORSfCKSXeU8cFqLN+mwe6Y8gJunAFaEoeNnY7ArqLewyDfRg4h2xDFIbzGycfzyZ
gYWdezkttvX0bGHHFwy/GKREDyIoHE+dYMCxgE822MhOuOuiS4bbmBdTCWwB8MM0
IhTubL5pETncTe5oV6pdN8SrykCZFaBZjbL3mXocsSfsCasqULstZfsj6MwcOygj
7dQFMYR7fPCgBCJO347vCejkSgZwpBw2utAwQjxKM6FKw3rSv6kJWM2Db97RvYtO
aUX0hh6hCmfMZm8WUKyR4a1asp8kF+lHukpUDw4KOhsOLHK1QdvGjHyl3vLoxk99
rVhr6oLD97UWPDd1/vtGAHLFFeNrhxOTujWuYVJ4pCquTrw13PF1wAIx6ucnfMw9
FafbKM19cSC4AA81uAEkThYYRCffNO4W83sI8b8Dd68sIwTWL3efH9BvGpzLQtuK
TEi87PLFM5xpxKpUVsTfXu0eJiA6J3PgueIJLRwFiJdMxd75+n/M8Wu3Lz7QfUcm
bfwjLS2CDz6CMcU2riW2eXsoQ0Mcbm0FCBD4Icm8iNiJ5vWMYAbjRctIJD1Ia5u9
TaTN7GJ2vI3A12tapVOV94qAAd4hhEudxcj/f9Fko6aFrwik/3Sz9V6SCWuNfQkS
WEbI3Ci60niwb4USm7UxrCvQL00wQbw1d1cOTSbFgZn1Edj3xVkUKM3odEYWSUAj
`protect END_PROTECTED
