`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3cwk+Ard+3oJoxcmMMdPrqMGZVIrkO9lqSE99XQPnWImZ3NyJWuN2zYYS1VzTCuV
RbRI8/R9NGjyT6YjGFz7QPFqkVUEZBPx9kIs51iW76rXa+9FcwlPz7jN83YlxnB7
JWJDV9O1aSB9Ai5KjwgPP/Lum6kNyKhlJ3/0P6y2rMXfk+3287HQJGV0OxvNmKT5
BYkMnThJo9JvzqnxGEWUBHTx7x48JUPIRByzAbOCzwm0juLmNdBay0YuuxhYWDVf
w4xXs/bR4ZazmJDOvQ9wA/UbMmMNY58tMO4oGv0huV54AzSIfYmUGDVenkqf622V
Vk76Cnyi9bmNTkvugIv2P6btfQY6LcMtLw5qExIhrCdKlf2nrs0VvVIROFzZ5dZ2
JHy+xyiVK+oqD7rQZE1ys5Tc+YjGzsD1DAzC1vURBS6u1U+UAk++dS0qzXkcILEg
Za/g7cw2fhlVHlocy5R7OyE6JXYO7mlQJEEYbXHICm6ACELA6CatYO82GLypu546
sEh9f3zUZYwtS0XH81wjPMxXvXz8OTF4DrRoLQOPV+uzZGApk35iPx5VlMDFysoo
tHOgUaPSGQlnsxBH6MEWnPQaaHc8M14o1Dnw3nPmKubFZELI+6CgciIKX2WNqLH6
8+CdRcZpEvDllqyChskp2rRK6cvuBX6Celqix+XWUqzCg2sVwt+yL8a4LAdVOiBI
FNWO+UNEtgrNCuNqILwKFfzs50U8UO4Yu0c9xQujZ0MH9GZHC14JJUxZZ1KyXAUC
Sg+RoQxAUX8pOk8Xr9inPteiSMSBaSAsMd4FNl37FJUIR5EZqt7G17yNpNR68KJb
xyoUuHZ4l4Sv2UeLLgyUchRWEO8Tp2g8HhFHTWQ/BajiTq1MqQSfLBlxqiHBArEP
YiWmd62BxvRDhR7R+CBlfefo7fRTXJMDP9Gq77F1saT3hFQ9CdGlyBUbOiRnZVj5
FqQKDqJmR4hmY7CTMNMIDDCpccr7fg5T9Az560jYmpqQui8VzAWRdr0pwnCp6WBL
ghus8kUcfuwszc5x0d6hKygiOBBybKmQVnWHuAimPc+JlAwbcKYZKtkQd5aYw3LD
8imUoGn7k7DwWKqrvZ57lu8Mhxvlg6HKSBnh4r07yautjXgxZ6/bZ5Os+COu1xRL
W5T9libxhILfRfa+syO5tH/ZBHxYFU2ZqoWCiBWL/d1k77tIeVpXv21P2X3aVkE6
bZaJupUrGk6h4lxqFiooHEaK3gzUbsOD4f/GbNjthnWt12XhbTh0qgN71PlrVLtK
sEJvdJY63lIsZo+rqKAy2vaxItnYb42+7xgCx+NwHxO99QXX+CFKjUk9MJTvxzNV
+lwWh0JXdsDHmWzY30zbuUiLTUeR68cJkF7kHfp5Y36TvescTgstBo+rIzZFTYiW
+BJrg/QFkbT5mmrd3VV3KsZiMzTgc/kyHqpQ9y/HzZr9RLP40ZMdubJrEpSOL4Ps
8+9KsUDOrIhZlmRMOBHfITsbU4ZXz/064Re+hoCjsJ19tGiKeCou1b6Gh/cbGQHm
4jaPgtYE3C46zDGyG72WZJyZc7TV6Qg5oM2VY6cjx/2WDfeeh0G3gH1ivA5Ryamk
TTdG/dbDk5cHLcz3ui7HGr4bxTbVDxCMzGZxO23FMgyAgbkyVCGxHb9rD11+X8Vb
EgzaiBQ8JTGd9YO2p5arthVCfi7c5XdTvBMW7/k1ODHy5OMoBo5x72idvNPi2H+z
QWiOTva+IkSB6u3EOpsoTWtjRn7AWOw09zzoXC+bl7Jax0paCAxWcaqqoaDqK4LU
HodNO0EiyQOv7aQI7pNwEM2SU5QcPH1vK8C1WDidk7Hbde4yWoWfkhln8KjnEUHi
xM29Y6m4eVwbb55OxJoUYFNnQR6bmzRm8h104PX9jEpWqMGYL7aOIXDpksEMG59K
IiVQ2ojsADfFVKwrTossUnS3CH2mMUOx9Xx4xDNn44qb8vB8au7UwLfuZMxCqBmL
VXsakjiGAiodVapKbNFJbBkxbLkMi+y3kZt441GZvqWVbGTHs1VqHP+8ffe8fobY
NS6/R5Na7Ozkm1Q6K6azL2vYzyiPglyxj8UAmWGy80t2xxoEyd95siMRU75Ov9aG
yUH3jAotMZIq91p5z7g/VExy58T+EcDXkROOdgHrEOLcjFxEUjld/DrK9Onkiu3b
N4MHY/Mr/zvdErVptZzrpPII5kQrs2AFLSHAvGS1vp7kEA/RgWmoW0PcXQs9r7nF
WU4paLPy4UAcXjrD35QDKDBn9EeO64S5tNwDGWaUkTj0hpkehOsPQtoFvyjwOYFh
6M9mmboPU4yZZv6hTaXcIB6gYOQszmJ3W9Xa/vNqxjK0s6OJpej6i3uUiUkng7NE
KoONI2zzJ23SqH4PaBPMOZ03VEwcePEhf2safPzXfteaK1sDAAQL3QVsn2RIKpL/
B5yXtbtDP4DPZ+SRDePFP2OIfvOUEmwBVt4fCFY4rtRSEN99vtZsQVNzd/sXsc5N
o+I6T/KEp32L5NG/euAAqWojY52bT3MXNhhGckuQyVRnR/vCSAoKyZRSj0Gc6tDQ
w8NDUlKkQhlJXtmashsxyB6yj/edHz5/vsBk4LJpRGaqmWCDOIF/jT7RYRKFRAnV
Sa8UUxx+HHjLhhbATVRy45ma93sz+5/UVO9WuobgmeqokVuCJ4zkwR+tpQ6VGOUw
P9jOw8yS5KA+5S2nTHK3d7sT81CcfnwRsdMUTP+Ib5mLodQGQEERGHwLgmO866CM
6iQX4RNH3bW8sLH2vPUv/n3GiN0z6Psk0If/02TSyp+Lu4MUsl8LX0V5VXIph8po
BgCvLvcRKg9xWDFMXVCg3ZM4LmlANeP4VAjIfiw8NvYKQZWFJspyoawVHiPwz5YT
oSJ9RkIgwkpAWSrqXTlpTouyRH+/82ptWQsizfB47F3VbVCELLnjAlHgyJ5NAPaC
OAp8z/RiLfrrwdOFZLjogw7iQ67suWoMQf9BhtcQlK6voc6UU6NjChNTCfH4FpOD
ocDZLDELdlGySvX01FeSHCZwQ2IHg1iqWF+15XfbrPMpS+jkZlBzARZuIuJ0Eql2
wiJa8qitd10AI0lSazbhCO4R4qknvAfbtoOZBdMFEwRm01qZsljopOw57XkBmFyG
V5TBTWhD64np+Rnr4paEIB/98e3pzF8LsT1jOag+nfB45nqPaifKubWb9zchi+Xw
/dfsXFM2Rwt61lstUuOI24xd4alx9+VrGGWFNw27ljwq7vgWucS152is6o76T1Al
BdAb30CZWzMzJZRPW/tVrSy5atXdLHNYpQjKfIjysUBGiZ+ZAPhH/PSrBRUjwsNh
qO4O8ar9aZSdnQx6bEonFJafs1V95EOO1fSY7/BWQk4KuKzTLcQFouysTMlALIEt
zPV0SJBlCvUlh2bifL3Fh+j8ABNE6zPYwa1xSA70Z4c3Tm5KZi9tU0RERg1ZJLN8
FOki9PBWSLy+2h6vAwiYxO2/B6uFDPygkcNHYrGx+7X4GmmtIhnMWxRG1sYEaVPh
4sXwDhtymY+Eb5S+0g2fJ6XtTniBe7X/J/n7/KCoctJI3FOMUK4M1Y9KDidFvajJ
y0Uh8TFOvi9COmDQDyNiRFsRmzV6Oh5aPDToQq1rc2kZJKhuq8xoz3v0W+RWUK9v
ksSjJhuGH24gLKO0STF6BR6jEqTqqZBm2p5jJL6ibvLkcADfHDIiQJDTesuGXL9Z
JqfhcNYFQfzoASzEmR0z0nXXrDzvRVZcQCK4RN65puKNlKUTH5wkHcXGFZGxgs2k
i3PwDaIyiXpD5o3L6WBiG5qgCJQiE6WnSkS980yfZnB8bBNQhU3YYztxzNQG6/vh
zLPYZCrkvPP4AG4lbL9bYSxVTclwG+WBd2Shz0pqPVLucZtawmJIy/XhChOQCpJ5
KGxIyN7V6e4kqN3wVRaUSQi5zqg6HDajdv9PDu+tDVdeEwO7Y4HFjnKSMDM6IFZN
ssFrnKHaDtygi03k/5D+dHdD4ZoRRyOBgpXcVeYP9Ory4vLJ7JP09GTqJJZAHMIw
YvIq1jaKnEqhEDFRDkGmMuir+71nK+vFLcvlNsB8Q8RWPZXj9JhXvVSAcsWhZyNv
f55+ikaU+DstRjmsX8NRij1xqNrgbHhUMIV+xYhkbO4MlUedi43XmmzAn62+D4za
f3Pw97zfdg1/lEVx+hWzuP90rEi5n3m7/D8IRmfen22sDGbUgyPPCs+ro2oa2rFU
ndEw+oyfeBvzABUZ//3SU1CULhLQbZse0halQg4JAE2EjH5IfmWPBkghRhHoJPMw
JaxDoCrRNMnC/9WXO/8piq9vGGtaSpMs1gduw8MzrWCjaQ1GrVF5jVpb3y+YZfsE
dWS6oyZXG9+hY1Dl8cDmGSQoTA8KPqkDL0L7DuI/lHdyzw6X6J4YhzGjCCIiGoxW
OWh4YbuVZrzSTv1mYzXY30W241Fl0rvUXarBoHNRM5cjbxiwpkNvZm+l41KN9zU6
zwvYc2gc7q5udyAB5PQflTfGGhLag88+e6185FOy0MVflEQbwh6uWCZLoss35MaB
ZlVyZcLun7y3yN5Z4b33GbONlDBmRGANqwAKiGWr/GJN22Xcg+PPZIeL5h1C3hx3
J/zWoAhX20laKRBOwFDhYMFqMQX6Xt5Tplb51x3Wphah2woSsbO4nxy6jn/BHErL
zdVGlng19h4NNU8C4hF1fiQKGQZ/obHgv7mF5LgRZwmp8io+5j89PDu7BYf4lRSp
MRBz+x2ihpGeA7wXbKexYUto263vwEH0JBVSSCsxIX69u54eBspmFBnG7Ktz+I/9
ELNbCLwlkvGniR2BCrI+rEFb7kRU/cV2cDR/f1IuSVjEjLC2KMKP8txD5/3OC4h+
9ZCnjP04k9OYPvZp33+1vUefMsqwLhhxftitIpKcAib9LavlnRcB9ZdqUjYeLtlV
I4Jgsa+VKRHxvX07h0JMSWHSo3gJdGD1skTeIcT3WAhgP21zgPKUn1Gx//oZ7TDh
O0Lk5dHSKXloHsB6H9aNfr9VXqhws8oWa95D92+kM+LJOzoGWarM6y2tAvfMN3r0
7Sj1jIpeI4nugjqEq0HXfYqjFB3gCNppGUXnk6f6sxrAd9dKwtx1zq06JR6AYVsd
qc6w9anhJCcQ1xTB4MQ/6TvShw+A7BrQRPghBhlkfmKl9iol7OMqTHO0koGBuxy4
tV0yq65vBrbyKYrASGGG9agh6i6bc3gtbPYBJIPMd6HDlfGuGIiQZg556g9gteoM
Si2EO2SFFc/h9/GI22UwcwP4beZGeQU1UxFSHGq3B+syv/YXhDu0swHS+nof8pHP
mf1uDrHYLK9Aq3sr8Vv+ePrKcdIC8dYW6ZnWuiXpOuDUb7hTPd5Ou4vR0PnbkulK
A6Q9QLHOEq8PMhnlsMv0p4XpY5h9t0iPAInjOkmJi1bhSI8aG2jLxhE8ytTdPGft
kMYDbDu9cnTRIbC9uwnbXRiMZCVtWIJ1My+uK7JiO2YAOr+7yXW72OPM10DsQert
blJB+6K+f10e1qTc/LD/twOGTUtsi0WEn140h1q8ZDaPrvpNrOfhXIYNWoGMS3sx
vR1Af0GYOpGKRJHJzn1ia/5NSL3vk5yqWG9FVq9w/qA8ulOUJW9haPHAN9iH2WGS
PFUwv5zefna2LoQVLKT/95v4CpelDON8GxpKYIPvLBl/7HQzdWEcZMrK/k33aJsP
sWWOlslw1OfeoopHkPllAQuJinqpi2LC4hHmtrWRujuiTZW/TTEuqhIbHoBdeZkI
+3z2t2vTdhKtrJ+J3txaUhv4wwmYLawMSbHOUPTS2P4VWsjiMRpGkCPsQ+8aZKgq
+kO4n6z6TpdNMrN5YU1yn7FMFUArytMQwFdFeVL1yO8sE8YRpIG0qBMM39EihKAW
f7jny7vUgF750mXbDgb2fe8gAYWDkhwwf0q8f8HV5nDzlUeN0RrGzO/PvPrRtCSW
pkQ7JIhWCHksEYiB29e7a5ZXJIfaQCqkD4IhMWp4QjTAAJnU2FA6tllgBIDmocf2
VZ4m61oqjqk7y/6W74nGxG72+9H5lai5EFqI5Afj45oJf+d7FnEswGWJTKyJ4ZVq
5FaYGij2PXBQpsPQr8A5TnIRHLTvNLKDY92LFQYksnVesAPZhlii4e6dcLDCoMTT
5awJm8h3NQq/blHPmH7hbGeBgrUVscC+pwFS+6aA3lT3I96OkMM03z+6BO9qpJwL
YiksxBcDLEew61X35wLwAosZbaOEE/jLflJlAv38TMnOVSNdBoLhYGKYiu7TbqDT
yhxuFf3JGaEuDnJ+Z3Sq4s4kSTyJYyEj+ojOvS83jJK5fV7ddvbGydPXzWesA5A7
ldPfIMfQyqUqG9PERXwo8CVg/9FPe6RSo9HItB7XCH05EiNyNTC8mbGyzi6HKkuW
+RSkwOSIiVhICAeCIuIUKfQJycXkjgTvAEbYtQjKvfQPY33ovRj9E1OFX+XCG/rB
qaNTsxJoMvbSzlmhALhm2i6ao68D1s+Sv1jDl5m9WvFNy6ulmJZRCgrJGcy6SjwQ
4VgilmdqRNHtbFa9YXiElaWekrPmesIOVMgUcrl625bF8nQ43j6IRzg1V29IxHM8
kiqRHFZCmNbG6EuYYC2vo5lsG8fz3m08DSTmk/6Aq3NvIq5NnMoq42keW+ODXGVp
X086rKhscZDHwTwga7Q/vcVvFGf7wA1u/aMFyLAaN+3qoyrVYtlgCYldBiaMSxdg
kcz+SMQ1gUT3V4xGuCc0nHXPXDH7NE4pG6ivrPzoYcLqa02WGXBcuZkTFS7wx2lb
WN7ojQemQvUrqfdEXlwtPq8TOAu5cdIeyFBMPX9e+b64HTQ3UAmSIRL94UXzzTzW
g57Nwiit66IYX5C5BR5L13qZUTtbGKbv7cl85Wb1Kh9N6zAprSWNKraccud3ebc3
FATQYzNEBOGtXSWTgiKDYW0LmtR0HJUuquoXeEtwjqloQpWJ6leDBtIkYZG2KBTw
qGLohb0Y5DvEt3ZDNoCWHeqyDKwJn/rHEf78cRNtUVUlxC/96ugr4fjaSLhWuCvC
2TCruMw3Mnkc5233bz9IBTS6B9Ml+SE3aUQaR1ep4LvUBawyoX7X3GBzdrCbuPfC
srQYxcJdQtZm/4M0vEEHigIM3ie5ocU7Dq51QVyGEWgiUGwUwXwmaRpQteEfPerN
DQk6p9iLp7G7d3TWcj13PKqkJnfezqvumEVUUt2PAVnu9YOSMTkpEA47qp5ibOrN
4nFNn8OnF6Yesw7i3JtA0d4rkUDnVed95U9WJq5EOl4VpjUrDApFvFpRr/DrEnFf
qe7heOT8cyQkPu2OsXVeY+yEdBC/DJY+QkryCrhynVz0Hu2sjbTHJvHocuqGptwG
ZNFLbY1o0su17kE73SUXOvaYtkhxLG/fvDVFB2AnP5Oa263bF2A2ZXLIp5KANrRl
rii+mepfl4XfF8mxiDO6/h+6K2tE7N+pS8tHinR35skSHTCEx9PojutN4Z2urseU
3vbj/LnHUHo8TlKVtoc/f6mstq1B5ZoKLg0yDKspXf0UPQok6tmj5WGtNkc++CV+
WnL/kGjuHVPu3CzA/iUPKGUqa+lzKdy7BZa2CNu6LqagG0AwsmflZMRR9/5+swiN
aO5lg0iJSsrk6UD/ZWn7QjFQ4dpgSSAhtAgtxVkvjSyHw3nInI3NaKYLgU8p+Nxb
O7rqz5jU2Y2OvEe+ADlyyizCnyfZcCJ33LXSStMMMSPeiOfEwxJchq8Mk4nK9b8V
sjKtTdU3HBcLYKCMhu4Ne3JqXOB6IAT8Yiboml0dT+O/ShXvpJn8wSJDrV/ejPVs
i2LRpAhxqJF0C8/50zkaX/YPpDc6LrRWntKLN+PPQETu5Xbb9oes/TSsORizcV4m
FfrKtII3Q3jRdGFgrfY+M9QBahFg0CAMOaI34MgyZtKGw+iKGpGoaOboy/07Nofa
GvgtdLepU8isRAW0CwgGd2Pizhe62nUxkQ9Fe9nC26AHlQyfHIAU3YNFJiVBJZDQ
gNSJtN8GBiswGkf6FtQRuI4DM/+rRPSR9c1mFqhPK/ja00Y49ZocjWpsPNueSd3u
7XKI1nXwrCvPYCXQ37LSEzI5OvG85o0bC5W43becppMS3Uq68kz9c9BMIQMWMUTJ
p8moKpI43msPz8jUyCHPKwhP0KoBa6OzFo6ONDMpJtxo0f+E/VgeYn/X87v/fr/M
uIGSkcBtm5AhECYO6CCixWRMdHVHcgncfQEcCgB3Kg3T8K2bBntSOdpB4bfbGpZr
qE+uvSERiTH6caL/TffveBNkyC4IYJv07R3Qvk7eKPHbY1EL928QEFJhZKYpYBiD
E4OP3xQ8LjZyUigSSzRDPl/0dO3zZcQ9gDj7hlgiojkvcckmP2vkYaraqna3JPQi
fuqWbT55DhiCP0C+S3Nty6lBMiBZ4XyeK9mKAnoBjqEpOsqG9CjwQ4EloC/bgSz0
1nXDYxuScsdGBSVq2x8EhAmobwUCOY7AiBmFhAW9MVlOVrTg33LxHKj8dStG+P0t
J8BtedjaazYVyZ87H6/U2H+bxmlky6iXXlSRnBqy0mF0OONwBQmAwzvgbE4iDH08
zEfSDiGma0WAZqTgG4hzv+Bs25+AAgE1D/L8AsaXnIqH26RHv9S7PV+dZT0Un44b
urHrYkZA4D7yv/Oy3yFJqhNGZBn3fBlUR98Xjk4Gdn2llEhA8CPP5UZV7jblarG5
7/1TIuKwzpv0g1Q4yeOEsE2APKBpQQ/P6wFiFAp3ZJXKhlnMHHteOE7FI8olAThd
59SHk8ZwLQx3aFxxqsqZZkQ6xcWacpYhcsmpa0pVqEcKkV47Pa1mo6WOd0BhRnSR
sM+yJVmEpGpp66xXDA0FVIWGkhmSkj+YkBw/zMbrbRWS9Pf2ozFZke1YM96n/hp3
C7uimI2ukZf1PmgHq2tcabtjwBi8mpyKlm07wugU+0VeIiRiJ0LJ0KWY86alJ9as
k51IfimH04gqnMmBMXKk6rTwCBZfRsGLpQ4l3oKuU/aO1iDpTme93DcmR2CZ33Gw
60OO8CuRiwpyJrEa8la879k+vAsTnJbVQL5CEZiQ1rI92gYWZVHfJRD2iTPeD1XY
ft3kc3EeLL/zWtNm07Aapq/7J6QQ1cEkq+3yGEjz4AHOFI1JONb9KTbfxYI4Kwng
q7Xqx2bc+KWqs/Z+LaeK774OyAaL1yRg4tY1/jCBZ753/ImdPP3akjVSRZ/eMDO5
u2hArcOIql/SdDb/TZIkRnvPdVFwyTZHdIo5tgyyjeg0vMjB7/g3B1hmr1Ue/7yJ
nwlc7fPvIDL23lZJRd4o3oPK1J4D7HeMWkXgxsmwfsaaMTx7kHsrVJT7CYeHvnSu
0+tzQp6gnIJC1loHcxYULxA2s3J0dHafK4pJjMEzBm/CWPcQ3+Xd3GTXVQtfiMR0
tHTA53fncm6VOMFQbQZQoTLb5BN+Gjf+wNcL/RbIVt7WFMHSlQYOdJ25QODLAQg7
HwjIHy5nymOjRd06497l0bEwmLPmnJzvFt9N+s1PGEX5OdKYUmbWIB5HGVfd8rhD
eoYmp1vlldISptTXYS+xr253FkA5RQsX8JeAq7vs3ev8TdoeuufrsTTTGTUO6dXI
0GZ4s3GDUzRMHP2uzb0CowCSxsdqTrrP3iVir64zmmP3IrQfLH+yBVnZujncI0SD
+rbN7EACZXXw442lV9zzM+TfOPh+J/pXBgcwgujCCZxCfeYtP+5JtNnPGNTE63+V
RhTGz8SjOqRyjQrVmr6WiLddH19XKNBZHcSuI/i7LK45SNOTObH167Qh8VR0x5X0
ijJAmyWlJ4+XbUuIWNNLtfsF4Sfwlmvhy0M4cNteoEGTuh8tGbsJkbxtTFSRtYx4
K23/PsHZiw5cfU6TUq8i1uHqrsD9uZkqeyYpYzpGkGh/n6ebKvnVPGDO7SGwmJ94
rv5P7e2VHK3FlAFSeRmQNH7CoOJvgVkvJr7xUBM8mm+j8a17e2DeLa8aJ4sZqIaO
wVviai8Rbbn5CHEAYXXYLbxvykyqUsCWc4CPcnm/+BCbI8ovXi8MX2vt5h/yCkY8
LajghjhEopEvuwZqghmrhzHmzoRwIK6dKcOsp1t+u0uuDE8ks4H6DLquPcNoE9Gz
dIKkphOUxVUS/0NOuWavNaL9oxdLOyAJri/vj158x3tPktYIzlP8qHG8Bg1pFJWV
oLBfZ62oCD55oEmlq89Baw+tSs+aY+EQXFYGiH/X/0goLAhvRAKEQIIfiabDCIjz
7vwy3XTZ74uDeo93Pse1yB9lRZurLM0JO7WtQ/S2WbqcyhhtfYVGvKLtviXD4qi1
BmXdgWz+yQ95TIlZLtlhfT/32gPps/71TthzoSrnpZervbgbXnoeIa14BRapSONe
uMX65ayhZ6KKyplWJ6qV4T1P4Mz1I+blosZ9azcSB7KPtcrgin0Tzc82mQLA6wvt
E6WmCkXp/MmCkNIvTXSecBUtO4WFkm8/70mViElm3GQhEo0BbAx0hW1YUw5rgvfi
wYiQZPIcmc4VVRcnYXrXn8uPhAWGkL28M0K3g4lwbeKPGQk+bAUGwc2pzHBW0axE
wAT+xkDnIlCwoRU3UWzGdXcyMjL8AGppzI2SUyoHng2X7ikzKq3ZEq6VnFAnaOu3
DIkVk6hVn+bNWDbv8TS/S2vPlQ6awF++6UqDDLVQA/PCKStWLlwK5u/sBvhe2G1c
mEHbuEcszdKmqlK7w1/f8gI1zUFq+j0mrl2gwmqp/iT5duaMT2P7DeH3k8PKxHQl
bXtG4EQn/bByiWgbZne36Gx+Hvecv8UHxHKA/qZKIEu/2GCsZF4ixLITnDLUe79o
nRjsaWrwdfZtXpyVOm+qTiDR8ZjBGhTsXXatbFKZzq+LUKJL0DufjMgjzMAYhHUI
sZ8V4Jnf2C0AYkLJAvCcuc/B4pOQ02OWGEmEZzXL1jZB+fK2s2HMaWFbopPaWrL3
K3Zxhk2UkGS/nNM5W4oyydu6S4BkYPZRrkHil9e+7JZXLjsIo5Pwwmczq3mEwhng
DNsHmGAidUpX04DCV5DGpQQGzD3SxyIf9HQ6DGXw9H64PrUgT4CmdqciOAkX5zp4
nnAVXxHx1y5jX309hX+bIAd+nhWYI4ghryJZBk5KKxq3gKG8pRM+NTPKqfHFnT9K
bVbWzy2OnkTD10iHB7WVRYw6nT5jjGwPS1XFkUWm2KepaDDokcffxGcFLqwBA6XF
LShQe+sGhuu4n2dr0N/Idj0a4sGQP9abOXyFiURjtwRq3H8z8t4psdgI+9wHlFze
BoPBkKStpGAMUSRU/qsDaZ7rFqmtNVZrnWSlf/Q7ROoM3WY+X32BeT9qgz/b54M6
TH0HEolhi0v+E5of6b6xnPwlU3JQeulHmVetAzseghBULEKl7a4wygUh/NzL/r1U
54112ltehuVqDgj/1sXQ3z3V6TXPw6p1mn412AAHhD7zrpaQBjxQ935hs9FEwWN/
Jb01S5TDMCnv2r7G+oQXtHDRrbZo75lluQMybScokLS9ZQY/8PZ4b4+rEgOnd9QJ
RhjnsRF8wvjtzJXEVS12KBFFedT1vUzTORo2qEeNwOSPOXD+RI7rrN0w2lUUb1/E
MPogfnNUnHtsa7YvmuWzBCUmZMjbHV61dJCQ7y24GEJkDs0UCjOAQfr7a5FXwoDy
Ws/FFlZrV+9EAp+O/coXKkSAv3tHgqNFlFiwcE9yIr6BL5E+5poThVgucb5vWVEO
awHZWgqahyXiWb6aiG7WoOQZfBw4TUDl2shS/wcKYIuIf6dBg0jZJVRG8x55p5qz
WlHzwIaY/7XYb+kmGHSlwYtM4cn91sJd146zqDq+GEIvRhLMenbQjLdu1AZmKJwP
gn+FERtuStiIsZlPICBQb5EqjDpWaQJAaPIO1rXGqVUhDrlWBK+nPncIFcp9Ny3i
+EMg+ZmMEhhEkw5GiDcK2glxhi+JGCPyV/wM3gflACLvEZzB944yDVMTthcg91oA
0TWo3f8lV9FDhJXlhtQpxnOi69VaG447vlgnbquXMmxDjdxSfqwjRu5zP/Q/CWP8
EYP1mSRG4PKcPjggNddtOimZILakaG3SVtZcjPIwS1bPXUFj9r7XVmad21bUwrgB
vEeAP2cwPwhTQdZ/bnDPAbXLsb8UOcVQ67vyDUEcP11FIv+U9FYHYvtxmSU4+g3G
iD3oFzUAJhH6iJccQ1EjfkbeBFJ/cPY1rHaNp9JWKADAPSf1ZqXKLD6nuPW6BO+V
Gbon2tNiL75Sxhge8X+2oDnlYuu+REyeuEJU5GKKNHoMd3rl3cx0cT1uD5nVcg12
jejmZd8SEZ+EbNm/rdtyKFQAQXs2A7guIoM7CSTlaMAHO2WE1/2+oVAe9lhs5FAj
Pv2lGfve/CPvxLN5+/H/Cortvy6BzYiTmhN8rIM3e4aQqWvILb0ODBOKy9GsDxQB
yKcRkhf1uO86JnNqAvv6DMYK9Wr3sXLCanXaCIPqEWfagtZ8L+O3KqZ2aFg9frlw
lJzFtIS55HyMXEdURO1WtU23FGWZkxGzW2CfivjV2uuqydnfvMtDKxjK63aaeBNW
VqvonJAjgk4h8+e92Z9j9+ZZbUylS3C6IywwrBfoAaxRPvku1T7jH5SxAFDKRgxs
xuxfMAHp3HC6MpZtZPsTW35z3uAefRHw+0ducVMn4P+Wykm8ejSfoXBOLTOxTCfo
ZITBd7YEUxenDEvYmBIxcaOCFKoyJKHAA0EQ3s28hyBKGBxoYWByzt6LHKD3O4Ai
VfiReYnnpyF0OaLiAPNny4Jg+svH5sp6tu/9t9ixVGuPW4UXIkhEtHf6VDMy9iOj
JSTeS9bRTmCDXVpfbbdqXqlHv8oCO2u1bTE7N1p6iBswhDqhePaGahF3/KCA1iHY
ZN7UkA8+xgxT03n2jl4v1tDMxRh1AtOLjQSWZNowsu0LlXSrDtSZ5smGziGLvFlv
0F0fvBJZgkyX3dIPJTwl1aacszVxFtqWjabcIUvRxBAf0G0W7ygB2vJ/n3wQtX4z
mP9Ypl/eJrSKj64eddVttR5i14NRyOhThBrxcd3rOufZ/OI3qt5H21X4EbrFcuQh
5BeGKR0yyChAxO9OlvAgDYlsnFM0QCwebXp+ZZN6Xtqhoahz4Pn4ZF6WDgXcHQbR
wWmmuoSM1EBz82zpnw5/QD3ypHGG/IjQgp2Rt+3is3UcYP7i0huV510vs6xpGgoY
ruTswI82y7Y712tO5j0g6Ce9+C+vRKwINgNAXusrXhuw9ePyudbPMakOV3kVHowH
zf9ieiruEe8RVUzXwioYYY6kbBSB18RyXWtC1TfPS8UVqhFReLX9octSNfYSD2xw
RAxy+bm4qgea7fx2Nly5VeyexWDtAd7pEAAcqZj5abVqRp3qOgkqTARz6AW7hoaQ
GIIwFcvpq6nxtZ1dVKrIbhr0NkmIiXO4CKgMREDVocsKtUirSN7nYyYtSgOqpKBv
5N8gF7/NxEHH9h7asEaXGLQ5EIj8klBGFSgeaTnuqpMglCI7oPx0gqlftM2S+h3E
2MamjJ8FdpVlPHIbT74Il5MgziuCExoGnz/pmCkhcEHjPq5o+Bk508vIVvSB/HDc
E1ltjFSYlipSdtPDpmogy2F9B5ZefTpUFM4ZmCjsTae9OWIbr2iwfnhiVKjGERIq
AW7I2o34SGIyZHAEJj1t8SZa91rmPody8C5z++EpKRYhKIeqt18rTXQOhNW07yTw
VvEyzYl/1ei8AEqpknD5PbCs38n6Mr1Ov2PWEJ70DfYUvatuTbMFx9nom1o0P7zB
c8Ys02k24CYPUGaA8sOH473fgERSpixUUTz40uajzVxq4z4G/hOcewm7IFptQgwA
b8SIZahy2yhnzsqgqhQ4eq5CcCNoJNK0iAE4Y0B3qXGR/PIfQp/1sPPuYy0R5FMA
TORzyrA7bRnNH+kzdq5pjCa1tlP651PU8uBn8cccPnwlP8/9CIdMoYQeJebSBL1H
j3oypMOCzkb7DkClrI7BkdjFOFu+yrRu9WKwbfVBnxzwuZvXnnLJpmOewLMeDpgu
o7PNhtHXZ4IEvpYqFRNb0enmAsTH3Aa3E4fKkXiFI2tmgR3hKfiKQ5LudOC5QeS6
UX20kR/PAA4JLfILRB5nDdo0OE2MKZzo0CdvhePPJVIIO0Z0FZTGUFZl4xVTpkQ/
dGE50jPly3YiYO8i6Gs31WNZHNzTfvO042uF4wkLKz3/PJ48qNjGCSiRRr4rJ+JR
NV6nXnJfcrEybIGbeL9YNAW2h87NQbX4FGAvSrHqujDA4+BGrvVQgAXdDqlwErVo
48MiU1RdbxdusF9Og9Bex64KmosfNCBju+E/5yt2mCFFKV2o0zWF0qHm7ZnGO0Fy
8cXPgKNhqNNctldy1TPGpzSvcQ2WHHox+S0vhs52S7/VZQ3Hyf0TNjur795buxkN
qHkw4ysSvPc/t/fsZINek9J2RwB51n2Nuv0gV5bDsMBAo6/ag3/1fCoq3S/PbUcp
oBHWD0Y+QBQ2AQgoLmZ/HcUyf0yUqBv1rHrdSf8hJnvNGuZRVNUaTaoKWz1881RC
XhSFDQY0R9MMD37yFynfuNPlh7AZFmh6vqTBrHhIbC70NElaP8FAy0yKJs/z/iB0
JNZt36ec/gYmpgxVdzEZTh7D3eXu1YbyG9q+uzvs/53ZAZQo+UeUsPayMDA5loCF
mzD1V70x4M9gcmcCbUTyEv5vomB1Xt+W1AmsdjqHDN6aET9mQiFmLTsFfO6Ad9AL
K+uXHQtMMF+BeHttolbaMPps3iNAe2WQvWF4PhS71rGgnsp1EYfvk3gVyYQjz71g
5K6TX5/kAkVi3uQKCpmKgg463qXlvfzo5p3KBqy076abH4GWuLG8nbV9e7ycuFNL
IShtPditp+NEb7tsdn7WYLfPP0tFs4NahzuDB4DkqueJhcuJ+LJdN9pGxFQ4BX+L
HZqdO+ZaLhhO9D24hYI0ragKV4qZb3hlqutPuGmGjPDqcO4Wzld3LubyKiXsZeLa
kOosR41CbbmYC88K1GjDqF9sfSv8WqEoq6GrpN+aDAqxyBczxfHsbtldCPIcQTF0
Tc/J9vv331JvZF6kBAF9R1Evt+sBJm93DRlOasIWHdGJSeQ0f5W1OJdzNqrIGzAM
UjuG23t52QYm+FAudCQx5GpsV8Dr2/mwYj9o+may55PcGhyc562SdcNm0yPIawjl
1QspnOd5De/4P+hGez9xm17AP1mOjgFlsBbOfYf4N6zjCVOcgV1Zc0zYPS1vs2RA
ScX6a4d73yFaHG+TKLXU4Jxq5QXj2a9Yt1TLzAXC8wHyYLcNo/hsnIiUOnTg3BUu
C9JGsJdcbjQFOIctUAwrnbQ1FhQFGn86WcJncodwd+IwCEIyunN44fbWE4sxHnq5
skOCll5Tlb4EGPsaP8qA/l07UFKKAy94GCnOve9B6rZ5o8ZwGAftyYW5WVQUpp9F
i7jkyL8rWTpM8IHNRsils1tMhu6XPd/7QyBAe9xJjW3OIplaPPqex+0+ZLAOZZGU
ARQvjr+SGlws1NUm8kTmf51iMu/eQRkiJJ/QgQMdHXXmR1684fDHCkIhTazWkcQW
HzEgdeByu90NyxCOOExqK5Ep3fnT4STOfKiCrbExUB99EMRYa4DhAhe1AD9cMpA0
K8JmwMibPBxj4ZDWGnBBw1GRqdVA8qZfF8GpK9/TmzeAFw6OWHQ8XmiWYEQDBxeN
aLoE2PuiLTBXxRZprmV2e3U5ricVftkyY+Wi4Uz33A4=
`protect END_PROTECTED
