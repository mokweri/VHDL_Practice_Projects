`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
omQPQfs2JJopCShcXFP6q1YInNV9ot+i7uzO2K52tuMTmtN/qTHSLyjt/tS025nq
3QNmo6uzrQK12TLez9P9BiyFfj8dnolL8qZIho2q8Xe//oaAcjUD1p82aYgohB4q
uEvoUdgdNskLVzJU8s1B2QRUiT2sM5lx/SsrrJp8Tpr3cy4mpXMpZEMuLZnpwrT2
Ak52Xr6J/80kifK4ldKffO/xbgvGE1C9U/di2YatiZ/fMI/M0X2rHi4xz7zE+M6Y
Bkrj2F+vaBUadXdpLD2SSLCRcVJsBre4qSYb83iqpv/eRG3Uk0KsBkiU/Kwmlavy
rjLx3eT+WijNxKtbouQRMzEuGM9yWITnGBULyrrS+ML+VqT63Z8sA9gPXQN1lHqM
srm2hnnlA95pyDPLpwckEsnlehQPLHxWGrtNJeGolYm/GFPHU5iV9suCyChR2WDq
nv5osVOcbwavBMjP8s+Adr8qEz+cw+W6FbiULSB4kfD+w4xi2zkCGdowXGu3MaoE
c3dotE8Y0sD9SEOpt3WdpNFAeu8Famgw1JU8MM/QLvIEgXxYqFlPbHNsvNMHuiz5
rFXh/erzMvYQEz9IjXJNWmFXVl3nIcovF5oXQ7IPcKiCmVw3NmUFOjzlh53o41Qk
bGnlZ/Qmow8wB+OYIxk5yrG5ZQrZltWcenajVieXXiwm+P8I+P6cXcjuplA4NQU2
H/Gvin5PH4EyTn7Y/2+eq/fDYzUmQDVileIu+C2FUWdW/KMXraXmuShhD87hAlfY
Nw+RnvjvBOUb00HTdiX9Cg==
`protect END_PROTECTED
