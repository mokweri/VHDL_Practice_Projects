`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kmKA5FB55Ydto1DBvvSKC0LGT0cTzz5LTtixr8x06RTdFNruljNUNufiP9TfmeKM
WxETbPhHfg5Yl29ReMnbEgSqyNc6mYDTSlfA1B3MqmJx3Nuiufrqd30lGi8mAmJC
Cu86Vr6AfwJI6IuumzXm9F+rQ5y6WssLxMoXJNvw1aj3f5+1uvGoDTFtQcup5upK
3oUNxhDC01OAQRtpCd6r5O2M+V8nsYUN9rBwwFwxORdGLkI0mxG9jiO99Ha8W2r9
FYGh0dAR2Aa+WF9EjcmL3KhtfdWySCwlj7psxb/t24W7ytYMH0kGHIpdkFLe8s0Q
nDUa0iu8zBgkfSweHmHQ0BrR9CVViJr0/Uk6XIly1WMIv/z9foPNy7/Eq+k3E30x
3V0PdM0QSH9hmoudOZy3f6UxUzqhhaibjvAoic8wu2E7R33hWejYghw3rzjeJbgK
7H08LEKWjHgoHQYFwcx2j1qaYMN1yI9YqB/8GaUSGbp166cMQ110evnPZeg+Qtyf
hpOGCuKXLrIEa/Lbj/V47zjR9UpcVlhV6ePFvHeWyFW7XqS+bl6/9gNp/zu9Supn
WvM/w7C9QyIGwfyyvF1ypWfU3c4GYkp7qoELKpHIjZNyqZmXviRQb03ng4oO0Oa+
RlnlGhjg2BxndaAEXf5HHTtar0o+0q+ZeSOBrwbdV+jMAab9uSc1LDTtXNegyD96
1z9seNGNggPkrE6JcWun3kBubrIqBWUGn9QmdQjfrspWWd7vnJA9It5D3KBrkUPa
mWeDq9TYC5h+rsSzIJTJOm1+EbhQcWumi4T/Tg3s/Lwf+LjY4MhYj5pJzuos6VJ3
zKIisG+KevxYCbdkJD/lIBnPCRVqkSaQY168Er6k1+h9r1xB0qtDVZ7z2JjGrnBK
GAHSWWSqEPjIB/h4MGld8uaTIqPqX/OlzwicADuZoWz1AEzj2J/l8yNLQTdg8Gus
mr9JlrReIkZKKiMP+ffkeZuxZi9xt/6j92VP7BnJGa95XU+GTWHdWanuWJjW0vFR
uGT8wrJj1dXPUyMjywJvTiJ3QSMUHcE+YQUTDfJ/n3WRc06DvABTTlEqoX4N6DRZ
nS9ElnesdG/5kwNI3yNQ7O8FES7aP85Z/Ab/+Xz4EzfTvvnGgU4PgFmUQgy8ygSq
Sgsn97xEfuebxPKvqXxFnLGhXd7fvMLUAmqBOIi6LgnnQknWzww+jur8qEg+acUp
XYqWcEenSEcy0227CIvYhy3fK4nQDQAp60OKmS/7/Yj2eimI7n02lBmYetTZa2h+
ERPv5cmH0iD0oMzNuaN0P9x380CC4zeHBIOggkeyUlbX5wQeNupCZgUkSL/CwjqV
bwsG35Acta2k1ohmtRORqj4CoatHt3FLmBLiLPvuOnUeRtklzxSGtg7u/WDFH27m
3k1FOecDiXarnL2lIV462tRMg+X6Amq2XQ73AAmp++wx5oNYbl6QePMd7Co1tdTh
s4gzAVM8MdtH1mZY90CSQapAxgOFU7lOSBKDJr6r5qm86SXsUzcb2aybmndv+uge
WFz/20J51NUplPybOjOAjZc6aJSnq8YsBMzjt6rGK8Bl6itSVN05v6XtsSNQ8gX4
MxxbWmZZq69XscCnBiYsx+7rA49NAgQ34OpideN57KP1PC4P+O2UrLDCeF0whANg
GDDIpblwP5fuwQ6FgCe1BaZp3sDxsaVKXMR41U3yzwEEUZK4vCOK5lYHfswZRY+T
OuNwLRAyy2rXY2mMF9pQZ0Zjv68kTBdfkSJkyg2iZjasybzZmgs01w1kY8TZnnNI
hocFuksoiG13i1P7S2QOKtXVsvRfTHFaEp1p6z2Gs1KjKdzUYK4aD6JQO68lkJBy
boRWvP90kv5uCa7zjdfhLDQPGTEtpPBaPcJDBheBoN6gfqaf1zaTkrphXSNJCIGN
Przda9dJZShB60y0w5DbWWcUBR27ew23/cUfDNE5i1Aq2tPTkDZ/OKwAvl9PDUPW
Xvh13mzvgN6/UC3MdDruBqJVY+vz9erEBlPWyM9QnrSFNOgxmCFG/jOSkgVpNXds
nZOqD9go7rYZihQwRoIbncJGDn/00OhOUwz5oa3LoFmja7PZRckIq9zPHKw7MC6L
4TVTA8vjJUOYRgRH9nO5DejwaSofxYwaRZWV7ULb8oSn46Bkcs5uLs1dBrZIUoLz
AlCtVm1cFEicuA6CESVNcfLa8BYnMCHtETGjiykOAR54xB4cT/fEljEXxtfSB4dR
ElFXimyMHDoeyeiv/BHa7hiVGPL0mIlSfIAAt2EgebxA2eYk3doLR1aS1b8yCHrK
120L4TyOvyHuUOT08WEWgmv0Z8BBZSTcNcFmEigjIYs7IXHLbDkxtBiiTYm7xViR
Bd22Jwx7JyepWOJXnq5VmDIaRtskHSh+ZbB6tIuWgMYrzr40RlAR+eYcuY4l9c2L
Uu3qFOqm/rZCaD09lSTyJvfp30lfbcwHsKPSuOxZ70NDtcp+YIFpczd9gderM1jT
90wvXCbZsgpDI8Vlxpuju1E0TzMhJ1sZvo2hZ6zMZIQhScVHxQubjIm44y0fiQSw
U+IMwVGNJWMGBcC9Jvjn696oHejRaxP/8N3T3T6jzTARiZFB29/vHN4E+ZC7NIZF
Hlcvz0/vtHf4T9WfRe2L5916GPLWKM0YEpeEoO0DdQRgNksZX+dCuoHCZNAUA2Uz
afkE1HUZ1cxINVQSp0WbSe3AK+5QuVUSDhbui4spHC331h0YsrFh9m4VcpnSMOj+
FIu0hbvtAD+bVOkwr1Fn2BT5LRpgmXT1QMuwLH5Q4/GkQRI/mXRbTt++ZAuoelBj
zMDQ/nqrFwC7hXcXkPW81cba14L7ryIq2/8im9GfzDfz+PgYLNROIhaM9CCpTcvW
tmLImM+wJ3flYJld4I1/LjNeEv2cLl+9kbkV8/aZsh7wHEU/q81cQp9yV12iglsS
2oxqzGOrVlTLdxhwoyBGA04241WclFRPxoUFoNbg81uuK13yoviAk1tvllgPoOyP
uSM0vgOcBTmlO2LTHX08KQHY0t2j4q67lazDMZ5Vi660T6opJqO1FRvoH7lqA9GM
o2X6moJxBjE78TAfmeooZ/XT1OdO8kV5hYlZ95gbIeXJ3Jjb+lP9XDKCGhWxAHIT
Oxc+oBr+7t5dtPuCcBrcKsV5QH5VLd+C4JYeCDvtfFqTJ8lwqzEE8Myw3F8TKyIu
JlBYQ2TqauszFQWfXb3vWhKz41XIkgRoKwFmvHLRhDZy1pxP0NpmaFa205wCccyc
WDF/jl565S1cWcZal/5RyjW4rS6/XxAemxuLRJWJWYQb+MjRFzJydW+AXJsK6pKB
74T8yQCOGyTihOl37iy3NhqeIOAQUAl9Co4xci5evXwpUilhePONAumC6m5GmsQb
qSdw+JursUDYyqbDl8j49f9NIz4cDhX35I1YRdUXZzISkgtv+Qnq3aFmBWpSdpG3
qICyiYsBUUU0XQDldsDWduVGNtF6gUvFVccVBnfFxKBWxmU8arx1efjmrPr3C9Dg
H3SPe0qRnjTT8CMoZUJnjJKHHUFIQEXhqv9pPmZHn7nCgLxZeqXM//zm2G91tQTt
7UR3smasi4/7VDoTjK13V6vMUqwnCxafs1E7rLuBEn0aml5prTV2JbVGzEC70iTQ
F3PgWz5b0sAS0w69coyIrajtvOHrMqmsvj3lz77EBq+B+W+h8rws+lewObSHAXV9
krc8ZTckSQ2It+V4dMfpYhujyiYdXNDU3pblc5YYMqJEPzdnaXYtIsYWxP9Et8GF
6K7UpFChD2IGd6KiOf0qfkp8Ksx/hTxkkADFkT7FiD6wQjUE+TzXWw/xYbBuXHTW
0/pYeNCJWAWmXsTfBSSe9gWu6kHxVhsTtbdo9SxMfZMvlNFJRDBjUYlGySE6vmQP
x8JfUcjV3FrVndFyjNf9YyLlHXNT+BMFSNMq1UsK+ZK6PI1//qus+IsluKL6hUyl
UHVPRqY63ZylZrafcr+WVZR0zAIxLylgQgmCeqRch2BGmxpMxbPwu7PPMfCYVkjr
9U6EaknZawEa8irUAbUIr50n5tlWTHyhH6qRpogRE00I/dGaVp3tldpEcUxuTJ68
uO3gYEfpgbVkHf2yCsdJ4TAE8cUHUpZBRi61G0UsDGSov9y13OC4QOb92WPluHOk
+EtXnFHOr8+/zuVa/TOycw8rqN9S9iSXrb0cmiWOdgTxM/o2fAChYeEKr1GqoFio
X6lf5lUwvJnwJ+1vJ3kEBz4utqQOMUoJFu3RzHmP+klFxVaj48ie70fLCm0N3sDD
0xeRndewpfHi43oC9uPQufsF420LuMLxpTkcsQ8GAhvjJpnckSNFZ9UxQzIOwaGI
cCzz1+W/VFMRiZ3Nu4cH/fRbq0wBkrAEqPCMADR+LecSeZX/EjUI3tNJ9F6lMkRL
30gLb5B+fcSqS/ndq6mbhwMt152+/WrnI9jZxz0N1mM=
`protect END_PROTECTED
