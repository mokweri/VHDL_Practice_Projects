`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g11S2dUg+Fpv0ZhJ9XJJNAWqwp6C4vTgvMCWG8iUNAyGs302hmucvGhO5sKQQc/Y
I+jGk8gMZ1J/1CO0YLSiZ7kyrMmaoZEOhIy/bU6jnD9nQqtsL5MQ+tlESAj+zb7A
Ih8GQ+3s9GaGdhKoElyXzDMMY+LyxKZ2rkdroqkpZHk22Yy0BhfdBBFPEjV5cafv
d4FYxfxsnedMzd7B8ZGqHKZvlM9+CcnfgHHzzJgpcfWvTyo/xEpYdN4yG+F25uvq
mn2ca6IDwjNWMYWnUsZIhcYGGqIOrnIVW41qsOLJr3zQtV5af/5dNrpG/Qf4WNVu
1gAKzOrC0RSE+KJvv6KZZ6NCl9HjYOK0xnsRMHHxETV4ImlRnb0G+bJludovDLAQ
TSk0v0k7s54gLZspLRQuShHYa5caKsrwm6udMtk2xfIrq8b7pdTINbNbGV2iWBtt
iDQJn3BhFlHRjFHEnIR0m3Jo1hoS4gS+0TNwyaIhVz3UhvVZBDlaNMf+IK2TWHhU
F9Gki/fyp6uwxQ9Vh+Jg3ApWpBgVYLOyG/gF8mVo0Z3H6JYduqKtX1F8TOtldS8X
Y+2jNbiMKaTHhyjX3cVIhJIAjXi7vy0sJKGs2IOjaQJPH88zI30rcvn1p0BD60VB
B0vu5hjKNhzmlrFzN4MbmJRbjkgFjkMrsX0sEgfutTZ+Puku8Fa2NMieaWMTh8yI
iwewQiaOhGiQlHQyVC/KUD2Poe0zv70bXnWM/YOu9og15+wvBGXn/O/YhD+cMnvu
YqxZAPPyhMLwP2gCWZ4tVAmH5eeUrOjbEf9ovgAH6+oHig5mS2oJMxR1r1aSKWXd
u5TCDhlgRQgmHYTbVhE5DZdFgKuGz3GEOmnIA2kca9nloU1Sbhv8ayjnB/T8hn4y
HAX83dHuU+c+hkw7lZnu+bEH8IbKr9eZ1wqc5vJ+ITSJa8FTu6rNOB+HKzu2Fms/
Il/53KVQ2TOo0NMKB4xRuYEcaJyB4o1KRkVf0VgXps8NTr5SQjR2fOG5Um6JjdY4
U+XbZE1m+lUpLUzabbKJDubPKkdMErmBnR2CCQFZoz7CIa8a1S6nw+2DiMBsD7cU
GhEGRjOAMP/KqdCYz6kWZlKkMnUKTsIiDP6IDqF3PEG+x1+yx64Cw1ze/7gdaorp
MrbCO9D+ZQXyHJyXECH8gmfEBFqTwVP0Sk1N/rfoEQ1fslft3nIVF8juUg7XWRJb
zlFj99RgFQ1ouBw3fwX3W5tQ8RSjM4N/0yfF3Md6d7EV1E+ZFYI3dE4mhZU2vkwC
h23RbuoJaFuvMVAv4ndicHJ+UwEB61l/l8ssIyRASDoSik+3QjAEKF7Ik7cCSnWp
qh7foDLqv4/i1Co0Zk/Qb0dbQaePORMP3i2koB4V2/KQF2uSNmLM94S2z85a9gu9
3WBGSBGD7+MyY5Aes2SiUkfkCWXgjeaQn0G5wXgiNthJToHHNuph97+GKVO53cKe
aCUQ2O2uWqlPdjvr3RaehOy/Yl5MvB4y/ahkJDxlCPVdmJtN+rczbkZGWRlEkjoV
XU3wuxeOXVTcKdmsRFtLDM3YYhqPnBEhlwT3Remc8Kid84kUC6duW8GhHUZJjOJj
XJLS1ylbVYDXAWsvl3cV/AMeJKtUpIKhAHSOSLUD13tAaCGhtEHFpdVhax67JjhL
2tA3gKg+9erchvybeoPzfJTI58IbojiOuqsgBXMcerdj3qHpDIo2T06r3E9bmOvq
fsuvhHt0g/A+NpTb7ebwNyu0vJcX2EfyXIxMlqx9mMwjO3aW4WLrj8jBkakwnWYF
bmS6a1Z1vyvrTSsxxJxII0AkoX+4z/KJnaTfyXsTc5rxnfAWTXzdpDi6plLWrGzN
AbmCQuA6VpfjPQ4MXu4V9OdclzYcUk1clQsbpNwGSZq6xAPoHUDzaZfns9Kd/EZu
GTpGbFQT7g2OPUyVmOweVBRfJPVibs9y4dq9Lq6c3GnsZEiR5yvA4+xM9iQaMbgq
zZw5tC6cYVpz7yAbfQpzTUP6E4ZAUTQ+CKvzkVRoj+jJXfhdx/2+HHQ80BFVTVpC
u2tPEf2PD5OParPwohOWDY8a5rwDka74919hOpXsfYtgj7TqdKxySf/ifOmJEinE
AjuHWty91kjCPAj04XS1EN2nfoha3J1Hb/7bPzcnIxDpKoNSAgQnHhaIxHOfTX3g
mRYVXuSg64k+QpuG68E4fRpupDMZEzzeL3nosvAvcpkr04eGjiS9wYYFGXUH5gD4
4wIr+a4u72eqzyoqEeZS5SJ+OVCldan65A2Vbw7qx5zpHZCT243V1RcV1vrL8GY0
LF2eILmk6T7cMMjP/1g3TECXVuoho7HxZ5cfW3Wqmod5ubQE5mpkbhbxZpGxC/qT
`protect END_PROTECTED
