`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N5cCL1A0pzhQX0oMj/4jDvmhJ77FSgfJ91lXottQorLYVe/uT8fWVRkT9CqFF6kF
3saswOLs3xyaJXSYzSFVI613SSdTyLLY7kV4aaqGT2qazwetN8Rh2gxECAOoQYdJ
+hzkEmRhNZ/CYpTexh3+ERvvzh3QUV7uPt07D+CwNVCKHjSnltHBlMsvuPyZpXDU
iEKL+sSeLD5XBXZ9Kg1ETVqNcTQ65caHRrd0gBqSMZna0Z+fWEXb+PUdS2AZhhlj
m7IFYvwoRcobX7Ve3T2ZHUHZ7Ig9MP3uodRJBUyCwQIcEmg0XO3hEd75ZaLWydPi
uM6QCEP4LVRB9uwpbkgx6NMFA5jtZGEPsEe3iUpqby4qTXr/nVz++b/PBwEHNKJi
7iw6Phf4+pj2b0/iRvZ/YXIMyPSQV1YwXUzm18saYtN6fzxw2jcTd7Og7+OQCGGi
gWO5QRZ7qKo/g5E+F12j17qV5EjH/6OFw8E9A79mAEUSPbV9IwvQMTKNIemcHZdC
tu1c145ulj21Eun2aPT+7lecvj5nYzCAuh/8pdONaxZDWyaBmbzsh35X1WCiiCLH
7cXzJ3eAzN7VoLo6YzaNbRhOvEFG8/MZo/qQYj/yft7nJon9Y0njVTDpB7moSm4B
YhSGBUSuuSYxSqFSDfLqmpbSeS88vzMQKZHlZ12QR27P0yzS5JEs2Y2ZioL6v1zM
tdHrq2d4XChBrrquirBXUZuASPitw/KT2afdMf5SPAWo6LJsLq8Voo8US9wrQx7J
qr2jxzkq8LzOXNwkR6so5zWcRerRGwlAChZcjRaU7S72tXIV/v/ilvkwrUbzMOyP
NEQPnxLxW5dE5IMhbYAAwTaymzV8VryPLEsLzvHzfUf/TjqO7pMZUnZ71pp8tsI6
6VBtxfxdfoIzAlh7eTYnOigeO89v198B4le1mh14Q1tiCSmtgIAgZnVKns1aLVOy
DwlyvjHCnwKnIi6KdpPhvTYVUa6JsyiJMpvWXzzzHg9SsFCSC66+y20Q/9Ur6LRW
rzccLtseS+1gRyQSpyJaScQ6ZqMLRCesXNKQtcjamYXncpllngmp5t9kWHRvFw10
`protect END_PROTECTED
