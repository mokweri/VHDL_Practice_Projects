`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rNEsvaOCr0/rKS7LlLDUEtjhLZssfXNDXwcccMBQuzV4K7IOcWGHBEJl8ruIeXUA
mE4hhqVJFRNq/xJ3L9GuEUjm5eKMNBenPJPf+CO0dMWMXVgrMqYf4iX6GUSVCrUB
6+spRagb83RA7Ws3JrDgHW0/AcR4XE6ZMXO+h+O7Niw2HG4RBeYB5rTi4vQEJYsh
c2tbB112v5OxP99Uvv83qIDIiXC9bqVMhxmUpFUG+91rOltMpXBU4t3UHjKxfq0d
CK6KOdhXeB0kIelfloD+DnrjPnpQkKea5YtHiFyrGDI4U0b61xZeETHUBRAROkBj
t1yVps+grp6kXx3DQwfxKiYCO/TVJo5Ta7okaxAhf7vQ014BxEe20SZ/+rRGnO3Y
kc/FZE7qETCD72IM3UjhDjcQqR0HPfwzsXh+L4jMdOu7yxJRtHo22/xHPCWT4cEm
+vlCwgBKdQckhtZvJu8a/+kmtR9aIaY/4gs9iYVCHW8=
`protect END_PROTECTED
