`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbVkTNA539l77mWIyQtvUx9dx5Z5VaUg/0mALGwoUZChIK1izHG6GWtoCOKrxCh3
V/Gmo/DuysuaZ4Q9xtjryo1mhLiJAUsqV+Tt51dRlauPHI6uq67QWNOtCjp3Vt2v
qggit/KEtiqxnB8WPaxq7pntGQdQDUWGAjCVYQqGebmMjVZhKCauyz4ebqWJlNJk
OVqEi83nmrwJOctmNeqmuWW3y7X6kSAqLV48zHbUYkvIibr7hfFzVLs8TLtVwmKp
8UHNnrM62U/S9B/SheCz9CZd4oUq1g66I3fOPTtRsXFar+tRbsGp0HImCYQMtud9
1xk7c8+ylHYGYTiCxQR3IXk4SDSWGyPloC5PvQfev5tk90mZJhW9MttBJo1TSp1v
xPbNv4r9ucODrtEvdJr0BuhyXPjOlNt+mKXSQ6Q7eFSQIikm4lZxtAEoNHAMMaVT
PbRb1Isx+76RNhwb8INwh9zPsmRr3ws0enzNbrYRT1UVLZ0pzRtjutioFkAh8eig
PXrzNaQ+AbTRDLa8PbphLe1FdEB1JgE9dlqQOjnPyFDTVldiA83y7JX4IN5IL1tG
xyCKIyajL39m30vDuacuDz3HqpU1tPI5vHyFrlOj8DouM0MDCMvDkHDJIIYR5V1U
0QmPtvs9RJDhfQhxt30KtnVp8+agGk0J9/Mz5VMe4CFo7J/X4Rk3giSRzFV8v1Zo
GZibSOf9Olnp+pWsa59aYm+1WlJwv6lgHKlFiCcnJciPh+CdqzGegGgbWrAHFX+t
/LNKD5CAasU9jJzUBj5WzdOdwKQG7YNQuU5HRRRaNnSrWlyE0Zcb4VAYN/SrK49k
rKoERSoJK8MtoYjq92D2iBlvlm5o8qmHjiy3q4Izkof6X9rH0IluLydczF0zDR5g
UwQVd8vRV5/E1Bb2KWyw6uB+Ev8HwcTR4eqhKrPkd95XB39pOAy8yRhi53qjnw0t
6cZs4pEC/AypkMKBYvgQEVtoUTkhDTKDPgzROWEDn38IXyfmVFRIAn1s0PTwdMCl
bvyOlo4EExEcV0FgQTDvQZspRehovYcMQweAzeSPuN+YYrqjjTcc4vgaBuzqs8YX
vAeLBE4fYWVH7q3sdEn9hLSFeww6sjvZhvhsoBdhVBDglmFp0+gtLCABRA40mmmP
nfWRcvZVYdFIEcVA+u/v+XWBIwfwHuZ9AS6ucyvYAzZngezr57hp0DbuJHdP4sjv
FNNMEp5a7Le0mCA8C8zs4fC+sGt5YDJtfRthVY1TrbsRps7eU8noY9agZVIV6HX9
2wpRa96Hwc90MrqBiYItm3X4pIrSBJuKOoU1ABVqaDTuCbs3FHXcWmDqeZEBNvwp
dINI2ohdOzV10gFgHT33AWbla1p/8Phy1lbOHdUelTSiunkJN2IhaT0Gp8s9P5aQ
vdZ63mpAg/ospEEpbkKTdg==
`protect END_PROTECTED
