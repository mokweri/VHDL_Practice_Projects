`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyH/TbkqVSM0Dzy0eFxyEMmV4tpvGzXdOmvHIkagEDDzlkyQqVD82AlzsivyUTYG
YxNACLkXhqeQr87HFObVd7y0ZZgYNWdsj9rujGUY93IqeNuDIX5egSBV2mIpvU65
H7gJiAUjMUP4Y9II/4unG14QL3uUy2j+vfMlm0rHD/puspnmMVut8gDZuguUf5yF
oD8WWE1FhmaAO5Np+C8UEsoeejuISBImphgcZ6zdJH4/iB962U8Lc4YTGYqb3Xmy
RgfigAk0Iy7n8bGKD2E6zBDSrmmVWM9ZZtp2rDTk+1/cz+7Ye5LeMbGnngMVWdUF
qrBwZb27tPOvQv92cIN8sq/8I2GZq+1lLakO7Zes6A7BVVm1soDOHg9nKPfOKD+w
Sva+RZwCLBmV90cbDLEReQdiTaF2l1wPzZiU5PaQTGTkA6F2CzNByrXczIq3GAa8
PP0kFNQeOfK/1Ktxt/bLej/PeeMA3O24Zi3v1fC5Pq3YeOXnh/1O0qZpJBYyhI56
epy2xKk8si8DvXemQhCu/SRZP1seKov6HzAP478p9vWDr0qgLMt4DVAR1vdhg/P+
2OvD/kBlambhWAfKJZs9BHTAkjQSbB+9M1dmzpj1OUmcaQO1rWvxNFIjJZd/blAx
5eFFizjZIlofE37VGt83Cg==
`protect END_PROTECTED
