`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7KwQVUku6clUr/fO5G2zAVwnB69H/612bqiV5AxW8WYsf9SCWOPaGVczx5Tl7BIZ
AO1xlDsEHTKzcMWakYhkbGr8ZeytCs/d1mjZKfa1hOW2MroTjXGn8RLUdlAon2WE
pnQF8M71P3zGqt0KcoJ8j6bPg8mIpX67tuTZI8X73aNnjn0C1p39eeX4oc9dY6N9
fcccQXVZ9ZzxdA79ANDCPMtDSrOCcU6XTA5usLSKf7bahV2KaBuTYjJ7U5uyxTfj
Q6IOvzRE5Z7yJ0jVXUp7QugFLyF3r1ZmIrRWN8/BoVCLyKEgHHYMEBR1s5hk5NIM
NOVujVf2r+RNNxzKp1m2sKkqla7SNpfCB+mQ1rOxb8GBfLRpdbVrEM/+jEv1Ffdh
6mHmKZO5lzitdCtIrDs4g2NZfYhltLQVg4JTOD+LjZWEcv05H9o4RXshgmNojwbB
Y+md0N4t0cVAZUEu8ICXZQvgVNVp3Z4LuR6MCZ4qfsuW4KPEvlFDpHu1nLrsvxP3
yWF9qBD/mOBwn0fI0GX4t5Ga+DIb0kRraG5l2b1cr6U1Y8vEGOq9kGIB7x1VlSKq
mwCNEtD7t1bZmK6VljrKMGndEY63vYxYUVVz5EuAcEIIPmKhRgQ2UnILmj+UVLBn
pyrDmP2fDus3eg8BOOzMeg+RiupjGP0mGo2v6EEVNgB5uwljV2mFLEayYkCBUsxu
+5pPBQHDrCRvARHsrbO9HcCbu4onAdC+qroncWedMBDOYsBnnDlOnlaNhjUXuTxK
tZxamkD4H6OCHeBS46xfgjQBdokVbGuYh+IuBeZlLwv+jFPp/8sZE/HOS/DS+5cp
lc5R/5z/zO4NhqM3DuAXG4KGVAoWtwjwx4lpdJ0AOqVwFStPtrC583QJdIUCnhZ6
i7VS3/2mNTk5w2EKt6VuYc7wtQ/7i6oKIL/xtIXApYNY0AiM9756CPl34fv0dTC8
pOcTt8LqXOvpPHDsU41Po6jsgTBZC8/vTi451bzcxDds0q7LZEgd30QsoQR1VRCz
40cEldeIC2F0BaTyGcqE9AYYCr2P2EgI5oO+A0RUHZzOGWQkrPM1cQNPyk7JWtDB
QsgoT9z9bn6dtyXphtIzX/sEBnrfQal2YWSVeptSejBM4y1XxJrQRQDP5arY8oYv
DPw+yjCKENq1Hu6QIO81NNISF6LFPcVfI1SCB4H/ifdEd1SA7g+PiAkNriqt8E8V
U/T3vXcciuE2NIDP5t4r5n/FrF+GGl15VZt/QEc0w54svRYJ6TpOFt/9mURZNDrB
0NHTB417sUc2pm6cNwCcBg==
`protect END_PROTECTED
