`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1cYoXBbx79hioeqgWvnpKhlL+f2eHPOOu9lul8+mNtrA0uqxArAz7tkppQhG/4h
xPXTTURrPrqq4dbE3F0qSo1cVMUt50REpnZp3CAHF7YgW2nwvN1vZpFrBoJpjAyV
NNDWWo4kDDg+GDyuiAMjJXjRggzh4Bu1fAwHUDCqE/8eD1z5gs+qU0owzk7HAcVC
rTvAuFkrJOVrzZLNhOJY0KGJ0XbZTKULESkevUdlhUlig7ne3eaeSivOnsgA/65P
Qr/aeZFEFvjyu8MWoCHY/jnJAqTAdW4j8LvE+0aN+ax8Ye3b8J9cSfaoLMTVBNhS
uT2+7uo16VjrEWrh4W6QqG1ne4xAzkYAS6tKvvcF9QQyndZ7EnR31r0Tdy+HyuKk
zWBz9cnP2zZgP+ZdCWJj+/uJYB2+evEEAmNyhAGr4wmBcfeF1OzvhUBwemkib9Mi
UFGNWpK7uLJkzOMKN0tCcnP59P6DxUB3ypA/at9ZkH6lOVWq2YBXTy9E1JBQJksx
5d6hyAq7jbNBJ+p/pWyIZhvapSQPUrgR3nLvpuTN5REL8Csy0k5SNRjowwczH1sX
EDzG619NIs10jBG8ZyEyMQbkSlAE5aJSROP0/782gDToJhcMiO9g6u9MYm69JRNJ
jT3vTppCnv7aMbYM1daTVHEVRzKLu+NL8mQmX/rLxAoFYjXlX+9KYqoIxhBBXEkn
35qpsHjQ2PGR5kc77MsaWUiZOm+hMS64hbr40gTMrzA2LEZsaMxUo0wS+ZS1oFgU
c//ztAYGpv8WiCBe18820fCxVlNAJyvADNRF5AO8j5gqbYmhKKa0UjIfPtTzF86j
n9mZJqBjFA8+csgcHS4y/UrpsTJNFGmA92D4KizC08OSDcx06ehICmmQUX5xIBhs
Y5P3OwxEoGFQIMxT6q8HDUugblG7elK4CbQfTag2w5Q9KhSvMC+X0FiE06cbWQ3R
besiTWX5GojYro6qxTVNYBowQ4Do6kYU2ZGRL2UyKbfEGHGogKZ5ymjDzMSi/GVt
lnkTY4f25JMreHR7/zb3pWedxdFdlRUe5UCFePkpRSvy7qgPDLB56a+3i9JZduvZ
dcljUK9oYf3RBOuUTKD2PmfLtn48yJwKIHS6CtvLvTbShS4rC0HqHVT1q9t7fYlY
2ChNYO/p6gGY3cpg2ZYzQu/1zifGazp64BlAVapaZ2+z6kGr/2z3mfuduv+AOq1D
ShVlCMWIExx6DlZ43axlQAI0ng+f1ETYz+FMgmknTQLOy65d2KMAq3HXso2mbQzB
Aa6oLZJyAptgMfeGkIKYEzK6tBCBH6YtPNXx7BGh/hS1IqxvCpo9Ohkk9ej3b9xC
rTHD4/vHgJXojX+Uyu010+RTepJaUf2lv6qeuTVnRq7bdXWQrXLE1xpvvZfvlV+U
uzRvYL8+I1Mq+TgOKEsJA9dGKeV5MR2cIRc0th/dxg6AKr4ClhxQ/VdOCYmgi0R0
PyEL+HXBfP2EE5lyueRR0fMZAaWCpSWmraRl2JnZcSa7b6k+A0Xq6Fvlzc60DyFM
7+mJ0rYEIUCf50aARlCoV42vjWrM5b+bmh1eQhB/fw3xxTsVRF9dDeK2e1+AgRdJ
L8N6ajTVW04nxDu5T/jUwhzEEos2SWfziLZB9PiJMUO5Zh5OPIqnUQqYrYv+GgvR
+i+m+f4CIB+xFC2mjPkE9WCLin6AwKJafPbA5TmORFgxq+g0Ih34vk44lwbVhHvM
6QZzJqD9KW27HZRh604Bt4OnqPJjnA8ip2fpvDLxoNT3MPpIZL3JWQmyAsl3UX24
iyM7HEhB9FSIxiqM9U4d3YP9lf3nVysoEu/jLwNdowwHwx5qKWhzJrPQmp03d9gZ
t41DkFIuisMi+VYr4WkEYwamiIdv2BgkctkQPP17bHq57zchb8OLxQN6vqtVlO/9
YmgQRRPGU1Kln6FnjKcV7bo32ByiV9r0GRtZOsR793kYzeuEgzZLYehJDkJZsRwJ
JiConFPZG60tKOLUjbOcYInO/EmNdj7x5rzXYYGXKf++LcBUtUEE0plZN5cBQJHN
AUzYY58Oii8WCmWKcawKN/x5Eh0UmSoOL1SwSHc9ssrvpQpS1Gr9JHD8QZx5HGN/
f7tK3stl5QZbAyQD1/NGsC3MbUfM34wy8dFx/AcBf3jSCF4ufiwx6YI+YmCG0O7J
xhys83wyRlNs6dG6jBHPMgsdnTe9DZ7DrLniC/WqBH5+A7vgJtqbwdEwTgKfJkqY
7VtsxhzFlfdoq6EPNmNMjBQTalkoMZwXhZ7DN7LxKYOhZhGCVqh9fbSnnJY5mZ9P
CCKUCW19KvYA3fWeGHjGuT+4J7jMac1Zr8t2VyudRQX3MYJTiE+9Y7d9JzVemsbs
i/mwhBz60HfzJLTTBXQfkC2rWaWLZLWXiQbqmEjFxiYYGxmLTgb6gdW5APvie2IZ
N7JnVAOEFQiGwI7afVbfJmQhN3xFMzNLyHuLU7vyXcoasuXA8Iiz/qUjr6uA0hxI
nt6ruV+s9lkdOPGQwpCSZ1ed/v1koQSv/MrwF5iCYazHpDMYAGQP4vFgYOq7FgkY
ns3uvLOnXgnuEIJksPI7I61jcWcMcUJPz8+xKvf/OL5LzrpIPnK66UK3RORIBUqd
cF1Ell34uLwIqw3G039elKKTFGz8YyAx/qfu5SAb0kd/qdWQ5Xd7GDKZHrNYmFWS
r816/h7Jr01eH5CIQwOG5pTHetZsElgSK8IScoqwUaaWh+RA+S5OjmtZdlXHWyjo
BRyoojFryvCBHnwBnLgFj8bMXIE1lzXqt5f29XtuOgvsIg3qFCUqoZuyWhOA9KrH
59Ojy/9h4yFxE9NegKNZpU88IoV+azgI2NXKYS7QSnqv2yTki7T/3TZd/CesB7A4
wnnLgEtnY3MuJh10bFyQvXuEY174npKVUTqd9NqqkeP82Gm2NLZFy342DTwnExBm
wJiwbTZiueTEn3MEIw65T/eVeHP2AogrgomylkA8bX2zIFTor4QMu5nv7N2OVXId
aFiiKoZ0v4+U+dxe3rxgBiRJkNYEyO5F9uGMZ8b3cFt7Gfae3CcQycyw5rbZisB9
i5XkI3DQXSci9Qn3q4uQLHS6ZSS8bnpIEZ5WPySi2fNw2AC3YNbabR4B3qBx9c/S
ia8hGuIQyPZkaFIP5tvGoBIhNWYIdO2MY5ni1ZbNH6YskZwZpRvkXoJNSccBdMEQ
ncgtPaIrCkfuOVpOipW07AWoQ6oGTJc+YEVymV9NLOU2mWi0/YxxFrFJtCpUltpQ
gC2Q1KuaUcERMXp8ShNSv6Z5WWMS+fgPk+LDD8iOtlSNL+ZTCZTrW7usF90weiyp
yzopocg2uNfc73alqQJI4tjCa0V52d77w4nsft1XnAlfZUN7jHWAsaouCtJuB1dc
VLfwdC/95wPHsSfq+0Vkx9tykfm42tk3lOqoWGD/mJ/TMSUqZTGy5KJ/JHyV47Hl
YDWOShGOgqdhIny0rxjfcGOeOS+Ow75EW2Cx0Ge/MhsphwKVDXteqwne4dqjGGJy
/HiIsPJEZ5q0x8jnYofIuF/gej+WyGlWV1OFjolQktK3pSpQjC0HwRKeuLWszIUz
dwbkGHxh9qQERqO7jb/eOfbU3ehHhuT1w3AcaAXCUbmctxDKJoX4lYX+sEYIITru
FvYEGTF77Zzvp32xd16+gct6Kzo/TFPd6QvMuAH35cHXsAXZIghCfWGWnP155Pkw
Xt1CFki2pzP3o0Q1lKKKPtuQo+VuhmqgU1Y6UULtzQRjyFIUQnmgFC66tPPptfht
aUpOqamY9HKSiulYu7mYCSYIc/j1ewThVBrmXbWG4Vjl9gUCP7UN0DhGydPFeDgy
PPWOUPQbWp8PoaHkw+B277SRNa1k2pl45uc+8inMgLjnrrEFu+adnb81YhDBpxBI
c78QbluWQi407yH6GK9FmhwUZyb3jb1pr1MAoOvYL9UOd9MSCf1aMKTlabTlb++J
Q5rwkjJXVSiXbkf5sKTMrLsODrINSgkgX8SuiPO27TFwn8XofAbQe2B3qf7gx9Cc
WHZP0WRyAcve0Lscz3YZ/T0tMtbI2FBiuN8ySiAm0giOyN5KPskZbXWXQC2iLT+m
y0CiV1bAwI47ETuTDdh9yjK9j5Fkm08OcYu/HsiUkk/A/UbsM/CZR26OwUTSegUo
AGamJzOiE2HGuOGsR1VxF3XpM9JYutEm1jcwBkp4JOJ5Q3gkDWgc5bCttGBN8Kjp
hv6B2b2DxAe5ESK5DV2zabXYTfS5qRPujMUfBg8/fK0Oq4QdBH70v2SX1Ud9Mh9Y
+eIF1zpkNguEGqkJAx/MnHITWIicToKyEAXOuhQBM9w01ekr+dWyZx0p9yglE8A9
x/XwuRFoNfL9fgXSe2x3VwBIs3mgOAkPWkXnlSc6u4EZjI7H5SaiairlbZJaQOea
2CHXcmuvtEzrhRGGBOqiRlUxBqnZiN+cBfBQAYgMDUJuQ1F2T7wHChrsqizJfMvq
RcRnjngYxABG1EHj0K2CR/CX79F/lSX7er0jk2PnRDqKFGD4Y/p/WdHHKpRZnpBv
21ZRhFgtNUsisS5nBUX6LyrTrLH3Ou/QBfSqxVPrTSitMaKYFnu3XeXNuVA8QgmQ
3GCL5vs/dy8HvmxI02TuZ/mM6QuT1qXWPgmWvADanjoNDNZDivrejMJmbbB9xNkp
YflOG+u3uUSs0oubhSGrc8I2zN6nQUw1PyLq7gSwMEgsmRQxZCtUvPaa5gDc3b9e
cpO6zqFD7cuyxZbgjzv2FZQNx5LSx392IRHhu4Jm9i+LOLyrn4BuCen4IyBvoCvL
UdPkpCiLKaIQQ38wUzFbOe9y4bvGCDCzAOyyX7/ilD71fBMX7S5q99A1v7U62usw
64ov2mt8azG6r14OM80z2nLioNso52vPtIW3IRfS1svw7BU/b/exCnFt8/HFyEOy
8WbOftX1J9J4yiZLIrfpLXDXKFJrwK/x3YM5P4LdaIYJ6N1fuk61qyigiHsCG79a
gdXAFX47ukt6HztrQIOE3WHBaauj3C+3RP8Xal0L9VzU3o8iJFLTyHEsfDLknii5
V7dl7Mc4EWZusRkhKy+O6UL7has2xZayyit5oioa1N/RgkahO7/ea5n2if/9ePHY
EungGX6wkBofjCAEN7Na5thMD+YPz7CzCaqKxjXvNxonA9k4Tt/xBKIw/64HNgI4
21C5asCgmPqoJRZJsan8EMrBEnr4QncRHz9COgLyg/3n2tFdY4S4Q8iouidCLahu
4HxukTYIfswR6mqfDo/i0TTwqgMirE8KE3U2rSmAIi79ouBs1+QmrBJsGwRdmJL5
UEdzCvsLDdDEJL74d9Qt8zg5I8A8zqTGc+FMXivY+VocB08sRJRx73V/iIxTETEG
GbQrf7IY8QnJo5KhklHZKoFYmcBXV2Wlgc+HRFuI8ajY1Cd3Y1anrrNeBOKxXhae
WTAvzfhpFlHVH0KoadJIAsqiJ4TQGQ6I9xO3JGTrbc8ERcOnpm0+ZOZfoNtk7Bt3
F0QXgjqaGHVW5a7Bv4Jm6pStTpwjqNZFFWofdCXGjRlOryXi5rc+m51BB/fK74Hl
LwhMNg2l6YxHQ2dwEv86vrs5t9EWL0tN+YLPz6mJjhCbxMe2U14wN8+6gmqPNAYN
e0SD43jvgAUST8ohC7JPuj2ePjYfDuEn+dkv7Quy6wK0BdKF7aZqRnqtVNknHl7n
U2UTJ/kHsPUg8apkgD0+UDEMDngYagp0WCm2mFAUW0XqCAtvnYi02OJn1Ws0of47
e2Ievjt7K6OcLH6aP1sFVWxemAOw48ATzYvCzlrQ1Ok1Ds8K5eKAvBnBkkhnmK1q
gOb1Flafc6Nm72DMQAGGPlZIUbhCvPjwUxL2CBKnLkgeiI4PlktLwpomb3QcX1bx
J3mivU9QEN59v4O3/k8skKpSeO5UkpdjnDwFeU28J0CKhSnknIkX15yM+moSeN0y
7HtJUFG163f2BoF1ItZeWqHTTy6K8r2jUVnMnJk/JFSXdew2j1f52qY6PFSjQXVB
`protect END_PROTECTED
