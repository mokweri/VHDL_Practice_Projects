`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7PUtRtn56edsp1jiqV8L6k96Poy1DMezUR+SJ7w/nhEIO8SAv6yy7KVwi24ATmM
04Tl0Z0xZKJ8AaA3VPZo55mPIPNGrfHHu/L5fI4nJQJ8TO8mHzlgvsJoqmytUH0s
Hnc2+iTM0nYDzVfc6Sx69roMSNMHwtTNgzxVNK6TFuzEgSnnpgpB1n3T++LeOEa8
bvh+6EoHLzqK0wlh+GTc4+qJ1Vf90Y1Ui9QG5lV8J0r8N4QcF762iwxVa2L6W7nG
50YJVO2eL+HmUnm3/+mLUPbTwv4ZVGGvmB+xEVbROgsILeid06R/auAvLg6bJNCv
hAyDYpX/T28jVILyyJhy6Cm+RrTYx7cax7/rM1ZFoetv6+Bn3Re8F8Y/XTCoiNwQ
SjnoK0T8BoFZq5TZ4Zwda1+LHKNfUtqMj9PQzho02VFLZ/zZcQrpi/7NqZsQ3Vny
HjAKsgtSYfpHRcBh6iYhVckd36FIXsKh1IikdJBHtDqZW2r5DOGC9uFhKhvJJ4LL
I5Pgi+wQ6vpJTFwc0wHPmfAZ7Vz7SDVyfMNek+go+BWWp/4sPOc6NyyrczDaqRDR
GVEPKnt2Hp1tE+qWXUTHZoxqZK81+ETPkHC/tPMrEYcYACAkDsEyTx8pLCp5JWPe
BIBqwclptvuuzG6XyzUxoazt71c7ZgnW1LFFuIcSKrkAJA+bcXe8WIj4pcLbugM7
n3UINqMZuARu7MbV20y8TpIdcjB1RnhScd28FnVHCPYLwpAvpbjQmA+jYyVtAYMa
tcCvHoYP4jqtQCHZNVEYAZRPjnfASQPy5yIB284khdQIiuoocG7OxPgvDtvx4DFF
fgeTWPRVWjDy04JqXlGkrSCqJ4XN3yI+A2v3AH0rjv+tLjQyskIolM9E8fGedN8s
tz/AKFtZgk8zYfv7KXazIao36FeeGr0oi4qfTido2lPYjkqc7cmd6043S/XmdtKT
812bmgQl40Z8rLSvfdSV61tiRCiynI/7UOeLp4ihbcKljnR/vxgBlkB70bJFAYC5
Kb7E+Hhavjco/DAdE2iTdGUOnTVstigc92PMTz8ML8sVDIGkVFkCQFY5MpxJHiZ+
NeSmiMPVC6v6zMRCuxQloI0WNgAy2silfw/Xmeb33mjRZcu5rnPbTXsSrdT0xjC3
o+hNlikbijieGN72h/y7qNwweaa6OA5zNeO5uYRpXq0riPsv/uA689jvz+EFuHM1
fyf1FKheM0Fd42Vry4Cmy6qbriJMFJEWJAmHTmzFN29ZNAjUSEOowSJxD/N1c7C3
X/mThhc2Fu8JsV908msjp1MrF4Q3GLf7E8U2l3QFHmy4Eh5Wr+HTslRnXj4t9gcp
Ew1jy4NuQI8UAUTVASkTXkrNx3nUd2DsAK5m/4PEYvzykjrktyfWyxxVGPwPlqmr
`protect END_PROTECTED
