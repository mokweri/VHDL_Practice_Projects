`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8EW18Sq8j1r+Uix/dw/Lyqg3h8L1rELme2DgY/hH2c5BD2cTs1fJEO7MePB63DD
EYbMbQx2K0mcSD1bXjBwhzLZhp0loqJPwR1FBgJ5Bmh/BashSJ1bbdRhMl1TQbJZ
gEv7vEyZ00kxlQhyi5Q9FU9DDymn6lG0ioJaMmu5DWn5txgdP9uTX7YHOGmnMpnp
mX3EydojkGTMtXvqK4A3dXVxFu+6CU3/QIS1zT1Hpa7SClvCRFHBf7r0ZlRHlyCP
FeioZTirxiL99J45gSIX5m4c9ID3Q62E1M+wX1CFVaSXdHRjwInm5/7dx4r+DMmx
dykB7Ng1NQhCF21dAlZXU5JS2WdlALliqO/MuG64EpIsq0WX+LnBIEFPrS/D1IT6
t8S8sVpjBKdgHTonmhEokaxPz4AyrctTy+1uCCa3tMGZUS2uzzkFx1T4jEANlNFR
3MaCM6qwkV78EqrD/PN5wDmtOwjjElwl6WbwsMGT1t7i9a4UvCX4iTYexGSNufuL
jXQZRFZrlV8bW/4o91QFi2DHLHljhTNyZO+AM3tpeYV2Xtr0718Qht9zVFMQhs3f
`protect END_PROTECTED
