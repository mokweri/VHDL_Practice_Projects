`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yflu0Ay9IQJvlPXcEfa2BSQ15g5ApMmgQqMkUeBcDJfuyEYLg7MceF66GnIkGaVG
mXGd0eZEHTe0GF18zlppMTb+axtqyzfmt4VO0AoOnfdSskkYnCWWPM5CsHr5YvlO
Z+erg2Uk4OVdzfzjd5vgnBMeViREAoEJv1ktE27CXOUQl86MVZ9Qh/bb6NMY2BOU
ySXR8uB9M9qJJqezdbpvYgeqrjQ1JyvTjMxrlgDhxfOPUpx+DBTtRCZMjXzAQKPR
r3heqTJnkXJstzxVG8d2xbE0qyS7gpY3c1jW8rX+QkobGx35iOj9rRXI3Djuz2RT
Xxqfe+SmeJjP92WpP5zM7VXhsWqimSILzs0qhF4PdynAMrVKdovg2FvMKUBJc5Mn
wSwb90Rw7teVmDcq9H5mMhwugjXJF739B8BNLGkZE62ByBSSVx9W7rdbO4pWTIMm
MeISZK1EG4VoBOQvOfcWUg==
`protect END_PROTECTED
