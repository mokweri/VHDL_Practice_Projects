`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jkxhi2leBSsnNbUoEEtE7ZMnjH1FX0A9v+Ry2aHLb3ruzkklgHchqvGWWrV/57kS
5sgHlBvzIF6RKpZnOgbVaHdrwnb9fU1Qj99GAOLIleQrcLkrYloii8G3HORzY49Z
k5VzTlXpx7eI3x4kKinTaPoGgmobT0aBXxFdo+KWNUMcEs4lISuUdf1UCppddxZn
Sr7maIEycc7shkcyl4cq1ETUmmr2I3JKmiNyQ5A5I98HlWl2maUH3XKeY+bn0n+r
agNixYgs13pxhduFy1WS8wta3VAXnEhySBH+uQiqBtf4CPBfeyjguBTOofgP65sy
UX+3njdd0xKG38+SmhzFLh3yPmReQF501QQdUSiJcwlda+NOQb1Yh18wbd8Yr+Mo
yB2EjHrpkKDh9r5ZUmKu8+94YsOcBa2ERFydlTD5tfXSWkjYg7K7gjdoRhkT9TSm
ETZcb1L9Y3bHbu+CXsv3y/e5mxwiFX17xdxkv0IDU+MI5Ibh8xw1xLL5IWvgcNLg
L9XFpknZgZBQWjSzU6uIVQU+V/DUENHe2i7X6NK1A0W15f7flb5aiXC3Le1E/mUe
BbTXaJhal61NoVBbir1LAM44okYvYVU3fv7f0hguAYOe35Te4rUTbZCq7fxR7p/r
c9l91yoZNqug//lFX1PEpznIcTEB7K/uhmF3FfDr4rQxcMx4rzTsQs+LA9dt1NJN
/wAxyLKLFeZtdTHOLbXJW69mj7LA7GWr5YoOdbK87/Us4Yaa6Dgqw3No5UI7x7XZ
vXHSg96gdLLjq7SNDQ1UAHcPgyMd6GwzPYv/mk6D5jn+wxRehaNn4epLalIz8CZD
UJK3CmQkIx616CpilOTXCZEKqzAHXeIdtr7LIoCW34lAb3qBiLWXlob+YT1yWliZ
z8AcUYeCHuz0tWwwpGQkn3vdT7+hIpAeKxxp7yTsuCWi5ZSRQWO3Uy3gYoyw1VIs
JWC2Y95M8InR4ZAbtY0hCEP8pEqPb9GWF9/1ckGoQVlt6aB504UYVIjSsZ9aJf3p
O/ypgtekCW7OGzIItlHWFh32zC6lOFLWs6SR8a/O2WtvrTS8G/SK0kfh2pzyVRrx
jUwCzXtgTexRw5+INAWjLP+EbAPk2cWbiC6sO3L91NGEMcabPoLqdhibxPFr/5wH
SFbO9xW9anXIB9/2QRMmK+6G5RyhFr4mZPVFfIlqq981e2pdGktMIadYTVe0LE/t
Bd/gkg+q4+HRiGPzAFiPvFHBsPXE+blSGDoTddkbL0p1wDzcMIZxdfvHoIXhehj9
NgTzwoHvQKBjNHIGqZH9fiZhuCltrX8LDx/TMG7wQdPuM2Q02K3ezw0MKQvSGzcm
h0WIbpT0WyfypT/ZPmrviWx4OcSe47bRc00Q0MH3EaQPyQX27c96CGWqLriXV81M
u3CD0qa/6p5WmW1gd5brQGk+LcnAyEa9dEiOs3X1q83NJeKrUscAymBLPQqlOjnh
Z57dYKX/+RdjhWDaUikLWK7vRa0NaoYH6qziAV+swT7nSHUtJRyXMfjg3tgiUUEJ
n/wjYfYBU87H5MkiTFJpeESSALX5lHyGjvhPW38xgEjorJB+mHsfE8JfTzGZdMet
S61J8ysOkLQKCOFAxGKZ+iTWCUOB3C4r9tHx6Ve7YAsyC1XhkCnfEmiafnvVbdaM
G+nBAAsBsEgLVIAAVa8xt3qr8+kzpIMUGQZsgY2yGRQBB8eMzXXiyZcM+ZUxBDqr
OvLLCQjg8aNIOHPjoioqj2Mc0gtnMn5yCcSR2IUcwsj/XPCn6B7Z5olTDSMwsZqQ
zKw94bSUjTFNy0SIZG1ZIN0D15NsLkQwCXdA8+JT9MdztLWLnIbO4uw10ZhXqPwx
UB7yU6wqShSAGa25djNePI5P/xDnTsQ34v0y6iG4xXTidWSRoK31+F5dIusrhLbx
4MqvYAdN3RpRlhnZyAXuH9OrW5LCQKa384150UgM07Wypq2/OgLFTK5aHxEdsqie
M5D5VjwYFlB/pI5s3MtrX4awSPRXuoDl3pr9XgFXNfPgbdxtb6/CjaJTSgw8TDM+
bSoZrCAqgbcZf0bbOvYb8zyCqobMHQTMzhNmAhqmbVt7h5JRBxSUtruQNT6sZPZZ
hansnH/HxDe8WYQci/SZ2QcmxVzZxRhMDSKu4s6aNITSwLPalSMuZfqPY647chyb
tozJQw+OiA+1+5E5T0EKGdVXry5DCw2mQWL/nc8VSHdWHIwtecJaM9n0uq2mMn16
VEmeK8qs7/UfwEHf02SGL1q4ELxFtK6ieMVtYetqULm5KMJ+Tp8oNwoKa+Tg+Yd+
tYcK4u8E28F4Z06JJEVhj71GTfQuVkvyqeDnaGm0ro5rkjWq0rBcZph1Qtflhac1
MqSrw/y6oZecgpjSa/SXyPsxBnP2u60CXnCUfh7azZFxiBmht1fcBtn5Lz2LPKTD
jSKxMa65zb3HnJqCNSCkUwM5pdCJ99GHuTgIW303A+15Pn0P6aQTgn2TgyaLtgVs
cAHChH6JJccNvCNlZM+5+BhoZcL1KA6ccGhutuBZcmeoMempD4OKT5wZVT0Dt262
SSMOqNI+JY+w+3w7oasAc0jjNCBGL9GGHaEdCQUq2eXDqgqGr6SqeRWDu/gXeJLi
PBCF5p5VqtMgYAVZpLAOsYurvnW363DaKwYd3h1w86Dmoqo7Jq40EuDbYtBjXK8M
dfTNwRa3hCeK3F/mu6+mZ1kPu3BnNe926xGPl/YROnnMadxY7p/hUc/EGKueVfMC
sm3Myet/jOBdAA30qbHdUmVxRhHBFgmexY4OaVlm8NXqfyXDmZk53D4LHPspdkmR
OpASCzGxXf6MNDYNoW67RWZwvJEU9YPHlK/3LkM5v39X+oaBFI7an3xLWXIhLNZM
h7mD5sXg8G2tzR3mk9EWTMMIs4B2/3HItye4jWLfzW773E3sMeV+X+ioY8/P3pcv
THCY6jaC82Z6VH5aUD+FPsBbAgXvzByJrbp0/nyE+KGc92ngupCoV1c/TDEu/pZL
WMchN0ZjhthEXqU2F8y2A1h9cL3NowPT7mw360A5yNRS8yVygXYiViokyzkOQK/s
7NDY87AvKCV1znlONlplieig0FynaVfKSB2WfqzW/Q+SI5k9KYcVdXlg5rC7uk4j
xluy7j8mbEOoQQKQ+E05NN3EtWsxSSgQsPeVKIWWtfC+i0shlGwwUNUUtPYsNSfv
WB15e8B0EdbZKJtwfxAVZDcndHPhXpD/tkFbSBZf9Hs4tlrEyPdD+s83Yypv3t7D
pGL2BYF+zYzARWjr9+dZvtfjZLtjC8mp5WtDc9EZsmtFrn0VOvOQjSeaA0Ynr7kS
fheHe/L1TeHoN78Cv4hcp1BpMEljyaE8W4bYwHFsp3xFbqYNAYPk/+mUHp6gP1FR
0fGDgzz7i50oj3fUYmDuFMw8y0DuhLwYd2J4vxJYDba5WeXAi5H7yyQ11SERc6sR
voVzzsUPX1APz+bWsyrvQVbJE1HnYYJRM8xQ9VM9a9ZFl360Evo8eMkQxkPLxjDh
`protect END_PROTECTED
