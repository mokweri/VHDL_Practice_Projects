`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
su/ZT3JfQs6s2rXRqx+kp4prP07KSK9GAvUf7nV+1w05CV15H+RW7tOF7Pt4d2u3
3hwZpAkD726Tnxa39+T0mNkBraQg1L/Q9tNqzdH0Bt7bjX0UxjkvjU97GQLpx3i8
myn9tgEWMSv5tJXzYmbtRnaGJqrt4r/6HdiyvWoISIn3kNhiqaSvfQj1MLxbXodo
kWTAzqZVm7OhTQLF6tVw1AiKP1i5jw6mPSJ70c9BkIgeZEwfM5OQN4IxpA/6732M
9eos1qXd4RPi6KxeqzI2F//OrKlheuxQ9NXIYXY52R1vsuwkY8sXi0ktg/AojCfW
iyyda0V4+b+Hw4MhoD213wc+Yj6buEvCGPe3j3nsAnaUc1UKLuf37DTLgDl8vNyZ
3KSqioZ7crpCPczJIO6+bk0zB3Wp2zDr0vkDIem8+iSLiRnSYwaOZ345kij6hJKU
p9N4OOVLA4wWnSiF6Yk37DpthR5DHqkc2fnhNyl6L4gfciYiNnKAgedKIDs/9THq
u3b7cHc9P56DOcr6Eo+GC3ux82LK27aqdHVhmINTlIIiEIvvvrybz3qjPyi5ChNR
HfYaqpkFpttI1iifhWzeBqYrCT6afbBJjFd5omPyOUYtbJ7SNzhsNNZXoJXJGUbU
ae1nVrNlHefMzM+AOKm+ILnjetI0ImUhjIaVyhveRZxkM+IYWVBYVhw9+Z1AozAL
ghq21NtH8PHV31USeVMjhZIdhiTPv3AsAe2ZyzH/O9Fi2zKEhNu1U3S+jdCG4xbW
w9NaivvPpXo2vHFEY2CkAPEGkhCafELG5vYTUq9R5HISp0umwVeARiUgjSU9gxcO
ZGsoWh+D2+QSWcEMKULgVScysQ2nOZmdvVy423hKtFs0vU/t3v+X1j0Ejkh3IGzS
Iq1YoXx38TuVWJbQsue9jYqkuLmK4NvjiL29osG94YVQJbqHM8m8X7suYxtnRkSO
qRbcgc8E22kquQe5ljjG1RkZ2IYG0Vjki36ZwIyWqJRvMna3kCokEJAmEybaedm4
4d3h6pyIJnrW6G9GWuscWKHFO9eZ8e6KMZgBQYVHMd8MBzkbeFx6rasBWtwAobDP
MFLF2NYGdCBFfFcF1k1iLKm3EMpAfGzRzjoYU/wzPcz0TBttxrd/o5BDhTm4ST5x
DerCb6U4QB38XyqmWjsKj5uYMMYYLWgrD7LFwmiQoEGcPNo/A+WFnDQ/+2C+mnar
WLswvSSXkKm56oSGL/VtFeJ/aU/xwnYXHDfv2jnn210PM85ZkSt+q/KFPbbiqWw0
6NLhmA3tdsvd0TFuuJm8aheVdzsntrQK6Pp8Ep3kZ5CEXeHc/KYqxZalx3KhCPAX
aTJ5PxOwe6yosLBLcEIwI0rWChN7geCQV31BJBHJcEL+D/9O4Y8Mztrwsesyr1Z+
/6OI5EJhzVWSzxTSfBBZXT/mHVNAgtn4npa5A89xZt/Tn5haKCR15UQ2OAvl4suZ
97zjTfNjefbFvjIBlS/S39CAJSUswZQoDi/50Qw4zUz8GSze7DkdyD+sFY9XM1uc
PpjAG6keEvOBV4A/sjvPp0o5373hlRr/kYfQNtic0SytiLAyRisQb32IkCFIBgqn
uu8jrmKf4ChEIK+6uhOzCuYU+TnNkfHQLa1uSYI4xTKoHpY/0iPYdhIodgWP8c8F
/qE04GtA2ugLbyg1xJ12CXC9rwDX9DA1xUi24PRecAoFaTdLo+z92ed7+D3bUS0w
uwVNeqsZhgBDJXETNduK5sdg603ULqTT71J6wPZ2bVoY9asSsb/lXcp8J+ES8XnH
2yaEGEPrTPaf1+TvTrFCUNMxHSpXqJHbkvJ53QUDhoy2UZCpP7X8IPn2KPREP6Nl
4AEHE3hx+mBcnglHxW8QJv5jupsqgw52L3eaSYyHgZ++DWDhgMKx39k4O5VxlEDf
kjI85eunU8r4Q/nDvbKvof4bCmj/f9ns55pwgJRAWqPoLLKMZI6/r3/04gVBt5FJ
NiRz72ila2xy/rcryMoTXiuRfcEvQpAM/vGMON51fx/6k1mdMYNmdGgfRMM+AAkz
URcMRLk59jYli7uuKKqP/IQaoKO4kYifdf54qQULXn1/nHnIEeMYN56IuaaxNVDu
T5vTqP1GABj18EH9fIlsU2gPVspueMgC/HeQSglJs7aQJGZERzr1HyV0l1BM2k6u
5KrX13UwhFiPBT1VJ4i8MDSBlUvCum835P5biEC6wkQMn0mJayNdK4PBQfFqgyg7
3AHKD0RiQLBeiE/zzcF1rl2x3kXkQOrxEAopMV5XBAzjf8tnWHvv30r+S2DV4qzT
sy7M5jSSgwBn9gH07FeeEAMU+O4t3Q4e+kEgXZaiZpsiGAInxyAsbZMk4cKhaNS6
Uz0OZY5nsthKycT3xbmn/X3Iu+/J76uvcbgq5onzmE5cBGtKqajYYrtYfnynDevs
YPq4j6KNUw1x6l8vFBCnPaoc9dfi152i/vzTTNyXkucGf6b4NhNxbFdo77TN+64G
+nwpd6l7lFkOPvnp/smDaZ1Y2/T+fRD0yPiER58RC3U4ECgZvsE0+cgfFSvRaVmZ
Qn3yE7nQx5ptMxaetJrn8kuaXeqOsRMn/YhGsINJbxYjR5cWgdbtsD2Bjg3X/ZwS
H7CQpOsxTKZer62bXzfyk4K7hg700FDdRuFy+ATqckw/6VBKwq0ZIG8ItEFbdP96
LO8KSgKh8/iIiUHN3SjMOV4ZiOfke4+wJz2cMVyPrZXXI3TRhZ5ZIOCWsB/s4bRj
qTJNSVBp+kTyY/URBV6qA40vPASaI3b7Scl3un4jWIQ3W/uhXxarXPGhPg/gCMBY
p1KtwPCashsprdTSXR9gp/oZO6umo4VY11E2q0tK8v8P4bkZdoDI5xk9SbgWUoG2
d1vUe7lYOpFKyaLjsSAdlE1f+cxNaqIP8+Fh2ium0pl6iWF6DFCD0eYknQO3wIaq
8zwuL02SkFMk4Nj+wWo6ZadMPZ1JP5ugntpNsst+3Wl09a5y5cuvQAQJoE9+xWo7
l3FkcMP3CG4gkLDEal96kcMUrlNXmmfdlcEnLHXux4fLmRiWLN18mha1ZGbvgcu6
pLbSjwduFHyj8kZLLTmWOfmY5a2xV39CI/wKlcctK1SAxoe+iFovvsNHx/iCYlU5
gJlY3SjvAFaRlI1LT+G9G6YkMeYcrS7ZLK9pbkapmseS76T2//DeN5YGGxItMyYS
JyVR5VX9TNLT3iTtaGqt3jzJyg7sIKiOOpsnhQROedWFxkRxvACUfIQ1y8ePGecz
ObnaWvLwiGSYysp53/mq9dtpr2POh6XGv73xEjKKbNUcsQzu+JeltlShiDR59V4c
JXLhYVMtppzLkkVXIRXfsNNX51lvsKgl0yJ/DBL1WuCBd8dcIIP8FQfb2dLFSTeo
ZVgBnfXKNyc5mJo28dLkwuNzL+7JQW/65cTyPZNs4BExuUGf97iy9dCQaeuqJqsf
2TDEekzs1LR6cJo2rb3Sd9HSwlGPK1Fz3wV1oOtht/aDRStqyD02dAgIzXXkLOyT
yxvylCI51GFXxIcllrN9AnmIc1poKrnyq2THJQBBCu+vFzYzfhD3SYyCPg/wWlvS
sueP1pYGFdSkk7+a9nrdx2nuT8NLKeC3AnqqX13UMyK1AZxal3SvyWebky8uze00
1GNSze0R8k333+B6BjgNxUO9T9LRIhez+xccmjPqln0gnKwePm8/A1V+gNgYdo43
ZtwxHQP5zHS5eUZ3vbkxRCFy75Au7WuLJOZIsrCwI+LxNSKwLvkELGxf5nsbzALz
ODglFSESBZQKvCyDnJJCu2/mUf34X+eJSbgpLtzhnoRd16x9qtb08vsk6NzKo/mb
yl1Tzbco0gGtu8xnVc0TOR4NGrb2suczeez8Z9zHsnuAav7EUQHDU7crwzbuH7Ka
+UiyauDsueM23H8Le4wKsOWV7vL7V31i4nlzkgdEdHxEAQSPQi/3i5df0xtddD1E
eNCN4tB7+zfqkfTm/I7I5/HC7/70P+x9Psn5EuaW5Mk3Vz4ddvYirlNzI+0OnFP6
QKoWmqJzhVzq0h+IM4GJgOPPNMNRT2JR4CXFfNAtY9SyHuLMxjVjSvuEgNZi7HyP
7PuBGQNIYOvS0AZTrZPvwluGB+WJ/BQpjxZ6Fuh3gvDej1xYCA+PU2Ryvi4sNd0+
qByfyiRxpHVeiKTrYu8VtHCfVRh2Fty2iEYQHcTee/G51s4Gah2e1CkDV/MkRVzd
G0cevQyDDJ+G3167iFs/wIfLgeMEhCDzwjLaSXVRcRvT56PIw9hx1/4L4sKkzUsk
QLi3Ws9IpuJExtjb5YX29Y9z2hmjmArCVfdDigVe27sWg5xd3gPPrAd+kfqOeRZl
hku0XvHDKvE2sY4InpwEa09p09mWjKG06+y7bGXqZJ3W5O2MLBDGBtL6FCwGcGqU
oJO2tseHJwpAyyleLMhso8A/09076jfPCudHTLnC6o9HLNIfU8ffTSj7qG1OqnaO
1LvNrHPLj3qmCYK9NI2TwfO9MfXtz/bsh81c7GhfNSN5KeBYBdPJaBHxER/QCFIm
i5BlhjYbCxAxd8yk2gAGijSPbhyLIFFjV5MGkv/K9ZQiJwsar9/qHxq2VECZlWA1
6s4MGGAiduMF00G5nx9hXCrdCCiOr5HYOVtpCi7MX7QwYDBzGwx5iXY0hUZKXh/k
aW8YxacxC8wtNHPsAboyDQV6QNkYSC3aGP2/egTmrRPNwo1HGuCogWEkthULGaAR
6ypoqfwAMNjKfFIQkDg9++apnQYypmBF20g+QcadbjvycrcRk4Dq8gZzEljWQB7q
pagwaU4AafohFuJY7ZDFBLZusZwCx2ZZfpZCnt2Sq8AInLad0S1SsaLWll9eWV4v
lxVDVhgs2Vh09v5cZgS/3MIUEg29KqeMvOhNSNMAMaesyaQVma6IUr2MLztan6C/
xUPei1lL8LoetpeP9owZ3YDSMd7/HBew5bo5I1CL6UOaA4s5CSIceH6H4kYf0UOo
nLtZgaWCrhhhWiUjuXYO9FvMkW3PB/lwuJfupLT+1Vjslwq/CT4jnqOBVpJB/zbb
i1obqoZVU36fqzIGysgINAf685xwWgS5n5pVe9ttnIZQZClwoX1GWaQCvqUOs34M
nb3ne6GQcIOA4pI+bfdkc5IXiXsLg2eq1x/f/Rbisjz74BBwmk0iFYmYUbM2F8JY
KN+kABgrYRuvFQOwPzaog5VKPIGGol9mSTJ5gSc4c6Q/GyWlrV4GmSUb57MX+23H
EsKZ8roUcWyijA9XCH8tBbrCsvzShVLeNTLYy7m7OxjnImuI6GsBYC/sIK4UGWi+
F/sCz37DtrZl7AaVU4Lll4mNHrhZBwZLUEdCk4xk+uBlzsghiosn96jNB9bGA+0q
tf4kw90xrjxGMkXk//LVfkB0DxbBZ6nypX4WC7hoGBQL+gRq393FDNkdma8OSHQO
mySnPtVvSS7rVF7vGgUSDfaD/BuRnP4eGyVqmzd7YlnX0+I/lJml3BMaSDGuQs71
be2g0mphj5ympDIpuR/xbbd/wxpCmaBP0vN9lhzan6zFY8Ia0krwQL37HltMBM8D
hNvoPj0HVK7GCZPD4xquPrMKvQUBaO64MOLNvGx2/sm5YQTs6HVA2jyFVFtS4Lnt
8oVlsHhnMZjBARzEzKxd4RNPhVqblqRYfzU+faObfe6TPJkXCckPCYxBN+cZ9mPr
q3OFA3PZ/RRaWg0UABNmpVDp6ikpd+3R29tselhJXPuhMdiNbD6dMg2T//rLX8at
FRkALWdLrbBkQz3W5+VOTGKoEIA6N0KA+qWQwCsSMPY=
`protect END_PROTECTED
