`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5118kGbiEYaVLoF0p8DvHHBLPrFWvAUdKNDdljsGPEHF8XJHBODCoCG0s8Km9gZ
m4l98bdXugOQxB0+4N1djTNRqfV9+WwFTYVMT12dkQVMVw+f+JHvsNz4RmFj4PVj
F2SDViZKZnhm2Rw1SH0Oro3izaaxQyqalHtaDjPuJDIA45pBUUdqrCXgoOB/hiBD
Tf22GKvp1n5iFLQysuqwRAJwfpZ6jXLlKGh+bp4Lv/TnONTZeKhXAKMBiX6HtLDw
fWYJV6urYg2nSTj9ExO40JgDO4VflGj8ExiDhjX2i6IPq5WXtvyDaadWESpElkRp
r9iidsp60ZaJrl1bMhZfERKQHACqcGYIKUxVGKqPCw17BHG749MMpeFZOLXX+kA6
g1KGn4j/CQRAXY56xTnGN6GA8tBYCWmllxrIE1zA2J1XL1uMZwb8lAv1MZQswbjR
p5BabGAwH5KPYiRM/HFXWI/BY0wBFn2V2QgaV/JMtNwMBMi/95mt9i1ITz7+SrL7
C6KkWGd1jyTB3rAVRHIDdUK+oemLKPI5Wdn69OZIP5kH3B8mSUtqCMB50Sz5VuA6
qOh0n3vENnWabRs22Pvfsv7KeqgaqsoFrSQE9leD3GrqMhac3gKoqE2Vvqjwljbd
hOW+bO0EULSACcCQ0kgEtrYbOwhhaukfR3mJJ6MsnzjUg2WwO2NNeijlizjxTg3G
1c7P6OS/70l8aoweHoEckRxNUpk4vmKuwM1JLhOj9KfpXFW9sMCMvcgdK0w3DtUl
6JTOY+fZcz4upe4zqEsuon1MnLoT3/mc8s+vohNZ/y4HDRcbm6bDyQ5LQfhG9hzf
BK2ioO891mPA8oAmlgwisRrD0yfbZtB5zw9qakRS1z9SXuD/H5U1cTR4gIrLMxRj
WsZiKnDO5X7vIJY01/hzszgiBihI0pbf9EVN1c8fyZcddg/mH+MLNHs3aNqok9Eo
fHIdotB0aZWehlHmA3qxrouZvNxwF4ItnykTq+ELH2FobM8Mn8M0kuZwzMV6UWtu
60w5ZeoEmqzwpxxa5S5LoZ+cfyqAprPMjZ4a9b1To1gV7/M6BUsJJpHLY9EkP1wZ
ABcEM4aaZoyOMphHGJfgaakjSRwPDVXas45YEaXCDWiWmnQHx2WPyGUwf8h9MMAZ
Wi2srxeAciclheALgD6QMA4QKoWghQFAP4qzVjYaXFKvys8coH5RIWpn9CtKUfMr
xrvJTvqEPP0Po/eLgeV/ctlP4GzY+xtJ9dqoAmymmV8+2aBKU46CFPWuWickEY+M
quiJ7UuBF7va3Rduhxr+URiziRcn8KPSqtUQVBt31wGNqcop0pzToE9pvXPoXP47
8tk4RvIeuQTqrjrAimANURo4jtYmfmlKlzbUSmTfr2NaSupXbggrCL9oLxBO8goJ
tkc2EjOhPofaWrrD9YtHg68Dwun6U7ssAkN4oiacQUxze5aHG7TLzbGz+8LlYgpz
BIs2Renwrg5aMhGRElPiHxG8RQrZwRuvez9SOnBJ+sDSf+WbeGS+WOEbvm/y2PxZ
1QkTXw5QE5wuSMurb0W/Lsxnfoj0kmEADQZ0vdtO+GfYoAy9HC0HtOmWubj/Nhuu
ZdJrtAcHFDPLUxjCxaPZIith/XdvgUQiYfY+XO4CSQ3TKQraXzZSMe+rJeXdYBGZ
BH/ypaXTbzLzda5CvyFCBTwbyY+MH4/1wz+X85/WITSeuT3Z76kYl3etpFTE/C/a
AilOSLBCIomH6M07TUuwXfhaf+BdWL7w2h1UTM1/FNMUamP+mdTg+om+Bai16W6l
0hq0TvRca4ICNzzPFu0ViPs2aulJZoQFXwY/Gk33XEP4JSIACbo4fFair++he6Pn
Mk6nVTXezlGELL9XrwfAIv2XkcQrYTpIOT7xu3tP4URTuvCGd6hDl0XTNnyR3UIw
qMpkyIcXvyazchpopVyaFu2GXsZIuvk1gDqJdmoFN3ULFNSjrWAcAbjmCIdOp3j2
dyx0xTKziqcRtbByAB2TnN6lN9lwgpBmjc9vZG7CdDKo1AaXsMIrv9zufjPT7amB
Xk07pTVohnlOMwbJ8L4cnr4IQAFX2wOh/IxuODh/vhhMCjK+c6y14yBbWCURkmsD
39lm5uR+HuXrlydmfJvXaVSeMknVNaaUx9shrhh/ohaSYv6P04WwVyT45kb6MROZ
lVWKu1hl7OSTswBBdYYtqxTJqRg3a2knaYtkuQtwWDVkh7dlD2Qzjpkee363lube
mbfnIAbl1twe/snWjGlTNFrgufucxfbNW5aJNZ91tP3Uf41ZQOdUB44Z6KOXK4oz
faceeS+xq3iB1H/hnqDHF9DiCbR+nntBg0ixaGz+FKhkTHPTvbfOZTAUjIxyhn0L
yk0Xdz4vtYEWKay+wdj8vrPW2CSDlVPprLeZXBXqWpp8U61wTZjIONsUn+yX6Wmu
c+bwTwrH4CZBB8YxRLxLwDM1avWeja8eeTK9XetU0C0qdPWlQhnw4K9lYljDFNj0
0TxHYiEP3nGBGe72nsEZfA==
`protect END_PROTECTED
