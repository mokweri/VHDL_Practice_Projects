`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGUl81fgACmEX+WbVV1YRDG/feYFYLZQIp9DwGNvk1aHFlXKi8+xrX+XwUYO8d6/
Uf3r1JFQIIPcwpuUHHJqPZlSsOn9VHGnLqmyMiYGVcEFyxCsT/mdWWum1QulQmWu
tIFj2/jLJC9yQqYOFegzLQ0vtzel8iFVTW4fCqjpn4feaOrX32vO2uRN7PsUA0wm
DSVyzLCyDzzIwoJ1yKMjPv7Uenx1XCArfrJo5OO9Yx2tPptgTy2yeGnn/HwHDsxw
ue/F5hw0sy8qVeBXL4GP//PuXEoXz+wkabMrWnvYSuaNL5AYQweXvwwCHMlO/Tay
Je7AXG4h1AUKVKPm/xxa2/5iJwY9JhPoUxltH7icPE5TRjU4cQDG0B3Ctw3vHWV1
63sdMIcwzlsWTh9biZoYHbg58tVKpBs8MUrB/1V4F0MusEJnK8CzBCTKi+BC+djk
rzmAPoivAYdOb0vzsiGoHY8bkh2ZsENeEnXZGLlKoYFIZprdKt0yhHDzZHGWCX1v
s61Pku6JuRDeoqn2JtXqLLESq3jP77S952+xduOx26aiF3PURzrKDqhbxVV7RWxa
tx+Q2FI0CFxaUOBpIKoPmA==
`protect END_PROTECTED
