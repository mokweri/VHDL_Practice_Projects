`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcb3mKWHmD4CWly+yYXioud/C036KTRGhhBb5ok6iEjpFfAzr6RskiYTIlNSxO/6
zNAkijGTmpAvmHuJLTLwCo7gHsWMPkxVOtL11RAMswpt0HldPCjP/EuVR5vr1q4n
KMOUdy7a0xROLhBDNS0lspLZeRJrKiRwK0LA3fOM1v54t8A5gMSxidwLzVRZlhFp
OGR4skubakxKwnRE04Drui378N+TMluOlM4/+eTFtSDE4xOoSnmz3mOQMk/sc1I2
mZV243dP3BnNeQd2eq2kMTS60vPbfhMeqXKVgtLPNnGRA6BMctm2VJgVzZsRV/H3
Fbpdx50eozYpHB2sodVP2SRH+J4WlnO0WFUwNH9yn+Nji7UIRoVq/fTw9Y0Cn8zG
O7eMNv2Qa0ZnOq0MSjpkaRFSo0qU5UuSgDAqqkFa/pVEqFcZDvvKzhMxhVJQ3UbA
kSvb3qsBSwrCaIar9WGjZhlHOMvtp9/u+JtVBuIUjRFZraKUQOC2RiB9vcetJbk2
UhbJjeBnm4TGuhpCukZR09w/q8Swuiwx7CLw7hpG0s39befai2g+woN502G+QHTC
oNV4v7vj1fy7OR8ow9gbXd2H+05K4ry+4sCzHBaq0QqBy3e1N+z734A1PmcyEoOD
WvNGzqCzD5JVLpfD2+LjW3F7fxUj334RmVLc9ahSTRXiqOCtCxE+38NglHFbGbcU
nObFEEINg1pUdsMuR1BiCz/HKKBulrQrXdMgSxly2rmVGBhXjbN0V3oUZq8aN4/n
ZKIgVKWdke5JOmqwU5HvACcffDoFfZr/0i/40CzfWU0NE9v+Reky+/Kudyv6rBxJ
q4Wp0QJnUaj20nPCteZUz79a5dT5PehqdGuiAXazaJJHVH43BS1B3BbZB4GwgLTV
JaWRbiTHyTo6IcdN0b7au/WyH5sAixjOVa0gWoMKPy0qjbxJ30p9r16RA1vY8fTz
+J7Z8JmypgeB4F/uv+vXy+wvACmkI9ag2w//J6zmIgAi67zUchSu2aCMBJKhqgDR
Z4U7qmuMZZupHX7Md8/J6X/bNZ+mgMGOYcccAw5NaXY/fT8926Zb5dL0865ROEB9
uNGuVaV0FGq1ixZSvH3Vtbne4r2mqI7pHL4PvfybvZ5xm9qGZoiy7hT/XwaIBEfB
g5aSMx+4UkoINRN4hU6wOpdeIexx0/uppuvS02j4YNFPyxoloyZ7IE5NdqYNtLT3
U1XUmmJZRHpeI9iIYL/E0zs1YPY3sQUkdTNy6xx3t8D2zvbEsTTaeoUWlelLAANQ
R6U19HjSxLxbfAuMklb7lSXFWnzAVhsX795s76TeAH2yM3sTickCB5addbynvoop
hHC7PaGojHXN3wmohUSqh5ruRBHe3LDzuyXXcbTxCDAEVXBqxM+JfTlanu1gAS9R
V/5jKhDEUYsXxnbObb60QqTHuxLWVHbe76xJGi4wqGEFrGVw1YjCdmhztzCBDBbm
I06Stya2xQgxgNIlJSo7gQyWKgcV5RqcX3QaYQy1gVYA4/PIMhkI0aCsKNoIC0K2
3dZNBtZ/Rra4RnVnS+NFN9pbiAE9Q6Tj5wnubrcEHMIIE72F41M4j8s5TmuJx1NO
gEcqd08q1QljfbRB2Cefls85uN9claO1g0SIZCQkJ5zBr3ie/BQRKJy4b+nCOemF
SfsJN9fBBb0pTPZZnlXQjefxpXqHvd5BE+ZsWFHeS0x28KhCiU58v4AdvjxI/563
/gyZrb0pYQUzZo0rD+RImp3l3JUHh4JNER4ATm4WXEsQtw5v3loBZA6bFIYHTzLC
dzEZwM1CIr043MtfG7X6VL5/Dx0zHjVZzyCEyDhvFLDiySFrbSCzGy8gUc497wu0
v76WoCXg7wF/XsY54FRhFkLW4aOqsDOn5T8DwNLpO+kpXjyVH+pUyl+OYxyGlMEa
bKbs3qDrcRkl6b8sKSRo4D4yNV1ho4mRuHmmJTnBnHTFB69SVUuM0GceZ0P+uWcf
ktN6+99evFm9PdNxLqBmWLt+km9d5lg2bHCPUn7o9d4PedAiX5MqVqZwVythhZow
CyqqZfE9AQt+BvZaw11pgGAcUw9pRCGmGvHLP1tcI9dUZdQNed8OJM9syu0TG2rf
465okCtTpUrGoS9hGT1ubuigl/xq+qrEX1YnaQwFBO3G1PAh6VG9YW+55Hxptc4Z
zYWKBQSKyKy/n9BqIJ+7TerjarbnLbZ9x5tLOPEuahEJV0Pl0XoZ9m5lqYkiuq0o
aghENdo9xUupvZPY0C4q+YDPTb+w0oFAz14TL1mfcH1NixPWSd/C8tNkroNbr82c
ow8qwWFaC572UusrH2brRYh8Dkv90ZPF+UMyRrS8J8E+pqfsv5Mte9CakBJhsBwU
pgLecIu4oPMtUiDqkgxSGZJItFfZmbnFJCVNrpneD3QIx4E3b3CUdxcUy/bWJT8X
hBVtgvoVlPu5Yp6jML5YDKqDwS3IiFJxUbEe++VV2SOPX4Ema3f7t+XxBOqbhdjb
hLUXBdh8uLz4CoRZXR8u9fv1CiAsKBp6bsYEx32PrEQ9j9snJIafGtSnum9mF6DI
p6T1rfdnbMr1M9nc4wcPuuAbFonW9z8hWOSvL3lTD/RAezHw+luImcfpvR5Jzq/U
9psO6KwuD8b/yeelWxm79A3Vzzqaujq9EG5ijw43PXO7f52qGgZozN4eW44fu7pz
XZnV3NigmntkkPGrQulEm6Ngi4vfyqR70XLrKLJ6mE2UhruulLx7Quu9mZoGwnH7
otKUrTHEQ3SjXYG7zTky4j1r4f4RWWxaPOL1zzDsXsiFVdOR97vqOlBrBSP40bvE
khJoFMMBFeWb0TH2pdD6G3ebj3Cjq+hAzstx15RkOh554rxN6kkkKf6Kyvatc8ai
vlIQaVe0VWRknIDUtR7H7FLKnpKRuIr96gvPvU2BskzjaFy1/l2Z2KeE1EO0YvqK
2sML2pioG9O6RQK66u16P6MTRRFjKfrrZEUkFWbOrXC/yUOd9cKX21Iu73xsm82r
XK1nLa7eoYeRx4YceYIbHx17T6qCluDz2YD0GCIU5uQ1jAcWlv552PQKapBvOop0
VgHDpruWkFQ3A29HNaiRTm2IlSPJz/sgVM2ssfgM5sELUxD/DH0JbhIUz+Ogn8ah
1A1NdCyVxy/LdFbJq7YQBnyVCR9AwugAsbJmOS3yixmsMYq7UlgozOHSLJ9yHnwE
X6sy1jVT/RcCWDHmcTCkixcGp2LZRQt05fF+TKMj1RM1Rss6XR12UDGLVzN2Vs9i
Tl1G9xMX5UndDW/8I2JH7C+lprc0lAKPoIB5MZ7pI5ftir5KFYi41k4WPOFZDlmU
no5IYX6409/pmpcyRhKt5vfXxGkyvIrbnknGku4WsMrIY9prFYP0UvvF7LPprAAG
3d6Ml7uh3sM0ZsN2AD45f9zd88g0k3S+WVGavHdos2Z+a4c0koNP6SyLakMDf8yT
pTfStmmWzlT4Wm3KErpZmdeiZPmSEAl7NT4BU/WywlcC7I0B7U1OGVBT8izP8kDM
f7AMQW2IrxnITxJNAzlw9ElGdOk6/ZMbSnQxKtn9NMzHn5OLqJj+uxOlxrVXi98s
FbYDww/bWzJquIH8Um1zT+GGOyXj2xRyCBYSa0ozTLMjkA0h8aIv8FSnINFes2xZ
/BompZi5SCti52KETe70HPz/wyHveDC2tKI1Yj1A9jODfpzsALLfzR09tnlACRgA
33g8AtRcqh01FcJ4Nm17QDwaVIxijC62stGe6LfkWXHe2Msu9+ehIaubWMFm7yKQ
rIDvjUkVvt/9dAkSmII+q0kK/52qllwEiu2Xzbgp+jP1xZx17mg1x6neU3qjOVew
gAJ30fEYyGVAUBjJ8Y3l8FtFxjNDP9vuZbe4h/lMaERSDSK+CoJXdTCcc6e+dvm1
DqPOzj2vWPU8dTAvJd5pXgrXOCk5GeReIMT/Jc1rEiFZRB9t2JBYekHrIHF8qiOH
ywwtjWbENpHjueQvC9/URwOWEh9BOm1o5siVMXyj8pEBWUkls8dF98MJfo39SADg
1ZtBVs0Jnfa5mtUmtq3SdQsZyStQx7JzJL19Uvjdk4xg8fS3RFkgIshUJ4PGUKST
LiSJ9VYMkWZKGgaya6qpK4d7K/lltkFXxcL6B49qG96bmNwwh862P2UM97Vs4ox5
cgsm+tmY7fYK6SvspqN7+AY0/Q61R5KUF+BUhhx8jD/DTWNT2x568+miWA/3rluW
hY6ODGgSHOGieuqjC47SraEQC8DvZ4LBaBmJvSP8E2AWk+JDBsH+LIKSYE8KW6PU
hz0eNX2nMgMdP562rX2T9OcUtwB2LYaXh6bsVmTR4b8KRe3X0nelhvx0anHLN66/
jSnD5aml3egzwegicjGf5J4Sb+h+mj/1I6zvK1u1c9Mia9vCxnZ/NB658FeX98vU
P7nr/M4GVKEu+OBOYr5pGfQlsYj5dEJ2zl2eqwWFNJ62DXwJpUe0+lNLnbj4e1bj
LLeFXHpkBcA5G7O+JpVAhpeRk3wPX8JA8rsEKGEYGTl0LjknjkU6Q0lu/S8ImJmU
UYgpQq/Od6Agt6K7YSezoVoA27skqiaYqcKy1M9T06yQM9Hc7Ol73EeXw20sNPn5
EoI+eYMiGoo4OBjEa9T0Go3cQIPLM6Vl1SouM5ysdfhjEX2GOk8sbav8MkORRuoy
8T6fzFQetni38Rx/OXSgjIAJaJDmTogDQTrl+XXgcVr+6L2DYlJ/dHKgZ06LJQWM
3lTuBsc2judeI+yEzxO2joe1cQwD2SVQQg/ssprd5xdvTAb6vR3OiuI5KaSMB1R0
5o0u/r6zC3EINVsSKHnbErGdX0UrI1TcKHKeA/iX1tZlZ/Mx+URMLxSz21hrW4YM
QKKuIZWkNIp8Rk5leBGeb4pWZ7TDz6hdpuDDSkjtcxEExqpzHrXQNfOj/Z3OctR7
QtXBN2Hn2DJd76u4Rt3Pk/iT4QtfMlFBHDs2nQ4OhzlmG+isS5Q9SsNB/1d3KVsO
bngJEIx8a/QdvNSHU+kLwLvl0Hb7iqi2exFo8IEj4Z+mRnG4Nc+SR20Mv742ti0/
jtRht+d+dL8WOBnu69Bpah3irfdZidhB/PX0t7W4W64xKPH9jIlWtSZbRudhhDp2
hXhwjrxw1dgCvFjEToykZXr9NUymWiLzEXtT3Gv7C1FKTIbNDEsLO2i4u9qp2gjD
n1nfUQ4XNxDAe8DTM9UaSi6b5gPubDk68Qw7BwekMc+EXh6I9HPCnzKdQ0WPeDDl
T+5uBTuS4QH5fdI9AWHeUqdRMV286gPnv+I8AWlMTCUeOjBwaBvDt2aduL7+/3YF
ljU2XiVvIK3ro4NfwVzVyxMGpG0F1todCJd+WX2G1vzRQ8LNGrRNhztIjhyNvA5H
OK0yOQ3il+yGn90KDILyjVP+tlK/g9kqw3arTJ9W/sFdTOfJcdy232BFzDtfrz+/
1AcRTAZv52bKRNTVm8Vchr1wwdhSsefahzakDfEEtkOvneZruhQMSLWR6cs6b1+n
5S31Ukc9j5rpBlJK9y2YtHHYD5F9ltHPppwCUEEBCWKBoV1PhHljEdOOOaSMmiT6
IPtnMF5sRuZNS3GcEI6eQf7uAcMwXZOA76AtBqJBkx68nWRWzNsD8qOgHhTCkcUn
RNe9t4hLDgQxjCY6W6P6gdMkLqDMFDDMBpIptKOfW6riE1MBVQl82DwpXK58Dnwu
JhGRH779juaV5oMybwZ2C5TXb1x5boHijw0JZ6oXWSmtlCNi4Lc0ND4WOr6oKA+m
yUJuaiC+hQl3hoxX0vgmLKuQ7V96T9taWG3Jr2xoZ/AxWoyGGfSCEeo6CIyyfgDM
/kV7jqhHPf3KAaawjNz0JS3Mxqsn+TsYyuEEgB00ibo7WRyzX1H7hkHFIqPs59sH
cIKCV/44wS16RCrwv7pmW2QEAktBFsjoXLwUoIU0+4NfUm7L/vQ3uFwxlUsJOgMl
9HJhFaTFzbRdpphMWTnG4kDiPa7Hx21p85Rf3QW9od0=
`protect END_PROTECTED
