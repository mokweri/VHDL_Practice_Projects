`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLQnsOjbiI7dtBnIxiKZEDNje+WdQu34Gl95e4sROo+G5U3gu+xHUGyfLjgc76KX
2MMRkcURd1IPT9trH4I21tTF79mpa6KX96spC6eFLqGZ0o98ZkuYw5qBSkZC+xvJ
uA443WFlxeY6XuqamSdq2g5f/Hi+m88/LMO8TOoqIJfNzFyE9dTm3k3MFlOu80lz
soSrFOOKb88BXRlBQmThYKDo+Y6h8SqDLe7GmQppaU50SOiCWCSCbhho4oVEGVHg
x0SlxwsDzVHFfdPaOWYaRPvt4XJY93r911nM8KfBf8dGIgCCWdI6PlGn/01PH5fM
oEByPvPaKmVvjtFqXzDoqLaYEWA0iKF+0EyrsaOljopz4Oi+E6H36c5shfRxDikn
8U4qIyr1LBUdGrFn3R/tsFinSHpa4Sw6Sg3zA5ZKaws5xCuUKHmjjKwaQW5Ax2I8
w7AT7WpUC/tlpgasfxvlSryhCOhgYZJeWtA497cZubqgOuhFxZGQiobc2kOLzQ2p
OPtWd4I8nxsjgXhP8ljz0bx/uW8ypuOAlfA4NmlymprE4MSAEv+Dmxp5EB297SCL
Z69QgNajibrNMVyI8k7Vf9sipeZ1J0yY0w81FWBTNTWTELRrPOwhotJ0ZMGlRA5F
uVjQV0zfCzmr6T5duRa/VNNwHz93xwThgyR+S2Lv94sUxsbQUPFmcCKy2XhMzDiz
dbmjRfHVzEwTNR/vP++68EgU+tvfpgBgTXXjmp4nAGO1Lc+P825pbclJNKpL/WsC
4Z0QGA7P5XPEMJUuNeFmAfU3DjSv6vpbqZY7bnGaJsIwABc9VQDbxywfkTmP8jMj
H/HLnEy6cfg8LsTcl1DU+TlCNjd5Sc50g6SUA5ckSZH5P1btjCf+OFURwLuXCYXJ
u81yOQ6mP2tLqCbv5301Lf0IIjXOyk2A7WZLhiZzTAx23PqkX/XyNnBkok1Asdd3
qGhTyYSG3JeyvlZRQpG8bVEnR+sNuSDG/sgSeoSTAy7Kd+aJMFe67WoDpskasDMr
FWvAveh4bb8vrMLpqm6l7QscNMYMGsgGTaYllUl0UuWF6LZr2pn/d/nEJM9Fh9ZF
4EDOcoFt3vy1X1FWSxkVGdgKOBDz3QlKsvbkqKGTPQp6WA92QO3c7y+uVhN1/9Xg
X1KBZvDYBtqwKymrh5t7yM494n8hYRApZtKUpGnjWlYwCitysfzrEFSi+AnRCQQp
VrkTLw55bNlLaQbZbEg1cNf8IxTOT3ok3DXkW/KuqTriGEbqd81bZLV5DaFUewCv
hr4hC388ffDg0S5+HOpS16PRyMk5ehE68MocjP9T+1nOuPVuJErjp12bn/PsePYa
Yk92v/4zShhd3K3DcO+BvO1rQi8o8zymRt86MXG5onHJT9FJp2oahdraeTCZGu/X
F3BzDOpUN1u4dX/OhTZ4bYW+D7e6epWTUqYAEkBjQsGapThrEqb7jOoIb6ZEv5kl
RhJA+VR2lFq0AbC9najO4Myw50dDwP8PUUh1Im+p9CKppc2RsBoY5idF2zAUAL9P
iqgXOG7rTgQd+saMXSkx2frTSzJDxzqTODAn0ZMnHN8wGxWCPtLi6EQ5QLvNegct
`protect END_PROTECTED
