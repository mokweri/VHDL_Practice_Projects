`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MgEgboe6HyQle8jbyWbsMhNujD8tKl5W8CBJCnpEDu/BW5WniiUpb3doWa+mLyLn
3Zw4F2loEIdNC5y7nh8+5IdgTI699DsXwybSwYPWuG5PeS5JwYvOR2mH8FE9tzIa
kAYpdYFMl2YIRnXvjJINoj+o5jrHNR5hDIexD4OPIFnfBWUoAjTcTUJysS+jnzqu
x7MYsHz9o79q8bOvgiA8sYBJp3zJ0uAun5blHwAAnwa54eofc4Mjyl3NzjMBAFdk
+77ABGUtxIVcuhh7Fg/y4nEi1PhJAbUg2hvVdQTkrBqmvPErvkdLy8Ojik0zpb8p
kksu0f+MmhEOvjqfiE8MVeTfD5WzbHIBjAbF3aPX+G2hN8a40SSbWV01T3ClC+dp
cvEp3oFijg7V/8w9EmZQ2ReDVFOuLBNWlv6QbxV3h3d1tSTJtv2JT0BXccj6PWqD
T1KfcOAKr7uqtW/ONWa/XTf6TYoYVp4wPcranOrb6XdvF6cFweDQxdVP+sj7G/uW
MtyHmXRd0eV4UORA7CnsFHLQ3EEMfXgVYxl2JaxZ6rY6HNW/joAfxCSeyWfHkTgQ
Wqkay1fS5qoov0ama13dysrCwPURuSn8VyKvcYAWDrmvUjKb6LqruBFP9wkaWbM4
mG69/pTwlem4CzY1eSARhgUJRU4ZMuFXrPq52aH8Iu6v9/p4fSeXruTJtxyZT/qi
QkeTuC0JH/n3+q3yx/9J6ktXoNEmsoUa9aZdVPcFMIy57X80J0N/g925+ZCGreeh
j4NfP+5k3mbslxpcMnTFtKAT5qWG6voeKi53Wv3VJb3/zH1tn3XRlAW0Rl0H1XI0
cwX6C7UnnVWzm/3GYxViqJ54AThirK2uy/loQYeVqWBHVJlvbRP/d+g2ifYfJlyr
MQ7eaPcs5c6ww8TIYrh3DnCHADb/WTEG4seU27ow3hDULdygZNedSzgKR5ifOkTk
oB5TXsDweBf9E7VGViJAIIqLdacN6dpIBZz53PDHD6g57TbvGW3iYm1vyCpHWwFY
M+2zKvmDD9+ad4zroGOmszoYFf7SLPHl0g2M51Zi+BRyBD9dBHecchLQAbRKr4bQ
mfj+Pc5p/opW7g954g2r0+d98EwYJdGY54hd7OlSnojzWu964i4bWYs3NOhkbM8N
Y899kDtEqXgoqBfDooCr7UEnIbX8SSoX/AJImyOw/Rc3a6FG0yuSj9Nr+yGf0mpU
M1SoUdsGN/D3x/rQxpeSv1wH25+ouv3+Rd3gMPoGB0bKFc89hwEnnnxFNjv2NgUa
pk3knDRnx7fOU6YtNoBYRX1ZxnRu7Xtuxfgj2/ur4yFEK1Wrhzs03f7qus/KJMef
oQ933vITlllW5RT1s9ab8urP8eLz04Wb8Ad6gsRZkZMCUjcX4ZMQcfDgcTBZHEXX
17Muq2pIJlx/UeUnjpWZAGbv1Iv/S9z+34y8ZGWaMfYN8B3j+XZyay2vDpLCByGn
kP+FtLDGUUpzy136jY8RLXfRJDeYA2Y2l/2i5MfMzH/ssV/AfA328xUqGAot4bpm
ZIfvBNY8fnAB9UXSPowiXVysze/osQo4pyPkKJfRPwC5I6knBl6Ovw07ZsNXmqLt
rrasSUBGgcnZlgMmU+vgdNbLjnF/d/yvMW+Ozd+N3UJdyqoFLGrqTYpLmxPfa8Io
IjedAySTFt/Rh+cwDJuI2Y9RaM78e2nUBy3upgtbDBBzK0H08JQJjMfBHJUVT+PY
nmE4uRzEFiVRrWHqqsRJ4v2rSbqH/97OecvXMO2NrTEzmvIBx3W41qQ6pG9E8Cna
EKurds0b9T1GtvrqC8TQ4V5pq0b6kbXjlQLMZyuXCyeOIhRTrHvQ7y+hBrd9Mquy
a79qptgPNfdsllWhc7o/R0skWQj3IrUPAjXMOPZn1pkstfHVcch7b2HeftLoFWpY
1EXtesv4q/q9qXxtakHLTKCxEQ9o5+cacUsclSymvDtFgx3mpk0MiB4SqBhU/Mnk
32acCGUMPln6gfOwztUrYGYMoeYtEzxbcm+92Y0vBX7WopJc2kfdRBJXFC0dY59x
O3Uyq5iyZUiZn8/17TQw/doAmrjcN7Ix2zSVJ6SjqAa+r9OaedJU9MmdOiqWGcYI
k4Yj1+DoIhsAw6cz8UcVZNo9DCHQaVFkgXONglNsVrQ06D8e6L6Q9xA9B6Dkh/G3
jkzOHUatE4tQwcbSkQNz9OjHOgSFXoGceH7y6B2ftRbzvYLIQEP306oCSFmi62t7
dR7xioDcjjCOszS6vPo7H06Ym5vOLf2kt7qc5RO1swHb4zuDlNaDoS2N3NzYaPiP
fqLNm3UrNzUj7jZRILc2iIieozqrvQSAKmgL6VurPFMKliiTsvnvtjg1oqfUUcuU
U0pAL9QzaqWDUkKsJ/eJdnwZwQ53g7+b+nLQG7XmtCUOKj4zShKqxz5JxlfFszGM
7kK7WcGup5FFq0yiEly+as8wr+2LeLBXhiQDdfdAo3097VgYGR5GhvJQwQLsKyw5
3SJwAWtIF22NjHRvYGXWyXqGDl4NnAYl7Cpe1KzeyaXF66l2r1N4pDb8T1JaqjMv
GCMYq1u4n3E6e29Qm3nEgjuoI9HtnH7UmoIPTpQlJ9qeiu0wrvDIxtRgrAAa7MYr
f/AFliWx7Gl3RdxVD9W1lQ6LvcILw2kVhAwday6uVBX8zR1xR+mBOWsI7WD0GQN2
`protect END_PROTECTED
