`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8z02RLybCE/dQqbsJmvOKlana19mMId6rqPLknOPyxIXIlLVv4+wJWSvm3LNOGk
8EOxCi2wyBn0TCOlNpA9bAvvwUovbSMVEf+CPRQOfrMYAiRinOAHWyGh8td4ve2z
iOHBjcNAqAXgJqg+0ZUIRTyK+zMi8Epr8XT8J5UJIuvswnUShtiIbSPxrERgwUvB
T7ByDRs1y9zj3U7OhSJfxHGnumOBx91Z11iLI5OpNf4QwpsR94jMHpzEU/1O5bhD
uT2xWytY+Oh85UQGvgPtHji+YYSH/8iecDI4BrXzdhxj8is7BgE+m/zjrDbqq8O4
TI2JuTJAcf+lBHg5LpZ6+OF8/2PvkDZfR9/AyfDfsjRBzJ34MUxaRqU3RCYAn6BG
IAb1FejYqvoVu0ZyoT3gdbnjBZlW/AEA+T6KC2zFCPg1LZ/RaYCpS00/OVwynd8p
pps/jXXBaYUeEeZQ9m/9rteZkVau+i4voBgOBC2y0LzES7UJNDwa6Z5CHOABzg3j
ZBV53nEyWtKFvY+JBQwdYahG8A5JKHZN27WLwCsqnajkh99+gD9KR99fqQKz6q+K
Hb8cuUu35GPcDy3PlXul1DpF6woAD8xULZEjvJcvSgU6DDD07tmHcH7yjpCNwMxJ
GVFj52XIzNk4ALX5eADTW45T12ZIqPtWGmxaHMvRRVeMSsB+uXLJh9UCm1LV0+eG
2pFK+j2FPVbSNon+Zj+h1p+jPMr8nd/BIut0MjUbm/crmNhcq4rKINOz3GYVxnkX
hhR4PjZ1Fy41iREG5dvjJDPEnHnziHcla5tdwBQ7dbLUMLih/JGg9C4YaYf5VCEx
kFXf0pHxtzPFWoI98kC8I6G4v7qJ5CaXwqQ2p4o02+rsJDRtVcnRSrZETM1L1kQ4
2QSN6LrY2TQim0IwYeiwieuBLmMdJ8gmhk7L4fLnViYc5R7TZDIvWXE+WTMDN8Be
Xf+kaQbouw2sqkxUuRazUoEk0GGA0F5rXFBy28t3cngBJASHLrKQC9YiAgmwKvfh
khR8dV8mPNloetHst3nUWw==
`protect END_PROTECTED
