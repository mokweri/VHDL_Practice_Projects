`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+vb09jqbMbV6OwELIys9pzQ6A571SCjZJ9Ti+hJlYUyAHBzsjunQadBxvxtgKBc
l2pXQX567cDNweHy2vQsG5ne3gK6Sr0hgVwsGt964Qu2nh68S5vQxHGfKQQXxCep
DGAuG/9kzuA/2TnlCAzLr6tS4jDMG12K/bdJtrF2m4mKMMV363I0bLuGAGjUzI1M
YoIoxMMvE69wKyHKUYWg0Jbq98tymGNn1ekB5OefqNkM0I4+8XTLnEj2a0afis83
U2vTuUT8wCJtabwJ2FPCjoZDBs5g71lIRYnRytvcdIsFNjKFNPmUPrVUH2xXn9i2
QCzzRC0g7Cs10rQnr88pTvPZKuiHvT//77OrhIHJZFKA19xZy/eb/Zi4FdF85GOT
Nzuwrt03T44b7m4lbsqjk9LKUCOmElxQtjOaPdB/dNQZViwXMdnLHJ0W6kDMf7Fy
ToNGbBDqNqQ2YAqrSpFvkg3AHyXDA9MdKFqqIr8U/GZeBc14ytGAjHTX1qp8LNvL
kv2Smx0jp35MMjlHBTVTlUHAbKP/A1kyqLEnRfuR8CdC/hO4nyPQQ6G7NznuVHQD
3lDfODa1ENivc3f1IVujyh7TzLJwfCFIesXvDPf/LZUAyr0xwLprww7PuNK1rR85
EQ4wvaKt+81TAtCvmKojKaz0r39j/BOXh1ybxc0y920+Trw0TLa06WSLAXLd9JwC
PVO4diD933DfbtCxA9bQL+H+14gIo2R92RAcwhZ6Mk2/ceG54rKNdWmqEy4Y/yLc
UZdJzHg/yVdR74Ma3StCEuEqywBUILPowY52JZzmnnNUYSFVNlBxo/A670d7l3TC
/9X32yX6Mu11uPhq6mRUVJulcxxbhv0gE1QNFZigqttGSyntyjxhNB4+Joco4GEa
aOCE5MuEhvHOKrIt3HgYLJXlkveGd+SJ15D3Ivp01SoHBC2HIxBN5ozLSBO5Qmmt
ksPKZ5QMf+1BIuqv6e0uo7c+DK7KtQgbamxmRLmR2199T2wsMBboskRahquNkq3h
tLMW5mTpAsQyZrbxYAr8uP86WNx/KvpeyV2dCCr0zFeKtSrUoUoqQJNhPsC1+h4Z
h9GdR++gz1SXtr8kJFLWmeBPiEU4pbQ/YbXpxGaTSIkJ5zZUvfMG2clRO+a6Alsl
BZrrWgnG1yIxl0q9Dmn6YtKrYhVuVxgZCCSabsSUFAaDb8U9O9uQsZTa8ThEE0Pu
XILegInW/WB8tTSm3egmGqZZ3LY0w6Y+Dx5KQe8Q54NBrpzorKAmD09z3MokYoyR
VvgtI+8BAqLEUsV52demUFPMSs4fdXE9MOADzg3xSPfS8w8rk8nTNHVvo2iR5zu4
VMdK4DbhRLUyWw40n0bXqnqMoh9AfxXsMVYaP0ucfux3PcLszocYd40QOqx1LCXB
1HDQLs7iK4RgrxeXykuhk3c0YUnlOVr3EbU6jtaoJA/3GYN73+L5g6FkQtVqOart
hgGbYkxh0R8+2PVxwLfeARQbRHk/tCAcUhe8l5gF+pE0g/Sdpl7cbhT5Vl4qSHFM
OEMqi/KGAAk+894CUp7/JRih2U1gUF0ZFfQyb5T6bUx6chmwRvCi42VCh3ejoPqr
3LnwIaZsEXVQI9+KlH/RFsw3kknMNa70ysYxfagkxrnvuhmKDbo9T49DKOrvv3+u
9aLdHjodzyyzTqc7gNhgsEkeoCQ+lJPNFd8VDRYeAFEQMMEoMl/1mDqHF/sLshoB
qO5NNRntqllUAZ/WiyzfRZHEaShqENqVuqaepZ9QdDranegWYUViVfhNCO7CZsFF
xbU/Zt7GzyUtitkHYOuVg0xd+L17zMxiTmkdFA9h11czNTJTXmiL9NdoI5hC2F8G
D5v0ZL5CJiM4znU4mVduc3N/9wAUOQWtCjgDARcUhalfisWK38daobYojhsJjHaS
sbtWWI9PTTwxmjajZsst7frKs7z87B5R/922lB+AfiDofzeOPfUxMdpiAd1Hg2X8
KhPiNASVBdcF2NktUhpfvuiNWb0SridCkX6E6eiEw/WWesCvyrPVzvLsMh1O8Saz
sE7BS7pPZgtfgB5Xy6xS5IFYPZfvk64M6CjZPECzvabRXbaccVR1qJeqDoX9U/g8
EoC2gfMM9wsUSNSwpfRjwBeYi7m9XU+wGcHhDxG/LAMTgZKfsKctA2aYF6pqQOv9
Xd8HgNaIFVk0M1G6lcRZ2wjG0Fwc6rRHfNoFOUVm4boqLF7kVvvQGXP4QBQZ1KWy
p3rfudeQsmtM2ppCM3YP+qhxqaabZU5Aa9IM9JS4Yd4+NvC5tcUEmO1pzN1P78jr
Tv86hyz6koyyEkLov2BGzK4dOVokZHD0bIUxr28ABIV3Qxt8+1TpW0KHN9gP8OZQ
rePOsFiDcKGwu2L66rmyuoUbND4qjEGtvGWQcuptM4P1SNnUlRU2cljVnyRvf+gl
H8clUxGkbeiyG327tIDQmOOu2LW+rq0BsOpXxLtuiWN9vDdnlU8Au7NtnsZf3Ud1
bPHS6L0RiA9gC8IGavnkE6oPKhB0Z7gxYDjjbu5djOsqXcF/t7qd9Ll7wOY5WuVP
DKzH5QR4zxjMyvTqOZLR0E7pZRmBn1MyUyfyMbqhMXmdVMIJ8UZW40BBprDuW63F
hDKxHv5IoBZ/UtH/Z5iYcLA8NNRcJ7YtF+70mAyIFErmrHweFZWjGBZ/Nyn2xa73
1rJlX9ISZW6g4AKYk5UJiunlmZb5JVzcHbIekB+whz54l5KSu8j55r/Lxg+Sw7UF
vL2XU94IFB4JXeSq5AWLGmjh6ZZfljHKAI0BkawluyIBz6onuvrKEC/MCghmLu8u
r/kagmycjJXMW5fREG33HUtnOjc+PPqlN0L072mHfkqVh6CznM8OnnZ/p1Eg7PWY
lJw8it5JGqAF6rbSkDYuT4xihxMcgA8FiFocUR7NSziZXMXq1XtPsu0VcLAF9ixz
jZ9BpK+3kfJRVHoRcU2xpLPKBkFoj3F8X2sOi8+DHSUyIa88SJvg811dNk8OJzeo
7BW5MwJInqM+Q5htuFQ8TMkffwUXxMa0dS6nIc3BxWi2m1yXvNd5TvRJmCCpofFD
AXP01bKsWnS4u2WG9InHaXSxHajapQ4N00Y87nOI2JJK7b2bEsocAN9R4YGRmnGR
TMWkMSS0a8WuA55afwX95Be4uU28GGP2WDBraIubCnnXCsJW/p+VuvxBEOioYXmL
YG5xMgZsuQ/DpGUgLZopF7LzRHRDr5y7EQKvDbzXAlsuenmIvJQbOTqnT6e5L2AS
Mn5+r/2aJBtsmwixZJNYOoHfEtN5oABmICudHDHGqJw8DLchkkVIUbUZuNLsxO0h
uh1zw6HTjiUP4F95B26ljC+PtnQVbvcoINZsXLosYb8aO5YmROzEr7//JBTK+Yjk
XP7N9T5Q7DNccgOqVjw1X0yq1oF+q5/QBHyCOWbmw2YSLB02nIKPAHMf5xpK2OMl
uLtcMTz5ckr4Nw2P62v8FjfPMT5h5pj87iREnmp0aRuF8Bs0Wqs/t0M0LPyDGpdC
BPRDOWNlXXiunkmkOwpfqyESsUkq/V6EcVKSOzStPFsRvZAY5RKhzsmO2K0JwpwA
vK8l7ZGsFRrodUVs/txhD2pgick3Gw6hFkbIlMMX2dlghuEbaNcPD1YuansWO/1d
m1OuqyaFOHqsIJ4i8t5TgN44PSymsZZR8Xo+CKtplcTwTPhQGHNac0QXZwd2SuJe
cK1A+Esqy+MUKEbAwtpVGQ==
`protect END_PROTECTED
