`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LACUA8MKdbK3u7lBJzVjbR413DMZUoQ8wnmalBwzA1B2jiJ/vOeT9l6aw4jOZ2jl
Pdx1L7oi4SiG932oDfd2pTNnvlmAalyu4Wxhf0vZojsy2/dCt+aaGd5Xdxog+hRz
0ouiyT7hAGIMUxN+66qSPHbTNmNtGWhsUrShCI8j9vBBFedBt9IckFweIqKlrjes
/wmEDlJHqir4Svff8EaH/mT1NrFb57fNRvHN7CoBJGyOq/82OUOQ5SJ7aWuBocYO
HOMDAZvEDYaOJv8TQ3WHiWNa3JSwfkP1kSdg5boRLgUbnE+OFdfrcYv2/c3j07lX
c9np8oTzWz63W+03K8i0w9Deq1sPaB2hY9SVUGWe0o3FnIU0m2R3Ys1lc+XSkwCx
TZcPmuxLYcIYW1MrRGej/LaSHKISsjPxyeyTNtif1OCrm4NkrH4Qdwpqps7H5jPh
wN7QSKibmKaTx8kriW4ewoBaEO7SrUww1ikQeINZWDsP4bqwlL5qwIP8mwNyhWbN
QIHUhXv5uTmK72c8ZhXNY/0uZMO/IpmA+2FIwWroJL+OFBSN9mf3lBHtsv+9HLoV
WHQdwFSsQEJRER1523rEl6PUcm8qG75YXXagPS7MDs5Zpyn8WnNunHyMUwvcogkt
8OYzftKJPCoWZamO351HsIIxvv+JNPMvj4x7uWI9fE3UHls48qEGh+kTCV+yKZl1
xjnbe2SxBK6B4aDb6v15CZ/FHFpzh8EMuFYKMeIA8p72f0nr4d8lvvglq8ud2P9r
vheQqtlp/Xr7ltftbamCFGBfrbw9bd+CoFQhXwznHCv8cUWHI7P4xRc9gJzAKNoy
/KbT53QrZ6ttGXx+je32/wRqXuWbUi/6w2tOp+ZrbNg7ODINC9cKpDK1x2AeuQnd
OpEhBE9Bm2Mlt/V86FA8eWipopScJDUpY9pc6bXvTAM=
`protect END_PROTECTED
