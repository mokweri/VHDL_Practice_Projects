`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdCgHExPTpJiiHKotaWatnJ31NaMoEmAqdtlio8RkmC6s98aObGCU8wXftWnt+/J
dPPnjmrxIdsFAc4betNCP5iPrkJckiH5pY78FH2ekfSL43mtajYxRtxc4JbO3ckz
em78npyInL26f3kMIInwJ9vRBXGOMy9hTA2elVvzlKCOjs93tm4r2GaDN//8dPak
TtnhD8mkHFz6SQqAE9mexKnC/FBpbF5tyEAnxhzcXWufX9NHYU3NEYqFQJZImUuT
73UvraZJvcP4ERNnLJvbqIa7E0r+oHMuMsQICVpsqGzjdf4HtoJrkt7UI64YHjHU
czSEZ9Yh5BUDg5/o7Ki6gD8ch8njGFob62b/Kf3agPU=
`protect END_PROTECTED
