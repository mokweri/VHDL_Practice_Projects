`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vEIF8g9yZAXObcElpI+BwEfBamBtANHp17osvFX+gz3UExbPwz3JUnhptQDgntC
K5oyZO086Jb/4M5qn7T8epHg5JzmllFNGBfpcCpgOmdgUKFzFPcIxSyyMNyD89+O
DIdePtOZuYuRF4+xpQ2HqhjnuFr+3/Ri8cMVCt4bZslQzMo/OFYuSC/tYd2i3LLF
NPguktTEeXp2cX5tH2x2TLlogQG4NIAS0hWRkQTm3lpDDAX/yF6Z2IlaqVgPfqP0
tc/t3qtTnBEN8GO/QvW4Pp5aiTJbCTCLNDcJ2ZCnAcdyqy5BxFKRv0W3oqsnqXtw
4432NGqIxGzfWSoLM1ovyJ4btyY62wEoiCl05sX7TpeG5MMyKvaHXu9VsXujjiL5
rPgPqZ/mJfhc3sWtEks+nghgcFWy2YDTgtsTFLGGeGdb21VhPY1URmyA5HtrhZ0u
LBX+PKyI6zO/9mA+ylQDEi/uaP9rmh+FPOQqsVjFzX4=
`protect END_PROTECTED
