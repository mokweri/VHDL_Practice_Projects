`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvJY1fm28tHQM7pEHJJDl6SPA4wzfQvV13bLvgiP/XvzOV83lM+JTd6TO0a2dQUQ
RWHaXgHmtVAmfc1imq5Bs5Dad8PkS0WHBvoPHUdT3QGP17yFFpKf/MG0cNLlzQC5
BhnWv4A7U/atM4Qw0X99PglLbHTcifIk1c9tW6z9c25MYa1MrDJuQg3LBDJDyZ6T
BT+lOdHDoo8wRnbq3XerAgBb+HlICF6EvENfFcVIaEAjc35W0wfk0G2mhHidLDi6
GhHityJKHDI2khX3fT7UEU2EYR9OxuZRhTKwdWQCTMNnmJgI5fGIVhwe9cPeDJFS
7pRgEGn0LVotZNahCZA5yx/UMOiuvry008pGxy9wLDOBEkS9w+tPi2rlRivNfWXz
MNNbrArSu5X78W21FKnRCjwb8nbfhlAeXfc2VSX5u9WqZUT4Wl6+EB8QcijJXQbw
ISAQWlFyQAU3q4/LUT89zXaYGZOf6Fc7ZHVwsEurknRJaf1xbiGnA5kc5wWUa6Pc
IncBeRZHBm0t9bNps7Nts0uhi/AIVpw8uyCgosoIGGLRytHXpXMRcZB4gC1ipMRD
HfvSlJQPiOYD0xx4j8KBdp8FTaOhDJFUDT4/K6h98D5tGsC0x0svFBKh191GlFp4
ex9YeC6ywpwZ4NBi03FOCXO6Ho2HIrVIb4XUTiuAI01ZGYENJullsFoDw1VZ/qgc
CctjhpASaRiFBGWfNdHZK8SBJ4YigSlhiz6G6duuA9zJFOhgxcLxsZ6rot5oFNXU
qRhgMmjEeftY4uMEQkphGwNoCts8bJwMcyMl3WCthAkjP1jGHS24KvPX9YJlf3OV
NI+hKILk43GUWDaPGoOrROR3UZ8CMAoSXBZS/+cwufX3XTfn3zcx1XYI40+QazjP
XGbAUWTxOkTn4Dxk7mWazTx5CL0q4nHTa+/XdNtf6mOTTqYpD11tTTXBoiTBRVul
3iHhz/O3YhTfIcEh+gW2PC8pC6DjF73UFpCwUXLwcdWKg/YaK2HVcoE68Lpjxbvw
0DmKqFtvXxvEX93k3boukJwrJiTIyY2NXeBwYJWbSINUepbSQ874xx23I3v6p1P/
ykXK0T0Gb3Gw+3xuKgT23g45CxvbAGSgirYpQOfBqoLSnUCMYGvDjks8to1uqmTl
bkr7nJ+yY4r8DNexkLfykYGyEfXx46fJFStBx1VNIVfSE1oTCEQ60VCsWKmeaOfi
teSyp8zFR6Vae9xT5SCXhCjjPoa6bF1jBNfwyBy3xHZYCW9CMzRp+c+O4I3d9hfy
JApfJqnWt/zUQ2MJoSHLQjVYYCX2uuqrHrxfJJgQgqkTdIn5KKgcumsHS0obn6A3
3/LsAt97QcA+9yGKlITJIA0frXhktaXwmN0oemP+ZjU3tox+c+LpWyV9bnn/gwGX
olnpvmK4R/qqFVy8u62WfmkTE6DQSGlbM9N39OL8vyEhJij+AlTMFIUN/nexUeBd
k47Wx/qiF1G7DSY25fpnYwt/S4apR0JsI8CFO8wvOSjLDjP598L+tZBLnSQEqYzk
z389ylODHznekltby6R6Ej7hM/mvnxpmxj2EWoNVOqCbOelX/h4LOIhjW9NLfyr7
8DQ3bV/ZUIIoBSDqd6LcB3rYQkehjjrmoz5N9kOdEkOBqfloAc/5id77Ruik51lw
sh3VoYS2KJgR4viu0RlzzxAR3Qxf8rvzSsGQLvjde7VRJjtZzVwHF6CtDUfvoa7O
zHFcai+UnQnUu7fR1nWum9F72vh2/1SmRfgWrgi3CcQ+X+GhwjSX+Q86VMxl2BHL
f4f4M0kzmx7j1qbGBlCIHfK6uc5rT9dwSUX0zPi5hizbaVCF6BvX/SWg7OnWO0pq
ciqkJC5aszVIsjH+UVzu55psxYTG3Kzs1FJwNdOxGk3EPKLUyeaQa6jfiiE7lcKJ
tS6adB30wbMBYSmgYL1tk8sWWJwQEQlslHCVMO+gFTtsnWnlL9BDKGLCQN1LWu5s
Co2t5FXcbzITNfiEvOjiWRupYdj3/tn5ciZilbtMSbhID8xOBfLU922mGZ60joee
OH11JA+IhopHmCltiO7WYmficRwjW8VPJw4J8Hz/7q3sFf5R0xfi6AWQxxmnxAD3
UURUQSTspFn0tv4Gyjb7PS+zMzTVqXXsime7uxCd26Uw2OEJXK2EuYf4oZ+y1XQB
5GJz8W0RtaWmRiA1CazRSRpM3JM9gIY+uhFpA3DTm0oYrrodYhbpVzeRvj0D39pq
+u8YMxflQWNCUsJDVIUGpp3pznSq2MSZEu8ouAjVZfBbHYjsVqJM0ioPNbLEC99k
2dXd4Jw7iOBSZaKZLNhwOnQ/cy32cqzaZK+67jEb9bJQpCpMPCDgQDV/kYHbR5b1
gs1UeZgEZslB6X/Pvklnn11V8T9sT8DvK6kNkwTpGjYV4usYN8oKmNTlBSvYM1bF
+3WrQ/YK1fAHdw+Jozldy6ouER3vmMVxBbdwpOTD8GiiZ19haetrolSzTxBlUha3
2TTh7jzOo9DcDh9I/04vpugmR+0AcL0c4jGP/k+oMXfnZhxUKRQ2/oxslhRaQtyZ
lbFt2U8Sm+sY8VKrCOxpAuJX3eZUlUefTLGa5M9PlkceByQsSw4F/e+PiKt8bxY1
ZTs9moAWwhOBwmRAs+SGOf4k0HBMk5OsxX5NxmZYkBy0D1qJZa/dEnq6y4nGJNvz
GLTrpVXOZDrSupQAhcwZE37K9H7xGXEA26gEt1mEkISEd+3aiSsXSSBbRlG0cJjk
LQJuU/b+kDa/IQCA4x3HBhnzEr6mQJ+4uTSWbq0eTx5a2M+DFV+fTcig6wJmYmsA
TRcg4Li17btSlvjQ9ZurwtYRyX/aHvuzvPa1KqzZpqyBbPTNsZ71i+PXTa+GdSJK
OTadfkXWzk6l3e5jVbe764vdLyTbum5LbVVNHkeDQ4/9YRXCy7uiIBeKCd3gYi2H
jeJs+vEj5zFql3OlrhR2E6uNGkJhgH8zUDQtgi6mWq+VS1jJj2+nncdRPsFCMxNU
893dOsK7f9tMSw/P3aJ+gsiphYj+g3H7I9y67iHbP+KClhwkHeNA/Q8wvFhO87Dy
Fn5CDBCE1EARxQlcb5MSV4LCzSFIyTPbzHUuFdZCl8W1OZTJ/J7clQKSAS0ve7us
E5VWgYEtbgtVVsfCrUFbl8b4SsNj3UehaXz045pvbzlO6UOW+dnEH98G5We3pcWl
uuC5gqmVsHnKgh+hLD064qTYFC18bdux1M0U5diQsKIjiBCsPE0TnGy+/NY7PL/J
DWGEQ/1Fio4oHg+J/qlDi3cf3R9AGPf78hqQaBUKvBQow4pyQPqQUbnBQG/pHPS1
WyvL7iVZCXEFAiUcn3AajYZSPqTaPHnGZXUt0o98wnkQp/k83XY4i0QKDx8D14fz
EuELbVLAlDQjgrbnr0LdOVV9pN7cleBviy66bVcUmeJuDirvrAtSK7CHZ+JLqw0/
sn/g9Fw1Mi433uPpIhMD8qSxlfnYWpPVkAAyCc7JvnpqTelTFugTRH4d2WEukU/m
H9HGIgwRpN4n2rJcAU6k+b7PmZ6dEe4F6dgVuwE3sMyJSsNEv664JEPNfowLgGR6
ARJxF5WdkNqMPtpVKZ47IjYpIgtW4JYPe3bncIMIIqZf8+Jq9BZx7lFUssc20Mdk
nX/jq0XUoAC9BcLenZvbpte3GvsKUjEMWUzhinx70ZZRja6x6fSvKITqgUmnYYxO
pZ3zCPXPM6tCzQ0JKHcWI7wF04lpcOFeQ8GEeWDpfsPqEL0G+VNVm0fO+8jC70MG
x893IIUe1vZsI4T6dwpmQ/ijWlqX1xz1qgMrWNgNpOA/4Yj0wcqUMgJckxtOiuXe
/9HzcKhRRsKmaFC8RlCly1Epcm5AqRh8RrQ34dTTuQa5eplZtWq6AJrpiaR8x18N
8u41H8Z1Z5RqfJRMGnOedgAGblvEjngUbFrX+Ca3LZMG/MKJfdWSmux5eLdb7Pj+
jgZX25GCZzCw1GWxI+tVF2R57/ns5a6ePWOTIvAgN9nP7x+f5tEVKFwRfUoX+xLr
J2WyO5Nd00DpNfq2DGn7CKZjinkxd2T+8RWBwiLA9gvJQINbC0XZkc8OveuIkHYw
HKcuqNoHfjLx5HjUTKJOcV1WE/bqgfsDvGfrz8bf37AmCvZMHcKhYYPSzwVupDrG
qbDL9jfZSFjtwtk+eb6yAJUckTeVQr9HvM3kGy+yIoBblFWNKOJINHBhbzVcJf3+
U6bNND+LfwzqBQLy8BfDWzmYbsW5EO1NpY8966n2RqoDurUO+etyAF8vIBX6wzrU
X0qx3Ah0NFFv4DRGR92DyA9GFsIqG5h7yEaAG1P7HjzC/PDMI+JOtLbFZE0RJ2Ac
m5hH4Q8KhgUHtk1JK4PDaJDvjK5lAK7kkHQ+xJ7q4e65oMvL8zjPEHPAhtAyNaZE
NGOa84r0TbD9hf4oUSUiNoQGSv2TlMv6DLHZvj7MhmlkceTzvJhae5a6go0/J9X7
b5syh/N9Q+97a3Th36t4ssRMlY3/dji+0EoWgUSBeSB3In8WZQkGVw5/zmyjhDTd
QD13Yv/lUK+jV9RGKVG4ygz1zPvMH5OWO/5ynY2R90/NYrQ7n6XKHAWbvC3aMpOb
XjTcMNUr8tgd5bcrmOKl9bfeymOz2kQXMFubNrOuCzohwjwCBpAT4CRPQKfLYQWK
P+L9TMlYtHJBwm0iIO4hG7C0TQqabprYReRzl8l1EUXt4PwMpuJLe/nmRefGqq6g
iaPexgSdHwpGB6rP7GzZp3ZpoyOMGrsF+itTFzaeFndd+9F+Ihgu2dN0CRaan4e7
/dJH5ntDhgG/um1WOISIETfOzKniD7Qiu++buwY7vJSite9WEr3He3biW6thtA0E
XK5+BHp53weNKig3n94I/hD15EdzojQMnK6Y53FlP+Bp/bc8Oh2DXnO1Fv87XiCX
uUNC8vRk0CqEcU12gSUEaMatl0zvyQdnT4cEc2v4O6GnR1h275SVe1Eo28X1Mt4u
2OBHYVVVIykEfZ0Pdyr1ea2HF0DA0sq4CzJgDQPyOd9F0MFqBOOPjdxfJ4V9ObKj
xXncURS+skE5TRr//DqH9MNws8qZNz0XJEoIR48SE3R66hk8U07HcIuMWvFkzTt+
4OKeosXbv2cGETRmj82hQUeNRBZ1YiHAUlZuBxo0W5Ad6UbJ2qxuPbgvFVqa134N
C3dOKDh2QdKQWm/O+piq3f9JFWX7uPZKZBKvyb06xrK4CjjrBbqyxc+kmLLshT9E
fBSWc5zI4BAHuQ4f//98RhH+dfq3U7MwuA+RKKMmq+k8oNQJoa/lS4xvIzeWPzWA
wQNZz444AyJWrk50QiGpDpHhE+neiYpFOzHYpogMoe7QArPfKwrOFYTwHbE0QMVg
WqpoUX4eW7wLE7+1XCg6rIyRyQdAV+4YpTZXpXXESm8kbno8lsWQVRB+BlJUYE0U
01FPB4x280rHJeExd9ecdobMcs/vEcGtIraoZbKxayoCO52Wu9h7oDlXjfB6EkYO
FhclkHJ0peRGDZhuDyV3oNIVOx8DHF5bUjAPhrs+yDch6uR1ZskPGMK4M6GvcfXN
bLIxwZKfHdwBY/VCjAHjf1b6UlRzd19FYqDsyyo9HPthb0bxKPU463LsThWbrJgD
lw6b8Fp1frJk08dUwdJQP8ce6up29TBmcFyKV6n2R2PPcrHcncvYuHYAoFbcMwlI
UNAMRBljSKlILE/9pEu48/00WtP0iZuDSnXyg1InUblCwrEdYqPLBdtxycnZuE0N
Mrz/dAqqEKh+srTUgLJqMK7Zl715pG5imb8j7pROys1qon5IUbXl+3lpKknNUzaD
cOFkUNWhREZf88RzYwZwQY3/+dJE2S477Ly7rmg8TS2u1CO3cZa6Qxj+ZRqFviaY
GQpOdu61wn0frUbk0onvyFvqkbJjAbmLynCGuhWLyxaxAgtfYtrQaI3ABK0NoRye
imtyoEAmIDMqg9BgMqQzGBdEBHmbT0kMjYS/UbvT6dmVLD9mDj0Gdzksz3htG+iJ
QpamxkxemgFyrO1d47+TqUHCYKfLvGYnSYe2CVcib/aorX6F2JohHiOG+EUBGFms
/aXw15hbylD+LmR95MVVydDoBOT9hJPqjLPOOe1a2//IBl/+gbbKBXWFONVSLmhr
SFXH3661vjpVMVnzeXk8dX1hX/SVTwisVcKsDp7SfK5Lh+rqDFg9L+dFkzrk1q22
iQmTJ0So2fUzdR3GmMIBJSmtoXMwk/KVngBIAa7+ZYsdeaP7fK4L/iflDtjv3vZE
YAukYxvtr0Divs2e+v/lz4noR2H+SsVxlbpPvShCU2sj8rJUEwS8ej+zE3QfQY2H
yr+wXvyOcjK5hKxv93GHohrtYrg6JKeP9lETywroBcts9yuys2PXp6r27yud/yqM
/u4TjhSp+0x1uUfcBBWYa0Ujecv/avdQgRM+4Tl0dcaLaR0CdzGA4p0+OsYm0eA5
CnOVh8f+A1ZiFwdvaWJkG1KNc2uU2hU4Qs+W9wZqSqixdJGhb+gtJX7Oh19vCWGU
jrY36mXJDCEaFgqy8FqVIH2bYRgUWYmFuDh6Z5qxcYexNSbkwEIl2hbDDeUsU23I
Z7vrPp4rgwyCgI/gsMrICrBSijhPywJLVLbWnZoBQl+xy+tZl0hiAGGwe+qKokoG
jw8/oqTzrBdb/as2DNzvX2AOSxPrbgGWPX3E0DpRf+3+UZ8beXjupB/pboeMm39i
8gnWT2khuuzApa6+4OuHZrIHSjWCshz/f72FIXOXkxcYEEqYoirv2FdBARkUace9
3eWJeLluMbi+SX4RYELFu11ZgZoYWza4eNRP6/udRztKs7wWB+PimK5BAikOJMEl
Z5Ij0x6Psy4SCMvxrBjZJn6OMEeHm9Yg3rCXudNfqb4P6q9yIQFiuIisuyJgcLH8
j0i8X+zkOHqQKJrt9EVrveAzUJoD769gI4JOoztLjQsd5fEGQ14CKVpW+wlGCWdG
RCMYnfiGZjl61XeCG2k7jSC7tkuqHWRpuqkAQbJonERnnFmcn1BMMgV0lgvSG67R
Dlbg/E6kR8PDwbvBHOVGDaP0Wtqorse8lW93xsGYn3fSWD0PWYxZFVCksJlErJoB
cupY3ynBdqphOskpMUaa3T2AX8fEtaKRwBo2xsKBeI97rESRhIRHra+7+Diqhf+3
76DsnkYN136HvFwNaNotfoa5FO3OvGnUah6Nsq3GutlN5f20uf+r28L5B9gioDfR
C9LDYc/nX7AUMTWqm4fU/zYUjwY+SjHYbdb9hiiDgM0w4uCKhlcRMd9i/YG4eRzQ
N0uyM+fbp7YPDYYXW8ENGneFmdAh8iYnRJ5LaAb0N0gYIdg2rDxOTTVAH9js4dz2
TxEoIhKVBqQlAv+YbSWorw4x/qaycQVrrU5bisi6HfWlXjB93jXyaJ+EiDLVn8Mb
LKt5Ly8LWLuV/n1MlrGdAgR7yIqGN+sHHrW1gGvai/sqyUhPA8yWd3miZxT/4SGF
9ua1dexy/d4XHC33YiI7vgbSCkzXMVjDzWsNS9Mwc0sysUAfQfJk6X5OSfzwyK/E
mjAYpIhFwFGiSPfjwVQBr/+mkeHHi7kJJdM23EqQis3G0IP6w9+KPC+Fx5MvrzC6
AZrDuWeckbSiZhN8YsI+bHS/F+XiNHNt3ltLhIC1GvGzgeKVsST8XD9ksOeSLWkm
cBsHqEfOUumEOnGBLrIePa9dFmjFjH/zRb76CMhvjI+SD2D73VT3yeSlFcZO8k5D
QwG+OKgdPuXmwoSYBLsQQxUm4aur9nr9GNe9rOrHhtV6yq5tnsS+jWzsk5B7s1Hh
EN8pu5hiiu9LbqkmzHVTDAr8DErMige9/FtJDe4VQemen3vscYrGlrQq3lFuSAEh
Ku2QeWLWFdGcBIQ27WjHDsctvX3UjgZ6tlUjUcWWXMfg6AC0Ti4TX8WytqhRQk0D
O1jDeLEwCPCXtt/5T+9OXoAQbdyBjosfHdn0oZub7Fd1cIh59NLSR5MgYnfd5iiD
FRl3ETehHEdGuTh/buHUyalrGzneoInb75g2F4H0RNxaK7pD6tzeX7ki9IwdPguR
GXwfA3i7V12x7Ypkxz88XaDl9gWltiTp8tfFCDooo+1q8jMUs+9Sl42sgnoNqEm0
Q/pYsVnvgd967j7kH2dhgKsIhFGoJLcjS7gGPMC/XPdSi/p71MWvokjF4DnF26xf
bfsOQNVr4zTFDbKaecLy6NzWUF5C25BGIkIhq3FQC1uGInMV24ngsql4dNdbCIkz
072TjGgnrPAWCKYNqBIo7iq8Th+CRXmJwYYsORb7u6gnv8eLgyXPSOgeIRxEBO8v
aW1778qUv3aZBCuDAaHlJbr+No8sW2FTFnUJyVu/sFlBFty/+q/xhxLNIzrkin2w
6MWY/7VDMvKzI+1mVP/lu7ZEbB5coD6Wy44UC/3oj5zbhZvnFqjyLe1BC3+y6nky
uoSQxJKB0R6Rd6mFp78XIrtrgtmO9+KapaxbxrLt23DEQxew/U9QArxQbqJ63Tsh
+zujwso/VzHf/tHyAeHy+WiFiTcQsOjfdPoZAcSnp8NkxAaM0UlZMld9BY/N4Oj9
h67yTSW6rfb0kk2UmRGZvlloBjXyiA2/oiS6ujVe4H1jobi3uD+bFxYzCSwiIw+s
cchbCUVCZK3P0gwgFd1xvpDWWh6NwenarLF9h7hFRNTwiyhnZZDD/Od2OgAdjV0m
bAmOIq19Iirm7g4vkAS2wtKBt++3BqweTPeOfFWi9ZbS8crtJ3wRe5VCQ8wtWtZL
H3MKMcPDYZBmO78cH8NEnZtm53h2kHDGdr6FYrFvVJ938ltKOGioSnn/6VRPcOdm
OBddQa7Rp3ZvEA3PH8PoNspwrTvApu/qlLT9DDWkhVyBjR9qhthBYQsEb55Vf+e5
FvDN8KFV+v57Y62Bv1u1GsTK0Bm1Yg+k/XFL/RtpGyZU8mS+EvvTxu5BzhRMagir
8Krg4rTyHfBes+xIwyw4k3OJFRxTvpnff2r+Cp49VsYk5g0B3qpDtfZ2CWA0S0lD
DrNyfvhDhOeO23IPnCmpis3imvPCTgs29srH/ukGg9dF+gfll5GJOww7ukfBdn+x
eFccVQaRt3KcPxjOT5GzrvmeahylLtnIWok15jJRv4O1QwlYIyo73Sd3lo5vl4kz
ZwdBTMdP7uvmapK5doI1hD5oUBpDTUFUYCVw9Yy0u7s54t+1xbhra42rVMWjaUGU
y/yCO0NnZWogZ1kIwQVJnXECdGvaYFPgS6KWjxFlKoyzfJIyGm1CyCBApg0RqJnx
6l8pc7x9hthGFbYHLr7vrhC7nb33hNlfbCrt8HEHces09R5ZAL4qQgRVxT91ZZaf
+Zgsi+sKRj7Hh8x3Sro8K74ZFzucuJV6r0sQp5yZZUFjWnkqu955LM8ep782+f3/
LsZCk/uoAY+66cjlZkTaShAPv2OKfVBXPG8sKeWHgt0wST3kyyRfJ/Bz3Y8qBW59
6ofYJLc7cfxXqIWSubvdA0Ms0lsMp2Q/ZJQV0yMJl3pA/YIMoqv6hLny+xN7jjiZ
N5tTjEbffRFIUK4Mo7oR5QPPQ0QnT/qGGdqbBQsWnIXcsFaxPOiQIF5qeiaTkpsE
hs+/3F83aki5DusFOyoyIFvkE1daCZcMyJGKLzLpJ4t9489hGnYQ9XtqETyzUsUU
qdStMg5Cadybrd50eov5tbna6HbWQ45nwSmFeCH6qbnFo/qA5aSimLFVKNL2CtAC
C2aPy040jCukwnAvisCpVeTBq3AtznXunMnKdJM/nC5WmCde3m8zIJUrP7jsvMi0
QjngsUdYddJCMlcsf+WMWMxGFrZ2iCemakHJW778uRgk08l6NqxZLHAbDDOjsRTb
s7km1NOtLXonDky4mYlut2I3E4UErLLkzkbt9FG8wTJ/Byu/1aOi+K+9TBzK3I0L
ljhB5M62S0pDUC4VEzdx9Ss6ffmSNuHiVwD7ngmL2tDr2TvjGm3szw7q/SKdJWYq
ziG7GiMdNE2vX7z41Ga9vOqLA7bwycilNf40VY0B5TwkF6DjrASfNDIKBvcE4N0L
4UKskyDcSoK0vE6+fzOf5cyMsHZmR0k5vTFNhkDj1Yf0EGflmPlpzEOP4mkraA2P
x1P4VF5KPBWNi4yTFuiBbwKt/x7IkkC7O1ytkQm2+7ffvw+79vuzr+OF9LYhPi3o
hFjvVsPu6GBgEEiYKlhfYksEqL06SSY0guzIBfWihh4xqejzT4/fEbc91kRa6uUb
eWXtPCnsS3oUrwuNPlM6KtIY+Ac/9a71Nk1aknMQ0CECRj2qGSHza5xHdlxNkqTE
p8aqCYstqHUfzsF5kLMl4MnrrdzsFmJtMrVpwfmGQfp5zHZwfpXEzMxxbdFsw1NR
dVjcU8N+ugj/yf4d4cmcwGIbM2SknsGIRzyROz9rv5J6PBDT6f3YBzzxPLhcaTN2
ko5/IXl3y/LNQw0Wd/ygFVS/m7BlA77+Tl1FD10kHliyYsG/NyOjIchvSbkyR2Wx
OTgAOEWmx4U/nF/jAsg+jdONYR+DIqcIPkugCjvaljt2Cy+avrdebWxiI6nb1XbJ
hBdObjVJrE4BNWtOVSaNerEkv2Wxo9dPp0k4DEViOLW7ZDV5YsZi0zMq//IeLIqC
+HerASnTgNZ8bVo22kBO9A1Vv70+4ijWQrveKzh793t9NOsMV4eTADJwjCp9l9RT
wNe2YjpRMpPWoVurdiKl+2chJEVkE0UD0gkghX/qHBqjQUn0jqwkfDFBA9PwY8jg
9pJGpKgbqqNpavql7KcfWgE3lbFcOyDZ3LresfOAST6QvPy+dRu8bdxrhseaxv1X
cF2W4trMJLHDFpvH9QCUhuF1ldftTWK5JtAedz54MxB3l7leLy4Qj/b3lZM5pRdD
itz9lR5ghWh5vvdBBdQvkqZ6WCh0vTbFoh60EFQf0IvsW+GJq4wNyHNJhR9qehvG
Gj4R+F3TgW4RiZWFonIc99fJokXwqErkhYAk9NJl8ZOXHrPVnueHEUW+upjrZ6/k
56Z8JeQ2h+x/3wimoqvtYP1WTn3clPDUf/8fCRBiC4R8/WynuLXVarEgbmk3qzEH
InJ5Sm7ha05XS0sc5rYNSfit9b8JEtF2ldJv/9AX625frmzNknrPFGfcvlGYhG/3
HFcM0s5Nt0E4pBKjSfV53KxaIDZQQVKM9wHMCJ/RrQZNx80WEmWBkC7JWSmYQxGJ
NvgV4kcXGtvahPIvk3Lkz20k5BUiVK5bdyMHTmTY5YGiZH0eU8/fazRgxszUoWoA
2Bp3HCjABG41A6dYrpyozme68pxREwNGIK44Alrm9gFXC1hkbNb6dWptACVmRBmc
dyCz54Cmk3R996TnMC/JpZL4C9HTkPKU1W2kHB1mOPvxHwmYIq78EfdzRsyfGA0u
TBzNPASEhDIhjxsJE9zVs6a8NQTiNlvzAi74ckuDYJ2ZrOaGsgP3NCDBfLpkPFtD
sNmyawkFLg6edFyE61qZkMc9LWqZHgOyXpxzgS2WqoQVo8oy6e7iQIJDQhifjy9G
kRFCkWVlM22UoXirg+ja0bXrtGQPDRu4WplU9qUBo3cd6f7GcBTNtGEp4vkKiel9
DEjtlh+DBeBamDc6icSYf23JnbqWx2rIN0QrdAB8PKwgCeaQlIOGbjtoW09/o5eC
W1G1iCheov4AS/WFr/T2pOfoNtLftBfzJLVFCIHOXJZ0iPGPUgc7m16Co0I2ZEqd
7MXJR3ruHJhH87CeGBIe88A0mNX34LyJ+cQkuQXyLGahGDWGZyDip1FdiD7OwBgu
bC7eP5K0EsT2TVsy7roEIWip+zV2HuqTjfb1sS5EZGmIANwYm17jGJg1Ya3Ju1+X
CpR7dd4YOkwUjN0L1jAABzaIntCwkjwMLxSm323EwNlVu00nLFOWfs6+Qg2wbD0h
g1d9sqQ2z0EjK1GYU/boFr7WYzYWSV3tMAKFDbrq95DMGMBgHuaoKnxlJi8FKxsQ
QveEopG/HJIaxIGnRgpOnwWZsQ0doDryBmvbmEMu9ygZuSlNPpmJ+jCxWb/XUNjg
PQCiPC+3u1P9o7W9zhieNlJxh1GO2lPGo7qSOMhuqbnI2JmcUquMRT5MkoQwwOev
c+KysMiKN2I1VV/Rvw/2Rnq15a0ochRBX3n4H5+vljeWWIitRemCKEynryP/Rcsp
VocDHBYuaERc/qeRVRnwOSE6BBtZ/rheo3Bhjj7/rQSejR3ouSsEnWwCPxAvfpM2
7zVuqiAcktbi84gjguJmxR1y8MKJIfvKaS8IEDCun/acNDEd3k87M4PIO99R/XY0
H/3L97ROt/EJNaPsWLk9148IIMmdKeSqhp4swaf9eAbQTmkWQqqptbk0cjRw3YFs
I0+wgi1mbpsN5o4qxddFlPvyaYqsnA0RLpO4L/amwPGDKl6wdugE+R77Yzrn9xlg
Lf0dIvaM5iVqLbObatuvEB8ZJ860A+BMMZQYUt5bnEkkoZ2YhILgMibk5/gSDxc6
Xaqoy/XMj3YE/+K7d3/aa+AJ9k6CCTGUuMJlqDz8tF70LMby+E3JgyQCM94ZyDPE
3FVN5RejEwuYIz9sDBVklKo8E+NFZC/r5+2L6mRIusscra7ixGTngz1PYb0GLa4X
VeqH3pqHaC4d7yusTN9XyJgOKxQphqgaMIKfyIgd56Up0NQkgW/nFx6WzWyH49Rf
r7XB53wvtY3egHV8pQvPytuG8QcfudQgfQUqElq1JX3SczIJJZxgBC+4Jw5UC25m
maT7tyx7fIhTyKp81ncrN+Y7joMKnxJ0rPnILCNJiCGOHzu1d+C9Obb83W3g6Lya
TO0R2kJv/uypvCRP2pgMYhmoDHP/W82KPHCSNpcelpZJNO2BGH/jOz/1RN63G17D
FBoIoi/xbhEkc7LqeO9BePq4VLvB5CIJ2osm1qP1X6cOt4rORKL26QWBlJhsTf7N
hlH+5ecWA4qju8q3iOJKV4pmpmxwq2aGeWp9F6UmqYfrMNmht2IEYFhi6Gfr1h6E
xN+ry90hvtLt8xEF7XNZcTj7ZeX6bJVoJsb1NnMK51HgL1D75CHc+QvSPXCW46qT
y8ZXTCcYBx7/iHnY14FFF8JdUD7eeBmkYjJ+ifqJsqRGesOPF9uPAqgILl9yJoyt
kFqD0xJcZgVmwdUNMRuEE1YM7M9Xc5Ukge/Bkiu677qChFS9iYM+L5TEXli8PaxT
unPLT3ldgRIYDpHUPgrDd2iBaHChy0BZLEkCp8aaFq4XI4Zc+Jewxf6ZPp5+xlPx
ZkZB3sxOJQOi+0CMfYZlhPN0vTLA3sROEi0WiS3ckjpJjSqYILdK0LJNIIGOAElx
Bk/UnBtIaVQIf25kdf4xF8fmAB2KjGhAwRW1/QhFplKK9qiNWaF/vnw7yI4ob8hN
e9uj8kFZFnRhUpUiIsjTStwxGARsBE4reBVARDLPHZWfrLybNga+FZcqiSjt1pQg
KMgMCKVVTNnsLtcEPRmmsJdGKpwkuZ/IMNhBnVnq3PZZF9rJwRL8Wly/h+85aZjW
wspgpAFH6UjdJuIslH/zTTPBAobDdG+aSuBSWkczEekbQWQpsT+38TyUxJzp/IC6
So0WZPzlsovf8dfyuC5nZsvKStzLNdJTgmtngollXQEoV2EtJaA0fEFyqXqom2VV
s3Dt1HxWJVEc/UrRjdXqWfy5d2J0OBGsoKoxqUSWH2NxMGWRuA7wMjmr430sCEQa
QiYWRF1qvJ6dLXFIzh3nrxhhN3XResSZmQzFPbO9hA9Cj3MWIEmH2ZPxMrfMZDVZ
xvzllHOk4hq1OwoYJb1ie+nlF67k2mOPL2R+q1rF4gjoIGhBXkskEGBe3/SWnnLX
QjfJX+ytf/kqPP+TR716lEctdqvv2p3G7pBj6W8VL4O37ZfTpyA2IYe8rN/xD0wN
B6jXKVGAGddRxLkJxSwomqTHBk4/GpH/5BStqqe2cvXCyTguU4Rye0MnDLkc7Fgq
FCgieLtJFPLCa9bJHzEKHeL0YghFobFBi0vKHBMR0f9MDMAmpAAF4k5t7aKwJLK3
PUrm/bEDuvWtWeURDYdujjNE7xjtz0bWk75yizC4P/vdJYWFF8O1XheEJQ/XGJtD
396DZAwIt07XkrjgKf5zOJsNpr4aOAsX71YML6NRptFgjUAy58TixC0xfNrPXrxO
AnCjwUny/tkTQiVZcmwRhcggsDosTkMhVrsia0x4UJpZg8ppT4ufA8e50yiEM7aW
2LwMC8cISB7fs94/Q9mKBaZ53m29QaZ2glgQEgbmBWeaHIK9eSY3r1G+nvI+DiR5
EcFjvHg3WFTAvqocOe3STxVqqdmCejArDS+xKG7RpjgbbW5/mDymYCWxIHerLCuo
ysZvdjI9qn6XKqK4IWoP/KbNnkyxkslhNgNi9DbFam25DAT5Uv3Ygf/HDdq/7wMg
G/J5Q1oX8hBj29lwDTUc/Zoqkftuj3xNx4TGAJdmrKgNXHpI/OCKgsSO7SGmLuLC
eOdq20DCTUp+Bg2VM6Q+o/MV/tjOUok7/qyeqJDba3O439gQt4xONhBuKPkgub+d
CvLrxInY+Wnhv8x4sJJGNBxRp198XspTeHtFXL7ElCEiHDVdbFwoqIpDvDHA5nnB
sZUSm3QTDhXQWw2vNZFPSxe2JbRvw+zDEDHjd5fTT2Ari0h+7zzPtp/NacWd54of
SjFCkVVFgP2Ycxu209UeRgHhRvGqs4GQOFDchNpspnNutNuaO8ZuBzzaOUGvtkvY
+XbLv1Piv/VrR4mkwiAxhCJdVY6xC/dbrgv2/Fkr+lPOIlgH3A2hh08uQ3QHp21C
h6a0XIDTUYYi3ON7CvO7gd3n16SuiCDdkFkaKE5wrkUFeMYHEbqt9IIQJ9HcoCwy
1JNcXUVZjIe7odAn5BxmO2+F00QbYopkOznFutLKlzlyDDgDchiMAjObfoxigaKr
jgmFYcLrMPDEaNzs7ZN9VFeqdi6QaCK8uZKumDi/mig+OTncImwmfOwhz2w9OqQg
oIvmwfMmWuo3asRJOVTtoJTXtCwofPmBckyTHivysQrd1Ul+PlRXWeCKLqKNQ4Ds
l2HblkRtHJvUXe379HEW4QlECIxffdG22inkx/lT+4af8B5hlP8bh+Nu0j0iY+Xw
GoWBR0Cum/aQS8JaCrXC9WPS5zbPctgZ6sbwK4gCplcu03jXV6WQSukOsbpADJcJ
mqZX6SI5xQz82qV0OFJFyS3Rf6gbFZ/Jmvq+BL5AqK65vPBOT0HNZP/7uQO3GMvZ
btmpiHTTDgpo7AH3VdLMUo4H5wWM1X85Y7Lx0h0T/bauaAafqCqz9/s0PCJ8D9wW
SRx4jCAnN03aV+C8itNUxFoPQRnX4WIoiUzye6tjUNCFXv0Bu92L8LRKmwvpojEG
6xpSJWjgiOPGyRCvLeO0ifNQF5fESKSpFwtW7P2AY47x38O29YQVkqXul5y7bD/J
gOM9C1DD6HqaT34bKgUPkIverGaBrUX/v+XjQbAi6voHyxjxju91CWq0w2vtPOGV
tatnYPKa7V8g2ONCr0jYbHbldaTfxvrAPW3be8+9g1RWdt5UjQiN7zbjjLkjFL1p
FaXHZrvAJEZON8zkvNYIId4jCxFi9xLjhRze5iKyz92raFKYOQASrLds6b/cRmfA
q/FtaYfUfJcVNmyiGCE15dugzmmo4Rw5tJrstPuJiY5wUx6BETBGuH8B4URXEw2k
W4IhtBb6JG4vJcwXtf/AGbQRh16WlzEafNdci4ldsKLp2qSwum89RkHb/lX1B127
THIfsElxNsiJmaoMQhrZfbl1Z9QOszSEdxumBqcQrL9o1ek/8uXqDz4VMOhcUSaF
N0VfApR4g9zMS16i3CmLUVKpNQNtNLix2lz9hWK2SJXc+SZzwPiXqNGtDsxK7LmL
ikqcYAdD/46rbxfHtWDQy9VOvLyRoxsRpyBe++rgCK/Qklqu/M4C6i1TL+FnCoe/
ynEsUPXAF1D1CqYlEO783B3cfJICyGFpsZM2nq5DlfHDZsGazx7M+dE6ThQjbkAI
keFYVQzeA3Ok3cxVKkhBjjmH+OPpbETZYqG+XMqFvvRpNQMyhsbB1cx5xKyi5wwx
l3xFjA9nv6RN++vANnnlNBbz9ZyIK5ffq6INT3OQ4OWf13X0GIbQjvNQeG8K7Ckn
82ulloNyvuZhgmav4r8irOq65UKvHOw3A2pG8f82vvX3W+aGxIscgdSSQiM5VC4d
S3q39jrMGdQJPZwPb7yHfJv12Ph6U7xQb3jI2YbnDTGigCes5oidV+dEdgCq+jvW
F83uNsW3YRUtIQAhrEtuplSPcoLMzzr4XSPYhrLw6pqLg8sm/UyitmU0WLkEchDE
FZZGTpzQvwsmWxgcb440P4/jvalukTB3bYNFnIljGDYNqraI4ShHJHVXK7GWnOzH
EpAk7TisS2ozb1A2x7A3cIxbZrYCqOwjWCBwNDsrZGJqBYyzzJuUQAEqvqn0AT50
5AU7tYEQ54ExFPjezz6G7BStMX/JcDOm+XSJf7NhfU5xoNjwuzJiUiaDXg4OZgdB
Lgpowo15dzCUgkSkivVCY1dUvl65RpkaTopDYywZk78sEGInR216xMLMPWhuDcWL
ywrXYF9aKy59/lJDYcZFF29X4AODa9+P+xu5ut/6pLPUIGRIcdYl4ytoSW9CKXDp
jV+Y/j44y1zsUvY5h90kahWtMHy8WTUWRbf/tH4UVvmLpzs0vFXAxHdRcO9Txkna
A+E7YEQ0qBQoLZazwyymcVfQGMf2gKJWay2K9RjSQWghDf5xgad7h+8AfIJTUqBD
aRTch0Zd3wEjP6ZxlhoT8P00VNwq7WVWLU7jvORo19OOdm8HDduIvy7Naz/X4vL8
gUvZswylos9SXAXIEB+q272YM+Qbgs/J/IqWTlG8gw87gTaxn5raUqllBzxnrP/P
tiMG6lnCsC2kGTrNPIaBB8rrum1QhX1whB/HGUfZId2tK4DgiEJA27aMBMBmloFX
tKA8Qa2KGgILeIuq4HwWG9aWc+0IMflQOa2uUCsTQWonWCiUYdfhToCpL3/Hm1JR
Gj/NRpePQ6XuRpLjabHH7Lu3UH8NSAtnTTJq2Rs2kmz84PFmaXH5wBnVo3sEsFYC
tW1tGb1Tdvk2/PCezPtyzrseGusQaPF4iCYtRiyzK5YW/cdTFGx56/QOb3qJBjsI
8qgo7kP2MTtOOr0km8w67eAl0NtasSvQIr/LPunWn72KuF/exYASldXSKem5F3y9
xPfEdyNK/lFvvzw788u+RaWgxoa5GEu/iHm+RylIwEo2zfj87HR1h23Mxse/MS1o
Te8y2bpWqZs+AKbGq7O35W8eVkAoDqSYWaTSv+Og3zxZHIdvd0rm/0ujDEUl2c72
LSQeer8Ld94xhOTZLPeDBSmKIOPXSiiAqBsld2laycDW6iiQn9sdKezPzy/OIm68
3RveJsanJsobIL4el5cbBd2dvrDdcUNezJA61DdrXv6v7zLtCfzHOpDJmpr+jgIo
oyM5NRNFZGNSoFvsJlaVE3dwY7jVgO3un3MOUkds/VwmYgmQdmIThPxR/ItIsCkw
XsETZAGDETZ223auPs6jb7uxPojm082tE3IXufXmwcqxZtEKyQnDvDu8q0yXRqHM
TwR/gMuHfch9Wdt7Z2+Le3fIdQf3zsiYndwwhv9KecufKVOXjK/+quGh4RSrZcMK
1j83Hqn3aAPwL+Gx2Olri5qSumvVD0F99appltdqgOABOR/g9RTvUJ1xJhDH/ZdM
BJDx++Ekhn1vcoWLHso2yEPS1/764wl/j+TcRwBFvP5GdbzcDvW7TVcUP3U6VXip
EuRuRnJCrYXABCV4VHM0q4TYGO4LlI9AvU4/HqoqFv2MlEgEqH7gWd1iXheVs5VE
sKdwFF2ySeMA6ZdlUJFOi5XstiIrz6MbAsiekf9yqedZXgb4lvRr840+3HVMqrjN
9YnOAApdDjSGY8jAHu73pLmA7Oaue0bNq5l0iLvYd16NNvhjfajHGjKr0zlEfZ2c
UR39Qcn1USoBcQyjDUUUy/wOr5TBkJptnuKEJQOzwgg13XeSSZG07RUS8EAzJ5S+
5JODSgOaxdVnMQh0apbQbJRJCGW3TAALa8NUuYPyXd7596gNSEmRBbPPbBpX1nC+
kaq+CfxF/Q96FrqOerth5043gZY9OSFvD3a+7ghhFqbMq0VLsJVnY6AzxHSpHo/3
r8wGuMvHj299BwFmEO9KulrNkyGyv/t/UdnUJU1ilcMUpjItqn1tqJpwtYluz9MR
oam6UfgR2cqjc3Un2TU4Tw/PjBKl/aw3aRDOvvFvFY6rQiOqWqjmMh9sHhAy50xa
s91kGOIXFctSdLp7unAR+jTdPaSQu/rpyT0e6tDsW8CkqW2CNvHhKi++oPZZG6Vm
xImYr5g0NIPfQTWkpnHbCFjhZqeF9iKeHPMqeAI8Cmq5MOOF+v73VDXD/MhQlM3J
Eq9qR3BAlq5iM41cuJnjLqqz88b10RkYN7/k1oNoGOGlQbcn/I9fO6GiACec2rM4
M/PCWycpq4KC22A/xiJPpxczlOoimFetXuFK0acM2WtiSHvhw0LGsIRYB90oyMrt
/q6ZEdvQwrOhgDqyETXGwMya5h2Tvo3bkhzRglAw/zeoVJTdmpcJfdhzEdn9VHjJ
FjYVpjllxbplkFWe+Hc3Ojt+1rvarTIi9GDvXwl10/IzjpCZkoS802OANe1a7bj4
MIZGmNVSK6UcUkXYjdUts9UddRVZPoL+rrKQxEH9PnqTInVTghFKO+Yo2bVsB5lw
jWqtITC9EHABYvpLgBiJTDI6GA/rE2yujOwsXazNnciDTU+57+pQFELHYrHb5uNe
zfmaooe2V6bRFHQj8CZG9W8C6St/rdFb3KoUeJfGLV7Rv25XId8HY5oxTJCXz0he
wJS5ryKjpDboDJ+gvIWaCDpdGgqFpUiVyO+Ml0U7bkx7o0uEKjNHo4exx3dCi4zE
Nn6gPCe0HUGyEORzb68f+2HzZzyxcQ+Ur9dhR8b4lZrVTi8WMUPFKEo9eNjwT77C
XLcGkjen+mGvnTtXYFgJJEvdC6sj50THdxW5umd4fDrt0TcZsMziCNPg7LTFoBQv
rTKYcD1QLoIOOBH6ewQcGfGGdXY+jcaHiTSzAER/KzclB2WOJxcNUCwhZJG5dIBL
jQ657C6dcycA4he0eyaUlo2Jb7t1A14YF3vU0EPWkjI2UzJ3fi6dHHVhHKNnkr31
74esQnnadiRGd8CX6aJ8hX2zKCT/OXuFDfFv4Q2v7ukM9QnUxKgj8ajAqOLNJeLi
hkGxWv+Qc3hiP0c5l0JpvC2ey/rA3zdHrXq6R4963gTXpVDwzopz5Lw937IbfLit
wQQ2Ot8aNJbQ5rBspnHEW7SFCLxk6l8/jA29acrEou22S1zfw0mVVycygky7RklM
JgjL6fzFmyJYtjxbRWYZQ/m7JHAL2QVL2R1fgftZisvhYW/henupfSPMAJhkzR8R
F5VwRoanHXq0hfCxx9bxogI5JAIkBb6KLrgSIwOVC7YHi0D5F2w3w2Nrz/bGc4o7
Aj5NpEZI2257UJH9nKaOz6oPoTd/9yPQwP/O3NDKUZ436qREYkJOK+0GjqzVCjEh
/vHksgM8/cqiSIcfKHWNFsc1gkjtyyP92hicMTZ+dcuDfNzUwTvlwsbXxbCiY4BT
H9ZCFWz5yoljBuyaBpsHZw1sx5433niVCbJDdZhj1Rmz13VP8OJ7nfE/Ml3xKdX8
vzd/q5zRpVylJ6Ni6CRxuhNv664sGpNmtws/iKpriUTuW8MFfCNPSHm0GE0DVfFw
zDq2g54rIuXZb0glty4NgG1tfqTRJ9jt5ZTcWPLIEWE/afUNXRyfMJflyBFV9LNf
32bFC1QmwhTTsOmA/DhwEI4NnKUN0GtLgAmuZNwaP1m4ESyfp2ZxEnYm5fBSQA+F
vhRp1zAF5nnSaWIvAZtPaG88Ns7ccpu2QBy3nUV8Dt67cWc/UgReBsf7fXGJHExK
uqU6DcS0UwHVC2Ml+ueyGrphoYC/wf7eRKu2pbKEfTR2SEJhd8kMsjzmjMq2G18T
Yf6EZEEWP4wUoT8xXQiMcieuRfy7ll/XMhUV7A1W1f9xS9Y4YiEgskJ0hFmiba3U
EoLgHRt8R6WW6u3Ss5tgb0mRpTH463MfLn//h5DD0B+hYH57vWmm1JBxoGrhZVsx
v+TsXH0BwvasCtZAJWQ1CfBxrLS1/PFt1QCcRu8IrrREbmgh1kdR5IROGk20GSyS
bE+Ujhu7THwgEyXkmc95UP3zHmZFajD5OOzELX1pq7sA8IJQnwU+/hzR5sq1d4aC
WiiS8I9CcGvQO3Lq3b2e9/hUu97anTQzh0f6t2x+YDPTziOhKkxSfmBGMwkEdNhl
BaAbm5RZG4TMmKQdTwtVem1AF1zO/yk05jQdc56hMnHqmy9ioGYZEE1Mwc7RFMV/
79PRLCFXcS+qFrxUWZ8Mk4hXOwk5/H7fS50csAn9Eebsfq3bXukoK1Ur2sxFC/5C
NYjqD1XExIBNk6RI/uhOD/ytTEU/Dmu5I/9RdSg5SsBPQIa/yG+cMpeBKj0imHqz
yJW1+dyVuT0ACwW0LrmI93LRMgH7xmBL8wQppwQjsEM4TU6Gdv6Yz2SgqaQoWzrB
bLaa4R9zcQeWc2MPj20Axlkl/HhiDauH3xHOMEQMI3N0z3oxWIjzfjFLKoTlY3ec
2Nr+Uz9jSQ9jiCqOOy4XFxV1X6kOtvk/q3rUto80RX1x0y1AGgK96dB5ZYTUadox
QCKjDo+VZKLYhzJJwFnYviSdmxjML/kYlI0xo/AIZs/SYVgf+yeyjuxDNQZQIFMm
hKGTyvX4hasODqEFKcGmB7LVelkeBnxlp7gSdupqMJYPh6xRqarU/Ozn5AjCoE7N
Ml3zCsQ2Ydv1/rOhfZ3PbiErahbXOLcqGV4Xv2QmQEdEiayb2eRmJNMfgzXqbFYo
VhkRNVuHJJuvyPb6DC0Jm/iDCwaJQ6EAo22kdzcSJdRVmCu22BdLc2I7CbnxI1lg
eMqIPIvuv/E8K9JQD9UPFoTn1B6XOfWwgWldFkmffDv1G0HETi2sYooVPlHVXyt7
SMMvjTWfK/lXhmjh0HyHlu8BIOPVWKvvQasSSDkb3xqiOvxfnQR+PEssJFHn/cR0
yECTpzs1ftanBvHgFxdYJvVz05KbvXm6/G/xEn58mRb7UEp6+pk11Oz8SsNq/wYI
KnLQ7UEAul3CvP2bJZ6PQ/SYQxPca9VIoSphRCA49TFDV6dlQXQWvXAdcHCRXpql
UE2DJ3q7YtDtR6+Pe6PLBJQDCnn7ds+8SWAV9SzptWG2FIe4pFzLWbEmCuvpqOtL
xjHFvAye6HGpGtaffA8J9Fdoc41uUw7FRBghfzTqRSieDz2wg8yuAqns0x/x+9LI
bOMU3aEVBWIuNcIUiGwqVqustx/7pd1HiB1tW4ylEQZnNkKYZjWUn4rOchnNUy3A
R4NfAD388u8hEUPQ6UppXidVdf5Sg65zImPxx55ZEkUJqvmWRiVy4FyJ1rQP48Uo
qEKMvQHFN+0mrJdfwM2iiZPHpiEB6UKQpiFjqMx6bjkTy1OeXk89Jbu3A1uwx8zm
cJ2JRpPl5jy5JURRSKMw9ednDj9837X9g9r4h5E8AUcG2rzSs5+ahm8fAsFQaSY2
m+F6+ELPF3B/WksMbPzosvwkPxHwBfYu85wszo0863t8OGM2GqCfvi2Ra5geatar
idgZLZQsLfKhHwSOAXBtYJhUMTlIBXDDIn+QHt4s+MvcNEUs5H9JB/nmjWwAkgEr
MNrQRG/XEuNzDVwUTuyiAs98Gt74atzjE4WLr2hF1jK/F+VRTmHR1JhrPgxbq0P7
yAoTVbuvbmgwmDr+/l/vp7iIDpCgVAcuZ6Kdw/u7qLLAX0ZT5bXV1PQ7OFnKBdxX
QmAUEz0yQmMedpOOEPucK9xVXFOXUwtFlJTwXi7EzB9xuhPafmRAsJtaoXCMp9Q9
ZBrRaR8XcPufTDL1y527jffzRdM48sdWI+rwHsCad32WIbcyjI6moIFpAQdVkirN
GPPnGY3NLCXcbsOPYOakYIgCsgWTWlmeknlVv5MbbskPJ2brQQ+He9mkpq1nvyRZ
8Z9QE3wdtjHwS9Gz/ChzTHZ/g1TgSKQQbtWrsGJETW14gLUe7OA5Oth9eiK48cg2
rJa/Zfml4upxT4nIVfvbIidAGmXRYTkLBCmqhdKwOUB4hZP6FtWr7KNZfs9X3S+h
oU3iJoqQAUDHSwwIyHuNy2Od/0dGYvssr/5dIa7vkwQXhsc9RxLQbecD7U5ty/Pn
UNL++JoZRfv8g0UuV2PgYcIUIW3AmPec16RRNGl1yJAdiVXDOD3igSyNDP5K9ULJ
+/HrTRFUn51ouAOkvkP3qoCazu92EIrvlilLJi1vW3hFSRYkCyZDHKTbzTyET8kK
WuV+8DFLFrp9JtiUv2rH8gwPI5lQlSQK/0m8O1sK6pWxgNWn6gt4XJg6r0zTfVl9
380uYg0GPyGY28RS1kTI8hgd640PRS/cMj4wb74g9lAswcHJNiAsaFYI3MSX3dyc
+2WDYGb2YITEIzYeRNPSgEf/gMVWdlBe6duaxOWmac6nAzYuGLrWZjhU5i6+oj0g
JQdeXyBSvsz3eJ+mAPwuD4sv22n1dU0x+gTYSfhe0slaMOFojd3wh46mtEVDBXcW
dpmoxOWovJIe6Cir6NvNc0/+uijZiTFrlkUMd0sLu9EeVakEyP0YzNkeWmcyFzXs
hIANIdKWSm/AN/phk6skPdWWxoEQZrATE98NmKVKQTWU/eh41nR+AKtjSHoB8F5s
pCAoCUum10HHjiUvhoyxHJhVnmvffgkcoisR9kbb1VBtB6xxUTjoHOpqRijp3baP
AhhvrZ5k36uJFwJ+pM8koLWLe114EmPaj47gPPP9vqfdJrISphSgbmOad3HCD+cE
rce5PecjIY65LShZP+C0ewV04Aq9n4ys9pxiv3t6IUBrP254z9y6MyyY2c+3R/3e
EtfNm4+OEZMVP0HM1Yu2pcabkt+OMS8EX7BFeCovjZad0dS2uUH92crtvqp9R7fK
+XTI4prmg9+VsY4oRUL/842LsI1Aqu7ULY0jdwUeCEzAw3sac097zrawyVB7h6iq
9E0IC6OH0xD1M1FtrvSW61qpr/kwq25h0yasyB6LDFxI0kCqAVbCoHJPQRhDC111
qVHCG9AHR/im4ZEmIRqxR7yYvzx8ntmUGc4tgJEWmjetGQG193TffOw7iKLclyb7
hcFwIDER4goPPkPveQaiv7HsbEFi/Y3Pwu2zStvb19AZPe1W7htjR1HHBoj1HNBc
DJP50fn+LSv6HX9jvGAtTcIZyv+Py77V861jn4Htcpt1dAu+5cUYdlY3xLGl+iVx
whKgi4M2boYgtQl151wCaM/KNZC2+bjAf+Orgla6dzdb0j+V8piOaPSsilORFARJ
FGDBX3g/h4PHKkB6zavTt8SjfpYDTJ/qMF1eM1iYVvwK6LcYMdI1hgwMWgQQL1wy
njYUg2ODj/Mp8w95JVpoMPmSlS+H452ki3/46JlbUIPxDeMT5OnnhBttgXyK1P4w
b4yyLEK/NgbcXc1VlL8ZXH0akCS3A4geYS5sr6HY1npvoYVMt5nN5zebDFoALD+9
D0TFbDdXcc9R/J8L3rgGCIJjLMd8AsSdIv5SJrNQa/HE8HWRIaEZmjs0JKCZv/sM
mZRHzQxemccf3lWvdDNSNdGJg3r4m6i1QcnqZpc5kkjj2YgsYBf/yZLi2CQjgadM
R99hYWjKq20O7xo1DV4eMxgmwmOVUtLBGWN8Vdu7+/ao+3WfOmaopmkTxm61szZL
xnC9v0v56zXLkSRUr+jLUQnCdi2q4E+CBJUjnMqWyLprMYGSCjNdjljXgRJZlqcQ
lgk4VomxGgq8WJXGROFyLXMPXnndUz0pxsNaFLUe3kWkJB//yjYMSfuOSoUj4tvP
BdO06JcBULzYbjn743BOGwsPuzkSb4g+E3kN/CharHsAfdKZW2SPgxpG1o9oBu0K
761t1ijLwO+z1nK7gj7Jzw+LTSNxlw0YlIL8ZStGgmaNxxYPTVzmlfi1TP/Ik3ab
LVGDB/Fa/gMJdbkb2rvxbxHJZHMSEMKl7an/MpaDFphVYlaWVa2VEfrOhm18RczU
iK0QtEUiWo6fdEh1JsRASC87GvjjK+dX3gXAd5KElonXehXR18e98owL3BISs933
Vxt6rSaHItQE8z9By0xEo0A8b7r5l4oxH1uu4I62LeAvsTaV66pAZ/XU8jnLDPfK
bYfkrTfiR2k9hHo2nB+k1sCd8kLcwgfaXCe8sEa5l1WyKX2XP3565IWNwHjALftB
yYGBb6MYkq71S7x4o7a/sQBdP+Ksb8EyuR/RIYgHBZ8Qn4d43/GcNd96EqLMHp5c
8yfzoKCpFGO5vQzvWc/ohUYiyMx2pHls/mbCGzUFprIgQSo8TpBso/ZMKB1MwsIj
9a48kwdkffzpIwACzvTKQmftJOy/s4bhZF8Gol16hV4fcwyzcqv6J/bXPGnkWTr6
qhVK2ujFsAOKv2WPxlN0K56zj5oC/pJgUAg/lefOQIAVcbvReHOl+HII2jo0Xmhm
wAWhjM68K0lcQE8+ZBrAYJaGJkLETh0LCCAT3QuEjulR7XM2ibwfDfxt+b9hSPb4
ryQIg8JGHZG094mCkruvo+Go6acCoSAcIhieVW+2/Ry9GkNJZmMQcEpkN7IG02a4
rPUWIP8nrAeoeW4w7tCRimGly4dpdw6NNgAyF+XGSYB4lvo77skpOPH/aVlGqQcn
b5EXvm7TLWv+ZFWZbQomNLAJLhcsYpNdrP5M+R+iAwEXSpklEU3Lyxrn/PirUiNh
kOQPa1Xlc9HnJ9i9jBYYdyuabWbagtIwAb7A8M1q/L4xXz1QwafSN7YVUe4lhGl3
vrr7CyeIkoyd1x5KUzP9fPzFYBo1zThkPIaFYZw8IQSlNZVl+aVsEEYT4fLo0iPL
uAn0OQu//V1a7SaENnAZOSpoyjVO1gAuoC+S111UsqNyJRRf2Ppp/b2I9hmkEZHJ
9ueA3cC+Y/9m2BPBvsvd1OSJadX+ydBguCENUzBA0wV7OQjITsV8sXcAWwf3FtoB
1hhGeldSamENpmzpl9lIsD9Kl3Yo48T//uxNhObldViNRZ4DA1ekaXq6NSDVhZ9U
KwV3SRWaAlmDVN9tfia3pzLc6XOl4xsTsCfjw0s3QXOcHnHRRB0oSQAJls+SLu/x
45dUbwioD7zUAJgt7dfoM/oxKzee6zXTCtLe2m3bTIOI4yKbuM3AagZRQk+23T4L
LfbdkbknTHF9yqh2+4gRH3Ew7pLz51PM80AdNOlXKlORs4KO2qOExipzbRRh8q0s
ptPFAeajUEor7oBQDjusrchd8JvuoW+EW9HXTsnK0ZVWdCATfvVHzQSKOIo8hiWN
JHlN2iWoR6GFYTND1FhW9BKPRR/pzh2hA2R91YsiYl9RxAZZIirk8RpgaOA92u/R
tCzhauvqtOwmmbqdwZUEMUuOlblMldSeChhl1QEywrs/gm3ROqNt2Rfkk5ocXQZA
SlwoFgxzefctm2bLsP5+cOxXs5b68lhCrueGj36YLuqHlRtg5FbR0oLMRrwCeeF9
QZuj9kjMUqGzkO+qjoENZbd44XUqYcaDSEcb0atFAs17WsgpdwlhN0pC+QTr9h4a
xLFPebEl8uNVhSq/TiKARzPYXVKAhbraEGc/3Gf0zNUn7jAeMjxpDlWiN/TWMLkp
EqRGGY4QSOLEYZQr7EviGxyipMhnc6veksJI+PpK1GxIVwkFi3uxt5UxJ+yi3Sj7
qvYeTCogrqqpFtWnHitjPR6iF83HggfCDrCK8EtV6h97XkFa+whbFBvI0lvw1IUt
OLYHcsE8UCLxkDbPkxMHzrdwaUyimzfW41CSnzhMDPwwCCSo30NnKhd1Ro7ZRzRx
PIGacuzon2TvifJ8xA7X7MleTvDHXP/Nihp53b811oSa/+6IPCx6kk5HF8w3zmvA
Rxyl66uFBSyk0x9IGx2EqNp7rVZU884hGDQCiJN6VLfRRHG/5XbAYhdxrLSuu4oP
n5dMWmv1vIhHoq1dFAf33xVeo1wUrVBm1aiYzX+EY9jk3Yy0sMNVjvFKfAPt3veD
tQokKx/Y+aMb/SD/oyT6Xs8o78xgHACibkQUPViVAumR6trpPSxdjx6cUfKxDEin
U1mAIu7Aq5naW8zLb9RnGjjO0MwP/tXiuuidPVt2KzMmnAY3f9rg5kxa6fkoBPAR
fXxuPtNLQ3yg6v4EXvsTI5aP+lKxpeVaGfYXw0cwlQVIv94TVxsO/xCTd+U3d+Ah
SE1je5jS8gA1qK6zLyb0FgQNIv1xhNWp2SAap0AkaSOloEoMDBtIVa2Vo7xe+5Ga
dlW8w11HucdW1XdAP3epIHqH5W9yKPK9qIpGNxftVXXFP+eb+hu+p6cGo0NO7TA5
dMldsr+SoCcAdU/aoy4rpIeNhqx01im5bW28QPtHfFsCVMu8yMBiTneL3IEtncGL
vGjVTjOzdTyVRoA7fh8JMheyonccm/1cTQyamTcWn5YKDFEwYCHeSChM1lw4KXeJ
okuFPiwW4ok5gn9aZai4mIlyz3CQdy7J7hrtxYjvsHew1TSGnZQPWW3p63ZjQm88
QzyjYVah3JqOOAHR7wwzBV1aoVEJZWlO/o4FCzyPFzKlI24xHhD2zfIviW3fO66p
R0xzFe7aSELE0rgGSe2ibdilD0HqUwlY9D8uCxZytz5R3EzSqjnmXLvDBADxPtqE
KIGDaht/sIoqRm6NLQKMAQkST4Eq5qLPeGu4qiguBabRwdm4t1UL+TXiFRZ6uVxS
8fT3Tt558gWd0cMWIaXwiLc7fCUDfeM9mkw7YN+f5gFxBUeEq+DdTFahf5Nl3Lna
oYJ+qC2f66cc0QkQfA30s5Hz/mrIxoTVT8156clogunOp2GrSm+sxJpK9VyEgRzu
LYFKohj7tb9/VWhEF3+g1VTDDIL2FKM20wT9juSxsszndG/mL3RqfvctZwtK6K0Y
aa/57I9QBUWnZYFwkFeGHRDEdiukL7jN9tmUgNxjcn4hyEpSBxDKyZ0ko0JWfnbs
ELpvFs2eCJq7wz4EQzs4SacSHrdmFqhPqVJlMAMdGKNJfdUdpFZbXnAeou8z28bP
tVnKosbgh6+XNJ2a+yENHnaeKFkFSjcUky+1vgSrC/LyANupm58gsDFXJW39a0lF
aH2pFxB/OA7PK0C0R8GmWGQQrQODXtpmpyf1cgvOkyzeFV8CaXyUCkRbbkCMNox0
eIZbvK7FOhJxvNorFKQ4zD3vlT6TQHjakilX6bk4ewQX0SrgwtKpGN0z+qZYuy7E
w7MPfdss18bObJBGzQjeUzskKgshhs40r+PFoQ4+p3+y/+Q/3nR3VrdtZ0M2Xgky
54+jWtL9ET8tqsyCkzV9PK5syy4NdtfmrWjnhp9rc9B0Y76fTKhYZjmtnYk619gX
wWutGSkBP67t6utPQyTaAiWFPIsU7Ct5BM2wi1ZLCv51lxuIz41c54K0cujjVUgU
j5O1DrA54oOVenbvi1DxOtOj0YPBpoMULT3RThu082f17+BHfX5JludwI3tHiM97
NmKMpQhTstSvoYA7zCXkogF72dHvUqpvJO/afA5oRWqw3oZY9Ng0XobnGcTn9Lf9
+z6kYBnQESNGS1CHxoLTZS1HiTjvb5GlO6ahnNXdAx9Gp7YXh7oRjdHHRdziq6gV
qNEITMtIXxiiuA1oQALZI0sJV0HQzDhY9Ew9BQdfoHHWMNRdlxARUbiEHJJJcLIh
f7K0oBeCqVSgikdm3ITJCcpRNp0difdeLe+3du6rd9MM5Pdg8YV94TbkAhJFQijb
pQat6jQmOI9h7lEN+E/ZIH7qDSGZhJWH6XLBa7NJoppIvhMdXAKA5ZgJNaEvbzb8
mBs6eDXD5G4oY/3y5JkNQO77B7w3oltqTzfq1zW/ZnSudodrgUkweGH216JUa1Rx
VF6vEohDst5T40CSEpb91vBc56Blui6pxJi0ccittfrY77QBvgJ23JdIBL35I4C1
RWLGM/vv2knFCR9XKY6Y6A6YCilSWRes8u+TqCH8GZFJymyaY66mqLtfKXxZCsOV
1Yod1iuQajCD8jj8TQxR5QqC/IuxuHcFvaB/kd/ak+A7zPt85lSBZfQTRjHtx+Af
oYcGAPbLVhZMJqevfR9J8ZouLtY+szTYRnrH/ijGlb0iO7KZhCD8sd5MtT6+sikC
Oes8iiIBoSCvMJEGb7ogLZF3m33jfTtEk9+JilaTYj+Tqk39z+P2T1jFIGm/s8A8
etXvxex3mMyK0RnBgfJCg+fHdUgYcOC5aPL1uGHqB2hZb+J/iU7bhrw8BHhb+JGE
tB+m1VWdmqOvqo9YJiwvo5pS6EnSCruNDIIteMVsJExsuw5+BJT7EPDHjS41sfmC
CROs4ZVQFRR8osoEQyMpnyJk7PKk/Ip6TGujyNYwwu/R/Vh+o2wMBVfnMgrn+t94
/xB2qPI5suMKnCEwnqYHTY2hhPE4VZG1vQqMtcl/H4P8fSU/WiW16EB3JlEb6vf7
VMPq05rhFHCt66Ayy8emEmLdMHUAFh3xbibT4bX6ar+qkWbcjEb5PlVtd2tqv8pe
gkVJmCud4JcBwCmX4Fi7MElCQ/CH2abOZtrutOFKgdy7yc8eLTau6+EB3M3Ziwad
E1VVvZ8L6+hC7ghHL1kD0h9F6bWUqeZWo0dv+OKRiSMyT33rsq2nQUCz61TwbGiD
W3TLEEELcOXoGo+ap5T47phY9aaWeZWiIXaUnPeNoQ+QkQFl/DviG0hURjZlsjJv
/jIzGHm8gf6B9vWm8Nr8O3y8M+p8bbByI39oEXM/ZwHeVFI5k3Z9xamotQTWnz0M
rrwUzqk7/FCA3gVh85MdghSBff6XMZYKoBYMVf9pqQRndd0Lnu4hPg/83Jsp9SVu
p5+/r1uUfyHFzlkXHj9J2bt1WSVoMf4m99GFV8zFTProyJDd8nIARsdv5x3Mpmq3
nYXKFqGpANJVc/NAdVirfsmLG00xLS0nij4ARpMeZkgcoLhLLhGNZLU2Q+lxkUQs
NXz7cbv2zEAiS+ctX5kODYDFSbSDOGusvZgBY/LQphaQO+4YfQ//aM3HP6UfrmzO
QfW4EEk2JUH5R2XlEsJIw8C9Pa3wxx/dwoZItr6d73ESG4Sqedh9irT4yDzlEI2K
g34iK6Y1G5DPS2qGSQ/OqRuMclMy50BgVqXs81lDrQR4LoRzePBQJLANevwivuTI
3+RF588PmS9/RZn9G4IYHaZat3qvEiqK5vKxN26ErwaCoETslZktFBCvxe8xfc1r
FqetjNGlci+9pI5+yokEZu93o7MuiXpdrv7NWNbbumz/Kli363OO3329ebFgkHoM
EPZPAYBuk29EIK/0Qc9nkmKf0N/yFr4+qxeq2Dwr5LYi6i3NB0fcViABni1UcGgy
vMk1jxI+bjBmQUuCrijLmZn2z/y5cxF/30Q9WkNw3uiYRcektEfa0z0UQKz4qHko
lphclG7gk+uKr4JpsUpCnOsTeFh4zmah2ZmHStSkSeM7zSOEI0yW2Z9L8V7vc988
ayNA4OMAZoKqc+iuytcJmE/ifGtis1V3s/8XUxcvKlH7+jZLzRQWJpxHeXLhpYk9
Ht7PbEDgQgaS6jNvTQnX/JQOuk8DjQoYfzar9vzGT4vt93iJ7+kDLrFXecBZKfzz
7/n+d6dCae5smQC7Re0irR1JM2/fwXV/6bmq6A9xI6ObDcV5lDgve77XO0pnwcx9
MsO/tJFb+IlXawz48wMtSh2+jgBLOB1MePL+aT5JKmYNqaSDy42052fzk/zkODbK
MZL0ozwhSpDSIlU1gPtEIbjGlP50KIefj6K5Zhf3c9hyBuA/E/+M/wuwJzpxTs/a
CwDF9lNSFMEtNJOs2EABhH/4rVcxC2SRkkGFKyWvi5WDjPdu8fLFauyjRamfeWQI
V4qxSNR0mIPyJMbG2r/uZZ1HTBlCf5H9BOFixAjVVPHNS2SyuBbgS+3HAl2E1Gor
yWwsCVdhjQq9PeTVTr96lWTnvyGrpW8Rps7B1pRD/o6RhwrN6cqFdIW21p4C4dVU
VFIi5FSXOo27hbVnmuD5s6aUQVUi2ED4oEf9GYQiHfyAH+YqTuX6IBTVG/JbsAPr
jCEJJBDZjP8ID75DGqtwh7zj9/pRxpj+7YknoC56DFZ6n4xj0biGOWTkvZ8oWJCM
SY4is7lXWb0/oySo0mnrprC0RTkUGxyneo3gfyW9FuVW2JqfL+fRvbAWgCqKugOa
vwFi6Cso8Q2gGxeHam1iISUEAoDycmOo7JZ9p2Qqk5UxxtGqeNf4NRH8DjT2yqHs
+bEtscF8CG+3kH4wQOy7xm0GNdpNXdEEE+s8rgGh5olpGdG6aSMpmlNkDIQwdWj0
aoS4KfP9mJwFSupafzzZ52jDXsxnAGiGRSpP3mxhmFgyrroAHQ0ITFfJtQ6WQBtN
B9L6P3Oh11q9IEtM6J1Ao7zT7EYuANM030EUEzHVhTuDDWZ8rTrpKZUGO7UVkl0c
G2i1NQsqqW3qLz5r3XCwEs6mChUsmDqgDTFkIufD4IlcoZGnJg0IGzNT5AGKQDlc
ugREcdAY8pTnqwd6t7K2+7sCCS1BlDyOwb6Hi8AsVmAT2XDm1hKJdgCigspeEY4j
gfkAGmNI8ARQmEsZdd55xaWV1lxl1DFDNMFThrsvyb5OQzkAQuVE2XpE0qqTUABq
B0v/x9/5hPbFwlwS5PUrHNje8KWDqrpnx186xG3lJSfaOsiaWHcXmZYEFJwcHMxR
ZRE1MhC7gwHRl5k6y5tzx8gRXEbc747L9/kodkBrCIbn3e7AFLDtWhdxbSeti5xc
nnhgKLtDRYDGFE8QvtkTsi6wTQeuLcmXBpteMvI7PM0GehoKrwcofDxE+Hf9KjfX
WnxvJigL6gHArxrXSDac54KFAB4FkhYwKhFUxCOcIg8Ol0SPocrAkjXIB7YMqLY0
Ugcqe5coBxMv3l4zM71Dus4D6NnMo5k4QGWECLyxZR+P1mlEnp8/L0k0ZZKBmATt
b6qc7kjlprb86Qhxs8rVRRDzNgTax4o32psU9jJaCcfq+LG7YHZJ3u56AH5OcPa2
sh8BKi/F3qJDsoLvmKyr3FvdHxGvtxXKeEtBP59ts84/MpVDbf4MY+NcftKflaZx
/1tnu0uN+hxogFpQa9LPu0va74zAa6OBtHzzwab8DxDperRKWyEyvzeMk4YEiAV5
SsJypZz7N839lnnQo1rKPD6oKwqyBADh060dpZHtt7FjHoXXbTqeqFqgnorVUbuW
YhEnnSRpUQBlVWPF5uqbmpEEQv0MGUdLyCLr5AZQ9KF4ll7r0cLIHo/askwB0xvt
LkEgd8aFgQXByka71HsHaEUy/g9j5dLGPeiKNOEvcVvw6oTwydqJtTqX52GiiF+u
pUMaD8vP7Zvw3WE3AHy1tU+Wu432+apRKfL1G2aGvTWRrjSmU2C7Nd++Lx+jQg7Z
Cojb1xYVATg4bSOYXQZqjq97Tz/Vh6hjQA8ckWXI87AiJZgKHwg84eeSkz5rm+UC
QhNDci+gEpwR/aiakV9cMo19ivgoFaxH/XG2ld4ms+DkQGY2bvtUl9bUjHvtY2Pn
CWWrVReMMYkwbFpfSYsf7nOVjrQGITIUyvBmRBElQIctKd6J+U9zV9Gf2L4NWvFo
8tB34CTYlNCtIBNS4lj2M4yGCb34dNb6B7OPI3kfDLzmjyBEm8/JZhVLFo9Dy628
wxMkbkGaVPJmt6KlG4n9Aj5DBWae3AvHtOedZfMW6+oZuiOVraWxao0Y4I/KSzmU
lT4n7O1xLuvbIqIbk/czxERdetG1LGnBKrhGY/ZBHQGwTbk7/bTYE5YeXSbV4AlW
Msvzet3GUqc2+6D8sC1/Hmc/avkbsMgRAeUtyagZNhsOwvMnQ+V5xMkZyWBkeI6D
UJy98HqSuO+umg3Wg0lWxOJFH+9LFcW45GUvt59LdwObJRrMAmb71uhDrqbVb1lT
8VOZCbkfXYMGB3uynMiMnWVHDHEfTSqhgCeIH36d4LL1szJONh+piV0VunjLT+P4
vJLYM95XXZZ5cZu00w97JDMN5IzNNJjX3uT/W8zm3v2oa/B9xGL8QwnuycCkGXp1
U2K1KcD1PXF0KwEVxSJgyMJIkowtytxRbvruij1tveF2YhLpZpnieglIwKhxATdK
wl3YdVCnnwagv/h03flcnaw9WOOuzF8z4i5atbXXrGK5kKQqo1IvSW6fDA97ocbq
ioNr6CJGQGCacRtOAXgscoGZmpJ24cMusxKTopeNIp6Bgsmm8PvaXLdLgiQTuFNK
VpvFGxxspS1IjpkFTQLHWrQSLyUKcPHzpw/3OKB+nI/KXzPvjoXlwzc9ZMAEJe0t
b3i7DbIQL3n5dFTPImp1PB0wm4vPnecYyJxD5o27kNzs7YTdhjD+eP+rP2cWI1Ur
3ty3RHVDP/VSwh3wwS3whJm+UNdhRDJgybLFbm2AKrtOTvPXaTyLzJo/jOQ9IQE5
j/DOdkiqE+tJ8lU+3cRSA1lf66LDNL4vRUUyLDHrTJO9THEyBNJE7DkUDhVefr0m
tQekcEM5iapinvZb0lZeBPwQ31t5C4vgR1wPS5LbeEK2d5+Po99IqqAeYGj1upqQ
AzmAINh/sjhxsHIJfS/zFa8Zrf3QvJW9hJErh9up9nPrL9p24FkWpavVxNKBWK8J
/ttYgnBzV9a4SZfmtJfXX8tshxU79ccJUTY954qGiPqwNQzT7NAfmILk/L4nSD1P
bwSj2NxiVWST6pLcJ+cG26TMsDKdGeeoflj59gFF6sTMd2r/WjoLCEpUfkoDK1uw
li/N83Vlo6bA8x5wHOtilr1WQu0Fx5HaMI/owLY2nN+XapsQUK/0fJ8bUVNNkcnu
s8D5L/PZjMjx8kh1LrEHQoP2oNuuKCvkotd0JbOl9hhY2z3W6JbIORMQWNCOigU1
SfMhEgnqY21JIIqxoakGlmgCclOJZy6sIYyQS9r3aqH+tH7qYbsA/R2S5KPpjoip
Yuxn5fKTlz1i9/vNKPqaGeLPaEQfgsw97TEgg1p4KBuqd/sPfQF6oRsvxXg77Wrj
K5g+D0D9dltHb7epHMsHKhl2Yc/pS08hXXtxWIZm/ckSHfOMr3/KgEFcu3Hhqyrr
mBI6FC0MEmZpXFR4J3bdsH27KEfuhiFgPkZFJQFrM/z3QzT7F1OMu1rjE+Ou70vB
SlIPq2lq0gh3hwMYNM4hBwndaqJs5YQZE35fuBJM0WyBgn4/coHbMX/tmXNsgmnr
RprFzZxwVLpRKJU+FuD7KshkwzzklFpHdTKxORkC5cmHaqvwJyISY9MJvazndmJk
WbQbSR2t5C29R4G5m4r+8WUTrc53x3KrRY2Op+t4z4TFdl/ExLJAagLH5nwfkjGv
hMT4n1YdlURWJRVkIav75bKyKaOylwrKbSqfr36OHr7TZgdS+2qvlksOyAZAYsv+
slZVlFI6JALMElDtaePJWeDfYftrOY52l4KFCP2Fb0JKku7O/g21Lz3Jjsb78Y2N
ggJPw6JhSXg4ypPuVbTmcs1mlate0x/Ve02bwKuudfylT+9EYMvdpINrDU1O20DJ
rfXuF5g8M5kqigcN3TMZ1S5alh3Yk98lKDWJsXgAPC+xooRuMFXZCI9KiA4FwR6K
svvpf9MZz5+pvRI3FU9bQXw9IM2YAk7FD1gzmvYgNtrWGwROBuvPKNxJvYGtzQ7C
7OaiM2f+cqxdxzfNemRhBMbNubPU2mHe0ggajjVa4N93VnrxO7dDhRKMYLF/luhj
kyC9YDH8EPEZx3O9abaVKX02RYHLq1H7FUkeBKXbxLdUqN+Rp/hZBL+BrrLXUoQh
Vwt18mvkYjJYbzOJUlWR4KKb0KOcvDGvqX52s4nwIGdf4knr/LoPRlE+ts3S4LLZ
dkAmu/Tfysm+jEeS0TWpLIffOEpgZUtYyqvyCjM4ebw8nOrK7i2NyefREU1EToDm
npPFMfgAmbJcYE/uRAF1tV27b7CjkHHfwCfKZX2tZKn4BUChM+Fkh8zPksTK+ujU
hWJ3T1CtHxp81kbf0Fy5LGtVeDPuFrHHv/duFIK0aDQFF7biLWvxIQPOmex6t7EF
SHU2ohq4aZC17Un6ebxYLdO8z1Rwu0ZFokyj+5oCqHrnuhN62atLiAKgxKVpzKrX
O7t0SjPuj+n1UOkLPqF7QDCUMMQzMOT8huIdv+LbJbiZxzIysIT+y4NAJZX38s7D
kno6FdbTphM0AjOnAiQ2g3hBB+h7gdkdtvwWSEUzbUJXC9heEwDQSfEp2Z7NN2ij
z/bUuGSnm7IpbtILkPk1Zb1ckMQDiKkFmq5/efzwufU8cohRWpuyf1Hx7CEh/rhT
9uXpQUjsiqn61Wih468qUqPYJQ5tC3Ccn5QyXWKsf42sdEoegsJDzTE6CWFuszES
dq1sbvNul+0r0cy0Ow+66ZxptOgBeD88KKhL76qkIXKfPzhqytp+hUKffnhB1iWI
o6/u97Na7tdiBM4qpQoS1r12gcGq/neqg6cURxiA7DPOdShlKIECX307IWOYCZCp
sG3s+B/lDFMfj10p6IxFrnGcD+LyZPDpXSnvlR8tHKVD/uL/QwBn/GvVepHen4NS
jygLYbM0Qp6dybE0MkJpzt/GqTUIKHDEqzncvJ14wDkeiKTl4oBuZ5u9uoD5kR3K
CclqS4LjnIC14qWJcbovcSSXX3CkbEZ1Kc7jhcKY/c1qC17um2A6NLIykkvqNt/c
z8lFSCZi2L+ucrzOqzp/dITZ3DvSwKrg36FJ5MUFJn+iJIfMEamUm10u60VfxrXa
ccHfR6ydth/NS1/3zEG4X6Z9+2/oPQJSSVX+z0y/rrSkU2Nj/y8ANt3TC94bBzgf
W+ldOGaNachMwcC7b4VOqxD0pFm/zmjDHsKL5SIjxrP58y2KbZ8LrAPvVRTExFIF
ZcqCCam1We72eDaIXt2q2PWvwlIcR+qFi+VTT6ztpw96qPlpZOpUMi0XW1ZgI7CS
WF5QtBLjGQcnCgosUW+Ux0EqoICiYjlvN4pEARkFQ790q7oyZ22weNBYxCAw2dFG
6V0PpcQG1Ej2IxYblNC3Rh8QdH3cVJaafZYGergLTFV0Yr1eWFMNqbtuWERfnEaX
KUnuQr1Cp9UTAFSDj3jZ3jImTT78JCWS/eHQkhaWRCvpE65+zOGi9U82oZNeuFIM
oNU8zUYjr+vqEA+BdOxdv4ZwZ9dN6jm5ZTsfis+P1i3Iy3m9NkNuAqUrJPFmtywy
YwRFwPrAQGfAyTL5g1d0WGeCW2b8097S1fVWf47hP4EG5UlSdn7oZg4VRrRQee8f
+plof4GuNJ2ejhleEYU+uUCvcFaF+WVrxP9BA/T61j6UovQ0uOJv4uyoexUjSQkJ
ecXXlWdOhDUO/8QmfF/cOHlbEeQrZOdMy9IFSn1B5MKpxZyILdjlBgCfERSsQMNq
wUrb56yJswtxqSDwMx2pG2xgw2BLEv3Vts4D6tuUTT5gIfSkR+ziuw1h33isEz/7
K+Sd9hUfiNdE+ju8vX93XbC69R+XrE0e2Enmqx1ZS57qTPXfGkoG1kKg5I9NR5xz
a1DlqBpTzH+n9EgPcCz6dMtfTQfflj0gzFE6jxsmwVp3uhqmDDblkdOlomJVGpOv
c2lRsjIUGwkjSmcIP/lrQ1EvyGWWRZ9E5qQAlEuQoQjArfpY5j/U2HxH8vl2rHm1
vb/JSFfCZHLD6NSelj+fOeoppL1g/XubovZSfazfeacmMH/CPAXUM25BzUDbR159
soV/yxLCtcuFMQwkFcHJxF6WsB27vhesr1AcWzC4y6G2edNQxtOtVwbUe1LQ9yKW
JR8yKVzPp+Q6gXlpR4l14RpKpv6gYiq5VW2uHoOBPVjraEQloo4bOVL4JZXKLd3U
VYsOdm9QmRqlu+d7kWnKMGZrvpV//J1P7ZFQPg+dY11Usi0SIuN+Dtp8i/4LC34u
kyiN3iBVpwyAwEnYkRr3XSYe43PScFhTqw/xtuuJ7taB81OFeazOXoUL88QP8ien
YJhkifaQTqNnzlD5u3LSuddM9nyO+sxFlPpzb1jnMtmecsvafNlk4cyk60ngHz+Y
x1sYOoG0AGnf0VkSSgQjQkdKRbrx0iCuE2L8B3U8yzvNHEWMSjfMYxikDFcqMSiW
c1KFuo+KaiEU+j0q1L9fIwj+2Jcvh6O9Njdt/Q777uAets/XdYFhUev/ecR1lG59
1ZN47xcSuOBYgt1QpNZfyz1lzVasibWb0wm3Q0g9XR1w2tFYFiG811T3c1WfS0TI
IATbi+OxBB1F12DGLthlLXtIyiRD+CRG/ZYNNSi8zS+Gb39mfemWmmrijtgPyznI
/irGH85HvRbORtHihH8GqqsHEiNSzevB7w1tIC1hNIfZT9JGm01Z3wWsMXcxZIHO
QbvbQNMxsJvopc+uO7H5ZT/GUr/kOnZidSUEYL8RBsOxrjwTzqKyrtf+zDtnbwwz
Yr0i5aDu9cOm4Pqh7rIi2/EFAkS1sXIDqNwCMmRgVCDvzsJtcRpd1NrbhMtFilC9
R/9sy4AVwSiC6UiF74mDvYf4Jv7sCK/DRXH0n9HFe95HQr/yhssh6qQC25n2gXzz
lbMjyM3WoZ0uCYnFDstpBtpVH4PKyF7EBGgp0AK6UHRU9U5ivx0hte+/xkoQG+VT
z/Eii4GLxBeldJhu8uSAyTbDHHRWKQmA9hJ5Ct38DPV+ATlySI5wZXTw73R6PWhT
CyEccXEJhDXbgKeYkMfIVMgzvOItNLbkgP/S1AUjp9TyJakonFdF6mGiiLXKnAjS
Jw5tDJijNQJrgqzh1tTqfhWzqMmATub8XDSrrnc4R/+t/01BDDZs7Zh8uHTw2VoR
CFDXJW3H0hVSLW2Oti4mQnWNPnCY0wzwQGpWk1fgmbDh1TX/ts4JDldQCrLG6xub
8SqyDBbcmw802bb55AxLJ+omz90nNH2h7bsZZJkhOnaiw4lLq5wq83FJTb462s5o
qAk1XUBR7UvCDxKj/xAcB3izHq0xjYcuJ2qzIPkUP0XBSB8ESUpHa8/3ffwFPElY
15AAtj0Y/ZNDxm7CpA7QY2zvnQZ9kzHWs6DkUyPMqofT5oI20r3GvRGAIeIYXLJc
rh4/Uou29PDSrOkAgSdC8QiN78PTB8/K6e75jwcI1p8fwHMn2FwY9WLUk5ctObac
sf9ZSGzOTDgNQjZFhNgTT7huIdZx7lFHBHoWz/FGz3qJ7abJ2N2rWs5oJM78HcVe
qPf/z7TfsHY3ldT9/jjJWJuiXUAacpnZQsecVdZ6lzoaiFrIPC34zPj+Cw8HHD24
oxfjg72ucGebtyUjD7iTKgmeE2rs3Zrh9qNcC+XKSeGaPY7P2OzsUwAA+LboXZwr
gduTZWT12REFH8BO3nH+WJwFNje3y1IYE/o+9j4AJrAkw0+nb7F/NTV4rAuCjxNw
iau22vUGvQr+xK0wgJqJNyzGCGAtCDihpPZI2tdpRO/TVP5mqMwGYAO5sPT4fQy8
n1tqeQlUjNL0C4VLRYV8fAjVpQaJjWE3lCLpsUjlceuOGGjnaBkqj4eUJNQuYj0e
3RbfoU/Z42rQA4i3/Sc9iSWtUwAM98s78dOllXyfKVraE6UhH4PkCZ/yGX3T6zRi
2k6zmZY4KNWZCoTtAzPgGTdR0IsrOhB8oWAp610mDkdgpKSejZi0CMroMUas1Kqh
SZmid9iSnMMhX7h3Dzvw56XuJq1kJse7gxoF3UrS6I42RnLFm5wXCGr7waAf4vuX
diyU3VDFFFGhyWvI4rN5caKqF9v+Z8hCyhk+p7JPwDKisXNWUEN1dorB+Ua2nTHp
LPyWiavF6puS8WYvXPdiS+xWZaLSo+3Vya2eu7qjraVGq8rG4nDrATWbdJ+BxSFS
338qugVFetqGKXTBx5YuqPooNKqDKAUOyclcO8d8CZ4CW9udAPtKcjVRQHBoOmcB
PX44cD/HvT43Y7W/oNtHxMEqc9+j1EH6G3E2nPQaeTB8CTOA3dvgKrtULtU9WDI+
xcP4O39kU4t0Vleqzk1sm5rNBVQsaDX9FXFG5tK2gDlSmEC2ykOrvY/IpjU8ZVjH
Yszq7JHCvpW+SkxWbHFlWO7cHKNYnx5FpP0y4x5zi6f6ZuHHdYZUl8Tkj3P7aZr1
Xvt/mRgnVhEjfQmwQ7PHFdUUAxiILyITkien7/pETH36tkaI6EL9C6dpTr2mI6ng
UArNnE3R6fz/o5EUXn097nzzkVqgSKYqXzDSvtvOl3BxHSCVPwFxgmQlhb+lcwI7
Gi6zVDuBmzmRS1bX3rzZtRyRaNS9TY6U2CpjQq69zm7XCc9Dz+98zFWg0abef3HB
HNmlYJS492PpWVvcraulJmdoCtf2cWT0WlMgfZzynY3ziiA+Oa9TYwpMoM3T/1lh
3qewB9gmoHkd8H3I2C72RkLMZvlXt7z5HzSXR2lu4LZFYjC1HZEjoCTgv4vlCBQw
kNImQ4zkxbAhFWY0YXhqX08qX2lACh5cS0Nd8BNQRL06im3hTxrKwHN/5OGKzp3+
GZK8lcmwgVrDyzHg8AqAsJgYRQd0tiVRtgi6VZBBBwJwdVETR00pAsuHxPw5Qc2q
mgHjYs6rU4X7oLBMibNjZM/t+fem18xDCH3ygTAaxoYers2O1182u/Yf0bX3X9/s
RX8ufVPQnLnNbCmCZaVHEHHMD0RFIPRvqwcYvUp05prX9G5/p94WfaNsF24MrVo0
ZL1QvzkqlyP8G675TXI77DA8iifju/Ysnwb6gNTWvZygKnFHZdwoJEfLy89qP/UF
yZQT9EuEaS1H4OOES3cdIGDXLJ4cweHVyfH0r8+A2zKYE8gQASIrnaQwIHcsUttb
ronIfYcAN0BD7SBWEFUkXL0LD/trOiIVrdBnYU+KWrgA91YId5VR1lmzNM25j0S5
YjHmEUW4fBoFE+7I2WiwC++8w+Vvf+GBL5Gzo83cMFGQbZAEK/tRDbPU3gGKZ4vC
lCaAz9tzHGvA7etVqrEHrJjLNntRQ9dnwuOza1tubfLqd9pdMozRUwaGG0jjiOJa
k6KnHEt7pv5AU7XNrOriZBHFrFSxmn/XyW4QaktvHffBe9rxmhzrhBchXVH9nYfh
WbAS771CHFf1H2MRD9EegcJ1l35xnSdb2x0Muf3qgyCd/O05kXKET6wo/NCPZnjF
d3GG2xdOq8vXtdhQzBxWnVww6WZfhZ+XXjAXGwcON+2A8X06Iax4mGcQ5YfBRky0
x9BtnFqZSWRcmJ1U/lZ6GY3+D1HTIsxSz2qjs8sTV/RhmdoAZxjI+syS+h4+2JKP
xLVPZofss+uLUzh0EFdwJWWsgcIV4g9fOgePNbXwf0zkq3bxJEcW2Ng+ToujwZjC
Oe8SthBw58qI3DGPZR5CypfAgkIVKd/mOuTb8sXhgH2UoHSjFlopOwI2NQq2qEnP
61+x5RWJNTkQYegYNmonXqnyDg+PSxLPQ54jcQMudoGw8b+aFqNTrONLT4JYxtZe
e2Wy/jFZCsZJ327AyHEbvBiNOOm6WGvGQEAasgggElqkfHit2+CNXcONrDC9+l8h
U0bEW/e06eGa25QNp1nyepffJOvpLFARnqQeWXz395j1jvMNAdvn9JpeZSRyYvJE
rJbJrryTf1HIzPGumsFcsxrDc1rAEIwP8behL9UR+EvWpZy7TcU7ze0C9ug/R0aX
Rrgi0SWH+j3sTGPEaFayFFIVSsSW5Cm5Wr1HJrrsh+vKSDpeQu5gwnkc930wwhYQ
XbdQ7fiAUqjXsQOJT8/Lu4HS+pg7D/Q/hAMEsJlKe0viz+KYvkd7qrPV1JxVHWEX
L21h/DJOq+HTDOZU8phgp42GBj/SaomWhhVMW52pX527WvHWuT8VJuF87du0mqbx
5CLkTM6HzNZH5hqh4nDf5f98I7Tg8pw3P6NGowbpS7sEVrwehsIcwOh3tCftRGJv
hXuGjBTlFGvb1dPw5HdYb7gbR4CSGApRV8heLurVBdLm9FwNnseYSMtVoQQckuTz
JXuAIVbmcqkj67mhAVDdmFqxp8BCOb1t4UxBVe0wKl1STFAVZ+axkn0pAzWplQLu
/NizKzeq9vTkMQPmK96wH3bxWx7UG8tfjvWIYHw4szvFyL92bvbWmhxZoNMhH9JH
yQoNq6+J2N0GLrv2sscPMCAV1+HaaFnPmDX30Mh0Ed4vQEeMZe4pE7pKoSWLBfND
0OmbkGZ3KnjKciLv6Tlre1FRJ3JSI9I7MeT23YET5PPcmAjYGHWoYR9NVurrrFVR
eRTDL/vlcfImtxASlgJ+cmA4TbWIJuKWFhi6i0d/cYAF37LQ8KUl+FrzEU8PRr2R
krfEIoSiaZuKGCOmu/HnCA677hY0fI7TP5iUqZdVKpCcuH1EiunGwVbXeW2ZcxRi
5vfiFqaWB69cpit1wpRBv2D5m+oce8NryRQ30ME9kNHhUfCRPcUVlnoTL6M3bxxI
Snmm8fc9B/YgIZexq3CsiteUFL3nyKhwhxdJ8mylxtszvJiVf1tVxt9zkBnSVQJA
56Ohxtul7cZObMIqC/KXXzTR3HPKkgArMeFbQa+G7QfdyeP+gmEdog095SZRqG5n
1oYANr7GikrqCSOdyHEXoh3X8b29GtF8jqva03Ac2KqzTycsxLYLQygJkosawo/V
v4gD3Cc4W7tKU0oUB/rhJ1SCgW8Z4I0pQI7NHYDLNvtkdiplq5vmw+VHz/ygo8n1
WgJtsowxabpU3agRg6mBk1IP2eBHV4Qf9qruZN84Dlkib6PSBbGfSQvsDryaaTWq
L6qdBbcJbMBvf6wPHnqVQWwiBdyOMlAm9wu25tf9tjA6T8r1+0ZGMCCdDZBz21kP
uspI2bbNEfAHNhPWvgNOnfQdXx7KXmwCkSo7E21umIArCq1Zk5EWtVU+jfdJP9vK
6SChOpSXSvsiZdTDw2ZIt7qztQYh9vZJ1JM7+RgUUH6Wlz7JEv2ubX9TIcn1DYwC
OKw4FZEIQrRuP8KrEaYC1P7ZjS3zTeXhB/R/O3gtvIOsqBM004Rw4HJAlXRUuon5
VOVt2PdvG4zprYvK77ueO1Nz2RnfCU1pq5PLjf1xn1L3VrpdDWcaAjQihS7BaLLf
eiWmuSr7k+leuyXur3ll744yN9Pf17K9Oqnn5CjXu92fbI3e+2on40RCLUsn6aB2
hdZ5JDa1G3a2uVUUXUJhPQEczmvcU6sMXPQq/UEwWaKqbVQ1frK20nr/ge6QKLbu
8ohghQTEqDYFrHdl7tRa/jUhbP2KyGaTskwv51qEog75c2hSCF6pqfhIdy2KVzoH
1df1wIN2kGMGHvEtNYx85DLvFVHDYnYg2/NzH5y2oeAzEJykvNeeKfy+otKEvzaU
gdPyIhw+b8Ssz9qmr1xHRSWUapbYUv/EqTNMzw9WzqxOR9PGvOhcbCA0D8/CB58P
Dpgt3hGt/CRBXOE759ntDZn7/uMmq/bNFuscWkREJRrfbQufGr/WDtLazAclTc8g
UmzXgoHi9RUOIosobQ9wuLDguloskOb+/ZAP96xjp6B+NfbxwXZn3gAUR6L8DlZD
34TEaCXR9mZPmdWCcwikpfUXfM6n5ANxCdxRG6ujg5DZNHI/QCtt6CAc2y/b3a/S
ugV4KhxZHYGX9fjkrhReZgpe6MAqcabsaMePtCBh6/oHJYiC9ocItOdHc1WjlWbk
UW/xRAYJdHlJpaAif8KyH/H7yZqNKFJ1dQwu2Ib3fYcI/diXqX6Qum19F1k5j6XG
g90liQXdSyvDJZ2pjDegf4+GlLPtIpsiZL1gm59cSEnp1rFlHpTCKIR1ONXcs5+S
Moht0/o+y+YrRoLdUnRrLRqPxj+HSl9Ei3v9VRbxgIQ9LNFGlr4UsMZCHiSouUAE
uLxlh9+shMbYY96nCxKZkmFGzcQ57tznJceVv2wXU+bDcLsfL5XIikCVFBGAerkn
nqEiPXJjMPSXXWuG76gF6niaIvftaN5ZU6unQEu7B1L1+6u439wGCNo/E6dDOAfF
N9nf+1DYmzmvJvNIS9oM48jIJCfNUUxFF8pJbQ6b0D0Um8DamIU/zQ5X2R+sb8fS
4UHvEAgqP0iTb9BgT1CL0yW0XYy+UxJM5/98i40Px/qdiogzrKNo/qOYtkKbqgBm
i0Gz8XiJJyT312iS5GawSyQwqfnwqTA5HL4php66F0m6yM8SDJjT0VfdU/ahl/Nj
kXkES8MhohS3Ds5QDPUtPV+ybCMkSKvBnUUVijJhkB4l2Bhj01ym1Dctx52gjaNa
neejPIwubHZ3JTVDeRgekox2L+CuuKkyRTkq9SHrkFlZFTqqHV4J6HWZWdlc69SZ
w5hAF3LLPT1JUMAl9eTbTkshYYrovqRkFbLO41/QF3O5cA1k6KopdGSpNr6js6uS
NTHIdifgAFNfYtioWFdnDuz20v5YGZHXogi6tH7bmpare129yZUieaOYMAXxasv6
kq6c4qX1VbegnbNjmwcGRSdPwSHttYsd1MSwrTT0CLxFG38+XICveACbNOivZ8RR
BToMacFn1iDWRmosFvDf6xcT4mqsxccF6EZnrFt3Q8qTmJPJFaVnYgx685PWk2DA
kMT7VcRH+qtTYgIqS9qhNdFNvWRewvINiWoidoGrT2Ue2dg7NWUqBpshJNKa8spY
setFIC6jQaVgY3UjNhtS8I10W2jgE8q5csJEg6OahzE+fMA+fx86w7dZC9E0rwN5
HOmctHI+45pBZYb6DdYEy9NQOx+eRam43tY1qqifXI5cvRRzESq2/REAyCHi6VWD
h9071U87UnFuI8vI/co8jUkNGuE7lkTfSy8tOxizezLIQg24tM4LRBXreZwgA19T
GpEpn9pWsQtJgZ4VxtQzMlnU933CfmK9ZsqRIveP8CaFwdMJzvW8KLADG/kyGBjE
iUbzYW6+4D8PhBdBQrg3PRgBIOEu97PUhmmhQjhYodvU543qTmCD7l5pnVaxWBBU
9uClX4pVEiesBZfC7g0dLBM04C2dY/XLGIXA0+7sdj4ANk4X4huLitiSUGRDa9Mw
3trb+FpcqwgmCbXgA7jUJgIwGc44MG0HOnEC8g48QLDx1n3bS0yiwb1VKEwsW87k
qGoxgE35NYz6YcQYnQ/6JFxhxlDWq8qcdKAD0QjZdrInIzKB/L3B6tcM3PNyO/Cb
ZC76p6lhZsOtuNMAP5m4bXOiqms4e0kLIbNGULFMzXl4cDDyrRC0Eg7vnDtV558q
vHLnFnev0sgztDrCBfewc5Csge+JH4p1z7Jwyh1YOy/sEmTZTl0HP5v1MCQDe7qG
YET+9xHLOg0ZipEeI8FV0uIN+p52lmMpsg9n2bnkMnvw2zj7/pZTh/VnqdZyABgk
oYNEUNm45AYMGDKK2vH7bG9IkLy/lqwnYm2qm9LVWtEcL/oLJ9Rziib+976/CH1y
WH0eonPO4kfS9Im3BcLK4krAQqYORE7B9R2bswGhcBBfKHv041bQvHFq62Jhzfit
yZAvp2y3HMExBWq8loJH7rS52w4J9MKOc+jHGNkre7vIByfIZ/wZOs89db6OCQTD
O5jXhVzAoRoEoIZGYf3AwAFqBGXxxBOyj7rZeGIytA21m82GXVgnzyCB1mx6Tocd
vUiuRxQeOMWNZyQypVlBDJ/6c0Azmd2/1gm2Oi+dg9IplbLTcozqk0FUlltBXvZr
TsRenp8iZjbxafgazSxNhRcSw4F5I6CFQB0EHjehfbXqazxszlMjVfivPmG1AOEi
GnvFTvygYPC3DdDci1sakqalVwlO/A4dCSSCDvIjvy8KyWfgbMRd7nYuzM+3NUON
Qv4G6z214oZra40oTbRxaOTYSxTKol69aBtlV5KdTEYFJLWIYaRa8q/Y3pT8/FPr
WDvj8LIHdhIafk83d0yTqhogHis3yhfExsqRWE1TarGa3hwGtoN4JySCJyKsTE7C
gzP4N6SwLo4wquA09W3UjVJw5Uwls+0A0amEHIA0YDkqtFgOC/5zHb5GSHN6I+pQ
PVLjRXeS2reUTbPJkWRPxv5/IL0CbP0hdrn7yL6yowEMaPV9A0DiPCtafWSWW0/e
+mPBtlwI6OPKpbZEglmhEugoGjdzsiA0mV8UumeeGKSv2xN4dzlB7biIjKeVmc6W
3U/QzaCt42HGPmB1OZJKiqrD3E6EsDabUGjkKP0U6FzNvDBe3uut5wyHX5MBwpg+
6YVi4W/hoqXGLAhnSyWt6j1kSE1bv4N6QzeP0dBsn3r3kDpTdyFMvALW5cnXU3vp
bkV3Be8N9OIVxOxeFl8diZxUq1g9gbQtqUw4Ou7vU4PapmmvanZPrnb+VnXJNedi
+mtZCNa/IWm+LF4YR6vvGgDBtkqd2ajCoRezcYuqwyJAX0pu4NqAuXMQrkz0molI
rgx8L9rvdcUWjGuVokdd6ARFm/xoMmHBKr46VDooeP0fLCjT92sCSfLWDflhfzJ/
dfJrOPRsykWFQw+fhcg4zJ1HXu2W57ZQDCGTeRGvnu60ogNcS5bZYiFP31JlBFWe
cKNobnhnMp+3HTdsQUkhHeH4HTnMjZVD/QQmZHb0ljDELI9Tof2C614TAWx1tjHh
MXOdiXrggbD3tl54NIOk2opDJZma/E/b8Ze/9GNZTJPryr3oda/EmGGmEwwKsGrq
6Qf3w+bQuShWVKCnXD25Chq52AI5O9BZAHxdfjwcr0oGA7lV6zRD+i7tZ+ROoR+u
dJxFseiOjwX/cUKpHss78Ugv5Kx58Gaxm1239rEqyXdcs7v35ZEANz7Y8TLFdv7y
a+qJt1gS0dAHdw3KwBhUdCRtmSNo89r4sb4M1lDcmknCmL22qMrs0tQCGU2Ud2jq
6VX+z2y5qARbKjsVF2mod2BYQizj0RXdPEGaZbSAmCQ529xbbrH16IJX1LXSEZx8
YRsKGx0/8QUMHbMpuB+fVSWiGBnU5D+vpDJNB0yjkcrjzfIN5DhMoeo/BgmkEnA8
33Vf63SnX2J6JEBKAsEbf2QD3EgFE7nyeH9GAInXqwMHjwkdeJ0DjT+gjSKsVwVO
kICzbe81ek5++P5KEYgSnX88+X+B3IHAfqvKToXc4cJv3jNBbM24k3denYvGgLFr
GWdDO+S1uS9BfdqW/ywR7CqWJir7NCwgeU3QyQ+bLk9o4eyEb3Zu1huI6hOEraox
fJTyQajjefr5FtBY84AmBS6sgHy3aqmKDlTQfPG7+55F6RD277S/QECnf09Clzyy
D/DBuMLnamJbFF+9zAJJ/4tOJdbENSRyns2mGmzkFQyO4MKG6URGC9mfIQv3eTc9
Corf6Hx5N1QUxext5qjpYNuYZGGVrfos6PA6ZQvDMFudKCMP3MdFpIriuq4OwtO8
VEF9m3lwHGbztprufo5jneknRvOOPzMjmKSTzMgyhr9rU0U75TG2R4Q0JwOlOAhX
ErUQuP+6WIHse73sYIv0MqnwQ/g8sW1zt0Z/KVyyYL8tQ4z+2wVn9E35aJK2umFo
UqLuVgHscdy7ioh7m+b0pPJcnPQDezGvzg6khBE7hbXqH3GpESoZsh0rH5TL1EWi
eyw5dyP4NAn9o4yiyJ0lHhz+sOw59OTCF1ZkwxATM7Z4irk0aRbVdJuY9hGFnujQ
K7NJAJa+MhmPJQjhgqgbvBs+b4bZl+wFoaQjYEPaWlTzgNFYuQ5VpT3T2c1xg3er
UnzjQp4h/WtFcBvq7xAyXKHhyYu05zi8wID7uuWV+Da8+thDGN1+OnyoKo+KtyjV
CCDcGZ8tMjNseCXwUzH/2bPlusb3DSKXWrkrskb4D3xrnouMRmxUi+BndPJxsiBP
Q8AbRwaVpighLOWNbrsbIgpDZE/hn5gxG2Oy84S9EY3vbKlfvoO7gBp+nCSDA6UR
EW7sz8rdL7UHBK30O4tgO4fd+uMBe2DH0ncQOoGGCjci0tBhrpbeAEjSDIHj6wVJ
e+9aqGAHj92IBbvCITuyvbi70WbdOhv6w5dBaLGbdDm9yDRxiZZKqdcPd8/igcgQ
F9iUV0jStdRAvWrLtdcq0Ch7w4Uq5c2fVMghkRV55j8wwYeITL8pcTb+XMmfVCLQ
6vhUg1ge6OZCjuiE0pnpW52lnRNqTsq4RsziA5gdThsNrt8i41gGifkd46vVPk24
oraLLD6Wke7XrmtYC3R2VceYtAnzI36mM+5CNK9kBq8IxvIAd7FwQwSIJ7TnPXqw
haT8K8BamiAX8YNoBc9ElL7LI2+sdoiXhW2ImxgaKQfhJ9KEyNhA9dSalrCUT7SF
s4FtvAqFY9AF28BNoGkQHbl+iDkehA0rU4dydaaB35n3C/p4w23fYcOV0qTScYAJ
wYaoBCm4roRCweEirzH9VqHl9casDJm2TeuBgHiSVY2n2/RbMtdGPdHzFaqVJXa6
g/pXYPolu1OXNN674FuoZo3M5fsZ7KiZZhKBGacpOkQ=
`protect END_PROTECTED
