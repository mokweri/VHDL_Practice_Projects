`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yjo0p3N8YVSj/lfJbDQZv1aMn/NkqYlWyf1HPSwG0Cd3mMSl2lecwKS+Le44Zl6z
pdQY8PbSRuB3OFtRxfWccpeoIBx9fLuV1bo9lINIyZfVe8QPW2ZQxaeAIKbsGgUc
YLCfGdgRbbJEkgmz2QsyVEcF3nEqBtB/nEp4uc+2lbU2eYrAQTPrm/yfxyfQ4Ay/
UVpCHLSGkzyoM2IVQtsZ3ZX2Ym/w7QYBY/sPUdz6ipdZjHyxU3IGZF5tA0znkWyx
zbBT447ImS2B6g55Wp+AnFBnyr2aJq8Fs2L/sx5aaS7T7iDHJO428tiQCytq+B71
ariVwRO6HZkKr/NUJzzdK6B3IEu9V8gB9w8uxwSTCV2TPK6FECB30lsJ5paKp7Kz
q2xDht1RF22JpYd/5DwTlGRgBoR2waCTf6r301EckFCIa+VwPhO/gCfBNrktyKy4
4Zx4Yqnlo0RzItvd+sgpC4b7145rXDMZlpOEqzo1KzZ9wC4WkSt4fZfqTCEcDi5W
N9cUIXgHlInUyAQXjeRwdwcCj1MkR6dmkuKmChTCiczB2//JosNAPNJPgdly5mog
FyWCgUv8Gkrg9T30AdQWh+Jnxe+zxGD+i7iu2gXrJIAAXpZ73kcg8PsBlUd6QO3V
uL+3mOuS8I0N7APBtjnjE2ZbzoYqaYUbp4w35HivP8ORATOZI9w/AiG/QqxtgEG5
8ZKKC/YmBzB9X/rODa57OdRzzYWBpHcodmoJKjYLDMXHcGSFdRf/uwMsG5XfDKf0
hL7Yzu4mm1ksjHwo0zJlLgJVWG7Vfq2UD9PZwsNvm9Kq4Tf9R+XdGpRWLWpyWf+A
yffCMbqALR5vdu7VPF1E6aMRrkMfi/TjyZAxMGUeBO5OuiQ8OUKsUVqhySI3jFgf
a/KdmASOxVsvGBOapDbhQZTiF7b1s68H1X10fXGZOMUt5HUlqtO34/zCG4W1/WfU
nTpDZW2IYYjPzGGkg1+6P4Pyp9Uxuf8bKsTHD6LKjrzEpP3R3v7t+NdjOdb6o74p
CSYHDCz2MKKLr7mVzsa82N0PyNYqx2kk2WvY2F7zLAc3DF3Wl5H9HTYwATb6x/wz
VCJ49YZUwyQxt15pku9mLJLLRACppEk4eTDyDHZpoDSH4WYHVRy05SEJB4oHDAdS
1ZSrO+Si7DyNTHEUpKJC+o0YOmPuiNpMmtIkydkIrN/F4C2694eaEyxcX2y9gVMz
mhdhBKJNO3OilHAGJOl/2Pe9oKPPSKDElvv7cTwiGuLYNvW/XOdUNIp2CefSAWYC
EcFXsojF+jx0OJO5QoZBdlf/kt0kJwiWXMrcIFJOsQJ4oLjyovz8CU6IidpadNji
skG3InzD1uESJP0c0imBGHIMFYJ4zFwGDUG/Jd+FyYwBhrBxaBCAjPa1Qzm2TDQd
P5aQ2UtWM3vM1gsN/Ouxm1oA5/EFr/ugbqEDynQEpjKOANvQgfogUZs3cNh7zfjp
u3ex3i/5aufwEfTq2rg59/FBJ5zECLXmJkCUHtBD4EqSZwmAJkIsi3hzSOyHyXGW
2FqSpP7yI5AN/6sWVJH38jNfh8ybxNVcZ2K64bQuoRbaVGPQeGru9y9VoCvC/MMW
`protect END_PROTECTED
