`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3bv/lFPSwXh08evfWti1hsqBd8M43tdJDNiMKeL59cEaqoZV9iOQLhjlyzNeKx2
59XylhCqbZwsY3as0c5+4q5KC7ReOG886pPih9gkx92e+wB7FwksRCLe6PuNTCSG
zALiUY78/qu/bbH39I4EdZExC1YuLyHVVP6OCmX/okXCBsO1aXTkkKrc/xt/dyv6
Zvz2YdBUv6JnKLPJ3emlOH0R2OwILDW8iDwQ168eDE5DrxwL8zqYMewb0Jzq1qD0
SfDyPT2VBbzOLqS3GiD3r4w5SMQCLeQ2yQyb/8e2sKZDWnZYHjI1frBjsPIarLiJ
fAYKYpOhk1tTOyOhr3C+VjDQH48UrytFlHDaqUFblYhInEVj74rTF3UqRBvmiZBZ
Jz9Z/nEpYHJF4kX/z7ARE/vMmjamesBWMTPfv0eA1C0LkB/VJjBwZZ461Wr0Dnck
uRRjlKIwXGjujbm3DQxuckO8Ht3F3knzj4qyy3RHfjY0UfantnSNpn554FX0c8Us
O3AyqbI4CqiCC7x3N7/2rxI3JrOeeTVIqyA+/PVs80P881XRRx0TbpdXbMDqv8L8
Zo5zqUSXO2HCWqr6Gg1REfOO1yWDurG4wP7N7bMUJHOLQgvoaWJJZySSflq8QrjP
MXbAbnQZkYqQNtOKrQ0F0jf3mrKU6HZOzDmPZsdjhmzRha+x/rXnmLafhVv7y77X
aRlqLvNidr/yS79F2d6/IVmzjk0NuzaTdg/7kW+Bm81zUB/D6GqHca3Z2cQPINxS
B0R481efGFRqCEd1TZTjkpRe2RWDzWwZmBDQ6Ep7dhAWdo3Gy9bz8KsvSJGOC94I
NArkCoMuf5ejiumGEKTCVxwonc8iMLloafOxZtnepXTI4LuEYwwjPu/Lx9JiOGLT
uD3nljVcDOmhBKGoR/pIjWHn1Gy7UC8lLZQ4dFkq5LRu04R3JzkaAExXWgG8haVq
daXdEjCS4XsuxnyA+L3z3eDNLCvbgp6sDOANB4ObOPgrLhMc1FAFVRimYa5oTThI
FZZgdpu0e0PmSBzS/kzvwG0u7zoT8pAl9M1caCv2n/2hEM2g9RHGPsoYa8iyfJTC
EavIEOUOlRyVxKrYmsUemKt/48q39JE5L9ieXUq19O1RdeW33SBVPEkmaDoLoj0d
6c3R2XDFcEETQgXhtsh4y4UNOFkh9Z2ZC4GCzo7JdDaQOEKSMEaI0qekWo92iYUe
aSux0XMzJdcund+ZCrPbndySAOD6VPtJFKbp++fRUxtVZ+3HjfTlLpTbDet3MORJ
YtZud85G3R/DhD6bDNHHg/oKuzQkLunMfnakzL2fLrEoQyZVejBOXAll6qB3bYzj
uwNAW1+LE/ic6I4dvcUBbKU8drRgxu+vTeBU3Xamfv2IwH2c8tMmCg6nMEfqf3mj
a9mwwGlJBot+DlKxZsgewT/L0jxRUNbHKmZ+E1vzrR3EzIEkVVzRFUo0vyBvnwQ9
`protect END_PROTECTED
