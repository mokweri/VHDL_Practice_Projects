`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcxAJZpD8uJbwovX+2MGM+UBUEBpqtQPvDUz3UbpSt7dBb95ld439QW+V2YyStZ/
QRyp4cFzIXIRZcdS0CX258q+Q390lsUFr8VSGz8ZoU11fOq57QJ/4JMKN7/UCbHi
SpJlDYl47pKmkGtJnrQVLBQZONDxaxKdCmYO+KbQE8lQS4ur8iOVR0pxpPqiYYEN
6XdrJiKj+TvKk3PEvyM6T2Sf16oc8aPZdygM/Yi/GgeRHVabuoFfB+M8jDx9yBr8
0FpY7XhytKBw0TeL1qiFVUVkfjYr7QkNRSELZVIkQ/mNWAKh5LtElNYSJF6UizoH
pXrfRFMwlIl5Jqvco/cvrvZQaNvqN1Yz43c7vPlReF+4RecYgWzVTxgJ3ah0VHT6
kpWAv1n+vqscpyibIXD2qAtEWI/AoewtsDloKSHy5WC9biRHEo3QzM8MB+N4Z6pW
b7izxlIvTHPz5TOhKRFbV99V4oMQTauJ83Kesb0YAaJMYinTQUzvowYt0mGxWAV/
eW27a259TmckTNUX0d0AURY5T+uyg1B4dt7OedT8DlkGmOO5NC4+TgFjM98Nd/sf
PToq0d748stEp6dK0AFIJwMLmtLmLz34KN7p40yRchjs28YflXHUlZRdrvn+ZPC0
OBks9sw6cLK9v+4BC3JkUiWrXB4kNWyGE5H4ZSl8Q64SeCDxll0hn78OWlNAUN1m
2B9MERPGLDinNaWuE2hAxKCC8Q7qJvKK6nu8CiEp7QivRQelM6oe9oP+oNekZhRw
D0WAmp1eKNDhM3xvSNSTeKt/J4HEfnOdQpCoizBRQ2nqEkl+Ou+1Tg5G/5oTbuG0
4wxfEMoaPfVH7YX+aCIUvmErgW5E0jVUbUtFaUp2wu4bjpC1Izk7SgwQ/hrttaqK
vE9Ssq+HoBAckRy68VpGsUS0yjDCIxxgdHfVyGmVZkuDp5Ugii31o33USlH71DDs
AoZXpC0ukO0RvAhQd5p8sjPw6/P3mOK2O43etSxlkKhZiAD4WMqJVT0zMJb3h3Q3
y+p6ieodRqhH1SsHYnp0kIlHFUYB6I1HEIjMpR1xMFif9HwvtKGx5+c0HjC7de+c
KfOOdUJyKuQhuRp3qon5zVR3hPq1qBhTJTtyTSrgJsJel6Qf3ROgonh1ZlBr9WlD
ke0jcy5sC+Bpetvkf1vTpBYxxzf4SEw/sVw3grZ6cbpLTq1JehEgBeCDXvzysYQi
wGCCKqK4HVzsL/jwFL4xunPIzMA35pJOjxZTGZb7+bY2fZxy4dmUfb8mxG1DLQwv
`protect END_PROTECTED
