`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8bqRIDhS7wfF4g3HwwY8kf9YMtmhLFyoJlIZ/0naurYtldUcXRfEJhv5AZtaAZo
m9FSZYeepokdAGcKum/wKtixD7P38c/V8pKjW+3qV83PYBEq9gfIocJzcsJKEF76
1XzxOwdfCpcI4Xjppz1XJcj4Q9O5kxC1fh33A0GIBc10yqfBdMjqCxYHTLu0PTMT
2rHOx52c26BnqWde4XWhmRL8ePlicjvyaCoxz0MqwL/UZe9E5H4SAiTYNbSMfRjN
iO/rhso5E9dwx7xCGHjcvai0DBFVPIZ+ah9ei8yt0yKA35oGsT1ob4vhmraaKbBy
dbnGixdAXxvunxLvLzbIPeiGustzzrIpdOLN1NWLD5s8WgR7is0sIN7iaT1T6VSO
hGL5v05tmSV4r2KcvxcGOuLwR1zaY4EcZkX/UnlL3c+Ssw45WX04LyJL5vJE03d6
M21+BNAHssC6DmdOh72fuFWL8xDdTRd3O9ljPeQh1msHNIYknjqlD4GQlJrXtnD+
ug0Rqs2ILsI7ZZpS/mnbkNRcgSoI7DDNO0/WwGsXzZ3paGnKOMbF5uc59Q6IezyR
VYS/rslSLUqGFeAycRH+dgstYc8/aqUm6LXTL2G8pAsyfahXJ7AeXrLK94DP+UDt
ahxl1S8AFAeKxm7U15PreAVuUIJvZEkYFi7TkHCUIQkse//ulNJ28kv6oY+1LFdN
nJeCnBqCvHlS0/vvgcFYqbUvmZ3ZIP/kDLvLmOkcFL/QKGnNbS2MJlbAP3hp9yCs
S73f/lobyiwAVNjYmHFYc0INGTl7tF5YfL8E8i8x9oap6v1pvH4HJvkjnHKOCpRP
b5E4urtkkGRgZYy7ddUx57lKZOMEztituOKBA28HSCS5Q8VcybadHMyTylaxP/B5
HWb3N0FEt+/tj2pcs/agsSYk/d5d0h+PeoLZz7H5iGCiI9FkC/0n70hyzY6KIpuc
zJURG+AHTiQ1glbRL2H6AZQpsFBHz/wLFx1bXGydgSXIXJSwEFgxINdBjqEoR23z
NHov99rPoUQW0cnXupKhbgkoEtFT0Ki1BAjr31616/bqdNhsb1QQIMhd1md813IF
Qf841YoCqfiQ5xJoyo422S5Hta/GR8FQYIaFUwIKW/ABdUXlh+ALiAImlxF2KKSb
xOt2HHLJgKjepaRXFQi5sOyf+By+F7ytPTsQragTzYvvQOEiTdSchH+kDvMwzQKg
UsvPU7Al6MGVPKJafiI+CeVu3Bb68CaKsiEXVyooDXQJ28OeRKF3RfLGePGTl6BN
+KtC0PdIXQ/q9n10v7TUs1vMlVLD3ZgvdohPd3/8qzRWASfg0ftNx46/kPe1WDb4
nUtnc2onl3q4ZImj88uyAzQ9L6u3g9JXMQFyAewK/bS0JUe5GAhl489fMfu2leDo
gVT2ZvUN4FLixpv/uolVbE689S12xp/jNvoQGmb2p5k1trx2OyvQPTodJKBoaci3
MK1S9SpABXUgRjItmrX6qhd7Wb5N4YpXgR5Z9QzpLaoH5Zp4haAguXmR7yLGMPyl
sbaVobupQl1Kt5na5dLx8k7yBal6KIEtCacwo0v3gzKl67GH1QrMYT9DgPSWrn4g
0QKIKr+dY/HZBXq+cdOBKPqfuoKKHcE0kT90c74hhtmbkIDNMnD3O3PE5vsIY/cx
ZR/k0Bil7W8dqxHvKTwCBnHtn0qSNRyuyZ/GPuWYwaQq1kDDzNd5VEG6tBWbREbx
fHJBrrugAaC/EJuer2RR6wER8nb30dPcQjgwld5Y7rITRYxecTm1PlXXqALN8pMv
okH+bZIEdnsT968mkDrA+dd+PGO2JX0tiQfx4BqYkaz2o2DoS6J6dKAcu14ppjak
uPKTHcUKBWL+T1zUJWyxocr6rOYzJacC46g52mSpum2s9lagJMk5ftvjms7xjEKW
eHFAv38Bhrqrcn0akdyfEzhZCYoWPam2rcHlgBYrr158xKTj/haSftAl4iykhEcR
aL6aCz1CQjB0gWOWblyz2OU8GFg4Ts2Y8Bqs4V9s4eQH4f2RHPml3Fr1h7grOa+Y
ct4y+uGnP9GNi1wsoepeY/4p8Gh3pSZQvamaD8aKLUaAPLFyy4oj/v1ABFq2sg19
ISg0TVuGQtj7M2EjjuKhMgyj5ZEYlasAc9cqg6QiFPnGeZ7De1AQGYfAho3qm1yr
MboAa7RNC0eETb1OEuJLXU9fR/hbbC7O0Yj1Ie1Fnm9ZZQwgDAdO3MLM8vFYXKdl
EQFd8/5lIihWAat5fy5eBusITzyO1c0E7vTIxLoOlX26GXtW2cvf3hfvq6w8D0Mu
SbpcHT8hYzIDGjrFYJ9pmhL+VO+2MuDn4Nj5hjHPwv507VyegGeoH9s6QqPIFgEo
349tt2LW66BAWaAjmmR2uQzYdeLmPDUvWOWhNV6lO0FOWO1G7dW3n6kGjP7HZ3p/
3cLYyvrNU+9yFxBDHF/9xKeT1gUEl0W+U3+L8Hc4nTIFZh3k4k6/sJc2K/fJi1dj
X5PR7p9msc8cmGnJIaNzT6E82soKpPAcZsm49Ku6O7L5PBooO33QC4ODmwu5UQPh
VB9E3KfAlPzKyKQs16/AIGEx7Hxg5DClXmCRaKDBWi0f4UuoxrEwIwL4b2+k5zpz
TPYqrV6wpAEUHE12pnFsotJ69exMkD/iyUzW5KJVzpH9OgA6vo+NGMfAGqv5kJPb
ylwvl+JaNXZ2+nCVQ+XAl+u4I9IEh/WuPPtx0BHkeTtQDcoippEhBPL5N5vrSjcv
wEOQMw75aoJ8haY/r2IHr+7Ogde83IlrKIkVxyobVWWucPCpLmKlYSxAoQpU7bhf
GKioTd0YFttqebT5qsirlxn4klE3gwxV3Q7B3OPR6uspNIkqMBK4O1qQPZ83LO5S
cEiNKsS/75FcZmAfhLJjruot3dNeIDLjSBPTOPv58MUPpGKyCH9jUr50LbA2PXcC
mZg+frAw5LyRSNeISxeTvH6j8te8hPUEcuDxLwHR0K2cgPODSmtmerSEirziBwfw
7F8T8bmYG49lT5JnjgvO4/1WMe02m7FYZNa6bjgfeYJV9+9Lu9rRPkQaIjO+NtDv
AJZb+NCAl+nD5whAwTzAwz+iDp2vvn9m+y2bTLJE/el35DDB0Nq0kjjX8TpPWA+R
ftcq+bh7FIYVro07QaijQ+CqwH96FciRLWZNhMQipFkY9sXJgkROcQuhcupq4LjL
+CztA0bDUQSMHEfaVj1x5figmK8/XwueTEQ+Qj/KhqYtR8Q3HrYtXYsEwYo7ytmd
F6JCX1Y2WKtGz4ZU59VSQ7bBREtLzJWWtnrZAodU3fvnmJwq1VmmruNxWA8uGGpa
osz9ezYMgY2duDwMcuDfd+zobgjNSQr75Oj2I3/9d9uMSW89R0YzYbN/Lzfa0EpZ
EUAPZcdyXP7Bmr+MC8c5lSUxFKCy31e1ZJyWofxfJ+8PeJO2gwcuNr+HWi7S8aC8
vaq8OihLaetQLcSp9enBoQDus3gJlhCRD7U+oEG2/JNEWyV9V9+XxyVxyJIgwKST
2DwPqvBhDKYXn5hl7jINPrEaGxk6XxIJSrvTHV86mQMHt1dSs3byT63y2l3IfhFi
6TASmMTBepfSCRdqiICpaaTJZ0lJtwFsoB6etIpIhsiJM4PROfz9cmKB2EsYnh00
vTd6YE0ek1uLMlhO0m3z7uUCpfmT31UUOXgwqET6oW+EWiBSyXNJMr1Ppkw6HrZO
bv9ZguAgTFYICfEh490QYCuNmW9X7whwrc6bz3q1NaiAAT9s5GAHb2c189rTZrVe
jIRJF9jepgmppQazuUrEacYfiehtYYl8VRqfFXWkqouHnPUXQMD+O4QAC+++2HSa
lRGw8GBwrKpLQmvKyCokTtP7FgdYjUfEnaJWXYXw63amVsoIeUpyPL/AbxRS4T+I
C03ZALa8r0aMPy9mg+xW1YQcERiDW7JtMtGNSmPFjzRS0VCH3Pw+sTwDMrq9U7Sd
mmDID5/M28ldoZ5d2Y1bojWctyRF7N4QSqxTcxckDyBbJAkQj4SZpejq5GeUvaEF
nyAdQOy7ZFII2xKQ2dY86Gz/tKeNbxrpDsixcWHWniz535WZRoKqJJMtQd2PjX5y
QJhhM97r9rCQf0lwKECYdF2fMjVjE6M/65yChDq1Q3YfrsHT9j5ztJJbVaMq94H6
sAryuMm/CIInEckLQfoQLM+DL3Ik9ojCgLM/MgmaPeDLgCcMAJ4BA+kSAE1pCkaw
38PULtgWlkgZ7MRUVJ6xrhmo5bzdhbZQPHanYHTtbs/9Pqq8gKUgLsYgG44KSgPx
gP3Qlb3eS6dQDxOsmRiVTd0hBxen6dLYFB9o2Sz40V0VwjRZZUouvzpMXzf5ixyb
vpbPECDsCtjKft00YmW9dULkPOsffgaPVjICi1rpN1L2AT4rqBSNbXwI8mEqdnGO
hlhXsF4VWhATIvMzpo52ps4tNOQbhGPuXetzKwsB1yqKQ20Bqo2IpHg7uL7jO0FJ
pGlmgqS4nR7DabRGRr3A/cNe/R4RboiB7CpKugZY1uVlanp/x1RR0gs4awjQLVtT
bsg1pftEFl/gPyspKjJMfQVhSIBwok9H2J/mxWp+fVcIPF4opmOJhgOAEiRvsrMq
RR8zbQufyvlZlmPL9plb4lFpDnyuaoaQXITPrm3Z8OBfqeAaasUBVtQBy4z/qziZ
nBDRbpO3mknqLk0AOeN45z8rzMojFvWRrWn3FngqxKKEHXUK9dBvjN56V854Cl8c
vCphdKp8RIs1QbiEzjNqu5xP2UrjwR6fYHqc0suQNHUzsi/kCEwCXGnzUD/luQ8P
NA8/0WMBGEtFxdRRFwHqJfz7G1/seaDqPa+5MwBvKxQ4zGQyE+WScsSzuRwFSCpM
cwNEwM3n+O0k22OJoa8UriBt29QViylKIVV40g/2/IE9bcENF8CSm9p928iatUGa
Ol8AguCGsZzmYetAA4W6ZYfRUTgJMB/ItI3E+fODZiRZJfwEhJkUxlwxPKiEqD0I
mH/arv/l0Fn+rgDsn4aHXLUM0mmfBLxy5c81ysBccG87IBqMSzRhYwhO+6HH9Zr+
F9QqnYJBMDKByR/MTQWr7oLLzjSeV0qQvPRfJIsMvHBPo862eB9bw1vn+DiEpdnf
ez5pD62w279Oiu5lZUHYmdyfRWQmsVDu+9fAg2OXhj+2EZr1VSEfuRcva4EmTSfb
AJxYz1sZgRu7637BNKncHEJM7NdmcQBDfKEtPVYMzHGP8PAu/tWzmRSWDCKKpGfi
+3tzVScgdR3Z9+FTXkim/jQwXAZ/QEQL9uXIRx1lBMg4WiyT18cFTZSCpTgoac79
srQYy+eeoy486Iwx3ABrH4GLaa1CkQwLvVVezKNTNIcHViuG5nULY163rQYiaYKp
G4BbdjKll455oO1gb2hnrexbSRzdlaBEfekoPXXB4KNBnCdzbgElqRW7hFpBdO6b
wp6nG8bmxmSHZMYHJNdabTe4R/r5XgMLTLrEEaxcDAMC1gBzaW3ee37OWZXEdJZQ
9wZziLtNhspTFUDKb6Q5X8e4M+O1KK40YaExkVGlckrtSdiwuqGCLraZ0eLBoX+Q
r97UH2Lj3bUMz2P1P4FFu2Rjb5TQ2Uc/PsJJs2BCSJh3wYirBLkOY6oyQa7wCVXN
RTGxbc8KSZu7AIbkbCiubI88q9NklzV9hUCkQE8iouK8deuwtKIHRK+3hfbVm0ku
JbCcMKWrCL+s6XBJzvt8LDxsUFhe1GZj1aILaw1OuA8N4oucE3edFsfzpTI+EqT7
wqUsSSVoBNrUpBYVKcFqlAm/Pp88ict/KrVq0YVFpETvHU76qgnT+MtVUjyFaebH
8K7OgIYD8jEU2ElQO/TpjB0UaK3sh6yi387E7uei7zsDcpmO9+lNii0pKQ9dcyHf
xtnJsrauyElqPHKdd0oVFoRqEBp6YRk/+mU8ZI5v6Vx/kIKgnGt7tdoqoe/3VE0I
SqZxccAvlG3VqbFnNdBx57+mZd/rAZJ+SJ+B6WTAHvmWiS737Oh+0G0I8nWMYFzW
jbvdFfZ01fyvS7Kf352dbTej/TuAlm1yzd2ZMXVohdkgtizJI6aDJwlRjJeeiFdU
69xh/jx42BMCzAfhFZYJ+yg8DqLUZlB9zGgxOtkQAbmhHig8zfwrFdDMVnonIH38
LTlTIBoRZvA31wXM7Tghjev5zq9fK3jLKcPTL5dAQHP2Qbhq0dtpRe2NQycQgzAv
9kZZ9RrW48ojgYUfuEWz5W/ChBDDVx42zN/eVDF+eTck+Kt34Xjcmk/uGHXBv8Ex
irUrN3YV+BhbXCc6RxNOecrgvJC5IadGJTehnw8rPyBS6aTNSwET0BD0be2uCROw
Mr0WeuQ9SR9hL9el+T2l5pppzvWaNEzfwLljI9cXf6c/dZRYquq1z5PQGFYyloVL
iMIOAIGBYfS+YSlWMPUAQO6PXLT2LX6FZF917voB+oPLVrtRgqWr79nS7o/HSxt6
uoJMCccqT6l1bmXOzqxZ7o0QC5MfQd5cOMyMITBVUgCl7v2EOvPJzY8f1sAGm4r8
n2wG+Bp7v8TVpW4N8i6u+h3d18qaQ7xQEJIAbA+GucdbiE9YSrfcJ4I7jLu3AVVx
oCXZJSqNwMjM2xVkzBEEvJYOWp9D9dAR5vBe2kleGHzTPLCEoryYaByiGeReoZRo
3qs1Qlytfm1NJM6y1FByH3f4mDLeMyT+Z3AFoSmeoFy840bagTJ2/VcdZxBdafTH
PVgJy9zOs5TkX/DDLvR4tag05RYomVrPQqfvduUDvdITe6zb1wAXc5FNAdtWUwLb
WrfQ16pfLYV1jqodcNG3Z04UGyNV6fuWWcQFB/mSQHul/Sfs1t5u4wi++QwTakiy
w0muUYJHIPz/I+OvpUZWxHwXSOaHHEQCc7Y0ejUNZ7HqmmUlkTRFdkZVADTwiCCK
ZmKArbxHkDjtiIYLx8MWjwn33tb0/CPlRdsMmYTTiXEsj1HZceAnCsgSmoj/a7cN
ONwC4BEsVo6mZxWkxwN7oLZS9lGi9Pd1rx0MZe86chB6W6e/dUu91t45YhRE3wJb
LPhMz23JC8MGMLUeoTwWXyTiHv5o1ukmR1Li29KFWOvqCAR9Ut0DtsdO13ZcMFbj
UgVRGoRjn+16ROJNVt1GiRD92zxxbSup5eB6byR9/njgP8hj0zNGa2PV5SoSpEgE
etBhSoYa8o7VUkuiBa6qxFfQ9QLMlKFQmf8zRUKQmHU1vDYA01M+x7wdR0RG4LU4
/hMVE1b3RWMIWuPTGUL1nShnpYjtictEk5SIAewpnil8nS2cgulJ+pqhYuy7HzKp
HXTL/EYvsLVlzKOLKl6na/Y4hL3WXWifdg/AcRf6YYBFlqbLf055OZRbv0FKf3nJ
J5igGvpvHxiHGiMaJ5V2GCACP2Nvhey3Fbw+rJjfWRxKfKQDtCjvuDD+wvKebyoz
xkYT3j3QSa//5q4/EzMpqxQQt72aG6yCd1bRYAo1/rYDQClq2kIGhuRTGuxhHHQW
8YsUwfCyFS4vznWc1Gx86sYt8b+3I3eDyVtg5duATOf93dwf4sMWoWx8roE5aRAm
0IqeIePNVfhavCoCtish5EBYgz3vrOllaV/4/Y4SjdjZXJjdk+8xREKqahtIkKoP
3cv+Ovez5zqQJw5JhPjCiF9uTVSpZM4JUsbzc0GC4HD5lZq50RNDiOFutVZjfyk5
J1uxGverHGNcyu7eVJI/Pl9j2r9lZItTheUIQCObzn+T0l3aMxf9UTr9GnGz3ive
rMBBYW14OqkPx1Ti8AiD0NgxAltrSijoVwT6ra8jksp44DFrdCFUSojni5hBqZxj
briuCTmxyd6BIWKtwwuLqU8d1G+TgiJ2qSAuUDVQvb+PQeuDW1yQrxFBEjB2Xepq
iyNlFoorTpY2uQlbBo7pygG3emChFMoSkUS7vYgU6NZBNNZfrcc/JSKfaaVUHNse
VIHBhOIaAl+tRX07EErtPRQDKzU2PsIoBGxkmorH3SLlE0WvpF7ToxYDMXU0TN4p
geggtI8+y8y1oCfjPsliyKpybWJyW33W9v7G8Smc08OHRl9npSXuwIgbBHOugmo6
9iwFRgOB3amT07naWltFnMO/QEXYeHCz/pDfXSrj2YLt83+NW1g5lnLz8NpZ2nEU
KYKih4+dLC1T1zmtWJc99HgI/DA81kGNoIcEwnN8RZQhY6w5r+aLFWwXvsxRdr6N
pdabHoVY9ujhDgGUJDMjFcBqRRJpZMFFaBmAf1LxoeRSlL3lW/iKBVk4Yh3toT2p
FXcYQj+AHLl8bJRSznmcGDvziy3Pt5OUr2d8SmXCSgH2tYuw7cav2kNJioN4U+pF
6yj+LKI/sP2hLFEslOavGoYMuch4rQOjnUEpTPnUCqy3IJWoAcsF7Vpr9IdXQiMR
NdUMhb7j4Pu5/CYgyHVOyEsZgG5X/M7XUCTHwWcTsRyCATfGRSERyFF0+3yen56B
7OMzkdrmn6EncH+s7mHgs2538Ox1mpOmpMcwOxufwuHf/2nzur7AR3Y9FHR+l2qf
krX0BqQp7E0vog0tMxqb9/fs4VuWhNUX2xR9SJPb7B16akjq9ajcko8vUaczl/KJ
5DgH2Cs7ldAVoPthojl34/hAJgJD0IBm9vG2otVB14hSsGJjZEIwyqlX+37J4Q/4
PkhMV+OMtgkSQ7vP3OznpQSrNnu0RiuFnZeXB4oNidoqmeenoWeBAT9p+1J3K5fA
gifXY/TZUmtER6yQqGPM+tshUhxHDJ9cXIGKZ4uX3r9fKU926nwQKZcIKwC674Zo
oQ0KURUJhj3cRVRz4x+W8yHt60yD00QjuFoTNZxfn6+cyZO3JciIyk1/RnLN9xdx
/XJG0LvxatpoKw/8WiZy/+pH19NEUY+Kr//y0i5Df7qg+4bBmNwXOqH7oQdt9/M+
SGqwtspIIK0ctgSsKJJ/fkB/Rn0wo5HGU1huwNalrJ9Z1MNBiEANaKeNOslGbQI3
n/JdhtTc53PFEXTuzeVTgTu/V5fdZeOM8TtC1DbEsTPpK8Pw1DXkA73RA4/5zSJA
izSRiaWXSToCy1QqaK8xG3PSYnVx67cL/aanqCqTJaaPvUby6HFXS2/vW37TUC/P
Rs+BwSclujQ15ysrDZr/nOHFuS1MLG3Z8FA7VKLuTRm6+7L1brk2XsfAWtkGsz6W
mZpKC94YIHcFHwna+Se1Q4gYkcFrZsqH4703Zp8QMM72AuBq3VN6uVSVYSs0sjzm
vfYwfVxTnaWohaPkaAF/T0uP3m4pijg6OHYtmeBpd7usfeQ9T+PzPEMWKOggYFwI
4q1RJq1jZjsR3QoBVfVNbhlFEDFyipt4ka7DZWZTNSUeOMgiXN7/ckxxRT8VKVgo
c46+v1BUfzBrV1BWhg41L49fyw7IEQ4jFwua7Q7vlhrDGZC+VMcfsRogxSxO3fyw
5B92DKLCyTp388XzxXchVumWRSLFVQqgI7fdfgZGANrU3yvy0zrOOt4Gvzgm39QD
5Ec72Le5Q0A1bXP4e2La5GNZLQ31JCu0qQ8Yc2qyYZJMgHzmJMqw4zP3iJcZ2m9v
jRQGygNgwcdDF0whBb0U+S2eECCaSt+PAr0/pqCygBz1Ah/Of/kVYHsJP2DXu1Qf
Hp4GhcceNdyyckdS3abfGMA+Bs/6KMIYRI1f625VfcNp5J05yC9yZj8y9f5+Goke
ersG5DoHVUNQWTYH0vkkmv/D7YEOQM2h2YGzOOjBRJnYcFN+LEnhYfsO3IdZU84j
+TAbtVNwqnkF0lKyjnHRnRMyU34AdeUNsOQvex+xsc7wK/+ZeRKmfQz5S3+sGcjR
sslAufS+nJq9dgwn2xmnwnyswnE8r10I1Ad5AlKgtOvCIemtr/74JjyZuZCyNhmI
wJa/qTbig41XNVN2Kgo9UHTNGx0OGiTuDKySbHNIv2iYHN/VGgBf20kCR5vEWkXE
B1AueAuwEJn/eGDQH++zubQnvKrbxahgUJcjc8b57YwMQBYg9EEQCGvMZOgHNdhi
wh79ABNUOt4rzpW1YDzVspNd2u+U84EVIttA8FDLlxZFT66fvZ8ba73IViMiz7Ap
e6o0nepKtLM00HuXKE0rAYp5Na/x05VkbLr4H1BxMp3lyFFYR3Cx/gMHAMbvserQ
MSdwGdcJhg+Jg9SvYVH8QWRI8Ky2oXyeUK7RHmDw0L/sB7XEvob1L8g+fb7J+4JM
91ykzSmdM8KQ7B+fPxRMYSAU3kXh0J0XNOgrO9whRqaflWywRPezYtTJskx0KmuH
FjgtS5vFrap0EWMgMs5CelL7fg8haNZZ1yqM4Bb+5OH7TZDYtqZQ8QiRoGYdhQmB
y9gMkBDVj6sExWACXpbBYp8iiZkXRBuHQR4EYKCq+oNaMEze2Jz1K+OoOXmHpF7B
lYLZLv8t7baIwYeta0DSSm9Rl3JSYe7wwE/KrkAS8BvbrysxuFbhwJ1SKHq8NU8e
Z9J4IQ/P2yEOPKav63MLZziMXlfMUglU4MAqjbiID8cFo2FOQJg6sjuFk2GJo1yv
rCB2pVMus17b4JyYPcR71MYNtHA5yLuPTETCMuMagrT0A6zU85SbEszQwixWojVa
BLQPsUKi2/sYv39gmiBhDUurC4VYddkx7QWefrgPg3tVqk2O5v7D3PjDmtFTngn4
PVf4KcE7+05oLhxUoIxEPOYIlO+AA4Rct4HjEr4gynKqgW8AdSvNLYo7KYPLThe3
ILmDAGDTUE2J7AQUr3Gw8CCWjhWN1LSv8k1z7V4H2SyA7ajl7JX36gqqrELxtqX+
Yg5sMkTGA2cBcBwQfO2PQeC1WmvRw9mZX+8op9q65ExPZ17X8QqnumdZro1JODsv
FKtXYBB4g0QMR2j4AZ04FhVTM2jCnYUWERfRj3PqhUBK+t9xg3PEpYBpZGNhwwVo
LQHH403HStTUJ4y4FNKU4gr1SYFG/3VHlwmvhVBWHqWpsFebe1bjSKrIdSiXuLu7
IwPbUH8eYkzWGiXtmBWLY4qrgrXqF9tMZ2gLXNQCY+r66Rrdhd+JGOA+3Wr4l9b9
ct2GbmNKUpjFPKxpLyn4UfL0b45iTrEEBJ/UXy9L+s9MQpr3Utf62GvXfxfvuhLR
nHtgOlilMp27K7foah3rk79qa+XLAw9DCJkN6Fj67vMkbqUZ5LDlFsrIvN+9I6s9
i178Ds77aORBXXFcYvIZU9dddi3lPW1w9Rx4b4PZuR6ZglN7je53UzbTlVYjxh4l
zNMZRGB5ObRPbHzPgmeV5txK9qYfxCqgFbWc5SLXM86MOKQ2ZEWoEtiZcgPBfCNh
awJM5JUIVwANDWT1YEuf6WoONyfYCoUqjW7Yl6O6JDoz/fPK1Rw95bSvM3fXbnBw
zhdhCgaHiJleuP4Y2QYjXpdT/FSBGerJRJ/NXaWOKLMUiO8Jjy6uMIADMIPfXtsa
wQt3JeQIbkU70BSPhEwkUbbbmf/z9E1NwDRhsgQNjW7whLAFolqIYZlxiwcajYBA
sc0Q/us1lm2Cs8VpunXTBkNUazhzx3Gp2MzAxGnt46ef4L028DEnAH6hXCrRCS53
/3BNmyWwdAMrtSIQ0vNJjNbGWJHywu+B9pXhFdQG3BUKZgi4F/Q9gw6kgvB9QdwT
95DmHZfwqDe84XLqOpx/6piGg4vAxJZ9h5mhZnCAF2GhMGNUtqvSovzYf1Y8pp+H
Qn5Fpf5mvqeL0iIb80Ns++z2bMxu2dpRrb124m0m2zDcQ3ytOmMj9wpsd36M32fl
c2t99ui7rMLggO6gPodFsAaNYQQ0NNgS8XIjEL/MVKETlt9KfZeNxyHgoCYmlElF
3O4mM8pS6trb5+QNDDIyPHZJTuNBA/lLsfY/dhAnACIIrcpDIr87qYMHDRPQDs7M
wRJf7Aw1kXlHY6As8AzeW7MKXIHoqR0zqcaCWhuB7460E4yEtB69ZPeUE0E//6Hy
oHXFWSrHXUMQRc/Tr++q2IM0DLugZyywap7JrOGPkzHJyscPTpx0+NCFO7tGreVi
6fEnwQa0Fq1OM7C+yHUinKnkY7p2aNgrbZnAypy3AFD2zO92Kh8Ijob4aDAAIS3U
CQ9Ys/wtqzIH8JDw8qsrhbTij/LC+ArHXbhF9JfFH4DrVg7K0Y8fdgh2SRePne6n
l0Wt4eoZYoU7CFe88wHUbVFU/pVO9epXbSQMkzHFKFIMebrKAvfjl28Rc6FN0qYm
Mnw8Nseh+TuvoSuDpegalxS3JrAmr36cRRKQpr8Xjor6CD6v87EmLtmddUPpSe92
BQBjPyg3Yp0pcI5NaQgzbHmMLr2NFM/To0XZGhS6bzchGWOofpDc6RlPSv54dUhI
1NF0ixseG7h0fokHhZPJIR4L0P1Ba/jxNDyRp3Hng1XUQLihfpgUctnCitu7wqA7
q8IEgUDlO7dsr+c7V2LPoGF4YOV/Ei5+4UTnphlkr8XOKN8+3FrhvrlftPNhoFQv
SVWba3z0n8eLZRaM7aNIraURAZvgefjNf7RwyOpoj0c+uZ7St4Kj2qfk3U2nDuHJ
Aa40JtruB5bnVjNh1PkmCqZNpmZKYT+JOTvSU4GM6Huzoit3f87QB0cGjQHdvwKI
dpZd4loC+7SlpFA76qYZclUVre7Vn8S7DJpMOKE84ATNpVHH+qFkk6FHEdVHgfZx
JQZifdfKTzkeKx5BsX5aCEcnX/lD/vnH+/waFnxhPBkTytQEQfjUI6lu7h2By7SO
GSvSDAIP0i5fTK60XdfcdFWwbP5oLmaOyEZICCeblon2ZC61XRTjeEQo+tYexNbc
j3EnXh25NaogOK6gXmhEoz7YaDtZaRYoi7BdoZHSbyE3cJH+1JVE2gnTM1QzWuoL
QLBLfbXOaEqNzlO2K8p4IZWZqjLz8GousVtmEIC1QwWOVXtQMyXivERNxULFzVJc
HcB1XdIdMnmNCHV82TMPUtkeQLK4QESr9UtBn3BgdH+9XurmcK4VfncgVoeBWjox
dpybcE6lxpJ1l7790V+LGZzSjCUi6JYeE3m8kn4o8D1XtzRkkt/1txEdrMVHP5KZ
NrtaMMSbMod0X798NZ6WArww2o7VDdFcnGMRKSGZSsuUtd2JN2uk9AvjWF34inTa
PUxvK9em+RZdNq4Jug0B/6ZhyMOXn0HDrtv9SKWGZ81MuXVvQ8OvTkTE/bUab6Fg
n0yEld/I0ey9YhHWdMcwSKZ3f5rQMVxk5O6xDoeMPjVeVIWP4HO9s+qINdFv7J04
JHg65f3m6eqxM9rocdaLcppfS4gOUx7Ls3P+ddff4tsrCU2zU/n/WQhlaj3oajcy
K8/nLCUu6GbTIYC4q+YWNJQka/yXSAErRTfdc7NTffEWySzUk9PGuk4671Ltp3rv
5aRd47ECvBk0/nHv8D4IJ6oAhhDh+KY+jC0/ZCA2yusvQPlUYkAwAG+z5XTEbQfm
M78LED9UIsP1Y4Iw+e8ClZ9OPVddPcqA2c1FVgYHtxxXXMNVjmj/ml/LygIIlS7G
wDJwFeswquzOo685kLUwKIB1YzyNjopnjboeeArPJzbDWZm924lkuUC5amMpjQFs
6Bggi74rMag4HTeAeOyQxZT8QQHPAShP7gRV9TpYlUEmH4L5pPskZ0DjlnjnzZtb
h9MmJs1oC6UNUVC+I2LLTUhRWQdIEkxdqV1Owy8MMHuqZ44056FYWPHXrq6J89V7
x0piSdKkSpGxdiX3LgZv85UAR9iYeuCTV0ro/tgV7tsQC0GZ18mYPFw8ilwqWEQI
ITmxkGhhWLv9Xtajlwtf4AjfECPoWyYnXgtTJgqnZOJa13OcgFZws/DH0AtKqSlA
P5A29bpqO48XT8/mfLRUnk6grO934khPia9Xjpz1FJPWG6LkuSrhsyb2zH99o1a1
bHQ/NH1PIVIg5rXTyU3MZOlRoXXUSlbASBImlWW7hroFvzAhqTItAti3q5M3yO54
VCMuNcw7ZejU2xx3uqcIZMUtzEm6zwvP47ZNFMgxaKbxhp2IGGVF+7lFsn4eI/C9
70ejy1gm+WII6Kr5l1X2wJHD/dHmfptTKG4tAgCwfbvpNh3gRQ5lE3Y8d3RDdZqO
57uG8IhK3CqBK1wrLXbLUcx+9DoxtinE63PXUoT4XSnrOYYLq/ai8CzYkzRf+iDJ
3xGwbTxmrLXiqLmKLz2Tvyh0EXXU6GKrtI8wqUCE4sBTpiGIxQsmbvRtI54dcvzM
amdyNDk91yV4sC/iFBV2QqxcGxYJTcKePW7PhCjA1RUHc0mk4RJ5KXHke+gfv/VC
Ard2jaJPV0LXm5bKjubEEt6H4dIwrSeUdspg4jvb/iV20izsA2cZ/g5e9Rlc+aNc
`protect END_PROTECTED
