`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMULDljPehrMRG4e1AHG+qMP+9roOx2wpOcFVI7VhvOKyMfjO+WkpAKkov8xhojM
1XZzhAQ8nbBxJsTLtWcbmAniys7HpIUC47LlR78eh+DjoPy9Ruixkx6UKizoMjC2
e9FxyzXWzb1uppMemyPBvcODVqfkbtjdHkELuiapJEzpefVn8lbf1qi1/H1blOTW
tY44Uzg7P4bxHjo/5Kxga06dLUWZ73RUcDfm/BaRJP/+1cIgJWx5dWTO7QmdtP+d
ZW07P1ojQ0sTrfrgZuiscf2KdcK/lqPqQCUZ4MVBp0Rh+5N4t6QUai+Xf1I3FdOt
ttXB+9etPt40zEKAAb21LziYfEp5i/P3Bv9qNefq9NCd3cRGYRF4foyrXoWWDiMy
cdjD5fChPTGeBR2MTkV8/FsUo/l+pVzgoFy9vxBgJj4HzutMim8+M/mMDadDdwqm
qEdAZHoOYwcOetOsgyqB1+yfZA0F0pWPjlqEwgZN8jLam+c8CqexbOEmWVfFbjut
disFVTyWgJSVr6iLnk3PXeGvnUzenY8+6UhoDkiGd5f1Pz2iuIOXTfW+ycdvkdyi
K2/az8TeC8y9O9AK8ET67ExvMDABQUvffDviuBT5G6mdt2FtypRb7XoPEzlVHEA2
mEFpTyMwIlKxzihaLOKjU+0MgChnZEGZwclx1NOV0qrHUHR2hEDUhCI1goWrUJ6L
JJdQTt9/rn2TWDjNK/4xVl526Xqp2UYeCCBKI+67FS0i3FtiSVfy4qRoY5IOwW6X
cjw1U/JLX+9LHaeVaLzfh2VpLkMkKpZxb9esxz8bwCO9ifoMsGudlZNfqEsG8GX/
0mO6A9+QmTuMo8gcB27LJneu+9kZ4ZsWSWM0gBr/gweC5I+K+rk2TldEkCKXKNWT
nTjOPcJeVkOa/DLsMIOqZQ==
`protect END_PROTECTED
