`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c7hi0OKxASAHC0lW38C+bBI/zFvL1Vnp7AnGeAeaU55fAV2haeJIXCmYkiW+6UIQ
7WWmqBKS9qxbQBvbpnofnOOOfgGdQvx5ThtzowXhOJisasHpUBEK4EY5NImCJPhc
uOsBNxzJdt7wNPB7/Q5ktk98XTE+w4IR5Tj9P5RY0yOPaLCLz3nRyDR77ximnP1t
W9QA3v9T0aNO8ltWG6d2hvsYy+EyPd3NXTjh2SWltqDmFbvTIkAtt1Vlu3B+tokd
xM058kagJ3CSKrTvaDUXQTmFJD7YxNDHNrqkQEEnB7ivVayuzgdTZby7I3df4f8e
qU7/yH4Bp5KaLop3zSI/WtoU/LZehVUhoQV9ktbvcWqWFw0YasHCadARMddwlaYH
YdYrO/DNhw47mCXpRi/SACzI6N2uOueFsjSriRTRMf5zF4UE9Kg8ngUzpgT57R6l
9PQIyAMIWyvza4yS4HLdHIkPY9+e70hyARc7wZoQXDWzSa6c1DAJa/XbjFffhI7K
zdMPPG0u3nKj02BkP9rvrD+L763VA8BF60GKF41f1OZWbIiZY87rDmSgLPRr78l3
6dOScb1W8628+xyArIjjq6JviKYAFtLY2Eh3BYDuigFPR5GVRKre29HsSC3OVYyQ
CLp7kB+kIic+ebZxfONWJURSEmP64gCrmw7t8ncBeYYpvkoW7t1IW61/aLVN7i9G
Oq0HsSPFgCWnLfo9++0AkWD8qPs9VJaGtS+oQkZFa4jjm60JEFncyWApWEJUjtiu
6GtAaPkTM+BQg8OdNDMImrYsPGlHxKjWXNIdb1Fra+014FzJXwXcJ95mNNPoQJCy
DQAw+WJou9jRQLpmgtxwLfVSEdbeJd2gOhoOgYQPlS6x9kuvpAPiGEk1V6cgNOHs
MfIZRdpPKE7C9i94oQGD6175P1A+JkLc0TZ+tRap6Cyi7E52xdO41NX2/zgjbhHk
TMiQKhcJHElI3Q8ghiOtaOXUiC/VKC7t89z3m70lalVWJ77A2nX7ixIn0s4FEbvD
WDL9fxeYNjZIWR6o90TN525UCx7SAF5iEJYeTdbR2IifDkhaEnnKZ5d9HRzoB25a
5vSg9TKHlgIbSLQH9Y7U9yte//uNYXz6lT0ith2/QfP2NpYcHK64kzncGZ6pVibb
b1Y80gtEN5a9uXjBOBoEWfm2DOJ5VD4wzqbpY1iXceF9HruD7wlptRtTuNMPYlq5
`protect END_PROTECTED
