`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DRMeibZln1unoHQCXPfwJBQqhVjr/eakVrBaD20HiE4JxjGFEnkbftHAgDJdW3n
3jR0/pdOrKk89f6Vy5wYTgIm8+vte304bLr+eXqgVcYTWqqCzvGxdpp5kYSSX2vE
YVd79iOjVHhbjWcGmFoxHbTF6rvzXplk0ihGp+5t2EjDoJm+xKZZSCU7bPSCgJxf
WSH0E/PDz1bEcujRZOca0w+ZIrbtlgZO41T+vwMaAo8eEQYRK5sPRNTnOOurJAzD
p22cugdZcdb3ShuXZiAe1EDSHZFnE6HWb9H+qyI/oGvqPNb2KHqh5g+5tBAlBnCe
Kq0v25+SBx2ZUd62v2Dz/Tigpkf3Z57Szlg2j1igTADF6cu/5IYyiSFG0JlsSb91
EF/VRoAkyd9CdTI1OPTbmQ==
`protect END_PROTECTED
