`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LiEF6dTilfYPRIiM+bG7SlQurumu3lrZRuwkH2P2L3a+S9kymi2QfFF7k7SAaI0h
CNgJmDiOq6hOmxGDAnQML9jCmbH/vO4p0LlCAqTg6sjutWtUqbWiHZ3o5jU5m8TE
jMaM8VyypccGB71EsTXIKe7BecNgnIwKdadh5ODQVQso9vD/+bLNOpuDsyztBcxP
g26idvpL5Ov1RJ4I7grH1YPQWuOs5C7A+q3qGgNrZ5Q77s+aTqHRWKrGd0fxNyhj
gzgrYFx1Sdp2T09wKo378bxI/pyAVKMosWfHGQ6u6Wy/R3AJKP9TqwjlUQS7R+LO
+rqozyfRtPFxn6EGnAkV0EV7210arm5oitsFt/qTOEQw/IZFkIngRCbTsKYuRnhq
hKf08bmvQf7duVkhoy8s31VytxDSFb1cJ5J4YpzP9Wn3XYBEtPoRU27B3BFXeckz
Yu8Qq2WxvRYU7nGVc/jGYPJc/733SRra9wA1CADDVrJGtGGYsvOpFkyitxDqu9P3
AG0qGzcHk8ZzAAx7OMuLamhvr+0ZXjta3k71QnwQvqkD+jhlApwGoiBCByfmEQt4
oB4QizkB2TAF8ns7sLPjoqfnvHSwDjBdN520JM2D4Ma6LxS/qmEmSY//b93Aoe2M
8EHLRSgBaa6U9mGJwXATyEwVWeIYpim2/3gfXeB9P9Hh8ntTL1n8gM+/Le1boN0E
MosK1WbJEq3zqbUXmBw29cyD6azs+XkEBQHWZuwXM7Kguvks5gev67arrVFjlew6
IF3rtaI9dtTTsaTHZ4auhw==
`protect END_PROTECTED
