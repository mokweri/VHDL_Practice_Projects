`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zj34Pa4kQvXiQyvdZ5KwUSED3cp4OGiYF++15JtOyW/4eyBwFMHqhxDTuFH54Ikg
YPDi3WPiMFlafAuczXETM9bChEjIscfYRZ+bsnjaCncaLpFdOrzCZTiFFeukjPVK
HRHTdKUjF+3sV/RchX5aN/NArZ06wmvsN92F+/Eaum5rclFcXKc+opuJ9yEBKn5P
/x1qnmJeZ1KJoKxAkbAZhNNYv8acYB4rHh0dJLpliS8TXFs2wtKZYOWaPOZ+jwLY
zQGdFqacsTIFnlCXjcReUa8rnIm+gaM6K6QuP0gxOChhg/LDmmei/8FfNAgNHHss
GISx8VP0e0Bq9Addgw0CUEyiA5hgZMbzmFH7EMurXeJOZV1k78ef4s6sVSX/qodk
XsyfRdY83ycbDJx1S/WLJuV3VPBx0VlTGyBG66Eu7pY+ovj8l7WV9tTaLc/IOw8T
fAdF2vEzi4CnC/m4uM6nDId5Zz6U+nsTJdJKIbeFWf+oaY9ElY8Pi4m5lsIe6Gc6
ZpXcZDNgNQB3Qf/JUzviG42AvMMspxU3EprGjJLFff4GbSpVpUwQGrd6asbnmFOX
aG8eXOoJctXNrxQEAYCcE7KVbXCHWWC4//WxxdNAG6a9e7lw3p7iLl6Cl7ApAzDt
ySd8Qp85cArUAN3E3tG1/A==
`protect END_PROTECTED
