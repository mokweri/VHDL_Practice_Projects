`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2uHPdzOiQC2YHNufqG7WX/HRjc7zZuJDS3KZRcQxipB9g0WjkfxBuMCObmgH8BEv
xDEQbkanJZxxlzXEzTd1V4aUvj+ln2SvVlJY+M85PFqB2uEkDk02NRqoObK1V3sd
J+j9ocIlEsYB6ZkNYT1Xi1Yok4Txwqpa0DVI3ExYVi2HvHrt108rKn3rKR7iJBav
oh4t1KtXWGKcOyxwWIkaPQn6NCI0+zrOAqM0EO4kUeqquPX5WyxBZ8eNREOncGjq
txa00cb/W/2L5hnMpOWQy9eO5+6/isOD2xlhI9himWo8nTt0UgY8GTg1N6cdwwrA
SzG47TulzEUPb2PzSAg4iy48lehUuKSBewttaHgSFTEtmEP+aGIIvWDMegyFb61z
BKeNpSLTFtMpi4FRV0ExV6gK0hlPvSezoyy8lehIvk+xhYG2LdMIj1EVtgU/IG2c
h1D/No7GnElTFEOMUfSYQ3pvhwY7QGM2lg8EqvhhIoMqgiIDN7ctGYMoHXF3P639
o8MxeUdU86GRbtBFgVwqhQYurs9R8pi1gvsLXm+2EuXA+q7dLpznUhW0kVXLM0ui
POnzF5z/S26W9c5LyY/XlVZPt9ZIINph/NXpy9tfYey0+NtlsIsBth3N474n7tlz
9csfNduKbGiMG36GAG9aQ+F+pr3bQaJp6D6Dg2PZ4kRrMMJq1qOxIHIb+vXP1tGN
jsDINmCuZSY0unzvh9FZW0yia/cSVksjjAzMbV8m9+/j3oSaDliYNyyeoX3xIya6
4qr0SIPlF7FXTRchQIOMF7fsR18FLN7HCsENU9FujvbLWcLcxY7Fue67aJJZkJiG
lslqZIeUBxpNbTL09Kk8yMFAnt43kOit2Sj3jd/w8+LJmrCZvwInITfiHYbqfJO7
tiIqFgiFcR+6K39TDkRmmwttmMFc6WbHUIyFm5p19/dOx64qRraBzrh2WYTneKQB
FhC/6wgudMXQLwXS0zZcV++Vtz7jp91FAyRdu0bgi5/cmrtXcWLfxusjK2Gq+I92
mWcNITX5e9l3I0Mkh438PBBi0TSS2qsF5JcKhmGSQTY=
`protect END_PROTECTED
