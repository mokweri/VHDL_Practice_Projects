`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iK0U3ZJxkNa3Q77iIoYV3puyjcNLhN2OvC8O+CD+nHj+9jubXiXatPIVYqZuuM/9
cl3J3uSjp2kGauMW1sTKyaHXos+xmfoBFmFuAD1HKQNjqebWoqFYxEZOBiWdc/5f
Zjb3pJJw+eoyJXEl+vHR7LfXhhYF5Clztp7JEnxa+tK6FYIrLK934MhFx8A2hBxu
wbQf9AzUHYxk9aa/QC42ypr9MEYuXmYEnfCHna4RGINNQCS6xdQVWTxt0UzoLpvt
/r7ow4Yo39zh/Q3ElAGtX0PDPdVQVqhqQEOpakoJEaGDjJhUtRmHwoOlYgYruaxn
tedfcvv7lt7RtL1t++P42qJXrYmQr8Ec9YRhAz50kHCQzN86rTSjfZhO7pNajGmo
Zpa2FtDifAHE1EFMKA7N5n9o2/J5TywckI1PXTKSyCWLjjnrvBCfZx/NX8ghKLj/
pa7j5QuHKbjK9/7b8D/biPD0gSe1L3YsFRt1nxg4aYFGdf0p5eenM4KPMDWRZd09
h9nBlaCqA7D010gS48I38AMX45ils4D7yWwWOw67HasXLTGfzl8N7S8iUzFioDlo
P4aqadQ04lWOsAVaqpJ9bPNpT8s/1fjDT7ra7enKqFHg1ybxe8IsBihi/d8d3Hzo
lC7BvgJCTYHOigizk8eVt+9Isv7TmjU7kmXr8GE2xDY69GOpbYt6oDJOtzhz8qLq
w3BF6ZCUpFaP/4RFoUOdrzleGGYII88LUYNGL2YJbfmdusmtQcRccrmdMY7U6WrI
+aojhO6rbxCNHJXdaaEyWtwZD87bc2AhsNn863oFWHr/be55VT5ycG3nQkVNO47P
TIDIEzm1FlbStHbet+48nZTRkc8YjmCifmfeAq6m0hw=
`protect END_PROTECTED
