`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X4mLRv1HgqyKhXVDkeqmM5TfTkg+bqNf6EXTkTTIqVDhI1/a9s5KeXhC6ICm/UvD
MS2Kg/ce0eiUQiljRC4nQn8UqS6MsIIYtwtIUEuBrkmG3yskdzOVm62HCWZOpbIO
6+CTB2P0Qwi0nCCsaPptwR9+TWdg5otCNoENPG6/GncO+3/Lby1PZtB5nSJji2hg
jHdw0XXulVt7uHEU0OQWbHbdTYP0dPh7PD3NVaR9jHykNr/PGonIbhD+60AsUBRF
siWRDzh3kU/Yh269VpX99h8zsIki50Emj5ye7cQqgkY5nI+Sqf65kw3UBsfJ+HQl
fs0h1wYNsJEtXpFfH3fQj5uP/ZyIVvCG0fSNGwtYZ7/Qba4GNrCtJ456dDzSG006
VSNJymBRiIwXquNnSuoLSVtCR7VjXg/3rLK4Kmvk3t7EIxL85DwTLjSN2teG/Dta
ohiOhe9FNZlLpzBqYGJfgMn+US70Zvf5NOvXGe3nzQaPoW2vXehN+5LNU3eH9X94
EMrv/TH2SvYhTIUXqsb2UYmxDH+NwNpReajLlO6agrfCX6JZ+XcD19+TUZkp59m8
sQpnNtntZVM4f9JRalhO/NYp+mmbI5/y2xEsvvHZKRt9xjUfY4sVIlx344GW2DLO
PUmWzafqkC86vXFvatbU89KhFiee0BERrPrChmow5rv+MXfpZ2FLurdDTx5nYaiw
nM1xZY96YI9gzaaNqnE2ul/u2QVcwAIBXPXejUhEdPshG0fQDjICf135l2cdxVwu
TJSoq1vmImku64gJirXxgGSn5KWWXbQFGS4NDQzMRtMEfNv8W5OsD91NKpvn0W/L
n4PS2InKO63fsLP7dgWROH71cNS15oIt5a3Uphd9uJxddeDX0Ga2nsl8TW+7Lf5i
Cc+dq0MOp4X5omtmV4mYJ96Aa458TTXrQsmvmqEQYffeOZWLE7d8TNBDDBN9Uvzw
Ii3ml9aUkKcXy+w9WH6CyXNJ/JuGKA9Wluug86CUNBYzGLfvsFCLUWzhBhRwueWG
EXA8o0V6KIo/v2Q+XefK7r2I7zy1x1t6Wz1NghSsEl+NgxTSf1gZ5TFVZosO4v0E
DsKnJNVUdRY3vMD0z33XryKVmG2yk4HrFtTKvBteDIjKPcHqbPTTcnxYKYNcsW4I
RxPsH9Y7JwjCpjrM7GQ2wu6c06OI13+QBiIw7o4IsadTVEL5Wi6nzr7HRN1YDyrB
V0YynHk/o8eSyrNVc3/wb5CSDWcxSNp0h6UxAGpUCqOpPCcWBnDPANN/7NcLAcuW
0jwa5/eCC/Or6s3vvfuwu5q1DUPg8man/fw2NZgd9L1j4YlbNCX8Oh7fszeFAjo2
YQpsCuJxk7Dg80vdF0wdlmCsB3Ffi8JcyE80MwWkRUKHTKG1zLgUHCot95epQU/B
2oAdiNDxvTqgN0pQnx7tySEijlEoKI7inzl4Rw6jZg414GkDFOb+7fEr7haEKLHS
MH8Wd/QF7vTrJycYiduq9gFEBq/EOQVNV3rklIB4D8ZeWZbfrkEljvT1yX8ETPvh
Qw3gShV1QEv5NB/LzZfimIE62x0DkWhcLbi9rXQusvO1vgS8tB/Ihg+N4blpXSL4
IehFZ7KbYyJkItiuPIMwf8zkOavnKCpEwwWkJ1k2YXA=
`protect END_PROTECTED
