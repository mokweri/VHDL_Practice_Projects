`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ewb15z0Iwta6Q6Mzs1e+yvNx68eLGpRL4EXfE9MUpF4rPjEAGy4zR3nmlRPtyTi
KhyTFKczC55hL3+LwG2fMbbJ4RJ+RPIJJHrJ7uuNgLy2f9tHnhm+HOV5oHCPvsW0
SFuqEAmNrn8j3U/aQPkhCWJ8Hu3Z2pfSaolipyFP34JTWcrYq+ZqAJ+XoVQqSrx2
5qHsDvJDdekG0rCqmd4948p0ErJMKG41Ehi2owxWmwqi2CDvzKcGSH6cYAGR7R+i
G6w5DSv+DP0lV7P61He0uNcoO/mjTJSxXinwKTExC2TFH367afNBKcoOrVUk5oqF
MDLQsZwYVagms+cVivO92+k8Kb7tw/HtCoHg8MlzuCRS1Q41L3P3M2I43jypi/8D
I4VCdvoJrRSvuDCSmFxkrJOqBCwCntL4WKBIE28YZfdTXKjMpUhPua5Nvs6KMYPL
GI0cUB56XU0lyfrwUM6KbN5HivpUWkpmp93h8PY5rN1omL2fBNhzKyxfqGRDD81Q
dO80lg5mo4b9FVLQN8v2nBP8sCz8BFH84FYqUSxalF+W500FKFz6dD8ql0+18NaZ
fuO2x601cK8JGnuRWAXPuFrzf+ceAC9zZLCzrHPFUdbiTyNLkk5Qqop/JJ6hW+je
QjnC4Ako2w9zYacqhHBJ5NCLBc10NEbbE3fAGz2tSz3K0/6RBfRu9bkc1LM0bxhF
UDt5EAVVy+L2Pbgx4cGja2MtAsrff2Y4E03M13YyxDUZyxcr7D2L/Z3AnGPWd4E4
JDwTNj1USChM3IMgmHUfI7YXIL6VsWVeKUCR2e2HiSKZcsmcR4hZVgsSoSE9/EWr
6C9miFAZhXm1TUJ/9851UBCwF4KHGTLTam1Z1PfAcbXuPYIEIXFZKNZsXtCq6cza
QlV9aMP6xR2+DFojj8oFrsoa5/1qynglWh2JXyOTueDiMHlSwwycL5PIz+WC/r7P
`protect END_PROTECTED
