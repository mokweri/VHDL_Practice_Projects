`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lvjKLXkC3MS9/GqnxdWy5fh3qePCrHwt6kZOBmKfamMypgY/V+wxb0Ap7T78Oe0t
n7g7QYsDFjnDWxDIJ5+uYVRhH39A7Dkmi5z9+izjP9ukYTgghRaXyfMqm7229EYa
qjITcUi/fwIRwUqVDz7DQhsO+9J7IY4JqruyIitDZpe1yPPWUR2RFaY5s9KTNHbs
i4i1ysY2LPYqBlU/90pdFfjIhghTh09Hh8mNJiGuT7Ai1Cb/0NzCLT1UzvBK9Lhe
uh06nZgY65NtRRgqcKW5Mgq4XObrhowzEBbad2omrIe5p14SYf56bWdQl0bsWXfQ
5hLfBXzaLWyu4pmsaMn271G7QTHn3abPssEAq2GXh8XMFusEeWP5a/2t2FJCdTDs
ZZv7DoPx272ayAbus0ixqJJnJfAjY95nrMwesE9C1l/IzJcaZx5IRRkHlaxVskqN
JyMH9xFciCdKUqc3sOdJAhwoGlWm62ykViRQ046jLwJlz+U20ge4De5nGU8fImNX
0QSq5VpB6i2KqWbnYOUZC7Qm51eWhsAr6IKgxzoNEg0iP7jQkBhKuDtyBP8p/mQH
egWgJyDl2yLujX/DFvPJgnT2UU8/TiCMbaFS25zecjggI+OiZzo9XUtk/SQFkDHt
WaSPtV9be5i2qcrb/XdhgjKWViBT9kl/eDAG6viOhkYicOfBJOckw4u9OdiQVypR
yk2RhAB6a85tpztUPef5zouF1Rg9da8u/LQsCNSgcAmSltUdinCLlIbsmkDlqhNi
2CUujh8axfkrCto6tpiQan6NiZNl2pzTl8fJVjRA4eyPfVa+KZCaWKrb6m1JCc5Q
ihci8DoRv2x/FZfrL95fDUGSd46I8Fbhs0g66VtJA7dIZMY0M+F4+3HnRbbJ+p4G
v5RNzh+9LkYAbfv1uG75Bc2jUfxgIPFkEAmb+5RR0ZE=
`protect END_PROTECTED
