`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wzfrp/r45wCmLGzdXjH3GKNInsAnccIPSQVTQWOthoJZ0RUUl8QegNW8f++KSIVI
1BfZz2QK0cytzo7RQjbQzK/Rf8+zJlb0rJRekBxPQRDdOsTWA4LZ/exV0JWo48tk
Xja8i3Iq8ARB0e2RPdo+ZeTMF9qK71zLWoUk0huPkrYtJzfYUlWkDQFmzG8v/0EH
2R1vOfKkKBuWwEN5SaEJj1qkqIA4/ONIJq+j3D4QxpYcq30ZJdpqht5yqDnUtxNZ
X4a5xVHtc0mulpP6wP5WQh2KMOG02MB1A9rbA0aPK+1GWbCgUgRh+oout32YCCwe
0fGTwHX3pdM6pBioK9+sytHXq7cLCnM/Yln/f+Zii1U+6yc/uZzzmUeTunT6dZml
337ddkLpzPv9Rvl6/4TpiLlWZHz3gy9o3xQ9hIouhUZadRkXr4FqCuV5lyD2YfqK
JcCoCZgUOsJ5bFMjCREPWugYWYmEtj0jnEOXN53nmiir5aaBaNU2ny/T5/FT0Uhc
bvV4dC/r54Q00DI/+paJoI0ZMvHIKKo4xWK38x6Zovn+xZpxlOdlhf5a+z3UkMdV
WspCsjWkAI5WPX8afZ3LA/WNWstFU/IOlhZnWXh4zuBmEXli8vzi+cXTyGApSvak
p//KriodISOvqkqGEXj4qPA0UPUbjgey6X4bKB3vSpLEdVxkJL3rI8ihrrSvSP96
Et24+4XtA5wkWCv9T7vTaVY/V7KPVDTVURBetCvDE59RvG4BPssev6XsuzeeBxDd
QYp1/0nI/drkT/g1p1IJdulQo5k6UHryjp7dnV7ljs5Pzsk/a+CLzBA0CNQbESKm
Dk8yBrfOaqfuLNEO9kkkCXHoBPmsvDiK5dmJEfLDF5YUqzvW+OA46LgrAuQnC/pk
gPqcShB6JN+FRR6hU3bHLL/nfmVDAGk/b6/HyBJZJMSqE/y0g8jZsBq/K0QFi4x5
kRxQfO3nS26J9eB3zHNkx+334T4y9h6z7Uinyv1llTUek5ys0ROfSgHfZcx6HPp3
R0HXQVwE507gT5Wvg6pT69uJmuKYiYH1Y1pDg2RUi+pdTjcs0o1XdppocHTby579
NcwNTOHTJKQL/ndPq6lSIfN/4JHx9AbrpCpioQFQBN1emLAlbb23qJO7p7bJAuIc
jlOwAxL+gc9IwGIGnh465fzVeV4UT3bgldShD7jbZan0RLAfFfyCvzM4T4Pth5/c
CExV2/FfvbZ7F6wFgMIHaSkAbLDwhyiKcflndSeKCxt7+hKKLfyGR9W7zLJFLcAT
oEv5P3kFWMOPBCRKZEaUNGsiISOtf5h/doCD2B+7Badc7EHghxA1sdSB+MidO1VP
RZ6xa1p0ReOILjzNTe1c+peu1iLJfizOGKTzkLiJ3f3AOJHCdjKMp46wjAtkIg6T
LRkt0CrZIGJ0MyIix/jpBxPMfSi8tDq4kWXXv4QPO1RkVDZ8fAVNfI4RwJTErIel
RUwbrM/NziqrtbtJKbgI0BAxaHpk2SECSBDqQpPmZuGaAzbRKy4r2K5oY/c16AGt
RE7zzx7kgaB8F4OEDR39LY/1mJYgQmhbswcMDbWVAew=
`protect END_PROTECTED
