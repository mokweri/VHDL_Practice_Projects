`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cf5oYU7U4o5RJ3W1IErlOk9XTIBTNQhW8w65jOUwFwubL15oQKzjGhEqOFO6Qgw+
U5FiVFtLOTTMgt+pJ6b+2MK6rJs7kRkB6MlVl6rMw97gCFgwx5ZrtvREimng8q8q
1AfY+wiDhiYBjyJZpDLsp4k5xNf3NWpPFGdv7IsDUESC20Xa+NOklETffXLG3d7p
oHrTUmOkEls8BAhB3RXc2c6n/WIjcdJKvzwPAB7BvqUG96QNiPMTcEwX4CZ0fljm
IUGu6AyZ9mj4WLQJOu8cFSUWKHp9YzIr+hfvZz2piyWRloLSbs8HjXWBAYOfi+XB
xvy8WuK5ohFNkEDe61OelafwjL5zsfYI7SNXTc6/9j16aCduOFJ+C77CYXzxVy7D
aSqa46XYhXjPKIeTTe3zxRLxhHnjiHYLuqkt+tNWjPLJSEVNQroIjlk7NHdRPE+X
LVbLI/4GlniHXiXTofgQ8ZMoxuHv7Ahbcsx9WlSTBOP6hBmspVZZUW+xFOrQQ/lr
6H/hrCphldceEkb+dEUI4oP4Keqoa9LMS7aB/3CzsGLn3xjZyvTOmntZGZWEgk2s
Lll/tvFPN+6UX8hV4Jfs/g==
`protect END_PROTECTED
