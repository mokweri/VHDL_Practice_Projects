`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oi9GatZiWOi/Wg+Am81GH0A8+12/qVcJaZw9W+OnYzROlEiWXf11q6jXVnTtuMPL
RzcrYKDkdaHCW7p6Ur2U4dcOf6U/JqHx9VD+ZBEMqfTulzXmehFW+kZPu1vQvdK8
C2AkoxVrOS43HlSNqiTUCCgLj6Q8HjK37P/7nE59d8bjIlI0HTg0sI2XxIwEpsEb
7p6lnXqC9Rw/GJR87vqimvw77ynbcZaFQUb3Kyd2h/3PU5FHi77hsPzVmRDzlBkv
Tvy0h5NYc6wgCwjhVdI7guC6M13fMvO5YRyuxh9Neh4bZJtRaCKxwpAIngvo3OPX
c89r+RBrztcabhVaCSyxWcQ3pMRimpd4IqOlZh2i310ypvYexUVUIzivjlK7m//9
mGfyRuxvcz/2nISGpOUQSJlCn4Cj9mEzz6ASpA0G+GvwxZjAc2/A8LLXpXhl1TVW
yc+O0M/0GnkEcMWasZY56tIUTn9zEFZLVyRctudH55eLPp/UawpofZvmEoKvcG6j
c5hzeYsPnFYX7VSQxq0RnQlfz4IoTMEdAzCufojz6Z5A+PynNFXmwb0xO6RDNrlc
0IxD7b0c3bnHzcZWzc1bQQFNSny/OI1ZNQxprZvXgpfd3ss61F9f8mHKJopL/vOw
RNMzsH1fKfLZGZ6GvePtxC6bUrN2snqE05/fjRVzBqk6XtD3kBPQYLxSZZ2eyaj3
jQlDuQFJNlL/QHBJHAk/0Nm3MCvbWY3QFfQ4/uaGdKASstQn/sHt4LRYLn10tkHQ
uk14oij6N6/e0NgS1TZinbhEI24YJfa9KLzAsLyGh+MnGlF5JPDaiSVrT3cc6MH5
1YCNMsspOsYA0n4aEI7NTwfULFjnrrZ5ypn+kL2uNoZHsb9Xmbf0P2cBsJ7e6yye
J+gNWwaAIAQgCDWp+y8hPhrbMiMdy86WYFhzIgqn/9Q=
`protect END_PROTECTED
