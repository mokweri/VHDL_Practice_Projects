`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aitDbSeK8oN56d4S1bUmLKf8XTT97FzxWeX7p7zh1UhQsWkDdj4aQ0Oxp/iXsOKO
vX94o9r6Tw78T7DDLZWc4EEzmhH3Rkg344dHoCsNQZGrvcUbbs/Dvpu88VXB7h8X
iu9XBBCuh1Zox9ywBJJFSf1BQqf3Sgadf05/wBjfFZhnYG1Hn+xDsQZUlPfQA4FL
4pTLdLuZ6h4l3iyDJGh/b46tAM4uqHyAhrLSTTaya4Sm2XhiQEcHPVAucjNXDptq
3nENuIUSM4Nl50Zdoa1OemwcEmbaOXJlT4FSaJD8iO9Ph2IcD1ScM3QxlF4hCY4U
pV54FSGjUYlI6GCbMjFsB5ZNJb2rE+J9NvqfPCdCootAJIq2cD5jA7mjFSQnB09J
NOcoWA0h4bi3c7l8YkJcN5aT1R0iko9BiMw1mUM7241IYI3bu+Fg7huSwsaVtHb2
ghbt6UiavAD8vCSBc9h1+KC+K6NUTLPLL/9JGL98gl2zKZS3ABE/cTpv/nRSCip7
mKcAPlTWsZXMIgD5A0n/L3qjH/DVOUqyVsmGnPwkQzg=
`protect END_PROTECTED
