`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCwSwWxukx6V6NqCwHoh9VlURwxe0QG11fZ98etaYwux0f1+8kYT7Y2/FPpKGpkc
sBjdyL+aDWxsRiNekk8CmTy+DUKp5dlcMrebY6c6m0/nN6PYptman4rndZg6P8+5
FnaJzosrkVCCTtRqyRr3bWcJU2V0HkfhTIY9NLDh521Ez14h8G9QIkPn1eb0axNE
kVWBlNJ/95Lzx6+0BwuII6HTe/2jOye8t/mEfcMAu7I7Yk0CvZ85CIV3euY34ZdK
ng42ZJ0t6eIebgSR1udJ0LMLYUXXirk4NKAdToaazeTdzPYkZLiDgrQHWnnGWpva
K2noG9ygjgQCQeFo/p2yfWOIDD7jni4g5m01rUszN7vt78nZpQgKX/E92cXMB9yP
cgMVKdhgRVJfXjy13rBjP5O9gqsF+zbOhChFUMQeIgypgCdcSYsWwjA6Ie0ComY9
WNCqzHLHArQ5ku+tcwlsgtCHWE15LJeYOfrtJ2mB9Nd/HYpcRurdAMKt8kc8G6Jb
owIAIIv+3mkSpawgA9yHfueF1ygChCd4aAlyZO7MR8Zv04QzLRaP5PZircsuZXS6
yetesNdkD1BEw/60Hd4kVyrAEZUVf+qpQevSHWia2NkeB1PPX96mtXMpNjz43K+k
jAxbLyEyh2vIm9NwpdDkug==
`protect END_PROTECTED
