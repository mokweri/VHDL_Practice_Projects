`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbo/3Y2E2W7pcG5sOm2o15XCx9ZEHd7dirPXcrDWXatvQ6TSzoRm1qz+BnztK+/X
uYFevuXE3HOH3LuhaNPng2qEVgm58iPT9WvqQ0IMWGMvSH9BapnnDUQsN5WQB5lr
FFbyP8vEtdKLBCERrpd+KaOGTlNwyz4/opQ5beMae+XMNzMTh1pRM9+7eekhkN97
+iFwmCyQ8oJjRokwfufiAETKsHleM9r4MxQVeo6bz5KTQinRGVhTF8/VVJBsXFwB
Nd7AadeMRtxjRKre9n4W3qVq+WjeKEbgT+tIi5u16VbdWnG3XTSVAgV5vG++RLpU
SbD8kIRCQEIIEqr0b38hIpRcFcTcYzzrRLSR9Dbpg9hPdU7ehgG97qKAwck+QjFK
XKZXuV+oIvDOWLQzuAmAYGg7sIp57GlhtOAPgR5Y7q+xMlcwLjvOHJ13EKv2gWcE
waymt44kdUKNBIz4qUlcSJuQJDgx2fYkymVsIJVWPf6TyR4Y7I7K2kFXScS7nfUv
9wa1yi71PCDLCfSjlzCxnqE2dQQhLcB3Dr5BJ8RIaQgcOFMYPvHTn2bRr7C3fKnU
bCBmr7RCMLyC8WQglwI5GLdwamefExLqT0pbf5IziIaU6SVeCsEdb003UvMUsT1D
4dmp78PM7Ybf4xc5eYmy+/8SyrUpXdgS+SuLkuyNlHtPrZvJHJu9cbR99mhgRd0d
Jf/i83Mpka1/7Bi2ishJlnbwXZQ2IQZnmkPsY7R4yXecKDMqPKcfk0veA8P86md/
3+zUhaqa/3kqNs7BubdPtU71lm82il3Ibelj8B2rKrWyBcfKaH/cmYDmreDlU4u9
PKifNnD+BzALl/ZKBaxkUBGB5Vz6TI/1KIdDWJKmI0doQQpj1IxUPLk1lYOTjEwi
4zif2/QcqpWM/FbaItINUCkYBLTYh0JJwYRH3BitUwNx3NuhSfUKt4ni3J6Zo3i2
HDeshxO09YIyDfRMgUK/mbkzJaSiPSeOii+BEU8xhtAIt5TW4j81vnwkeMH1M2+m
1AU+/PgZp7+QPvGdQcgTw5bvLrrHxUSEMaVVBZSZCHobxzA/AhpYjaYKcX/bS5ZK
UJ7vVzkytKrBCurc2S9XDGRoXNbLDuKFBgWZJrQhM/fNoX3WmMvj9uQJXXtpK6GS
MEk1Ac2C50WgeEoL9LtJCg==
`protect END_PROTECTED
