`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FBGykTEHBBS+PIeszHzFyrYTbQ+AXL5mHMbHSsEwEkMXtPGgO8wNTARbdspFz8+i
cpWueHccw0MUG3CACuUbWqPGVGfpLPjvUMDxLc41v1gSLFqAITx5F1UpUuRUJ5qv
UzYCc3kd2ZCgIsGtTnYUR95+XtKvZjbH4CXl0tJQPtA2joa2AYaMa/WWn8kJTBYA
GWkxqazOSPvxzC5nC8oqrbxvxwI+IzDDjYZdLNt+0X1PmqVJplIhLT/GMwhUrVOg
wiE2PTnSQTiRYNvmlxpIIv9JPGdQnhQW5M6NmLQau7jP06gJG0oN41w0RMaQ/U4q
di4FkfgffosVCZ//vdXIN1W0sdZAWTp6Zy2sLnBEClOWyRcPbXsZEU0o/fLtOg5W
rOQoaoIDx9IRsRO/HvFHwH2DoGrsPSvtKR+YJOKnUVuXgYLHYO9s+NUYGqw0kn6b
XvTlL4ANHjP4PnrDLCyZ8tA4ivm4Ajvia/JkPpY6ytJsRWarhF4dzH3dDKToKZHW
U/3WURreEgMJEzuJGe/ORGMw0Z3Qk/O0HAVadCQ0YBoCH1MFcNrzpNeo2WYnG1kc
IPY+lgcxpDu+40lS3e2EyqfZNtJciUbGn/t3Cfo1XLr0SPfYjC5N+DEZdtU2ieeP
Rw9m6Qz4FmwZ9xyToknHC3oxlTQVk198mTDA+Ss9TeuNlOqB9yguqZKHFdToR3fB
sk4u8poLiN/rvfRJ1VReoctkSsSy5IpnarRjUai0WlwNg7FlyiU63e+O9bD2JLGZ
bpXAXmw24avKHkOZcEigg8uPvNuCYHG/Y5vedYG/q3hAF6nzZ5yG/2rNM3nWFtt8
P3xYompyP1+KiHIDHBGQubvdvHvoUCktSU/oPvzPkar8gvndKS766TqmEUqPkGc4
0wKZ81sf9Zx8NI92It45mBh7LSxVur3xi7h6Lpdu9dF6KuopB1FaJw5Tu+XWy7yt
ZTK52dZvyS6vcvciACLxVEgviexVSMTOH1tHchpH1tdQJ4yxGxSjAU7ofhHBRakT
k+Rdj3dsNTsaTg0wx567OXtLGuGtC0asRej453dKC8BO4q8dfpXOUP4caHw+VWJO
KbrqLkuItR0dAN3v2dHT/ahneUZD5SdFInRGT5F97TSn10Dh89Exy4VJGB569pCk
bypNpNIKtBsJekXWMkWKnkqPZLlxBpSixbl8Pif+YMZrTyMjeQzRFqFAebbexrNz
Zu6rSoFB8LTtS64NRgbV9I0pCSN7s1yZockQklyAfC+9atnNyA8PmDzHuksnviAL
ywKl+Zd+gpFJw3LxO3k7LxMQME0sePKY41eYr38wPG6GDGZiYwtG+f/h2ad0k8zl
AyXu521IEeGfUyku/waBN2yctLPZlKvP/YBNeH7JiaQwotgBlWTFmfqBvWi8BeF6
1vMYavidlRP//rwjFvePAVzXB/xlOYOO12SkOFVAM/zohTD0HJ/NH3xYFbjSm/rw
st7x3wVNVRKcKYEkHRq6vh++9Nt+zW6TyWA4c+EPv2l3Zj8QqE0xXKDdzjE/1Wt9
B7cRQj/a5fIN8xieSO1Dgwtr7SUbMBmY35pdi/Rw/hMI9C2SyM7GxWYWUiPKKTg8
mFK6Psm99NRvwjaSt999PvoBq3nmnHFHdKQceOJGVPPZFgoSd5cu+MCniHlpqz0I
ukTkXpSSebZMqPoC88rLnxSYsZxwr9uknLL19jGjJncYp0t7VGlbNQyGQewmNn1w
f932ks81Xl4BQxhxwCyJUBY41ptGwesZ5C7OWzEHFc8gUR+zG6G1UBCconwNCZwM
L1ryJj16ZK4rxJqZyWao8lckjwOFT/AKJJWxBx8tdePluw04cSJHCs+5YGe92sZq
Z61C82NNQLFj11Y7uv6ZN6813caMK0nYZJHU4nwuOR/5aYfkI1i9cyNgdAR9yqRr
sR40bS3UL68FE0ZOU+wuj4pf0BgFJzIxtK+UqUnAigVO5seN9ekWkAluSX6BFA2C
FC886D6kLljOyk/2mVSmo4H9ArJpdnh73XjTdGQgDV8vJipGj62zf0K0azNQrsva
hkYEax9fxSNFyVLtjt033FMIICFmF6sqTBcAODs3z1iWblxw8kpiSj74PUfWurr5
VoClLsUGXccKDDEtL0eC1nSQbl8uU6qVGI6mH6QZ44bg7dT9FG1fsU3UJ4Ajz0wM
BNCv9LSdi85lf94oUkIsv3Ryni5xKi5Oox16nwoEgG7c+uG89EicktMwJGbZPUOT
XL+sVMEHMLRjDN8TInj7OiV2dT1rdk+Zm0HVvWVicUncO04/hyiGmvZxDhz9ONqY
uRzUeCja2n4mtbWvYu8AVzby48wV0hWBE7Jg/aS1ab9y1UalWcnj7ikcPjhjVsxP
xUCrG+yqF3A1KlNI9BAtxpM2mfFz4TSfxegHGA+KVCyG2UdJZbnJllhWDe29+oJ9
BxNZSxUAurKWdiPzm6NecC3Nbd4BDNemFMe7kSv4hUf/G9MeOHy1733Nl7cZ67c3
ooO4YVs9NBru9qdcBkQria9Q2vexSRnKr3ij23ySLXWEDnnC6q0HTRhrMdRJQfKF
dn+RXPzctaYNc22S4RCm18PKNYEhz9QbeV9TJPBVQifoN1JQucasBO1FJtAqiJ6+
R8EdoZyiKUvKQ4b2Z1dKitUbnPMD9KbXRdASPW6q3fgrbIkpfugNMWw0YshWTCwh
UTiHrAc4f+jwjzKQw5qewVibZzH6YasSlFmoLUckN9xNEPIYqUyxE0yqNfoI4Quo
BNWRyjNg7ViuS3iHqszZIogPg0U/AOMk2rELqzwSxyXu6YviGW0/3wg5gXDtd2gR
uTGo0I2LXPTA9o7jdeJC+6d8jqNM888wgQmAXBkpx18WoDktp045VNAe5Eh7E7i3
Cr7HPgajHaX4FVeAYedjDKCcelX9PRKDstyCWQd3ZRNoxiXEy2hYkqHCY/mgkbx+
1vbgxiCcayYSEmX19gL2Zalli+G/1lhmXDmMjFMJxh+SK4jEv2FDmBWNj3aY/dmC
nJAyugNbDu03dLQEaYvsunbWcw92J+6EcPmT0odjOyiv/v1Xh2nlFmDfZzdnPncK
aI4/euit/+g3NtnYrPxHd/yGg9wHhQ2+PFFQ4XLVZaM/Qsn81ifVqSRj0OcDsiE1
y6+vTFa+9MRu2YMBFSDvMtxU6TaI8984R9uV4nwlTCmdE50tquEBAFaswtgaSLND
yb6S6yG2HuSiwQWxcz/EgxGITUYibCWSkxWnkBlCMME/HYseDyy92n2BftOshNdu
pnlb89tSymApwQ9AUpfayRxzsEoqYgO52LOr1b797CFe4CfbHzA07U5kogY06qzm
GTDRnw5q/7YXF6Bfw4m47OuRnJ9Gp6zpFm7VcLYmYgaU2R0PmAxCPf0buUs/XRwI
6aSPVkZST6ijz3uepCaTcWfmxewbpUF1el8pHwx1rFyZtV4SK3UiD2mJAJAeUlcm
uQMcnJsOVeqQWejsOm6ox8dOEvt1LQa8oO7A+63Ddak=
`protect END_PROTECTED
