`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXP4G6gI0C1ySnLuTh9a2+ZXDSXN/adh/C5Ph5Pv5ZvMLN9Pb/sf7y7QHet7rcVt
jlIKBdVShKlnOtsBRd8r5p5J8mcOVCMqJd5pnhUUCJZp14rB5bc6vfGWy85gbVIM
Hf+d70ny8MTgro0g+sdtuSzEF8pBlVOyr7MLyCbPcWNOU3k0lKSxZhFZjyMu/Se1
`protect END_PROTECTED
