`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wp8gscGusxfHBu714Cxrp4AZ07w/rANg2+eg19G1Tw21gpK1LKo1skWb04rNNd9c
xkjv078vJQQyz00HI7uAO2qikaIh+twZIvu2CVKHJXlbegzbtc4tsq+MxSx1EY5g
7LpbMLfGJprj4bMdziw9Q7j0D8dx2ycXKhPis3rlddYJaHSlR02Tt3f9hA2xB2qU
hSTaGsvofVzsQIpqK2E6ET2xJ6MTyEe4AAIyUONp+MV/Ocq1xl0kino5v2Bjz+5r
RrJxEYIq/4lEGFCeHbJSNPp7IuK5O/NHahydlS74Q5hDQeL+WBMTp0F9J03WdIUm
HWwSMJznovAiYzMqJQxPDln+QknYt9sd5W8ecNNw5UPKUSwb6QmuHUaihNshvZ1y
Wf4Akwc8ZN8vAj6YLuejfTpv9MEbs6PWb8wwuOzHxL8ASFc5FNYeFCKLFPhIctst
3vSO2Pm0OX21usyzFPsUod1Q96nMJACM8YGp5ZQPuG/1/ppXHG6nkR53z4NYhvbp
Tmg/TipGytI/NXUZ3SfLKeNMTPWl88AyV5U/lx7EcyypMM8x/pu+RCBPlcf0rwe1
D/x4PJR+FHA8LRq2WgTw+jTRm1+PbZR5YTlJB0fFq9e+aaIXvUGJsPPT38VAp4p5
3O7CpuIGn5sakDt2ly6O79Om0Z5Gp3C/gF9CKb8nubW06/QLMiVTtxphp+iklzxy
W7684H32DNkVj4pQEsGDwLv59CkaFe96KxJ0E29ujOTwxI1cX47/TK58n5NnKjD5
DQ6gfjjFMLpFH7J5EBqBtrRoVtTrqmpsFgTD/+A7YMstscPfiaINQ6ZhP+2iUAeA
JOJ4lDz6uKTdRDXZDL1Ffm78guEd/7Wt3Ksgeo+si8zQ4Y1zTLnmP+G4dzGTWvOS
Ge2pV7tKlg0I7bDTBa9NGOK84zuydFliQ5HDl8LNDi5wwBrKqUu26vJJ6O9ey6v3
Din1X7ByLN71EMIbmLnaS8buHYjUjiUzNmBLtfLX+DIUyfi+xbYQc7l/HFeZzMCZ
ESOj6DsVqXCSXm6c0X3dhlUvsRCG7/3O4lzhz0qybY+h6mCZm6isApQXvgLQLHRt
h/dftNFw1FkfBlC5+l2fW0rq/vuoH6g+yikl+mYFPhKAU0A00MBenH1sQ/swuXNE
rK00jmgATqlo4bIwmzFqv5eGcRfMs7vhRDlPijjG8aL54ghdAzJQM5SbusWppo7g
SZ5yg7uf0iEe5qC0YDdpicKNlHcDku8aN75hY+aNnMar7LLvaUiWCm26k0YNcihI
vwWmW3ghnbfuIaTnXjulTY+brTGFbzEB0BJbdJV1WMPEkN7gSAVzunS36e/NXOwx
LctX42REC832OiuYWaHa0blm4uC7dLNGjFNYAlDO5cVmEN/ATr51wl0hAgoOlkd0
M0clG8CLUcheusK56yCIufYONCzFNE66mvE9amRr2PHT4TJ/z5yP6IXALSG4skuo
6NDy8qAEy0stcf+GETMnnn1MNCujPa6HSF+TK/bG3GgOIDvEi6y415Regutarrzd
SYNgvaRnajDxj+tQJ2vDZ0Di5/kjL0y2wtZMlsjbKxxBrNO+/AKoz1PZgvSvki8Z
ysOhVjLqunhBu2U8gkCIY9p6Yk2R/9OOMOi0jKH9vPmZUbraFp7dAbqrBVwY0jkx
JsQjBmasIGa2Ko6JGgZeFxH5Bf/er0UBQ9i2FJEez8cnYx7LJvFm3B5iggdsFW0G
HNXUM+mOH9I5DtjOFtfQlhQB6hVWP98akQvQS+tmsu2zBBxaP1vCeoH+bGkbvo8B
CVmyW6x36Lib5nUE/p37UCds+5tIhrbF9qr8pg1PGUFr4t64+kDvbAh6zRLxgzaD
UI3rDkQAoUFJOWFjLTTbLjt9tOIP0l7/HQg53VGTuFjFNttDj/hZa5SkZ5Xch4jG
gyd6mgz3o4vjgYmhZEsEG7MlTxuYRfQR+wQEAJPe3rHcYA6SU9x8QJDdPMZI+Z1l
T/LchBtmZpcJex2cLiUzvF/fl3l4F7BWML3H0jtI7Vc4JGZL1A6sl5kmKdN5chWs
QeZGi+WQ0mir4w3VYLTAv81V+M4XVXm56h4J8MXOQ76kPUxnfpGO1iQo7b4ukD7d
ThVOQp3tQ8XqX1gmkfITKvIvq6ZsmGLHNg7Q8i92qRXmWYXB0bJlp2fc+k6nd//n
UGLBotkllAif6Iy69x3NAJgdunvsvGBkVb6k6/M3dxNbx4NsPE0lR7ZswFUdc+So
CxTuuZNxN0nwJ1x86bJ7jv56b4Ka2GE/IZI3IBULiDOfB64zwvXFDBY4hQK0c32Q
jIYUZ4ojEQS5LFLTbuLY/RwHDLizCOcxbWrdzsiuMb2iyiA7BBxdg7YvbCL60bWk
DW7yiv09BErb8ktd6nWF4NyDXAtukbiVg8arxcw6IQzfbzPe1j77tjgeD9J4bl1r
o2szz8ztL4aKdRSmcZBgBPwC1LqFibODFLCitmTz9GM0tKUg8flghzOtZwaYaINi
RdqJmev7CAg5e5fWW4/t97/Tlt7lvVxZuMD/uGPnFXZ1uubxpOfQPdehWWmf4cFQ
CqOnI5K5jsQEFSsXES+xZxhpXSH8MYCXN2s+ljsNrhU2LlpeCeHNZ+Uqqz8EpqKa
K59WkiCWFN0OuCgaU4om089Cdj1sEbE4SLYoK/T/PC2nyfHhaR+ZqQ+mrSKGlUwb
eb35e3mN0PvFlddBj0f//NL3GxT4SjYHqzioH82CXJBVK8Cm8Lx90jR/pxGvXp2l
OypQpGbXpqrpMJx6S1M9wYuxS/6/AWBPN83xf/Yvgmn6UAGJfdtcNoB1XLXPxQG+
JtSxbAqSgOZrYP8jPvi6xML86vy1e7uv9FEVdosomq+VWMGSgEUA4WLiAXxo2xUX
cUKVOZNSk0eIIsK5aFWc1bAkbAOEpbPT1FGxyDzayIRP7ySKcmuUcVvWrVkz+bN5
sMTHu2qJKxSVbxt1Z5w2ieoqrA70phvKdnAOrIS/x2J+i0sO8nbpaTVuogPE9IGQ
AiAyw9HZgaclysYSOf6FY2UWdrtcVbL8jZVRdv8rQKiamiYLy227eOCOyEG/xN5Z
n1uoeCafM4WbS6SD0vTyUazEibRzZzcdhpYfz1LqJeJtOYFLNYa1NBaWrJot3FN+
m3BDHR9V4uurxOLmvsx1u6Facwn0F8UpavPHqPQXsC5TFlnXRMBjbUPMIx/ATzV1
7FsrdQs9w7cQleBdPuBsEpndhncBH+RsqQTRFBuEmzOrwOez7zaSDJ3hvU1DmBaY
d25Ufl6bAb1pEviejD3xBJHeTqeQtxI9f2Fj632nuwrzSdMh9mXIu81ob8GpVqh5
FkZ2t4+3BY72dEe1ApQ5KrcBi5bhqZZlJubAZXAzYOu+ydZP3ZUiJsKW/9gk4XTZ
+P61hqzwLILJ/Z+HQ8yWcJhCq/OzOuNexKqLAkc6ry5lavjnXwfvE7cYf6LdUopI
SQt47bFpuPMIXBX6MQdpdLBqxXbq5nBIoIOHpJcHPU69UNTRAsR/x2+GxaWPhnHV
2ceWwe8r1Emc6ybiQGv75zMFtj8Y2kGBmSgi/+lkTCkemdTbzXSAINE69yZGInvB
lV9bN2zqH/ZNZKmAz7Niz/2rr6KFhuDW+D2Xh4p+cnIT9v1iC1oTyRVKpjSZvCWQ
dxGzAIy5OMPavI6a3na/HSCr3cdrMwCzT7HWi+72le9RNIEa46jnQfqxD9rmKF4x
Qxpqy3D8MTpwx/KQgJ+3BabTJYobyS0kLnSiAQIzsFj3HgsqtP8Y0+yncvfC6EJq
qa4WY1aSaU6IeqW6ZKCyB2/0rlxxV3mIyRHbzyFnsCk9U0t3jlchvftu8x82gqB0
FaZrODV3D+ALK7BA0QK0lbAnbC06HMTjXQlojRaOeb8PMbcOiJ0AgSiroiNZhNvg
xdecehpT9cj/ap7m8LRJ5HAJourdfm61K6Q3XJHPugJnmCWon2nNdSyU7Uk0phvO
3ma9dv+zx9qMV2P81BLYVH99hnfOhHlXHvlBt/uYGxrQ0mP9kqnIcHLMpT/YJbXu
a2m7Alv7WAic5w0x4C+LeBS1g0mmkSIM7Kl1Pt+H7iK99Gdgbp8MXBTufaJXclcF
o6xC5+5uWVOs771pBjqK+AnfTjGX7vZetNvFpU5lHN0D50zf20HOHoIe1CXMi5/A
ohkFsFW+uDbCbsT5xdKQ/2fmE2+EMQVx2Z6KJiWbyiTOgDsyYGkAfX80yIwrN8xP
raXankObzp2T745pAghdMlly1cmPv+Oy2RBtgd5yKL4bVb1o9yqtCtTN4FMDCPNr
SGAgTqg3UzHYICoDSfBBiswWy7bgf65bdb6mCg0i9SNnFD7uRLp6+BHqo9NNInV2
Y8lJMNdtDAY/dG2y2qy0qXlmbX8fy3HlAPdmxEjYmyWzxZXTQhQpGhv+Z2RZl7Kv
LHVA/Dr8lPvMV1hLB2ubj3boCJBDMjeF1h1T0EF+1GjEVNcevI+7QQ4CtNipSM9X
7UgeySftJVANo05h/B7GJx1ihKcYM6+HbCDBg6yt6FfdgsLrm4NuphvcdJDTqrV2
ROyIbgeGHUzF9wzsd1DyI66OMbccwQe5Hi75Bs/Psr3D12XCG7VUhPZRvZJ4b+SD
ZXlw5HkB/tjQ1NDMNe5q9QwrTxcVWNUy9YnluskGb7O1a5uqQ7ERH+BZ5BLo2Q8U
72Tv2YLKfSuID5nEfiYdFb10jwlMHtcOgvTF6A7zn8rR69+Y5gkf9eYSD2b7gIFv
UuMIGTkq+hbW9Vd30wv12DDlXMk/DBJa3MWyCw3/kGlufrIdRK5Laj0GwAUQBaKF
vYVTN7H/1tYGVXerWfEA0Gj6uRhSIKtqdWtxjEwew1uEkMeGnnkEGrBux78+8/Dk
eYdp5sjcUTeVER4gBva/AJ6XLUqYhWoNK8npymfFpwm+XYV/kRB1bvN8xzHwCrMx
aEqEGr6MMUEtl3Wnd7076PLFXleuGFRpaVVro5EpSMJ2A/p/SjrbvrRmR2jlDvA2
Lx5heFWshEmy66GsAAR8W+qaoG9P9XDkUam6RVDxNKcoOEti/84t9PNR9b61/0t+
YC9s8Sri6xe0wnP/hK8wvbDyVSHo+5bI3H2FZ57rrTluXdH4Ro8mc7iYSHODE8+x
Y6m14ZqF926lYxTw3//OSJVOWiEzIxhPhfXvbJgQ9iHoliPVD4yqukCzWrAJpDhF
u8QoNPJIb6ftli+6z6tisQYMBZlS8/3Hekg7BIzTux3xyBXUikqc21k2AkpnM9zI
CdLCl1cfSB7aNlSisH85vaFEEKHYIrFOcyZYB8D3OUqSybAB+KocrVWvV0L0wD9K
NhmfJRpcyL6IgN2tXSrkHuucwYgeOO5jVcml9NLTA6B03O+cPO028xbTImOV2ohn
YaXooZ9zdBoyvuFKYWFsgI4/qIQlfMc+GFFcGVoZpQ4TDR2n884motL2VYVS36HL
j5nRnD7LGPi+S4X/bNcP/6jx6pPBy/u3BQydlzb3fz0hsgFgGX/loEVONLhHFb1D
gTREEowcz7vE4BZnAX4h7N62SSdf0X83lCO7PexNo3qomky0vETHJiFkSJ9bAe15
fLn64kO5I/w02UNF1kQTCyT2uE3H/996+kG4sY9q9NTIyGLMwjyGhVpNnR1m3xic
oiXpZ4c91k2ZyG6ZafhfQg==
`protect END_PROTECTED
