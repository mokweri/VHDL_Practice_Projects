`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBJ759vbpnktT9GhQF4gg1H7VaCISsq1vrKCHkBYKzGTYDX+o8ZSAwT/AUDQmO1+
ptw9svbr8OJqrRrF1rnFVzI9264sGQTg6ZG59z88EUMurCEw8d+0ysHEs2BYW+nL
odTLJL3+LZUGFY7+mfEDR5O+4DGBPD76R7cTDF5S/l3WX3fEFMRLwC/vhP5/JqMk
IJLzvGIYLFXRQrwTtu9WygcO9gxdgvRFJFjOETVROwZT1F+guqHIugUO96S4bS9l
4dlo+nGAdvaI7VpFCDhGkwty+8YSGFpdgboZ8er//HOCOJFBA/jV4YchiUrm0ADN
hTwfH1kYmO0Y9Zw3UF2xmNu4FO4cpVigIcCusCmY0Az35AENJ6NZQ+SEU4VsJdZi
oiI26Iwx3KBuJv5XKLDguTNRbPuzrqx+8Z1bm/TZ7BT5aKfQNrcodQUhaoQV4C6J
qi2NZC+p7ZPM+O+F5m07lsgh3Ks0/RwHlStuq6aXLfFvd9qVtDEOrTq3ZP2mP004
lELfJjbKk4+2nRAw6+DPT+I364Guq1jDnvikCruCoyaPZBV+1NcPRq4Lnm/0QAqS
70x7oW8WVDdZdgEbZq7H9cXW9gLW12BREjoX1r6UB3eoWZ8lZecLe1bsOLy/c36I
CMzVAVX5aM0Wu7HaOUVquM4RalRIX5AvLRsmYDw4Lopt7DpqF527nSXV3p7rNibJ
OmbBNnUzyBkwN4HK0rG7JI2B8GQuElDDwdFsT4pf5+aSLkAop6WWatDvpHli1DOn
eXQDxDKPL5H4OzqxKik9eKWH7Gyv44ofOnNf/cZVWt9+z+0cdu8Vi1Uw+V399PkQ
LhJhv2Qj8UEeFIt5Znw2H8RxNI9cfh+Jq7AeHX4ygc3ejwGxlmJ2s35/PjSwW5MO
Lu/tJXGf8pV1ApAUNjjil0g5GgTTTm4YnF47Bn7nFuqIbA7/eS/s4kIRoTccXurM
CT94qBBgtTdCMqNVOIRcwHyj0jWSaVT+zrQQVVsr+7f3K3dxkn/C8AXdkAIopJMb
/IkAvW3NxZZI5KmhHY5bFlWFOa6jT5A+m+vvTdINcXk9KnED/JKhM3zVb6mOM5TB
LrlzgYAqi7TWwU9j/4icgIuGOPfqocHIyUXWir18cpqlVjZyrEKO7IIXQu8eyZWZ
hs9vMifPLdcewG5mKUBKxgPVo/kexe8tTCosOEcnD2C8+T6iw3hiHJhz0RxghnQx
lqa/Ak5OIoiU7LJP8JzADLOi63Zia81xi4L8LrqXWslhD7lcDUR9j+DlwPkW7ZI9
qROcrLCjDoeFHBwRREncmEUy3TRTO7PWAxFNTlGCJwn4W8/VEcvrbP0ZrtcKlOtD
PeQgyORWWulqYi1mDyz8DmDtNXNY2QFtaHJKZytkJCEc2VUzMEHf3uCUFXuQWyU7
079l/q+hr6rETAxaxH7uMNHfcaLclxO4cZpykFqoj7hO1CUGAnxjzaj4eIh33N1z
J5oCjqAer5hskl8W0GXzfNXqSVyj0gb+iFXri1OIdmyIlXxaTnfr/K6Kdz6k0W/s
7swT0Qxm1ZQ/v6Bj12LxJPos30pQU07lNVK+N21HvP6quUH9FA3LfgjaEE5VF+Lf
EPgNvO6l2Wt5qHNKmQ5vwE3UWbEbN4oSq1dXeGMo1fmj7zR/QlV9r9ume0WCA5e9
fBZvmIxg3btLvqD6MjZfEzvqGP3f8H6Npim5h9eXF5awo9ZQh2tzrGS4+eyhznNf
tHXigpGoGOK1Ud55/VVXHboM8hFgC98WO3ZeVZN23ayyR0cEG5jdWH0cnNkC8iJD
JfbtvDOzsnRLGNvq7KbIFLmDdIPKCf7RIeVjPwTVegUCPPRvdtFlqAhZ1sCNDjBi
ZEpkWPLITH2bmu5y8NsoA+pixZLgFRr7wj80ETJZfKolnDuC5Y92mJY8H52EmQFw
mPNE9AcZpd3YY2TN9ITKbHA2zKSsJ6vsPbJTUEWzA3KTtjcE/PcF+5wYm6Tg05hQ
ehIQyx5tuA1Rjz8w8ZQL2FhxzkyxYUpQVAdBSjDKUd29Piag9p9OUU8dpZ1z1wd1
08CSI46y+UPzWr0JZjkjaQA3VTgUfB6WqkmlCII8h8i93tkldLovqWYVLW4xcT1I
98YnD0lxmHFSFtlUGmSQ0/Buf2s2AGmqfIE/v7eMm+gkX3zbJG5Vzm2qCus+5IAI
X5JYhfdb0u1oK+DxNbEhCiGAIW6y78X7L7OGiR8VHkynrBDxf8R4ViKtvAycbUjV
N3Gc7TaqIBMR/fv0wGnhX7cJmJ8g0KiBhZPCpIb9SGy79xgEbcSeYVlLf1YOyM1O
Q4j2BgWSqkD2Qi3LJDWcqu56oMd68fff64r1lQWuyYuvkorkRrr/3FH3zlbxXy8t
o26QnqNlDXOv3JFdAHSLxWxwd4sMIrxL2zOZdCA/k9pukNwaIs/MQa4TTZNEPBpN
VQrOjED6u/y6PDgop2Ru3rply73PJ49Cu/eOYf/1NbM9MTYEssbBHck1C+8jPcFX
2eV6/DQ8M1r/XpfLzc73pqEq2a9fmS7gq5ho2/VOicAtfknVhrajqVn0O6gRc1ta
3A/JX3hXM8ehHcXvtJHlQb1XP7Gx4hY/y3uoAk9ZuAc4QZPjv7aIOBJlBZAhlJmr
H9FOD9eTCOHxZMOicOobNmu2+tD67eQ1/dr3ki3WXDpEFWUKFYi2KCChMckIgwvV
V/h4+Gpfjc+p+E4ZhFzljnZBbY3nhOK5X84OATcgbqWgQDOaaLYVUXS/7fH2Pif+
8UQEqFbpkfz8OJerIO01lpzk4x7LpkOKeX6eOKxlHfRs89p/7ti+E5FZm7UkfXpc
+TjGTeznO/WmGQCt0aj2BHfNRVDrBqUgkIoWmkWxEg2homtVo38EI4FKg9zD3Ygq
TX3DfoYYLMqpZ3db4bA42VtRDA537Ru4Pcs6ggLSzMVRP8m1bfMfYg75mVGfk98Z
XmMfhl3xzMyCQIrb7mkt/jEriFzYGEeA5wUD8PfRJRKaQDKJSR0nzeZlg1GaidF2
nPVJstAEZd+4rVrThBUbWfW0KTVaH0Ytvh0cvEzYh+r2lA8qBm5aAI91qZl1G+/0
xZ3lJcRzvnRyHMeWF3FS5a+sgglAVTFUT7n+zH7OWbcYyiXEP61bvyHNvSFZlwf0
5UT9cCVIx+9homjwomo3ywt9ABIVU5clf0wjyWbZO3ixifl7Le0h8OjBme1JI5jv
nmcNlYNaX/A5PaWhBHVPoAWtvUDZodMvJ2nxHOzZQ40PUESoyMIXkelzEK87lrGx
lQSjTUMAhvElFwrlfVUkhP+gk+IYQjjgvuR1TuAGS4oqI5a/ry0CyCS80GQDi3/c
tqoOCqsZyO6af+NuU1nrdjLQgtACJELtkjmQ4ntEHWWuq84vflzqs8Z20prySF80
94ttLGAMGpBccqd8aFxboD2NlF1dGRKDBmqOUw2No+owyCqUyzcbGJqXoWJwqyE0
d9xHQxqnOnJEc/GbvKsutTaOGCOPNsyoYFe5G248AjOfS9VFMxX6pxVmZNiq4Rvb
jASp6HXbj0vxN8OhhbQUiywF1dJrjOT+8DPzON0Pf4/V+ZR3FemifGPORPEfiN7V
bmypVeeASHof8mprzTGFCyovNgfFNiJJBhg+HMUTlAfN7WIL9xBmtTMygmfBZ045
P4+2XR+PAkC9IsSZWxM5MWtHv3jPkbFrMhqjkxkFA8/4sVM4nUfv5RsfKWz2a+3M
Ey3AotI6MCzpnH/wVxu5uP6hn5Za0p7UA1BfitcKF3ut489RmoZLMgOSkzJUb/Hj
d/ckCkeV7zRcbrGJ24O1XgEX88+tko8Y4AqaMFS3s/v+0ZS20BrciX5lRJL94U3+
5ueAMIIOiHqbC2SpOEtRFDEmtEUj77J9+33/RLsXrusEv+ZWi0NJEN4jcjp7M+3z
HruzL0GCuTDaXnR+iUlVcZauyf24pLa+U7tUb5z61Gx77fM2oMSbRdxK/VAHG7ar
1d5XBezBhhTyZLZghCcF6gASMe+y67nizMhkNx8TB7TdezYDuTCb/PZ/POnsi6cR
64ITZ4VOB3vm9DhNRW5vAUbF3tp6Sw2deGlHEa4jaq+bLbEJzflNu3n+bqJKom69
ZJjTDGxel/gbDkGwagJKypKOjz2AW2L7QEEIR55p1Enp2fbNW6F7NN8MWmD2v3tC
hgFah1nIZiiQvlt0ysE1cFuoG3OpxK6SJw9krhZR+/RYKIwol1UEBkYNQiDM3eVj
8HnhWjl1KePDqyzwyW/KSSsk+Opf1XaIqTgBrDxUyyn55DBKUCWsaMyUHm+K8u3a
1mz6y2Q0FVkDbwVyWR9r+65Vusvd18WOxQ0MxA/dbqJldQSr7coSeX4Lycmp5eeb
oW3K9kBY9/9MgYSqP3csEgKPLKRFOQWi9nSz1VN1BVS61szY7si89JIXiiO4oFd6
AIbheU66P/IqjKNUejdlhrWx3TIuhJ5m74Uksb7DlEa03zWvGuPWcWXRQOx+nowr
k6Ah3H9bD485ZI31ErL0L+NYA045RQnbDNpNLhiUfDyUm1pEBavnOEzVWZt+5XUb
5LvVnNm/uV2DKpdpGvNq9pRPD6VHuugWEkSPVMlLtqHG5b6CE1Lgy4Ys4vzKUhmr
D1glLKsPdbfeDWP7VxrZ0qHDz05qdesuBFnD7P/+y0X4rpcZZyFmXZAI/7P6PHGQ
YuuTJgYT/iE9/DBVw8k9+o5m9QuVEajF3JWIIWpdtRxI15HFnYyYGyTS7QsQmuLo
cEuWFlE4EOmtVauiz4t06dsf4DXBVWQu0WUfTIpemzm6wlF6hGhe50OGTMynPgnm
2qwD2eSt0cS277LTU8Q6WrSjJ36QRm9yyrKetpgJOtFrG8bNJbroIf8mM8/7elQm
7BDQ2GssSpkp/+GXCDR/s0SwP3yQgPQhOP+l4rcspsCcUW7B4XQUXiwN+3eeYjQT
86KoyyCfUdNu5XS5QxSrNCeusBw7ykDzABBgXV3+NYFpAe6OLRM9Mlua/UP6ExpV
xsc88l39afZ/SE/5oYtbEqdYJTA1setvM+C2sxpF9SyPeT4uSbHHxpffVdS+QVvV
fepHmCNxhXDmIlfsMlqRjsCxBt9zZ3k35GfBcUgdMLdgMJJRGfoQ5pMJaaxKxosp
omxCWaMkPGxrfQmF/pLIFd3Bla3vccoBegTsJbtTgLlm9onUWtzPn7UrBUl2lY61
HPIvmmst+AbNEre1DFGsxgg/s4lHp7paq0Oii+KaQ+KO3S3nPkF3GIzCWPIsfhdI
Y7dbbqaU85tdCFApYQjW0CnijMhBwOp0r/bGqSEgwUD/e4sHxG6BtZ8XRhaiwHuy
6uM7bb0SNDcjb75tWsfM9wkVTK/j11o0ftLCCVyKctpogwN5jEhQqiYiGGQXTyBI
x3ZnWkXqYYfvLWNouNk/MESx0Sj53ATx9eq95QCrZw4LwPGNrnY38ITopsAKyib4
pmgEJ5o8XVAC744ScsCH8Q+g57xFEbVi1oG7/sWbtzJKQ7MJ/SHlyAIxYGh1H4lo
YPJBzzMqZPjv2QbqNVj1KDYWUma4PycpD7M8WUBCS2ZrUTuifb1OOQfMR601uYaA
pw/H94KWp/WnQsGUDkaZs7ETOy91PUQNCRwJrKwmh56cMbuexHwy6fUkD7HXY8Nf
glt9DflpKCgvDFf2ERCZChH5aVzle/Vl/AuUjRMyv49jgkOWgl7CYUY8Pe2mw4Wa
Qgnz7eSS7nYRKTBabZ3YvPWDhdGAVUyDDlfd/hwzpeqxvRoIx8aiyHCr402JoPIM
V8Ws7TCaQGNvLbNCod+DgdweDHe0sYlv2bbe0x/6IuSTz8AissmzD7OTIIcGU8dt
hMvzvUMdi5qhmvB3+xxlN02rFepSjqybqWLVvWLnoj+/ITsl0UV17cvbTsTPAl7R
+Jr9JXJbEFOd7oQXsSKvI0z1i3CVjqQrgPkpQ0icRPX+puvy1RmW0WaPlI4MtHT5
ldGIx6B/4GzODcSlEF/YG0cQEOIEOmBaWbb0zFANAVJ39dBHftpDzz8AM6SHYbuV
SkZJaS4P6+OYnWldKZ/XE9C0yW21VzY40bqbu6iCCV6HTo3Yc6n3401kImlNtWQ4
Qp++Sey79qpK2u2eZrNc342uLN46dWfV6HGuQvQfHnjRSIrsEObcH4uETQUNpeEB
pW72VSNGfltsf15b/jWm4J21igL5nxT04JkmSws16nJPwjjrZcANmkQz75RPuXHs
1In6QmPM3r5UqQkcy1aN7opBDw+LKf+cTCOG5Wljs9t/F9XDT4XQQPQ/HcratuoR
7IVRY4jKODcHUqsk/fOS8eR11y95pCkIQsh2vle3m+LseTTMyUJ2qrJ2cu8W+Ye7
7MndTWfUgkXIRIChKtzzwubxu8KY15FsGkEzcDLBsCZoneFIxhFAZNI1lr2oOt7r
jPt3BzGYu+5Ei0pjgjIOTWwsxvwwBSIGbWFKscFkXjkPv/6qGxaLPpFekrQNBcJn
47om4t2aP0UGCnmPSzp9ITQwztDx6Fj2IAo8uKTkeBS9FCQn7BCSe7jCO7M2z6yX
w6GdiV7dTkhUw1aV3A16BSoVUBVJYP+c0GPsWXFdmsvZh8+LctwQBIkjnCR+0y25
RIKD0V9MWKrfpDrdqeQ3Sru+kDCgTIGQZ9xWnvJULMZF6+F6Ndmihy3xQKilzEqS
lgZjp+8jxxTsRzfkva0l9+jiK4lw4IiQjkgrvUZlcY39o8nb8HUImBKPw2py9Gmx
0MO8VZ2sO1YTBT6yqiwjoGRmtOINaBL/Jz9X3+kHBsaHPmx4j+jOu7yV5UNKNpQ1
pCgPw7jCEsz3pczPaSHVNrgMuGTNJDvT8YCvNXYCgUhRNr7Ahd/CmVQYI8NZrL88
mk1tsqCwt4bNjv0J0w/JHwqQUKiLnil4cTWCOKF05oEpKV3bFUNX8EQ+rMVu1ypt
9QTbWMduRAaKzHjuk6NoNJzlU5lOqorSe68fSzSW6QOKszBvlFdBTSYUAdx8/gzZ
BWTq4++FjmZ+zkEJ3+o4pynmdhuUC3wMllKTcu7z3w9xyu9Wq+7Wm2he/VwbIJnJ
YMS4OaZaHtdMSGwbyRwSpBcCanir5tVCsHa2Q5CF6bZqyca34bkjNp0/2YGEMJ/L
t/uQC/ig3qPTSg1GA4n1EQphEJjX90jR+bD7Ty5yVPNd6/GNFbO5goHgn24RAPZP
PPPMHWoB2Qq2GzmGCztKR5L4UTKhGy61lQKa1++QKDOOT2yWkqjdXlJgu2fzFB/N
eU7zW+JxmwWIo7KUvCTO4/3oDvguUc0S1UfrR3hyRI4ALIbLPcXuO4OzUVZiAP2a
0/s+w16MgtNW+knedY33l5jSWvkAmr0rsNTvxY0u0xQCP6YNVTpZxkDsB3tfBQBg
f2sDa3dofiKMsPZIZ2aUajuM6uIv43Ks5hQeSVoTHkVXX16y8OjKT22MtPvZKEHW
Kj1i7CLqY5JMGmMylGWdGE5WfBS4RrZ/OP0tD4zRmE5lQhv1+LEamxpSwS/ewCrL
v/X72piL9EfKihulIbfG4d//WEegyxFLH9VGtdgEtUVWVZUT193jmnPFAxzX6kC0
bOREN6hSxONKnRPjGcDOhx7fyZmLuSesBkOEGcmly+DBSKLF2xwGuOjl/021IoiF
0CvL/31I8j+MZIVH14a91NZSBfP/ENUBBDdaAGeeHMd1L66gJXYmQhmNa9OqxoJO
5EtV0Wz3DvPbRxVpszOAe+ICGN3ID8y9rghRQQP9xwF8u/R+rCuMZ0g/6Qs3TOKs
2KW0pNe5411x59a+6AnFNIbm9TrztN3fY1dVxWGjKaj3piYjpoH/S4bzhNup8yRK
QImayWFCWbEdYXfuhfdQxE6G8HRQ7GPPU8DSZBm52ymSSXElWq1/J8eiMUdPPc97
xf7HKzZL9O1n22KtCZTeV80LUXaVFXa5IVtyF8GGVt55nYYKHR4atvrcsAcjzp8O
0/zjLzO2lU8XOb7cbSuiFfmrxzcgki0O7B+tu9RA0yoJYrPxzBnZDhK5gghgu9tp
nfKm0w0mArV4lsO7MqstdmtKYoCrQz8IUvVqQjS9Niob259ttRwYjiibobM2+epM
Kjng8zqLGfmU1UDR1Hq/TIe6eBdYdN+2EeHTL84uOOazVCoxwV3ztL9FdNbySDNa
mmgEgQWY+e/3BOhl4TuDI/TBzhTChuYnyCwywR6pEodgjUNazbk+eDBhOjw+7RAd
zKV+0Sgvuf3KNX3nHG50a1d583SuimkHUQ9Cbuw7Hb5xUTREmgaCBPcR2xaZq7/t
esg/5q4hHgDOdF4UJLyeh+7BVVI6s+y9rkyDa/EGNlGZDFZ1F0W/0CnYaQ4UAdDw
a0YAeiCBP4z2VU+QikyKLrfPZpQLm6oAXlfGoStmVLUJiOuEQeBNR+4dvj0lnePA
MLrFz0h3R0yYj60JJRkEFwJOsgOx5bmVhTObn5Yzba5Gqh97dcG/dRauFgHijik9
FF5d1LvcM/MSoaTpiTha7Po7m+Z/MzZik2NGaQhtfP8LBlm9AMuFBVRV7DwxgJWy
UdiAYYu2p/enFl55L72QR023ITn1s/amisAm4SIAhBTMwN5abwdV8rP0blpx+EA8
cEnJpV/jC3a3lZ24jNakYlS9ni6YKX5TG5digh8vI4djwSpmiLkAlqMouDvCVJh1
8EW9EzqfB9KxD/IMRz77ziwq4y7GVVYlIOKeJvlZ7dFUZxdC5u87IkjrELOcMUvF
eBCdqDBI8J8h2+eKC6mp7bGqlrCgsY2E8hQgQniuW8XUNvyxiOTC7VfLqGAftnSq
NC3Fvlko+GbJruzu0ZB3L0fC1d1JeR4P+3B6SHrduIPEZ61uKrFh2pq26rMEaR6/
qaIr/hqp8Til2B82c3gOl06kId+BGd16P3EqPWHPmGQaIoOGUbhJsS7TcjhJTejY
mcsMmJBVytGyZGcuj07UB3DO9w3sVZDjCjWNcfV4Lt6HNbe4p7rDOGuxlfIUWDzC
cR02sco+l5slq6oDPWPjcue/PriPA8bYjutKzW17DC/iTN+lP8ieLutVT/h3Qu/Q
rIV8ifIebmeQh2yJmg/0Cvh9i/W5Qt0dpRpjoBwXXmmdhqt0TLPLoOmvvSQ6ZfgI
DK1XP51wPGk0yIlCiLeYxENqYij6Ak077hT/xc01kojAgSGgwN9kT+zaBDYYeM74
pzcKWPug1UgVBCtFIG9+6EsCW+DaqiFlv/sFkPs6qh81nxaIe4AyvfuAmcMvtcuc
Kt1FZfSUtr7lPBkbV6ePUGkxuNX3eWV3Xc3rBhjvs9ZYk9J4aSZf2NbFYQbeEKxi
BinI18ubPw/hLW+9fNpTS+PV6v9i0r6oIU+E3csAfnTrqMMrIrn0fjwxZGrBiI/b
kVikMRNtl4BKlG7UJIdfiqHxUmSrCAaPfd8D112s1lWLhezy780mxZCwETeDXVnS
5yCcKzgYyH0kqDcoaLAstWEO8Wp2bv1Frl1oDpIXeCgI6r1CGI/e8/pfAIrb6Kaq
sWFBTq99EJcmZvfU4uJYjNItVTebXlTo50tUIxvPalwkGt83zUYyLwpolx+dHqfP
SfsH6mMN00GK9XbCisc4fjpASwWY5sC8WfZK7GViS9f1ncjQ7abxv5XMuU2GoBvU
VxIGLRDewbgaCkZj++KZGe5G4xA9ggTLRHReoCulHowHQrGeAuVdFyDCaUGOe28A
jRmOqIZeFYjx9xVVdb8RP7SDnAOR6YpiiNn7Xxi3My4IvsfDIjFK0M29iEHtDNrC
+WrRI5ag3cSMgMbDoFvGQ4eO6OtxAO+DlSbeCm437x0+g4QW6U/Blrw6f72KzD4f
Henl7wlsir/5KLNxR0QV5cL0HyudPCfjvMcq3meTF2eirQRDUssPqtyWYuosAepc
ZwdVAAC/OJilzpRqt3qKPq8SZuah0YuInf1X8vdZw8+ZRyuj7nH+hvQhXM/DCZ6Y
XiNsYd0ei1U9IURdzY4ViwejKFslY+Tqyq/WpwlY+7TzHc6l98UcAocVXtrAJWIQ
k5Rk3dIAswH+kfymihwLyFjNTcq5uylfZsQOizzZZZp4cpeW1B/TOMaEkDg9jH02
1pCE33eUjx47OSlDBk1orLf6i6TM1R+mL0FZqc36p0QGJ7sr+I7Grhw3mhrIVD49
DcGeH6M8mDRVSKjfE/nEA+bHrmpQ1EcUzspLizgyIkoLe8lRuqPJWOJMXBgwUQh8
79G449fyIh6/LZ8ymo9GdvfRIz06LDMDiK6HOT5C57M7ZEtwXzW2OrooVDmYX3nL
f9qI4/3C5Mrszb2KR1TXCckgKqbkkMk966akYCLA8oZgXEmCDpm/iXjLOM1gVorO
s1GGSphJWrbZBAxWrDAfuMnSBU3BKG9ip4o4vfhexIlyBi/pWiOxhgsouzP92Ixj
//EhwWsr/FT/xMRoSdDkW5rYqyrWKrAM/uGqhoQknDVeIq/ZYhUkT9nP0PkyFn9Y
srhXVEH+1xMJ9Qz+V6aHtiWiaKx5wRVRUdr6ZUJGSI0NHB4QvI1bTe6kL5yMkbJT
dhxgrTBdfBHs43Y6/pB8fFN9sjP/36pD15udqupdssP/zAshWJxcX9zNpA45rGSW
qhH61w2yBxZnurtgmB7RNEoJyQ7V9eW760+G6YLSLurBqvEjcBls9o+cthLpf9n0
EDu8jMux268t4iGG+c9cDxBnB2YEgUUVWn5RVRSLvkXKsLwqLOdgSwzRXdb6hpYU
C5jbQKZU860hWTcXoFuwr8q1wlX/Dr4b8K8DalRsZ2/2ley14XRN0cO1H4t8fX3Q
FzivUnZbPDVGtucNBRICj18JGQ5BJGrx2LfMZeX4juBuJKBZ3pnND//r+SHSVRaZ
e/5dEsnj1F8BiEbn25RqlVXZIPZjwd3WrimAYgn96iZz3U57GKwT/Rs0ErFZhZVd
WgTu0gF2L/knN5QM1ftwuAv11z/FQez34QHecCYx8j9Vof0HfJfDPX9+v2s74MP1
bsd3Jdk+zwTQrnVAVYCA385f8gF2Bmz+T8rQGGX6Eg5v6TIL08gKHzantvwzT0md
bY5hB1Z6mNsWSvQ3Ce8K/Q6jmdgVA3pwVZnOBocL7AXUvbSizKomVd6mLAwC3X2K
kxJR7t2umY0yZnCXAO/GD14ghf3LeuFoXMcJGZ0ng6F3d6C2BooiUMPTsH2bpWwC
p7JLibEGuLxA6g5qzYlr7tqBBGJv1js78ZbH5cezBFAryB8piMy8mAExzZbm6PhG
qPYWLk3EhY9RI6e/aAd7nZiMwY/wrdWrRPl5qYWwsJeLWlkDw3n48kT38OIY+xJV
wSQhC5Mj7/6oWpq5DRC3jgiCrfgziwUzkXpqCL9dS7IZErzN80YLQJxIFXqIQ4ik
aTEMAzDJIvU9uNU5aDnf/C4YgU7FH6iVG9NKMKlY1tmGsleVQUUmW4BSSkg1SuMX
HzcNmrN95OE46mSOcPkopTsLCDRFWk72+xU/sQTPJnY2gfrIhboIjo2fd329/WR+
HFc046Uj39bnHCp0T+QxFD+r5/ckbhfvnWI7/51kBqhqxs9drQ8orXksRd5Q+NAY
/I/kHsp6DwjHDSs+xmPS/zEXXRZQf1OvQPDuGUmTV4neFdJy9nGS5A4geZp8zllH
Wi0tCRWmVvz4wh7BnmE7HQ0xIDUlqykRHuJIntx8Niz+wb++DDuhiVX98gkH1k9i
JRc1rnaPEXMbMFxYCau/KHPCj3rp9FrdMmeejvpLDEegRXFe1R8gK1KmpeMwYMGa
2Un8bvfh5BaGMbG6w8o6a/+s9mak/TG3evHJVlk27FK0ziuzuknhiandn4+qUqhC
ZAx5aEPAbtwgXbh5+HRp8KT/tDKf+YyVB//+Bk9vs5qu1AGhG/mouVQfpUi33E/S
FTWZ2VuSOfDgpyn9zsPkk+6PF6xiDbEg9FnxjMnLjJReV/5wh6rFaglxeXwoEJgw
n+PBQPkmiwkeOCu58BhZR83zO0zuszT/zNlI4cV6JZXukqSwSdWKIqGNTt8/hRL3
FaygxQu3feBbGxwpWQ1olQEqAoU7TXng8J8qmF9V0BnFz0rMlgAVW/8gmRQMa87b
plgxfOCvLUk+WwkBEwD7k6Ft9b8sv9aCi60ZuRbFPy942oPX5blN6mvsOxPOvhr5
Ql/KH8dEfF1pARxBSOggUpWgPyTa34kNjKjmItXvlvJxcjLw+1EZ/1W9lYqlCrfB
AuX8qEwjIZJ2Diqwm9oYxYX9wnC8v66IkxFCMv9hKZYxW96T4X0w1cwWJ7/UTSma
likE3KVgRzC8YSg8HI26RDQFK0PO/PDzxBhK8HnOAi7QFFrA8Zpa7PVNAU+FraLt
FfIkvUv3C2td9r+kOV4s3/Q8iRgSgnXiDE1+X0Gp668W3hs81W0TE6gbA8VypTPM
GNLHiXGu+HdjaK2o9M7h3zQWA9HWPaMSiWTbJXKR1ay7EsoBnKIBoyapi5mmPV0S
40EDswif40EOnyC9XP9Kan1nLWd3J8YaFKeBxdnrsKyt//GWPHO1M/D+QiwYScG4
PoZrKdB18uvAyvmVTur56hwyW4pYUs+Vf7T6cEQihnsyBYN51GgyHdOP28UJVbgE
hdGWmZcWn1daDxHCW/xamb4yjMCe3xoO7fN0VNsR5aZEHQ3CeXd+p/kKAo6Rcfg+
67m4DUvG5FlnS13srLdkCBC3EECv/aVgJmTxX5onyyNj+1syC31+gJSj3eZWRR15
s7MVl20GXXyAlcnCcKTssxY4VPHM2Sxt9tPxGLXMlmK4qFyGoNxrmZC4Xzo16Gwh
qbWGcTod7xsFnrZsrq0RQjG8tyY1YormVpkjFmvRUEGD1QKcUlH+LrCOJOz1HZCV
M9QyB+dQrJQMctFoJcgA+sghLx/K1ql9bA9XB6w3rNHlB7suV/4F9FDDdBmmKazc
BRh+7v5lUiIekdRgWSZ8zrHZTWXU4M4fNrOdg8Y3IZuDUphsqBsH0GQ1tUwZ9jQ1
Jg3UedGRe+6zCKF5wUlg9BINtbPXuWfE3NQVT5W/la6kM5T9a7aTQ2qa3XXCoORm
5yBsf6Y37pJRqrRcOf+Ce8WsfDSGloq2vp++469otyofeQFvQiaqZBuMdsB9HsNg
GGAYrRKnmNOxchcEABNrxQl3AL22BxRPwm65gsz57hD11ifvOry6XWKjS2QQ9qWD
AG7PMmX75Xr12ZBpMFBs+YWz9jtbSfQylvXn2wEgBaCb4xCiiBxTrNvZDkozGDtO
KBIE75NUz7vxl0a5iwMTapUtrbzjXc2nN10H+7tgCz3onjTSRbOP7YSR6WSQDj/g
pp6GyDEBKztVFV0gfOa+7K9IpBUdk/ZhonpKJ6ijwNPIZ1Pkh3Eygc+ekwW++RwW
ECybbYREbWsF4KuBWU6a4Jb9n9eGxG83XxntJcCQw0VuC5JqS3hCzmwTKjEXYX8f
mClcrGdNG+pL0C8PIf6luNUQ3PAQi2yFMlvtrJ/01mqBl2fDOsRU5+Y32DL/K1xC
R3xJ/K7siBJJFLigSB7xZjtvivo/7MUSsVb74Z2chMoYKCv9qRUpeoubYt4i0b/Z
l1ldqBJ7PGLLJ3VISu6B5fBmu5h41s2ww60bQgLhsZyIBESguBBXQzVGvlHUcv6A
2fyLf+RvLd7cetbxDs498V4YxepDz7abXs3W/9hgAJs+LqBxPEo677FiZpFGvQFz
19ZgyoOHgcwr4ChZ3OGDn2plOslPpDVtDYqN1yAlybqGaakUcH4xB5/FQWajv9bF
KwFgag2x5cUlC+oLi22Vdt3dasQwtkBNv6fig/3FwnRDf+GTimZSqypQx/WxD1eo
cdMNDOFPFP5FzWJUtjKHJ/h9LCgUvuijZHOQKyD2gkJ1GnMhD3/TuDSV7qYSUypo
mGdUqYLtWSZ4eOFQ/6jwcSAGCdT4LbE50+bCwHRIWAhENnEDqFpwQpHekUgEr8ed
urXmrP2MIHWK/n1vIpUvYO5h2uzHjKrIGqinrAVXrICgKoKzJBbXfR0oZQiw2r4p
INdbLjKAObiAue/3wNN9ifvScHoBgeQRLSE7UbPQxRB3AQHyie+kQPVr8kOR0xmX
jnyjvOz8SoNk2l7XZNCunZ63O1dV+ZDTp+8rW+Iyiavprb6TrC4u6fW5TxP9FmUB
f276hVIqajXSrVENfEFHZeXvqCXD/Ts8YAEqehQ5HkDJ82SPFdwWJyRqjs4E6jaE
Qsu3FYQkAdNRYip0BRV8Ouhvx1oMZOQ8bivfxWuVmu1SG3ihYwc8bjAokbvCLkAt
5RqJMm0BT55oiT+wg4UQ6kEhFQ6uykfhLFSCEc2rLvJh/fRYXOHBuzH6RGElBiej
BwWemaojVg++aplaG37upr57nsrbc8sCeR/iI4HWs3v3OHWaOj+SGpvynzutbg0R
39gb+SoqxQYHBou5r7YHeScntknSvaVC74LOccz9fEaUdLTvLkgahv7UgJ1oL1hU
1Amz5veRenhuE2c7VSjw8K0B1NwIERKxy81Vl2jOru3TgS7vKn9QwENF6zU1ufcC
yzPAvkEBnHwlySuwK2+69KL1O8LbZfalg5CInfYBAczx+s30uCk0mEM8XwwAmlLE
7xRWk6BGNx07f9552k5FDcsbVAsuoHyApGQbRgFYgpLHduh14Cc37M4h5L/qfk1x
WsxrieiT+ohnf6FKEN/rQ+z1bchcQ7kTvNGu7hwLk2bzeHagf7O23xiNie9SUYhA
blEYazh/0wqaTuCq4Ns9qFQLjTz5bdfozOsBYc7RHvwWy55tKtRsVKYT/iwYJ7VS
mm9KIT/dphDY8pMbiS/TvHxtGIKJ5mT0wy/K4CnWqzZEX46GK845sp/xRtMDAGVx
vvG/1UZT0B6D+BLLlTGBOV9vHSpOrqUH2T0TBSFaDrD3jjJDU/d8YbVk+FQl1Cre
sPaoGDSEzaIL5cX9RLpkar+WxpNYOS34zklxaCRiV4qPzJ9JGjRXrxq1HPELTVrZ
nXd0xUAfUHon2vl/6vy3jXEfvfiskXXqZdfD2TcVTq61HS0JytuSWMcqkroPrXCS
zY/aFFIes0pZaqpNHk/8sK+rjrLjyb0Nlz7buR0idYCHDSzjsnepXePVizqeN7wS
MQlQl6KZHxe7miWHbPjkN2yAIaIPNtYEEonBGrCoXR0BcQ+B8xAtFIrNCjiONdjk
wYLzcD3XJvqRF/dMXcFvwl4EGXqsxKtjZAFLCW1WA0fRX6EmpXus3TD/qgAQmGSg
k4vBj/sNr9JCnOKU68SeoOEnaqwucwGPnRJWAL2fKxG5PSLJhqflNc1D4Ro7P6F2
14qJHe9ZAIwIkCkVTKfXvoQvoSBoS2/7Y2gyp3ZswvMJUdLmfEeirRtStf1mSQZ4
99NKxBC3kxjwNBhAkReaPA34b0vVYdZLXFz69Oau4tVV8JP5CB1NY+sGgcU6PeJ8
S2GXAEgfzckb6CHCzWgVnZySPQ4uECernu6/3T9PrUDVD+fziE4NegOf5DvITIU5
v17BXwW2/PPGbZAZk/ZXrNm9rEfK7mR16zRWdpQ7ndbEJd+cmqqnWgcmr0ZkxpEe
D2SiAEscUKiEycCLYB/kfztfHcxjPo5Xouu7dCitmIXk/l/TftbS2m4lyPWbsNDT
DXmwergJwtHezcLzMgNOgCkb+K3QOMaYIWs1nwYqYSTPGXDaqZ6DxRRCBLCHXnh3
IsKDszQDqb3eHL2XLquPp3Z5fah2ZULCRvsNU9HMEWrULDZcOF90ePDqN4+wIVDk
cBCjDIGQdXAZB1EOoBNLRcelCnG0qn+8ITpOXjUYPaUDBPnBKoq/tTgVcvvM1bqg
yipDjCJu0kSBLEu0JsV7ndX0j2dvsIOIbozlRH3WaWqXMhAkJLWSxQT9fAJhWt3M
3qCpB72rNJ0bVMzPNMeLx6TENIrleBOTKanGKy65P1n91sTBJ5Tjic+BQaKF3D1P
Q3N8IesyGsORsgCyuxWP2WE+1pu0kIHA5IevJB75czBKfdnEAhJft5FnNRiD6T7f
MZnaHHoUssWuMFEcl/qlJ3X8RMYYSVZ/bN6+HSYp2M+zJIgYW0P2bz2m3KYT+BBt
XekgTvNnME4zpTjTQ2Tl8Uh4s7kPhhc+ndl7YVRmHzf7XTj3fLmdFcOqklo/cdRl
SQ6fSjHDXmpr4kMwoh512By5sITQkbUABaWzt/cU1255bUM5M7XEY77gIKMnR5oM
03psFTn27zB41rdyyLb2wtKLvd3JzDQ3pMdfiNWs6eQIeDRvcAg/IglKAZUz+2uB
X/x3dTks7KcSl5ud78hW1q0LqQyAKyYKCMt5zRE9pMitykTemVtnvxMDmZYBgpkx
PFiB89I1ROZ3iajn3RJf9dBzo69pl1tepRVaGmnWauvWQFvMi/AX/3pPJC6kmgtX
jYLFs2rcrI0Vmi/uQ5u4+7AyOF6r3famPFVmeRwB9VuSBdvZLpbhG7gIhGs6TN9F
eJ15xqNxSkHuzA0uk+GLsHXTsRT0KZYo4q9+RYpMeukSqfOgrvN1fwWMuIVp1bkm
nzUnv3iJT9Keggz9AjPgW+8ULnws3MrgKzpzgaL8cZ3pTgh0dJCh1OoQrOn9qQfy
3RbKoME2EZq8aDaESmya/W2Onje75LGKWuozxI2oRl1LQf+UGpXQNLWz4N3RrW7y
DCfzH9c5yg9vKZ+G6JzwIuJtUrDhtkSiockqS3Q7gGTgfxCgudtpshKtDAf5NM1y
76jsLxj5KvAvd7xM7mZmuRn3kVE58mLhsuwxCSb5X5cnf9O0ULmvzvfaci9bdQ+W
nVb7xUf5nzt8S1bxMloRQtw3k4ebG3ioSX79n3xvda6UqM3i9Z+eHMnaGOw53REq
6rQWw3awVHhnNukjIKuX+ZljV1qfNV3s0BYpPEm+GOZxYwG0YMlqQ+GT8aOlrFZE
EsWE0pc/rBnewK4emndtXzhCvH+CZ5McuoAyCbnDxuLU8jNHEBxVUghpdHFFpbVL
VF9ZNRPlr/DzFqcMzsRndJMeUoypr/CYSgANzbhFIfu2S/mhpFRGkmZVUNyy6sv+
DbAQqoQshaoStj5obmFix+6X0wZuDzE/j1zSwcCApTS7Nhuabtz5fhwm43+w8bkB
vwa+NyqRI7qCvCWXlbYrO5RXdBiry3RULRiSviMP3AA48h5ByZ3fx3bPS+bMDL8Q
/UNR0m8r54Pi9iNK5DXOmjWJZp6UncR5a+72s9AA/mTeq5vVCCOWQ7GX3JjxfH6Y
SWP+Ciz42OrVZu4hBfVLkRfZuFYyQOeHtRxDuwg1pfYXQUbzGNGlLEeo/vaELF+8
XRcsxchZbG+FYQ0AGqw1wgGL4jEsRgM4PLISM5oxb9zCM7jOASP0OkVRhN9ColTw
T2X/oL2tv/LrExLBQEWKlI50aToB7SIz5zeD/3QBRVji8tAwzuAwMi+9r3jjFgeU
R0PND4VIFkre6cK/lObxnj0wL868dfa/EbwtzGTG18SjIyksRCVXd7St64mQ5ep8
4oGlpzDbj1SoCJeOpVJhSYv1gIJ8DSjaN3kv4Caccj3bXW5dEFqo3I5Xb5PaHBJm
GqYxdAsPswoImeAWg09fzInFE4b0kNfxc2Zc16J5OmG/X4MOeQxm4aq6LZw5KFiA
1fjLnqQhduzgIB6kFrg5+WNKfa7wd7Si8LtS3ZqWGlgqS5tAU/Gnwk1sd/6Ovcu4
9qAE68rbXcFYu1CTnwwYyUz7b8F0hbRDFzK/O+7qc3ceS6qAV5QqVS8+DzuV0H3f
rWTtKYXf4VffgqaoG/h6cloJxtJSww+olHqLR1MHTqMuLMc/wU3DS1G3ePktC/Dl
NjU0448NwgQ3Ir228Ar/REw2o7BxOqvgEx5s/TgYYcnTxwukZo7LgJc80pw8Pzpp
tXVa6q/FbF7KfvPbaIu4tUuqJpU6EcsEOsZ3Cm6Z+dYJEQkhAgGT44AWAfymwAZC
XibJa3pWddASczsmbn8qm4/PkfgbTAacnnTIxcbrqR6eKn/txtfhkrwBPPLksUil
G6OCkLMAqvjMJLQ8tzjp7rzOOBBitD650ITcUpNsA1xLBy5B3D57FLmdSsQzLuxF
Bn4i97YqrQvs/gnADZilF0KmtIwTx7ztDhVJk6i4uG2qDnmORXuBqj5biR0+l+gn
fKn5N2OjSW4n5ged6tVWw/o/vem1+8TFJNnyoAL7HISYzrjIUdA4eGzcrV/7Mxox
PHtVXuNVMBHiLw4jnkpTS/rjiZfWJFPieH1GPziQ6GltdhHGzkTimzYi8lcfygiG
DhlMVa60+RyRgEVnoMcHA/moud3h+UMf/aEhb0Tx/2PgcikcCG5ECio/KzCPFSgD
wypw1RzIbR6o6LZ7MYDnMq4ycCgdPLq7lzSi9UEzevaAMBNgwr2YtuBhAxzYGY+m
zhMjVBjykITstbrT0yft6cSuFQOqz3GXbT8TBehR2waTuuBsnnHtrkTuduQZy93c
I0aJic03SV9hhDLpf+GQzXZD60Oii8LOMzQyCoCT+sK4m/IqSF9+UtZxShDMoefA
1JW9Zc93J3KwJFWWiwhLc6wSW/3mvUHG2Of7Nx8keIyckzxA7gTb2oR2vIqwNlMk
gubZ4SpRkCkYASWD7inRHEoDn6B2N9IPmtA5nh3e/vs1+ZUuQ80znpGoAi15+n51
YOxUbDoUksGAZu9KYNjZl3tHravMwzNAbk5maFckrin1IzqY8HMVi3xqdqn/je56
Ck4E5NtPe9nlHkGwNvJYxO8/vi4CtkFO+/e68RLgwqB6HNpyezwZFiecqCEKmtzP
B7aG8iiqs8g7XFN9tnQTjhDPsw8I06/ibzg9IiAH5bpva7123+evwet/oMKQb+on
rLJlA8ysFzuJ53t0x/nbgjhPKT2l79LkybLdWD5ayAEOth8KLQBoQlxBEDMvq3KG
6wZTVMxB5Bpm7gMvb58mF/4zVb9JMEB2C84HdYzyDdaNcUPZRtONbNvRtufZ2fO7
AQuEZrPHeKmFQQVPQocDLAE0ZLxFI4t7jbsLwT9bH/QZ2tc/J8yZ5R1/m+JyI5D1
fiDSncFrGtMnEnoHhK9JP/gx4NSF3dxX2rXhHtpWDWom705WdgURk/1z5kppgUBn
B4a4fhFqDFg7aPhJcLM4QS1yEQFY18Uecev/N0S8rJJ9urWS7248cqNHZar4h6T/
2/dWmyKooMfAPvxbjzCsDuoGwMmzGsUz5UuId+2wmuZ0MOfD8zYqY92B647pfySR
Tnzy05WDxtnhIUJmb6PtvrKfvFaM16WrlG82kCEyUM0AcEHpwPDamx4jT6X9KiVW
1pQ/BUPBG4tNM72pp7Ce79QVqNAWDRngLSlsux5PA8u6UY3CBSmBRbZhJtdzD/E7
tUVNUSfDxbCFnCvZ2ll5iQOBpUlu/27nIL95u1FW94zyu4OCFkeJz70kps3j/Fcj
U69UIFO78MriaKLY4calI4ZcyuCfzFEaFJoLyIdE63kpdUfze5YJQRj4Vq+qKF6L
4zDXW7CQJD6xybgy4Zm7aFzwcpgf2Gp6KqPh9V8j5rO87pPjZyvSGW5f95Emb5bb
lgrlo/fTkQ/g08ZISwkoyNQlHv49A2g/bbTzQ9bKhDYXR7hVa+Gl5rKl5K/22Yzt
qUO3URmMIRrRGaTbxRkUG3zq9PnByoWC2WUULVTQgHwYyD/10Aoos+LlbjnuLJsi
ZcqrxDWhqOgupmaJ+9p5Ove4+LcRs0SHNx5QRhTXZ3kwnG5uv4ePIZFi1jCZVl2r
klxpKcUpkvT8o2HNjiOjUlKjAqKnwwZ44gYr9juBNfd2WSprGfbOzi5K+nTFTiFE
OvDU7c2D20FdkGB5RCOjGkXcd0TmTk0uImi+nmhYcFEcuSswqYZOiX2jy0q2x49o
A3VLHknLgubFrPy7+dq4rJPlA0zC2EYJEMphIXhZQ90XzCYvVqT+6zpxNAhw5ZFQ
dmWRgBtChknVu+UH9uzYHOjXkJE0AvpRA0OIKZcLWa+H1MSWVOyR/I5OA+pDXO04
nmrPELwNl9WwWZ4eNezNnZO8t6NZQ017kyVC5PUmbgPVN/12wxQrcBT4BL5WMEyg
IndfeY8YO+CUv+pD/iMyb7UMKy7MUoXcXfgRh7EB7M7d/szqEJiHWQKPFfKrDECh
pafcsyFIKp41j2kPGg85uqS9RKk+g3SYAtWPCBqJSoKHrwABEnF6/IHHYdzwksUI
iOxWXJ0mn59bGQE+X7CxRdIzEWGycP4qrWjfk7u0Vdq4JE8IwVXa3xvTnwApmAUZ
+HhW+j2YeUVF1RbgNYM9vGL/fcDHpQlWp8s0Lvdn4g4apEEXTOOciNKCV+L2QYA/
szzm5gevHbLycpdWuMivVW4kPN1p2XZf5dPYisZz1DM2NZRg8K53MI2XLdI8ehla
cVbMMLA7onc6YA+jFBWsHiRLx0a3/GYCcBc/eY1gJtDnxDh3YQ9XwzqPbKdjvFgC
pDddNZmlQHY3DdTBST7G6lst+uw2ljEoRI6jObPzY+MLHgbxzCdMLfVzFw6ttcpl
fO401mTiHjqaj8o/GQ724Y96Kzb8UXmM6cLy5jys6NjUYVAfDAUU7HfVNy6AjOFn
gZx5v9tlS+KdQPIvhxQmq6By8L3/EGOyTShGz5+w5uVu4LrQXe16iWPXA7mOc5wX
YPD1h4ZwOS6dbg6h/sJ0Q/1gq2p7HsNvRr2Hv8SgLMevK0jr2STHd0/iM8ViOW2s
WWkSnY9Ro2oIE0m+W3KLM9vdQ4zYnaQ0wjpzR4EK5+nUUP/njR8I5Zilp8ZgQAs/
44CjBxD2RB/2cVkRJKeekpsbh7PmofFs8VQYFxI+AQLUxArDlsSQi+OKmo+sffEM
IeJ9je5ZYw689xFIjPPQUh3JgS2VWpQtAWB4MUbFWXcOrKrZuBulmsl11AGEtLYD
el4Pisz05P/mxsSDtqJCILtVvidtZoGyxRMfqMc9D8PhzEL3zXDA4o3vVCN4Qbyg
uJhstW5ir00JVUB7wL0nD1piXKJQ61WEgzsD8WJL0oDACUxhNR5VRAi0ORXdHmk9
dhsvGJ1L1rgZLwLcY8xyD3mtAGmWbzCBwzXboJWaskfysN4Jkhi0HQxOMdSYKnBS
WIoJtF8E0NEmEHOhNqacU2lr285lib7qKo0/DuPChD1tItfT5ABWy10jARs6UHz4
RCQtt2WiIUoPPFmklFFo7hLzi3itXTGd7vesLNm/XUwB6r1TzpiDGopiYCnN0p02
2shIl6L/ut/FPsD/DeQTJ1CYSDfmzRgsEKW2ZGwcA5QiZhz0dyz97Oy7YhorfwuU
8234g+NLoNIAQaTU5QTFIrBGzumrClIvfCGQdXCY4G9wBuRqq6uqKF63TBPoVhTZ
QSyRmnF9dM8i34mt+AKR0Wh8Nz/rXvYB5YdmkHCOOezdYZsinmHSJbgbmiWo/lvg
1lFkPoyanhsIF6tKn1E8GVK5OprilS6d5gXsn72AUyF4xN7f3fwhCZ5g4UI6ujFg
tU2ZIa+xve1lfDGERWPFrpmXmvEIPKr5mFbXScX4qmzUbinDp/bGFzDBCmAxiD2t
bixVYHPXLvoBdfIvAlAvYrbIL3iU2fmafCWt8kmOADv/yoraMPzs265r5iVWSX6k
PsTT7IZXWgG1BB8ritMnr1rGYu/zvFTvXu8WNvwnTdO5w1ISZj7LEZkmwQYPy0RR
deAEcuKR6O3I03+m2pzmt7HFnxWPhC7SuE65TzoCReZo4YP4L0Zu5gtf2Z6fwavz
6ljG6ro5444Iiq2XNLzJZXtxpEL3fSCX00jHopGwuzz/LQC/SrAsRkep5U4+HEg4
i0FLBjB3qAGG0yBU5OMY5VTQdlnjDAxQGTFwTSZMv/ugiVPRLAzLlNqoAMTgphM5
6E5GjbOUnBOQgPGw9OJpKkQUEyLrzSA3jJXdFWNS/KtDSnBf29Gft7n9Zyo7tgVR
KVakiFgVxWcaiLS1lIBUkda11J0ZPhgo/mHJZl8h8+xVFBzZlRRPpTEzgJu4dUl0
w04MOKbWUq++oNS0+Jp/nsuNR5hlQ13C1iPFcGbD/dpdzSEXzlsMRI/MtY9av5LV
5o9zCigiiFD8mZGMp//nirbHF94hJ9MivLOMD9jgLC8NTitg/ct09JweUC7nzWZF
GrZjjMeswHnW0ZQ6U5AoKsSKpApFoBYjrHWdGEH6rXmXDfinetnIeivUVinKpRDi
u3f/RkcMW1XykDYkJT7FJFpRFh7JqqTxQqSnAQpGusZxLuVMUC/eot2JUJFxmy/E
cK40TQaqT+s1DJajtZhYwGCkfE3FAr20QZyZtf5ZnJDOl81wlBHcrGpNa713KC/a
+X3dM8C76bEJg9SemWZdxB4+C3r62aPl0ePe4uIt72fneATXPL4NmlVZXBTthZc8
8SX1fDywtDKX4jwdC1WB20p6ONqa2W7j9TQ6ieqS64QvtzFSkA52yycQfXUm334z
8SvWb1acCEG7u3U72ARfY4q6m6v/hAFGmLiSQE5fwQYthQEOkbsJcCv+zUPI9YKr
OuSJOwBDw2gHOspNHTksq58L/lHgQlFFClWvVOqzVQ12+Bx/ypDLnDfdhaEOPXdG
ZVVo2HCip5qCYYXdefuhqdwXjcScyMLAou7YofmcHKtFZZmJShyl3PcARB2cZ9Iu
3hDNTTzFUtt3EWoKHTfVc/m4174QwsBV/qOo47/AxwR15fbGFMN/vCVoRAANarNu
Ub0wcko4/FyxxZICPHElXm2nzuCu9xEGZGSw+QnsoXdhMmach4SqPyY9fx/YFWdp
KsAPTcU4zEpa+6hzmGS3W9cnR2SDozoQVRXBEA5iTo3hEfnrG9LPO+48Ms8gWBOE
S2spTFK8P+4GOm7/52PGnmB6HjOctjL6XE2OE8lkI7K0fo/zSHDn1hD/6EyMJWW4
QKhtuui7idL9AM5i1lSS4wegs3R3gXx4nOsy7aPmujox4L9vIyDbC+DZk8IQL8gy
bZP+jk7fAZZ9wODDyFtpx2oQJ2JFzTSgrh7CjK9Ra5wq8MurmpLEV1DhpVFH9I4l
kouffsZZkfKQ2DrnUYh1U3BLCi05XEDlbob7S1pEM/K+uvIKSyhAMn2tI1YQMfNE
2cppVj5tyPqIRG6FxO3WwnZI7FbCEZd4OeUqqYpRUTWQ22NS79VR72e8sUW3vEK4
L6Ys7Ua9REFaOrHkvrgoMMZdwbM60ehIJMxJq4q1iv2gDj2ey4CHrv4X2ALDXMC3
zY/21iUcgWz3ylJb550dkgtCgrxfjQM562BRJcNIo3B7LuFEBmVmYEHbz0cb+1Mt
oFT2fUk882lasWem65uQFwplW5HCqrKdywp0H2od5M0+g8akXeaiFHspWBBgf6YM
IoaeAV2eJCEWPeG2j8GvNC4FdKynEVuSfm3tzcyVWvz0DEPOl79M+xcF6PIzDGTQ
vVgE3aWxYPcwcKdmtYmzL9F1932onlea6G79nnfOHTuZyzQJo2ncb1lhTtBv16EH
AUYBWecJ+NstL++6WqfTtJp5eljiLczfqSwX48Y/x3vOhc7JMKIZeKu+FajSe6vR
9GzM/V4ohskf2Kbk8rujt5dyc5ShmnMj1lI11qjyc3Fqiu29lSeGkhx1JTeEZwHt
G0TMvBqxlolD9OYllTUyII4syYtxI4snvWwrI+yh0AaiRZLGei1GTueO2OEDLeSn
zaioNXCpWqZtH3P9tWFMF/ucUt6OKyrQddEP6lzsPYnuyrPMy1mXvXwTHx7l6YwN
cYbQQawhnGOYaJB2ewp4MyMSa5uU+EFa3azIkLXukDyfqy4fSUcfquvSoKQDrCVR
OQ98EW5dXEOxrGylbOjhlbfHcKv32w8mK6/PwEYvybUePovtCVao3sZHs5C0eb7I
dJsWS364A+i6kTSHm+4AezJ/kegQ0/crdjYsmUZE96r9ZCbdwoUrCwQBI8rKop42
LX4RApjbCgC6NfYGV6L4lYjvxBlzDcBaFeuKJC1HeiV+wC4eeLDlg4rxe3LuCjfz
7N75sEigP21oXdZIWtH8A8vK6XXR5I8XfxHixoyLGs9dl8t3r6R7DHDsRNZgfyEi
u+zrkq+aniYYD1RXiUmDRVwqmgMdpJk22nQnRshWA41V+zRNPn1n+aAOcQb4cWCA
zuk8DDBhQVzNxSK99sDzb1T3b1t14IIQwbRaJ19xJSYCBv+oTfp5a4rLMKYbiMzS
PdFxnOPiOyg5eqM+wHFdobszynyTkWV4g9U7pp6nauE45l1ckx8ZPi2o0TM1j+Fm
xnFr10+CX3nvZkg9uVxdQC+96YKHO6ZlhI3NOJefxAlLLVcFqY39bg9lnIvy8nVJ
SCMMWGHEwNr1zzvjh31Gw7dPHz8uKV61OsN+ZKDG1QO3ntDCb/hnPP7WiSixdpF2
4rYJqDcdynj8kLqLxzHj5ZEtvXJ6zjABajR1TPjF3ZrXegeYNgz3loOSJ+wLT61w
nJNsqoOvyOHoRUy6PKudsnEcAcNHLW1bzrTI0zE35vb2Xk+wLvsWuVM3GQLN4ySj
z1kLaAqCAYcvB2f/ldTDJDiqL72NUMV+SrpriJ8RePueSdK4tnNa/h03pUwAITnJ
Do52EaBRvngpd3FoDQww+1Oa/VwFt99R8y6jexchyeAEOpuei90Pa/lSfLadgSNs
/BQDZ6kK8N6UlOEcrQGEshghNSyCNsPflAeXIOBbhkonrNTR5j6SCzf8HyGCBPJc
mufT5gVH7X6o+L6Ml0w8ObOZs5O3xmGTXOtlzLml0kkkeBv9i5gF3oJHBFzXUQ1O
Ay57mERHcNUtMPkvIPyWau6JtClmMrPOG0Re5x61OKPIDwe1VTFEdE3/TaIqh2j5
xgwfY2I6e3CtF9kHTUEhO+hl305gwpKQl5F0l1pKCz3OpGNAIKD2q7UfuYWSIeOj
71tD3vreBUnztxfI2Y+NltL+ki9yVQfScN0m6gY8f7qCMf+9p8t78n9yLwaYra+n
ijbR9ehMwNJaBaITc85VkOft4ylNsjf9NWtKf3JunovGyJYctnUw2829T4ILZx+D
Nr/Q2cBoWPrhTE+EQ4kRNFazYLYMZJ4wAmqlyt/rQgnWPkeUStOeI5FRMf6KaNTc
dTd53h1sTMtTHd+jFiSXYQqZ37A3XqDqgSZMRzrl495QtZwblYv2prqG4JNB/H3n
b6LyLbkngZLuYY4R9bIwOb9LQukYiTtKgWJUz/lakALu4RsloKqWpIoGsV9R6YWK
HRrKoTMkKtNTbJmYzKmaNS08ypsQiJlqM8eAXvR+f2WMv5D0rrh6aXgyh5JQf0NP
vQvGtSWVRnBaLiggsPJOik0wqh8QyEt7wANRolFYqeDfYfV9aFENGL3vbF3vhzIC
Cuyspp5+vb5EgUL9uRqKtknLfIJ2lgltjg9FJrXluNFD0c11OrOsaAM9ZLsRyeBU
S0/h7sjaZON/wzvGMqCxVEqdLgt4Cvout8/7wOJ5xUDjXDHALzOxcHLekvrcl1kA
sfOe354yEjjlLzm0rGbN614TGS+q+de8+JrcSsKLNBtaKZRc3I6AXfu+rpJF9MHz
CulYIPOGFBIIW9P08WNFpDk/LMdIMNHYol0RHs/SZAEcurlHNkBxTPSEAmHHmoxd
pZIHNiN4zNOVgsoUHidpszFEzz66MWMcg2X3OHrAa5y1IQoFV2PX6kU/axI0M+ws
k60qTJeCGKdVMRrYItGaJPIl33enTBi8n0thPylBJFOxdrisvN31ta7kc/GwEDvy
LghYgudZ2kDSXEPELM4rl2qkEUDQJqXfHeMP3z2fPglwlB8xXl5jmozzbfrLau81
bIch8IoREqCYkVEkTva7DOHyw0zbJWdNa0gjyl9x1NYFx/VIARO1b1q/aTGN7Cjf
E3bh5MyJs93MgFdm9j4DQwLiS2qhmoz5liXoatgGppE9R1hjwPhK4sYwJjGfsVrH
qt+jtQnsrj/ZFaUPZP1LLTNU8j7QRhe7oF0CvKOiLHcxNZoLpjf7GcF3WEsBtcGe
ekq4K6Tohiie4EMOJDvNF2bAhzRJ7gHqKkqcHmBLlknAxjoRZssaMMMw+OqOiEQO
QobNzpME8YT5gbWkum2MzOgY7PwVGD2IS8CN10ybITWxRT6WKV8KeEsfmk0K6EiU
I8XuqyPDV8vZRN4yryzC+RK9UzQdO9D5fhLVrK7YZX0PmXL+fI8ESTTwZiZwhcow
r3Y/647d7nVN1oOhHRrDPYF7rFwN67MC3Rlc/mGWUFoL6lJ4Az1ymi38l+5mIS9b
RrBscNAHbWjfb1vB75CSNq6RX73L5Lof32tOAMlBBlEcZYMc1H/T7RPrJpDU4akS
zHBCHT52q0PF9nbqNPmo01gxoZ8Gi2Lmpp7QGue5CtMlK5eymD9SnDUrZhvusHJK
MUTOUE51ST5J6giwMEgr370dWauFcz5Km+3fbdr9UgkZXnpUSZnZovJCSC/YrzIx
IozaA/9w/PzO4lr3QVpGkCmv8CP4oPiFxeigCIptpY2s9GfWzQJx/k3bmE19ySbe
gufvrPxzn7fStKLSrQYGxLKhudXjN8uzNkQNn6esPqCNCMckzm+4PTAGgOr95yrp
D0arRf2JWiIi9xcjQCyieST61BnOtyVg0kS0+uPnT0FZbtC7Yb7Zu7zshiZUlGn1
fpM+8kBFXwpp7rHzO68B1+KxraYx31Z+x3MsMaszKxE4JWcbUDaAmYelYDG2b8oK
MCQ2CmN1miiZkEt1ekXEb/Wkzn1NIkzcl/vkiDjXtCkguJuv705GZUh3iI1s+X6a
4vHyOrmxN2+qFMAZ0cgI+kh8Z83RdHngO5zkI1v8p3kjAKqTUiThxWaGHB1kPOd1
q2M4/XUsrq1wnGffImlLNScHtqcJ8WArMtxfyza18EOMwQ8AYuXZIrwvzcBsQzmZ
8msjiuJMIwBja6ksow44T7VKrdLjew9mavj5r9nNH5oPRGhxrfuVcdPYYFP50LK5
ZEaEsmhe65gPajcQpQ3wOyUblOJtjV6quIoDAucECTdq+rZHbuSGEJH6X08zkFMN
KzRckqJUfcTcVrLmTxCh3ngchfmpwOwNCwZoe/IiSeUmBfp7lng4GKE0Vs3JjMTw
3b00Be9M7tJmGugP+QzaWgBtdywMB1hm1/pbFrEDcIKwO20m2eipE7Ed73gfaNav
s7iNS9VAsjP1wEgJtxizedcvTPMQwwkE2wGQarDHuZE5D9YfOlNpuXsHfNTT7S72
R283ceLC8lYhpofYnPlS0KZj91sXXM0UGlZJ9XckRGM0C3CL5pSC4iy6BYJAo1I4
cNsmlLpnsiI5CqSVKflu0zmCXLv3vu35VGnF8q8rV/lQFaaXOKqNJZFw9uytRDhh
AUtmfrIzyHpwdJ7Con/2JybHFjbuXQE1Kb2TlNPJQuecR4pWuw08WG9JY3O4d4R2
ZE9p3FLTXs978bABmFIpvNCDSvCI8Qt+mMzk+VGP+Ne4+Npy19zogmsv0C5Bv/ze
YabMKq/bGdoihIxEJzEvcz3sK+myZfxyCfXM3QbuTO66U12hcDNU2q2yVJZQMQZt
TVETG1MVzRFAZBb4quhMtimUTSuD4j1WxSOGTQFNyMfeSCDljE0NdlSyOvOh5pW1
6eP8wuexXq2hu5AbxiSu+IUeVV+qllBCC1VBBENj+Bs4paUcOsO2ArsFkdawXRau
Z1zGHIe5HIAZN0aufkca0nOmM+3alaolpEnjeRy51CuTKeUwQlbY6zJb847BanFe
MBkkazzg6ovZcAA8PxCbpghFcr+IJxR9RjCsBDUPBiF2g889USorAFL3UsqlLjKF
ffOpXuuHaHB9RweVxwnF1cIFm0pe5xhemP12oxw32QivmmustF8jcfF409kK2u0j
Nr/PMNOtqavU6bCnJU7ohIPNsMNsqWMHhxxqzCnPugox2vdesusxRHS3mYm6EYX/
+jaM1LnpMf5zomsJAItqvkCYFlu9mS2xE+1azJK+GW8baRQ1bFyQs656tIWy/vBu
+FfnB0QPPNxaPeFjwilKWIENoYc+CScowBv9pEtGH1V1Exqryq2EMnyOjpE4YFiN
PA+AMLHC+TVCeE3YZZpzE4YZIAm1z1EqKXZqfNaSUHPMPL9yPmFycuP1669X+9FO
QGeoV2KAFgRP1fvAbXsQ6438s7qtqeWUmoJz5ieJZo/0Ct1ttqpJBCf37wUMbCGV
XxC3f0P16pHhMPCQf+zbalgDgEwt/0qptKufB0mzZQiA41WlGD/fC5vnBU7v2c6Y
kAnYcQAiMuB73n4shK0xuf8h4dNs7G0BXYk/f3KOy+lSq9HKKbKHHG+FdOxOYuV/
hQAy/dCsZbQP5BRb7ijsQVKIJmTeuGGoWY26HtiFYLKlQBE7XUtMhWRXs3TPA+Jb
cWlY1Y2FfQ0NnAu1bmkr5NlZNXAXH364vTsW/voc/R60jaTZzGIl6vSEzrQpuS3Q
PGd7q8PQRpljKsXYMQqMSnMXjzqOUusg4eEeExkLSdfZkUp+USRh1Prm4LJmlG0K
tib7q8g1J+yutDLzjA7rs14nCPipEGukMj1P2GG+QaNL7JPQpC4qczo3fU0yixL/
l3ZL+Y9mzuLjIUr8CLqkp8aQ2zRlJXKHhtf81h4I4hTcdbslw+Nt+G1et5HD2cP9
Rs9okRJw2lkyZOevZ8rI8a6sxrxUK4+r6TlU6mUXb8n0rga5qj0ltb5XhqDSE4vc
rsJauSOfwje9hPTx+i4oqzeGp2z74x34m8aD29FAAL3LHSyLRhuLIOsTOsW4oGkc
tzwn+DIHHa6H4CbQR/QHq8nJRwZHai2etNm+QpYzX70xIKoPqg3WBCDseVcF/UKb
lfckRopoiwQmBGBw41FPI0q9ziJXGOZ4DjIQsqqvZy09vPnmlNrXEiyqrvRPC5si
ri8PX6tAgapbFAmau78pZA9SlbvDtkXEWNI1wYVBREaX+kqoH1EGoymQ2ytnEOJJ
/+6AOytCfw6BddBiizFZ39vFGrohv6CmVt0xu64Q2/evFhN/wd+vtaq/LRv4H7gJ
NZyra7DsOlZ1g35SI3JsDjm0yEIv9TqXeEMAKOyXY5jmi+qQgWjn22EGQ8gYWCET
qOTUmFH7NQ6qoCkyZrdf3ozj/v0wx4IZgNV2MmVg3qwq8Rqm+5a+KJYJ0ysyoHfL
IAGiAxU+2jgW+eRafJ5pyl3mWGKrMjO9ii2qZzwC3q3p1OdpiYylEROY4iUDgmhM
Y4h36EgSrI34BDfmqHbPdHJncm0zu2uCWqFPZgFhbASBMi7ALp1EDPzYV+EnFJ1d
Jr/X2m5LupTyztz4np3oeMbasPFdvRy38RkRIUfqokLFZyqmVIzGJHDCgVTX+Fsi
M5Sv2dH1fdVeqts5QYg/XJ9eYmyDQKzIpG75SMf/CsFSl1r57eaYhryXrxMMbRf/
MvVgBsgS4NUKPUoLsn0RmyyluEI+QDKHZJ4cQIuNwwBrgRnhdYGrcQWO/8MbCioP
KDikC/SoVEP4Z7v3bdP994WbCeZzk04jbXLRTV4KjO1yUZw0CEPpYGfSnsJc48Zg
H+yJ+9ewRpCRsjcj4ZLHKTo7EgM/DshIUZsb1lDNsljXgUgAF+APSz30UXRDCu62
5a/LxW/Q+yCXlrW4Nv8DLSY8FedQzNWfFkT+kJuRZFuTP8sW+eCWzP9yHlVA9nei
CnrIaGmgCM98zoXPXCfNmnWEYO6A4iLE7YVXdkpX340CyKIJow6hvMGACqwlgYO/
pIxJTRoShgNvE7Koh1bhpiMr5KUe0F8MKg3Duh1jEKysmfMrZ7RfCIXbCOSEx5mQ
ZhsPBbJultBsPeO/2LDwmy2HDZStjmlWTmdRzFhfa3zBG7ZlXqDg2b00uPymlJvl
HN70QzGbSL29CtzDRQzgOYgwVkox/F77ciskhhoa/JMsasaJ5s7GNlUXP9Ahd6A2
QBV7Y1qf1FB0Pq2gaivyhRrrGsMKAgwPIphOwius3NyJxV8SSCs535PQvwAK0Sm9
tTUnaXvDRDshh/tB2yZWu69BQ/L2gUvclzrkLebHO+aoFpbj7cdpUG0nWmmj/enG
7YOQxh8Mg8pR8ze71uPt29G1L0oDliuT8uZDtYcE/ha0w0cp8dycNRev9Qs0WiuZ
eCicVYVEH99knVk78GoU2X8sHI8er0FJt/xSZHehnWn37xb7zUOviIbjJE/9r7na
V64B/YfCDHFa3qWShsaIfpEFOGDCVpF8zIH7L1u7RjL5VVnvIdM8wqTi1yS3Vlx5
0Z8YFgNmCV4Z4bTXkdF3yS4/KNywhQu6f6AY5pjd7aByeCj+BTfBFD2wn9/WHXYV
5SDiRJm82KIAnOVa03lq687ZXjAxDVt00CCDebl6gV+Ag9IbUONLnm50OgujB7HI
kXe28OCssaJ76/jOYcvmb9wxZG2EIIuUoRL3mmbECR6fmwbZOq1DN7f9RUXAzVWs
7pK7sSKVGns5UOUbU8UUavygS/F1c6lAkJyg3Y7lERGRMfxmHBWkTuZqwRmvmvYF
XWc6gjb7TEzfQKG6jB8Dli6mFW7bb8BkkaWYiCxroD64Yntxi5fmE/p1JAUmwvXf
BEq4xx4PVub0ChkZm36EpMV9XT6CKw1eKM7tMgxQgXSe1Ps0LknQPP9vF12cl3Pm
Qni+M/UyHr2st5oBNK8VRMU2ITeH0Os1wA5OYyXSTm6JYoQ4m90N+6ZxSkTo4FGE
o84mG9A4/SCZgiaQmPsSXxql7KcLz0iqqjOJ2lYHM1tabBmGmdOxtAYSZ2xVrilK
VEhcLMaA+zDdsc/Zh5pxCAtCdO8cP1pGyLxV/rClklOBv487k8yZdfkBl7oRYgKu
v7JBsDQ7Gh2x2XV6ZQCZDDgb+a8AThHtzPfkMDFrq44k5fO/w1Rouae08naigm3Z
Z7np3XmJ47ReNMVyzaEMX83qMqN2Ylc6cg2HH/X0K73hgXff4iZmOEUNi3FWndLo
PosVVoKP3+xbS1msi3t03Lkn2qtpD7krSdPQceR/HyuJjkhNlTkJ6p4wTloZUf/W
EXCQ9lMbZuwoJ5Jwu/mvuoXu7vV8mbmkIRi56xWwa+812P3pF04LNdUC0mWp2hkN
kg0ZQQFvAurKI2D7BECOwPlZ2To31tBqTC0l65tC0Q1Vf8fSK22nmHOfIAlV7ymq
p+jJbdvEF60dw711MtLtuAWslUQFXJwJ2RiY7hU7IZSgd3Gm4px35HFL7+sq4ddW
CH+3/cg9yRnM6VtnCZ8PxtrCso0BpHSkHA2H+Xv2lYKqPJDZpy0zf8FQ76oruuaF
rrWgxrDV+68QYiv2DtETIfoHtil+IWEVZ+4fkQ1YmFnLSTMZcKzH+N5DsdO6PMKT
qLQwj65vrDw1Usabo1pPSGhBoeZVDiP5zrVLuzsDmiasdgSKFrum72SeFJaxuAjE
7k4yPI1uxnkVVkWNTp39DpaWOER+E0iTxBxBLQCcf4KOOS37xrwJya1SJIphJG7J
Xu9ogAXqwWmmFu8B6q48C/ADS5pK3sLnddhg7gM4ml3mYUUpPgLF/XiclU9IfdZq
+05lYgN1MTKQlhWW84OVqpUMX7lKBsKRNKTgLRvimn2KArM5lKVOcoRdPQvjMZe3
8JoZj9dWbNZ1CYbqivKTJHg7yMuSV3LjoGFYbvzi8PUzx/hDhroEDL/Q9/ZTyb2e
MQAId7jvvzdwlkOWTuGKTkmoyqNVkKDj/0hjW2fVYChdwVAwqJMGKosHsigo0umN
XQv2UGXEPe1maoN7E+gJC7ok4PxhWVaf5RmiW25wWu3Uz4Tb+iU7yLtOUgWEr+36
daU3f/ycDzrQgKMk6rxFVsDcZC8Gt+b+dasPoCsEANbV0tEtutJkade53JlLjpQl
emoIo5nHE2Ro8RxDA5YjP9S65sxlI8sfQ+6iSJwtYig6Wjx0XIOdNqu/ziP3K9Gu
DHONUUH8sCSNjI7adLqqMpOjwEqTG3yPY4PxMtN3LxQ0AVCo7s4SVZJwYdNqGPFY
306MnXNOKFLuVqRwUVAsJHcERMk53YyYksIxyJWGVA9aTCKV/lXs0TxYqnIF8Sgq
5pwwzj3GpQTTDenhThteG4fBylDHDQUoCq9iPY4s8zu5bk4aHT5l42oBa0yR4rgO
1OfBbio4z7Xqt2C9k5i8Hz/AGToH7WL0IrSPWr4XRjtPK353QoW2TpIjT4okzqRj
gi9W646gE4EZLDfipHP1TiY0Pz5+AHUPp4Bd99xAzvd3PH8Y+Qe8FnQhulrFlTX6
3SMwhGafOOHTyv9oubNYIjBM4hEBVgCBreva7Y7S5dPXFkGG4Xe/pJDMCnscFmh6
CPHSYV+RCTTszSYPJhPRzP9D9svw6Fq26cFawW+W4utf1DQ5StLAyCqBHt2LklaY
CWSeFB9T6D3Ogfh45HWp4j498sSa6kyBFqyFn9HyKfgzEWOB3Us211R2MB/Zx1yz
sUOHwByC3p1DT3VuMa1vLYZRBi8TV+ZTCIRvDNMEEMEhLAkhHDrFKUdvKbVExRgp
OkdLPLGFNbj/Tk3p5PWpCmLaeUEK2jhEE7jBG88kOeGEwBbkw/uAuyE7yNhDLzN7
EMsOxEjONfbzBQQpOzHHWcsKd14T4VEtISv2kNo0lv43KvzOFI3NJ8gWXNjr4cJr
J4IWRd7GxYJiqo3RjdqXqfpwdpo+6+A61O1sk8KDBMIKFmKQRLKPo81OdUko0rbt
0CvrcmmmA5uSKsy0DA0GBgMmV3i6Bt/6UVe+m+EknMeqm1C6yfQn3/JogiUelkAY
0SmMxrVWP39A/iZAY8jql63zDuOLOVuIn+NixlzmSxpNuTjxgeMEmUxXgZOt6dwu
JMm8893n6kYsaeg9JXHLfW3lKIQ1A7SyfF6z3T3bgQgN7JrC/0HZjYnBBh7J8iyK
CUFQz+HtZSCetnZbCbB+zkP7Qf6Gr2/QG60RAxihKjE0Erc3QU8w8Cx6pj+kiw6D
0/RgR1J8DwbiQMHDYKFCRaqpc2YUHyn9rP0M5iEz/0EFyF6pWbTMy1fDbp4IDgvG
yxVDd/rDl2NXkEo+/abqu/s+Aaw3e5aACGlmiT0/pqs+/x/lzgUsligfGe4tnddt
AV8ZYqlANzA2hH+vanfnyl5AD47WBOd9VcdujerV+MB6LkCDfaAUkvIdC9TAwy6D
YSJ4yKZ2POtijUaA5IuP00NMkqXAIU8vM4brXO4A3GKaItrMa4xNsqh4TC7pZHMf
Oc3cD1adPiVYM83Ovp0cKOpVgNgwN+R4vNihN4vkcSJiQh+vti0AGtWIB6pkcnNs
1sGCQr0sYTyIBJZCal8wOfZXo78b0hvwmNZwe3x/wU0zLrkgg+Abb7058VIbTCJV
QSINkvft63QOQbFTYbKHg/YHE1j035fZHWfqy0LKkAGeVk5/2ibibd5HMFBYhOP/
e8V63poQazwonbNbzgKAfgfSTB1jPSZrIPWlI6wze+1Z9nf0G2EYk+HLXRS5zAPH
H8mKocGvvrSChzMOC7ergemmxMxpteYU9pjkndkHpyU0D8jmQcbbeRNZr7LsA7GO
gtxVYwKKDqli0JHyNQLjODs/68kjd+i7K5oDN42flqJzYbNmK5koZb310OzouOqn
aqRjgQ81Ag3+geFpJh9LcTz6GQn1RKiBvOZhkwtmKN5t5Z9a83mRbg0HzoFoufoX
T3UfDUCow2M2T2+hZ/7T80yfcJV+5ZtzJVl2b7/kehh9hRhx+sGtFbsdzCnwBGus
PgS1j/qnhqboK1JizIpcBaMeMRPNLqXQ2C50RwcqU7zbnILfTTCkJ+/K3IW9/E9i
68sngIJFJkNRTS7Zsrok+Vk8Jq8BzEHtPKKWWVZ9Yhb4v4vVtIeyzpVJHo2TNz3/
z3XocnEfv+ESIZwAE1jsoCFnRzUn1U5x7oqtgBxtVvfIRycs0izW3fau5KTVPCAd
6Fd6KvQ+9fJ10DlvA5cqjtC0f54evzfvME9xi2UadYqDhowa7RWXLNrNlam/vao/
Je+XeaeQ6rv9QrqHFHUDuRlEGXckylCL1hXYh3NCRieyvEgB3+vw9irNYf1iWMO0
JLKW1hagFUsMaQ+q4ECT77K6GvH2fDaAU6LhHYGoDY+krxxhcadQPCRnl7/qJFih
FgwJf+U9TSroM69ncHkNlZPPHctcFgcaEfPRErYPtPIZ3l9R/90MFB/xu77C4VP5
sNl9LH7MCa1TFErYd9C/qGHIOPlZlPG3F7UrCl9m0RSB8ThNSTMoUH4ujKSEIiGN
4usFA9qdkuSvaTisu7+T+LAeuzV4ALn4UpqFnpBv6iQEE7aPZmJzj/38pQKq8jDf
iE9gZhhikY5iEqrMWZcp6K6XmOfy2/Dsoc+lTl3szHLn7aJ4O897fozSBNtsm4dk
bmHBhhxjawJJF2RpAprQRHS6VG2bE4iZOQMMGhy8cYkGud1k8xV6KiTX5uOFJhAw
T4Po8Rvq73BVkQdILEn3XQYS9xMTGYcphKs9ziE5I9ed9NbbyR0v4TUL+WwRIVvR
nD2DbEpPI71wx09EadXokx1hukWtf8W9fgQs4EDH+g+5hLje0jop06qogZswFUG2
wMEcuW2/Sv9vjkivHorysn9Q3IwF+Ov6++ObAXQWVtuWU0eXasyg59uEY0KoYgVf
WNJSt313HYGhxUub+qD3XbG7qQHN2mz2aTUDeWSM7kwj2FGqj/cjmsS9MCBM2t5m
46Xz7PHcOyXig/MMEES5cqa+8pZDSIP3GBrkZW4Leqk3MxqtVCDVJWxf6IHNYZxu
hSnmbVPGhNv6KyNaQnl7RMqS8yYroZTFh6Ta4VplP7nUBDS5Nwk00bLZ6HLtw81o
z6YWJSCi3tfTPzu2LQNSNOn1ZzmH8O1MK5AT41+yWjFR89CO+KZiziYo3x8GERZB
jGlpF0a2l4UcMrP3kPTcKwgwAmAO8U4rWH8lPYnZ8CyyOiXxDt3Gw35xj77Q9Hww
y4VyagkxNQryKqevKP9Ot/AljLY69VbaGEhvNui36p5n+18UL0waTAy7/EPindvp
R83SByYpmQtA2+JXXx+CwSW9hwNhckEUNDBd8/Z6gWJZ+KcT3icRnVieBBQhZd4N
+/uivlcT8OxHzSE5Fn4X9vlj0OdAuFdxJyDYy6X4VY3sCsKWgf5MkLLcYXBLNjCB
xMksItSfMFi2abiZLiBbXJ6+eFd7kCnXdNVPci61/ro4heMFQN0BclnHiJauUwkd
1gW4F98vfzO4TK+FMkxgaupTz6Rr4KAnk21ADUI7/j0CtXhUjIUuo7v67MjP3e1x
b2Q9HmtaEyAIjyL5Z8Uxv+XvjQuvohxAYY/XXl4IEml0f3dWDfkkK0cHxAvFLEkK
ZFWjHPfMKiyw1HXv5L40+BZ1a7eBHbHRy7nWtp/XY+jEQ1utDfRIHT8dNKnUYVF5
3FDBKmGAMbywXhS9CdALCAhqCLIl1IKAG3iqzIwJOeurhA2KosJ1ZcbFtSX0mCgg
EOyvA9YarrE/JD2hb9zT7zTZOyqaQBS530yQ/S6+ksFZG27Ow2eSjAQdYgrHamwe
qDK3+ojczJc8uGIyIpt2UYJd0sm7HdS8xWEheKEmGi9pDU+GallTNahKWpavCHbW
ygc1ZXihLABM0CgAU8PIRRRCIfsJAYLyt4/Q4BN/jvVqY9nDcbHKQhmF8vD6yo4F
c4ek/6Quf88EZIgCce7a9AderRHZu5rSdkwiGYx0jH+GWgFOPsy2dSW23iYVZS3J
UQa6R6jG8NV/2aah00cOaBMPjKP8JFepDIGZIoaG53DuLatr74HBqMGaP/Mw9Ntf
NQYOTWi0iPixZaNtQi4VeMHlRHSnbTYd1nk86CbDG9ZVgqASkM8iBO6sYWBwU3ng
4ZcXP7fI3VEzSCPcVO+tVwLsLuaxc3mZK1yqqToig4EFArZTN6AKm0JX1LWHrpcs
Ls3jrkFlIPeyLjB+gqgC3dBWiwlcOPWBxaBNmI1Gqh7OX20Ur3xqOOlKT1QwkHpW
mGGOOXuLU0+MEf9AHLxT4A3t85JtemG15bZ/ojvhfjw/lFmi/HqjDRJeexYzLAjT
W4WVOcepPSkij0rFNlOJKKFB5Ew0rUMv8x6hhBKtcUY3mb5/3NBySZs4T42bBCL7
cLOaYQQkKXBUb0AhvPZ4jhATGgSqFF5wL43vqUu5IDfZb0OiMTy4+gaJRUrOkBqG
pz9cXvvh8pmRa9U797ykCdONoGspGpM7jSSeRJPBwIA/hXg0Q6wzuTwymMijRV6Y
ESdc6e/nbag+KLnTrMh5Cl4W6tCRmbIqAxL6fRuuJEVabAWtfB2C7nN7mfbN0Zq3
12VvGyeAI49a0D7tu7r7oHsdgyRqDQI53NMQR0hmJQ//IhWVpdNFX3NuaLbXJxmp
yVPkBgq3ZxNR01b1ruIh8dDC5d6tqpTq26yZm4Xpdhor4WPC346RVJrVPgdKZSdI
jDswp7PlWJ4ijZP7t8QisRKFBiRY4DedlWDf1Uqj2z5yBueEf+G78zLmBIalFqVd
nJzAgWa9pKlkB1UyItJmN+xPzW5xX5lJ9aH+UqW9oKxdbXq5DICi0qK4hfF6o+GP
RX0hftpfoz1ToVnXR2xTF02D6bZtK6VkjOqoxx1eUDeq1Gofw1X39oGZ1QiuJ7AC
bkU9Ji5cvGU1tHDNTNrU7iV/dxJvz7KuZWpQoFqvXzZHSYGsDNB7CTJvFkAPj4YL
ToTDvLbZstI5+QD6RFHOWl2TVkHW+nAx960gGX94IUbwTksWVI5Ae1kCy3ibQzeT
V0l8eL+KKD3bgGch+RY5tTZnzLOotJpfz4pHugQir1lrL2EYSjkVWagtJFeHXAnc
nmQetx6dPtW9mujeO2mYD7VA+Jymrqll3QZHXnjTmyDLYciIQk8eGH02cpX4v2Y5
8vm6qX7wf9rCLin2+P2QgQCjGpeDElSaiVrBoDJmasXinQGgYcqU8lH86xtziRUB
6h509yCBlEvzBw0ec9VY24YCNGZXSTnavHZ6TRN1+PCbOY4DWVxRgs9MAgnH7wOp
KTyUVLGdlaesJhOzy+S3r9Fhgw6SnhLYfdcC7fJasuSedi3S8qe7MYmfGL8HSYYG
GyPq/Ontcd5qlWZQfLU+PTf+m3Zhac/iqb232/KrjMelf6e1DB+miNh+WMdQkzRw
O4I3QOl38j1/bXy+H3f+F08B1/8YAPi82FRUv8FUQFezB5aiii7Ltg4e/HhW+XC6
KlG6S8JxaxFPCE2v+EKftTvW3Abz2L+LrhwsmYPncR+Nmds8XV3fhCXtvJMjmsSh
fWZ+B+HLoQEyU27y2Yf19saHTu9wfQxxX2R+Q5I91l7/YE9yKW/8GQNoM357/+JE
egJE9LjUq7ziE9Tu0NW6nZ2NA7HaSdp+y7K6cuJEGBwc5LuLngRmazWJrXT7UueW
s98Sn6hq/ssxHrHme2RLpMKV2k1mGJoCjY6nJnpOPOz2Ro/v+C1kTc7W2t+yeYR4
JHhVvjiijkAIs9tnJbzWD1ZCSECUgg8Yid7gkQL1U+XJW7S7zqqM0yIrrr+fhxE9
jTrrBwWtCHVKH0SiZ4HrCsr9K46xnHLFOzfs7ah3w1Jiv9kMuriAuTNy2KiP8hpI
OMSdBzPfQ9El3hjNTSFkIPhUo9jQHS/JToADTz9xX62CMQoOu861wIDRgklB77da
qhQmf6l3lc4e3D2lzZx9ylQeAVj/1hVcDFaJRZq2SeYB09C+clK2/9Wv+xMGLUgI
qgRJrkDZRcThSu56lDi/C026Uv65gqBEoQ6KtZmw1g9I3XJC06Tl5KyIQBF5vv3V
81Rzp4cHCd+L2HcKqeXwx5AJMA11VU8YEC1USlXJhOFg/1rRj2lTho1hUE7AdXtC
U6mBWebQf0Xjyg7YTQUpjatB2iMufkMfD8eY5p8BrBIOrIggk2uySaykYlqAidYh
PKzDyu9acR+N1Ktd7iqhL2lcRWGyRvfS/davNhPASDdr6ut7eZ2C2t/XMZYUVyyA
9ibYl0rL2jXs7cKdY2s5L0EFIpygisw7tj/XwAx3QDT8uaRdriudHExc9BQIFfaU
2b4GppbUzsAYPEfea97/nc7GhTvyOH4wJLKG2BsFYRtCeT30VqoenR/aMDiLou9u
5RYZwFNyz4JoxRVKNkaf1hpvvXFSy8fuU4EpPOc3MBMi9lX9ke/YK+lZndT9w7mg
kxiB9OlvqDt1A3H5VDOSYX4SRpmk6EsbqXIfLiVZtS/g+SloFYSHqN+dSb+lbmyB
5dVS2PjhJX0a9OYQ2XuHiNTFZGpHobq+51v15AqdSWD30InkQoIQgY8QgjaewkOO
iWaF235WNQPokocczZGMwxwlI5XL/oq52rwPeRB+2/mKeRb3urTJ9INzHviYX+uh
rX6MJKcnzFTQzYW6wg1IoFK9xHnHttlvTycU0/3er22pmPfJzWY3XNz6HVuKZkRr
rFGxLDF8PfD0TOvRtfGcrCPpJi7vv8VdbkujO1nxZH5kJtjTONp0cbqhAUToNsYK
yvmp8tGZ+X1qCB3yeFYqQCBSiNv/ApzAZUySs047mW0ME5OS3iKf39mZmwLkVe6F
SxhyodSSxdTTaInbKJg6Vyq8DBwwBNi7OfLxYG98Joz6B1NDoOSKx868str3hu6p
PVkYkF7uY40DENCJovSwQ3WCgxGtrvyuJYjDG//SdazdDU4n31tLg0RVecJOx39B
YhNN2HK5D9vl7izHtSXtbJQ+kG6gHsKSagR6hl+cmVBxH1i/xjMsTrfNL9QjTob0
hi1TuJHC48Z3yN/oZyXhM2qY/ifCxBe40CYoYnVDIGLDpmyB0TdZRnGvxROGBb+r
fczE+89ktDukPrRHhXvn2V0f9snMhPPaepQfgKTNwSck/DCDwd7VUr+kqgR7MqZ0
Vn3YIrn8XlysXl/XdKMWIjWeDTdjwaX/lNywskf7DK1HCvudV6b9afjW42fXLqxR
lwbS6sFB1jWEW685hjgVg+J4AmlTK0WjhuUc77vPY74Cx7g5GmxEVb2nXDeNZLpo
OSVlHq1ePV2MCxvfvvshhdElMn6QOpsTdqhUAU5gcFyjC7pdEP64nJ8MteAb0NyC
GN+lm4VOWwr0eHsa5m0INO/RHtsoXmMQ+mOOws2vhWQA7Ql/Ywo7vjes+xHOM62j
TYPB2+/mA76uPqFyeam64GTlg8PNUTxLp8AauCudd1WM6F1b0y14xAGDswGP6y+r
i4vrkw4w3kffNZrQyvN2B7butNfl+g3JScXqwu/ZboTsQOf6AM+NZ9z3rpCa0D7e
hoEw2vBKm2scTJmGqed+ZtksA7ny0XBQFzEY18RcRPMeK7LJpOiEqRB9fFugURsU
pZvfRozHDEUhOyGIBB4rZyfuQbpV5AtUoBPmk1Tc5Jrwbw9pc7Vxu1QF55+vfODI
RFd5KlVg+OPsqRz85vT4CNFR06TPvKCy5ttR1JOayjowVuLhvW4kW6cmw+rwB5lM
ssyoEXHkTcudaYVIfInpJpcwwhOwUFalhHVNTzMYIGEtrxzzPQzGp0Qa1CvrYTAO
dXzmlJDePXN7+Cx2QIuqVSPsbYggUhy/ucbP8pkqEVfRc/R64Ku9zoSl/W1hIZSd
tro1LvTi94jop905hUO38HKdUsX+Hp9JBCycO123+j/h0HzE1o+ePMTNcraQwQtY
KgdlsZKb3KfpoUfWSwXTfeYi1gdxEYa/8abTeSXLYv9FhkYlGJ7qOjCUiimZuuJ1
Bf64rzD1IfKpezmQUggUwLW2c3m33qrlBiSK+MKruBWnBjg2Zn2tHDWdoTO7h11z
LFhOnM2stvdmmoO8lJhIHQFgrrFw0pxDabf51V16c7kK7p6YrL6xvK1TLC0mKd7R
KjEHvRJxlociNsfbaCxsz68J1YwFK0xOJ+5SRtgCaQpudf6VH0DffVPGB4QDgjr+
3QWriqecH0KAwZtUiAkdSVisTbV9oZQyBOYGD2gK58xfeAX59+p1rKAVqRXYIpHm
oz/uVGvWfr3qzP9oltOqoWHNeiCTvqD1gmmr6oZL5r+6vPv07weV7ztFRS+7QvBn
YGw4ZZQIyu4xYV7hXxun9IabVI3ZoaMTR1/njxDFx/1NCd4m/0S+xIBb74iW/kc8
RK+u8JyrYbk1V5XZpRYm+DbQwZcAia2KLwhWJRZ6HUSD/2PrtdGaVrqJUn3z8UBa
VWOGXDGJ00xXlTJRX5nLljlmE6JzU2ZudK8cl5v8Sfpxqqr3iF6koBwYorGQcSlE
9WSe7djF7aIUCiYCJh5fjtdLJGi7P0CF+2Fwqi03FBWs4hY7uTPw3oFbKIMS7ne/
arlkCk/+gh3Un2qqLezisfME29UUS5Qd4brCgXnE2x8MK2tpkyOCa7i81dXvAdto
Kt8sLjcK5Ta3ob0cwNW7fpPI1ye6b1Sh4JOUUnkVdWS04uIG3XYSb00VhF7D9tpF
XBYocemlN5miJIUV4TTUaDixdUXzukHouhKkRFAi4jVWKp8htXz+C+5gXyNZSkrL
hwWziq0d8qtpVW7Ha02/s13oMEo0VFJ/EtcYc/hkywB7yuqxTtidd8QN8GyDx18K
36mbMEDwolnOBJCrQUlCX+GjqctSNIsd1xN4NpOzxUYyTnwTYlaR0EBWH0/VxlQ0
+h4myTrGOToA2c94iEGG25gWRceyanNN+lc3fvcTx4fMe4ro44PzfCefnSc9dlEM
Pgp3KY6UHPeiIdJ8ZzCLTmqH5Rgr6LDrBE0bDNPTpcJfG2iY5QeDg5NuEXOvnYsZ
mpLQ/Y0+zidVRwgRyblaLmr50zdqTEjJ3nkzhE11qVQmJhrtC5VoO1WXl2TxazyV
bwR6e4uC1qqa4gFRg8xnQp8zp5Gbht/0QqWAgloIPbNmuk57FmaHL3pBhNNFGDRZ
FgtyWz1Rktijov2eBnH4d48tVh+wEBlAzAXCyhtgsV7lbifTj2t4RNwNsN+Pnzyc
kDNKIO1YHHR+TUQXE3LV3NAiIWiSQKyiA6h/1+sqc+M/LoZCePhOcgwOftNuvCxp
FdgnBr1DYCHECzDTY6Y+/Yj11xZNfZNm6Rlz/bJZKOdXIyTtbUiCt5OQbTKK3xYz
AjSerkovgzkuDXBKWgKIn+opRYHeT7F4b/0R6t2a+/kx7yC3hC3lrg15B0SDGogL
hU+OdstOgLhBTAQdiVLPwUAcSMrB/Ia1OoDgaTnRIMohVtjo+gMNnXVv/X38urYC
JLxK3w+MKgXbZGTaPsg94FPH7i6TVbcCoo7HfVtS2F1XH/GAjg8h3PpwBeDoXqfh
N+WWhb9Jd0YTC0G9w6p7MbWYUksrdpG2FGzI4AHHkD6RjMZ6+o6QXg8cS+2rb3z8
x2eCKLML9EVRN98gRFy+OvGmu+b52m6d9imI/jSrYfwYib7AwMx/IXEh1Zzgsnt1
S0LKoyL8WcpBJxBmo8T3glZvNkexgviEXUmdSSkUHMbGSfULfI05HxlgEesxRJq/
XyryAilt/b5R7T95m1i3wtgUe2uPYMvIKjchAXFPdvJVIY7+qTuGp9m5VqypLVR9
9PCdNjgdfhieSoIxhU6Rk15NdUpWSv0iRQCBV/hhz4gf3+Q9boOB5kRl2jyvOMrR
dQe3A88LxLsFPJNbOQSQ788nJSWlv/BmXycVVILubcmvhdkGRatOoet0O7l8057J
pP8IblkFLcs3HUCmbNbccfljdsDEIaqnZX9qrC5cnBcaS3Mr+ZhsO3tJwqtnV0xU
ijCsPfgxhP/ODEebPWNJi/597hMHPDpyifH5JZqMj9LK96miJXiC7XjZWsRSSSrm
yQvXImkLSuBj5+q/tOVnivb6ShIInVI1NVveFSendYIQR+EYIyg3/2SI5MycG3Vc
Y6h7ZKLrhef0ymnqW7OArUW2O7VOgn3LzaNn5vCyXpnHWXB6ZoTBb4H7BLbTbm7w
epKk0lQnfWY6aZNKjkYy//vtyvG7m6+0UL+CTPMm0a/+Hrj+CUhEDvBEG2sSo3m/
phRXajy4p181qs3GjEC+fPQVhyIxl4FqOA32LxNo4w7SecYqe8v3Gu4FbnSVwv6I
iDzbXi+gLJM/85jod/hO142VnYNQmMyqKWwlDf3U/Qm9hMo7zGtUVb0NAI6NMByX
gZS83z6JnnphCTSNwAtRDzs8sAalOB+NIYfqYXeEeh+f1mNq8fifIR4njbqjnST3
GNcswTPZITbbQK2vogmmfOAYNZVP05cFAqKTwzdeX0IhBzdfu+h4GEMsYKJxgE7Y
gLjTYwzxzCrTzi/J2uelbndTT3+I7ThHaDSxWvSnnggKAAA9S6l6fX8G68gCVFOG
Nyr6ofJA/Z0monDoy/c+SxYOGvCu4qALFx+5EHwQldtzZfMjD12UYIxymeV72zPY
JrzkMFq72Evx05WLkBN+aRbA7qrTRkPKEsLUwx61mjGIR8FUQ2zuy6wepVyeEvHb
F4UP3JVAvZN+DBJAfSJ8RIs/r7UjP5Y4imtH2x+pOrVz/Jxn8uAtaTaZbcxCFlmW
ekoTllV0SxWi5mygn0j+UNLVeBLsQR3hjnyqaQ74cxEBM2uh5ckp7Jxy2D7lM2jg
LYE0fMNDwfKtBV6Sq+xkkOHLo0VdVq9BVF1vWvdOPIz1YqkMSp4wND7RASDRxG2g
E0qYLygPXc6bxxf2EU3OV164J7+YpzsMwnjpF7ye6aTjpaWInaufXrtws1c8qInP
n0GpAlVuWMQ+MtoPI+PyAwvV72eMDM1FrzaocB5Vg4Pfj7G87TSaH3ACHm9veCbf
yh3Gy2miWfPfOxsUnt318KAwE4glD9IVf7f6z0LKI9BixiQ9zl+NvWyIxjYvBYNA
vMrA/gXUOstNIp6Y/cBp/n3649hbFHunK++oFqHPwRn/aOhIzPK0G6XyOCkH55YP
CO/rD7SmYPOf333BrdV+Wqsy3/IBxfxrSrDHPP/z96AxGTFL5QfKgRZGFubGVNJl
WT7WZfglw3nq9A6BKmER6mE/G7TPtCuyZ2GxTPv7bwxpZou+yIYuvQT58vdb3YCc
5QJzOp5n/GiKi5TETV6KQi2ePWVURAhI7819WmbixTfY2bEp1Vkhh3Rb4Q1RzcPZ
6uvUDpb8HXPLGNoeW9fS3BOjQHvCDlaoyb/Nt3FiAef8JMxPlITJfraXWOwGE/xx
SXpMKAWcIhXzxHkwq/45NzBo9xxYsuoD1kzVNyCQ7RK9Sd94nnoZKtWOClryDj01
rT8Xmh65FrwcR3L2mw502qpUuu5XycOTlyAYIMobIIgxS5oI1C406mZSypkf74r7
QaIBW3UewM45z6UZV7DgRrb2yGYQ9HdWJEzhUY134XUlvajMc08UQeNavKk3jKHP
WRzUqmrPBlXtyaVuRBjMJGR/P6f6qsg7RayhNwbU9hWbGaRe3spjuywPDPGnmzwL
yg01ZMgnL3cBeHTOq/VJCz04McctvNR7bxU2+95F8rBpMhUuKnhRRRNrjdoyL0jK
21Vu+aAigyIsGhYmtZmrNnb2RuCs5rT0B7LTo4V0IqztlUarLDFC255TGir3fZSR
TM8se7R95ieoYQJXMFd6EpX5DhKmuwp5fzwe0ESOSIs8OfNQB6tkKP98/Lq/97Gg
2Xpr4/qhQsl7oW/qtXFFz3WboYqrnEXBKqREgyq/Wkna8PGe+eOqYwvfEqd3lsYh
C1MxmM+OmX3E+lYNYmpf/aKc/bA2TRWYdMyQNy5JZfwHqvfFzs8h8um11VEAs3KC
WiZG26VsuvgAKJq5gARhBORXTfz6RmINsaYocDlsc2gmxDmabu/ciRuNH7LGxCC+
KpWjmwk6Lbc2vmFjJgCh5/xdEzXv0tk2Gw4gORMMKoi+jnsRkgAiSxFGhyeODYF5
vnXhz+HhHStg1ZHsUWZq+w1ZiUPwTBAF08T4qsHpUQFXC8ZqFOfrhKpNrNnDKRkF
rgJJK6k+cI8QKMb8TcKv+SawLJhwD6WbfH8aRy2qNwg+0Bq0Q2+4p7kO+I5IP6Gv
botCnI5KSGkPESGkV3vGvLpTRLoTrE9ABaiTtyEW3XalF7jT/3x9i2q8SL48BZRj
t5M2RBPHEezD4uxV6HH3ST0Sm/RO9ZOzTuslnWsmMftexxj2vDA4YfWx/NmkoAnc
LVYSA24iFpk4N+SpBBnO4cL+dGJxJco248590pfKU/nCdNVGXxzNwtMVqMK6Ky5V
hT24Zf9NJsSsV8Sut5ikdz3P3X4JWyrSZnJqw4LER+p3xyG+Q2OZnROmh7V2aG4G
zbfHkGXDzm20t93Qn512WdQ0DWqZsgX9ng8M9fHSVKsj/opYyUnj3uKa3h63Ozp7
/vJhmqDiaD/mrdIx27zP91WcYJUmsfssZCmm5klxjmIHi3iiDcA8jPpprLvRNxIc
VLyJRq2WVX1H2YOp8Zowm9hy9rfHpSqyx6CNTP20flLbIR4Cjvzu6S3cmWve+yQI
kollz0Lr1uDL02DkI+H8gzlGpVlp1xxx82TUyaDa8Vr1ElTaEQMGw0g4LuKKJHfy
dfd0Uc+B4f/UiX9FRTqIvGwJUWIgi1qGQu7ZuEAOmbw9EDzXjSYaTKcKGDxEmmoV
Y6tMs6lsliewR8bIHyD7TDoy6XhL3Av5wMB2B060asIaM6e2HkxYjjd7wB3g/R6C
xkUj779T/3+6yznv5RjkETUQWv1c/3fcWI7jDBAb5BFGQbxHVZRoJ2g9LKxjB38a
tuURD+ZzKvosXLQU9RSz4r5o0090e/RA4tW8IBt2TPEsCdZQ4/VIzlQSfyWZiN8r
aN9boxUg9NDSVfcOxg5erVeHlxcKna4Erg1d0pSpsuzYLCeywWnMh6IxG+EHCu4X
CsW57Scg9sROpjFHPvACO62mn/ys7qO9P1EJJSqH1JtNarWZQo5MsHAuEoYPJCZk
fC24cqRktsOzPGwoLKGHZUNLe2Y4AC0N/ONk9hGUqSEYumlbK222XfIkdoDhFs9Q
KWyPisBViEZu9HtkBXGzYvwaRVo49DA+19l8u9UhXPFThc9kzpaNoqWIGSvg9kPu
06KXlzyE1OuPUIO8ZmhSbuejLeuSQtI0+iaGTlsocWELSNAUPC7vSgzijy9QNzVv
hhbfH5Ki6LQJXy/nmOCT96sRoEEn5VvQov/CJPi9qZKS+wipo8A79+lDHy6HAjqd
Rj0cE0YD3Wd7Y98gZDaORAXFVyvfWcHcsTt7x++7BtmuraLVmW/H2mPb4Um0v1n9
zXWTKj9FKPSJ/OOUDLgsP1Rbb+921bW1NbWMCEiagSraWHDhSfcz5QrGaBSSILuA
BR9MVksQosAjU6iIwJMjedzV6K4PZLWNDTmXVqwq2lBS6xS/pJOnqqffpKO56azK
aFngt4mSECK0H1jh2lxQ1k7imqbop+D7yDajTnJi2JTh7aaV6b3P+8jg9ys1Fl3H
uubNXDzQuXkl0EYsf9q18FaCay+k7b0XiQvkNyyDxmvOMAohDwTx0PW7+Ne/QgYV
tUUGZVvqJszcRs2IN23kyovGMawRuuDm+xCrzDQPkLs2wcgt8NasGOLjp5b60NZ3
NB9UuABs6v8j5CJkS4cvvll0Zh/UOZgVEUJ0kv+7R1ONg4oGbVPfrRAat48uv1Qj
vq/zbRNuqVh3jBThYX4rTR9Zxf0oc+QdOEt2OHE9qI4iUGnpxCtwzyh71rBbfF2T
IiXn4R6cy9T5NI0c0AdM+z/s7TbGhAdJQ40KHDxXlNRBuvy8nQl1CJOjemlbdkgI
HYPXYCZTxL2HFdtR8aO8Xga8cUilII2Lz3A9Ca6ua7Lb81iUna+st5hdz7zoVNuF
eO8JWue2WhOGfpSJQ1ZUpfwHxwE+0AtIFsUBBL7mZdNnKO5SXrBXvEqwc94LocKH
0a/Nj8Vh5BSl4C3ERiQgE2x6+D3E0DW9QqRn8F8iW7Q3I8XU45ApWt4Ake66x5++
RUHMjLAVb3Kcz+7kj8UjTOh38x8jqzIU8nIZ5CwHHKmY3a/qJdYutqdR8oC94YVO
PhuB5QPoyEOeffhTbEcSufkacD3MT/OmYcQLOM5liJkDrkFlQ/GSE+Ac9XEcpiAu
WqUZeBfC27vsDaO+2qFrfZT+Lbyy+nHBc2a/syxIYc0CKDHqbIzArebIMyzsaQwo
NSZpIQo6ltgvFMO2lscSZ2BlP/uKYMrEBBuCjC/Tp++zZntzosum4rRw6e4UxExn
I+Si9AOnQ3OtnhOnaAcn61U5kYIXvblOMAP95FDrG4ba2M2S7kERfObUo1CJn/TU
xGqqiggoXeI1c39/wryklj+YO89RZi0erREBpyhRXaQwWwpR3fdKj/MrZi96QBpc
q+0kkRKi1fripmg5vl85FZE2U5rzws1nDldsxUswCFoEUrXwrcUr9LZ5dXptcYp6
dJlMnLtoxvFM4eXwe3PTXNOzgh8VhDraZraGSOm+dG+X5NAb176zbCG8kHD9YJTI
dzSHscx5pmGFFhEZUuW+MrR9AXXRArwWv/4qQsC7WneqAS/Su+ArWAVp8H0RzgSE
YyA16CpMmybj+W4bR22ZnLzvU5i1/IkeMllUj4N35VVxzAx7pP9pbcOly4LzezrE
Y9VXSgQKvPBQqc6MP+ldV+ocuFvEfJKqtBW/2lRNerFMA/EE9K+RVUeAIrswYfBI
CWPMNXe3d8qtKwV05yIWc9rEKdc+7h8LonPdb3z87UwqgjpKWCJG4nDofmJVelz0
o0WGOvOQP8tiJKuSyPeNKTt4Agah15vUj9b9xKVmh/wwvt+w+dulY/J4MWWVVINx
eDuRfPKXYe5MEnBj9tV+AtEiCo2PW0g8oGgozQBNKjdV64PDvhZJzUhzwPUMMQin
3/E7jDFy4/4rLqur3Z2IivdqhbmIBTZYx7IXcqMRiQUfU7PBQQSMSTdfQwpRgSPF
hrDOkzOu1jIpWvJ6/Mf8FJffJhVDwmwb6GLvPUIiWmAhItglNVsp2knR5zHt8HDl
NdToTQhYaE0cr4/sx1Srzhqd3ui9NrnJo/ziko9rcKLIoSu22ElkXNElyqd2Ygzk
Y5AanbA6eVFNclc9vRDwS2t/yS21f/Z5BcP+4bwoOhB3n32X1DBjrbC9jewTlc1S
feazwytwKmTyIoFqwZsXfWW5joP47YZaPFX+W8vY4cbr7M06rWDTemLKTu6NIh2X
o/HalW6JLzZAc12Ex1PSONHUdDDFmOfLXVfVa02LE35FqYJNfkapi6DxF/vWVDHk
IUDsCWJNKJns/lEtYF9r9C0Tmv45LyaIeDNV6x7SyrKnOjCxhj1+4A8FkcocXWVz
Pc5ePjxtIQFVbiHYL3WLBkh9/F27zM0ex5vCi9Nd9yKYRm/1i/U9ZFbhHtWmlo+f
aubk4YH94ClSa2zLz6AK+lQ/Zw6VZE0Twlgatt8lDnT/5otFJSyXfJ4Haz1cQeac
eIfdxuZY0GTkXtRxtUNbcFAGbDfCStFkuRwRn959d+tTI9fnnKwjAlJkm1BndHyB
eclYY/D9Abw+5ENJ8M/REmyj94M+6lm2ndxOJhlsoBp9wMZpzNyYCLnzP+qGlfj/
Fm43o6jZ91uqzkk/BRmcK8oPMIn0QI+yRxdFAh3KOGaYp8xjDpDCvfMXLr9IjBTL
jO/q/xjMUg/DLyT2h9vju7Z9DFro5+t0Y8W49vDowxtWLLXnnXLNuKrHLw5npYvY
Qg2tUoidUfWLSA1UUvVdSjWjM+2WAbFa9T5Z/beTCgH9b+ZgqgaisQWE9F7GSqE6
68PWFWlIg/HmFpt/lP7IczTCUCT0nJkWL17cCALcejlMuuuxaIk3C7b9D8invPzT
XR77Bo5zi3aDnxyzDMxfKe+O/p4JxCCXq3o7nNxm6hZ4Z4FoOM1v4ki4clUpuOxW
7Uzvq+OkRQmXsyAsNGTsiqJR8BpwqI+tERS2R74bxIEaJBoEB6gmPYNDF+rt3yxa
8ywbXSLUKH2Yzm7VIorlKictLu43Y0t67Gxv6V8o79fSa/qVBl6AL6R607qevq6t
hf7oSBMsvanCUyFWQpcUL5m4p35eNH6K48rdY58+Xi0LSQwozkNCz5MovYK8Jx54
rYgd4Fs8yY/AIVAruBm0nEXzxBbUvXrqaZJBOlxOmWosaZJPOK4evIBNhOLnbtHC
SICoJTXVaRbHePt/r09hAFEqkMPOc4HGn3g8MW+d+L5/LmnQ4FWaiBo8nCLh2bI6
PTRERrkSHltr+NIQGgBp/z080C1KWvU7zUwjSCeIOVqKMFX9D0dWZfAXPM9b9fhW
MJ3ftLpGYWpPptMe5HPV7P2/w2qgL2bCVLvfLoWxcqeHRhMM5Y47BH0kwEJkW73G
WC84PRAbEu26FPzL2FFTKndB0Ox/NIb8zylBF58KT6gGWNc0jeoH9S6CBv3ypPZ6
LhB1GpsQKGXCQ3OzRq5C0VVWTFfRPqSQi096sC2lLIfgrwcTeUZxa0oAUUMc3yNn
Eu8kxuiYM5XnLoklNkUJclwbC9F/ML0GZnoX2QKkTm8n48w9IyFyLnQa7Syx0oXE
6L+bG4aadhGcyi5saPG4ADGJi7GPVR6y6kvK1+gKK6tstqqMdY0h7r+ttLw5nLAr
ZKZlnAWakmmMqYJMHBH7vf76e6UjFkmruKieijJk2Fy1XuEPHgCE8zXwHE6yXr3V
RI9Qa0FpslJ2KQM8MYdtRSwWAPJpyaJFjtLEa4ZFfsEZk6Kc+8siYZ7cGWhMSuPv
/5JHkEGxr6GdGV0QzCmDEfvENTSkS0lA521IvmV7RdY9HJH7X30gnS6uKE9veFv2
xggBkaqyJdZVcLUXmuQoaR9404TZb4sQ8kZ9nyrrUvxcKaGSmwiwT5bYe278JngL
0YRauaf+TjLPTN+EYNOIvCc27g6AJ3bb0tjxgSFR9mMUD6pLxPcHnrjxQUQ2xLTv
ENs8scvTvurCdqrob4SWnSqUk7lL/BO5ynX7wYrBl+R7FWp0/gP1p8ZIGD38GrOr
8Y5ILom4zPZDxcvJ3S41HyzHLwxHoF4kWUndCZHMWAlzWrCqtcERwkNM3Xux72z6
abaHIXfkAbJ0m2wKY9Pyd2zQsHaRFPC4qHMI6khHyuiFTQ7wV0KmhtAOq4sWaz/u
tGFOzKn/4T+vVtKtMQf1jnR3AtA1B4nVsi31ql5vYUaQKGHgrpl/u1Ko9EojHetd
puixuqqeHH1LyxTwsdQN091exvh9ojt1a0MFs0Fexh6T+9VP1M63D3L3OwAk+UxS
lksdq3nw5iKAvxTSPyEF3adyMgjNY71cI7EFHi+jvPql4L8B3YfANy3KFMs7RJR2
hTeUMVRysOzkhcd9Hl9758YQLyxikLSSjNmw2af6QbcGHK1gAkqBssJ/I2bzb4T4
BqBY38GjeqEl/Vg4l8QQP72VKPTnUp1c78UsxMajaEIqizR+zGXCxKdrdr4i9Q/B
sIqeGZGri5PrFJsMMQAfPzsc+e7I0JPD/KfXAi5k99N0RrNXcxHAKVmDJRE1mu+K
vF2qq8YiTQJE7jCpjArJAfT+HQ+lm2eGTpQn+FFu/LLzooONMsZmMuxg5smOu0cD
GRrjgNhyDhi8vwUxOQ5IUFTxiIL5v55617kih5G6oTRQ4kC18zOThgpVGsj0HcN3
Xz23+JoEf3pW6IpoNfKEuF6mg+2NpAX+4UnGeti+6NA6bfZJelxP9iR5AI585PJc
8Una13SxL2u+ApBUUvo2SJo8HvU4+okucJA4ZpHReFO6nPezatkDci6Llss6YFhX
zuzm/ohU6XEA2OTXytqJsXPvxLd6Y++/ULwhcixGwsJ9iLsdxPoyyjckgrGfDixs
1gL1GfkxWeTvEV6iYKe3SHGxsqtwC2A1GDIGYNQWOPCfnm9/fb5/XQoUO9h9Nbbv
q2iVuLquuF99ZwBxFpHoB05kkKfkTYNZRqTwIzNhO6kdF0HPtdsOOQEKQX88P26G
mwf9aM1fhAXqvtSKIiAzxfiSDM3rcTNlAVyIqnwZMAJf1mmJ9x+lMXnhXQQXCkor
zY5UwieNtS2qAGY77ifSIJ5FeGGzanFpgJEXlZ2BxooNlimZq6G4h8Lu36zI6llV
rxsoIgEwNJVWuADPmaks5fwf4RE3REkiJ0k9mWQV8lRsFVKqsav/r483DnemEoki
9NETCPuCznjiElnNg3jqydozKWZH/J/lXo4XS6hdZJVDoOhF1W2A7kBby1XDFVcY
WuNyMY2FCcKsxeSKqFAEnjRHsOE/qUT/bwhXLyZhLfGJPPmovJLatsp2kLgrNrBU
Kxr7med6Xlh1i1VyDT2bSU5Z7PsVTWYQ5vDVzn5GK24tni7MFiiOSRr0M0xxh5y+
kXJurysEyuRcpl333ms2n9if2RvQ9aTMIvXfW9YgAEZEiAR882piCJ9NIC++OSL+
PbbW7ET8glFgUIPAgZ3j5lmJaoIzaPGBP5vInsvpPpl8Gtqmo1wYTvG5QlIUHKAp
XRcQL5de380jaimCG+G4L9HDC+Vb+4SL2E7jWf3qmzsXqNKpR/U4Ghx7F0N/IV05
xRk1pzC2At2rwA/QWnIz+8u8fjZSxcjDp3OzrYHkBdTPBMaTZeUDA5Y7Wnx4TTbY
ewySP1KWcOvX2XahAfRFpU8xkpWXl/l+CCN7Y2nQRqDyjQqBDTxD6wic/rpvjLEI
`protect END_PROTECTED
