`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DerTtvjD/YW9eXXn92DbMjg+lLjCaYC2ixa1Dug7DknzwnDQDno95SFATpS6qMi3
4lwmKIG1XGsu/pgeZfANT+bzhXCIHmnagBdzb2ZCSe4eB5kNVx3KrdgxZo5PbTnS
7+FevBfE8Nnlq3GMziRaf5v2J/E5RNmf4J6H6YxZfLiIHVRmmQHldG02cwNRZyqV
Fp3im17ncZOeUYK/Pu2varP/ec4OA2KMnEqO56SKtzogo5H3R2vvknM1gAKRcxo4
7Gqr9Qz8DH/54Rur4JWjgfmMBToSnBPt1cM8qlGCHEx37EFXstEc4cKyqTsQLnej
VXQnokJjniz71PZ3yp3m8jje5RhUSP3f5BvlDOCJjwS/Yy01m2ZJIL3Angb+fbgc
lknAfuQzdVBlO9NLp+KJfAioFmjr0SY/ToEvdpakgIlEPiaN1ipiIRtfWSAVkKZA
Qw6hpGy4IJMhaLWLg06aHWcv8lhdzLBf83jY1uGD2K/SMGcml9zu+YX5sqDb3p+Y
Se8jfveSyyJxJYevB9zub0ys6L2pr+kd/Ma28OM934h1Dk0Qji/6MKUxB0+LhMih
dA/2g9X9Wz8CQJZqwfORG+1+AIQr2bTAbLCsPThw120FS4NoWPhSfZ2J+fHgWEds
pnlqA8R8fveCVKYKxJ8ExDKaxoYJEKgFdYvWhCsjHImafKZkUTb21vIq/oXYrLin
yQeq9rbY+yW2jEp/t/GUkWCVnXp7vtxIOMCN6UyF75U+l/N9CBKeDTBZXSMeFvcH
MGj9Bn6BzQpy/8dAxIJoeOd9ZcR71Ecw/6i6/LXVc5H91XL3osKkLJSjd26/yiU+
HAC3LChUtfw7eCjc2DDzLlueqbXxPVCyTfR4FYz0ET3swRytmyonIkIWBakAxIzP
z7wyoOLrXGhM4y0mOADvzm1sEc00QRVxTcGlrbtIZD0dglxr3/ANl7lJAo/AsE0y
hXgzTkGGEZEfIUuUsR/aCx1h3QklyaSXzW3mQABeST25FHKDIuyUIgy+dND3Cl2l
cdG16ZkquTUO3OKR837jjXNSzUT5rjjEYlAJ3b2P67c0+BtY32dciJtNF4YTFeAL
wbxjX+4hTDtrQHgogspvFIz4oyHeOWfzMSkUINk1ddh6IOJh9z4nq+Fs7gZuHvzr
fD/M7Itubx4Ls8RxQXJStXjoox+TIVjQ8C9dQbdYJQ2zeJgtXnKDP8gbTrPIN3Er
Htpmk5LpRY0NFVQM4/jX2lOuQnHj9+QZxZqu8FveW+1ZYBod8aE+3E0aW0cIgQwv
WbkpVHPkh7Q6744p5tWmrnBX7wZq1RMfKXW/RcePeuRVc4mISJtVt19ynuCko+1a
WKJ9tMGuOr/4cN+DgMFjKDfV+2GNV5+r/f7Op6VJVUnCCdH8NUke/QYejiCqvHcP
KxR1dEkrR7HHy39LCRl9VsaVeWLvgH04DrpgmDFJWG5el7W53HbDkAiuidroJXE6
5GCyj33uiSlo0o2b0cW6t5CkM553Wj4qCSXuinbqLj8d788u5fbw61YpTs12fFYu
8aL5f+vxqKESppdX1h0YXEluWZfX5LH9tQi0giI9nQ8OA5y2alETXYLiRtSxtHwD
QbGvnnt4E/PNvdNH+yo1bbApdjX1EaibY4tm1kJfkmrcCpiKXJBuKlYMIymm46m5
S4Xajow98dKo/hw/f2oQ5CF4UsfMf+khh7n6buaR3mCSicZTYsTy2WnCzEol/Vi4
m+5+6wVlpsNll6+moH4as3po0aXas+tn1k1LffInNvrDsdnI4QaOPhNPYD5kkYXO
x+W3155BwYmeHavtETmY39MjeR7OAo7Wx5a35/PWK9bBZK50ZZzHwKFmuLYH1G1Z
w/TFMfWt3uH5s7By/i56IHUq/CXg11G9GJkiUgeRqsrlUHeOBWbnmyvfTlN7dmEI
c5U/dgTEBNsY8PYRIbRSCq2C8RyhLEi/djffjKWdSaFuobgmUlOG1zDlmR+vN/tj
ndcqyEgPkoyr2oZ/gtR7zTz3mbvIvRG150irxyQ2ghO5Yj1JjOpxgK9eu1BJ6M70
Z1l507TFhsnyafLaEMXiuWx4n4qKASZ3f4hUxLc75Ct74kf5UYAYEC1P8TrqL+gA
qkOx67+DYzUjN78tICeloQpy9U6X1WgHBt5VujLEQrc2fMRpC1bWrOCtmHXE4FdC
wTaJGqzLudlP7PB4nLX6bN2xTGdUputjECXSeP3J3L8quNrzGqaMtLINuHABheSF
MC3qWDuO6ADGGUjd8mCimJpRpaj3P+rpBU2FZ79Y+hTydHpS9dpgHfQ2DSw+0lIl
yx12yqjrxNcb2MOCFLfTf0DVAbHdLIquG/iRC1OYnQl20EJM0niYk0BruuENdHQu
6Dk5hnSpTV/KljDhNoyObgoHf7c5GMm21svh+il/AiP3VNSTiSHZSiur2saj+QKw
cya9QO2vUmfLvf/IvfADy/0cIp04OiFFFG8NQ0ZwFgjFSDlIfaIAfkTUlmuFjwhI
b0GRE5dyUdHGgwESntOjbA==
`protect END_PROTECTED
