`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFUPAOBgNRoMwzqYvuBt4JE72OwXvQayiiwnheC//GxMuH8r+OAdEz80ffoUqAP/
mPYuu95B2/BeJ1pxOO7yd9u5Y1avRJ6fnqhTfT9Vd+XfCWewOZ3grmH1kHuVoVPB
TqRpApEz2oxdyCyb4bNSnSmd4SllpcAr1Og9RqY0HAsFbcBzR41Jd+CZqPh/csgS
d4aPMxkF9K/W4teJh/HJ1mr3JMFPtElhy6JLJ3yCck9TNIwNZgp9Hk7ZFLXk3RrS
covQF0MByHKDJy14eBoqsxzUWE9sLrH40uRrIEkUmQDCbyK011oMa6i4+MqI48D5
ecbN4Fb4TwCt+MmAERAUgw37EBFAEEv3mGn+xm6r8Dk4EKMZMneYaWzj0Xw3FFZ9
kMllcCHxgxlFgp5EXbALdtGoUdSOP+51BJaTSJ+3w0hv2BJ43lIJB5vchm3pDc76
NVVUBMjKQ4/0c+KNSblVjnKe2CDffcmDP0XDKcK7aJ2CAEmMtk0+ow/Rd3juZ8tZ
xzRSeVd7yw67D09RFMo6k9i0q2QHc6xij3FkXggtKGubAY6olOFDnJ6l4XSVFSET
RDTzrUN/2Jalh83kWC98S7Uq73vOOopYYR2hLYOku8xJHhxrv3Jczxve9MMCEnjl
x0Xl3Ld4x8sPxQ/VNwVbzAeFOEwJ57lsi/4LoqO553fBEGMz9Vkb67AwdLRGO4NZ
s8AlWpj7iy/IFqSypIi76LZWbJjnKTgcZXjptzYXAwMp4rzx9u2wYcyxSQ+E+/DX
0J4O2V3m8OF40J6BDOQO+GHf+GTEujR/HlgvX+9m6W+MSMy5dxh7YlhKAYAe/jEh
Wu7xn/lLR7Mc1F9to//1LcQawLXI20NHG/UaBliRtGSFvku7MYO+YyuYlh/aeYmQ
atIZtxSCvNQAhdS7jlPIYhNwwo9g+vlq59qn8oNzGUU=
`protect END_PROTECTED
