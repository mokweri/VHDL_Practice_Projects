`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/pbCgOsE9EZKUOi8xlyEw1Ga5PSkgC6rwMpg9RDv5zPzcm8FO7bwcSt1JvYMwQYD
NPfoBWR6AUj9jiNhtUxRveF+ZzWtdzCpUbmVf3HE3XfGX3e1xEWwOx50/fG//r+9
mY8p+Ow0CrlsciSAW/Qu1dZ/gFGd4GNLkbvf+A2Pm9fyeiMHgstsEwYLeKMdxA/R
grvNLR5Lpr83NuiowiRgUaBVvT1reCxMuNaWDeeQ+xN7ToVV3KJyHXolvHCInoqb
2L8Bg/KVfxZHyy+1K4686YjHmOYoCBMA8JdkokYKc0wD4wwYYKeqKhFh0Zs60s1s
16SGeBrfi8gAnQjCsU6yurZVldGTxS1WAKkEkOSFul8aguHPcyJKl0YRzZ/8FuPd
HhrfSsyYPAUfDrshoYe5EFG7u1GjHvJpC62C7oSeAScYH9KnkgTw35sqltrpYJaP
k2e7VCEdrP/XCYQxMQDPGiDqreJiPUZce+oaZ796OhbDBP6l+vl8wyowFBkO+PRr
iHAHSUHTTPpiiT8zaE1KTybHhQXZZVN/q01dxZ/KpAZCEaRD6K3Bz4r1Dh3UF5X1
Sn06J+Q8tv7Gv2uVgIeqvQlRYoNBa18Q88KU+2aCg5+JqwtmMRCPu/8jCb5jv/wx
X2y4wCVMaZ5FDTANJxlFOQPs/cmsT41uXy19Y2t48zzDuHNGzudpQmznPCpg7wmD
mQ1vvjd3/o8KFuik31LpidO7G+85dWcrLFKllwA/V2pBCQVGto/G3CojID//5Zfx
zlB+Cp8kfBFqgw3gk3dpqZAKtFBfPf0v8F4Va7dzcysfTGqdhNhxg2IUTht9CqHd
sBXR2eOSJFdnN0do7tsA3SxKWd1KpB2L5Ci7pN8Hu0xLjwO+kkJupyXSs39C19ph
oZGNfsuyG+uHbwKk9kGEG14dByFpMKCr95swUxa/E/az1GATH/XyLEzm/OYdryPy
Slb1JZZjgRPGjs8aVrdo8/9bPPYJunToZJJsMdy9TXzYE8D1QHND/HiK19yjvytL
N132JTdSEJXwoAWjqblbNlTM3ocgVeAgxAHNdIRAWE7+ElU5+arfKDkB2y47Kssq
O2OfurQ2n8oIYa+c5VI710XuRnCUipXKbZaIH/3e9dNBkGefSjHj9iBJxBjSX6vJ
qMdjJ+7wlSbzJ8NTETXmvJJcHjSXJWqJOoqDbnC/AUrUdav0nb2cCvPE1SEAe2Xh
YQ+TyU3gZ7tjMa4+fBNSUiQ/s+lR1R3/9Uq+6SW1PUz+bKyjYg3INseMuz+oceEa
+NzdyZMBBPjqnRrenBvPdSKaMIkkiuq4gVtNaUq2dc9x6O2BVl6A66smS5kbryBL
ZS/mcU3w0jfpmaGwzH02dCze86QvP8vleYsdvfHOgnavsdH/9jUpBFx8+Tm334j8
S9DLvEkJ3OLH1aXhXtXjxGDhK1WsruVT3JqUTGI3yBzeKBoZs+kVu7clSe3GiLMO
semzYm7EZt4gFMSeGSF6kUYOLx03PSsB/o1ub+uZ4gVY2icfiKQBnHLY79S22ZQo
CTtkblQ+5LegSGfSrKVE9zgAtYqXeAplZVBrDVszXVY4NcuY6VQSopI6EiWdCBaA
HWHIuJTE3zBjVJGMVg0W7dd4KciYdW1Gaobkww2TwmnkeAbIdS2nBfGdHNOoECHx
HlOYnCkfCuMhMI1wp4bDH0k+xs51cCEeEJuYqlGumDbJWuZTDnHxMJLVIoZo3fOt
1czMSvksU/kzsHkXLvF0m2MB7wH0txJhqsJiJDxLArm3zZS+Gm63cnvDnkg04tTN
tf6zVi9b4ZAXBH+vAdz+0SMUB5X1mt4IV1cvH893yAnH2Kdy4qvxHClCAruab+i5
d0bODrC450eSS6ApL2dA7wqCLKl84lmuKfBI5ijeFpbg1eFnTD1VqJ1s+ZM0blNR
P+eQrhJc7SBuoNzhWAXrgmVs/DsKtlrycwGIXGkezHizbaJ1zMek77zbAi3qwwA2
3DOd5vRAzqV35vZ6sQhhakTUz+Jci3YXlOBu+6j70q/87GwmEztMXsR4qzr6QVs7
iUiwaKfGATXSK1AgoqugKmSHuREjT6RFd6tsfC3XbviK+mPv3xiXt4qdfqkqMao5
W4uI6car1OLZ5dsR3EGv2X0OLweH+XUWPWPAvb1jpF+P9/bxk3ZY5NZCmAHOBWbT
t6/YeExCiJelN+CwoDJh1D2gy3fDt4pTAXcFJu0y8w1eQXPB4TrVj1vfpxpJrxs2
rvMBKr6jg7ElBkTvZbgqYZhzkW8tnMyDA/hLMpXmUDv+65Fn37uymRmWBCB3zof7
BUSj2zGa+8R9wwpMCnzGTt5/YaxYwjJ8OAS9mCDzOJBrK73z+Ugd+91v+P15EdHg
24R0/qQiOydhNLTRdGEToDChvZhizDaYgCI5j01ddy3eu5MQnmI3yQswK3IJqSY3
d/iQBegF+JqfT+FYKNuQCCKTWM4Wjslk4TsVKrK1Y5KUVguf4roTHWOeyt9qcJYm
DC3Obi9KaIekt6ZLWpCyTN6y34f2Bv2HNAs1LFPmJo9eP6bh2ZZXpzVVwJVZtKB+
CZQH/5Q3Xn6mVlmWbnDMbeJvkWFsVppfKw+ncPqpPdVPxxoPZWZe7Gr/BQH6RCxk
4/5E29cJ1gQu8kiXGtjw/onPRDqiYVpZHj4/oFaywF2CyGC6XEAEgpjU1NE2L4NA
E/Z4QLzWaOmxTEGjw1AUxShQjBxEjstscDP24L5v32UAVu0Pq0YqKT+AFG2H5xJR
jGGJcDZ7yb2T+IW3OR1Lwe7N8/GauzeLF1iF7VvjBFyydYuVwkpOE1FJtnVkIwnN
y0ZNValtVf9gULfH4UEFO25r17wUKNRHl+tMbi0TT7iBX4T9wgr7tHDWa22vyL82
vgAuIsgqFVEGb5XZcNpJ0oSnsEg8vNlxLqbWpIEXruhqczATrpLB97ef42bmTJUk
iynH2in5IlHupzgNpxCOFdJCSI/rPQsJ7DjfMsGdCvyL3AjyU4RAvWVesC/LJMdo
g4jREsFg9eJtsQSA21iU0SV2vOAugZG88F+ovCPPIDq2BzjpTUY4U85BR3xUr+kS
dZ7KEEM9FlCfbtlpXGNxCV6o97olipp816OeA6WYu8tG8MSqJ9fPFQEtybMAM+t2
9XzJH6prOgAmDBuWJdv/7OhCw+22CwbBygm24m2VPCc7RuY/7xuNAMIojK0MDiNk
iWTD61HQhZC48LrQyDmjPuh0W75CyoMjrJ1n2UCB9KJT7El0ssfUSECu61PCaWjT
Q9ubGojwVe1X4Ky9D3LTnaFEexRGuv/Nl7sUzSPcNnZXgmYdP93jrPAuyZsxPgMa
/F0V5Yay4ZXTG2ORwVw8TST7k6dXGyzJr/R1E1RQ0RmLd6TohTmwvrqh3icvIm67
2p29TAL9OqDqPm0XAWgLNLyVFzwUaU44jRr9LdYQqzV+xRhtM5wP9HdHoWkOeksb
6MaHiSdKkYtiaKJTzbDkVEcUt/6D8+8FMZXUWWM9x0aNSXsr5XAr8uTr2G4lRrvg
ebtQFNWosp6JZOAAa934m9TGvjkIdnAmGHgDSRGnIfn3Q/2X3Utwdn/LP0gvRoY4
TlHZgVNMNAyNmMauxerwPFvTpi3ztKJH3O5GQjccN0yZ5Q7gKbAEsGgpqG1OlMtz
68yUh0oAfP0BV9Zzc3lhCQh/Zu9AcBPI5O7OxvjbVvhgyFluPBK36Ii2I82oe33I
ac2qX2pFuqN0BqzkuRRA71kr06tZ7zT2LOj8LwK/eFLP/9AGKyTuPufFhKz8/dW+
1NxsYmL5ZzLRKXL15yEJgNCQiC4k781hLz2mi1GP09VLwlhofa+6CVWGdyacFwuF
bKzopUsltErDB6S8VqJygTBmvCKJlhlMGSz+8fxaCovD7SjgK0PM4nk/Z6rnSfqd
P/jpAa6WlrOSwAkmSJGc/hOP8ytRnvL5Azzd8kMedQfqiz4jX4HkCa7WtaZwhdlB
Ck35fo33Iz/9hyGZgMuHUSwA25Pcirepzoo66MNkfuHRbsFCl+9/iC7GiPwqVUqj
Z84TBhvPuTdgtNk8TrEXXCU5blzT6Mb+J1L7l4x+i2IWaibOkRppTHlQrebBjzZs
xn9gabRKZv99Tno8M0BkvMECgMtkZRosv2rh2VAqZZG1e62je2wqVBLj5uagUaiF
61Mdch6nXlN8D4CPIoMMtESOR/BEFq0ymcSiRLfpQgRVlbFE+CgeiVyaXVDW4Gf1
K3FRlh97c5b4APoWIrVsqEMg98B0XwVYJ8nP23r/TDKAQR9HH4gWYj0Fbz6fCNHI
TCv19MSZ4tv1cxBed5K6J6+j6HHZKrhurBMtXvTXmRezTECuWUKW/1pHvLCuj4ve
3UvtwEKFGCw6n1+TcsLeVL0v93CAVh7DiWjQQozNq1WajU/BrvrdPfqtVPaxBKbE
umyi5swKG4YLaJOGEMU+QJFa82nXynBm9YBsnO+M6PUdfxarWY65h5awiopwDk53
WDGMtKQ9wP6rv21fCaoV5WliMMoD/O3+84CtheK39g6nKCw8hlYN0MZ21zGb8hTl
1+IWA6DTXSE/PI09Q8Lljf3ZvEr74Eh7Ce8mr6frXWZAxA/WaoJMeJq0kN6oe/MA
MRTnc8948bTOo+OhZrCWsjXWFn8iOINK3gMCSKJUdamJcI07NjR0IBKm9WJayb+r
p4YgNRK+2VJbXKWEvPAwrEe5ieD4eL2hZEZT/b4frbGPM8GA1D6J97/cxo/9qh5l
4rNvk0ChzbtKpbfQMkacItAOwNN3Xlhk/OQhIuqsy2rs4Xi5rSIJWFJXVOUmHJ0C
FWKMlgt5kWnEhCzXjgIVOr+r8Um2TFax8uThFk27Y8OnV6KySZGdzPD3U/tlexYY
tk+2y/48gMR9rt2oqbWA9KKHv3OY9lgMM4puXPFbBkNmne8zPode98gfVboOQocN
hc6JvyElQDieNaEULldMvnPixwhONDTna8dl5Qcv1S1iPm+V6OOLofGlrPPCrO0T
l56zDKi0bEFk2EZykr6lhQya24i03p9Y+/NMmxPWtUX/4Fcgxp9GY+6hRNCf01Un
esZ1WMzBxMBmwYVKk+AkeK5bJwB87ACav/Avfs8qqlqhIEJXgQBY9E4if2AvHza5
gQ7Q9INoLBY1BtYzTkw1Ypu88DucV0Fm5EjE3ZdsSqxZh+1wQkgfh8e8gZpax0BA
VMw3YMLJIaL7h6VmrFhII4Ie71vCIhoQBgTCd8vLpA7CoanBQV0DlmSQ1ecsH2Iy
+6BhgeERMtEPPC8tjCvMWPk0eCSz05MCOx4C+PK8NHtoyDSdg3mzbj9Xnjpk+ZOF
Si8mlu4ocuBuE5eqf+MdHhWI1YumXAznvjqBAMiLfWUCYLsO2j5qAUlNsvwmuuAZ
VAk7y4/EUHv4zMJ8P1FxFfGl+Yi8+fDrfsv8Cv3ly/nossxiAAAbfbxuvQWIcjsC
F001RwfT2oWSc+iorASF3n1BVhTjQSs7U7z1rXrWFCBu9kUKNipJ0rQksYPzS8Al
KdvhDphRV0gtf8zGBSi4tT4j63YrH5LUiKb/Ewtu+xaFHe+wlrPqh3TUNQwk8aIs
cHkL5pQWJOLx9tXvuWeT+MobnsEWnUJjkLLr0C+C6w8jFRdFOYu7nBqkasQhKMs/
iNOOIk3sG/3wa0Dwg3oSG8ee6ywea6s6zGW6vs9IOQEx3oqCRSJjLrvVe8GUuodR
wyNf+eWSQEspzUzqwNKqI/ONS8pja753x4w3BnnqSRwb/ABZfJLTH82O+DLRjwN8
l19ZLkFFZwBBvfYtrVKTrWXyNt/5UnKSpW1WqE+IF+PFNwrjyi1h6MsIFQFLfTum
5Elu5/Z9ckyHUt2vip3weUNHbINupVRzvyIxNzxvoEo=
`protect END_PROTECTED
