`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+e5d7aBLdTbVO7gXwR7n/16bMYUC8dQwsOeAYPgWitVzGp3/+S68Mbwgr8RG1gBU
2onygL8Y8XsjdzQzzm34NuWeMJLDljDIk1b9fAXDZV4qWh4YUpYo1+NXc/eYdigI
jexZ0CBaSWMH9glxjCYxTYPRkLnI2No3+3LQlpEaDceusEBd6T25Kxe69o7pwx/O
p8hFeG9+ow5GQm4SiHFLVZ3WtkY1mFi86R+RHJCyKpddcMDR5IJak8i8UZjhF+4G
ElA2O5UIomAZ7ZChbEpTAQI1pjOFmq5gx2bbxBOi3t2S0Tri6ZaB84cxD5BnZUCd
77OEl3Xt6Gl+l2WmwDhGO+80PcQdA8cACuGoSk30fDfaimwR8QjwasPLtvEa9cdJ
SrBP1yq9KK/yoPs3gkso3SJkjZwfjNyN611/NmeA0OkzUt1AXPBMarEJCUP9D3Y5
VgsV6lzxlt4Ah7YjmMKTMHsailN7/lmfj/t8yYTSLESUrdTus0pW7jn+iqSNl7+9
XSUzGIWMkdGQU1PVgRzWv/MfBBBsvUBEFaSYatg3nHQHpVSr+NQutUGshdgMWD0n
sQMtS+PYNJ30dtbyGujL5ujdS8vK+1U1XMRv4QAt0C3O6LzcmHevBbmiw5Cw/nV0
YqTCsKbbyLa5taFkJlviXj2C3+XR9od2kxIU2EpmmPb2nh8so6XNBZndgOUg3P0g
npIV9TSoEZlTQyQLaaQrHoo5wRkbtso/alnTigz/xWSorYlQlsc3flsevjkqE0Wt
yzmLFLjTcoESsvvzDkcKR2JbfiOifDBJKSIoSp2QJ3XpCeBFCatZcULUo6i1xGnt
Cz/LNfdU3DGO9Fnhp17VmpIZ2FSLRtH3Us5ax7V3tPfndYvN+t7qZHDFuTagKZ9p
`protect END_PROTECTED
