`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ziUS6HyUK183frebFceMrkyjrzuOr4DBn81RfOWjZnLrRiTKlfr+Bq+MxhTjET2
GBe/bf6C3yIABVDg5tIAzV6Qq7SgzbOXiFpeKARkp9hnfwc5we7tRAEZSgWxohkT
5dHec2WmcJqh+hhwdTBz7MuX7FIGiZj4PbRj4RDd+AL+Z8gul2DC7oPDWBytsj1R
S2+DzuDyuG6lQD8sGLzQ+Z2XqnDzVfzN8UO79RCJ46BQ6bujgmGECYxfPlEYgo7m
xLyuxOXR6yTUKj8A5GENHaun71h+x7B4y31lpAyVdVtG81/rmnR4c/dEsOgsLdrN
qlYslQslHuRacEm/GAt+Q6KHDZ8HQi91dRKtjpdZ3TqXFegF7cYK3jGgwbx3Xi0j
uLsL2sE1HjWEZ8EZbyAws4bdbdEeY1re9mljyxEXgy/JRrkgk9TaIIFXy2VrVdUQ
kV5APkcncX0IgzMYF0/hrykChLi+Zdzs+hcsBklO+B7hzZOd8lHHJZhRvsHi6UmO
qBMctvYyMj8h7eQAwesVEtyc5jC5KD88ovbaUVAH5tlHG1J1gSi8dcw70VAwvHYt
q2Ft3q5UTozeu3W4dONfw/jWZes5Yv2dLHaigC7NkgKVNblWVYLFmNMcWPWtozU/
HGYoi68z1WqO42YYtfLubtzqv3LvW0pvkCcGfKSJHFXaAxVJ2RTGLeSkVJvQnb3R
z6rCU/ja1/gGmJN9XR4u1z4eR40enH64moVs6g1JLPLff+tR/7QIfPmJjf/zU3yA
Op4696hFCVEtn0yI2TEjh8WxofiNPsc37x4ebDIDckDd7jj34qhdmzqcUES3GnPe
HUHuWkgHnOm9ibVPtMpglqy1ClETzeblu6+1YbCfhPH/C3FNzAb22fUDjM6j2p3f
nqQLVvmy99gWcUfRaKuQJw+cudKGusEpjRcHWGysaKwt9NK1mlfyLmt+KSI7C7wP
KXHvX8jP7Vqwxko3UrqU49zDlxOEWUy6wCaVFPnZB5wNSEy0IHnT3L5kTqP/PP/V
GiR2KTxVNvTMnbbKOj0yzsurju72/24DhWGaD8KtNU8/C6lCp0G8i6zuQrYIEpX7
sr3pyylYWs3ZSzxA8x7rxjMDlSLtMMjnvr3UG8USrpN166VOFwPfffSJ1D49TW86
AWZ8fwWU8tY6+VSu/K0j4BVjuujaFuqH2WNMu6wFMTtjUnzvGB4yMwi7u+h5rw/x
nvGWEipNmVG+0CF8L59+xQXGvCMAlHiQ+YGYXBdHqsUMy0wGBj45IQcs7MPfeOy4
5PErdRzTVbADfjPuHqCXcQPaWVRGRpx2B3MWovIMiuqSJ+W0udKwL8TsofGceu5Y
SOD3CuSnyXt5EDyNKRLZsdu4dKJSUyipshFdlb1Wr80c6Nsk92/ew9t/lZejSbDg
JDEWtvWwM4wpAUpZCs2x07jt8guESaZv2Dmd7r/e0a8b9QfoRYIPGU6xEAsMP1wI
PZUhV2fpCBSQe4/IRpf0sgiA9k1+/rCNyQu0NWCDNlOm5IbVNiGu+yjvz4n+BOBe
f2BCm1784LW0vbngZ25nyRerD1drac+uRcokE95CXHGKBoei/xGtGYkOv7y+WiLg
QI3ZQCYELmgx/HX27i+Gu97MGWSlCB6mKahAIrGdoOGKLjn/EQkNV4VaVE4UDRrA
A2Vqw569B/X0LN8iFYXATMagr6K9F3GDbXxQGW7srq4LT+RUbCAwYW1jyfY9q3tI
oxHixFn0TEn4hxzMyeW8NENtBy9dBRWW1cWaMkEGI4KsALCZAF3Keh+CXIM+biku
pjpZyvzxTPVmfZowIHrkgRwzylCIxe5sHOtnVbU5DhCVGX/m728aUwD6lO9ymBmJ
zryA1gM3zoAnGEucwBQ6poFrAeO4G/LbtfREaHosmPSTWpq4AkV2avrMtBKx6MCV
cc9nSl1zdoOgOPAyZWWvh2jPSmyQTjuoGUaX3zNg7/Qv0Mc17p7TiKniJfAse4uq
nBZImeIuW8VG+G0sYSr85215pmlP1evsiILqjDPMpGhClXPVRT/3S9rhofdV+Kf5
lmzSc8uSfeRAIV15YLyckkVNCuFeOVDa4sywu6uoV//vWbgDoR26V2cCSlBQznrx
H+Oay6RDjhYipd4ie5VJVq6snBwous+mXuREWKdEhIwSvYULfdpjcFFRv+aOQR72
buR3n8h1YJUBCqZ5vRt3RfAO+pIhkBc1D3VniaFuiyRVgLxmpBb8NbR5AIZB/daF
af73akYa4ChsbUoGj3tgKsxKpy5b+IcmJRqkDfuE5IO7HxJB4FgyRlhvXhF5fDU2
7PvaacR3dHwpFuuzwM1jAvKwa+3aW0hCDk1+6d0ewMst0ihjIqGWqRZ/826YvCG2
ZUn95lNyF6AFbqW+0SE7rbMkPfo4chzigli1g2C8cvsnONN/1HzDjKgjjI5Zi+Qv
YxUlLLj0rHGkr6Rh/OJT+H0UmsZVez40V2eIHAj8alHEFESI8kkEd3SyqWiJjbwJ
LnUi6MoluUAy++uZprPMHhkl6+rjEB/RRo6Sux/pRvsQK0T5yZ44lWS2S62+P0/N
10LXbJJ+yBmWyyrM902ujKC0/KjI1VzgsH/eCbVTcAY4bj8DZfxLi++akNvfa7Gg
VMuw0/HRnJEng5FUf2O0s9xM0Yc3M6JNp+u9c2idj1UN2bec9qA9ezznevAZy84e
XPc61tKF852OpkKoUhCngFbhuGQRQvBa2fLkYzvB19FRnx1+nsqh44yyba1hQTph
1rzgx2VowxIc45y5J6iBm/AHo0rhdPwd6WTwFAHbwDl8blNZOI+FQJVc8GdlXG20
EWURLKaGN45z86zwJHtWyExNbRdG1z+PJ0wryNSxPfM/jpb48KSo7hhnNcEAHUKp
yTC9pxJEJqGt2P2Cn3GNWP+2Xpz0I8cKOvF+ZW9FuENoEqbP98o3vBZeZu11xLeo
G/G7YB6sTi2BOvNcOKSbBcLsTo1In1GPx0bbsqbejcnFrpmq8HQrIU1BCwphSXXG
tC5naNfC72a3hCn8MhYaokm2Tw11EJ9LKQ0LL5B34nel24L3ng63qps1LyuDPMmT
H+eR3mj/g/+qPDWfNbEOlMiY0pJSI6WSt+CSptyj2bq7txTD4LIZ9cKmMkGEqLDF
TnwvGtU0WIMgT2+Ch0hItNWh7CXiLQ1EITCW3R6sBedIR+EWiS8ep0D0QkuZKX3d
qMxOm6vPR1Z8ArTj3QSaTFGHHkOheRc/djoH6L31MbAOZY/rw/pfyujAeZ/NW+zu
Mb3bcIMUVkJ2GsFgOEYe2Ow+jdnt9BeKbObqabdD4BN77mzSATKc8ZHokmAC6N9q
FwWkwpK+VLWsWZcSr6felKrCX6wjFfomRrlHsg49j9b20b3NOFiSFvMf82Hawrp5
OdkjTdkkLwmEg/xde76ov/QxpEMhwavHJ2upqMTKZhDpEzuvtUAt19fJmIlIW3jI
ycySRsmrzzOSRtMXtU8Z3l9MnLzmofxgQdJl3J6CUrQ22izxO42vbhrZUDC8FcOt
QexG5xw5p9jV5EtHz5zvkmIYfM6dnOpy+or8YOngRBFfPuI7pGUHkCprZWcjoEIe
Hexi/qzx0cYBKssex7VRua+2jhzBUL7x9nKPfAG449uRQtILZODUgOap9vX+UIzR
C3fp49PAHMcT/K5ABCIC+Pa32xLWlKk+VfO9MOSrvoMDJEG/+47ZtIpgu/Wx39oS
7W9aNsrQk1Fgc/UzToGmmyu+CUSqL6qq1Ix91hgrnVA5rKrGtVgJTwdP/u1tWPzY
zCGGhFVu9LpYObzTx+MrYkIwmPGFoIhpcgG81kGFmRniZYGo5sqi/GAz8F72f0ao
9GOXNhrrxh/V/hPDJ4tcV1OKzcxHYBkuX29ujVkkM4/npgZC5jvk8z0BVYTM35tN
zoRVZhpoF10gZ18LLt5GVZZx3bZklcjUxfJG/J7+hXO2rn1QabR7eAqPED8/l+Zv
zka80QvaAmmYAGsj0LFXav2O475x4Rv3qVq1vLUkuoVg6CH5wt2NyWlxDKkc+8rk
3ATAbyyNWFEyWkvkt1YSr40m36jUG4b96Klp6LyYGU4fg8ji2qds0Bn0q/+LYiwl
bRI6kxKStNUxxy7qjpwC+svHzph/M45m2h0LpF/sqxNVLTeZqoiDdqGad0y8q9i7
pQgFf7qmJFAPkgiW7dHsx68b6/px/py4H1Ry9qMiWB2FerLnK6V2HbXGMDwq5NuT
PqjgmgFqMB5ZrKg4rpuu9eDdhzuJcg6fg24AYMUQinhnCtgQI9cr5KB/ZF3dHGG6
muTG6CAsCb8uKmZMMgpk4KSSvX87FyLGsnhsSFiuxKrR81HXQ3N1qNuEjvFDwh2y
dQtOLJ736pA+L2bxjpzvtOfGgMHcwNSY5Te7ppzn4w7A9mYx524F8nEdXAX+f52V
SPjuSLcxeFIqD6xSfrmyU5Z2yy8gxErJ1/6+cLG6XZlWJmbTdqUVpf3m9dKR6Uug
KtMHw5FYmjoHZ9/9Ex3L7s0XrgaT/xc5edaqdqVVR7Ysg7CvTCh/u3hkhEoniNlM
85e47VmAxElKcZjt0rWpGROS6aBAmnlkrGBJ9AFuDVOIiADutquuSi4yj+yRixn4
1c4Qt7VEA/QlJbUSufOw6ffc0t44whkvD56AeiYpB9OlKfxmqU1yKMY/re5UTxH8
ywOKm/K5eRAQl7Ru2ImV6TMdbZBynNDn5vaGjRPf+vQG4SJPyEjsHBNZPTYQOF7a
GtkxUCKBkp/8alunK9PU+97jNhZah+57lET8abSnesBoAYvHJxLqGNQZiDdrEOlh
AjQtWZ5/CAfkQ7zSZ1lsXm0fawQDYUCbsZArhSnkCoF0sS9JhzgFxB83l8uff12P
8gTdMyEl3m10LB1kXTYeOTs327vaTB5m9IQjVbRBKtZvxfGHEYObvCg5O/0vpwsV
BumYVjRh6l1OsRUCt4fiqIt156+9XMM57kPYvHOhDfoCy+M+ubdVXjXpBOqqN3wE
SEuZ+kwvHygV+zcL1STl2yytPntAGYZDjxb5PlWtPLFLn5+KkikxnfEP+aONu6uv
SdN8ccGL+scDnmw68H3lL5nmSsFRAeQveBtlHk+VxJs/4WYzwwK8Exq8EbnNt5cp
rLeH+H/JeJvpa6OjXgHTlxB5bfH+2rBBh9nDVLJv8byaAPtrrCum+l0LmfjQVrOd
5TDX8xCUBloMMfS9IW+vp+JWCCeQ5IN6N0AS3m/Wq3v++ZYRiNw16vNaTpXdyFjg
WwilNiz67iwyaq1qT15SU37gi9eXA6RE0PcZVdmo17RVqrZrHIEu8M5kIE5bQ2x6
s4qly9vsUdAoaxBVGP/thpA4l1WgXb9uuhbfe7vtYMlaM4g3Grs06Y+QQHK4ja1s
uOcRSZ9yM5oVyrLkGZD4KKZnaDmV+kSLlEF8QevmSdbCDkatTZiyJO9RiR4xpkHj
3oDPckSfa/KqG4E7u2ukqYGe86J8bAX7RJXMqMaHrKjWYCOHvoOCwObIZcDHpBEI
x47LViQpeOsR2Smlt+xzGj/c0aZYnAYdAlYcn0mWQ5bN8IBkAFH+fh9plyeWOSFd
9X7ommZNzZMaEc/kwZiLD6ILzKJWY+K9+o0BzvMvb6ydYkj2fkytfz/8aIyLPUIy
bOqJQPMZ63KKvZykiXdT5fuHx4Ay7SzDrz0etbyUeErDMA84Z1Fsc1gkbMkAodV5
sQP0p8+9VNTX22f2LychhbydW/W2oeUksFGVr78Td64GnNzNxXExMm1BKOdrz8s2
GniC2Jw/T0jFtSc//+GpCKDKJLWCiPTS45dOtXNjNXpAogS+/+jmbWIn4yKFD5F7
TRn+Et6U77VZkaiTEHD8Fdruf7rfV5FFEX668YSM7wYeps5kDI0i5wLO6UkoeiN+
DBCdpAdNwRnrlkWRygQSARtbxX8zPzBhvzPPKpP7kZ86O0wlraPGP8PbI2nGwOL6
yr/AEOmhuiCeG1fqj2/3KzvUAkgAvn7O98G1LB/HJ/UvhFzXKsscX4aRKjcAKqB7
Cr7YgXPrDCFq+eN2ZBfYv+BIugh4KfRh+6IaBuyPgLvFn+jmRpSx/IBbHiulscSZ
SyFoIlptuBeZi7SG8JCvUTY3Ujp6CspcpIENEchIPlVYf7HIUiTSLA/B63AtHkWP
3RMaidSJQp/D18GCGf5yPss5XjRE43bpJkKtrlRidK3/nXsl2BPCinX2T6+RwXez
vDFSwL2mL/Tem3KYFC/bEyQkxSIQUv6PZvs0TQH0qowZRRaL/AiKsuyE1E7VPP2B
hgTTELHKKiF9kiRSPzKQSBZCCG0W81j54Mx1vYNfvbiHLxQ9aFkC6wNyeRrdNYPK
QGJYtZbwcesUANUEdIxgP+AxghEdO/qfQZJmWDfZ//Wzu50DiuQ5rHrXcuVTVe2U
4WOIJPYIqtreo30dPoShRoMSOHuMmAzSkcaPPm/S8VqyUZqQJPoB7E3JOJcP22+F
48W+Conh8LpoROLnDUkSPcDsyQ3L5M8nnZc+6/k9a5tWr6MS7nWgYNX/7bCFLg5y
obEL5iu1bJ/JB21427k8Qov9c2sOAHexPFr1Q1On/wIULClvrnl31DIERxV5sr4z
NC36d15jkF1cEIBE6U4my5BJoeiZPZgGxUfmR7azOd4Fv8+97kzVv2kbFCsoNpXv
lfOWnLHjXjFJ2bLwG+mPP0it0l4lw95y19ZQl9P5E6eErkimEjHJDqqB1HHSY785
zAHSeSKVIA2e15a1xqW1a4ilkz1/5XDB+HJnmwpExP+N7zj59Ch07SMID09kJd9k
YSOMrU0M7USTc1N2tW4fYT1otlKynPgg2caq4tXq+wtyrhA4F1IGwUpyFg/Bb+8r
MeqwWW7kovhbr5lyoApma15tI65KMWAukO5N06AFMBujNakLlTCVXxR+xPSqcRh0
UO8wEl2Yisqeuky/G+qNrulByQQuG2rs5nnVki8U+2HVzn9oMivLz6WmttdsOKOy
3gmwJTNFbgEmOLkkhFOVt1BpDG4CQ1IfJ1l1G5aOFRdW6yHzuK4MbxEg8/iT74Gi
60dWPix7x/50Qo2kmC2TWHeghDZTb34rKr+GU9wbG8kJtPP2WHYxwu0Kyr73at/8
oF0JU4pHtae22y2aZXPZowWD5k/0RL7gqrfhWAQEPNgxgxLYpeKX2/sTU6s4MZBB
+Vn4K4jmPXebAwdIfVNso7nocgyrdKk4EMuqZI/XRxNFcepA9EL+Ga4IizCK034U
txgkUspvni7hZyHGYvUWcX6n5e6Y/xHgInM/cNPEn96EsDs6cWi3F/f6u4aGKbEs
8ZMJ1tqBOMCOFiWvuvgb90qXz0DUZCm6GQTAja1MjmLKanhbqc96o1+ecMQfuttj
eJh0n+fL/ankFnDbX7fKvpheCJvpNPu1eBkUOTb5kbktnWbcznlIFSzuHROzmeBh
m5JuTAo10+QHf2RyIJKY9K0EQ0qcebMnkmUEWNlBUIxPdPgEqJ9c743cggNAKuhb
n1E4yLDio7dJ+MV7Jgk6W2+q+cMvvlVOpSuPDFb1p/l4WdhERUwth8wdSUGYc9GP
+3jpM32z7WT2I6zbd6ykZrbnzzJ7Ew6I72bSTok7J5HlJxEUg4TBP9h3GAtj6y8O
Ipa3/znn9V0vboRWi0rBnBK2XECY5k0Uy1ASi4VgA8eOnJ7isDE3ciY09mvYFtP9
iq/lfBI8q1EhVHWCS8fCR6xSbK8YqDo2Uk7pv+Jd4N4LjHCD0Dxn8DNjuEPV3VP9
43o0bbHH5Fp48Dx1AZA5a7wJuI+KX+OvQ4apGh0/gq6jbMTfPtGI0SNzky8+Eol1
Hb6stoHhiyl0HnQ9TL23KNje0WR9Hv+E6dv2SKXajEZ7pczIeHMMna/aLD7KQJSb
LxkXf0Eursb9/4iXax58t9etQYzYO4DuIa/LaflUaBCsxNKloKtquq5vcB1EQqHt
acxD130wEBElToPPNe0LWFsg/EYXHL1CjV0GSlxRtwwqz9n4xJrd0XVRnGMbjhOS
5t89BuBtv8bmIuMtlPbkfeDEkvTKOhBzb3azvaInkdqzias+3nJVcqQKOPIMGOJn
Ad9iVWYGlm7fWV7YwbP0ROk3bguyLN+VuTXxloTNmRKK4n/7+i0lPtEkcT80DPnA
RxkjWf6h5qsAJ7w2hhW1qDSYsV9JA15tLxRfgSvxFePppicr/Tal63J7bYhxdrBS
sisNoOYfp89g5ha8Y6z8gdNlXQ6XRXtbG4xWnbXOn88IonsAg40ZrhC/m3Yr/Ezh
YX3es/DLdJTvxSo6W8SxNmR+3+2YFviQ4s1ahUTPrc/B3rLZgv0IZrA3CoqpFGqi
SdgaJaZZIHrUFmSbpBMcfJm2tXvBO5nc3B+2Vqm4pxp2bvrwpoqv8tPJy+ZhTrKQ
Y+r1lWZEUuriYG7Q/rIv1ZIdrdSC1fvxtwAc/sdueRoMB+3IBmoJQ4dYqhf+4yJy
mPozEjcSt1b4iwWePB/Fsw0W/UbBQxhKfKrvlgiFteR+Z+V50XtM4kctn3Sx+//g
cZbqNrRHtlxJVRUaS1LU5uzgJ2TbjjGm4vaQjl/dLpS1K5l/06nTUqi/IRiL+37Q
vccslKoTUT8h/429Uynhqw9wdkw1FOH6RVwD+uT6tzQmQzD5grR7JrQwtV9cqchg
GjhpegBlad1WwMTgRXfT+WZDUCUL/3cCac3n0JdIJA44/tZdZRP6ZG8arPagnVFZ
+UZaVWhCCC/WZjl4WfVbdVWOJtagUlFidbaqgiZJTZyMaCSmRCHHu672Ta6ZQjIf
HN55vXZU6jE+N+qvOhpF4Y6v9edcpxx5/aldjBbltYXtE2fPCNSiTRLFc8mof7Dq
Xm30WrCHc+xNJaNlmEYsgKqMk/3jVyf3eOUy7S8bw5abfK+qlgiV35Puy0TtYWCx
H6Uk4ErUoZKCWLllGyoL5VIX4+Le6q6TkKguHKjiR6QiqljhybqmmOIXlnipypUe
NPU8blVO9Uquwuk7utXJwX7HRO+LW6MUM+zXHdbqWIxO3eDnyip/KRVk8gFl/K4f
yHAdWMkkXTcMEibOk95+rEYS7PyFKcKqahaje1U34tpqzZUM80CZYcR7++Tp1XkY
9eElybPXSeXJas8V4FbKcKmqYHTNTQa9k2ug1ywZsnq67ltvsPGPexx6VJ5wpk+m
yd/YnXXKtqFwVgdZBcKPfs/kJgC+/rq231sy32RetKkAWbmZs/PopYVondK0kdmr
NJHoHhsIemJaoAUw2ilPTZ41nSzBX7g8srBJihQpgqynwYK18ToWbsGNqMwhRO+i
DtKvDYT5L4zzXKETLzbMP1D2VddHgZA+S5va4eCHl9GbnaMd6l8s+T3vcxc68jhr
CsyJ4YOEXJLvPRCrqsrsOy1moDio8MzQLIKV92vmGdoYh7TeeuQKTdgaAXgS3b6w
PCF5wrvHCtPMb7Fxj6G2Gid8DB9zEUPFnXie1TL8kCq20p+hBfdE/SakN+1nOp5r
A0DXh+fkbAW1OrPOVAn1CGai0mGCz7cN/qr7nfC616lwsvW7n32gsMN4BvT+LZdl
nZ18G/NPJlOqJMR88sBlcihTlSAzYLU0BcWYIkBG/S+aa6nLLol2JGcscMv6MXql
WxxFc/UoeX18AJyaGtT3X6BoxO511w5W0cXzUA/RsWOnM5PFXBQmC06BebDhETQb
6ZGDGEO7SqBmy+ErmyTnoPEjCLWOQ3yuzYd5m9Q75bMEOeIzAV1b6cD+HUAk/2Sn
BNVaT3/pzDDLnwnoujgX9mrcyCeZjHb9hqhaqy3FoAB330BTMQFDLaJWr2yW3hyj
ES49G6zztrITFEVURXc5Rx8SFxkAhsZNcfRCb5q5nphSdgJ7ybNbarMg3jj2CHT8
NKX9NkmXn+QIkuSZ5zyX3eP0FS6o40FY+6UIR0bA1ZF8P/V7N3+ZbxvTJGTD2CfO
ZBmp+lK63Esflt8rJMOSfeWJveLBCa37U90RrkhUtpk/zWY4Y27VC/ms8OEcvmiM
+KJj4e/Uc54FZQ7FcVs0rBd/+qk2z8uAHlpNdk211GoaVuDUZXbelIxTlvzGKEnR
lB4GNAxvFyk4u5yMRFjE2u6uj3mKvttbp8rT7f+BxJ25OAoMlEt6FsLIfBbnVkx1
pW3lxifq5DqSKK4n67VHXxQ3xXkW/F223ZF61uhsdir/fAs/8sgcEz0tYEr7syUO
Rml0nq0LfMmk9yaL3y1Ky9Td2Rwdl1DthrWvYcErxTvUq9HId1stuM7UV1gb8FMk
H8kTx7KPKDPIXkPseCkn34tllp8e4ARNNMOPJDksTB9mm+5kyLbaG+o2cyt4Mm+t
dUDsfAjV6JXwX4YCHnfFBw38w4/XTrr2kMTOO+yMWyvS/FsRmMW7IcQ2V6pL/D9b
tVDH3OyqqbY41dV/FmPm4ojHlx59iom3i85vFsQNbrb46XuSOvfk4l6rz8xgpILG
3+np+eXHM6vLsnAap3v8waRkNJMtnRAwugQJFcHoFZewWI/dBK8mmVGc+TT588Fw
Hhe+ycnVQ/f9pzwwi7g26oJgOHs1wGnQ7h01wQ64mA//p2r+WplerSYgjMIihPKS
tXE5uez/0zRCNT1Qn6qlajOp6v7FyRBba4WdsPaBtMM/rt9tvpediU1DklzqfX5m
T+8dXLpIIDeGo4lBzclr5Q2HGAjOau4SlTkDjENpse45KGdUu04Xle9jJPlFsZ4N
FVhrlVT57sbAa0zK1CP+t/FoBrpegxphGCSjhUZsl8KwI4bTucTmqXEiRYlz9Jmo
fFO7tg2NQHKu3yW3YcMFGlVAAQu92nrLKGupmDdMGF1X+cSGm+LoR4QC9IX6Unb2
Yk+GsCy6EMkdV6iOMubY1b5OWfuiExR2sMc3zvyJQwGZ1sjareuLl/xomPt2o46b
/33x9jIh1OwubPKE31Hk+rZBtRLZaEZUGmV+A0VdsiHdUNINy7IkjvfD4sJL19Ex
MOM32knuER7IwZZXHPdTE7WgijeE9xLeoDsn/dH3JYNGwBrEwq0rh/s2LjSztwgL
BnRGl+LAP8vA6XiI7uLTabZtn6Z/0LPE0w0DUq9VnGYGj27nICcDIapeJIi0FLW2
RAdD6w9zmg9L5cvMODuPD/zA51u3H810CRabjLF4W6TxSG/jlWoj3qc5bISo957y
VcjiyH3mlFIULUE9y+irA3bar+Jd+zkK7AMNsikhzQe4AZFGIG4PUaC1EDAm+rJB
wM1FbA+hLwozNDkIAUWSsj4Mc2Tcp5zaUedVb0W0rp8GERotkOa+lpzu8Luv5OQZ
j/cmwvqwzmFcKjKTPiLENxShW+v6YzovRej8dsoCG/WJF/+yQ1GXBhELhemYuEMg
nRRg200SVuYFsIV3n73PIpjc+IYuPMjHvNaPpCqnVTiLRXQ2vyf73P3ZSgS+/4BW
KR/pyHBTS0gUxy+wPrla/gR6H1WUhaXT7abLv2Ihqad5I6RnYI/m2MGBY0MLU0sS
g1lh+Dq4Rg7hqXAKKuKX/Oft/BSciYLKEbkDDYdNFzi7XGVVXavCCHdgj7zTRBQG
ANYQDUzRPzzFpps5Ej3DSNULBa3KAYPtspvUKc0ejOpGHUCMXgIXjXNULkeUhsVW
tSo2DJ2duKh9pIgcsEghYo+8AU4/wBWOz3gm6JfVXRDAZyoCeazFBIbKWTsCcefp
c1yoVBkWY2Gg9KojcrtGYbjBPINHhojWcE3O47CzzRFE3QDladJvbYCoNEIUIsqB
zQzPgqG0TtGcvilM0E+8cafkf2G6PcwHAu8lAQB2yaxNncbBOlnG+wQTmMkrwPyn
jeg6ba5uVdRFqXU4JW92CxLDQX2TYVe9w2JQXQ15TZsW0ftVJkb0jFbnaLokmtjH
DnWRs4r5KQcQVq2vCyfo5uv4KapCwWne3k9/qyudXqTMoeOp6VFZ6aGc+YWwysAF
TzJKL6jBNGBrQmGDaP3sN/Q15DTSWeHE4jSNyN1FGZGndN2pWmU18Spz6d5enQPT
dg4xq4FPOjWCpRhxdSwfN2F7480BKDyZd353MStyeRZTQbj/f32WByRehc/jMfZD
35+n56seGQlSQBK4oc7ky+v+JVjztd39k7rpP+SH+mtGWF1BGeS1/L/IZ8F1NU5f
McOIXhvdAa/Z0XMb/Uuhx20uRzLDKhM771ANfNBlXJS0lbDq4I+e6EgLNdHwF0p0
IdMMMcmd8w2smz029yaQiuSWgn4ohPlaN6zsxmB97XV1+lKTK/23hQFJbKW5K+F2
gUmrnyMYS0W5Nl7Q5+RR0Aa5z1xwP/bLQJcSatyAkMLK1j6EIbYdBmrQVRSRQVin
Z2BG2Ic1bcw/mgmWMOlKRIuyvxrZaRJd47pW+gZyVPLeZfsKI3F5SuRNwhDEC896
3jazjeb2sWwsRU9800GUjo89oXeE+s3Qk5F/64kcVrLEUVWWdnL8PwDL+y4YFMKb
I/fP0tNWySC6drtcoh339K7Bxdw4WjfpiZA4PJtfqplwA6E/G+zlTufoC62EvAJ6
hKFCjoubeCsPdhy5Fqy2RrtrxVG/h/utD/8ztvFlCWI8Pd1wKfz/VTfQC7D6BS41
PWQwv1i3brfkmsYgUVHnZaEf9FIiVLuXwl7F1Yan5zk4SOpwpOugO4dFwJV+bfqY
SeSuF//w+1ve8zbHUB+hbgtoXBRMG1fAdFWGfuOXRq2Lzu88R+mry7WBNVbD8HKn
/xyg4ucFVu0O+lVUQkRqJ1ldriRwVhdz1S39uIifSUJhuniMbThzyuFENpuTgRGg
7Pn0auZ6LxwdpeMTXTBZNSIALk4Gw0ehDSPJXE5F64fFelXzsf7PH3lHaXBbudzl
/fkC21PXH0kO9/7ZmMAAWEKDo2FUmyeLugrqcUM302vZJkJDiyxOl3ZSje8rjOh4
as5L+2BdrtoT3ei5cz/3Zf49BqRqNJEfrxVTAk8oF7ffxeCZhODAu4f3BsFsZgmP
KSfbJA0lsrleDzf7apr+CPh1ntq/7xxnQNG55o+pSkGbNjcPSJXb9UYyyWibot2j
w5w+k9cHC0bgizer6Wm/7EGyCvMq3B2uiQ7YPZOuHXYFZZSdcFkMcRizhJdYgTLZ
tI+NyL9fNXVnjiO0nPAqL27Vpoqrx8GwncPsahLnCzLBLMvV9bbyCq+zU7ns4B8E
CL7gdXfkp0feClWQAzYoBYzclvvWtf2EU084oEGWOwmGlbPwyOmRmS0NF5WAwGkX
g5A9kKfyWsO2n5K0Vh/p45mofdBvepkwCR3VqIysBv6uKdNEtlPflrRZwmL5F13D
x+nazBIgFm7MLUeQQdJ1PSh6f44fw9XJjgWDnMSapcn0ZALvQDrnPvNx7Cg/iKsR
MchCdNEup8Fl7HvjsuL3eR/Ku0gsREKxnemDK/Bmwk3hfHC+BWBvMPLid7MlVRhd
bHPLwTsYMZvBQtpURBODy5MQjKLoBPd6Z+24bwVuTCqFG6dpSRH5ywJdOk1ImMLZ
R/SemazQCE9ZVCFdqUYTatF076GoluTj2T8r5SUY222vKPV+ZROKbg4zHbD1bOrC
SyZHlL7pKOt4MXCqHl3C1nPePFnShduQv2mV23aZC2be9D0Uu9wpXlSzF1XtHveq
WSj6Rp77uh0BgEAzQcEgWDDuF/Aaug+v6/h0WS7KaNFb0xYtFrzsHjZEeZkNR02i
8VFhLgEClmDq0jXQnodb/TGf/Y7NHIRQGcWoOkpS97XjNVeiZKtG9USya1P9ppeX
5SieRity0jj0xGArhz3wV9dlCZ01l8j7ALYjLF3V4QysKxRJb1UnwICX6GvSW6YE
jEAE8T7bPrwsxthS5m1VKWgHy/FeEvsYrxn/nNmXjsXGX5zc2oXaqHQdNIfTTYrG
Kd3fm0KxuVjwOUiE9S4WeRanzSX55+J9QtJYnTmWvujiVTuPV2DYbxv7KbhxPbDe
bGoToFDMxfQen/vRFwsZilL8vos4Yzi6SnsgQyWSMXKk/zafgbzP9htCIxc9jOFw
wK2cPVfTeOJ6F7Vmsh0KkG5dZmSRuUx/AIA/TATvH5p8tQbTOwsU4Mz3/pxAySqO
INfDReZfQ3hE9TFMqbalvJRr15j/Ntrs42sV4rc4mjAltmt6AbHdvSSD8BM3iSVO
ou6cO+rkqa6kHMhgKMOQmX4OjXX2M8wVD13NlhYv0fQSW8wHv1dIcRkO/WQmaapK
CPgUb+qI+y1qEdvfB2ANrKyg93T4rxmdxk3u9oEDsdJzFav7OhOjkU9xrd33BWxh
oyyVGAwu8aD5jkhObWkoPQU4/iJRQ16uiugccIBUisIwGZ3KpN+OUKZVCuf/WZwg
5VObhAzdCyEto8xgZCPiLg1sTRJUfqMNRkJjigUO276HBpx+2/dI3tb8kmphgxKD
RMb5Gx4me5IKi9s4Id79491m0DoWReyXdMMu3S4agpCn+Agj8pXGUh8kwguYrrom
mnTJG0EsS1pg4S50SSKDo/mDXrfva8lZbFMxY0RNMzdlyzJ3g0z5aEvQ+yD5/25j
mn4Zc82cw7jDloG+leaUuX9bZ9PBOnqSZ597HGg9YciYu/MEwNTq9DluT0zvf/+D
4kzCHaprKGT/hsxRMm87rwNrvffGFoyqYb4+WmeQuCet85gE5lCETIB5XxXU2vKP
pKtpEKLUgNFgyDkVN6VsH6Tp4b+mlxapoM86O2xTYUFW2pcvCPiIjii8DtBAnTIE
1TvpWbpilr5nxxf9W6ynRjUd0KGmdQraU2VtF0VgvjYb6IcwUYJ+54XL0CI0tE+N
7k9uuPW9fTJ23HgvAvN3bSZkn6VJyHJf4GII2ggSdd9aRlMYfbSR+E1jS7AszjFw
6vn07fJYyIJhVrRXMyL+ymxr7NFeVGleGUed3CTWsWqmSG0IAJQA/gFmhKUEd3nK
D/LfVe5uI30gMlosoo/NJl5JDePGp67dMxCYuzcENFK4tztgg1p6PNJxMXnQY54u
VnUee+TpmuRkVYFxSxmV6TgJwK+OObS3LbhpbFJ/Er2K7YV/FTJuBwV6zbkrAMqv
bTYa9X3IQc+1QGvGgPxozZaobqRxRlDe1Q0GmeBzN4u1wmhVznRdObqXVKT1vjIu
WitSQPGgwx+fJ722kKNsPAsoAE3S1+DR8DhKoFRZTJ9S7vjrYEP5suGoGHC9kBCQ
W8Q8gRVidFB3BR1cBjbr7Vw0cCKAc6Rq7ZmzTwyoDPtVPPgkXXBetgloqw3wbTl3
UIN4FRaT+CZljbujmTRFwBvebudN9KlyesdhlKHP+/ZVxtwWFIlZtOLYlOXPW2Qp
9PkyaLwOPR2mlHJUu404/6GVCKRj3ujS7583bFwa/Q+ovCUL75OfrGqY+cTXzb6A
1poP4YJYK6tJRaJ3OzrNOo6n9dyJsPtZfcntYFZKWtQMJgdcJt40NEsq6Wrrf5Ks
yfjRZL+PuulIaF0XqkXZFCzZstUq6djTjf5GFftj+KxaFSsb3GCZAtZLa8vPxw54
BoOTwof5+shptkNBa9g8S9+3NZEoSyiFpsCsrSqOYTfdWL3Azhz9sXddFw3Gv8f2
3HUT/4wUPpu8Mqj+pqK9KhlLb5/AqyjOpSFRjXWcID8VORfSZTPZindsQmNNvKX4
6ZOA5jAIHkLyqwj+YE6Q/na5gzMjShDeBOpFdHnwk8XfX1vBeYVxZfWT61b0VWu6
wINP1w7nNFMSDL4gs/2hfQRZ+uUSNWTHVgEzk/ZF69Piw/OwtudPFLnfMZKivOPO
smW407+VEAfY5J0LQqHuP+oMy06o1rBDPgMO9zfs0ZD2im0DuHc2FPPmRlfVaH8S
4wWmNbGE59tk6/DwfrbtalwS/Os1RvLGmPiL03Vdzn88djrOozJQzhgCSWEOTVgU
Ti5yTcsqI0ADkH0GpyS2uajNmCfmu+8jMr2lYmIIFcp4vsD6ekCdnYsFPJrNkYFl
HHsKiVBmhEm2fm/WWrtxCjLoeBo4fkmrC5T4tuIgpdQiIe5/LLjVZqal23PdJRNW
XrmKYXFmYM+aeL0WBWPr95cqkQY73jNGRM+SRDgIgGTlbRwzHt+jqjArJN8d7uOH
LVkh+rMCfSFy6DowJv9T99nGV3SUk2VbNvPV5DRunLY34/tLS0U0vl4iDU5Redn4
++D0g5tQj3DwVf9a7HRfs7GU/X8Ukd0Eo79n2aVG8gGaRuG/XI7aDCOdIA/54M/+
LzBrC2PkNChhPjDUMAHXx6xxn7kjMy5DEraxHNieuavT7Zaez0jvJohCo1GyK0IN
Pf6e5wKkimUS13G8LhHY2bE0yNARPwiCLjuM6uoWMRFZn/IrgUuCkWmR4kOUGOXE
2jGsN9urFyOuk2mg/jIi6aW6hxYoasMwwZk1H50fSLynFNWIrHOMqcSNAjNyo319
mOaLscF1n820fn8r4dpDvCjjwsE8a6Ivcc2stc/Pb/UOevpyAUS46YbyTzMtCrtN
vCjg3+uxnJ1Mk2F1GHjAylhJsfXZw7KQcODk8npgh8cnGAR8eUkHNkogx3BusKT1
8JnXxSPfgRL+GU5bCBcUgO2UPup7M3EmghHTPu1qS3qYsa1eSQ1N/ZjgBFoIoURR
mhaw9rweCCIGL1tvyY1XYuvmmCtPdYGmW09ms+5sp1FlC5j0LyFA0iDoA7eJ5JGI
lza5wlVtuZWI9MSOsbO67WQzfUWR3ehEb1e6SgB/R99D/bwxz5xI8UFAfsxurlxC
fZcmUzn3xEhV/0H9FGrj2sufLc8vWjxcq5E1kuMWSgnOf8a8kKvcpCGNftJ8gJL9
HiMYgxgtITm7Iq2J83AwhiEDQoyZ+AyCGpGbUGIbQLUT2ytfnxs8y5ADCv2zHwu2
iADDh2bAsuZnRsakjJJMsD9ZneJYlm7BZ0qzm2z7xblQn6qA/qVMrpSPlWWSuucR
LTvJ9Auu7l1Amdp1N99g3W8JT8UOSIGECFlICikCGT4IfdYPbsbXNPoMKHTSBb31
Iw+1nQO3zcEJ466wSqnOiJRl5jWCFXXzfof5KrFdOf4qzZ6WAWV22u9P9PMjV7DI
yL5wes/woyNgmtvoHvENlsW5AedXQcoBaw+EWmZZz2S64tDdqGn9/vUDkLMg9aJp
8nSyPWin6k4WcOM6UXgs6magRiH85Pqfh7tqhZb4tAsL0rg7PBQ8W3Sdf+9gKQTa
HLTQPyIwmGOi04E12smMGQiXtmm0d4BAWVQz1QM6RdhZUbGbGt9PpROHyLtstmMa
P8mAohakrzhBqMAly/nQEjPte69ftIm1p/EenQcBdzuAAj0JSYZH2DKqRaC4ZIoX
M686J3acURhs0VqFUmWBUatavRjHUpjxqWbMvX5UYFmDmdoDjLVsHNE8HOwo2xPz
qr7d35hsXtI56v9V68/sZ1W2jZK52BFHDYI3ENzSlQ/Phm19HooPIjqo5vbYYzWx
gTjACSCN5CUhziWi0TeeX+VDUIhVTRR3+RbEcIl6pQzs5xgasjkIXMAmXFp8fXZa
UVD9kiNDmuZoqoYG5rTGLk4kn2OF5SmXdGamrXiss21O/sJZwJ/5P83RoB2+KGav
d2hA8O3nNzQUcxyt4lh2IKb1JSaSKpnJTuzmcJlH6bAdGylTDJ4B3ca5RIq3AXlK
nLkQNKbjInKEioh/AH4K+MGBMNJsreqHAAg5nIh8lIZzzNQ32LuLYl8H7JOyVCcp
+1m43vCgCD9GDzTWSygquecWr/B1Dz577Z6m/x60Ca5u/671plTAaqJkeZgS5DT+
7EMLR3EvkZwCkrX644LwWiOmbX/0+Agc/IuNgTJmKMDN8gnYXSqJYH9C/qOkkU+X
1RCuHVbtB/46Pkj4iST6n+xFbltrn0dKiM5EC+P9JbWpWFbzZ3rBr6qpyTVnLhVI
DiFTp3lm07OnbHxFXVDmkmp8Mp053fTi89RVmd6YKd1QJ5Hj8fxDtB870e4WsaB2
zAZhITOzztgxNSCUT+LhxEkcwS2pk4VbP2/VBf+dAy3N6DKGW9yYCHT259zEw+22
yITXwEXEv2VeJAZn/41nRq558IHzUtWk+O53VKzVAlO/yZs31euda7a2ZcaoVVo7
MPeM9spIiyCd7pg18PeBGr04147GK5vIyleDidq6v3H9d1v+MFIFqiS/jfmXB2lV
ZsZij/PModCvkzISth/qp3qWKbQTTw9VZSijb64r1qhZCR9xyjOaCdh4uPvGNh7w
DRzh37xX2/DbZ3/R/5EtgSnT9Q+Es+WYwGigU9TNOHjK/xM74FfnSd0WYCRGnyfk
uGG3qvTSrPWn6XhFmWM4vFug42u+8FOMmkbcUAB2c16NTGWN1QaLc9sCof8nYUqG
A6EcDoGIFADPgX7eLNRYAFZ7NHSGBohRQTwrrINh3j1ipRbN8C9St0QYOFidqf4J
VrJlP52Ig3jN//4l5yWfU2l/PUuDFlMlPgynFBY+5USOBxTPgwnIqz9iw9G+e3Wq
yalM8qH4cqrdAswymN7M/6giZK963JF2ISvJ4PNev7LjGfACMF0Sf23lgL0yOd+t
hKzPMFkW59ZqQ3SM7BkbW4wmiuwwWhkRXHUi/RCMWG0zhcVtGpAziDS1V3W2KkBa
jEAqbgMoidCwOrOKqIzjWUUBQDpdpCbn6PT4JfnmgLTypLHOklY0OqjAd2T+mAF7
pB9BkE+ysfqveYRiOjGxaWfOclPj0EqwSaoEdR0IxN3ZFa4Yl62sBQ4k1eVYnvur
JfBXUvLIRmKpOB8AFva3RPsApShEcfxP31f68E3ZwhKg6tXqxdpzUkuvbN/42OfU
fcpWFkNNETG0VXAABAQWsd/QDff1e02VJeme1rMy7UWqrPjQCGH8t19g/+4JxyD0
t0BlSUvZ/8fdEZP8JS4feNL9y6V/4PeQ0ADU7+jY2UFfu73BkmB/JPXib6CfX3me
UcZABE7pTHu6T5eEUmXqxituuN4Nl+kbADunrBWoA0Pl7sAHEPFPaU2BM0Z8yORK
jeNTK0UaaAS78C2m2D18Zl5sIo2NlCTj7s15qfB4XveVbS+Sdtu0Y30DzVyXjEva
4pOHpWQT2XLf4zyLktWxMEk+c+xkP8NYNLijSWTdhxR22gKDV8pAGOmtwYjy7F5J
hfJ44Q7TpQ0qqV23mSFcFupBb4kRNixtih9VXmwfxnLEWUCKKJVdnz8ti4OUvR5s
ydCIiNcWugOY3NlcaqerRFviNA5HSX36odk+sOLPoKL9s1S7m3SEGegOJ/Z+C/Om
v65SmzdQ7g16VVnPbVBvkGiIk4IhhT4FfXJzRqn0519/veRBnRR6bXnvnQnXS6IY
pUKVvnj93LPJmjVsOh8QV51s6uZ0qLftj7aCKCmIzMQTYuJgCFuJQukmG5vKAYzV
SRYLdMnJm4zCC1hKqIhS1IXESU4IdKztyU4MNo5JwrwDLKbHlEAtZcNBJx663oDi
GtamtKmn3Ih8iDyYOCrnbXWOtqskFmJ5es6Kg51bOKHm3xx25ei/UebFoDVzbNf6
fmME3LgPKA1RT28uujBvleSkS3V1Q074OiGwwEgxuiQ5BBxwGDqLta1ydpmKrdhd
rwEIUa8dCWVfnk5OCua0u0j97CnWzH5NPgF/ECtWwYqQpt6+7QQ7LDvjitEt7cu7
G1nO3Kifbxbr4CUfpN7tSdV+JcyYynAvwAgj4z7+28Uv7+5ZbATg7FwwbXCI3hR1
pDVoCnwhgCRWoZszgxaiNZAFenv5P/oFUpniRz66IIrIsH+7EoAtNc7dBhu9f6Na
qC6e6ACOD0HRvzZKsoww6xgnycuR43YgtSHdc5KQxWOOXWi/Owam+2xlz4oMvNkd
ZdoXqT/D5BfsqJYV/o8bW87O3X16IuOBG+di6UbhvdN2/BOQWxFWV7u1lXyetdyc
vBOPeTe8q+QKb30meZ1SXxhurL8bbJ0h/9fXP8hjWdS5iJMEke6ypjCFGGwhygar
tPpPwaQdixQ0Unvb08PYAnhEbY18IE2CIkXjCS+cVVGvQsoWvBl48UmJfyIdALCv
+NrJfqd5qisoI2i9EES0HtsCbPj8+741T6HvTc2Mqy6rcoptnTy+HCOlsyHZ9DtD
LepUH3qVsIQ7jUkODdCgeGquWUjYxh0u0QKYDAMHQmNyaZQdA2U7SRc0ZlWK+UEu
iNWqS4gEFZJj18xHiwEh+OKqs53ais3XtfMCKyuCyg4f2SbpjhopxCNISkyLrG04
zEbJIwj0SbXhhhMTiLsLv/RGf1z4pcBUzQhSsrZuJ7ek6r4sIKLj6A2WJ4E/mIJc
+1Q909mT68VLwDllox0sVC2zi+qmZW89Z1kFO76/0jAqhhHCa++Jg1n541ygvoa8
2F8OENh0sX+GyS6SljUdh6fnhhY4ZwrZWjVZZxTvYkmH374Oa7M/zBmZ5RxlC0iu
rsG92f/CGooL8iRLBYFLhjji0otxH9TaO2p2WZOe1asK/ni9TWbqHwdymI+N5qhp
zkFlX/V0y5wcCNXWzN4SyOSEmsgA2iiwL6bJRudL0JIc6oPFjkQ64Pz3RZeN/9j7
Pqcue/PWEfP/88Y9zLGSG6TSn0JzDDTYnpiyzo+W80gHWY4+isHwX/hy8Re2pVac
CIdJv73fJYXq8GcLuaOvGJzBXjSa+U7pRN8Mp7zy+L2zsqUxndbAtim8F8E2wm/A
VfXat8uSeNN+z2NCxEXweU8tZgebiLNM44+k+vL7w7ZCDMrjwrl9U6MCpdmYg3vx
46cgiWTS4gHjwaJokmzGO933Irsc97xZssNWIXBdwJ5JClpRAqVg0FaRwZid/Z3V
pqFimPIqSIzUfjol5xwr7K/wBbEa207/DJ5q+44y98S3GBmvqo+7qg94jpjexzPp
BfYy2pw9BrUnpCeignZzd/atj8qkHidJ5s7eDh+GierjWVedtMFogpD4TygURYr7
Rbx1xpM8KA99iXXWDH+epDGjpFslCjv3rp2mg/+JxpaLYQgmiPJaYJ46HM2i+of/
7khN8Z/+rVLMqlr6w+uJrA5tFWT043HL6hy8iD7nlpnOPCq1AvLFj8TcNsSYeJmd
vme4P5eR4rxpDFFD2V/5BKg8t/aPXcIWS0R4uHosUfv8B2aX/w4i2c+WddWpq7jg
gmWJNZQXTdNDj1lCVBdJ6hG638tvU7zGnf69ARZxErb4NDU47Rt1+u1WCm+mc8Dw
HxsYc3mYLV38DAsIeXCNwWVbXcT3528bKF0qvPhz3t2P3QDQraykNf1D6bpHt+/2
1PggKxYvuvdAJe1Nv26ugF0g7OrjBQ+MCEmhNGnwuZqOlduZGWwzVPXT0BH+S6/K
4lWhqMQpN55FVaAnRaU41L6cIkWYy5gCbkL4097q4BnBD37mWBYb4QUtUvBtDXgl
O0E9CeN1mGxfHqCz277KaZzioABjwKwWq+tYMiMSfnlBneutK4LOo6xTFb8QwW6V
elQAjH4l8qtNgeW7YTglqpdkixzY+sOwryKvJx6q2ebeZQQGsSQjezEDzY8EKb4X
Aohgzb/gDm//TE5HuXjYsckkxoYej72pau66n8F+/ckWGv9HLlaFE7LXTNL73G3N
+OJyJewi1wxbV/B4M4IZK0eEkHo8tx6lo1hwTs9AJzSrwGbn0f1AajKBDPgJre5O
9hPL+Y91WT8Xx3X7MJrzfLDY8AS9wAnb7410BuALXup7QBsiWU478zhh8mQYJqA9
LIT3ZKcTnKY0f5lBjpSqt36/tuXQ7TfuEOxnsP4WzVRvqNBOtT4VGQIQy4KHrZ5H
XZ76csmMMTt5PS5vPwTGMUf7CgIO/6kLaWWgU2J79/xKJCHv6J4RajTG68iBgPbQ
l0xrOxIBEkgfRSkUjqwyI0rQNHNGtdku8sNcO0xcezhYruPzO3rJJflmPhhF2ZtC
Cb8Vpw5SezJ210iDU6734jmr3+Eyx8SNl1hli1dH9rY6GqJkwIQrw0OiuxywI4qM
SZvSuWuPVRHvov+uSKOuOPY3/xoP15WRLMZF8de4tqV3oAVq4I6droUParfZXoqU
96KN1K87gpz/80piaeYSfCgPySAbD+FCCrwrJurwVEycdXAKrRnZSDEbwH7eQqit
2OOXHOhtBOdKqMXbnR566zM1y3r6hkMX3t8R3UW4HOiSj9Q3VfkjL7GGHZmThCvS
DtAPgvbdYIrVRryflouWTozYfr/hFd5Wuz3qOaoZ3A+c7qL/HyWStOli9D4RTZFN
0tqD37i6ilfwPyFUs0QD2ORn+AMZ0mJE7tZNIHGOxJON9DkLaqSzpmsUwieuKHPW
RVdZjof+KI5A8kPxrpW5w6TeIw4+u+wLD3qOhofPfqCQHoS5Fm2nomi8kgtu0xmo
j1txgpfzCw/9xN0fDxemHk79vX12+x28lVFKBzXFLYlkY9t33IndCzBAzXWBV9Si
31i9Jk0reAGe9gdzLpHYT/6wOgHCE6/I3poW8t27HGhDD3eXIZo2sHJUw1cCZZSd
EtrJG4S2ggdSoydlEwRULb1+mWxZETwlb7LOLebPBW99ZH3IlU8eKvazIkuDFqpQ
GeMs0RPt5ahY9Io/CI6ToPmU86zoAK37K2IS9uxg+U2fRh5mSnuVrXd+eMfMInru
oADlkKhOxSAYFw61eUN88tAj89P2bnW9izC+S6p67hVCe4DmQ4w41t3SSdzzXTcL
NFjl344e4TOR2rbAqpsAltEr0FMYrQogbe+qhTMppB+hdpBU+COAMjiOM3BRK2Ta
CBsVD4vkji4bzWcu7cEoZo1nj+3bGABy1cqdlpNVdzOZ9tUGZZLjox5KzG1dTNpW
Eg7au1yQHbkKlrNFthLpysUwfEya12uSRcl0ZpCdg5Bzz6BqzcwdcHYdw6zcVSLX
KeAaeTPv+ke6n+uN0z7dsyD3YecX+pOa+vbIyX1Nm4E4gCcxZ2eNByC0Qdv5uItL
GIcfjm2uNxvSso0EWRCwTZ6eVx1zRhcVzEGlM7DTlStY3bPvGRoVbVRX4dTqCy80
ap1u3Ai8U1OnEbuQfrWF2ybjI2izxlWy7p/J6N9tzItRuSdWqlNW6jRdLgocdo+s
f6q+N1wrNpUKTXFcdR+0vRiQafIRZmBMniJgIQ2HPnRUBEno8kTwzWVABod0maK0
sLIUNzOEzrBpXU1Fzr911qDexdSlY234s4KcsCvo7Mn4MFpXVEOrh66wIddlOKRa
Oq5Uo5Cj780MiZkC0JKe1sQyad6Hlhcz+wdjVxx5ljYpLKKzJh4gBewpfcs5XChD
JDhXQ5lxJkgpwKBeVT3DYtbb7z/P7MbkRcKQXfCtHVS30Z91l8SmP/bFIWzO3AI1
FYs3bd73bgQXx8sb7C/XRtJU4FD7tN0u0ltb/zfczFFx7iGa6cZ8PsCe5by1yZxG
0GsY4wVv3hHgu3hHcgolGuzxJ6P70qL5xj4JqswnVCQvDEKY/pvhykI2uhJnhWHR
WnyfOA4fl42DnSOXm2QtMJUrRApHsmTH/ysOhUD7XMij+/puErSxsPbbKOZ3XHv2
BLeXUpEb5YWZGJt8mtPiWRwshRWHotUEpFa3ahLsQta49RqN4LW1ls8c7N4Ql0rT
JuVPbX2QhpVU4/qDw167uIDuuHU5N6gL47G+aqKNHy56dP2U9HBby9LED7/wHNtX
nmT33LY/YEJJv15AZe/a+4mR1Xkja/+qeC3NQUj/uuIoyFnouWdgvyOjOWlWiZSW
E3Pju8M4+m58P2j1whd7H9M0ip8qtmwGVX+nqOZGmWCl+jjacIAAqipgCY1nft4G
mAya6mkGM+jon8mL5AKN6Of7/SFMX9V1vBvQEpMKy3cbl/JWOpEsWBPyHKgkrocF
HTk1mOKZOQWIzrZ9qesjrPBLlk95OdTN/E8QgyoMlYNERwu2uNlC2s10QmuuvT9y
HI74IScJjdTmodSV1v8mOM5LZCC38xiAmoPkAa1sJob0h5XstE2SsUIfrBu03Duo
xRHWcdWDuxxOL+DdgIcMkvmcMZuozEk35qVYx25LXrV0AIfZjiYmIfJMsYCPw4UP
rzhNkTweF0uslD4yMPXh3HHqdPuJ9Z4yT7L30JPasTGuK7kvUbZsN4HCdxVfjJIW
JgWgoWdQS6FkcyzNS7rRgXDDTqgETqm8y1Qh60QVZMnbCwRxHJioMiPMa1WTsAf5
3EO7l6dCa9IuRC5t0GDvZi4pm8soHIwsaylirQMQQUf0/8RD/OTkUlLd6nwAIKEq
tAWA78SFe3SQ8vQeXcES2W1bjnBe3zVguF0kZGmTvS07ojhMGLG2riI+52wBIDdF
8ecQH1X6RjzYvU9dATP4eZnUkRK429vSGpJvCEX8VxuFoeHWlm2cwC/FI6SfmLjh
ZxGEoITIQf8t/LeZEOi28EfJXDhQmENuu/B1fsQaVg6BT3B9ourvtD4yhnne5f7r
Q+iQNLJNITMfw4YEs1rM7p9L5OD3j5FofUXn+SV2FR2T+Nm5jmF+9uDdPV1F11h2
r2rNZWIHSomegNgUgg23RLdfT56bexeRV6MiAklkW/rby4twQAhF+BkQoej9uwx1
5Rel6L3NQXhn3scToYwM/HjslKXXRrC3V6/ylmTFeZgBx9SU8ZOaJXi3iLSOi2pb
g+D1pEPv17tRZgdhQE6vfNYyaEDuSfj4gWUUBzB5zD+1K1iIHkd8HYwDyWxGcaOa
ud41+8qOTXMRRJz6fiQSjjPbsz1QgXfjBPbfJAzNdpecplv50jpzVcYr7VSYlfVs
XZUD3wdB+0+PlJyIsSdDEHZLZj+tQIfxQQYthRPWZ1vGFoRYl64IJAe+Jf6w/c7e
h0xWL5sbWxW2P8kBwWwyaYadOkRKJzyhKceMKMNOlXCQhK0LXRf2U1xjHb25/3AN
sCS+2Pyw3IacUwMfxZ8Ci8UAaXiHLr9mmSALYNnclmmyBCwQ8Ovsbypsl+6+XUul
uiVzrl1AXM8OXmhGoSnzkoBVCebK6T238+eptHwuzY+96XBE94t/BD9vrXC3llQR
Y5jsGYMpg/Wv/sWLRGJlPVeWB9u3ZEJe863SUWd5F0PbcLAXpQfyYu8Kx/3zGN/E
s1sI7oE6MqLc8/7MNkHWVaRWj5s7DU3YgGchY7ADqJYtG1sVLz6TcCntn7aSTyJe
8tLRfmC47gs6wcP5VHtry6XtqGXSdrNEZ140anNy6Sr7NBvCQZFq/xDvs1jMwBJy
wsFKImc5xgj6RWUUe0RlM+2nawDCJNBgDZlZWOtBKLIHbnw088kvGkVTA2ZjV6SW
MqQqUAknP9WU8PF83yuJsGn5nm5/khwPpIKYKbkfDg3NJpe1+VfW2n848C95VA8R
w1vi20+bCnHYnPvtT2gEwrhykzcUAZWwsGZxLTv59XHZ4kTeOL9z6i4vuVCJxiq6
eXNWzoQQ8TKAUimIUmWtIImcp4hyKfSV4z8fcZkTvOZQ7Z8ZEkiQcmYko7ZcNKMg
HfoTWK+LwUbX6RFmQQFXyvoBIWT9Temfq/X3O/nSrgoyASJDOBHdfpfcVqHRXDxc
vVsYhVyL8M/Oj1GD8qq5kaGsm0omN2+FonqwZbTYgoGQXTKLJyobShbC+l5BYVH9
nBC/6wEJRSbA7A8ClyGM88LW/UbjvkmpAhkGSAAP2E0jbkhvLjhEIjHHxY19hKnI
3759+XmstWtcRs/KN59HBqULvajAdSu5GtgirAuAgbiD7FjnMcP7/P36SsbzqXB9
rhuAC8UpxApBA3uNY+ATVVwyyEBJSiFUqIVF2TM89P/eB0V52Ca+ACF5/fZTT8y0
vSVEdGvfO60+Sw3aEhJ6lbw5YC/kUjRdTXhvEVYZ2cxufcIY+P5maLG4rtg0nvy7
Den+KfRkK2aO3guZY+Wqm4dtlmMznTq5k3+kU1uM9dzEnaH16pVfQ95R770zPkXp
hiF95/RI1dUFbL32Y43RNkchQyy9gNLNxIjKYDbEU5Ff3JbQsmFt7PIdcxtc2Hv+
Ab/YhCWdcKCoMNJnt23VtRHGdgis1nICigO8jbRGcYF+iVju5h8nQKNtaY8H/Y6h
FN6K3WQdLbxW7LhgW3s+tYpxXoqRFQlSTCaD8NzkhSav+jL7YtfGBfxNq5LeC9is
Kky6yjRtGsE/fDZuj/U86QdwM75Ia8Z7RQ9QLUOVnDkRBjhvSKdQMOI18MdwXt8U
CxYvevYJGeEh/WdTAfnRjlhaH5rqhG3tq/W0nskL5lm8JyRxdsXT2+Uet2uNI9ZR
DDdyojc0odgS5rIWDHYKWXnuo4MGwbKpnhKV10wSc4avbkevpHeaYVN3e1DvcW6S
OxnYziDejOLb4XnDFWUc6bqN8On1Mb6FeACXYCaZ89PTR0aFMorCvfDh3VtBxd+Y
6JW/xbEiHCkfGA6CEWDG3PLnNR6mukpptnnRhOelM8fN0GEYgaiKWmI/tPkK2TMN
GV0mLbG6+vAesUfEDoJ0VNkb9L/AoHnjcRVWFKWfTiT0LVCmTC/nkcVpWmMfzPam
wAqHjwQtrLXnzLQjP990/A4GiV8CaJz1rAyIHAohIluCQiNz6Nbt+QC6ObmHWnrv
UEgH9hnT+smHyWQB+IRYjqSS1PCn1vBMmaQF9YMjdKo5Qvy5Cuo9t8Ad5NOSV30k
K60TY25ZAyCmjmCuOYDrVmCf3CRJsE13T+CAIlWOm/EvZX9l5HdrsAnxDwnyz5aM
DGCMaQhKohawsrLxYFYq+R/HjkLugO5lug6RCsec5E50kcNj6FOpgqKayh9IpU3Z
b5x8h7lgRVTBO+r9NMgfHrKa6/U3A02P3TkHYl7PnO22ff/4zJ4bqYdUDsBRVLdv
Nv1+mbtKk4AIYT0oGg2X/mmM24C5i2YVc1jWYOSF+LPzFw8EJLHwyn3LweTEHpnF
ACBea415Qq3W6gl5bRB1Q9v4MiYF53XQjOxN3ZwvagiqrH9sR/B1SsTM3rR6L5o5
Ai6mT8ah2pY9jtkTIFL8Qe+E8fJaIn0CIlewtW9bFlK72zvYhepZMw+0TmWJzWVV
JKT8w7dvOYfMzVLM6IuPxpTo9pWANmGGVbwaYpcxNwy40Y33B1Oy07AyHr7pF2VA
vmTKSj5mShf34E6qzk6DdyyC/7vdwvOrlE7vgsJssajRl7mBzUOqQxe0q3D0ouiy
L/sDwyt9H+abQH6HM9xCm+DLKHbR343xLYnQhzioOeTpO6yEQg6CjvjnuJ5/ijmj
+bSyp17CM8o5vklpwL2rIZtIUmW7SIcxU1CeMTLtxSycZtygnjdLqFhygdXjaXmh
rF4asuDtpn78mUhRjvKfYsL4ROH6xkqgdYdeg+EdtPMaAe3eALniznPXoaVKU/EE
C1MBYTI3DVS4N2kFrkMri8NEz/S3jghuUB4QYq5uAY0QSJwCFkmsm3kC5URPwCPm
5NEA3xaomrOYwa8DRzt2Hk/pBnm+VkcvGtE0jAImKCGc91xaFDl5caWVGLG6NbPe
DP2HcppbfgU3ykEHK5ZZU3Qq430nOI3MW5qvC/jg2/Q20KW7KwzR4UnMuRtxEn3k
Dwy+3B4ddYEJvXLsRdaiZCktCcpi0EjxxBWxUuWC1aCb8dzEAtDWS7/W/e/EbYnQ
vzTaXxvZlvcRsp589+ca8T9yHBuaFN/A7+fxKnmxlI4xoYiBvDQQuL3NN2ebrb7V
x9u6oMGtWAgMNrS/TrExyqnBjXGBTE4Ax4JDhFCRuT+sJ3YS3JsWy14IhS81Ew0h
LeWoAMB02NfLvRzrGUH+vRDLTWPlFL0ivxYeDXCgvg8Hq4CczuVJuHdVP0noJTNr
lCGgRc6z1ljIg8THYbaCwlXtCDzPuid56xgyG4ZuMj1naG2RPiEGq+/0qNA5CPtl
HJuArLBJR5d2YbwQ9tBgNCjM/ZJ5Qivce0uq11u5yX12ID7+V6zSZWGKArWSWznd
nxgj3RjM4GQS6H6epOUywYiNRSBSPlQrk6nFeMokw7p0ECvc10QaFHOVmBF18BEW
8Y0IjnrfOYHi9FbWxde5ovJsLUsjTwbtX346Wpt5tFl6x1U8lFRZThOlObK3tNpU
phYM4bq30QEyDi2nEaTUIPt7VQtQmzzR/7VtC4ldH4qbFcIZSa+V4Q9AzmDuGYEi
ZwbfDTC+x4qjHqbQP33DGoPGhKCumP1qtXtbQOCGyTKthVo0NEKmtvPvkqcudqv0
vl2onQCfnV9Cu+tduj3JCh2pnVsNeOdGVdhhI5443HrY1mF+r9vX0MvcIMz8WSCz
E8IXigL91MGK19rAaf0e/qmFofeAi/CiXACwyBYwdApsREk9rfp6CbyZCIDOMhEt
uVttAL+XA1mL8/8ADmDp+eDrIt0QVJO1t8vGd+KMOYWbLbMr7kvTQH4Us/xKLTFm
fZNJZrOAoeiKQAdLTx/4kCnJ1rKyrChrElTPkZt1A9kXNgGGHbl34S1ptVSnAhe9
1XKj9FCznR2regyWiPm+5MsHDwOVcFEQkxO9E5pllrEUSfr56jvFMVHwOH+gzIAr
rzD2s6i3lzSEkRnCGujZx75MBiqlWdd09YRDylS4GUr07hCaEZ4tyUdtszNk93dr
cydcGGDcGkGGKexQep9eWyQjYbMyYIdudmE0bOmsl5VOn9RqFAtWwzZC2rrwyqpm
V8/OhSB2hqpTmrEplsIJNB2J0/tB2O/dEBUADwRTWV5Q+Q/sARpo8q5M2eX1OfAv
1e/cj1iZsXjWETj3q3knjx+ZbhjKVxOXA8sr0q11Cn79ucDpXwsSWhzRGThLv4q+
0MsZ+VzV9sx6wrXyQcgYZZXGNRapYiSG1tqXoE+5YyhyyWMwUW4+nlythi5BNEcG
hJZp3kfCRDB6Pxs7DclRgvvP40/zkXlpn2MfcJUKOOlFclV4W3MFVPmfLXvHyVuB
BxV4Iajvgjh8lTvjiBE5Nk1HQp4X5PgKsUaPAOeS/cf+7zQAYcAEzJzlgC5vJ8He
iqpOWeWUWbQ8uiOFZAOsgmk0Ek/qdnFhvn9xwXZ6XgV7F4QLXQqm7lwd/04/fJ8o
Uf6UtHVJanpOxbSep/7LK0HfFb6Va0+ZDiECYXQ1PiMIPJIkp4hh7VsXMfEA1Bw7
SeZo6hV6tViFOzQK8HFyHTETgsZ2tNokiyYacEFQgwZ0YYpJn2TblqWtAw/ct2Ec
DIuDoaj7hXpDmOXpIJLxdxF82V2rSUoKyQvjLCUicFOkAbnVCOD31r0UpqaFqIXn
aO3gnBCEuq3Bqgn/N3mLuZWQErtxGPMyjTeqoXZqsAVUMUdqms+PQma4Df9+RGv0
mRUjPs9Aw+hgVNgeDqOg9NgoHsQNh5YEpl5uN2Nk8doszc4LAeo+IvVFBLFpyPYY
BPTxKXnfiF1+ZS+PLCendohiIYpXEFRGGxOBgcDmXH9pNMA5MxUrEiHqi57Ne49E
wcmT9KEhMhl3bc8aqNzrfhxMd7ZOgAYFqTVpCZEk+umqdI6Uui9SB4K7Awt/Yczq
5IEsApitPq3oBIjxm7a15Z835FgkiFHkq4xD6/SDxfSfwIsXhwqon7JJ8wR9utoI
fkc2qAMlMlGmuGUL+7BnjRhnJrR9nqFWXnRQhlk/B1AzcUTs4p+MjElM8gl7/xAw
0JSj4oRHiUO3sO5M2itr1KUuh4FoO3Rut/Jh3DTr9nupLxoYKAJQn5lYlqaRl5JH
D0zhscFML6VxrlIDgZUV4T4X7/VgQLQouSLQARgrIuy+/QiOdQLBBVTrEfTcfLx+
M+4aLn9TNwrFVHPkO1J/zYZrbEUeQhQlWoEsTGjBZ9u9ahj4CY7ScgGzFF4lwY2S
MpokZispC0wEPsDLTRVE9LjVW5dNqTAvFg7s0ssO/pi3Ri6JjmbEcUMOunpHbvkP
kAprFgzrw6FkVly0mNidvrxHDKHN2txCUNN/iofBsWI37kn8C00zpqahyNjiIqR4
QuD/s73/0o8vhyA+wT824B4E1bQGChtQ53RkyuqbsDGnsYdYPfUOkLmSY8efv0Nw
F/YGBIbINsJ+/5KFGuqNYyw1QtipoW6M0Y3r294xSwWfbi9Dh/6NTuMp7m/UK+zH
TupBYYM5zpXIJj/uhOY6Zb99b4egtFJDB53kNB2LVYpD4tHg8MV07MHfH9OQ02IR
ni60fp+jUk0NHOiUom9YWdcI6oCqzg7DMMMjmMFTjPw1hKUyulS9ZEwIb3q3E0vx
yudv5WHZd8+VzOO6nFBPEAGHfkFy0yi1W2I77dYHY5iIHsrocMbZuP2Xyrh7+qY8
1RBtznxVM/sZPwukbFjhmhxa+VmGEZs7yG1E7HVzJQ+2KEb6gGpRCAqTnS40yoIZ
Nmc5RCItJBtaCaUa44XgExY+O4vthxpZ25E0TcER/3UfI8m3cs3kUzppPagNXkfc
wNU7WI1efovkfqS51NsEXyfOGi46E3XARA8hMc703Gv6B779wXjgCRB/RGC1uoMI
0iabQo3PjvRcjupnj/6Fj4sqqI0NcmSZDIHWw3/V+ZA25xVJ0n6zDYzfynqp926o
5zqJ0grQHU1+nUbH9A3RTyII9p/SWoWApParcwCl6Ekh/DgmYWUmI3Sgs6broM3i
bATBbWvwGdTMwYARLAUpEnlmloDJYia6XeKzQcnhnMPHec/s0l7nzgiDDULRHLDc
0g93gcBTx7VJjRjf1cfQeW4bYufz/OJhVQoE0ayyIPcCWKzV2MRDxWJCTcFhJSgk
Fg3wPQ12s7CY16uGNnDFrzK5qBKCGPc5wCdjQ5c6g0fBLbjiar3U7brGZh79+Jou
Icn3jc6ZWiPqfqmUXAOS7+5tg+1/V+I6XdjY01yIvX0+UWJTe2DHzKefLtJGuXMX
yRkX6fx+WlG56/pk3nut3Zb0FJxaG7SWTGVc1WgJgCignk+hNX4oooi7N4EERzn5
zScuQh/+21wGI8U9e1hrcoQSON+9cd6zq6fatRVw0tvXQPxZkO/ulqUird8Dk5gV
iE4UnDzoIzo5FJGvx/daf1jk+lZP0/YcQaWbgjrs0YOPDX55JINSjCBSH6CLcNOC
fLboTSxoj3N7cAhNvETr9URxLZfMZqerA2duqUT1jxlMRw3scphlN11NjrHivmhC
cUUIjzi9C6XAeW4LWAyefWNzZf8VwH3JtqUgoHz5gvAFf32TYjqy3okgmuMajfPd
hrTMyC8LB5oWt5zWYJruc2WMOjsppZua+OOpSHakjxYpVeMV9iQ5benzRmv599D6
9o+nM2kpZ9BLBhswX5gGq6NqtIZy6NASpBss1tv+NU0UdqGJHbqH1vWVbOi+9HFI
HShTPxgvnpRxmGndGERzNzGrDrJCJbfd96D9fdTXPy+a0dOPa6iDEtjXtVCIUgVA
1jFxX6MHPJpLF0Hpc70xRqlAdEPJSlVd78mO1DswzfY6C44j6EcwfaBH1nAmz4wJ
mqM75oXZDtzlr9ssryIfpWTvuRg02YC0EWmQLFx2OqwIpiOT3MIAPJAlHVN8f1JC
xcOhRTYNZJ0lYw9pGUUd9YJGKOvEqNs62ikXzXrMdiZbTFOTfdkTk5KUL2tHQj31
4ivvCryJt3Fhuj4DyWMpdXSsuV0hrblZigx9xYDjORzInQJgkVMn1TIjCBQoYVZq
rxrk6lew+tc0Ltd8RBDqfe0Ca70q1B4Ju6TzXwWJkgMpCOHWayls/PfL3hkmMNP0
0bwj5aEd/7s2Ns81ejco4HJDL0qjA9OSHHVgHgMzvFfu4SyG8qAoKTwQzRe8p+Ve
j5M5IgCxtiY3TV6XdHC1Ak77uyAbgzyiGIpgufFfFQuhhDjJhfLTNECq/FXSy1AC
rtJExo0b1vmWSjpbZkM7TeYSgb/M/zGosopaZhIt7rLvgrrdiDFsmkZsQhxFyFdx
ORWkWpXmXdXq/Bu8OW43oblLFmG9MmbzwZSGLs5+p9suRJvhE998IQacJ9W99C8F
9/lra/mFizppcW3TZo/dhpnEv1H2U2VSWF+h0ckdVE1HRrA9rhOLCD4Ttm5F7m8E
DkCJ5CuqchXB9rLYzUAPMZmHeCHykgSRqKjgvYoXIVFkpeh6nfYt3WSBnU0c1jTp
V0txhRWvOPrieoGk6+XHWkZruZM1UCFc8gN85ZW4I9zw9BDAOZdsJ01SvA/FBy44
Y9ztZOuVzBtKXhc55G6Hgib34wBhEX8XUFpR8z3Y5pxA1D65kaA7eUS5X7iLd5Ys
Bst9YdIp+nkF4OT2TditQlt4kkxaBroVefc3/fYzJ0bC/Kl3HjeFH0RSFqMZv1GX
zt9t7BuSBayAAQrOV7lc69mRH75M0W+vnDY0e/IkjMN4/31ZujJMMsm1m1HJjwO/
fgTSPxc6++7UxlNaWngIopSrPIpaTQJrOFLPJjSrjj9o/MAaVTZQLUSe6kVykYKx
M6f/WkcPPNmB/Uz1wkjcY29vGTbKQo48DahGXPpPs8KofbwDyA7UHS9vlWO8HWWH
dLOjuyXGb4peW3sCJUz5BaIide0RFeX63lIiOsnHQZ3PppyQRPuJdDVZwdSjiwTv
vpsW1p0rJi3gpjcloV8V6NmoSp21fuhI+7JsriH7RWmLdpZEpk9IQXghuZfy8N3w
nt4ttm/fa1E9ERbn4YLnw2iU+tR0FNN4qHmfXUKkhn9BpXqcjzsYGTBypCm4clU0
x59eNB4vsPd9OFNX6NP3ppDNTWHuZCSc9UFVP4fJOZMHtcB/BwkX22cGNYZDvITM
7sRW1alZs3LKyIi3mSgJ7nBe6RIc17KfZLWAk6Y8yEKOJVrbJeNDmeo7dMkqw+ru
prcDW7kcjflLxjgR0+mI+gntW185kXQEjG1hhBlxM7gomzmSQYcChb1XF+KHN2uc
IFD4AKmDCQmKtW8wBZFmmExqqSfvC7ilFV/W2sR8hASwH0AVLhUHL+5/2NjA3MnP
nh6b4I6BA0guuW7Ut2Ec44Z+py9w/g86cRnAVHeM6ZJkxPRc8REc50ORV0nz1lQi
1rHFNKE2ZZiSVE7GRYYNHbdt5IxUI1V1Y5KrnOw5tRm323AvSIj6mfEtQrSrlAAq
NH92YeEiU082C+4l/cwf8COLBqMMGpxTEVCc/Oue4tr19dbbJ/p5e2y20cU+IHK+
NRnOkPTT8y2WFPVlrnYvNaiOaw/uXxcGssAqIXtEK5ESGWHE4DoGj/we5WpcU9p+
blHPCeQgdhKzENHk+YP7xnyFN0xubwItJd7qOYn4acRUbsPBoU7fp6qbjs7QMhGa
G3smnsGOxyhgnCguk2bHGOUudVpHX3kOfybhBVkdJpTFXiIfHWH1Wr2Xi2YBRoSX
DTzp5/kk23SAApSpLr5XF1xGn/eNAgQ8QJcobT9PTaMOkjHhWCQmzsO+S4YRAxXc
8RZUbLIPJeJ/hxkq2kJMcd3QtrqSF/4kz0Aa34WEMa1VWWIFZRAQ7sE7rASeWAdD
vPlXg2L5SPKrrCtKVfFMpMNoZ7UgqI0/AJ871qPHY/dKI5ko3hKe6aqHTlLPZEfF
fpEOiikGraeVrVXWOeOaOkB9ojW7H9BS8edtIERscuIfK2xEkHJszbfIrKNZleLL
Ej1TdEfTmYulJazHawNNet0rEproA8PNpcxNEhvejeVVKWMN4jOwJrX8uJmFZx9d
lWGcwPb8DhI1akrlc/4raIoWQ9w3OZumb/m8vT3lsXPN4MWWOpcpdm5U3gUmf9z1
/XRQHni8TmtfozH8BYv/dn1N3WUuiAmqwYnv3SWp5M+nL/ModsxBbLZRLGG+83Cr
ZB6SBFpk21GD9Xnnm0IJvW5OyMncFDQiDYbj+t6seKmI3MeukpVFf+f1xMlEF1q3
9G2dFQMBVjA9LXGri/KbhknuY2Oqslj8JjRrRjUXnEv7NKo/fTokEzFhIhO6+yKB
4b38EdeGozsNj7VoT0PvAShvS4ybfLanekYBSH6elrC0Vgpb2QY6zzG05tsfHu0u
hkviqwJ9OsFyuTtXEK0Os7bdGQ0PCRYt906vzmHWckHBsgSTPFTWbut6xGILv/rb
Z3ni66FNJP85LQBJ8o3KoPxB8OQtVMvZy1CidEG7VSLjVh0/nR1TYSAMwcbR0iSq
SLLJuoCfe0iAkzFdiX6md4+HMK5qeVDFzuj19AlKkAz/4XLdu2mcT5rJHD93k6q4
dshUicPVPNJZyhEcz7bPjyABc7p4GshTIhjtGEn6rauUWXFfXBR1FKOBbD0ht6XA
fXiiz1x+pMHyDD6bWRo5XTud6TA6DJZ2ZRVRTc1Wo2m6sWwDgmqyXl5rG6QKkhzu
mBLNUlBVfLTJ8zib3vG4NuXwPRR+2Y0v82FDg1ShjzEPRKQ1AEGS6WfGXZnzoqU0
pMMdeUFOe84EOIsxafhB+Lx9BjRRl3065/18naS8yRcpbIYAvE7iVRuF+JRTBcPQ
2MNB1DB+eY96h/U5wdI/FPwqLiIqcLyxgqvP9lkd60Y6dcpJ/zGv4R6pL/BQd34m
12ocxKLLvQ/lVDDf5RuWp5/oIt4x/0vliQm2iCBgl0m1oczFxyrZJis8pH1qneah
HVB+vicfLVg7ce80Tja8YQVsEVqccg5MoAYO9AT90bToWYWM8naF5UAIZWjrSAYe
BtucQAH3EtOWMyb3Zv/5MCko4fFilg56nm+FA+F5UewqfIIYxuXQCZ0p8Ln6VcoB
kelDuT8aXh1KepYm9gsGML5zcy07ubPCczvm2rbkU4KNtAQq/hfYxtR6qGonqICk
j96QBhHs4p3jRSu/WffJjSZTg9CFgfjozUq8f7yFvEVqGQyFz0+S2uxaP9tns3MQ
G8ngQvZr9vDTl/8yoD6d+sBvRnbVm+RVa6dSnP3l8wh38pa4FbTFDdY/MvPU8cSQ
yj0Jm9fkehgHwCyGQ2/RokLvDbyQmoH2p5QO+nxanq72gyu1rbc9e4BrskS1MYSG
PJCjm1rsKqwxGk/W2lA5ytV9zZ7xqPYTWsXiBPCvRw/87nJmu+UzBiZZTbCXvVXt
Jy0/LSiBVzb5u3oDLfWyzrSMrj75MX0SCtUYtaKV3YzJ8a7bPcbGyESsusSqwkk1
uZgP7x8hpjFsoTfk3btVsc4iIwZxJstd/9jB45K5Y9XvbaOcKAhf83G2z0gq+k8y
7t7rismWDX7NsWgQDHlMhCD0/jPQExjxWI6/RAUJbXd8Gv/94SWQIff1qxBDEshv
gbmQtBwu7BkmyXZA0iUHKGg5REtQcF6qNwLQxi9Nhtgwvj7CmQjBpMZu2KjFGxmO
tcAEojJfwYJr/0ntiS39z5MjLuoEkKmSu6sidCisvPiOgXdB8DwHHeEunVsSiAvd
hHfUizEQvKK6XOkQSF1N4Vrj+xxGtqZppkfqDg5BySftO+DB4LHphJgu1fBMULJN
Tfkin9LD/BNfdt4JZ9/m7Eu22Nw35EPDWDfx+9VK08l5GXlSou2H4oqbaIRCB4uT
5rIZNQ4mneGskfFXMzahqYkqFT4VH5limJmG40atqYNwsuFgSYt/+KcErEcW6fNN
ndF3OOhUh989S95jrxszkHu6C0tWSulqmRHEm2M/vKiL+C7k/cKnFKJaCNbtgkHv
7sSSBvF/+a4WOX32Rhy7N2jOyrwBOMnqOzkunLPgiEX3AYpov3sAIiH0MhFwsT/m
DnZHw1WdCm+8GdEofUGktUa0tDwN7My6aFr2ZxM1LumElOqXOxkatBIfn9nC1sR2
/GxOsnTtslQZBet2QEutTWGyCBHJyPE7VryHwM6HAAnxJFifD+Ee4hRM92quIGTd
RViALbJfXyOyBvV3HOTpmMlw5Pk8U9LBYnocWW9LAXmpfhYnAjhGk0GfAfI/Ntl+
r4tZce9U3H4UW9ax7Wfr4iqEuC1myIX5f+krfogtH4Tn4fsfpAllbXgARnpBOtrj
X4IirgCpsERt6XmjlnUghhlzsP3OUwuvMULcgRhajssIYBK6HiwX3nDF7EyLs7e8
QXI1ojea3WoxpjueAP5a94CW08svv32AKUngGee/OjpwX5b3mVsjwei8ghf/ndrc
NYFLCON2GWmXZVRcNXir+7wgT56e3XMrHoyqw8DDboKDPi+rLkg8DwPIqw7JNQmT
GeIOUWjnHRTFDgqDZ4rHhjkRfJeXImKTLXGPUW4EI8ccnAp2Y28LKaABrguK0AT8
/cdiya6W4zepcKpn+AMghySW4lGgw/CsGu8K9/5YhC/F5a7PrKaTyfEXKqPcIEws
pSEY9sTnlr62vbTWwJe1MraD9/EqZtj3NRmP+CcbExCKMJAsW0QYvEchsEqr4us2
lueqdMMEAAJUKPDV5LcL1n+95Zf8Bz8C1aZqp22/YKmZ1pyQEGfeKPSXN+XVbIib
Cf+bdTmiHDpg4t+mKRjUDLatXGRoET5As5jqmqYoqLLqoP4L13mAFmt6SMtUrh8+
BiYkSTwK8CHPdtP5sXO3DSDk5wAWbol/VcWy+OFT6qWxzNAWuDq2Vslo1M3EJ+y2
gIP6qOJswhyGGiwyJGyiss9HO4ITbMoGWOfgW6yt6jdoIU2X58pmDYobSS7d8wBw
7L9weH43AaNCbqa+FxAfhqE3NSzk6PkD/AV5RwGrRrlGJhvu0fvQvcI4MS1XuAOY
IRgfxQ83hppzYufd0YidXVlyDsNwWsGLFiRyfCIBNJuVeDMe9qqBrfBlVFLZ+NlX
H3CeTnlJlcGe5cdhLkq6SrhKvx+qnRPi4ElfakQHCbGN6P+VDXA+hMopik+BJG5t
9STPZl3lGZ+asUMw9CcdjHp85XC9TRckKs/yvS+EuZNcmSHEOq/rPFLXoA9Ag8qL
/k1Wsrl5Zet1eUSNvSAjFNvcQtNxkq5IcDBnnUP+07OJkM7lTX8cBO7dPVzFDTdX
oNDpps0VTRbNztvXJl3QMac2KuifbeOysD45lUNzG7xkpNX2cZ/TsEWMpVHE2z6v
A3RZ0MMyCedVuHKC6AsW7mjmdglO2u30xQYyzG8k+a4hvboIHyxgms85zI/iPimh
Tl1aUUPRrlxKQNgdZes2k2cFR5txN651Sl0vmSYedoIzeu8fxKIhMoSFjcY7q2l8
2brfHmFoogUFmsPb6dxc54Gq57Bzs3kzfKFs4iG0wnuYYWplaN+XREojFkoctArj
bUvbL1uEkDtinqbi1SBZVtPDInfgPfiKt7aWc5YZPeAEjj9HtxpChirSpaeaWa3v
YxfUlwszJ5YbLlgadHPMWZ+BDlj9ZvTukW5am8ODLPBCPcsDe/0EV/+pC7iQLTdR
9LRgxsxvHuzSZFd7KGPDBcdD+RLIE4MAI0HCz21kXz+QtLTUf89r2VVakYDKrSIq
60+VEByV135yTdIvHKdZLc2XVgyWNyqIZ7kksotBLg6CqsmQj5liB+kWorYCinow
Sq/GEbZ4WpQntUigBXOM1wGg0bLRHyq+4T89TZhE8tv2GXgH6l8HMuhvIERCphiV
+9sEw3fXwqrwuR0jKxSBpltQDbxUzZ/BkE4bUdlMzU2SRxnHY7dkGTQlGae1iPol
xSjloTX2D+9bbMsSAgfDvquaBzuobCHM+H+cwrGGE6tjMQEEyjyLZ0yavHIGH6WO
8a7nshxyWDDPf5u411ZJRrDFN1K5eZVgR1RmbXhOpy5QCyp5djggDIFBIANi8fFv
hsordOC7I06XDCUxfNoITeju0xNhs8kDz2YasLXAywQYxQ9DGUNPbnn23m0/chKx
fJpzgalDwkaBQJb1wBDo6hVA8N3KOyhVpM+i6PlwvdGPUhOMrLLbLIbopBQA7iWn
HMvAH33XFSpoyIoVZyNK1EnAiRtz4xdzhDJ81/+bTcVx3XEZ2mWqTDVjOOqbJt64
QuSRfuI+QpieNjtFk9SHxOVoYb7cTlk744Jv/2JqX8hYDCXMz5LtcEM+ktvmfYAt
faMtOYDy/SRIEGigzFkdEIqEucpnn+Otfz5L33fHNM/nOT7fZ1To7JCrpHG8f2Ew
SPXttFz3oM8KbJXqm4RxaI2qWdZ9fuQhJljDeJn8umevsnmbVzfgh4ayErQkcyM0
xeJExA79Czy7m1iqMpFo9L1kRMgoEzejOnn0v7VuoqfEQ2kadfJDMOtcp5TXddWz
L08wTRAWeTNBLptTYrCipAeuD5PUzciM9lSNhSfdLBmZ04AAD9ZdlbWLd7I4WRan
LlvF2ROWfXtRzpsVHuBnkWyop5nos4j7GZ4+E80usVyeEwx60Ziw+hhBc/2Fdw/v
SsobZANB3JFDyQRETBPrDjZ09gS04/37eTyuDasIihB3+Qseqh3gXSeAQo9wU94h
gUPNkPRf0d9biCjMyclseJinsJsiRydZzDEOuC6yamNWj80nK5MaA/Q5u3nyEh6/
1+9L38cCbzXqlUmcb4paraEtY/Dhafbop9y9AWDawNcHIYyUX7ZXhLyZ7/Qnz46x
c7JJtqvkzTDNhJI+M7vEXf2BKS4oZx+Ll7FOb0Dqfm6M6PbCBFpNewFnqsfeWb/g
XfOvq+je0onKsPOBDQTDF9lMk3BP5l2xoq8MUvFYk9oK4rt7tzqf87mGCcQkYcxd
/41pDKLkckCY2//MLE5YMQhU9uI8y8qs+r/GlCvIQV9pBSn9Ki9gx+PDdL5UfxUm
sTIXU1iAVn/2+LqDsNP8OuDr6I+O7bvAGUkokzTIyBB6J+OUKr77O/PyBxNFwKnk
ueZLgEYwde9u4ApKLWsM6jRrGqC7BNpbEQ2ojz4pq2a5sQ+KoDhs4aXCq87rC59+
JZOPsu5pBVyd8yFI12echCudjUIye0sl6/CX4klVMcibL2C4QI0l6kCq86CdbmqC
lqM+Pd/UMJsHvM5Bz+EOGtuksaeceLVtbpZSoqvnE/19fEFE71K/qc9tp/QRnion
uOuoVKwGTmPXAnaN5acMSdw6Z/cU1R/57F/jqXjmQ6h4M8zAvYLs4fwfPPE/3MG/
ENknPw2UhLFJqxvlwz47YNXE26sOsjg+U+zvD5M7oNDisw2DSwS74R7CqP0HIYpW
iUcq/KFkl2C9FYKtCRf2un3BFM+4VTZf9Od5LRNDIKDEm8meIf2n596fIy6p4kxf
jDcclEZah8empQBNJ87E9ANFznLqgiGqiSEKCvg4tm+StijkepnuIWjLLcj7Kojz
f3zV2IPrtgPK8vEwfxxqKTdZ1FgQsz5lKaqDXlKMtY9sCr7hfEoBMgsvngeHR0rQ
+RWxDgwudzU9TWvXMr3N3R/9kO3Z42+pQvKPsdyVbHQ5TooP777ZE6dlaEPW7yUU
qxeIC7Gi9Qk/Vx3sZ4RCLtIWmcu2vppp4L74neu0Mb2CVc8HS0hgbn2tj6LoYQud
fH4M0VbWQ1qOd2v9rcvYSY/oSLWI6tMFqu0y39F4kT9YjN+j7DgZNuvXm2H1zZBh
TMno++qtGio/vvoO5nFldQcSAR4bo8kFGwylCWioNLJAhhKRI49y12XNTK75qtjs
VnmyjtQRXrbiRYI6MjnZbLmCYAXh09h13ND2eUb0+ePzgzMsreR8yJI4QyPOMbEP
mvpJEvsh986ZTG4eUipedWp0XpBQ1rEkEY0IToyeW/jKtMYuTTtwPnHS5Kwvl54D
nACtT8wX2QVmPFKW2h9CPB+vKNqFu6qGCaj3BpBAHxAaCsdvLZPCfS6MisZbooFl
UCGyJIhcs/OJZAv2BkjyziLtXNUxwCN7MqmShZms16vANv7K+qOABfhisZEOgRm1
jHk5t1L99byMPaTL2iQ1+IlYjZ8IVziKo/OJ2stPGoVcfYaVVwNqfkseTmGG4Va8
iV9JU6RY5u8McTY/KKWk5m0Q6zCq2K2c04QJV/TPrTIMuEJIuAVAj4nY/Jxcr/ZI
v/1fVhaKfe77/Ewt9ID+87lGsP3KSS3g8H0+ZLTfAKUdT/zeO2GCSUedOtnxD7Ap
uSv0xa5aH0m7QjJRYu3HojudUO0xBWjkRM3lUG8qKVsWSj6K6r6EukWNPYwqzeiv
enK39yJLVq79eTK7TdUBxGL1+SGLecipmunvV/Y7l/hdMpcv/xhmslnAeHx9eyLW
NfwsTJcs1Y+yPW2ePY0KuuTbUuQnFZHiL1DvA+Yi6m58sOsIhsTyP8vNRjw1wwuF
/pW2pyuGQharP3shTUpiCKrjiVS/6tPP8goGbWNCQUlESCsKp/2RVIUzerkPyX/H
M640TFiY3vOOcIcnfqEDzf/2YOnFjK+1gJDSLec38+1eZjM3Yxc43rjhaUZ3D/vG
G6hieIKuwkF/Bu6wxzZKBA3SxNjm5TXzS5HhlGbB2+FbHP+r2NPzGg1d9N0PO8Un
OjFOTU+O+NLjzVnbRiexSS0J30M1i4BS1g5w9RClXmo/qPR7U0fnwx4T+aV8BUBy
RmxI3FA4r3sQaJxdHV5pGUFASoSkqU224Orrw+wM9WF5Qpo6IytD7j0YO/sVhNOF
KsOH+CITz31K01euI0OuRRACadrIfOpUiG55yDPFReuo/o9rOeeOF1krcPBdkKB3
K4yo2mQ1txxLwYJzOHd05TycS4LVONGfsvPoyK1uqphALOQx4NcsdgPaJ37lqr3h
Mp2XozCyFH/DVCCHEy1/78DsBEBRA6ESo5KIxe+9aAydIyIPYUcfrIf/LOM9jYjX
dG8KO4bfTOpRf4JvGsTfvKArlbkZePtcL1+MCF5FH1+g3yu+yzZKq5g8jC2q0J83
aj6krQGZIWrMO56eD+AtBGzH58LMkGgTGsKRZ5B+bH26dgklV0Oyp4l7rxcdg3P6
DWJ3M3/dyhc1fZ0VzzRHNGStu/u0gzsmzK57DC+Iiva657HvbsDX2DnwumdkC+ut
vwqfdQFn1spt0ikJhX4/sWAEjy9Z+qs/UxlA5EPBS+6aKVudD2Co2RbRpdyVrVLV
hW8UAEpTKk0coJUEc4v0SLiKjhL/60LKSk7NISxzal7jYMkaviN7xWhO3f9aAKo7
6or+aFNVb1LmyT5WsZMUBPMCWPU5DaHORNqLS3JcPXdASbo6rz+EuAv174jeExXX
WU3TsN5YUNrn5q1Tunjr7gk/APrSurO3AwEstARaT5Aqf9TxyW8S4T7F0ZRik+o8
uOa0tjlH6pABGuILvX3ScWL0PDKvEy0lCZqiB6MP16h55Mm8+SeBtmqbg1rtv0yv
Nb/RQFdXLa7t6X4IasnK5em9cTHRSH7ay84lvLfC6ZuTRsKg7gWiQwAL8NvTKyqV
VDfRuS1DyGAMVoIhUtp3RkN6TpqPFrdeX36+wvTyd2bEYEQV/hIxweUwKIwP9HT9
HiSZI15X1C5tvp3/Wi5tZqMeNKBKe/TBdXyLKtMwTq+/zfRH4aotHyoh/K+nkDIb
nqgJTep9iDHaJJty3OZqghKJxnxP5kj/awEbGcQXa1sUMS892mnyrM4qc7g4T+5C
cw2sB/rtU/Ck+VblacLgl1a+YsiChqfCpDcESAIP67LPqMa7ieL0pCjfIy1AfcTD
/Qc+HJ4WccuJrFRmHVAGts5IXVOlkbruPaD6CCSS6QpelIo+TOOAnrqaUr2xWGpU
4v3cM/Q/2kzWxeq0aM24dC0oz0A0EWV5OvYvQiB9F8ZmSQgAFoAjPrw4CSdP3ido
GIv7kxjkJ9YRblr2ZBN+iv9ZaA8ObU4y8WTMAB+7IRqUxE1VvcbXgtaOu5GcSkgb
VgP9E5fKKHbtTJOJ23Zubye/hk30grxeRVdG8o1hO5nKi/IODm8jWMWLgCDH7P5M
cU3M2ZVeBDOlvrzlDqAd5Qe9sgjtwM64MehL40pD4ZLZ3PnkDBNGLfUrQZAa8gok
70VsPHHQjW5fs0oHVOBbTlUZEOmv2Nfk/xMecFiK2wbIYI6DvsG71ov0WLvf67af
a3S7L/ShvqvecIx4sQxQ/wRMOFbam00VCvy5kyHd1eJul3/3PgTHaTGnj7mFSDa3
r59Vd3e3NkcWy+loo81nhQ3mVrrahYGTbN5hzm0UIb1dSff4qpaQqXnZseWBkaHf
b/bweAH8iQKA+iVhZkUEAMj9cmub9KXiMYzrccRKvOVcx8zqJKO6/EXG2402Umfe
y19vkIBrMtkzjPT6E/KEQfyL1l7xKlJ8zDu12dwa1720s0uGdXRGxezceqPBghLE
Gm3MY8F5s6ZLS9r+uk3fAGcjxmAhtagS30EhA5exd4usiyYxgOlSBnT7Ya0J5JND
zkMewx7Fbrobm2+WPtKdqkWkAlMGtVEINH0rFV0m9fvllwjQ66meDhjEHu6K2fih
AoIpLLGPgewUXfA7jEYzM9bCkqK53QW1Bhi4ur10vOrO9es3p8ZSFR2cqcup3Cqu
xrMIxZNymTCm8VovlkOIT1Y/qItSKVXyG92iXextUBBMzZLpiP4mjSuwq0bg2+mU
My0rZku4lGlPx3Rr23skgTthQrpTlbajovn9smVe7wlVMMgDCKd4Z1WAzzgFywXV
mSC538QzOJLGaRwzSZLpKEkuG/24L68NCkPXs7yevGBplhTH2aW3osn9LUnPVHvl
I1llFzKeIJOKpUruL/N859OWhJHvVr6wnVjWrdZtj+ME+ByWpiWa/Vb9y7OQlSpS
WngDN6vLPm4QgUN/IZeSnEdYNtOK6ime1CwXD73yO4DLHG3i609pZ7dj5Z8K0Wc8
poiMgKp03xb+LrH0zaEcCOeSJ9dTHUwV0IHO8S0l2UgGhZkg6qkAqKBZWejoq4Pa
REnm6VRBkvFb64jeL3qhItomOy1H4rydZy670QAwkTMjwJoMcXnjMjodv0nwvr7N
5RNenT9Ybk+vqIeZ8NrT1UWsLSC1K5YuM6QQDfXp/jS3lUxwsZzkCtKG2SdEX2fV
Dwmlz5Jdij/ePZEGckoqfAnibb3cYq3XbCgjKo2g5OCT6GnuXOcqCAorEQpo/71w
cEggPfqvFjNfRxYF97LljRa8r38s45gItB7wh7VDYD91uSKtSb1fhTmKCIRjk4cL
L7wa4NDHGw8HQWX7k82/nZ88JIeJN8ozTBG8r90G7ABCJGGNjYj8lzUhJD53MBeF
WczTcnbkZOS8mg9sRFir018Tc+VwfQkDHcWtRY8C+beHknbFjfGakePP9vO3bg+B
k7pogmSa9IAQKJ5wB/R1h4zg+KVapCGRWxg/p6QyR30Hgc9GDzZFD5z0hWD3Ns1Z
lCIzihK1n54Qyc2EcV4M5KsVKkWJNoxEDj4oE1JaH3r/GZ4X49Xfy56P5NCLjTX1
IM1TGbQ9qqOgfHfUd2N1Q0IJaXn2BwcFFOo1eKZJCCxyq3bmxh4pca4cfOYDhqqs
W3+zDxjDRUnDdjex3nH3FtL+wGZpmldWegv4JOYSXgfDHryQp6KIa3412ae2yjfK
hly8ESjslHCEOF0Ni8h/3f0wLKVFyCTm4zCMz0+DWrJ9uHo+8UIPMyAdTLUNjpJf
uswMlQvMAXengi9eWF2FoGKqvd+PLjMs/qCGm+BeyXdeRxY9a3fWUCN4U71hkL4i
DwDw4LBLmoWa0vr0F/5NvtPgZ+7xlJEFBu1S8qG9rNQ/Y4gFL+AGMrTu72cB4BL+
Mc7fXmNruIiy3iAFRc+lsm4JWGaWFpcBUI6869sDSn8SXTYHqv6MeepJ+oiGHmEv
9RVsxyr/cQxC+ii8sGYXzFoniQO7iou80ydo+lbxagP2biQNdf4G+nyWZU7Nta9S
zfCLT2no8CL3/D3MSMtAAO0/J+lUWU/QOGRN53SnKGgmF9hJnaaWJKIeoRzSM1ea
74NekaVU9XkAjamV/jCegCWGKQNswk5S0dTmyT1u2zKU6I6tcEDhm+f0SOqRAnZI
T6kAElPbsZgze8qM8bW6CXhAcyS2swAKMAhaJgLJoevEUcddM6pAOYsX20Ha0euW
/yMdCw9csA7Og3eC3C+vDTBdA+n9uVY4YW3ERuAOIJw44U9jvUe3Iof82WcY8uZM
FtDyzBI4IwudLAVorqMFcBJhAcAdDGkAQO2ZjUgSF+3vPheM6jKJzmnuGThgvqFz
B3OOoqRVSMsDC/gMeUmHPJBDglyUa4qcNbh8ijHqL9nrhxQB7kB0zVGxZAXG5yWH
eJqGaX/4MfYzOkKWMOJA1+5kHbQDosxJSCc/ihbJQgyFim5mMCqMhyeBKxt9lJWq
mltOis8jzWJL9WAjobEL2rCHzM/E/YpwH0J89W+h3mE90xB7ZBLHJW/jstVfdqss
D3VkxoXGt7B1t/MzK0hlt/33T/KtezPE14BK7XlGLSY1PQfvkrW3Yn6VBXr+wK8v
5rCLfU+elXYEvGMgYNwqImb+WOOXxIdWkB4eRHfFn2zru+2aRLhIq7Zp18QG5L3c
LT91oE1LlwcYuvrtqFVK3+GF7+IzZiA6Jrd9J5gQKi8V2Kaf93fXjEVAYpDKt3gx
gSlO+Mr1gOFHP5gHWPQZtAgxnCDHJjNaf8Ku/mj5L9J2yLf4LEeG2pgvYjaWB7xi
QtySKUKmc10rSTcd0KRmVpHj46EZBSiogtMsJaeXE9f8auObTFS05oJdBwRHPFO9
PRYvX087SbibzZ136toRtbegB9nYVe6EjLkQ2WRRr9l5pC3uVrH4SYQIANEqvbJT
AN1iKEi/3pb/gsL8zmUdOOOEXTW2IjwNbVH6qswT83uA7LDSv4raBuY3i91r/n8+
dopBRQGBCgVu4LblvChRXMRNCiISqmTaTv3fLXheyF57RpDTFsNdjQLImhEc42og
gNhabrQuQ/z4puv4NfbI1LHwXKFVRIwvJsXxFQDKGEdktWhh8I/+tI3aKVWgyLPT
kt/zuUHGdr4FbgWDuGYqbzwLdtMjmNnmcPeajN3scjDuhrf1EAXItXr3vRnOUBUi
u2G00h5TFuBQ57sxEe4rrITsFtP4NTkqxTDFXGf+RHGtti6Fw04U1oXz5v2tC39R
YU9qjZYESfjIU+jHqVhQG5XxVi2Dqx/0x+L0ySv42g2NPjlgYAnzK5L0rjSEgbTv
OAJU/BGVt08a0IShuYCiGNewcDg3QvoclI/rLs+eElYhAiyif1dUe2bZzHiaONWP
kPSJJIuKuFLrHoNG23neaRDaOgApFnqZXkwsevRTOZHiXPeP/YN9RN64aoJdp2qC
Cled2yN07mw0gywQq0dKyX77kNyyStdWs0GollhjVWQSH+G2psvWJKkubiDOr7OC
ahjISyd/uwWfdOB8IWyC4jCiOBchTAOYOuZqWad09jJI2lRN8hAW25dTfhVANhGb
mWG7ftdd5fBQ7S6is2BDIDf26a7j3MH9P9jY7+5xc7ynxoKp1ZF7fcmTkoZKegro
DmoX6+YG8qH84Fdo0zrWhALzt7ZroeGxSmD1mxQ1M5icXsJDKuNV0A6uSe6QaMCa
sp8c+odvvl7UjAIKW9biBqh+/4Uy3XG04/IJ4j82s54jL66KrMkbdQCHz4NmGSHb
mAYx3R2wn14hnfjjJKr3BOmb+y+wX8HBUM2Ljh+ZWzYxYq4RXDivY+VyTzVeB4q6
79sLGzMRCOoNM3v7/GJQ2jKQr7JTvpG5zKAjuiXZXsAESA3n5ZzoewAxlJ1kExxg
5AGK8misAm6ZSQ8oK0MukJrjefIcWoKymoLlHMdgV50P7+NeoacvHQikuJfBw4jC
2QHgsNCkrdE2Xh2ZI2V7jISDMvcVgU1hTqTomaCI6aFXWyjLgdRIl97s0CkAJM9r
lgOO9Z1Eo/QRuEz6sTfbouZ6pklvdSg82fff2fduyLCk3JaVukhUxOKr+V9ffO9z
WEyf4cTjKqrRiI29CIe2tCKDF/1g31Mv6S06R5df3EgsT3hUJAOTMJ4V/aJEEnHt
/nEiwofyNB0PPs8wUaBcr/0iwtuG7SEOTKoOTdVewWbw9A4jTeZ3G75Rto/KAWf/
BKoIu9lDvQHnPAxnj13CEoLWvjqUZTs9DR6k/8tvd5H4jvcIres9r2kddV0mukZl
i+wi/bHH/B4Wm0mBrmSWr7aE4D9AQ469eh7VjO0CBYSC1DSeFGVtGFIKqBc8rYPS
NitLMZ8+0y9GdrBkJfm0ahu9rVTHcpa7LKqVSQaP2bQjI8rmS1qacbuBOHduK5Cp
V56T71coL/KGlX0dZFPrb/O3PGo9qssormzQ6lyWochKrtV9SQeUKLpeJlONi3GB
/nIEkVzva2H9w/8e5c74iOS9RhfhP8aIo+R8TAeHJKhVvBcEPf/mQ67xGOgdFoai
62mji2eLTFPQcqs9ZhcuArJrGqlq3cLXZdkOC7LgCIrpepER0CnHJIItDNuoBLZ8
2bj4NBMR1ezpSn3dEfGgKulk47bUfjxOJ50DUpP32j+51gafqER4zyAv24cHfF5m
9ss5G+vEbbM3piReDo5KTrLdhpZN116Kbo9kr2us8roBRjbfUzOT1rQMgp6sZDme
2seqX7sp8QZj/k4RNM6rpFu6RB+ZWEoVN/t4JrWwYMAq6lgqkFXwBgikQUPcSn0o
6V+MGlE15nuOWYzyjAEV4/66toh/LJoxXzERh4oOkuf+yU6o/nybJAxBkHkctwKG
LuBOr2JhahQuz6MFZbonTlQXFhAK31wiQXXmi3ppqy6YyVr8+1dli7RnmPsp01xl
C+c1fmiqrxsbvW7++nt3FsXnkzPtkwum4BKSSaYJND/SHJZFAw6USDsnDlLWsGeu
BHo7h4wVAbOYwskif5K04Ig6YECthbFvlTsLSSgibRf7cAIV2BHfLOZkPkpjiNoK
dbM2tkMIgvemS6qpShu6xkXGxNiZKcL7sVwIBzyFof5vWGLLLPd8sDelzcRsr5LH
O6wNxQOgebjHVR5nOW2sdFLfnThrt0k8tllldIY8I1IHme1fvb1MohzVJKFR0dsf
W3x0xPaThQlinr+B2bWzXP18y6xYljz9T8HicKmWFoKU1wnb/CgxlZhqsGniUebY
2Qri/gwlznZ8cgEYDg+uM7feRQBGyh3pNyokSj68zOz9mpoO52vRtbiDbSGX+LQh
KAswWApnfFIbYl3hJ6bM+EIgFy5m+B1XalrqfezKs2Z6xtb9RKRkcJxJS6qWgG0a
xd4B5AkEHiZsuRZ4m68Ljkhl71b6foJSuqaZGbweG00GHml/wpzsnzDbHxMvY3Ze
so+zCnSZmm1grgLUsXO6JXAp0L2bSRFe0XN7VMiQMNglYN3USLgrZFeMpm14ajfl
Mbl+7t/7JukWDtVRnR9pJySUko5DQrQFI2xT/fuaVzRQzymXkru0zvMVfpLclLoR
gjBzIQDUwLRYisA68+6uYM89Rdutt9+lKN68u+vrKMAoVKT5rzRHMYva4S27eXya
rs3brwZIowxYiW1Sp0IYy6mn1IxXQXBHhE8fh/+iMlMQ9aMEX8ApeNO61HzIcjGk
BD0yqy5knhhY01zK1z/m67aAY7uooIK4tNzl+UzfAktw6HktnFcXuQvw0WFVImTl
EZ9ax7EiFSkykpV5er8EyH6Q/PAr8HmlsjYJe7BaDAltxhR8fb+zcDvi32hLgnlC
soYaKYDHm1daOQX3DPC164ncmjH4d7zeyN5leg5HXM9Up0+DEOZKWaVsWcaSWOU1
J22wPRX71iMkDn8wTGQ9Z6pDTUbkE7pw2f4W1np6pp8RYkOZLD71oPnMrlq3P7Eg
bKBUIAdjznIFt06drCbBw19FmBx0ZWDlaAEyGnQ0KaG5cOw5dR7HbRXZfag1ICsS
vEVNNYscA40WGQ0/uiAE8hcjc/nycUs2lV2bLDGr3mBcEvqsZgFmWX5M2RrxFmXd
Ud+vOJMCNJ3v7TVZhtY1/hDfTtfmOoehS0CzRwCwxyH3W4KuZtzx6+vid6UyDWb/
4G8e25osakMQlqIy9zjunZSVOr0Toj8bv60fX4X4Y2OHNIUlRqRyFO4MTFn6s7DF
gYFjrIC/oS/qyBNpby54wlmc+i1IZmW4ylTrpjiA2yNMASuj7GCid5/Cps1OMWyj
3vSVQGA71ds5Ep3+KViAZ2BLZyHZDfsRChLsw03XupAboXyPs2VNTILZYbYasSd4
Qa6UWzqaVSBI0AyBPLn6JWNvOM7D6FsD3fVPR0HiWK8QLZdMv2GZQaVTKejmGAmh
7jwkt7YQcD/Z6NpKnK5T3wgdInNtgTsQWKPi9Y4e+E0f5nXXyLs9al2uLkxO5g9X
U396+fertVoqGEQjo/5J2Zjnm4ocuMEDbl+QA+3FjcKvK03pbnPYh4InckIgwoKW
olhQTW1iTDgdIg1s6gjAG1hfJFws0HSs9Q21iIbqBVfjVd9ff1LiVvugv+CG52zd
j9xhtc99S+48xbfT8u2TqYhg83LOZ5P8IdCfjqtNeaYrd9Y0aWDIpAGXBxec0MOm
obSINyu/Y8q/ZaRpjn2OSSHb1njt3cVgC+3fGmr+3CW3opbu1iCgQJSy1UCfMihu
Jnm9L3KYpy4gVcK7IaRcVl2WJFtJjAdtvpO39z05kQx/T7FbgSK3ok7jZqnv44iM
QjquKJwA8W4OphR/okWRv18tPisQezNy1qbhmcN9RDzn4bvORVjImwhXxIZDtluo
y/Ntv0Zey+2/ZPkOGcBMUwP1EH32Jbcl31INuu+U51OPVHRtucnB6TbiGMIf9ZGU
Lrz1a36osKAL3xfnNL4D3CprpIgA3QDed68fzh4VyEGxqX+wiTbRksu2+58HQbdX
OMm+x8djn0w2EdNWIkkL5TLv43/EKTQFy4JqGNEmHyOLJCUDmfHFA2gGVnXoDWt+
NjkS+5/GqE8pEvf1RXGgw9i2M4CJ4SbgcaM9ax/nadpavwPHAjgO1l5X2XGJ5b77
4CVztZq+zfrwYEPu6QEWdp3CfR7FDiAZ08gKKATKM2oRzJqYNf2ZyV95DeIC0Kfz
woSTkxBiEkbjGVUUriP0l8nmF/YIYooFrMBjiCT+SxiZTVxLmuHULFHkgaNk3hb9
4zYO4RuTx0mgdNxxZgbS7IdFmnZcNh8udJ0+5iO6kv1ysTowWZIf/b/+uHjU/UZK
Ybks7XvGz5tqbjE4fae0FLNoMPFW6gOPleY9g9b0ynPVr7R3g1UaND807+S2c+WX
CAGaKPpKIJBMsOjHNeDPQZl+cR26bZ3A0cwQA3CPXGkmCwwg8htWbYyr1/HbB5/m
khopgEzJKsIYzidJg2TnBerRc0ngbcXdiyhBfLNvt0mXvUTf/rGUj1Su2Ny8ubok
d/+mgtZDB5AXaMNf8ZjXiOuvHCsbkGxVBIkC6jDVjrur26c+iupfIKM7HUzwYy/t
OpLLBUoY2fzPuMr3AVzp+F26cuTfnbWC/ejCEn8slxjbiYPUcdDlqCarC8ZId2z3
3qP+VVsDDSEfzXUnj1q/C999iUN4ic+hHAF4o8NKfXKtCv/fUfON3O6GVgVw4+AC
Akl5IGDi9ia80lEJVUqJkd8O6qBte4Q5Q+ANbi1qlFZFfpuA7utM93P+Z2JduNsh
AOIuhhvPG2c83meotRrm5umkPOY9peUsgY2EQBVZzhML+6urk7uujSZC1uD+bHL/
GRNCgNpdCWIq3sNK1X8iWc+Tbk4WsjwnyopUqwjdrxL6I3CoNJ/5H2WlDBo7MV8y
jjYIa6nw/tbz/g05I3QU6nDxBKBKaGLvmeLfHQ/C9+ZH5BYdiPtEoPVkAxI6vHHI
kJTOZ3znbuHx0zkvVno79cJUiZGgDoUrCgS6cY4mnomPCBGbSZPd/jzfqt4NCSby
bPzl2cigU0Cl98uf+Pb31hLUKOd2JDL1oMp9GdErMXSdN31gkF7ObiKNKKZr3+Rg
J7S6lqUC1D/IYs+rofvAxe4G0tipOrx0OK+3ysDSCyY6Hl9X0JK2VFnPND5VvaG/
292zT2u/xfz2n7oCpkuqsAT/ohbv9JRc3vF2yq57Zc2xcdi6/VH+A5PMYOfkAjNS
5Sp2uZEOa4Nt8aJqahSd5pq9oyaKHPo0Gf5lofawaQle1ZSeZOj4XVcY0z5VHc4N
0uK2ApTX8fpGY3LspNApUlyjNRzM+lqwq5P50HwMDOmp0k+Nf6a6Zgxi5MRIAJrs
8d0zxg136gdyvWpHrYKROjg/fRT9U2/JKYSmD3i0WgebHNC8PMbZrBu6pnxY2tZq
eNS7vu5Dm9PgjHRor8z/MIPFFmvHi7RQUksjQTt/yazzFKKvFQ6rnf3Ql65Q7gCj
UQpSuWTnZe7FT4S/eKyxGH2wouo7Xm29VzgqnZGt7tnTBgVf+QFdFplME1lBBKXa
bcH8YsOTui/9I86qiE0lPL4fijdSZZi7kTdxasXVRIadUiPfCWkOvFD5sZXZX9XZ
GwaWCu1GvhAV6Hmn2vW9mH0q3ZInye6Y6k4PG9Y378CY3Ve6GCadnc1V5vyDKhZ8
OQxyjihqNTQnwOXuEoCtPePeBHEDBb3H5N0C3o4in1JAFr4qS9BbYVEr0Et/bx8X
oj7yaha+eNsUGMzCaTyeRUlxxRuWizArH+Wj+FclgFZmBlk9e2QyNDy3IzqLJ4A6
6/fGK9Tu327d8xBccoYetNWhgLEcuazyDlGAIe/y4xOyrsOzgf0stlOUuccnhpeJ
EIDBC31VBQ5eT/TJavR4ij+VT1FDVq26nTh9qiGmHl0kFLG1cwgdmZyy+aVJypZi
8VFJhlHaBjGhG2K+ODXg1VpwtAyCXKeiLKrgKB8n10Whgdzlq+FgA+qIdNm/Z2Ow
4V5Kf1FGS3F2w3Y7mYlnQOj+XaqTTkyAjMXzMwsMZ9m7m46l7+0mtq7O5XpNU1Jk
58swGaPz5BpSdV4N4s39g8qjLYA+/gSAoUSTqchm/K3s32WfI3DCS2O19THSq+8h
rG3Fd0/xPHu2l67VYNGkSkZcROheObllhd/i97fWLL8Av2hihsYBMjogHOamRYSo
TO4HMG3ichMyqTRs0CLotfIeDqLwnXzoTuc1iEPzg4K7vYiqdAH9rVVyC7uO5zpF
yxx61Tu5N8dPVb6hjff3mMj5apdg3nJ6htkCe/lJZheW0k9Srf4Jopj/mluzKdp6
R0k4vOEAEXntWJwOcvrOjF679WuE/E7JcDAG4qSa2bUCIIWJxQ8z0z5qcJ3qX3aN
9hFKlA3d0PuoeUqqOzbh6zUiCN9LWfu2DNNIsFmWX8qN7QEmhMrQQPCoEfhkj6j4
5eYroDd3c2ogulMx9gTfJboz4YEgS+RP8vVWo/sjZC5ZZJ6MlkEA+8qL7ljWPeox
g4N8gXTjlJRygyy12hMGldhocsORTJXUFGYZJcaW+zcqt/S2/8opfOsp43RUn6If
RN3cLQune/lBvC8EOE86hVN9O0pTdQ4vd7p4ZeVnZ7LPtYE0teH47g6dQSJHNRl1
yZXgw9s5pt47YY3SZihzgqNJ6Ko9e1asTndy9GgfZLvtQMb1vdgMHRjFIcugDpzN
jNbue6GD3yu4cGblLgdGMKlfnjlV3fXJ/Z+AZG6WRoES3d3ETjLGd61pxW8Xmp8D
bbnLYvf6244ZJrbHUZkDlPL3c4+6WruhgXPF9+mu776kdaQ/tK9EntKA5HX6Vwbk
ybWGdJnARPOq9+8JGUcURuAZwJa4DGnbmsdu1IcfnBieShvxnSqvNFQOpVVNKEzJ
chNP+PUVdLFEtBkxcr1mjG8Xheso4nD+iX5tAecwWh29vEekMe/qhH9RQ21sPcU1
LZRI9Us3MdDj90BVFR9j6LiT5SABHf2gEQchazqmF0KqD6uPck5iZUqq2My08urz
RR0RXDF3tl6rwDOT5JSvzMY6jeLbjX0on8tBj9+FTftRBsVPHwFV/s1MGlKd8tsj
IhOPo1PoaWnrxBII91P+uY28AFo5NeQRwHXixsakzHQ5U3+MXs80wypdSCHFa58R
IhOUfwNymKutZZEIq2hMBJNO+Den5x1xSDTbVBG2guZKpabn7Zwdfyloxdx9MdwC
FV22jwhDqN42v48r6W9TQrXsmOixdQBDcltSraUzBjTy/wsatpl8VJAjux91QQsp
QSCacnLZUic3S2m73+UTRv2qezD4MtGun/LccCMHVWbGb3WRpSfVyi6BGyQaYX/v
5krYQKHAjydP33Rvuaa57prrpVJ/PaEhAiiXMjKUYCpAVi9FI2UMbD/23sccos8o
Bf9m4VDubU1Rr9By4sUyQpbQeIrt0G9zn8TMqaUrfOZUB+Q618UzAg3b7VOD6ZTx
vhOeh5ewxvx1kvBCG2aVX15gocF/IvZDV7LnzAJZKGKc0fMKqPW5TpLuS2qkkuVq
YrPFZQHvONq0CuZ+iNUaGiQ97wXh5h6YvqZdwtkCNCKlGI5WBlgQn2th2Bph/bJx
duaLG4KnMM2X1Fzxav3PSkMo6wdpNtdiAs+e5YH2D/SUllNQZFLYVgtPR0Hpt8Sx
7pmE4kEqpWKXpbHiXs1gA/tA1OiJB7bomx464FGVBqktNNP04ff910sLB/boD9eP
tryI+WRykxf1X9kY4kOvOE+AJeZMcHDM7UWpRAP4D270B9VeZBAU5mZSDlYGHTFd
W6xcaXYzW1AUyCMNh3OY9VlZh/22OWZ2LndSbRDkugsc5bUgko2qPyOvW7FqqeO6
3RUuUKpHHAOGc+qi7WeiMBqfVbkP4YseR87cAEZTdETie1xPp1ZBnDb7tb+c38HN
iYZDQZU0Bx2w54R4HYtNlTUaquMFddHIXEBmxczm07BeTmjvsp7JTRA1p3uE1JNI
8ps/ZoNRQzRoDapF6wBS1xMNBfQpeRXdEJnEfsoIyQFGfMpmVyfRTURZp/BUg2KF
oaUGrXh8ZqijEgfKBTogF1RmkfqXIWuTVJE8pOenqcnLBe5rLMViaR/hqoODdHwD
LG/vPCixG0KtRUInTOk9flzbkENK6C/16W+5b1qfjzgiTl7MhzNPzJIMEkqUOJiX
uLGDk0gHAsaBp+a1yGpXowRSGAC/9/46c8NEkiWItebGBupgA18OCMcdQj6pyQmZ
7wVSMfjPrL5FbmhYE3bzdI2xfQ6cy6DWWEQ7Xo/qyDp5aKrzq9Kkgrh9OiiV5CNo
1OqCx1NdphWQ6yCDvFHzTNTOyVmCzSWjxMUU8w9XNiYvbR4eofOVDDIRud3ioQIB
/Wydw63myI3mDSGLR+xGITuVIw5r21Dy1zSmedXxyePInb7FuWLUuN9Eii74z2MZ
XrDNxdT4YnU8qGhhOpKgmkPkorhgPJoeynW/3gx92fgJ8DrbdwE4Wkb3qs2d0JlD
rtNRD9E5iGnoeBVZ3U0IvBYsQI0mXDUErURmShWk7qwMGgJ/vw2rVprHjY+IruRb
qlpscqiRvt/pDUrI0jDZUD7d0MvRWPo29Vf596F6B62dcefHuUGukff12TBQ9MGu
BzkNiIJyVZ/88htY8QeFbLO6ymUEHSZgUioV3LbxL4hNfu0CPE0TBYYppPibvsng
Tu7psSVrQIrE6+X3Vw7A/2Nh2Xt041X90XIjClP3SYfkNLwx9jcNNclxEAeulY2Z
tjFG+Hy5csaeUc9x5H19bjE7Cb+DFm5Pii1QOIbqO7abyXW1Q8IUUpLSMFopjoDR
6H829n+NpOvEVz35ihEfFdd9pqNVKhgHgyijWUbDYgC5AOrdFhMFuFu4sPwprNPQ
1GbbzW9CUav8OqvDiGqvfHFEXUE/24BjDwBQMC8k8mcDj4O9nc9/4xYtTkDTIT0m
MZVpmeessV0N3b29scfY2LumSAkmOXVY/GNQ/u21mJrXRF8tpEumEUy+O0WKCDZI
3DHnEI/2e8NxAM1bQETKMaZUSGiulamNu1ZNW7rSaF6eSF+yp+cQPjU2LGE/NVFu
Ql96W0+KQsJQXgCBGw/qXfaw/TBto1Yyu7GJX7vj5HcOwbDq66vD8QrXl1G3qsiK
YplMTnRIg2Z8AJfPnOSDKbr40TGxQxlO0ybSQOgErWIoSCi3DSrwmoUFHigz0Lbe
WPh/zK1xbZFY7Vcbu0KE/1T4iEPpe/iACCG7woz8SiuWb2kllv+DmoILISi/qhxZ
oG1x9okfNmj2/3tU5BHqqWELca3UW15srlurF9C6fjVu+A6Qd6aVs7QvjcfoaxVc
iD32pukRpSakDxF/CnMYrdsYu6u2KRlzMYoycZkMjyDIQUe8cfAqowCsztom+AFs
Z/l/OjNQONUZ7n1RYMRL4yqyESNj2RhVl1rbAX01kfILJ8V/mRI2yi5O/0QAIk1A
/i5JOCPDk9n7iQ86sFMZyUSiDVWspr4MG/Tm3dfy1dC15e1i/9++rze9CGejEREE
MMRZ2GmRIZy8utLIP5kw/sYxu6bGKPSodFp3mjLOfeLUYELEYj9P1tywqGBPazkj
LPNXff9Na1Rs4J+iMZTWcqdanZgxtXLtfsSkJ4hXf12EEyKbQqvLt3eGYE40KEPX
y8e6DmBbBEfTwka/5B59yjjUsPU/GmJde56p8wzogikkYtdTB1ctI61Lzb4462jV
U/YjzOpFb4F88dm4cV3dZYhTW+dSiuumMiuDJ4i+w2vVBN1J4dvL6j5OYAyc9HRx
LtCgy8dkZCZW0Z+l1Kj+ywHS1EyffzgT8jdkPVN9vpT9DdP4EDrtzIiIHG/U4TB/
Df3UjbGYjsWldhk4v+svIglImLHeSGaNYar3z/s3sH5VHkmRW+Bu2jAds5XrLvdm
CDyLnqGmcUoFXrrw5K7iX/8tMhbkbfe+jxAVudh/KW7IVuqOl/XCqovQJT2sQ8EE
hVZFZL/OT/u6NHzuS+zk4A6FVw+sz2Mgdghz0CoWSEcD9qUSX1+SOObd0dXsZG8K
hGnZW6yfWIBAxggHEnoYOzMZL1NfpsXEZHXz1vTAs0K7ovxjw50UBsTM5rWG3HWO
JixODiiuHo6TCwqyYanNeUTOTTyLc7JllPRXJ32Sg6ItCfxlUj3XLff5ZutYQBcr
ZjgA856oMZvWKSqmBz32Y/Sr5QSouU3r8jelbxc8IxIyPGosOQYSHIdr3G2XD0ZJ
Av1msJOK7+pSpXYDwcgOAZwKr5nMZV/Sftqagd6t7x0t9IbBznIGl+zxMRRcsEup
CVVi1V0J9Ovm05E7nRKsdVnVF6Gl0ZiF64YYGtS6xLugPk9qIocD3ghYdyX1ifd9
7NwVVWTeAbKHvQlz2gdP6Uvgpn6XJIzXnzDWBIAdIuoG+U3OSCmt5EGEbUs5RTFf
u7Zs8PLh0WlTNAjU/Myg7gH8C9lJTrzf3Y2baXNUCdwkZTCj7r0S2sd/TUhSFA7n
iNY8rICXg5nX5yJzX85TD6ScJqxj65PGj3VbUrnhCtAhxms6KQ7q6fswUVYBuQgn
2VC5BGN80m5ip/ETlREVH4hKdRWmfw5qHUU02tPI1czrHPKdQKoLe1z5TOYtTgTf
ID3kTJworyV4Ggd7H4s2GpGiXMnHbGmzjJ1+hI/7ngHrCxbPv/Mu6nHoyZwUaxL1
on6GB0l628A5VdQGYmVHoO64MsrFIuc/25i+g1yf53Go1SJUTomuze5/HOqGLMxk
L0HWS05YE5fc6uOdEz22at6824gZxKBsEHIqM26s+PMqO/g+boK9NajJzsgtRwI6
0mgFmIPkdW3k47bE54vS1xwdvZen3LM8IB8r2aBjYm4MRAB1lNn/w2QDZTLFmUxx
5B+gio82YRO2c67qHxa+WlSBL3dQKKgC9OlhsW6N2402lhu84mGACjzgEbdzFvhp
mDLvza4JbEzEBH1i8QSB8o2u111EHK8R6yR0XlRyTdp2isE13DS40XSdFAzEerXF
/F6xB1pAglyub6M6zQE7iEYWvbgWJee9STl3Sj/syDze+ZqCeFYjktuEAP1xA2rb
rHcJmBpTZrNkPrYN+/dVTHKu2kkx0syk1UjZYTJZx2xUHFh1Aoq65iI1c5GNUGPG
2xmZHEzZit+j9Ck8O+qt/KDp3OYiduCd6Hj5N4G4v9oNILiLHIfN4AfcnbKgwNnH
ZYV0M7uECPgkzjO/Hit815Ehthpajrj3e95opFk0e/2o2LzTKBlYt12uHR/8SF5Q
TGYXSrNaIrkJg35U4XyaLrcNK85BPwGGbV1bVCJonm8Iz19iRj6p3+fuQbyOsLtP
MIBI3hHbTzxJslhAZg8gg0L4vpKU1/l8ew+PUp7INzukUjOlLY3GES4xb5S1X1s2
gLDvNDShE1vTi+6lC/BaTM4T6DZu9qaqYPJ6Ee/w56wxuwkawsCAjRFAu9JueH1T
JNtr33zc7125bQOm0rlcb2FNXTxou3vh50V5FOOhMQzn3G2ohcnWYiKEkH4MbVhP
Y8+i3iC02JwjhoCgNRpZSXuv2EGLHx5k/zEu+RvCeifo1Xq/s7Z6gEWCVvFQcrXH
Yc5iMbF9LkGD/u/f3X4QJRn2prjzBZco9gDcrSXhaCWuP0QLcI5jiDgGxrRZxbPz
6nmNqz7rCarxvTBgKir0hj68y5tf1wmhVuHQ3bOC4WVMrRtuk9d+ae47f+P5VXRT
0wXl3G5PjZJ/X1le1sLt7juwJg6ghe/bxCTK3bonCrZOgrRC8BC3GQ+UsHyqZX2r
z6L+WLgDKaWDW+qbJnAoew5IPuZ43H13ZV2c9wQ24SOJPW8gd7K12+BfiWZ5AQK6
sa8SG6NYuNRwbKyKi0gdiyJviTtEjC8NmA3PAn6Z40XRZvsoVCOJz4cnTPoGJmbQ
oKNkg2Z13Sfpa3QoH9B2rR52S0ICpmsGTu6bgwGme4JEXgLqhvhwgwr6Rwl7SchK
Rc1oQWiGv8ab64MdpYFDuIUmZsYxmXpNF/4XDCkhwPka/JttSEUS3Vm6VPM09b5B
uJYb+B2Lwh0eTqFyHMnFYWG3DFM3q1rMVoPI17gdO27v5fn9/MNibdCDG5jcgA1Z
HQLHHUWMuvzzDPJVXfZAYU0lQWGrXcyVQFoj47Gc2/iF3iRZN4HxtZWEfBbwzT2V
d3MlemFnoxD2wx11AHOd8RoIJiB8pW0pqOfbb1nEWYn3ehZvHr86++P0j66EU91p
npwNGp5wWq80Oo0NIgFe8G/IoATW9IaCShqsfxDQ7bNmC+LpTMaVYZZ7wTct3oKh
DWRQ83f36rbuOdsdiXILCVdbvlxPJ/SmEdr9mnpLCsXoZxvBUeITwgyK/E7Y1qHA
PYJ0SAu3Ny5Yv9pcTUrr/lUpo3ZPf2TPEIuEJphESXLYQb9O3SodU42m57SU7K79
Pf7aNdtRfKrt2x/L+jWWKiuvP7LAFs+k80v4swahEmksPd3C7li1XxgCYepku1q3
yVHqutgSRE1vagxMQnZaa3yBrGa9T64v0VF2bgYwmTW1ha1+F27vuvxBe5Dyuaz1
rfVdnuPdcoO8KKxUQCrDdsOAsSLjMdoNLD7HZpYov9TKrGgvAMcpM8/V0578vwXN
1ykJYyEdre39EeFfLrltWHmbc1Hc14Rle8OvgAXsVb8MUu91aX98RfgN944LcmsX
JMMq4mDjzlZ8T1BlbpDke9ho++gezqUaYM2sC1VRwE1q4BpBL6FpflpgeH/lVmFo
y+mkeUn4KsSmYm6a83NHG/Ol1URFZZc/coEj5+JF/I+O+euh9Zsjsoajcwex0DZy
mm/9augD/vqArM/C3LCBjUP9cEB/sICojBs78xgkvgPGjnqlGXpldlQzJt3ro2g/
GaOsTVB2jX4zWIWBjYVAeep1AJMSutsjtG8NAtCxjTSmEzCm2iB/ZBky9sz3pFY7
rZE5vtl4hrDYACtlNCDXdHcrH5yLncH3CMcP8KJQT88bEJxFpCy1/lOhLyVKwJG8
+8SIWQlpyWUkkQwGmUlB+zsTkOwen1RFngU5zZA1pq92CgZuu2cRIvgVh3XMII+2
SewJ3Jw/sk2j1TbcwWT+Ex32uGKMFoB8zUwgLh7bqupqMIfRmJwxGhBTVJ9mkS2m
zfQJ70WOCuvjGeZerFr6LfP5sPsnEKu6sdHG1lJJdID7iFW1XDdvZIFVc27D23SY
LEcmz8/kO8SV44QLyWCXfpfkaTpumXiCDz9x4u5iZ/VETSmayMNShzZZUWHXCodX
fDUyrHjWXs+0/4xxwqSQ97WNpNXga45Q2YT4OhiafoMOsIfK8UFsGjwciQaMJb6v
9VtbXuyz4WuR2A9O8LF0JTGpQroVOjKo1u4SPCOkvgqUVd5BxGEOCZDBew5frJ0s
IT89kTNBPuBu8caQ/NeM5S1lBU4k/KHBiIUqvI0a8DmjPVTAuqOValGPMCO4YrVP
uRejXF9vcVdGh18Hgb+8vVJDlQCC90cpAPWK5JV6sOdzONRYjJBHubmjCELQUxxb
oH+GzCB0amsGeZ+VWg1Q/h1hx1BnzhBXmBcTKnpSpujnuMnSu0S4vW8Kfhq0dc3m
ZM6e689lFUIxdDVUlJW95RDe7IThoQ1bYtKsM4lSocO78lrtXWe1r72LQ3TBxpwr
GbF6T/egt09mvhaGuRVVBiTZF8Ynuxn7BXMC/vOQ6X6+mv/+8aAQM/IS+C2rhDUy
5xizAm3VFGqvfTWU3kCHjUCcS3edkE53ni4g++tFMHxz0F0jRPDBvZFiiRtn5kiK
xtcFRwGtxxbLelkj4ePxiAzU6EP9OcopK1lgLxrdeTV/Vg4ifpKbZfxQdmV8SNQc
VErVqQQf3A7S9UN/exWyewleACUdak1rAz+2vmsS5ZHw19721aCkQ64W1vbRmuYn
xuXRZPb+RB3tVvI1N6sbMoIvFIU7FqtujdryFYoe3UrzXV0nDFYXWmOjr6zS1G1Z
0Prg8+k5nGWsx6nS2UlJobIGBlHeY+n8pCPKkeTRBNy6k1h4241h/uURIvmCKKiR
cG6rDMJUJZ2PksoBA5xQF46oG1R74ssq4fRVjQWLN0uutmfUfKi4z4exiM/C9bzy
dKuTIstpbC1TWxHuZtbel3H7dCKl9JsIziCs10OKolLe7W+LOrJq2nZhGWnppnkL
XpMd0VgZvMz2vP1SFj28h3L2V4F3K9UADNEBcmS6F5XqwOEC4fG3IygMzBGyEWxd
kVvBNAktNwb7u0CogDJOyl0yqA7k/6f1iI9cCmOrS1PAUM2WZ7ft2m7CH8BnmY27
H9/ExM1UAHfeYWv7MbICYq84BEZCYTKSRLwLVD+R6NAhcySCe/RK2l//ARg7NQwj
5/cWmJpWQMr8/Di/Tz5xvse01ExRVur/jQw1MM32+fejO9vKHPkM4/MTOG9TmxLj
G0dFLTDG98XjrN4qk5OGvKW6nmiDgfoMn8xDgdA8dG8qZF1P9hSW+Q2WjNeAx6FW
2kOUGrpHJNdbGJJnCkkKhIvep249/UfVGJEoTtdkA6yKYmg6O0GpBaUBPYAmAk3y
23Y2bpljtvsEA4BtTPnSF0tdwgcmi4c1+OzsyD29hHblDLD6O7Q81COfqS5I1p2Q
C8FPrdSVotmuNCOPnOFyiZfx3U1cTwTUrjsfxVdcBiUsnD2joBeB9/sbEV3b3TTx
JRLY+8jJdrbCpKNOrzBnu59LE6qlan0RlA7eZHA77fL0SM9gx4FQJWu/4QO+4IT8
tmt521uIdZ90uJ8ilr+ZKyQw9jknpoLhuO7LREcfBNNklArv/yXO3IXm0C8cJJob
QgXmRmHxQpWiXbfcIiOGoFwra8/cWfML/tspkTuiYjpJAK7TyMQqHFzB8gWi61wi
M0U9s1zc9NUeajq2uDVD2mOhC5L7R6vuosHzpUQOi+C+OvdlE0OvmSBx74NO2iPk
G2+KFOGOKZYkhM1fE7LWeKB9gsKlXu5psQXg5qMR3mbjxKYkuSthLJZwUJGs8Ao+
imf8cCL4o0ek/oApjEOhporDL5MvDXvr6SA5Gm9XTzbKK6WfznbluqXhLRJDi2yt
9j/KvzpgKe9ZHdZIUMsnYM06UXIbI7DpJjAkDhkExgFlGU83InoSOhx5scaqZ6Kn
d1MXYlvwkNjNUlhUp6zUR8nsk5riXxKRcOpGMsBYLlKRASbk7sxMswuUL8YUEL16
MceGpROOM0u9+mlYkCr7U+FFEAzITQAGee7ie2qRfSJYCagws0f21Rl4jncMacM8
en44KsF78mNkR66G6KXXp0FZVA/JGpYZCFhs3Y3czVU7Hc3o05SwlzmBEFdNiwVO
YMqI2kS96rBIaEXEjwuye1vyBqUOeAI5AY0IXnIE4A3UcBzlP5Kde9eMuyupcWde
JDr8ENbuhzXGE5mZWYprzctxD7b2l+tKrOIQq9b4Yf3K0+Z8yXLW0284jBj8s/O9
0KYKgYpQcuipDm643t5LfUus0ySr1lQP7KJBxOFZncTwgMjLFMSjCffwVmYCRr9Y
e6JymlHfL2EDKnnyxewq/sm04vp4247yEUTPB6fSkhgcp2Bc/v6/bpVfoWZORS6D
r8E7t6DhQjsMkfelk9G9Bik8507ns9hTZITGWbq3K6e7BSdn/TqLgfCcC+q7PSR/
6MGhiP/yIj/Q8BQWPr7BkP7vJGulDCjaBHahYvKKbLlWDbSIi+I2irHBJXmtWBRf
XDju2Dbyz5in/CdxW5cUMo5ZXh+nKSsH46cPK6g2wfXV6VTjL2a6NmJnYaWwc/TO
I3cM8+uYpU4KDn9WMzUqs0zJ8M40kSVtsTnP1IcZbYS2Qgu3mzDO/6GrUdMR2rqN
XWnDn0PRL1L9agn0gkn3lnRpXTt6eVgAk5ujIeVpSUoClgRz6UBBzq8+IQ8stAwW
8nBElWkzf0MUDern4fi6pqtcHLi0etOw0aw/g9tyWBfFxIdPDtsdQkpxzuakLF0a
vNv7md7L0ns8PA92+vZ0OAzmY1mHA6h1sOzsnKvFx25NIyMIYV5WLNlDwAsGdw2/
E5OwHU106tCdYsUf2SHOil9nOi/Cbhwtp5vh7MVdvkYBrwK5bqlSD8yonjFEypPY
za8GScE8ZJofag3BuIoYi5Zp7wRjQ4eaOhH0c3S2TsU94CXWRSXszY+/PGeUsxoq
V/N473NX+VXPXA7hgDX0VrTZLumYromzagmR4v7cZU+ZTo27Ns7fd8IrEDhgGaBj
STLE09JSgAufPX8aQZClDFeAXUfExPqb/0y01vDziknTNuR/XB/gsVBdRsZD+KQ7
oYQzbxZZ4ZsWZIc8t8F8EFY3bnyt1MLh7a6H0G5uD0rIL4qvXdetAXnVjOIHokKJ
vZm2RP+cmof/+82H6L0Z4fDeCkGh6NEDTjiz3B97p/PDna9oeZxdFlMINPXlC/tm
t4awKlNnkv4P7bWtC3iqpj6el9Bc/VbE33rymY1hlepYFMRkc8IqyoIspmlQ8poL
+BgieyOqnHzuffdY1GkFPNDUiZcQ9hMP/m3vESsoFZpC9ceLeJvrNNarHBGi1h2E
CEzaIs5gFjBNsKeG1Kf8D6RZjLUzuWCcCmzyFs0DQ0vrAU3+RXYRWIJLnh/G/uY9
ATo7JkH1BzL/zm2KGE3ZF2ZKzn2cNUNexxCGH8bLgYcdRE4HCXPcnOfeCULyaWzE
4sJhkXvF2nNgodkjUn4zZ1z6bILkpHND791YDQn+yz28bbOT+JCetQRAnbiPHXQZ
J6xDlYUoQ5F5zQ8tFV/zkyfeYCJpop7Wf2v9Xe+B6YLQYkUeRi32tO0zT3f7jKVp
HTT1CBoMWfv7Q6b8Xl90/mCRnyc26f6XFJR6ckBuquIu0lh1QvszFj2uZJ1p0oqb
xIY1Ak057RJGb96Khr/o1/xkX80yAiZDw/9Ovqe+59l3s4BIokYLgaC1Ek+dUYis
gzwLbfy2lwYeHIOjycUDzjmBbzzIoYpcXxpKP15WYuCMZjMz2cfLLjamEpDHrTEQ
Jab7cprIjjrRW0s0BuNSeZ6qjz1rlGo9TeeKEIMRI/0fRIc5Weo4ZeKCdUNdhavP
Zuh9EW4WhX/gEEUwIn/8Q/ptHXZ+FmEXkTzglpzLJStbCMZGrnmOw7J814ct0Jxl
XW0fMzrNSVEg8+Xdl/3fBKF1ozpNyRFkW7rCjNXOhSDKaT0iruVRkHdhnp/rAqIX
9owOI7+L0xoqNC69ccKZWNNQh7fVyXqd/Bbl6vMO3rVOiR+7GoZxKtMjLdW8xDrY
cQe3yfwd6agOMDRMBnePZAhKnYVjrWIHKwDkMsVjvHw+WYUfxvKYASC7fZnaH6+T
dHg9ULSnzp23EJYnGnzEjryhMVXW+4mg50eXXKwQ0R2anV38gttR5+ufxrWMJAQx
X8zH1PriHZCmEaltW9vheKoRk2Yi4posYAUemu03poRmXsV4PwVXCXmDGgTHYPNY
gwGTU0HwKiiV6o/UEz77VqnnLrWvY8ZAucYd/mCUYrMzajrHAz+1B1N/uTjVgEFV
liko55atCPxD0iEGzg2VIBG9zK1rqr8yrYBZQYPEvikoTnyc8zshQRebMVY7rA5A
xCIJqZ+djRz57KQ6VYFK0UG84dO7UsTPbPKaih77zn1YxxRRBg534zD9HnA3hVOM
qMLla3Lc+zqVrPz2q9KT4+v8v1bcLKNRxdfuRzNy/e/Bao7uoK+pmWWj2hmNNFV4
87r7AcwWTjw08coPTBq2Zy+PjuRDh9H1qZ2H5eP46LX5oXqt4e6nJ9JdswyTbsAv
wCa3Y7wpFzp5YMAm9ZmCBuWZJHkVBHmSqV64kDJgK5JOQs0Wv1RqbfGVNWoCYYa4
1d+W+jUZGahaU3PdMfjqcrv+5Yy7j1aRwsygWViuFen38x0ZA/t617QOT9GnTFAG
+bZ3Wbf/WCdEqaB6EFx3/tJg70KCJGdLBooT1PDeBsREZY3aXXMgS/eRJVtLVGVl
OYLGd3oULTa6lkLGm28CbZVUcnjwqieZxnQHVoF0yU9Yn6R1nP6amIa+PRMN+oMX
ex7Xpb6nosdiFS2L7iyb8WBeh1ExRJF/lmx9DQ4BMlQCz8T8dpBZ0Zern2zybr4Y
Tmc9dMpbyM1ACg5gipTS/3e+ihQKofQ41kaYY/ER+k4G7qOZ2wc9/e6DOcTcDsUN
ZRjaNC8Bx5uUCf9eOUPQVagEsJMpn+0JDq490F3ErwFTs3ZUQ3eIEm10qftERLR3
mxBUTFcleyPk5DTcGOteyHJT6hwx70mRJ36KB55OV7AM/bnXfMQyY1DOM6/vnxVh
lWNwccs2jOUHGHZztc1WraElOVruaUMlNhYclUsdOjn/cc8que5VgR2pZwEOnGBo
Z7c2lSC5rH23ppVydJjPj6q4wD/s0mqwYkbPmw7v7Ah25RkLA3FYyJrbbc61YRWq
ZPd8VsTnv/la9Hjl6FiCIixmS7j71USv8rtYlORB+/iBlXoQ+PXtdvfcSblO2R2g
Bkgt1/N5RUJGOaveXg32yVihzEXZSC98pNvTR0DzffoIpfBe3J4nukmO9/gDqOIe
+kE1nXMcBxg2hUnAp3ww8gcmGNxn4CoMHo7ZFDwFeArwKAQnt2hwf47Ysa1aTulV
ZvzMpG9E/WWsBT3i6hhwEyvJ7fgGd+RE2YeCAUTOu46Y2FGMgF0TXHyWf5suj+pX
jtMvApLhoxRgHATYIxsctiMe4LHCzIlipkNlSJ3my9jioWYZP7Fw6GMuRMSATMIg
B9X55vhv0eLL7GE7M12Rdg+H3XnSUhAxwlXXIrjYpbux3+KBRZdAX5LPDJod2cZ6
Zqb579PGLPZ1NEzOxHhIDYORpijDGMzzISyUhc1yU3y3FgXVg0S9LCTJL1s0r2oC
Xn/dODfxle3eqL4AFFucuQcrQ4Ot6W5IcpQ3gCPAzKbj8GgKvTfTdfNE/TMejD+J
50vEf9UE6/SVdIl7Prb1WJBgVDCEMFqWUr0ztsSMn8P0yII0oZzsqtcyJu/KiyBf
ubffwkF2BmVfTKyJDTWvfxp8Y4W5OQiz9qd4o0kfsXe+na3rE4/FlYE7i4N++hkB
QMLtpEw7VdnTKA0bonM/Je+ziEkmamaRPC6sNWyBTHqewkcGPROcSZ7Fv8tuArbY
TqUNxkLsYHNTFF2MJAQdy+QMTXdFCwsqjdcKQycboWrfhp4S7LNPF0ND957isx/a
Xd1enYbha4EMLSvhEeL5xQ4jb4ZKFwLGM7inwXhX1sHGyOhvUbD7tIVoRP0VsQ5s
VDc9Lkh6dqa54gwIHpf2l0gzbl0rAeHXZh3Js6Hq8o9c7aIfIbBMUeaumzsS3lGL
MDS+ALpOXBT5GOi0JiSvHMSp6N4SOhPKYmo0PPXs+6grp+9vo35RnedantKOAccg
ghnB3kAbaMMSRCcvAb9urH5LPnfwjEAOU8D0fwILks4StZhiDCpP4hk5CYwUIIe4
rvsASqX8ZlSVDy9ajhmgo0H65XAl8JKw1d+cRaQoaWyYzbfdlG37seq4aFWU2EQ/
fKtTwRNSs9RSh9HbAPAu+WTeWvs45qbcNNfLBLHfljQGeEBkuQwqjNzhwluRXOP4
miV8vnQMVyIFZIXAtKXr5KVwDGFA5050Gke8m2UW+NKuEzqFrJ1jBbuLUGd2VG9S
u1EK+mghkeIpfytmLxf66QSLv1Z0fbYXfKpbWoUoMzpSwRJ5l9Jtn/RtV6uK6z9j
IG+/YIRSGla23D8aVI7ulu8TKw8BBMMbUJnIVxFew/8j5Y1YuafXS9Be6hkpTUN1
k8lGK7aYIQzZBCr3+aYEBn7uTO+6NItcOUPXJiuC5ENXVWBnaa+hWO8VQu2oqF8u
g08Bn0jsKHzUGiYOdSpxAd6MToKmx96/BtJqHCCbAkSRoccSPQQdNxSOPiGX+pe8
qp/U1EiFEjUF9gcpcNS/aSnqmtODuqDrPkRPNyET8hmAx+OlnzfukQlJ90z6RzbW
WU/BAruxHJ0F3oo6N76qTFSJSriT9vpirDCN5hjFy+RbeBTVLYXHK/Yfj7DJrAR3
kQgKz6wjGHhQVIjbJd02aZPw61ElrMygKOL0E3N8iit3jhKVqgAg55DtpV12xnnW
3T8NnaJCEH5D/rgvCR+AdCqBCf7f6PTHIytD5erYW7bRdzyPViRMc/shhMozojFH
3kXY+/y8sbnOjoqqzqNdGMN/N6iT+LLv0e7zuAFhrZi3nDPLIUENXARv8tkUwM2o
vyz8RQuj8Ki71gkFUAKj9kjRXfRdqA/dC9bALjCxY9O9G6q/cPzkr8fogc67mgi+
OMAqAM9qvx3BL0xhUtWbjgwrNkf1ZmYVHbJoQgxCQSniuTDWxENL9DkrGJE40Ptg
mVIekEsqmWKsp/+R9Sfpjpq0tHKcHXCpBUNGN1wANRT/wY8YBs6axfIkSlSfhFL8
lrwwM7SuFg8hJzG4tni00qrE9NmbQNfemQuyxIi+EX2NJyy/8uH6dbWhvvpW4bOl
SW/VQwaCTuaLCx1gXIXoLbL6bsmwyiJxatMqd7JsMQFEgFGBQ9BdC79/e10xRB0L
CGhTn7hyjuiqDlfaeiS6sJLHOQeObxjpVLzS2mp6ZPK17aQz2cLeI+WUTPK3/uiU
SV8rhCmiPuUYnC56oiXTZyIgpSiEQYjwszuD5d5cLC95TwXXGMbOeDvZqP/z4ILF
7Iaa5Z2c4UV8jztUsgFata3f4qm8B7q7IBfa1z+nISvJ1ZNlzR7P/+utuPf6DXAq
SYIJ0JD0907alL+4Q7pUxFu70/4EVrOzMzFx9NqNU6NGgMoy4PswCGsdC3R3v3Ne
F0hQmURqXIgc1WyCAZftUY5x3ZP2zABCzInYxpwexqscRSYlnmgEd0r6/pogxUZc
uLBVc2Up0NcoLSxs1bb2tXo9dOoTUlE45Ex8bHVLMNre45sPWM7ve/cJt04fhO3M
mZm7Jal98gwGwHOsbZkl7lJtQVxKaBe4VH+9iybi/TXJrwmAuKcWhUuNH7htQHOy
KcaF5PZyujrm0owo2vl1J7ZDyVRuRlANkR8vVo8PSFb2hVWitPa/V9FBhO4+zRL6
ksS9MBX0lyjUVZvaetVYyRTwwgz+nba4AKWJWETQKRetY27HraRhdD+RuKy9Sb3T
JNd53+LquDcc/0nSBFVsQVzGohH0zqRhGI562uXWoib5DfE9tizFnzOxDAKCJCVv
elnmi1yhBoJRDmzWCxGnZAMsOGtbgkcP/VhO+djJIdcFsNyx5NSiEWOUk4jF2RCT
5vIGq7Pqh1dZsO3cz3/UGlXnAFgGQNa7+fGlvog3VJSC7pxRdcEwAmwSXegAaFon
5qcCbARXlbxQOrFcG07hxLXuLsfOsRKpu/shUA6p8VJt2fKvzrSbmoxU6Z+nsItS
FQdqlvT2ztu20tEXYovHG5S5NqhRLBAcoZHZglJ8PqvaaN7yKbFIF82WtYDezbM8
18FZBo2q+z/hLoCS7yk1OHbnfHBKRs6g6bwnqFrzcDpyH19eRa0Kf4WYhUCC9gU1
+QzdfJTnOqQsRBrWiixdK9Ly1zQT81y6yTqrx8k9gB7IJb0yGayb4z69WBYJEthR
sObDfFAFPl/ElvAJNFWoIYIAfUmMGA5STgP2MY+HbDJM41Ytcka/BqN8+mSsq2sk
cGSfzih9HP3wkQEIdWjl85ZLZ8PSRRUjzutXf/vggXArB1/U9ck8z3l6BlrBDxT9
LWdRjMue/4LBgOnmy34iOQ6HRJJ8jhf/+ssyWOfmjJ2pJI9UldASusftz16UiKTK
HxMObT3mLMi3HFnbLDW2SJnsJAl01PU6lW4mtY6T4sxU46EZg3qT41dpsy6PY8x/
lKjXHnr00VmiutZHzNLfyfhdLOspRJ6ehCxAt/HpFvR74trV6P/TbaaZDheOymy0
6hiKeCDrUn00FAYJABcK38d820+SRvGuTIcR6pqQKts1TZyZfXDyZvY3KGAsc7sO
IrR0XhQg8iEBgzhYHUaCpVjyQCWQjoDgejiITKFn8BPE2lFXbaQB/Z4KgekWz5+9
6rSQ2TUv4vDqi1sct9zehxtvJN8w3pdMMN87qB6SgHkAv+NBgqVnycZn2dEuA/7h
cmC5NezNmsT2wtsZvcwQBNGrqBg9VmdYrHaNL6WVg70Y/u0lPMQCmHHOKW8Jna0Z
ncQ5yn4s08jq3RijK0HLlkLzNZyd9VsXBwTD2HXX1Rv37eK15W+8OmzMwGCQqHJo
SN9PFvj0JgaLcRmOeFwZQo6ekuonpWBby5s6mJTZVuSy8NWXnL8g8nbmXrzKUIBB
rH1P6UaLLzBo01cKClmJa/1YnfeU9d6S3o1wEdCLxV3FYVpXbSwbOn8OZluW8wTa
ndyx+Yntmc+eS6StKv/9YMTxSHej0Dw7dfRxXWdiXlWv52yx5fyPXXbQmqSIqhkx
CY9BMkzxcXtLh/yJdMCrPj6WgmEcFkyJAdJ5YUyi1JvV9jpczHIB/bSBdokr70+M
aJ5pSH2eYOmUgXLqZACbI776rzHYvsBE9REyMrKbNexO1NSwF3BX6ZO7zeVlie+V
IUgGH/uD2QRixVb+JoSTaGgrUdca+oKgzkPRGQQaVhzTonQCL15Gn/g98sJm/DwO
NTuRdkvfElMgZO/1X90EUPRtrYySrxGB/Zpue1kuy73e+9fk2ZB8SonwYYBUQ6r5
hDwEBQB9aovqlgZCyJw7u+ejMKuJQRZyQoeKZ8mYXoAHNHk4ESbrILtHyYpji72o
etg1lVum49CLSRrzeDMXz6IOLHzfp3etE6Xy2YtVPGjLkwWvzPSdvxivyXRoPQ2F
mg8ztm9OQg8kKDPTG6LIGSzKW70mxnXVoys3Ps3z3nqgTnZ4YbaprU41oGn+Lj8Z
Zp+7RhhbTyT4Y/9AHhn/CnH9Ore4OwDwWzbitw0M0xGV6ZeUzcF4RmtlR1bnYIOG
wvVJVt/r7vMsBiz+kPYh8EiCZuvaK5fE5yyfEwFXUXVSHqZ6grf6HMvdp4IY6BmX
pZCabo4UXCBbxPASEkjV3hyMVV6EGL/g/21aZBCoP4wQtoOgFJkG9zMrUYJ7Rceq
dJjPffz/AHwk40iEw/Dw2RS3jbFwmtRcqwgble+scpD/S6nsXoLdkyAUI2p3oGAr
vctiDFqvrvlERrsOz4Rr9dFcT0XFHzgbrfQD0aVpwhUl8xrgA4iJ4UbVxU8/aucF
YqQpEIn/Y8DFwMUji5Xgm3DIcQGCFZr5LcGSCYOXt0iICDqUY/fLZXV1P6JhW9Rg
8kvKmgh3Zs+k8d3Ks2NudWEQQJWcVjzxXv3x6MJCSwmEvASiBzuTAm4eUzHUyot1
Crj0XR/MKGbUSWTpzTCLlsBHwi+5YXNjqG9FJRMYHvTyfnIEJ6gLsqppDcsraWGs
lg+OwFSuCEjph78T4E+LXszTPPQpbDk6mPrYUaVYxYRoc/kY/ZXx/KSlpvMVNTHh
hRaUmguEiEQuSsu/2AnNb9ZRVBxJ7etzLi/S8+rpuV11TAFA4lgdJOITvG0aKAsT
q7r64fxDPGc75wyMFX9wJx8SEL02NcQ5FroBB3xsoE/b4NEHy7FLSEZ3fCCvlNx+
HHB6E9QJcjY3YjvutyfP8rtxiQzLmdxhMuf55KYKdkUmEDrSVCqvZi7DXMYr81zg
93Xar9sylfUfz5jb8sidKNzcsFTwAB4ooITgZP4yfOSqua5PIB4UEdSgb3iLtPMu
QSWMVNHgUl3yTT70FmigSkqQMGIPHRCr6QFJs62aoqfOttzAnp2GXqwCeCBHSECC
i50yGdAgAk7b/5pNuydLzL5m9C+U9QOJGL6Vz8vJ1XERs4RAux6d7BtjVVPNWpvZ
KpR3DFMxhxdl9Klw7ePnM4z8QXJTBRjW4fylzYf936oetFtU05i7RgS3BjVHtH34
1SHMd6eb5RNiKQUTpvWmtLIAwOxkUKvD43XyWASqeH+oXHv1x+XR7LDC8671sKsQ
qB2xD5NmaK5i4vUzF4pNAAYu8/Hn5nrva5JCxarl/aUNiRFz+JrXLCWwwOyi4lpS
CcWKarjC8HA78DZysd7YDJI77Xb3ZmmmrBCAvLYBClghhzIYjKeHt27/pNuKbH0i
DKajmFdjwPH93TPht/Bvc8/DEVmdM1AqmkWAgig+4oEQZdiPPEAAgE7njfgOWEHC
cQD0rPBxhQDisWuqtvFgIRkcOQCiXhk13Z4w1kRa5EXF/bctnQeqJvhNhpj5EAML
OZhvp/pPv3K+LVjARzEBB0MEEoDS6a+8JnRDmXUOQ1l8ga/PlCQArD5fplSGcjdn
nInc5fpVsceXtgAFoyvouME+oRA+qEQFjtXBkqxj0XORcpvHwZr3YKA1hbfMV8Xi
9aTQ3SNdNk7Vrn6y/xyXLSVuK2VW5CEncHxeZSyWMpBVP1qLnElMA6gLVuteqalf
qAueHC25Ik4XmE5LesftjY3DhW5OR/oOxWIAAZBv7SWvRJ1IVR5hyAY5LVfFXqqY
S/ULa+Ey/3KuWQ8Laj2Vdk3YsBp+KFpEGpw9rbBh1krS+75H4HwD8gA99tfOcvq+
EBCdp1K9HHZYqdeaOqCcxZC9UlAZv3/nbbiZzrFDFdV3erw6EkvoS/AC0lu+UTQ8
CKl3cSDlUsUHvUastRHTaEBvLkf8xZc4kTlybV55i7UbINXiRtqOxw/Hoo+7TrGo
VdRh3qdnNFofQ5sMlAOYLDj8QUk6E47S45XKNZr+quzTBP6Gp5aEYA4n0oAFz3Dt
2jiPl6DrpfAvSxc8d7SwRAjryOf6Do4mL0xhI1cuZemcsVPviON3Zs73bh2GHLCB
ofUXFaHjEAyqZJ5xLbF4ieLjayD3Fvf7XQSxVeBohbDV36QgeI52fFVezY+ZqdMl
O94rNYfmrP5CvHnFJ4vQ1eQOR3agZIs9BrkWFpGTLJ/P54WDimEHRfd5STlsO/hw
e1bIEHGNvfEGXt+lSorcMq5Gvy3Mx42n10nFfcnsmUFbl/8r6WK4Z/2X3ruDYJnT
Ir3g/BBFanNaycoYjNMTUMpLRHkAlEo5o0wAzDzifk7E9GWpWDeylLTwVEZJdtKy
7+wXiRaQjANcqFXINcMiVj7q+He+clo4J0jr3FSNv0pdkltICIXXbt52/o+kdCJy
gXHlssrkqD2Qfc5VudbzjGF3hAsphxGfPLiWahJJhmd2n8bKKM2xv1itb170V+xu
tk6y5x4oeotFk/eczS7GpCxYf9XTCn700fOTmUganyOFiperr0+Fa7PN/Aa8hOdC
SvzrZM9WfeWwlMlkYe3Pf9mB11xgZV0lzR9Il9dvdZj1Wv/rgp6crUepiR8RL8+k
tk8bmKzs5Yn8WroP3FwIyv8AkKEXatSvPMoapvSkh4D5R3zDflSviwsbtgi9kEq+
b4GGbxO+aQp4NsfkHdes5s/mL1gifw4cKtmVGQlwBSO4h++RQCq5yk/qLEGhBVc5
9pzaT7r3W7Sff3Ab2IH1MqeT9e4RjuvDze2LrE8oeQcx2zOzI3cQBz09TlTbHkpT
oFbJU5MS8R5FEdwTTGSkmqj1f9Uv2i5vFArAV3imYaLTLU2Ql/R/zOGnjhj/cx7L
tPSKaN0qCiNRO+VdDul3foh7psJd0y1P0o9jiHp8J/jcZGRM4/0k2OBInVGDN1rh
Z+yc80bVgAb0MzEDyoHGnwhbb94US3YT0ElcST2eJO4pbwfc63XOOnoZ9TRje0iR
lYhKcDrRasNoDCCsxAg5iM/LYyT4ibp119BQwkq7KcxkdzmZG0hSvbuHVgdza/gg
VdVYdCCp5HiFKwL6K6Sw/Arb8TrtNTQlSyH6hhh/M5nks/qMH2+/2peBXtx520JZ
8vqTHFVYJtNLK2REB0pqNuDtEXx8e0jY5E0v7BME5/0d0u6nLtQp7fHGjbxcn6L7
0P2wQ6OdQESl6Fo+KJ6dHKySl5qYpssqIZRqqPzJyNZcG2/gJ5krSjq7lzlpkSml
SxPVNjqZA9pN3jJPM8/CDq9jNm/N39vXuapkF8TCyV/MzmTGZV3F1DAyU/IH7Sns
+0XuFhFzHiJnQIfgWjQJRTCvN+8ny/GAf0L6H8PDXPtIv7xLDFkIZNppHqpxhZ92
n/mIXQxeWpgVLRO7+Wlue5waQLDPUO0aJqnf6JvLXxxSLh34Z5H4YEB7Gbwx4/rt
Jw6P0azy0VTpYP1QctHc/zS50l+7gQCfsUI1SzE9qTwocoMgDX/ZPTGm1LCpSfbM
rSkwSyT1CiLUftsL4KOEltDoYS1dPASmEBgljVN+WBIB26O2qANLh6oJAmaxTURv
PBhF3BxRT45auTirb8+xqQhEsfmEvTU0G71zLHi1Vg1pQRIcFsQQzPTXV4upXXsm
YfbholBpbQ3aj7O0b3mNN0Sog0hm/mRvBIHQXYf1CGddCcObDJ1zLfIvLt6VSRlJ
jW8HHZVK6tEB+/oyszhcK5t558/27jz2CsW0Wu1cE8N64w8wp9KNDETIBH0VL0b9
KAXKHYzQONes7lCRP204e3k1+h24P1bZpbrfuQZGaMfjaEVMkMjGS1tr0ffVKQnZ
voVULWsiZ9pvV7F6tKn2YjEseCaWuRW8Y/JPFpU0puJ4ylbWdgoZAGfbhmGnaOPm
FaaWAIXbnLP7laJKU5DPri6SMtrucY3IEpFKRLL6hTvoLxlEjO/g3OIY8Ir/heJd
4gd5Zb3t+iiHOT+5/CX8JC+5gSrOalH3qk8ST190qNbRkAlKORwJrqGZDlw4vDgh
sBLOWklnLGo4YcE7Nu/bkspJ3zCSRL8FFtPjx/RlDfWROIG9lxXayR3DvDbUhK/H
TbnWDl2h5C1qMx1t88jfGE6lYPLcDDi0O6k2KseWw3WU4KqV+L+SDg7f7n0ypuTd
i+YmXNhsN6fCDSj+oevCqJ6NM5Y9wd9s2wwz2ZLxC23pTfYxOqhXrONuNvkVywc4
7Gip00AIMdsh7x9oAYDkK39pNuWlBzMX0TmskxL19Tt59omz0Qo22ICZrL6YLDPp
Nzfgw65rCzoewFvM44D8d+r1mIf3f0F4fpvz9TlOrqi0+/gMwUHYZU5r/Tdww8R0
Q1hCHtjFOIT/uZRA+Vz2QJD4eHKfqNu2zCELY/lx+u3mh9I+Yw+8jEDQOFUqUrTf
7lbo5owqABldiuxhDBCX/NK7qw8KARsyTETdmJxjqKs2eAgCudhSEuVAsUJS6CKB
lvbwCVf7alSLkn/K6aLfECZVZxdrDLRwa0EpJgfOUR0a5WhpARGpaOz18x6FrIdC
As0J0c7+eDF+tiiuLaJKn2L3VXbT4FkrnLcTNj552oFeZGnqqUJVJYOlVzrBCTGH
8QXmdLvzeYhFcDmlCrTY3ryaMy2cSO68MGMtbrK2J3+BfxTVnkgaLcU6ICzVD/Jg
L7xeP10Y5pxlVn/5mPFrwVNl5RRFGKHpB+VQcAAGIz6R5zV6RkwOXVrygsYoa6Qz
uPDdhGqxV5/5eWLA/waaVQ7EJ4Jlohdzgwk6h1kPURjxaC0LJXDoJm+PAfaYFtbA
aqYcXt9evYSxtHQKbuOqIcyx3pU/33OhkcZIZsQt/5/jZ2NhXnrHT8WNhPP+Gidp
X4+wiQgMelLvkMqA1cldcOv/aef0qP/hRMVp53nc/F62fAALxuv65b2oAN+UeFUd
Qe9s5jP9lMxudEpYKEirfEcXNJyxLEjJEUxilkSDsREfVfZeMI+zsp2UHGNs3IM5
U7bp0sVdDLFjpg/29kosp0+Ce+8UdkaeBXf3voPb07/m05CBv4vq3JMLfplC5/zF
c0RgJcIPpz+ry3A3a6DvHsrW3+Mofv8ZxfcYJAaXiVLjFOlr+pS+gdNTUKnXe2km
NgwroIUhykGSuO3rG5e2srr7OJEegaeaMzCV4GkZ9pSno1gsO6oRKwTEnGvZeJeV
/9coQZONUiRkp/RQM3NUIGHvOJk3pVXs+wVpSKexUr7ew+UqfrlUy/YZk75xKEoK
Ukh10HN6HssbX+T6jh4lsuThSFe9HdcwcgYnIjvpAeT1A6wfrjjipfKIhgl7M7cF
PmPiz+KklU8DipBDZTaCFx/Za5/d9PU1SI49eLmakak1YtCahXEmXV5IJZui7cHW
dMCap6WWI1/tSONjwooMPsGxlPTaynBIXIIE2J+hBc10EK1fyVlpGfEfUlbxp8De
btDZUC6SDiQRwlPA900I1pMCzSsKEYl+d0eDvWuPlQpfriHZ30173GyLA++VzTuf
eVDvXHKZGSwXelMciYeJMEnghV7AMmrwEQgYolSviB1z8zcnWknFEI6EY0hEo3+o
IyokatazWDoSvN63OCsD8gyubXv8sty6Z8O+K4P3QfGCggvuMETKRIigH28iQlMz
UcfGhZqDXHgX8mdqWU7y4mTvpgEjd47pUq/EtQE4479qiHS/L57C7yfZVIHs7e/f
5RrvTmoTN6RXSzAPEdkelzEs6J9BDBnoPdCtT+NZRBQhTMkOkZKwrK8JAArk/uH7
adWaGifDYjgR2HgZ13L/MrtLfSusksXZ2sBeQYo8KssIJ5s6pnuCnfkhipRyIBDJ
wn+nvh4kI3cGgLvz57EdNaicJqI4oZ9B9rnFncPWGFheJgoE/dVj7Bwqasizz7Od
87ivenO1/lYN2mHXPBGFF5JYXj+4+63+XduRsnz+d2JLM7kNLQyTUgs/ogKM7ypa
VrmtT8rwT4ff0yz+bWFQLtuajnZayScXGSnzZFNJ4Xq50mKlqaiG1XcQwF6FfzPz
eCIYmnW9mmjM8O2O27QsSvNxQZRk0b51adXNZ0AWKYbp9RRpZkl0NgbYnQhQf9+4
KoE3H2Q4xweKqgbmJPKq0mkzgEnIZ2zGesJK3GxIvhLHIWdXkU6x7LCqZf3yvlU3
AG7jESozLl6EFzEJ5LcrKyAt8I7qHMZC00JNbMMOLsFOAwS1XFZR8GFJBBBvgFqW
sxOxVvIgfqg9ykWSTRyHJumkIiR4QtTOtcvykLNb2+DTQNfjBu3VNvatIiMtNkV2
iAIvphZBQKACu5PhXrPzOV/KlyhhhQYU+Ntb/ydXubXz6BF9O4cUzM1Lmm0UszqK
5qVlEWYR3JWhHoHO5Tr1EW/9eW9CaZHYzQdV01Cv/j3w49fuJH2LEbCegbOfBgvD
fAGcA8HPffVsu9pODguycXY8RHputZSRI3ghFKS0gNMCi4lC93KaZGXlKKlWUavA
S8elFpiUdMBEcm+NpSd0v5eMCVAF+oCIchbJHbjVp2WWfCFVmC/pYcvextAcr3rG
7Mn9D+KTjyUyzidH03LtPt6K2p9N9yWzqoEenjqsB8fdwLXOkGpQWu96iLDfYZJR
l3UM/e9OFEinWq4YM+nkUeYaCpH25mWPwfhgDuOVyT5vSVAZdEu+6WhdfipBh67r
EeamU1baw2PwXj2MbQduhYNQYVylM6eRyaEn8ftUa/lwqgiP41dZschIq/xETF1P
LMLKZaUQejgwMqbj2q73DQl0IvVTKkp2nqcUhiOdK/eCoNFs7vB+GBO7BKmqSlqY
lSGxIS6MLRKaRlqK4cOqla3cgUNHjjX5puIFkwSVGTA/nsKaz0WRUxGoWBhoFAl+
IQuXmOG+gkwL2kdpg37+9PWjaI9ZmUbF8ywVaeNGjz0Y5WkBmWD6nSpWzqld8/XC
Oiic0HCLwnk+ZlLqYhWHJfZVEHZnqLS+E9dvT9SkD1M6JkU2uk4McLB2sXJS8Gl8
7l+wu6dzcOZXVv4R3UIa4xgVyW+i63GPKCE/LMVzEPNdNQombdM6cTFRq1QcZXlK
t9NqLdo/6x1f5FzKquyNY+2MzfV/VMNDGQP0jCjxayp+BSgAQpbH0LIZK0Ty1NdU
tVHNnUwci3wn7giHwBRQZTkSJNnWepTkHSBuGuDATRV5bsIDZ3tUURQxhsn1+P+J
NLtzooybK9cVS15fqzyFrmfnVnRmTwRqVQaGwbqWyyJpsLIc14cDZYV7meBZ5D+/
Go6gIHCwilibvEurj1VLNbeBc5j+AZp6J/e+4lR6lxcFkvYGvVnvBqcWi/xmS/qZ
YEr72hD2zGJKxijcD0t3bAjrP8Ep0l/mgatn8+Gn/nLd1/v7ZxugKYAudFyUUm81
kbuqL6p6tBVaDct+uYF+nDKsJh+B91fsb17Mo7AZOEFtnsN8aFs59vLjCu4ZUxXN
GlgCprTtmwvZoiwTYkVsR72jtA1nsYn508h8hEAntEJ3U6xLLUI3Ei7fVdb8Oxsm
ukBCjKr6tXeQlRIRseg3qk7P4icVuDnm1k2kDAvzD2VvMajNc2YmTCqPfTqFN52F
fa4BpnObWPchNifci70/WBDIajzvM6sVZGOnbHXTrzBN67T1leMUVVLtHr5IIUu1
nD/79TOyo87MFL2dCtcBoInSsgP2SZtUVtO+TNMPLOOgxjYTwArpSXYBePc9ral/
nxfoavQ3Pbfd4UqhTIFgEQwY9oB95rXEDxJee+oTAJwNnSO7bgWWKzJkn8ZEx0cT
OOLpVmHtpKpqeqVC2zGIraqYS2QU9vu1IGuiUCk5PIPahzVbBqt3io7c/2oZBtfR
bFsQstgdpst2EOgdJInkm8alPLxGQ6/5vEjpPi2vNQ+Xcifz7emt+kw7jv+egUMX
nfsXjPm/Vf2w8lPsL6zp91ZGqHgAUX7iPI7+BV2j8uqTBXyOmuiXhuB75bTUyCm8
86Tq05paWAuWyHsqUaCQmbFMS8LNj6AYpmQyy2OQa7v+9Q5OsPwxNnjev9W5t91L
AJqySKuQbQWatuIOJsp2x2Hy++ayMhyixELPQfLsebGkwImkqKFU1aBPwZq1vXRn
tccni06M+0qrozBVHTyAj3bKf04i/6xZ3kTAISzLYQDKku2ELxRL0RkaINGSeTgR
6NpEZxMssr64650dYG7nXuz563mitsTMDPplzM6h2n3jkDyrcmxWO8mxHoF9ojPg
KgKnDwoSepq2hSkJse1VtxQ1Ij1P+SH2xt9oO3nF/JVPV8p+tq6hY5O+RT/BuGap
0YZenOZbK2LBNGqRiauFvElqD5+Dso4pKQczPqY18j2l+YxJ5ZyFtOibvqvaT63l
CkPS6Cn9X/FujHbffl2qURNONKZf5daQoIwmUB1yL/Vwr6vzuPs9T738lY7lMiVd
yz4VxGNE87HEPMJYm62S2UNiccwrq5Z22jBgUC+KDY4cSsMZSMEV1W4p19z2AIFP
hPdFVO/Xi4rEPydjDkIs0OUVAa4fCDV8cryw03CBt2GZkdL7AQb6MEhYmXWvoO0g
txkxBrP8Xvv0dJxJoGcratHX1CEg4k3x+DvWtDuU00oNtPf14zBGdkTUk4rB8PXZ
Y1ELaace6U0s3UHKrDz4E0Uqd9JM0C3EYr5Vq+e6xGJeFT3l49XDqcWWw3Ae5dCn
loaYtPtTJ6R4kEMtS45VRyw+3NCDqoeNLEwRqQUQ/FU0bBi5LrRr+V6Dq7oiUf3Y
BVD+U2iCriHpZqywkqavKlo1uMUIqWsvf32zcswozSi6TIgZcSx8M9ZJrSCGsXT9
1RI4uk2VHb2wnNpV0h4md0qfuYdzc48t0L1uzM8d3s5kyWOGWjq+rI5W1+XYPrOr
FVSM/QssQ0qUW26ocm1MO5cJNAUPI1cG3KbrFYuIG9EHPwGI1CfopMQYmKAb0zie
1g4KWR+zmLQ5XdUA9j5YR2ZfQJu0weFBtcXB1kwte3XdQmZR9bzZc91Gswk4QpHm
0pPNeR45izQaE+Mmrm9Cm50/Y/w1Q5BNn91L8qiT2P8dnsZFeysDjSDxVcqtFjQ1
IPVVBZVSnz8w827x8rwdRlpAPuxcgG9mkfhmW23ZOfA2FnnPYq1logiRQU0NKMbJ
ZJSN9aDVmbXnm4XrlPWBRk+2aRqYsW13bC4TFv5uI2dnz+8KOnZ5x5h5epxUv83H
xa4qtAYhDIGhZQYQBfM+6Is2AuhT7/4cuxTOFcqdWoQydgBYPeiCv8/lG5kyYTDd
xC72XklnLrD3alnjw5tkINuJB8O2wfTkKr8q4QFiWpeyqxEtz+Pipq9esqxJ95e3
C+dbxUpjOOTxJYg6WnPCE8T+jp8qTyKniNqn/4efI03WTR7ANw8GpsDg5PzjM0SH
+NpMUwYFFAdf+HpFy3snm6kXL0ZX2ls7zXhdHLjoffM3lToh9KrAceTsenWiZDAL
GQoXXfihn0F3Fruc97qeu3+CzEVWnfPzI22hZ/Ue+GC6bLKvGYATVVipFVQPuY85
A5E0Vag1o87ol/xWSBn2mEjRNB5Wdm4X4TJsbWXQDW/EP7lNDKcclsamIMuxVHK2
312/zaK8UcOJo3wdQReVPpfNJ14avPAejQfWPlOoixjNg70hKO3MNWhwUYNK0ZxS
scUktS9dlkWFcVC+YkWH1cA3ENRPRTNA8KizuUaG0giGqs2fGk+9nabsfrvDym6I
SP2GbbAHME59PwZDvH2bILgP8DZn7J9F81mFotNW5FZrPTDfWVm6Att1ZDLp+BoU
Lat+YkokHrjxhzqY3P/CXLS80gY+bGl8Fs4VMmKBl8IGsWEFcwScAwa7k5njkVq/
dz+qE4qUehs4hsOUXF/J+tkBG0RiTfFxcRjMHx3CDsVi+u5l0BNcFcdUugIuGvU7
1fTFjD446xZI3vvjz+oc+qFCWbtGKa0G/JQac3wnAUmEBBTFIpHcR/7JcrzDk3ov
W3CwIraa21u2HDUMWbIRnurDXzZMPUUgqYokmddzBnHBs0oECgLfTEBSGYz5Efvz
EMXs7OKHaJgKWHLD10xmqACk6yrsBxVT+q/+nKRKxPLRXlAkqat45RNY8V/yvwfl
wD0f6a/BrbVVEx86qzLxkpXRcvP31/OCfCjVBR8My/0Z+Y+n+uTu9ZQPixnnmKcO
tH+Gw/Dwcg731DqkeQ5Z+aNslt/0qcH54tkFlnICHMCpdF0TVifP5eWWCpN7Gbt6
xeBSPR6jcoYct+w6DDIdeq82pSum847GEr51bmd4Q9H0dObjyGJMBsK4NEZUQtH/
CNDyERv/hAtgBhrArHXEeA9BAH//mqfrYTrc7iTADy6d2uQK7KEglCt19vnA3nRI
71lXXCtMbybpIzcnv4IPBnOm5GdGvch/9NiK35rQR/nSMK/eAJXzqo2+trERqv4F
Xu64kzUBT7yBxK+iL51D8XitQpTjQtUUzshebsgSqN86AojdjFDlAlf/P5gKqjXU
QYDDZnqnraZDD+hLAFk7sl5Byyk1uhizqcRdnpnnjrmmIhVAhhgv1k4OIz1pkb8V
tYqWTwOUHXF0nJYpqfzJ9RiUKymXei6o7aBMJ3GpZqFjtxkyY4FqBwJe1NHgTwfe
XXUYGPQeRgXA3QS/ze9F/OldD+/lMBJY3/F1oOAgpmW2v7BkQraoiWAvEloNn+Pw
aOz4vKcreQ69muRO+DBjaiiC0u4N402+KO5hWU2hi5wE4l62H7nN3kg1oIgAYRQm
cGfBicfAPjjqz9vXOLyRh+nvppbYrE5pndq7ijfe2ywb/UUkf+RuSHvOVvmOsFbN
jajQ/k0A1eJpTCmzwF4Hh16sRKwx38OYlUiJeeDq8nxOi0FUHyQVWPCkBOUX38on
obIjuHw/XcYRvnblR8eRYxAHqfoO7TJVU60VJMgsbHaJR6fvGWNnVqF+hf2Odq1D
MLsJY2NTQuJP8s4I0imqAgMB0/V9tEcCxnkpWcvV+7OCdL8XucMojc5H/6lJ/k1u
v/F+5kufAOD6oVgAJ+fMti56gv/oG7vlj7lZBpIEUjtGm0xxuVgNTD0yqyVY6PpP
Z8XT2c+XR59XeJmzelGd343M/A2FsAvEp7VtuDAiHwFU/GiFdR3wDL7EKP9jLHJj
NSVYYnw22s4Qa6c21yjQyeLgxYJebCuRECuxw9daIjRJOAuDgqtvaZbGoPPNNFpa
d91jAhb7ebS4L2HYUMEIwjT7GX8d0J8uhBXDk08Yb9ApBHDMpURpNAyWXQsIj/RV
CeAlPknVupboPH4fH87vLI1xyzhguXvjVtdOm4D6rCJh2z6i59fjqVehk+NAodam
oJW2ngeLsa585dU8ltueQO/uXOkrEGdDKk7x8x0AszbrjcQiGXjVyixl8GKfzXfR
rShay5/ciLNAsffeVyJ6pD4ydzARghCiNS8h79/fb7ik0IaH9/H7CTfpdNvaqYQ/
6s7MaGDC8Lq7mZEgeI1CRlP3gTp+MTo8JLVRVzAb9wh7D+onQ/rbvoSHwtkMTjFv
Js3baWwv9U819xW2NUNDMbg/u7VDUn6REgglzMpjb7BhU5D05QvRCgZGZCK6bs3+
CCAEgIHqsjcEd9h78xEXJvZspHnY+Hq0TVLo+t4iuYGHmHtnm7WruE1MlXMEuwea
ZW0osqoNhuumhZlTBvD0+DPjim5i9MjNM+QfKWmogpfevacPdkfPPptUdWfkmNfO
VtEihueJv2cGTi3smzy/pA3KDwEQJDxUoV849+HIEqjmptZEHjvt/TlmB4eYXKZN
HR1Z2GV1C0PjNCTebBheoMC5Ig9Bma9UI5FG1y/OMWVWNMrDPQ2HiF23iGO51B2+
jgMrH+h5V7s3ZBeUptL4NaY9nSBsPOs9WmlYigK8iuR+KqY8m/Zcuk48QHRxhT6m
AGLFvB/aOqnaRhJixYjp1pEaQ7duEcibhNRjmGWxkSGcukqrPYTArOaqqbqGzH+c
g2HKTNCnHYuWNwhn+bUCxdXewRFSBQz2zEMkM+OzsHB08o6CmUkm16Vrl9kfircw
gdpBZKLD7bcu1VW9M2HVyrLnEjNBnd8KPUpwMjwKiRQi4r+X5KZPECzzZ5t3VzHp
7nzamPM4PPRWuVfj8rL7WDi1tGNqdntQQjBMcbrHpNRQsfmKQptadCuUBDtPTgya
7DiXr7h/3Mf0UWTyD9q0835ohk6FuEvabegunNZc8FPyw7sAnyr/HhwB8llK6TRc
A3DueV3OMPUxAorfNXh4MTtC+iHs4HZTIN8a8vnHweyl1FQwoTc7gmZdCm9UOJEq
oLwiwOvNUbQrV9iqCIwCRCw5WHr6rzmIvlA9e4O3aCPZwTReS8WkKkO7V7dok4De
GfuRi9nzxZ/hvaDZ9LDvy+EOJts2Y6vfyfTwRJr1SHlHZY99pDEEV7GPvCq43vL7
GbAWW5agsojaghzZzUqdXP145+Hs2vymids8z39lBmExbni9RwH+DK9ke7fw+cSw
BhFllMkmQge9Ku9LN/wjFpbmL7CvBU3UYYKwA4w/OxzadUCYU7U6nM91ASuxKnqO
dUg3CT36g7Ginowp/ynhorgWofe0o/AqztUrkVLvrMtu80ZfGbEBoxzi9Urs9HBw
POw+7agzO95y/XXsiSm6e5+/o0gA7DU6uqxTmMEfdY58HZplcV4QN4Pf+2xf5zUI
ohlZCHdRG/axFhr4HFp2kzMhpbkMOoIA5LdkqoMfCl20uhdt0oPGuiDNcksIqFwg
YJ10mowpIvICaehEOf1gbsiJb85OyES7QuIbKiq2C71MFfF8rRbF5KZjPe0XICgX
MeE2MQm1VgSvGrSLr5UBiP46n/pAikcAZBKqfqkFdS9wpLkKr+1+mBsT0xhibc0U
btpcjvk8DDIWoyV/CLTllZKRSa8mfp3r7JgylTQ/wYA3RHeI65xYI0Nd0QenygV/
aw6rn4dAPsUvv+GU3vYK5zRepAK95aIPSi7KLrlXdIAXoZ3B+wtsRhBgzn378Y3G
mT7BAF+Su0w4KolnYRr6j0y+maWvKJChsm/ACKBbAli6dn7WbLQVKXe7KQnZ1uQM
7tWYIvRnNPJ2o1k2Ec4bO/SF3pVHHFA734SzQgPss6rx4GfIzc731fH84IQTIayP
VotpPDR/s3WSKbZIgwl+t2BK4m+uJHUX0+YJPqfDXCiKcBdb2SyfWOcwOHi2FKPk
f8bbc8zKtLXMJt7ocFAQfU4McazJuQTq6vNUWxt7RcWaVdjyZCuYuGRQtWkR2P2q
PcvMt+54ZAiJS6171GB1p3iZIq5DUAETijOlz+9+ufiASJgIUcMlN48fp8ZSm1UT
2RKNcuBV6n/TCjajG/C6Aguy5bjHhA5ZSVz9w8v/PkPrLNwDYQKJcIeuKHt8tPBC
8PGOB9wNS2WVH5hb9N4a/6JTSv4V1Pn8yTVEOdUtlIabNiFmS5vX0yJkkfxsGczI
SqtatuHepH9iJSpDT8gU5UYqxhk8b6f/Uzh7kXdnIevSqK68bs9rHAT7HIf2f7X5
DvmaMZV55DdpDC91wa2B6ZqtIhaoNVSuF7V47qEzPzcpi7zKEvCwr5OxxTEBcQgB
Y2jka+KN6e0nIFrXdsYz9Hj5bY09lNKnERB5R9Md2fIBl8AL/S6s3IG8EDe/yH1n
TwlEC2SGOz7F259STq+sChOmYuTp0thZ0YC4jdVe+clHyWW2HkUx+fVQGA9b8ZbM
GjX+DuwgsK1nODrJTAdhbdw3wo6q22lHp20HMqlCedOw0XAtYJ4pJ9HK2wwT59Aw
0IvG7fRu7I2p+e+C5jUeZzyrKL3a+F3pf1Wuox2aohNzJbJ4zKP3yxhTIj76N0Mz
hdSU8tkLWMY3YmF5rINwIORkRfBl2/8Dm7VMgLAaTen92isowc8I6PGhc4dxJ3Ds
Gq6V3r0h8KVKNJQiYhc/B3wYITVRPFo28zQ4dNYsvSkcLhcUkTbd25A4PUU7ypxG
+6F+NKN9GDEXgiHB/oMOxZXMEWR2BLdh1AnBRvuEoG1ObyRfFzNSayZcoTOS/ApB
c9G8wxb81yxk8jSIdZvGIY7ISB9Vgqqd8Q9ixjLHOiq5GbrqfSLJsYXrutDKOTKB
q4nz+ZMnYWe2FwqSsfZF5a3sPatGGa//TvUgzvgwkOi5f2eimdgkpxGLi19Tu7hU
OiJW+ulkJMLLVxjZq1F4M4YVJP9RvXzwfxm2jNj/Or76vig/SaIfVfgZe4JxNPDF
mTIhaOs9YJ5dSQzaEpn9qcpKCure4YMOJwrlCrPzgyQbuUDFzPZTUrDnM8rAh/tI
0P+Pt3BnSUSwCLQITn9x6B1mpykvDIiod49rQ2mQe+aaEPirQepfZJ4AEATvMDM4
nIp1Jdnd8FvG+JYLv1xvE2y8h82cOu32v173PIttVag2SftpTJcCOzeonAOzF8uX
XWP6MJUPTyZBORhljdxziibm1mC01aj1O4YaDUr87Wx9BdC7Z9faKs+dMhUdNU5R
yNRtjkV4sXqDXKOepk5EtkyMtEAnDeX3f1ismGR2CSI5bl0fcEKanxwtBZzmIoAp
HQQvdyJM10PgxtE9qWpha56yatoIrRgvUMvgdLR73qpqIyqkvFBwttXWV6+Acf/x
y12L28zA+yU1VBlvR29rAII/h0elIbbOPBu1FkySe8su8tSpQfVtWACRlAkOCPjd
Bfvd5hgAMICuJgZC94B1UIxCqqkCm3D6wgHE++JsjHjLzHB0h9Y/f6mt1GLSqU7T
DfFE/zA9JFKf3AmMEWhINIkvxYZHA8me3bTFHXYENRMSNUbOpl//XiYxJ3QU1XCq
D18HXTekBKD8BP0qV6wP1CgXkHeo7Ie4ynhQo47nU35U/RlNaX4HVz0sNMXbJLIq
M5cW0aAlEMjAefVwX4hYk9tPEBlfrW0apczuZYfs6HS8CyWV9tm7aWncQaNfzmtl
2AxRzkJEBcm7+OKrq7vZ5CFakym99P/KNQ1J0FERydo2TQ9BQ7RBOzXz3QnV6I2K
xUyRA2iXcR0s8mWpKxglRxIcMcfw9EJohfEX516aIe+vX7eGH7pnjdQ7QxX1Yg/E
ZaOcCo/Sy2ol4ObIdBnqyV9jp1DBtWOegJnHwMf3lL/m8/GL4h/tSByPHjf667cE
7kz2R6x7/1ApxTefz/Pr9F0FzbxrxOGPRR/lmHUBWw+5wH0ttxgRAxFrOZ8nYs8C
z7O9ETFLiJqxVX9eNsrygQ2A63GDOs2ovxN6OZFaBt9+acabI7X+hh+KWbUGP5tC
jzAKUN5OxbmGtsUvp75c4e5BlT+JYlP/4kryzVERZCW+zcvrRWlGKFqjgckF4lPu
LQDK6w99IZk3lbNv7kmL0OIKGzf4sd48A1NP7Xejmuxb70WwWNsv9/Z6vYj41kI+
vRC5fKRMpNLA+bCQhYyepah8z0FkqrEendZ/YkPzjmKqc09834cBjfTWocNrsq5G
JsrO0u6yY/myTZfaiCBV6bq4hbIEBS3EmYHe6VhSGsZqRFGgRvO0977Y0rSv8M82
NCyiYN/fvlICfjwW78kWt/gKOC1wZL5yG7s+k2JBM4YWgy6AW47E4HUpt/9zhQl+
sIz8dtR2oJrY8ufjd95fVgB3Ya9A7P1GaGfTPnxm5YCSF0+izBzroKTzowax5zCI
lfGqSGr4qJeLku2S4e5g9wNcHqlrsm2ixmQSkGq5I7RwQeYBQ1uFohUHLSBOUo+T
+rY3hJooClIARC+cZyrdj6rkRv+1ZJp5+OWzrK21ajuJYAycIWoM8JS7rqjJT1qc
Yver1qEaUV4mhxTFZsKrcW4PN+fkzCQgN4f24we1WeebFxwfcjRui3opDeLX7EK/
AMZAQ3kLADYhgcnudRIJy7rY0R4OJqXd2aQFXt/JwwUGxpfReFRzqgarxWvyHvYS
36RFahPNiuZdbmTfvLfZS/FL2FilxWNE3AJspt66cutPNebR8T91hy7pqgwhKpxB
rTmSGgnFUquu8ePGaqVdyU7CnieocBlA2i9ryj4wWk1hzHnuWtNN1qh98Dwq5Suw
ut7GQDpTLHYYD+KdvooSuFJXNgV9tp9ajCI3bp536ibh06ZsNMirL7p1VAd+JTJV
KAFAYJLVRCgwJSXjd/hBjL6bq2QN7QJTkKET3cRGE440tkBJ4ZmVtUq11x8kLB+n
AslphX2GfbFUg6ED+byrLUYoCvUKSNFKw/TdbKizudHTxEURgbivedq5BpZgmV9T
NdDu6KSnhJHUgfjXObIaOW6+UIFjDQcxoIHBX/yzHsge/a7K1Yv5+Y7/P+kZ5UUl
eSg0p8DMQ7q40ZLbh/zzotjTjfxXJ/mgR1mmYZKEQaUDCE5FSB5qxBmMORHpJQ9v
TIsBHbvyNuMnmauoo29s9SVuBxQQXWeN7u5atqjO1Sd7Dg3Jz7p6ADm4reVTkUeG
PzOXLlEDERuJoxWQL5iT1mz0yMmzGm2qOg4sqRftS8lwcDbhlEaJ87/iY41r4meZ
S2A4U0+O+k1Ac+SzFZ8zZp/EpbIxTGNG5P35Mr2U3EajoIQA+QZm8hjLXGXlB5HK
oHAio7OHjLtBv86+WlJwrAzlg22qAdQM5WpkYqVBz0IqzyVPRs1g+sUscMRx32RT
n73sJGSvdRhepVr9zb5Gf0zhA146h5cM6wdyAtVfeTWNndPhPzSgmurID6O8vo8H
YlBPr+2F/7znyn+iaw82oAay/UIMxxmpedS/RNm04L5XLClGHmiqALgJRbkFOd/2
0tvQuyDVcC++xwGHETO2ZFyJc67IY0BACp1CG42gwBXYnfjjpJbpjtTJXO3tw5WV
ng7LgBuiK3EXGQA+Ct+XM/zMiEm44ZiqsjFKDcBliQaCxYaKLAhDVoThx7U39HeE
7CIbRH+zMLTdnA6NVUCIvdDjY+PJZ2qgy2NqDrUrmY/ntE/p7eFY2U1Tx86elIDY
pWBnmY76uCryGDmENX0yB5QrlzMZ4CQKGdylDaad1HS4T8ceTMtl4r9zDhXWKgWQ
8QW1Iq4X61kHEY7OsOvJhqbLO1gqDz7xwDKJ8F0KYsqcB9tCH4BjfMRPiMR/o4XU
0rfe01tArsfTNVVATvHlYpT/+tIKaYRJu9ZGOgwv5WVTBF9sMfckEUGTqUC8tAy/
ce/HUyOhMQAHU6vd8VjkXDVflPHm09xod2VzRYRxW/HljYc8odvbJGTTkzG+idf0
FksgMgLpG3fFHr2zw7OBw4hhnD8A6N42rPX5ngOBxGoN9PkYbsewvVs9h7+M5vae
cMkZNNhUYhGGg7khGiK0W4HlfedvV8DrDEvlZv2mjEF8lE+5NL/nKjOtCixNxT81
H39/WatOG+6pNrqZ0SrUo3AO5KZk+PucYHlZDx3IMBuQ6n1shxFBA3kQ8sqQbkMg
JToGp/w145rhF9diqxp9jYd0KsoUMwQKLjxTJqna9dknHdcGKvRN2wP9jlUtqgFQ
F7WfjG/MZdruCy0M921ZOmILCIF1ibTM7QPundvyFWr/TBpGUVfer8mGbdAeIh3+
PFMSQzaYb6gvzkkB0uvym2o05rrB2F7i7zx6bHRZHGRVaX12ddRGFouHMmz9tH6T
mblsycvXHmDBAKzZgKPqU3e/k1pCJh2PKUKrM5ZPnvDbl2R/LnS0l6gCxgE+hGPn
0wYEo3IckPs8BEI+E1YtUUiFFfk7OL+ZNo4clOiXDWDKb4DPbixxASU1kzqifLhv
5puHaYTZ9+eqSNkSTG08EB1lotHXAO8oTLlxDpEfPMX9NLBnduy7DJMze8b2NiCP
7ORP6PtZ0erj54wcAnhMBh7Onjcdwq9rNE8NXhQlqDjtMeYXQ5BcGy2D9ySsJ6Au
VewVe5SrCUdxO8cRUg76Kq4yuI0n1LhlqO9999puf9iPE6v6xGYiSd7wggE6ht2w
CwY5y0M/EqP0b6ifUvfDkKOeIao+u9z64r+3/AO7/cIwDlZaJHuhDmhEglMi4fVD
fKhkfBcfQ3PR6VgKOUoprfP5RXzNvAWY877y/Bvx78TsQHvh0weFcLFGBvXzok1A
Qt3ECzsD3GNK81mNP1hbI+3HT3PMypKOT/B8YJ6yyfI/9yXd9prIfxxKHRvVEqxJ
vFT05G8gX6xxOWpqdcVs0TYC4SoonhDDU4lwSbdLTtoDEttd/NDU7lcPfNhBwwwE
qX6VhUiBcD/OFsfER2MLvKDaUCtNh7QdqVOcnFrRnSRghrtmoF7peSp6ygo+7MYH
yApT0GZmEXcnBcRQZQBbz1/sDcULo2HlmxKMgO+cOS0ZkAal79KETPsYwT5V0gsQ
iVOTMYCWiY1OI6N9ohoqRkS4IUWhbBW0G3ogeO9u9N4q3gcfek1SeWeYTBgrfCma
O6ccQEsOwA4oZPCwvoEE5bQo7fgExr7vKgqCMdM0alJXmNiGDmLj3fmOe/MCvgZh
eYJ7plDjp59sqawBye8lhooa6AXQiRew69c9eg8o7Ip6xvuoun2K/0XHWiyVWviu
RVBGrlDVCPuLGXW2ZwarB6GJzNXzw/GdFLWWr68oOzMQUOpbXtXXa8HPhw/c4ykw
Ypoaok+HW3kcxc9Qj/5Onsi19uxWhjUrhaWyAhXs6l2lp0lo9YCKfzZGNQNsctFT
TSIntYQxLOtYF1wTcW0HzjCASGhYjx3ihIgjWZkeiqjHowW3Dtel0Wy5bxME9vOo
IFZKuGsQq+4PHjktHzWFkaM6Y92ygD4nF1GtbJu71wEecq/UiJAQajwGZvi8IHO0
XnEgYas56bA/Y8Iy9gxpT/vD+hqlVrWNDyD7mqEsNUgaMMMV4eUVtyWov+DkHfe+
fLuMPK7Ydpgy5Tt3mJMDJesWt/s4On0iPwGycVjVLhXIBWctE+EecD7SC+LWmlz4
Rm0rB4G3aOGIENH/T5S29gR/z/CrrXQqnlHMq/S/3Sk7fEXaxXb1J6VZPpFcxmqn
ZV74HXB4IhabU61CDolLp/OnYcJBlO2vpO10djcFB6j7jIfyUe9QKGdHbiEgoNEz
ef9Ofl1GgjkgzV1PYq+XjpIUdg+PNjH0et7XMtQKvzr+7CTFxsbdGspRzWxsPrxJ
e0aHjLKquQ0l32xLuMupdW7OS/9kGUyP4Y8OqHB50qh3hLMZezy3S3jo90TAWsTH
O+SQgkpzeb+1o3iD7f+7DDeaLLGWX3RsXVhT84GgQaMeJCOFPi1dCflWPJx81SHf
zKHQP9i6kQqqQAtrnaLMMUD/5laD8uI7gULyEcT4eekXEmhfjY851ASzFAnHQY9V
HeE7dk37yek4BPmIzuDdRG9i8gwDhf+5U1TkkE3tgK6aNB8w3jJbLAGIH8VbyYjR
hOlBM10mJBcnfXmUkqcyNlCsLtZGwzr2xUg5c8UwZ7fgCfHyNQd+S0fSa+VRKqbz
3pG8MsoO+bgfTDkl2iM7L3hTlCSFgaCRkWRGhG9ZkoDriPs7c8csdJDyKOpmCVp4
YwQZF8IVjjTGsfQGIOsWQ6UfGD37Af5PFiW61liLKdbGu0+0APcyLhj+Y9SRcNXy
L5smWAsH+QmpxWiEzz6MGu5R81v+L4DxXv7YBIxsnAfo6QZY1JCo89cOlC4kSTmk
o7uMpk4629/5k4Tf36jglUnD+IlGIDy1Cu7Ah2TQoBTlHsfsO94ChvnF2A4VQnvn
CSb4ZYl0a3I7a9AbrJHjUZkhgtGr59Td9vimYpMn9F5ENCuew4oB6/ahNpV5JMeW
KPBjZ4kQrAgFzlVVLAhTSagrrXaaoA1lF4ZgIzufj/LgPd61LzJvYPrjIWHvHeJy
cDgJRqlLkiq9auubbbRSP9sTTKaH8YrHLBk0RRj4EY2Iw08AWG66bqAZbTA3SXuK
eRy99gwwrETQShgi57f0YRgbH7UdlAIuvL7VU7hJkBQ0/wWZ3nBh4uz/5xcjmiXi
P+pN9XXiiFKnJUqPgklfsDRpespxdE9KsI8QD5Rz2JrtF+QmywKoQAwa1/ACMpMx
dLnha+UIBE5xK6LJ/yTKAl7+NtB2ZTVBoxKUYtV+sNarphTPnsVxINbLc6Rw/BKn
F243QL2ZVwBcYbWAIAEkBTdCU7P9ZNNu6U8Np+lmwyU7guMwC5+4a7I/Lz1tQqSO
hrXssKvmwbh+AboeLb1itgKp6V7mMetWoC7JHZ4tJD3FrFVUtKrWZ0YUEBJRKjor
bMvqj1P1m1K4aI31ZbQvPpsDpmCrk8qx2QLcpofrIRhGw8wwfixKdFmrWt283f13
tI2CfxAH6+ZSivnxoCxoFVAC2Xmdm7Mo7FWxv5HU4whOqG8EprhZoqFz9k90dznd
RqKwr1crTYCap6roLMzTV+Hhd5GOjyWBeHcCG5LVPvsZIpRmTpvg3Wfs3AEwlFSe
5ptHiGDtpOht1Rkxv44QqQWL6kK3bF3LQPeJ5HLkIyrE8TNLs0Qfyym5X/aXOAZP
0VTv6aRxZa6nejwhDufqCaV3Je8QgV35h5DLdUATOEDnkUDDICLINJJ3CdMvuHyg
TzvHssHwojIfCowfJsAFHnBSC9VgRPZgays4AfzU8wi0/JBSl8TAn1sF3wkP4UsV
k/rZ1QNLSfyg1QW6ozbb7sM7T+HgVvPhwEKlsnPQvBGW7bbJo7CrSlv19sHmIUYq
UVjbbC1mycqqaYAz3lWYxGUotd64NNbmJVTB9o8mtpz+FMtYAkqV0k0dUPUuC/QX
1q/vCgoO6I6QSC+KHzKOLQUw6IjorGvzaH0jz0IirYl+dK7PtIx14aIK2LWrHAGe
4iHINukXOUI+qla73fxEXK9trMozr5IB9g4R2dHsDzG0PRWXoyPQLnqeEQUbefad
m2w62ZDy6KPxDQOD4T4VAJjrjhuIoSBFWEE3rzem3tV7mc+Ntd5UimDhv4QhZjxq
GbpjIiaaO5wD3AFqXGWdcKmEu1Q3rPc6MSZvwwcBGWy0csG7J4PytFO8V5Lg6khx
75BNpxLqCRR1rkjau4xOb3WORHBng6xjd9cZmxJ5BcQTb7k2POaMQuMgxHPmzw5U
uOof8JprVMUo5I/SFn7RNShGrwY6Xeqm2p1tdY6zDCDFEqlu9uR8U6ZxvU8pTMhV
5tUbBEIr0Bi/B5EommVG/PBP9QMMoweVjkD5+d5O0viR2T8xQryLU2Cua+baEibe
uoCpCapdGvPnZxJe7xGPviqEpfOtZAQL2s3gZHbPqt9+mgNz5IjjU54JCBgOF5Ux
O3111qD7fq9Zcui+3Q3B42mZWQ4uYH8ORjzIZ7zHNyQfZtqcHP8APajsoA9DcPO6
PP4uci6EAHhX7Diw61usFpjjnm8EZASVXs4/Z84UU5kT7D9qVmNeeNIQWpo400Mb
eSAJ622whEK+3Gtn/nhReqq3OW3Dgv21ws+xKKAcdAJSjjjpg5Ubl2tv7XN5yAbR
9atr47IeJXRYTPhj6C2DybErZ/97l635LcEfc655TdUEEnJKqmDdTIV4175z3wSp
IKMlvwx58ivS4Bfksdyj+sgobASw89UBFW3nBnyRWfUXma/toS4sk40SXhX210qw
Tys9oayOYvCaApTnnlKu/tVImnHpGhzCr3inQ0wrolf9DdSzSyUnAWMm6YiJCBA8
n79JmDwoeLtBPh4aDdEWMjJJz/cmIjzEso+XFx2avOLzxP3Pa66/looKyLmhqKTL
k5TkTEsXfOEmRuehKfVw9r1cXHbbOIlJQprNZPTv9tEHK9C1P14XGC0VkS11Lx4I
IIr6qGVv7sYxZF0QmVIPrFbeOzFLX61Soe2TzmUKQA9EE/7KCyG6uCqas52MbamU
ivR4A5EIL+hiRewK4WR9hOdoFtgq03L0BAkFUPuBQTtZ8/kEG89jx0X1a4uaBVU6
LO0WpoKc4Qxvh/KoLr6iQDvkDoT7q6dsvAE04usoFWDtiz7aXc2DlixOpYBDN5Uf
Jzn2ZDABBP82cpvPXuB13vNMRBqzG5RaW+e4LqywPVL5U1Om5ygy7Oxc7E70K8/h
jTIN0DaH6KIg4mZt52KXA/z8mT7TPNfG4RxsT3DK6ccEUQ1wtJb9gUSB2S4ChyK4
nUcpmbbCbHbU08myBjSa627Zz5Z/s+W7vIUbIOOuI9VaGVVvL9s2gJ5u/CMtGc1J
HISxj23HWmqNWtGDbJmoQacFh3YBskek8Gj8a/AsaBFiEJdGlajU0/wyhHaX+WOc
F6d8w0vLQTGJGlt3PMcvhnpacdOLNyTGiB+8/M/pXhuENumlyreRW3OufU8Gc+bt
vmoOZK7ynsEZ7gKvNSz+8SStZDfJeUuFM5dR2eiJUDemKUgAts6xQ0epHZYwSgCe
5Qt13xFvxb1ziKytKtFdqHPz/ZwZ0BxdCKdL64Tfw8JKmm/EODKwj4Csgd65yW6M
B7C871SfMU80C27/71xAD7joY6QTgVFAFBm+fguH/2lKEwEkQN/K28/dTJfjfXcI
u25yukRPNa7YuaJZjOI7MJWP9HT37HJbYZ6TH1A8oIy5ABHTP68JBl7MAyy7WJ+X
pmFEXLYTqj4d4iVdbJCM1uRn1wcGmDDVhhzIjtsPxjBa7N79IRyn/yZsqoqmLh8s
FASBMk1rrw8jFcNYfKqLrNaFICezi6oOaDGrNrtKISO5QJcoGezLbbRwgYMi3SVJ
EoygzyduSAJc+ZSN+zSsznkSuEtzmCXyJSfI3CQ55TGqJQNsjxDsedat72ex3zzZ
RGvk3n13G/w1tWnLQyE/3l/mplzCXcQM+MDtWO2yfaC/s561rS4mFV6uPzNZhNHZ
MopUXiKlY3kVs1C4xuGe6+X9Dcb7+5tVpcAXuRGMO/uUPR/ShWvwiX2vTMyWden2
oOQoXJgYm+l6y8UL0eeG9J+zV9SeOxtaAfxIoJ2lNxDn86cVFPHaU87G51K5efXI
BsMY5clB1AWTDkMKWoZhzFVWHmXKCaRvURBauV2uzYx4dm6yUzHwWwlaGLkcj229
MTUOLZVQhoubiHjRPxvqnpU42OMW38awjv2FeZtTJN2j+FKujssIVM9+xH/nzCYv
vFmzqB0YpGyd5Gw1rJu3P1g+cvPofoytQa2kaKRyvfPhhYQeyQ3inf9mioFFAJqx
U5AxdvgA5PbVOWnet4LYI93bfwmQ0LoYPErDxye/ryWEYeONaBNB3XsAd8qk34ku
9L/er7VqBwHgTkWd9KSvdVz4Uo8idyY+eFlsQMdM6jWJ9gy0EuUMIZu7ZFf0+FGY
pbsl1g90bws9j0f9huWdEK1+PHQEjeeV+f5fqwtaa+wDSmnNkVhlNyrPlm4Vk9s6
ym67DtitAmP0DB1dfMxqUk5eYYai8jF+kEhlwSGt1g20i4rhlKPa7P7zphR7CvqN
WOE5tOBDlW/Eue/qgCljhj8e1Y6jPuOLuq958K0NdGEF4XvDMuj4IRuqRM7P1EZR
AVgswqRB3v8rKriTFcgvdyPoB0oUP5EzgPWl98aVuoMnCi1c2/p5apnM83YHfEYc
WU+6iVP0eV2PFBuNeoorAoSNh85zP4Uvp9O3Gve1RLajjD5xSEf4ay79d7AJI5w5
Hqv9rl/A7sgNkn2ybet0ictRngpakRVbJoCg+rz+NJA5i8jk6tRqneEN9HBuYFeN
+P6PJ5kvZYq0IEgcwmtXyUM7vYk+L0UHPQ40AiSbXqu0r6cyUZOr/b4GouDkwbOp
XWwOX8+Eyo4c7agg4yvW2DeNfvhMCfXtJ5BkK3WnhXhXDFmBiwGL2yGY8gFjxqLb
EAFZ9syfsVWNpK3i5bg1YtQtXQJistlicXh1h5YEiEhoYoTjfZkzFFysQUYv6sVo
uF5xgt/xXqLwMCJkQmmujE9n9mI58H3MBm/LvIQIZgH27U2ZMcYd4pJnALV0CSix
XfnEVGI6GPvt+5Nicoiz8XGy/Z95RHJZanlTO6k0ToUesC+uFk1OW3yzZu19CVVA
z9VxXLxwXZ4PwHoXWtlsow/wFFba8KFI4T2fcsY+Vp0zgX7XeugYTU3rRzdH9djo
00uRxqlaP3gR+mKkpEnsjRSt1kl1TN4XrYSD7nRQnPEdzBgzeFdu6cEq2J6XWt4S
X1+60WMDsNYTPsQsvosRin0eA0MDzZWZYME/LKOp64PKxUZXs4Ay3otARmXiKvvR
YSgVTBrwKBYhJuEILYqB01uYfCIyCBgzRzdnI22i6gbVOhsM0fbGwMItKCUrecnU
wVPU3f2hZ1vvKPBZjABnnQsw9Zi0mRwYSEykI7wWgYKgd/mVWKPEPgDXRGDQD+BE
ivFlLdAPoHprsfFJwW8C0LAcdqFHZcpQxqkJ612jRDSPz11BIpX5pHlw9/pwpSm+
opV6XKi2n4dM/CgznQK5ObBXwiMDeIbd0cNQkz1ydlaD6/1wkXUHghHnLIyyFzxF
AhzBDad7tHy0KBbEMjLzYtz6hNDT9H17k9IWdOzZUoaoOtLLF9cXUcun+ZwZeXeE
8SoviWGDHsy4/vc9s04LP0XXv2yApCMRWi2etV59i9Lu4u49Ygin0KFrbsht8TEp
QPxrUYQftAjOSM49MbTm5jDhoGeKLa+f80qhn+Qy3V05GXPDGyjeAbaM1+e85NJh
FxJq+bt2K+ThC6sVI2Ww7Sdqvpl30e/BnrqOtEqe8GLcoHsUtrC6ICpKQU764r07
TpZ7dDPyFOium+tFXg0tpOTcTquebjJOpjoNMaNYR/u1gXqkM7kG9FCqQjxTvJJD
0ndkFuls0LXl+2s0JLHeWZmtSJ2SabMwirvEpZJ9cZTbG1QGzgPZZ/DxUFBVCD0p
k2mTA8ybWsuXZfGx3pDAnnbeaNsia93GY0nVZ/LJvpMl/brJLVBUQEqXxEhsArEt
8GVouCdve91M8KrmSduBb6YytSNt5EBioWBE1GvESpGhknNpU3IqaZBxfKPlGw0z
DXVc8cwYQLGb8EBBMwtiWOqIjpH491ZBibpmTkDdAaERNMZR1Ejckx3pIckmCnce
kOxqQxyzoQF4WeEd/nn2FsbfohOjqXGckoBQmzfd68lWvjEXDz8Q5TYXJ8kpg899
rsWJZieAxyxSzIGPAw0Pn6eoznYAAiMRRR8fKSGSojc5i2FAOlqdOOn8N4PApvtX
2U7foKrRAed2Whr/Jc9vxCnIIs/SajfOV+nKeBoFtu2H/QYdq2HBacVzQ/Q7ZKu4
BixknZY0gT5d6zfTFFvXHRRuSN/0cJT+NdIZhjuNvcA4KH87XRo/LMmKMeDrSNye
WgDrljv6R76c3VXUOnePLCUa66SDwNvLLRgR2e5frKtxYCAsxt4nVzYJoQs8pGgH
ZJty6+9QGuPNq1nIw1HmAFjamxEg9QDu3nk/Tk3ZKbpfX15gEir3s9q1oLZcH56O
yeTxkZaDcXd95mOuoaD2bXPe/OphNdAtTUjaWU3DqgptswqcvjtLhjPCCr4E0VC3
ZSzS9OeYCrL8f94krHWq6Fdf6YIZDFyalKf4hkG7+kXDQ6JGJTYKN2psR2fJlmSz
/apL8n7S4oxlfTcwQQKugu5AHOZ3aLQQEyg3SHZYfyE+RPboLMnLvjMEjuq2CuIk
V6wQJ089xoOECK+Lr9Qgfq6ey2ywf2WbBzQKiq6dY4/NhZkhcDahqIHGGdyxRjxe
dC4e2SgHjxFobJ9NGKUMXXHtAYo/Rk8L1yhNuIpThsa2BQkIBuQmWhFLiaZxnN1i
AprMOk+dD8/CvMPmHQiSpCmDEIaTvd/YUJh7R/b3vjIOAXPNN7vfzHoewm4Q/WSR
GXnCxKNuF+UIHR+VkRhcuxoQTXl6lnGxiR69Ldprt3hqHi8TrtvZws4n6TQoarG6
D4Wkncbm9sMcTyl5D/Tj/HaXJxDVGFDHTAWkO2J3575MoYif8lKnIiht1x3sQcrJ
HkWHtG7YjqcvX+RZrk80AIuRbVzjK+gZf8E0cX0jVy05gbcjvNcYeRNNGIs2tv8V
gR9tv6Qj7oA1LyAGoOidqQ0bv3gsoLs9SVl9v8Ro+p04kHGUuCHW/nBmMPKUqGof
AwnZZCLA7T9nnQr/SD9mFrNh5LtkOwPoj8pI2q332R0by0KGRMRF7NWvXbOeCv/4
JqrgrqEoNVy2MQLkXtDo00udVRFZd7pLNIr0f2bCSMs5qOjItC4/D644ikS61Zuj
spivG4j3DYeWdwLqdF8DdtH/lgi2iI3VaBgHMbiSJN6SjSLQj2M0toAEb/m/F4Do
vv0+Lb+8Deod71kuT+8FcQloYlCYcHbs/ceiqr+sb0HqCaSdFkf6qs4I50C+dezK
vg3ERZncu/RnNgnSqBPaRME4LoUy3Z6mNfVAh8ObTRDiNl1/XMDoM9EenEzXptoM
hiqF0Xgy9ZJUDwn47eenii5S+UfIIzTRNpQ/0EjcCD3lMU80aIh6WbSRnt9NFqt3
aoKn05Rusgz9DR0PBIa77puFA90MB4UIghesCjsU53DVNqCKp+lo0gdWnf47z3y+
ky3qWwbftQH2P3MSlVUzfkKBFV7734Zayh4P1O00GDbGk1TEj6mYFgxmRCZ1ccIp
3EtTPbRu3imtUBgaRFsV5VE8j/J0y5YegBMHlmjemqq+C5spDzi1XnEM4QHiqRjF
3Ackn51rbkLcv4A2L+izO8jC7mAZiIaKBz3e4JvVUqLB0qGJazLxffntr3vhpeTj
LaZnolO7K5xKQQGGQlXTk0stibm9P8nIUEXb1IdjwkirrjlXI3WsGZmj9LiNsA+b
5p5ElqAd7Ui1mdfi1KCNfjzqy5t+/SBeUVvRpFsznsiHBX1DoPCeAzUxKO5psctv
Xj8kWSVBAgVOyyWXeT9xC+QUcMKKaKUteyDoUTm0l/YYe1I10O8sD01ozc/vnN0G
1LM8w+E+34ilUVZtuTS+CexUjINH3aCRXvCtG6pHG/sWomGZUbfsFetWPbqShiDH
ucCt58KYD/aLeBDQSHfDW0lthei2zzcqvuO9OiamFP/1EBcAV6o2oordzcpK6gDs
xwSkzvgETpq3UZgcD8NfI17Ds7QUknD8ei14bkKW/jT4xQWNYfW5W2enLxzYY8an
YCmMG0oxmi/iEMRi9a2rKEHCqlH6RuKLhE3XeMP4dPGqq/38FAwP5pZmqlTQYThW
RZ+H7UPS8BL0KhfO/ACpVNmAe/u0s+vWrOe8/EUPe9bMFjrjSiBTcAHApdIT/Fjr
IQtZpCb4TpzSxz3v0KbzyMZ5Y4stIOD3wm2Skr7DMLWU5GVNAXrTvcmh4ffKCskB
`protect END_PROTECTED
