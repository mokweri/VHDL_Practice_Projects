`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vpm6Tkbsa/aiI+fIJENhbkBDQVFvJTU7kqCmTtUj9fUrRl2bcDbhpNU41oLWsD3M
aqsJDF9nHxUQkpAKRA99bWg+gKKvrOTKk3Wg8JhpBKpUxaHgdZ/C77o1Cwu7wKiG
4DrBP0qKzCF2be84NzGAnjAdM+DYdNeH1We245Br4mUzPkjxJVStEXVdrawqpJeC
BobrPpSrsIsHcjzNrW6pyaVFxbGYScLXORyekLI7wDAHFGSGvM5lE89tyqUZntVt
06GjINPEahb3wQuTNIguBwAiM9p2fZ4MSUUHRvB2I2cFLP/gwN3Ty92a8kwfDax9
cMHyC9JbhCJLUxfkLG+5uAHnfz1Au6KgQBaDzJRfIUsE1/vV3Y57mbriuK9FH5uG
OlxFBp/48sV0ZW5BsEOHCkjFbwm4kavs8OnkY6XAnt3VRs6Qp+T445FkCSI4RBLM
rkHds8OnRQSlUF814LFzoMYzGdQIkgYtixwP+2pqkSnenkaO/lij3aECaDwucw1k
QKXywvpcOZYfl2V1pwk1accNlgEGbUSLtwEXEWlKtnoELeUrUQPDXaiWEKN+E/4L
NFwFvAXVfvS8jPY8r9XxzJvl7B3v69xcWJXvWaJ2w/JSiAo77/UWyyuTbGcPHyZ5
NicCifEHVzANBNfmrDBquKOQnMSOuJ5eLVDJG5Pvi+LQOIuVf3ldVp2+bYpXA2sX
+sv3R5B/HRqsUZyojF9Bjlg8YfjTXUP0VtSBQUlQE4sabW3MUQPborzF76e+tH0U
4CCq5KbvRHcRrqpSCvKM8A==
`protect END_PROTECTED
