`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y8hjTiHXZXq9lQrSKkr36Tbv4JouKf09M2V0fZ06MKtNzUbXbrdw6+XGQ0jn8MO9
HjfI8bYEXgcAZX1sz66NTHcWRnChephtg+y9iKKk+0Cc552Y/tEneMkKvTkLRQSm
XZKKhaQHvkw4K5mvF8Xav1QSkg22ffmHw7FFvPAAiWG1q7vHMQFJy4KQT68a76xc
F1X8g5DmZD56ccwJoFMcQRTF75sJRqcaM+h9ayfZWXB72R5x5it/HH+yTJ66vqxA
Zo12T3BGCNqCeaJKU+vUyQjMtqD7yCWLPPObF2uVczch7+s4YB77xTSdTSueAXP1
OaC1rukVHjI4FzU3dLw7K/KoTEcC3/bsu/LWZmQ7qEPilL1MLL4XRuWwr6QqIv9u
C1K4aHYqcuAVtZcdgDlQzONsTrp/HfHsxrXlu0wx5/IGZotTTVqXB4FJX6GbvLT6
4pIiiUFvJu0bb+mR3ZjbGnCXa/UjRj5SHdNrUQDu0fz2rIhASRkkjojmH91wpKRr
YI73c3c/CKreOf29UFvemX1sDZPQdpewXoJvRk+gr4hQtJ7I1wfW+zuiKXuMOw9J
tl9Q+DVqJLHBzZaaZWUEbcGvjPx9zyNfi21OQwniMPyjjMX8A9uHYWUoFANB3VKJ
PcV3wh8UnrQ349uT5jlyd21N/p7evN0QH4o/Tl3j+xcN14dj+MOqL7Y3bqGRINBd
2YxfGf7h1Qzt9zBXVq18UgXS3w4iFWMzUz0XM78wWqlfYXEHxGVF7j5uZbBzlRyv
7EpW15HbYuS+S3FgPh3M0Afy3u+a4JH7Q2Ose7RMuMTBVGl1FDRIVs5fBo6Pq90y
UFYnGL64qUoxXOEx9YG+wkt5WCAwYEJ6hwvw9cgdiQjA5eCfKkUTna3FWoOCmiPm
StgouGg7u2monPR8dVX16s09oZ8oFj3rEKNrLn2F6Hb9QOaWHGKxRjYMETaUJgAe
s1vX20oFeog7SzsdKPSRSc/G3JfKQTAw0JKR7wpvcAgdZEjgHOdNj8OxeExp/VLb
u4Z4lYSvFPcoKSlspjUNv+LKLeQui3qJjmSnYQkId67q9ywbPWgn4Q0wGwzZ3xGL
OdK5neKaUXc/BHxFvmv3Hv3ce7OYJr70lvhjvR8/x+xRlK6tW4kJ9W3qSdh/sHkO
wDw2AnZMnWyQQ5S4lRP5g00ya/4l4c/sN/tleI/+gWrPmkfva3+ITU/xBmbjJ8Gk
UXHUzd0kyQDxWZfQxua3FcA4eSKgtir/fKEJXl94NuDBnkaOEyXfWIYr9mnWXeJ8
sndXYFRti3GTq2ICbwexWQ0ZiVjdJ3ulbgMtve1n36Wrkjz6qT4Bi+XL2y20f8XV
IcyXBqCKL/JdXIDFEH4iop2tgfQVHqG0lFb2dFqFl1Qa/xjSArhmoYtcX9Im9nP5
kLjE344MZ+JBoO/oF6FC6STKDL2dQJFvus3iTKQRnKoaEbTaevhgSf+zaD9kvid1
D1p/1/83jsP/LtvQ/oN8y6uGBdaZwaETQivGzzLKZ/zNnx10bWbZ2/TicdJ33/+S
w4YD1noylik3tUDsV8sByqk5mw8mbCpKoAiptsNvbnAxZfc7u0btTplDdJjhOQYz
pPlVd5fsDZcl8FnX899KF/vXgvnEDXHwp51KkgKFOOXg9inlRDv3rDs27E41yAFw
5doInHvfnZB2rwyopLi514IIZf5HF1ZcWlVOc/n8dXfyYOERx98nhW7A3WmQjWqz
sGnvsEKcWOxcr/Kz40XfXkUtkp7JlAbK71hFEAV7Ushv8bwMoc6a5QsBHHOr6+8R
kGjEvBSr+RH/8yqb2Q+7HoL3c1VeFqAH53a6H6qhUuXKUusRtkZmolj/QGDFWggq
4Lc8MXfO9C3UvqVFFyUH1v8DtV+r6xvMN9TaG83AVy3jDjXsfL495vWrRG3g6JB9
ux1XbkOz6+d60EMOE/4Ol0/kHw94wd3aWuLBwB2xqnhE5uOCweBr4bKDcg5RzjHg
UrygT/MmZCksnnPAIeZfxbqDTwBIeOJvrHbJA/M4fc0lJwUmBE+MM6SZcSvLatfN
3LUc31hx9AIYfBXhOExKEB2Uwp6O1BvuQxgirY3WhXtMq7g7p7dDXHwHiqOIicu4
jmTUQP7gS+PWnCUGpRyPv7wLUmnejk2PmXPR06vtpPmDuMcouqunvahTiZvbwTkJ
kofAmqXvcESJ2rYW9QeRdQDNMpS/ajN49Fcm4xeAHJmif3qobSz+pgoYOKWpFPYS
/tcm5xCkA/CFo6CS7KXffVh9SgFI9pyisEqpCdSlQiO2uSY4DN8YYXvi9+HuDzxW
40kzPBGokVtMkaiIgbw0Ar8oEiorlJBy8W2JtqZ+3EZR6yqSbDOKU8imp40Tqguz
oCjiria0InvBGZhnGPV5Pu9Dxwvmjjd5TwJzd79fWO5cAfhM8i/sCdwldKz6jXOZ
yoy5fLIRQD+a/WAK1ujhIiZ4n3LDGCNkq1YtczfJMFtO71/oR5gM5JZLGEiofwN7
JR7oF1v9q9lbK2HHzKCi1cR5DijXXWOeWQj3VW2h2sWkrBA125CAqY+KlFKx3xkX
tQv0dPIrRwciPxhr2bq/0jsY2/GLX2FZexBnzEADkpU08vXHaSRkbfOCWQRczxVm
OqF+D/7p/+x0WyftW80eGR4W2GIRAbhed1/gNzSUPh5KD6HG6oPs1Tr+fjFPP6Lp
oQxvPqa6EIpbKbk2uaLQTHOuUIbrfaSwdMySZmQWghQIAIx+I/TgjIW3dULKDny8
XDVs2677se0iPjo6Ayihgip68wnACoOo6/nS0jNJPgmf0BW/7GDVqPAmW55kW0KT
tW1sbjbZpvVNo+Tltm1rB72vRkr6mmxvJMAHStrtuF8RaCkIcLghxrNOyyKutSID
tDQZsOmjkyvwe8DeqX5a7BEQLgFObbvNoIYbGjsX5lZ9ZPHtIgrxhAkYfTXqbh0z
aMsqEYgJosLYS677A6lObENNGm0QGUgiUrq5p3vFDRS+UcB36MR20PvzCb5fnlsA
5vbg5eF0wnhKUyLCzY4jvFcGuRD/QMCcx2Hc0B/Fmb54m5Hs/u8YrCqWcL1Xogeh
BTETFKdqLaDp1g2vRBPrUrr1sYVLKRYtVE7RRhh9M1Db/99A8v+niynA8KoynK2f
+FSuTjEmYlL+w9T5rW0qJBv11GaagyXlb/jntolF6IoLFwTaCNnwmszbcuEXcJ7k
WFaDkgVPdA8wlXZoLDTVmI+BsjEjCU1uUZLQIWCr1ZmWYJcs7P2MGP+3UVUx/tPw
PshLQnBKBwawtC1BMU2775BjN3vq03GuDvTvbffvSnX2lZB5suh5pk3ZaEQ7Eu7x
1ffQ9rKpUGnmUi/giE9FmrFyczCyPJdII1SkLyomTsDSEL3GHZZ7/80WFTOhjHbq
QQ1BNpEU5sxnklWKpWs3le6lL22bl52/xva8T2A2KhW/mVPC6pQwUJ44RTW+w0KJ
iQh3nIDu1D3RQT7mq/5duF63iuA7MgsXvlWT5PloAGlLC1a+mGD013jwbBP1vB2B
Ro1Mw3dhUCQbKpF8ayCdmZDMoRYF/3YNryXTOA6P5MVQ79sW7/RX9noVRwhG5JZP
nfpZB6CahUjEjvac+pa3Lz/24EjjEud0VB5sg7Kwlk9Zlta3Zvb8e0vLiQSJMhlV
6wFNmCvwzG6FYfxIcy9Hly95FHVeYYYZPgjRMLu5lT0AYjOzd+5oV561PQDuDHj0
YzX4dl1bD49+FhqrHwxbVUS15rDpD9hjDbN0EBE2bQTWckcTTwWlAWDdJwnw31KX
yseBztu+ZQD8XX/KovnBR8/Bahdll8o2g2A2QQkR6uRSA1ykm2vYMuMxakD8AfUk
i3H1q/STL2ZO34fgzsIfhntZRafBYkS+G6Kc5kRusvNvlEvbEBzrIziscPKUyXPz
RqGNPd+AXwr9IBTMsgG63uAXxMP1mkX2rrbZzuINL7sRt0IM3xDSkOpkC9kJ43D7
mMZOJ8b7A04xtdR5mAOpcWIMRjEJNfbk1g1twWrkW1m6kRRNYs7aa+JCdD31iPIi
MnxAgY1aUomI9DwwS3T0dO8oa4PrE7deGax8ouDwjfXBZbPgvb0JkfAc2SFnueBd
WuM74TF2gicF9xWSjk/9nJHcWiIN6A1NSL8jpAluOiFblzzXuS9DkbIKzfgRwpsJ
3W945hfLV9R5E9uD3Gs2V4NeOwrhYJbabrL/To1UOfntLe/XN8B7abSc4lLWw0Og
8tvDZ6fz0k+ab17PJwk4hstKW/ktNyiimcc6IdOYmApPYeFqn8BAxIoFiLWK+dtC
tpijZmBWKGggcsOIaFhTEhHt8oWemfw7cBuyE+pAmOQ5PFdGduJNVXg3GhWka9Zw
pwo2q2kqgwtwf3qw/s4f/AMoEIy5uQmjSkOjhVIZ8k/vsxNWQeDkZO1hSoSrKG/B
UcoqpJKs2dXwEhT9lyO2lfHtqR/BuG+XIHqKfv++OVRlrITqHRZhL0qo67Tp7znu
rsKWJH+tXWnmh30FfJuCVT6RYYGhZMx7OE3ofVvPvFOTFDZZef982eIwnxKQURCw
KBEX7rHWvY3S3e+k3w0P/8PQZez66OBrOPME6bnfBqYMnDDoojdy4aB4rbWiIZuM
xiVJSa2FUPkqUb3uQt02eNs87cdcPE1gcgzxHnSRF4Shg5M1skH3udtwqhVfiZuH
UDIqBmaG05dxRkMMxd3d2iCzi/Or7DcBTu+b43wZkkIeezNw+TcXuVQNZ3BiMD30
wgxA0+R8gKSHwfDF0yOXOektdbaU/Vq/LYc5xjD824ZIuO/IU0CDzj2CT7hMhxHj
oO3WSj6j+6L0iuDFEHasRigeEsfm/d5L3WPeM3RrqYPIM8e4zTZhwp9DOzJF0Fy3
lPSae8DWGT0ZI+ptJKp1I3eGkTxdKSRdsyvwz7Gv2GdFQ1KQ0pFXSwfbcqtQtf+3
ItjXHzXIb+Jag3PLP4FduoiPBNjmEYnTXNd0MAnPY5CqBt/8qH6JYziupORcNAik
yg8InkNAbIg4mcQuuR/hlFHHdECZMI95UWE1uM2svMkeLlYOmnXVFPwVrab2Vh3z
c5uqzc8mQOqUnfsPobz7qSP7fhpCfDQlQyxbBoImQBRaj8Yi7HiOkLzra328hhEv
0jZ744f5Pr8+t5vHaS6Lcq6U3m2gG0pWIvnnsYWO2cwvGetshSXvxxJH6/DRGgyZ
KcKfio9l73PVAHI1nhfsSuVO9T9xT3ud4k6Aa9b7Xb7LvJrWSDiSIzA1P9Iaz4DS
c0O1q5jg4+vCnu+TG9ovGlllTZO3Zdsl3XdfVbtgnwIcau+U1PerJi4n/zE1/2sm
0gAKZB7rVp6Yb2CJYTeXIc8BqC81Oy/J4yB016kJhrgCTctVvZMLzqRW/62Thp/L
QqA7oN/nHGlKvHKckl7D378jOW3jLmQM/JyQ7orpKJ/AWFly16z9STsBcLLgTWzM
pQ3fTufa8qompgQwkvLLnnMMcTnvC5zbHd62FcVWOAxoYzDk3IhDYVcM9h5oPVq+
MYAu65XCN+agoFIsEaiHfjUMKhZYA/GPQ0UDLGATjjLkhbv4rQ5sJVinHgQKgSiJ
jL9qkRqLCEOMM0ZyaG5EsG0AXSIc76KVM0Qzo7PnFwTCfdjCkVi98Tlias9SEZxb
4MCMsnMdL2IibEN2109ZkHsO3AfiO4PbbPpJG4w5AJ/eXJvFqpWw0OmXQs7iwAYS
tszNGd95rNW6MnwgJuXpwFEVDOLEll0qfqrpp5yD65npGLPktlarG9KgsY9epUvg
4LQ4pvp6Lm6EsUPxHFZY83TV9+YDCfhxcPQoK2ksCGWPfHyQbyoMX0SjU+RfVUmY
3c3bNLfB6jlRwoVW4DkMFXYMnF1xa0eKbYzAFBW9/33MHMghj4Roujp+KZcJPUx8
bMPiYVb0EHWuWuHuo1n/Tj6yVA3Xpbu+IS9/7pKda25mfvWZH+WxKvb6rCUM/++T
YUdyB7xjiW4doOZBEQvJuCOMa+kZyEvs6phTbv6WAy/QYQl2E/aYPqWiaVzKqoiS
VyyLwP2kp8KreaYZ4gw+JjN1hfbxpHwqDmw+oEMNGetbSTmQUnWp4UJ72Kc5W2VZ
3VR3aA9gDf68hY4x6Qqdp/FhGp4s+Ov0bsq6P6wBjFPoyirt8Mzg+qXq7if2wnzu
YHSzChHFHMKap/OA8ZiKcsAkNBWyKNe4eXIrkdheNJ1LuLrymPhVXRFCZESWCMIm
KVODQbxqMskuQ8uL3KUT33M/gEveu18F0IkhWpx5WwwXKUn4O9EiZFQLK6ZgReag
UvxTB9u96NCy2hIyM1EzXqs3TI0v2reKZnm7ui+TA3Uz9LlKwtAYmv9gftGmjmYp
tsRG3yfriUZuILFkH2KgCFPr+P+3JLsEcwvFGeGqnY0+ByVjXXf+JzTC5AvVcxuc
Tsmp2DcQg4xf6/bTp7O+srzGyVUSdZL+JVdhFQMKvQpPVIut3FXSW5dN5AmnGEfv
aUUH7cyjV3bhEIlZtB8AiQF0ObsLOhYuzBqHjri69FUP+26Rcz6PV4vA7kTA9Cn/
zp2h+j4b21yFQfsCkUf8uU/lUKujAUxUqyLR2My1iDDOKEcbTXT6ih09WPGlCYUJ
pqCzgG/Ifdj+OwjMx+Ew3t5RuItJoYWBnu7Y0DaFeZX91telLC0mjU39xIok2h9W
g/i3eVIvWc7DWIqIe5Ia5umi/7DOH2NTDazhe1JeaaFzhjA3dHSpVQGGLoVWFeLv
GRjkIyiNtgnQQXKlPUuCx0VruTgxhxWq++HmfBAwbPI5TuP/dRiSFxi+Q0qCTQWy
2c0C35if77Imuo1ly+eaw46/ZyUHoVUJQhkJerNAaQZvK4+At8TZwOaz3cBuM50E
vtBPUUMJSKNwWGjuW45awhH9ye7I/EepTNqUiga688nl4ld01DjhUjflOXYRKTq2
5d8SB+IseRhgmFVTjwP8JlczF32SWlc6uoLZop42q3CbRWDTA1rHlMb8BwNP34I9
vJczLDsDIt0hegD2wiIUj/zSyzYi/L4Sk52wbzEV17XZAtLk5VW2Jiu1lqgkMoPw
6hSn3NqKIwv8PpA0nRblqzwaerIBKUCOXd52uFms42hGD5s9tM2+sv1XoOLCu+ex
DkUnhDf8Rrg6T6eqXiq4Dmxe5LJnEPQrMIWDMlSz71L4QGYBk5YCVRrLS13wadNP
u87L4TsV40W3UZ7IcuA5z1S6A7Fdcv1OJvgtYMl0bD6AsV4iXx6XpD9F1ND2qDrI
OadnvawHZ/1wcDUpnq6Bw/r8mcPnTNE0Cb8v2CKwygSZlmBc8U39UZ+gzp1vjdKb
VY/d/qv3le+CKx1S/z1vVfeDN242mZyJrfqSL2dmEEjgOQfyvukMcobffDsj0gf6
FiJIhUlv2PzoAtmVQB5MxVS/4cIgbN2tCHAMzHK664KBkiUNCM/ls87UhLNfj8ZX
0jgSFHTzELPSEEN8SECrL87HebtkvqayYKwHbRfw1Lp2PTfRfBJudT6816/9PLGv
gqWP/zr827D3vHsJIKOvBj2ru4icGnqyxD0vDZJ1pkx3Moy5FgVwqo7ye2b+vGw4
xBl9PWIE9Sr6lpIWZk34lxPJORpd1SX3dY6Z3VcYCPlbE1Pb8gKqv0jafyeBA3ii
dILli78Kcw0EtqJawu4eDVwUa5N1UvBHd9ObMr3AGTqeu5FEhTQRSWi8Oi5fAcdC
XYde14dj9bfS6SRahxyUXRahnjtNeJvPqFDpM8dtuJLs+rYA5BjFR8Lhxw9WMWk4
X+yNKE45fKprcDITweaEMRcX0Y0ydRY5sc8SnfPOEejNHrKC9EMtmiqK509t6cIW
SXWRBJuU+HvGGU1LCzQRVTPK6Aa17S5fNYy1dHu8/rGeATt5QvXPBYMd9KSxHwOM
WQlpD8jxquWMR4SAqZ6alGi1vcccxwG9HQNdngwwlDa9ocEEJITVcVzaj/GUT13a
WLyScscPmpZ9x1wgyRrsk0X0FRPuG6sfQIMRoXgXL++AsAOWPdSwr8MykTlRWsUO
BZwE2ZKS1CVk786DLJtmct92VuIF7apfFntNzPX5r9Z9VZ/ysozyEdGvoT/6otaT
Q4Ao5sDRxWlD6F/zvAeINKILwLfYF5DvZhpvBctNZ2y6ATVczmljxc548gTVLYWc
COSXvcCdJA4tf3ABELJLQHkFRwQ4UeffWTA4UUZkMYFElSp5kETmi1m6tO2UI4W1
xY2/qhKYIkw9Nc+4TCe2Xxo9IpqdE94Z9ety6H7bB1lWVYZ1ezZbkVzK3/OneCNi
8xnd/gBK9wSGQ0DXFepemq4SLDFn04QBkNuWGvIxqPh7LEbvR8HOS743rsG75ylZ
ryFUGqApYZ+fo8d5yS1s+LJHJToxZFg7xQe+N5c9FmRdblVCj2m59TAMTyazkhoq
DA1sAaMRcWzWCCsncCetNCl3XH5UTo5BtBMGgoBia7RO48RM+WNjtJwXRz/V60e7
jbHELwAasy+u5MAJoMRIZlwsAwowQ18dWDZBvAZMPXFxaWro85GgMbJAaIvDBjIX
4amO6CAP8UUgqMBtgUoNellHCTg7L/gRE9VrGtGCdT+FHT2O+GDwHbFF6vqNIQzq
f0aFm0UWyitXGVi0sTFnVWvUVu5lMLbylgHS9BHulQ3pRoGSxmjUSQl4s4hb2Ajo
QsKEapiQOaeQbk+y0yc/GkrifLyRkWl4XsWpPr3zTK1PGrM338vwS+byX2D0/unK
S+TkJ/ylm8tTepxK6HL/A/bNWFa5XqXASOK3y23ECXaTjky1MlqzNwSPKLS0WyvV
HFtVaF1cz5T9o+48N3j3/BfBtSUk4IQV24X55tEht1J1aKq15PfnK0EeiMRL8Rb/
lGrwRlbXbd60BpCVvfdNEFT9F2j8hWLHey2t2B+3rBxUQDnjYIYuiHfyjCHcxgFt
8h2yypFEUydHh7ZGpHTEgFzl8TpujLgqAingdGCA9EWHVrpzOB169y7U5P6cIWmC
tALCU6J+S3k+SXNEvUP0idfFSl9S+MgBy/5b4kVCsVAe3wsW1URakPOg2o9PDT34
qzbg0tFzPwWGg3tXv419WDJke7k+mFxo6q+7YYP6ZxaRJOxhXDOE3rkH39Y9TRqH
RnRyH/pD9MG2PZMNsquDPwCRaSlja/Wu/t7WTCW7GU4acCGjkF+tEim2qIxzH6Zv
oPpxFVA/SfnVonBTmeeCkTNCXC3d3+/+O/IAfeBFQyPg0ey1PGwR4CU8fkkzkIDK
w8/HtaIC2A5fLtfjJnriyDnHsEeOQDREPAqdwqC7WskIs2X7TOFxrz5jAk4weWlI
7Mipi10XctyF1RI8kodjPZxNpeURpz/o3DdHGP3eaPlhIwm6p7QaVtLPKfnq4Kzb
y0Rp83hY1wPyslwAgUwEm7nBkzLpu0eD9+5efGVluqEZeF85DZXq86ZvL7B67Pkj
k5c/z+99QQYC4CfTnEv9efDuJs85An1vESmnxDkSHfVmVc3yEs3Pr81/olsbCULU
cicwskl6P1IZhtq+kZmc5IXMPd4jqiGNfmRHcpTkbx8IRRCuEN77U/h7sBcQzK6t
k5rh8f/pZkoms4DzgXyH4TP1lbeqkmI19kk74vTHUBP4H1Qo7Hl4xdZpJecjkMkR
3cavXNY6Zb8PITMXHtcsGutt++ojBZBn1iuLQ97cHtcGB5sTc6ilHzyuHLuQ6cMX
K6WPw1YWOGcgWe9HAqs3cle+muCQY9kutIRTM2RY2dlJ6StxH7yM4eTSGeA519X4
LD6Qgaoi2QRCHFKnkDet6SusJAegq7efL4wtcIGWyCJuodGl6Xxf+DoEW3LqfeWT
rxdHpCd1nLqfM6xLnphaROpOPEvt4ko/feqpYdQvvgXk0356IojvixLwcPpnIjLP
ODLlmoV8M8hSlfMCdtFd0GR44uapJFyRdrEUX1IUGMn4QDTbmhkGmHAM7nWIyaR9
WZFjuqVzRE70hryro9WD5M6hnWdFn0/e2GsmppIHfq6O1tuNLrWyn0QC3yyyrlZ0
FV56I2tKADburekOr9DhxT3TLOYgYkFTW+fqnrapk1E8MyFGfKujIbsUexdu2pZX
8TSXIR/m1/4zoLToYcPzvUatZ9bEwquJXVGd8bfPo3foYsrVz4XM4227wYMaZQaL
tP2kg/tIDz3P3LhbGizLkb5GYKo6r3N8qFkgfVluHPbL9aID4rIibmhEu4Rxan2K
qlaGvSorul9/OEIr1LUevfqMJRKd6UA8XNnwk6o5n9DM645+QWh7xAbfKszKzRJz
5q2ghLhdLDbdTUx0IFW/4h0tzi5reP51q0ZlwG4v7e8RHAFy0voD4p+wzxh9iVq1
usgRJ6+RMa6vflxjT+Y9onTMiCxZpRFACZuuBCNG4iwjgwFNo9oywo4h1LCiqEpz
97uEcRfCwbmJMTsxnToznPv60hbOeEbV9j8v8Grrwzic/1AYpu8lfVfTmIULXkTq
USNeEG+ytHG4Zmvsikzr7k1cFSWN1v9AudmzBYcSjyK9wTAAlet2nE63lgIv29w0
pskUdmfSAGrMBcaKAjJXT/+1Kue705rSx+d3+gDWwkYNWvpUSyJ4xWy50Bx+4zKF
NDwqsHFNSmRapKBCwUeE4m75e38WwqB4d9NtBYUsEs6WPUhwPbfuTBYbnqSSArJW
oW9Y/Mss4991mpqm/Fe5qCqtZMsJDSGUDBHWcz46gQe8oHBbj3wQCUNX5fxf4C7l
ze7cqef1LbMktYwrlKD2pveud+rHwl6eu2yBBBOp5B/sWxQkmcXw1VI2TMFfH3sY
cfpf0C6LFj5XlfOIMEyPvzG4rK/gbj9EGUZ3U0O5w6brS4SbF9WPorgxZua2I2wH
d1nfbbd24JC6PtttKjCIDXTend7Qs3wVCjJts21MOK1deI0OBGD3+u9L+/KOLlzU
4bDg/M1WMCU5yJLUApUnyGx3K97emqYJPox+fBHRcLy7PI8fEd3ymGAb9aurbZZc
5wCGXDUB4lWR05pgzpJ/XcKyDgY5ncm3qZdC2uB4+G6J8d40e6PuPd+TJAIdcvRx
izID4og1Q0S5xbUKvNJ0tMqU2RJhu4LnWGn3/eEG8gbi1ART2MVYTrtx12zd1OUu
71RrWARKU1nk3QaKtpB2TiYjXH//XewjmAINejzlIM/1pncuNc1jnkq6CopDEWQy
+0IcEKAG+yFiRpuE8PhUxpnMqSRqe+7NMWyfXuAxcnk/nUPypKqR7KJhqSjO/4o7
cKPtTt3kspzDsyWL91vpoqhk3E7jCSu0mqWl8QnAS5SDa5NdubDAWN7Nb5Fq8OQM
zwBqN/kJPx2HxKes1FZLVRZHm4XBxRDYSwi/3kM7WzQE+fZ7oZ8wrwGGiEhuPA2B
riJrdZmIBeokRiTWnBllDldGyDATjsqNwIlIQyfxksJkXF6ztLGpHMQvERCRH0tv
yrQwiJ1TcyOElDR+6qToWIUKw0tlgRBCo6QWz8gprUwqOm+suu2LF8nvGW8DbOpD
9vbduZyq2eQU4aiEng+7NRafMev0/HtMfwd3Re0fuIDg1CXkMncCGQEawUsn3ZID
jIImVEuhF5BKveIgLLAvH2AjccMtFF56N4R1G5wINHRpXlCEgnqjZ043e/mdwJjw
vxijkXTyn+GV109qCAJFEP8DD8s4kstlZYSXVu6Hz+OxI4MJEpqB/UhK8IDmNg2g
UYmInH6EmiXvP10QvIKlH/wTubdr52m9OYDSEYIGqZCVhUHpwRFXiXhiq6p2Tgzx
anHY7yINFva1dGDl0sl63dHcULJB2oSoAWBafzuEN+Ayn8PhKdtsCxR1D9IquRG3
mQvOYupedanv3oKUX8xTlyilyb1i83b/j1tANAmnl2RmgkjO58mhuDVg8NSQZYWj
xUEEqMgl82a1pnvTVMmWSYhjfVzES6WXjA4q7tYmcopH9yvoIk5Sh7IT2sH+6mw5
C1l5m3WF44M2AERFZcSJxPtROCb/kFbVedZiWM+UlJQQCUG/iGOpE5SEYhxx+y7x
0nPHnGEVTa9SViDHCZy6aMqZs+xrTe6r6f5zNmZz49zn+Rxqh80zGZNwpRu9LLtY
dJzoIJ9Wemq54lL2eY7uVmBGByUPoCml/ctikkRmURohXOETaJhhtn5dYg6YoAkp
5QUcFzENjzh5HpXErvFM2cxaKWXKntyQKn686lWN2UFUELEJvi8gGM7uH91S0VKK
oQgI8fVeNOI1wAZ7XdUL+fbFO4U+NUOuXG0R4bFGs1v+JUiRHdCJh6yekV61NkKV
34M/JlZgOZBH4cYw3dweYR5jiWBNOjipydNdXKqfVk0+6A8Lps3roT7Uk+HokeOz
B5SDi4v2uqIWVNquV0L1AYRb8vd7KWnwqrAOh8VGFw1Uz6s7hOPrDI0Dtsp8NHcC
RUargHzN5uzgaNDl8iWvw6sYNmGVtzxWkKQlQREdpFkRdO4MvzMLCvssJh47dyjB
+nYcSa0WUCHt7UMuprWu4Xf+BTS40Ux2anOU+u7YPWEsgwGCaDkrSn5BzSISeZX5
WypLQ/FPPMDojiBC38FsiYAuF4Jp9KyYfN7WQYbItmzNH6rhNAPy++VoT7B5h7h3
yz0avsYViXfanCs5rqNtuvTzm2g+NBc9rXc/V9aQUvnG3QevMpaIpYlvPvnGvtvT
VH5FnNOIkXsyOLGX00BqrSvPuZzu00qmPGE2djalxfJ2rb3WUnnDrHXETeP/3YbF
uedMHvmMLEVex6EQDV3Br4ElrbzQcdfN8d+M/R22TGARKLY3I0JeSmman/z2Lz9x
p2yB2CWaVcBrMuermQErVTfN8O4yqfMR06Re2NoPdK9LqArdf48SxazbjHcBNk9V
hocG+v3EhrkFozbdYsKVanDNHMOm36BF5CibRjXSVoMo/SwOVlMo7dxvTaZ2fJfj
TZjtVw5lRK9K7hkwnUClTKC5jFuf0dhEOnhB4ZQGbYOyrNbFhv5VAAkYpUgtbhbj
fjSihJQ5WP2MufyCF5rkMt6DTjfcTSKZezhA3y7s0B7gIzOhJARJbuObYCHnEfes
oSkp6cB8q1nY9TM8SBlm3PGJw9Nz00wDOmiTOCDmCVGrUwGMxdvRPQilkzUZivtl
UOE6dh/ryuhOfo5nJaBkX9BqrShGQLFYbx8qWZcmmKiCzfwqUSSUrSUgTk2v4ws8
JCXXOBpOk3p1HYPBRZXtieWMEq1AdCDm1zepWgXDHdGUbMszHfgC/hB0a+54Uwj+
//tFQHBiOYtNx73N1zKwpDmLkoSRWW2LlHxLIqTx7ujcelSUTQC/Nd0x7AerWCN2
jpj7wVRxexxRWgtKRAWRLVQt304sAMeCdDIctg/IqqgFl8sWkhQH5u25gWYpi3QK
3+wqbhhrXtKy+eJGcuKLUD1P5CinHx3SZRP+ROxwzgsvHGhxahLQ9qE4Duq9cCPh
880syAc6DCi2G8IiiluffLm82ApE7xZjtBobAgXywU1N1c8Qvqf4dqib10TMitJ5
lownlZIgUALLraMk9LsvHuvDy+onuIiYLVKh8Fx4YBXHVVHT2V6tUqCWu/xCqhEP
cXB/MvavL3qIeKHkW8HMLJWI42rnA9RqA2r2BdPg3E4ANkyf1XDH13gEWWGkJg5G
O3or0eo9zyBgUGep09YAHvBLk6OlWeHUgp10wqFeLOpgxMGH/RY0ETKS3P2oVQw9
qlH/PKiatX/PFHqWiK1qd2dO1gGJ1GG6wFHAGzj+bX3tdrMBuSWHbDqDPym/gZKK
19wbrmsVCxkH8DpF9YkyIMg7515Ze3ZhLrGFFzAZDQie2yTBMtZvWNGDouzgHiNB
bqXABaGDvg2eoiYlUEVlqF40rP2LRCVE93WwabQvDL1qEaLNTwXSY+M3BtVtnDIX
/HmPp89ug2ZBTfpjsR8pSlleB/h2k1k/kzgKxsGDEa2MuHizV5BGHjUOGQtKlgqf
MqbEze473jMeKT8O9uF0cicJRwnolS0EzyBTuHuhQ3zVw8H9x1ReGamMeITYAuw+
keKpyeGsk8XFphVUc1Lo0q8wDKR0cVzMOozoGcOyGZG96/YmqlfdE+ATYtblX0wC
gsrT3zl2tsTkSFLAH+CrC5XDAtBCKhsA4Z+P/o5HpL1baYHgmzhHF9AZwumRKFG5
FaNZ3+taCnYFGmApPHt+YAhcFSwZS7ONXQxW2lQ2FDrMJoFbAwzHa0MRR1k7KN3K
wGMR8c4OBWEcA1sGA28zl8Sdvvl5ERfZGP2JZoGpnlzzGuyruhlgF9zAGjcmOxFa
ZOGfB3IPjgBdC/Y2eRKT4uH5+RRB5yT9nHOomduPiUH4vpaytUmtJYRIbwDBj1yv
NFpeldtCzXB2AvbW+JFv4eoELzngTGJmwZTbBjOhz61Wndc9I/LLJnDrp3PULdMo
eZjI7bJMuabvM90vaBk2ZWH4V/kAvoVriBdZJ84ZWvvkmF+1trcM3sYVw+GCX/uU
sOFCjWhjSL5s2FZxUjV0+Ebd8SWa3rDYN4371mGa5flk0sqt8VEHDgz7WoYyN3Ck
kb9fEPwYZ9zhnfvOaB4/2e+BqxfTnLY4IcTw+tslwyx3Gr0OUZUvJY4wS9nrAlyW
Y/rRjsyXSBSXcQxUJ8g30BvYmWQIMUTMSoamiKJVDQjMxaP/dCh5haqWcsXW+yO0
JPB53pqY4XyMHova0xi3dheLn7Vxrj4PYDcrtBQmlR2Vz1YhdjvMMox7Sm8q65wq
lSHiOdDyhO3DyDMf4kT4/y6CEQImjRx38QVoejssqYNNG9bq+bqW6MsDgPya3lS6
NgdRvY7jFNEDibbH5OpGoJ952FInvpWnrUY8z0mdDSVHZ/Tzz6681UPyhL1GPZic
+1K6fI0AkZlmW0wSCwG4lU1KRBEKzi86HzOlHBr4F9E8ejGRsF5DpqnJ/9zBXrfB
KQ+Zhtog0xLFCWlIU1OQRS8jcZAqlQ3P7SdH1AYGzGkPbHE68/Qt1djKlm0ifSaJ
yJrIsWZl/WVLlJxLebBEiBTyuuJXgCzewXDo9IozWtrSQnGHI3fSvL3w+XBTT7V1
qAtcSl1gQVZ+tEELtCZhbw2lSvyKXTas45lxuSXuHa+h+ubJ5ZtRDo8TZ0ON+BMq
P5YCUWqgTGWKl4VCOlqGzWCG7+IST4FFtLsbvhuOFl6ZLOrTfWl3Tf6lYCZBijMN
jou+T8zS2S2C0s0Qj1sOVhdVnIKekzkL70S+yciw4D7WlR+NUr7NQH88TitqbqDZ
hp35Ib1MyXnSHKsreJyO+L8lcX2yO5vHFTEpp3dKu/QT/eVEGRpOJb/H4szC3zNR
opm80SO9Wql8uGUWQF9ChlrcmijNgW5vRLMpF/tbcSljMh56FeTLiAvUMAFdPxia
w0mKHnPX0hqUwwU2Tyj7j91b/+i7EO5+Wwst3Y3+V6SwPa0vgJYuyxGNhMNfB5FR
qcoWFprvd3L87e1jmBqn3Be0XrYd5jaj44KyszjdZrQHEy9OU44SXDU0yDHaIo/8
rdQl2ejHFquJusj5/zu2IEHvNqCWkiD0A+SAHkavVa6xD6I3yCR5dcpEuMWVuDSO
D1IRocyDdODaUCDnA+kXyfyJ8Rlg4XGS8kAu70xGjff/U4bzgF6stm55yCdcQF8s
t3BpyxvaiMw1o1UsdE71VtgXPW2hDIlbayh4V08YIpDt8vUySE7Vr6yNZSR+jAcx
smjnKcpzb+OxFKTS7pyBncLhPpOUkuOxjRkL7+ZFvQ04Thn/nVHOwRD1YqwYPMEC
eB79AEiVFy56/sLTiAmg4YwlYSlvwXJ5ERL1iHaFvcD5DxzOWIZU5NaoR1MBT5aD
G94j940rFlw0/ygIxAAyXqtpPBqV5MDWXdLtjIjITR9Yzb0lohgJnu9FdVRE74T3
XA7K4yHhGODWjTHmFnOt4/oT4BfmnJ8zLs62abXe0yp4bY/oTBICmd6T3kJtJyOJ
jKjm5Qp2+4wv5j+59aTO3/O1CAlBPWasp2WmPFOlUpYsq+WbTCTRp4OP2a6ftpHm
z4g42X4MgRT7kJ3UwMyBVJBKPlEVwNCtMJZpGnCjFFtP86nk83l7pC41H7y6/NBL
HlyHRbjBspeWd7ka79gPgiC0OabjGg9AmVqOtLvlDy7fGIoA+qYYh4af75cnvh29
NjWZ6BGBCfVWRkbSsAujShsl3RwCt40E+3js9Hb/8aZgbpeErLifsXJu51rx7Jjt
I9CT0YYtBzZ41XnWBrRdp/rD6yTei2xd8b1C584BuFMfgNecuhv2lqkC/VDlqOG5
VI5SdWgmeS+byNB3gTwuSzRhwB4Y0q3cuMc/8oWs9TkQBeoKUoDSfmPC3/VIXdVE
LFyrIKGCcpOmzse2daMhLIGoVMpKRdurC8OhSymrfoITpOyCzGAwRYaK5H/6ri4f
mkzOdsErSxevmNFSrAXi3iZXaxHimvupvgAHQZEDmOW8J7+q8y+eup7kh9FRdh6K
3SXn5tpLRExamLai0Fjxfj/YKMzXmMpECRwbgWcRU2YJedoNOdx+hGFeL4Ir1Mgy
celL98jtEqHe0xAlnTlfDRz/R5I6MVcwz0QnJsTRk0cKwWQn3XWwOfGBLo9NaQCz
gc+0BGg2ywodxg6WoV4AVfoGvagbH0p7n5WESQGoev67X5cEk4HDso6TLUz9jUWP
4CZYveRb1xkHgHPb/aySnJW4KuvOi8ojI8b/z3LbPvmOOjfzCBvLCC5cfTzUO4bE
TAppEFFMHqtLyYSvNY7ec+viilAAPyBsMEh+I5Jz2NCOSzfrXgL1+87dzZWPu2xJ
9Ab8W24ddilh8ww0XmOY83Xp0yr5B4Jh8NChwdypypfV+oTrJxQlwq2mrs5MTfYL
B4GCU0DOV5UazBr9D/KGINU2VeQ1D//sgllTg1YiUsqatdBFCb9JPdwkNaesynRN
mYibVIqGjJCXfBRyiVKEiCfncHBl9dUFwoBMDj57fX5p+oiFlOunwhXKu+JWiEld
1ThTuuAJDZDgrBATYOgKEOvlFOBFNbY+pdjIuPTz1SXa85eDpkm3EAvEoNu1XUnx
th99x2kePbzfEKMRWiuCkkFaS8VuA04Md7r3VgnlZQqv5e2ryJLIUv/rCYXDrpwV
NGyUspxkM9o/gaLKvjXgBdNQMWGby9kIF23WZFL1reWRJl5f0K7NfA5fu62j+AvW
KIyWF5bnb06S3ZzTogBaAWMV6RZZlSJFJvXc8jWo+EY32eA88va9As1t6a7gUQGf
niWtW8Nl4ovAF0s8EKFrEF/kuhF+d1g8rSYMmyT6QGYTMiG0+xbBTm2mNkZEjDEz
c6bPyrObkqvJzkTZHHXihHuK88l4Pwp0krMRQbsOf0guDHTZ/TULWTEB/BGk8G9d
LUTM+VV2eIz86oVP+GqEBJpg3Wrjv4GuQoPjGdv9qMOUufKZdUQQCkp8y/falrM7
pZDOGLEQMS4c1z4auhQZSb7SR+ZoNiPSy2s6k6PnTNTxJKNlBpJWjBxtYK1XWjPS
t1Jtrs2ZazRujWmTG0aN0rc/mSSPHfZnd0gS7dL2ZvAKLugGJyT0o2PXQq+/9Wsa
9ugXBNwdGXns/canpTEu8s4t2bzFqqjAIuM1LS7OYlpMciUbnL10R81OSqhDhVna
zzxtj3HGtZeP8QbX0J8W+s1m55jv/D+4nWNJeyAxcMYvYTCJb0jjkT5zw6KPz6QA
NAsXQOLLQFtAHubFq0ZsDV2iAFSj1MNqdYmu7WfRMn2aXTw8KIHdToxyp/HfhJij
yJ2aseZeHLZdKDEEkYsv4wHcXCXwMIHFwN09d/DEJN8SYw9uXrglDvbk+e72TfTI
8fAchFCkJ5n4Qv4WGFMJHNOKAwpA+66vVBtrZhNGITdVNu8xIdiQBN1Kt/4flyzT
Rpf5NMCtT6MAIvswULvVLYu5W5D90bzB3W2rDJj2jVCTlee6gDKfVMY5JNrOymH/
SlERJyBT34jLwv6XQOmXXOa++xhTciv9mOVz9p/I4iMYHcmJDL17Kd9Nl00n8mQy
ml1rmox1O+KiEKUDkZlf/eicS4cZ5ntGyVf3UTEcPCzKgSDuwbumFgTFQQHwSlab
1ZBksCvdBRblGM15A3DQuSePb7jdnI3SKGucNBlK8MP313WfRefnxLK2moZT+3pj
EC04Y3FVmqIQ8MaTaIlewaE5QFNuFaVAQXR6Ex2JBzXdYw+3i9IUrjfq4nk+Hf0Y
zEExt8Gfx/IK6k8gGZvC0CKix0rKPtmoou1p/UCKTq2nPrcVQ7sd11PUf/C91lbQ
iLllSIz5AJ7pOJe37XLhhL2kxUkYIod5XoQUZGGDuPy6gPV0clkMvHaxITaRArgc
8c8nIvgfZ+LwIEIGtujWjJn10QfdD5L3/UpXW8wV4rZh5UBWVsDV0j7vsxvt1quV
v7dTT7xXOOeKv25NbTdB9ogXDijYVodRaaoeScHwuyxTWIoivRHAzYgGwyv+6VTJ
dJz1GObH7fpQI/n63AGIHi+rI+iiJYySigfRSZIkaBNQPaE8IIu+fu0Vfxw1eWzd
6bixxjYxjS/ZPoajtHDGecEA/ilLAGfm4BgYxFitvezHBQzqZtnE0FDFsr94F/U/
YYkT3nJVpQq90k/aR4xJKyOlJpfTy+t3ZKFyEVYtd4Wn7D3fnAvWrd3wgl7qkDZR
D+rQm2Z2gFkIZpHHnNuZFmL7hlnWU26tvVwiHxSwcpFo1XeVdTbKSuODJCuSgOzA
NMpm9PDy5Dr5d2cAazhgB8/BrzX92ARwImG9FYeBwQeB7K5lVJ6oeSsf2iHyf+Id
wd4ryxIcaXDcjIhNQBzWF0dVuVnYlbBktUDtR+XlXx2mUk9rmExNajoeMSW4GzK4
xJKxGbYBIXjatqaaw6NcdLjjld5dMtffmtdDsEwrkfxCR70DoUjF3s30XKzwzaLY
C+ln2xG9IlhIL8P7Y/6puExbOP7DTxwYWJJaQDXRV/2McLmovhV2KHgKZJv63WEy
2ghHVJRGIHYT+mIjLrir0ocXWFZh8YLNdEg4G5khG2qUWaG0nY2+mWxIEaAAgizN
f2b8Me+w4A3tsO/VmBa1UlZeTdtkeSpVO7k/G6pLb2mUVzD25VQCAIE8FBuRo/4L
4UDrYFkomDDhxyuSuHr18Cii4tmX1Fp1l82B9PlfNMcB7R1n9wuL6rn/2ONW6DVq
7WMJ6abMYzw4zEsk9DdvcLH6KT8gjvtk82EeAeJQb153NCK0bfAbAInDRWQwEm33
8Y4ATaRPurvucYviK2kDrF6MnH9LI9ZllyDn53iVTl23BpnAC0r8FHvARWWToJHd
o1Y/s1TO6ZgjW6samJr9Kdxn0MX6XTwIrCPbsu60cSR2BPcBCAtc7YEC8fv5SqHT
bLhf+M/1Hm6P8/aoWTE/G8coBmIawtwGzV1/56P27iU1ZWwx31xqtTgglYYOOF+3
OhcJ2ftpScXrPmp/2an5ItpdfYsrpdAf6IefX31ydRd/gm8VvITOqUk7eDvkCtlN
od6PJffaU5IyHg3RrDZ9zWzuxrLOWFfROAp96qI9wy9Z0h6Wh1LvqYNdojsFm986
e4YKSsAqLS/dfD0AlHyZ5wK1iUK5TWFzfuse1WU2aZ8byPkSIRpACKn+JxY+aamH
WEd0pzNbV0NXJWGC3vUloxVy2kUIYDPrA/uiIqgNZxaNguORw+634A80r9qwdQue
UCcT8eB9GhoF4/7GMDpjRCp0EKkfIeyNqn6sPJzlW9vrBNNt/zwwxoWmgUigd+x3
njXzYDh0bxWjEUD54R/3KjduD+WwQRKYlbY3HCjPuFtQa2jTxQ49hvzpBYB0iXQl
aBlkEoPWz0y35Vw8mnfrJhv7TlhO1H+33Sq6ghdgFF4LHYCiAvC7AZx4s7ppxYNq
1uLNcTP9sMC9aAUb+rjK1MEPnN1u/OLxLy7WMCaHqbR09Sei769zth8hNfSa1J9F
8RZPi0O9cILK8HnxmJzzBdy9v3EOmwH4PpPiwE40X2acQgmj8v/ZoMJIk13gHPSk
kXh54zUQF9H4vPenQC52dj8y/5P9LCzihchKPCbv6YcCG5tVP4mx4B+DheSIPGMX
JvxQ9IUCy9XBWMJz/EqjgJ5XY7QFd532Y67xoEvIWrtxx+AsrVhQKuK3MDh4YAbw
CdFTq7tE1ckWZQmJQ4CnRL2KjLtc1YRqEyHSpyzmbc7Q3h4sAtBnk4J3B2VlulDq
IRGOg4mFp7iH538/oR2X+yB/VFAzfb8e4Dfv/fc1B1kkdYxdbERRMEiL6p9F9nWJ
c1XcKcGGeStjPYCBUPJJ9ErEhavKhkvpNRA67BtAtVY3urKCcJfB3ikrKxMhh82P
5w8a4fvUK795CDGgU4ap6r9G+hNOhZDQUjAe+UWVFuS4jLGEfYZZbUPoJcpMOFjS
9q3VSHsVyqSfGaqQMQJouWL1IJRfv0/UVoTMECjp2lN/2+eitGn574dVznba+7kJ
GlCgfuSgWAX29eBcNILQsN9JwRRBdFcP8p2zYKp9+ZnbIfHGNSdjZRQWw2VICga6
aDY1zvXCYxSa0dwe/miV5mazUPb+mXhcJg4M6q2/MASV4a9f+fZgRWrqieyulzrM
01KYUJ4o1wZH7hL1fDczP1IG24D0P2qW1eY2M48jbBhvD6AA0/z7ceebhAH16Nal
MWiI0ZYxe/sUgWU3NrCa8jRXaT9Bfq3VdTUsud1izE35O+eqRXC7nD86CqI6wjZL
xgwCefLTI1nQO9LvaTo1g2YIx83z14QgS2AARdo7Kys2N7dtgaPqF6P7OyI5n1Ef
Ge0T8rWXVolGnl4oKn2sU7RAJO/pq21E10hX8nCizuO+Ek+lS9b//kQhWbSipjNz
RJH6Kk4o2vQH0gTgxtY6LTrd09QqOsrPlMLXTUftHL5w4Vjc0VfZ6MSlbhyU6SfV
/GpiZh+lYRRp+pwH9HJCEbq1fGLxH3nOdYy5xDxpSpvH7gI1P8sbmfSL/8PLbvPl
rs1maGuMwRDLHA+hHwp+YLKNBGIzaq0J6eYbnrG3ob3kSdRjYbWSz0JLltHOuTfU
yPoM6WQCmaPBJjj+OY61uhtxVWPyRTWKzIcb7LBTJ3d6CarWKz9AHMqLGZbDy+40
OSfgUDiCpfWnt5BLWu0iRJ2doaUiQXclizzgZhcP+i3MDjoN6fzllJ5j9dxmKKCO
jfuw3aSP195/wEUO2flgB4bzdfw8LO0JJ1bgfYeXcM/7S1YKs3Ju+4WjA62M/mGh
GEQCzDitE6u0P2mkS42lGiU4ZdNSS7lxpg2n4gGZOTWld9Lil6bg9Nk0NqVsw0fd
m7tvTEeXBt48uadjQ1nL0xcURe3JAKlZjUcycQW00t/9vgnGzkJEXtCDMcg0Aag6
cr7m+Fur7EhmLvCFLJpeLlxNlgt5TyNAcaRVG8rcFdYFWm0UGC56fogS0TbGcxiu
bkFJ3Lxy7mi8coUcwco/beXIKWO44gtNJ4LVJpYsDgrf8w07Hjzbn98G+UOpoDX0
Xy8UOzmaaovffRMcDwZorrUjRnWt+pUfZX1fIc4MIGk8CJecfqd2+gKxSg8AhjEH
yoYop77wzJiLaFfH1E9Pe5G8lxo/WvrHgpj1GZqi4a+6FktX/9mK2P2X0tZr4+5m
wGAb3brPJjuFQpHEmfomZrLbih33MdnRF6DAxpeByER1IvlszQp6LftQaJe+4JK1
Gg1GlUaLhOIYo/67q6FiWISVaQfcN8vmOdOx79s0jd2Jk56pYjd/FiGSQ/eIJoJ+
wcpvSADjAL4dJDhJojOvbOzijphSRicI6PphY3P/B4Nu2Fvz2dIu4BvSvFmSUhXL
e/CAcfIniFWwbrDg21o3bcldUcgY8vy5q02xSC5Hgt8bfEXGPUkKwcqJFFmVYEaA
W8dRtV7Dl1CZsJGn/JyYRUH9T/RUIY0m6betqiTMTvp95kKoIVbyb+FBAfdlqUP0
SsrbGiW4DZsUV7Xh2H3mU9HK3rSdQVfsuvUULUR0wHrf5h+/taczI3YuVlTB69mq
vDvSo7F0CcVjyIa8dR+uLnkKyUaPf+P6kDvsMGSOTpbkkvbG8e8/tcvtbIjo428w
MJFi8EF8FnD9n/zeRRa2Z1ZX/HSp8f1sn6UdLLTJUwR/keqUXQwsU2DMM+rCcVYX
RfJC59/uaBBW4sHrwd/+QGVL8o0nlp4GpzBbCr3v8KCQFQ8GzMBX3y6eV3ktMyek
4SVNgOTkjDYl4ApoKuJN7x8LCexgAMXRn6dBJz/CxYYnvdJpBWs8qXiieuxEXfJR
CIN5mb4UdBytIPkPY+KWV5QwOXneF3jmvt+c1uvF4r30eaL13Ub/geCtT6dn5S1y
Ez/mXdJhE94LhO+T5dfBSv30kpYVI9opN8HpR9L91GQE+FLGneZIq833XopA1Ke3
7Nr738Ab9oQ4GXH6QGd2Yo17S46wzUUqNL+AIF27P0led9JhjwqwMDUrs2eAFKGR
iuPeLbaGtVjQMSHvGek7W8I5egWfZx1U2csfXRvo4+njz2eC70/z1qCsW2WtrS4v
Lnr1D0MI9bN4ZLRSOsvWMg9r5uJyrEMg30SYWj8W4bGhG4EArFmy040M/fE19oTH
gMi3hOrzq3yW+LtrH1nv10wtqvrbi9INt2NOSCWjI+VRUWs98fhloV5mmhoKmDS7
j/yqRIc5eo6irbJKBQhtxB5my1cZgWC0jyfHrRBXa/rN2ULDXlboEBfonJxAMXZB
7r9WsocUyuJ8P+s3thnrniQ48gE0eOi5t0oa/5mAqstCKP7PyH1bAEqInMbwdO13
bB93ki7BtfASrMfxjKy8T2Gq/2EHv3AaXsLiLAERi3qDzKuuffhFTvZq1FKsD1mh
HcZhxluRjlpqmG/gIud3JKa6bzz6V3p3EPAocb/1I2se5wgwNDWos3/F+7OZhw0B
wH90CFoC8lTXxnIe4HR9A7rGvUdxjaRFKZjNrjaxKGXEO0hzGj/w1saummFdkT8P
ZdNtH+H+nFOJD5hPKfmFASvAxfai3bNcvDVWJbVN1Tu0tPvz3Cl/O0VCEzhwxC5S
hFmwawgu6mmOq9+Du3uMRjCjE8BVJTXcoOqT/edGp+riOYrL4XoKE1xyVK50oOLo
TxRUxXndgcX143MGIsQj5M/QEwa71dmmAihpLuExiZx4VDOjvKKt2QNetF43g1XQ
kwZG1QoZQkhVAhg6h5ekX57Mm0Jff1bExhynfQzmLNHuLAD83N1gnrBm3fWUO6ig
71hyvnC2ub+2TW3WuAhWx+hxvcoTjbAHHZORggG9cwsxkxDFt1OQAqhCIKLcuFES
xO8F/QD2/pZDStDCQrxeIz6AsdF4hwarMlYMN+0d+lwG6d8lS6p44wpZp7wqWqrs
qLmXs3pO/epWNxATGWpg23t1yqQldxgCfTAX3uGEWwAVl07bv0qb2KFrQhi0V7sN
kr1Lsw+wLo6+WTakx9YBPRu/l/SKSPuHwr/Pt69rECR1NQk2vD8epzkiugXuK9EO
hwQEuqUbtZipgMSnP65NtNdw9l/WFMTPtQKGaCUm8kZ9o8GaBgiqnYdo5Zp5+xrb
bFgrIaDA49cRO2Jb0++pybZkvoSLGgpEbHGC+T3yabFE8LjpYFXvDKrkHI4e82jk
nxuThGo6MHvpWpW8ZMVtrvbtyPzaO4BOEhNHiM7WIDZWZsbbeHR3i7aulTd2Zt3e
NYMLOQF+8gq2oa90ORpZ8o3v3K/hug5d2a/ivZSOLp2LaOjW69iU9V3V6rKnnFjL
ga6enBerH6GbdUZR+MyUOzFID4tMrQX3mjPvVz4Pvl+k0yhSR0ycrLyNvQFbkfZh
MadrHQXiUmOsiLX23hZcoXUYL0xm6dhdbjOTUdP5pW3cJ9Omg/A67Yj6qdT4Uull
gSHvyVPHIbkDg59suWco317extoUpQzhPEdaPg6TPlySQFuNzprcVbKDng2iA373
n3bMaSW4VTH6ZNQ0/tIFiT3iW+o7ueX6Gw3IjOm0W9SXr7kosC83V1L+rtNZKgQr
0/VuavMr0vQ7eVzT0+oJjcpvQ2SAFolqeaJbA43Gngw3nY/JKCIgzQKW1H3Q6K/4
4LPB896vGnX5/s/1aD3DK1PKD6KatTJzKRaZMOmBX6oCL+QzK8TuwgTS8y2e1eQ+
mew4uAyZ62Bun93lnBE8FqvGWsgAeX33Qkh8xmDH9NykZtxBbnD84Bc5AvIVpUjZ
Ao/txJiGHu+1J/KTvve/jw4lDxJ+dIGGKdyC0XDZ+NCIouT5Qjs6FM6It12gp9Wc
4UQ/dFCMdzgwpHwuSdzNxuwTk8m5en++eUkarHRlW1Fkc/2Y+smVTQlwVvt6szIh
+GriPWVzjk7BQV8lIQGvPZB4IzCW+oe1xqzAvY6eAUHPW3fTBD94lJRInsKKaZuf
5aWlF/6HDzu2YyLhe+yUio83BEHPzzVoSjYj9493BIDotlbUGn4MtWmA10ORDStu
Ohv+x0H4Zq8+fiLiNIYFakGci7hfnuUUwEptzg5uwpQn3eEEAQq5k0LqWQXTdg2c
A90Yaibg000A3TkmkLU5AsbtrZznbr2m2v7xF14LECDnTqSV0I5jl/I2HZoKh5Bb
WOXFxDgH69/CVFNS8+1HWsLXNTKusBnPVgpOq/rV9IfZiJ9EBOFjbcZuj44voZul
sMrbMzhICLQW/+X0qOYJwQll3YngFjMiRgpTvxIDhqYgRoJNWkg8QGfN9pqXKkct
r1U0WaEwMaafa2GJeCAhF9nOuZB761kXmdsQ/gjLj1g5QpXyRY6ZzeJYE51kPUkX
EIhTXTCejFZkgyB0KDChZ7+fgzT9FLmI4chJINOK1sV7NKIhSUi4WzGsXgWlRIGG
uVFyRRROsHdI37JVxqoM1HywCBfbPCBGiT/FMuCspVLs3rzQhPoAmXoOTln4DK16
ED/hc8ruPNRyQJC6iKgXlvgDunBMOyzsp5IEo8kXsqD+3A5vlm+UhnN/9MiQ7lNS
VrlEknJM8RVdfkbtFjZPzJhubs0CHcEwwgERbCjLe1Bm/xYMHzJkad7QRGZIVYBC
FRfpVdY1t0b6mdOwlPenPsuyOxmpr/aXujV7/BabnRnAVEFoEAccxPbL0CIfSDzs
Ufrry1N4jkD0SWixSRitBAwy+4Y5Bf+JUJ257IGts0c8ZT/mKqnwQAcjoitOakAd
Z2uerRbocLSNmU2/ZFHRw5HreE6sCD+PHuvu5unpxKH+o5qPKePAfbRw/Qnha84/
4nRhTrfG+FhtMw5EdeyP63UNYcE5I25PvARrXbpv8zD6TCs2Mi3Pl0z8B8fWuUSq
7XjjGPU5PX/PuHCcLta7vXyVZ0MZxa1T37PdqieaOUUC9FX7XVrNHLSNpfWNE1wO
yWBXAtfn8x7tZo03jTr+aNWIYDb6/MBDfsbRGkisgzCH8u60ceOIaxY7k6N2bXBP
t7Io/atXOdoZR2EgQnU1SReVwdc8ozdG6wb/c0shJoY+EjICP+PrIyWtiVUB3oaw
iG/TQH4mbtI/uFMfa4j6hWjBEgNwoN636VDvwrJxZsJd2nIvk9e1hY92AtS72YqY
LwNkvSybU8R8PbS/I8azO7Kwz6XVCHuBqVD96EDDqAU2LYk5KoFjdoo4oyyIhkNA
znmS8rlyj8a7XguZoyLMM5ZUM5LJklAtPCd/sBni7Rl/t0emZGXCFBuBopxze0EG
vTOZHPIJXv4Z9Xr2mPZMPdZdjhRYLXHgU0ZdJQyM/Zlr+VcLKDvJkRCoTDsggFDr
rMikgHy5n2hs6ICjOxLPT9C4GRyKmGzucnYMLr3fPnFsqVo3ayDFtc9Haw4DkYkT
pltKhi+mfT0f1ysSg9PSBGnPoNnb+tCeqkjOcYfYSgvz2Eu3gzCWl+zqQln4O/cI
Ysjazv+fKcuB9f7hfaweLEO9L7bhHI4kcaMoqUEHLqDsmpphstpw3+KAg+sNiasv
CQ1Ebru42H6wzCq+W1S2OVwRl7dCdl/DR6Q+tTgPFVloHQr6uONCdbt8n4Vi/sv4
A5EJAVzIVuqbagNv6H78F4MLUlr9XSDi2ySyEm0k1GhWEG5kcNwO1KOyW4muOCaO
tEugFHMeYlGMlwfZEtFpWq0uAvcGjo6j5fqltSLyw0LZI7zPLYYNd2h/JQbri6tL
bggIz9rWNVBUiqfDDlp+1MV8vpf540E4ktSfQiytaKVvPZyyw4oYmJDa+58W2fzp
o8AD2DztYxCCmHsMq+Z8vYfqtcWwHmnN8JPz1YCCcLOXGyglBhXNzS8RTIgFql/c
whzIR/1w7czHCz30DWufnMdAsE8/9DgCdKHSBcDNhFX71k/vLf4yIxTh+NQa2rO1
Jdzv7HJChDigKg+/orsr6VKpjWqV5DIao0TInsacCTlON1s0/EbnTRs11pGM0l+h
FL5LMi5IGAGPpDFT+3nvtsPNjH5TBKY+R9sM2+8P+db/6jkGcCWYq/9p8OLrJEB0
74ZRXetFGCsGCIRwXTPEq5nUNFDKt6r/Q8Ia32BuzVHhJ5K8Zg4vYGYXm4SEtrhk
PzdjkHLfBtc7jdiKb3jM42AApVH8Z+OZ0b4sq+/zjs3WS9i9jF0Tm/sOCOs1UNHa
RaNsHDBsQjYLOQy7qPd6mhIv/h79VaTfekEWJiKln+QnwblBhk7spN5IqhjJ2h3d
4ex3ouSVzoceNTW/bSZV6qixFmNZrO1DYpXzsUqU2Y8q9Vg5pSNUr5spwyEUrKoK
aoYwqwGshRieOCwWyBfYEq9syBsGMqIasT5Uok7XEITrfDdYLq5YzSMRfNML69Xe
YzeuZ4w9OKnQQI1GXP5wMA==
`protect END_PROTECTED
