`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q24NaU1yrt4Fw9QPH7e34xnCtP6Mj6C88ZSyjdF/fzZh6hxjmtYmHRt578RxgBDb
4bgKa42XpyrlvBmemZbAxZMqajmAGKXZXqsJl4YOe4HVLhNlzsxiNkeeecU2kqFh
Vc6LlpQIKbyZELa6hw8FRgS6Zn5EOzeAh0gahtbFA9oNIBuok7QMFaBMRc65bAxm
Mf7zFowA1PC4/SyYFBrfAwgFNqPaGf+bL2N2BHDAD6pEL++5D2CDZuUDkUPhGpwv
WQH5cs3fOOvlzoWNhJeC/a0ZuyE5lvWdfv29+XSo14TKe5/uy8LTVEDEPeI2n28L
nUTzlIhxO0T9LY5xjhOFIPraMonH/TIaxTQnux6AMRxbf52aXNCd8lj5iniKSoGC
UdMkuKmHlGSzpyxaBH7IB4GafDGRp+xuaddGhNqSiLWSkvlXdfQPaOVCi/BUMFY5
aOW90/hv05KFo+zcqn4AdFcbFsnoPu/++vQK9BBHKll/3EbLIgqnSz1U5nBqe7kx
HuS3zyRkFiulpJTeUZI5PSZKcOnt2s/hbOEVKQgu9lhdzHA2zk06ifQJU55yDQwP
Qk9Mbdwz0RaP3dFult+3xnYyudASplVcgp2T2G769OB5085dhCthHgnd2AAdu2gu
5G0J7ZV85oR7RA2uv9ukrGWiLYti8qkuqj0BQqxpPaXMQqh44BxF7I9KK4Nhd9vx
D0r6qAcjBAL2GZSvgieakDXVTJpPohNnMThBrgTL64YKlaLmSbN1IONdJO2wKEai
TMJCap31ZVeuN7xWRLQYwiel+GtLIgTDrI47lVmP8TNC7vab46xkq3Zh9b7zD0Y+
DBaL3bQrP9G6P68zUEOneMnJrsVSIZZuSjwZj+Dwlyi/6mInEr4VPt1KDlFdIZmN
wpEcofRKsgvlWxWDS3sWjq23QIypKtZjGDMfWTWptKUo0cr1rx3QbnTURODJ509O
x1tkbOwiXnbeavdQ+P1B1rH382M8DrspKxBUPumcy9gZFkv9aPCmO/tu6gGBl4/I
Vh46OKQLNt0Rwp4u3u/a/fGJuyXcpnfKHbXtDWpj9vt6/nB756fomarnZqUE6UXd
9xYh3aFBVJ2mRLN1Bp21oP+/li+iNWBs18MFxjAErM6H48vr06f2s7owlBgPuUIW
41wKZjEKALHyJKHMJ0saFQ3fRYi9Bbul0aZLYK9uMCKS62jN/gWPiG+qbU7VoY28
gwbmPxyzcry8pMr6ds05yw7p0jS6bL3qvaFez+pr65JATjOemkewI/sDLptRjy2e
p4inE87CASigxdjIV/O14SaBYowg72i7DzMezksRsUW7M+QfFFYmdVPkRBTDpCdx
FjP5qHXG+cYm+ltFPzTcZhC6Htf/fGdt6OZkPdv837EdnNFd/FkU0gEzy6ibboNB
M8HBpFNPVL4I0X3bQXEiIAjXTjVQKkpBJkf3JQdARuKicxQCelro8eARRtZoMXsz
xDaguhS16nLts12+5aBhZ2gFEfwkUN3vA6EIjyACbSba/RIQa2knv1pB9yOIRWc5
yzX3RVyslH0IhzpIj+FsazZREUB7CtSepQyDR9s9pXu4aZ4bfSV9eMTKEcxR+Ixa
YZudKb3EW68ob9isisThOSJdWgYZ7xxkwK4CwldAkrfkQE8CeOEQFdyA4FTtQUve
VCu34I3qM0jvxAFX8MVNY0jh6yuZT46LsId0+YLuPJZieI6Dx9/S8HiSVxqTOZuY
cb/ZBw1161WjgAK45jPA4Z3wDkq5H5gqxE2UOS5XVILvo3LmaDNvgZOggSHQtS83
5ARQ3FZ8QX4jxJtyxpm1SGWWgkEVQN9koSWY1BmIIPNFy4kztGBPD+fZTv+dh5lk
WWWUGxk2jyRzy/IWt+83B5Zr51CTCrJZXwYiH3LanDzOYlEa4HMiC3bs03YbiZJX
Dk64gjrFa62eIhG1b/8Wtlqf2BWYjL5kc7vu57p2GhrvsKAVHi2qh7BNXgGcI+kI
U4o+LePr0++spc5jJ7P5a2vRFGFc+PjmJ1OwvrpOsO2Bj27Dk1ktGQRoB548gV+m
zRK2Adu5RDDwqKVPe1gSl1nCaB5NG2PfcRoeDYOoLS4Ycf6Hk/HjYSHJ0dR0MdX3
L5i9kyi73147r5JbFtso+NuFHW9cl7cfpgNNhhNcXYqLy6LLYgH2x5rIXaEiDoW8
YfeQo9dQbTlSIXcYb8wouRwdXD9mqRsaMTT1k6bzFld2py47UiSAitioPv+fsM52
BnEZO2paFjX5Rc5e8z5DG8wzcSt4BLPvo8UhuVrZqgIidG5xZkegWv61Vv6GyKHv
rEmB/QkHEMUVl1oQEPdSlyJfrBjSYZdyLmn71qFPn7q5mOHHg9LTL0SeclguqRBK
VPEDKQECpfrwUMlg22I6ppo+flt2F4NmFyb7PP74vbbynlpvNAiW3sXHNpycDpp6
0I/Z+yW5/inMSFCj6PiPyDvY5/quNHjm3BiuddG9Q++q7OduTAXAFE8ZikXxKsW2
nMv7oxuWeGz8XfUCV7WyJzSEnJx7BamUHOEseoVX1OID/du/xscOMh5fKUpYrYhf
Yl40uW6JGeUadhNwoP8LXvXWZ+51kMlDeMAe5qx5YdzJBDSERs9OxKV0gMGmlKxR
W0WPmxw1Vwgq01FNpyc8YBVfwy3I66JblZ1gvdIQdNnBg3XjkAi9lH1ts76lMLSn
/G19LMUmZQZYjW3aqxP6b9wjLQ1KbY5P3defFr1Lxexsx43n9l+UmhiY59ckLMd1
2q4JTZUnU3+g3QTS/UdO8ZdIygpj2cELtUkM6s5yb3PBQqZP0MchBY7fGGOlL+DM
VXKLJZNtqLEUhhou9P3l7Qymoc/aLwwxH18TqW08QcTN3SvUJAVpmp8cJKF6XAeG
3CooTuHTf2VPIp0i/n4xiJieD2YHM/ftfQRCJEcTmtZF5RTsgsZM/u2n2qmg8To4
73xP1RqpK2Y0PC0ErHsS5kaOoibNrF33eSjzfz/2BMHpi1vmqMVfWu13dj3lyE98
k9twdjkNNxwhUHTOA+mLBi7dQLxdunOTJifTuEgga/mSM3q9cYmHUYkHhFM3+Jsh
aB06hlJAdoC1Fh24rwITI6EfAIx+oObBs9QUlUyUAvLsromQwTVmvkt/R/uC9BTr
MniplNQ/A8fiu/+pw1PCbTunEuMGUTN8GePSdp8d7h3SuzrzM2X0WNSyLMEbmoa5
XuLTm0f+rQ7QvXb0FrCikHKaplLtRr9qgNWiaZPLjlbxUTrugp1vnrCjlFPQn6KJ
0ahcg68qtDBv+aIgzrnfMuSOmXpvXZ16g4S2QwmgPhhbvifF5MNiChn3PsgIhWCM
JzpqL+gHKFmJKnz7ukTysr60huGVMHEYXhskLhahFP5xxnQ2u3EWotcESX0PBHy8
X/L8RzMhVdqX0NxHp99ptQlHvVKCgVHRU8byiYGzTbsH7n5Di3kuxSvIXKRN6F3l
SNlJ/XOmqeRGhVELipVqM28itsFUsFbAeyaJF2NHe5XDd6CMjkEJ5kP/Ly01Enc+
lCWis+t5lkzrMwbI/vvPIiDc74cj72JMGO1l8yVlzfz5RwVJRCwxvppCwON3WiQ6
iE63egMEdu9Hr24C50CVyZlKhXcSzVCcWhFCI6wEXVpWMwYE9JL1I8XwMbxJSKJ0
CTjShJwMOqQ/Tdf6l3iSqw6mXSHCMZK2Bz8Zfsaf24JsysUIn98tOzCiiT4tZS5A
K8If7d6rjRefNS8TFoAtzC4T+GzhF3lTjMkRJOCKcKYVhCEI7rww/OfwYJ0Cdq27
0i4iXnMk+mDFplIr5behj5W4aGpWYxoYf0SuMvLmcN4QqH3+0LliSEncS7veb8Js
lSZSUB08Ivfp32hKK7A2g12gGfAn2Dc0xQU8f7smCwL3PsRWbeCUUk3ConZo6agO
uTJfp6wdMASjlCY9VHo1ZuryuPTQGvJxVrlhf1+T09z6QOp+ZBetc5fZK9PF4hKy
RdrTFvC64XpSqzz0iq36AYa7gSlsEHcdCk4xMwntR+DkfFm2POYaCoiJuiuqqmxz
GAW4ofXInkSBorrqObh0bWt6xQKE3S5xwqqH1VXFqocKZD/R1f2pMxkJwRUu1Bv/
rz+1os3/gP0nZ1WpnG2HA1trUwQCtKUkytRAjVFjSJznPaxVjBAcSOR4MOjTgh1I
+kJ5XBTKDikio6Fgj+TMikvXNtsdOPQgkJpywXV2fNKAzTnIulpkQPEq5u0ST4MO
NUkrKWSefRXuaVxC+OSPO7rW8aOO8F1A51z+JwKDKTH92ZqoKk4eq7mMx/tjbaSI
0iZB0WUfWoOoQfs0RIosjNPZXr1lbGUKEoMxPgEg5pgTuZst2xec3PGuN/qx9tWn
fM6zYs+N6LYaW6aHSEycFag6m0vgfIW7R4hyYF8D8HoKZW1xmeMRUCiMGXJHf+VM
F6jG+fWMgJ15UXSdS3upZo5vW+OBk9s1aU5nJBYFYhfWyPfG5mKAXcvYq+3cHHdW
OgSrHO2K4Cn4R4WEv9x89ZqyzTiZ09eMMAG70e5xNMsAUwQDQg6lXNTUsaunHAbr
c7/+GtLddBKxWMC4a9yfh8J1vYJI41hVemoNBi3uK5i6T35fmFAZ2Xsfl9g1bDi1
rMQF+N++L8T3gGAkmM2IabE9gbg8+pJPzzjqgaRNoV+1n8+4Ms5UlyQtFFASrXcJ
3QbufYcE6ujRBL2t3s2fFJVXt1ffnuC0YjKx8gt/tDWMHdsIWH+XJ3b7No7UpfyM
VClQCV3cmzVQXyS+v8NE2Nyfqx2Q0O0+kE62blIK3mXtloxMSr7/X8nTmvhwp8Rq
i2TkrnRc4eFP4HQnHWQoYODrKYzGLYKQh6FnmpKGDNKywsAXEyr7Ik8Cfb70EkC/
0IRysXpTuAv6icrf8mYwYm/FXWglJPo3r0GY4LcZDa28q67V8nw5XMGnecIkGqSk
kx9K/ST87rHKVCui4lLmpAxp2jsR0vJnRzmVhqEGW+xVIOSgsU8FqEdYE/o0l4a2
1GjLVeoVs4eUQg+Chd5U0INEFRRKyBGlhddBTv3O+bSt1N/72cA6QGWjr40QdYSq
icd6QpKEGt5LVYZan/W3DxWBm3CQ8GIYH73E+QC5bq9WJ5uH7aS2oRraX0q6GCDS
Wrgq01T8BKin6l73QUyGuhHPi/GB1q5Q4Uv0nyAUJenEWhZrgOZo+4OGGRXG0kfI
sRon4yNz/ofXizwflouIWaPu3m4zpP6QL0Hp89Ui8EnekPpM5sLgCkpG0kNtv+NY
dOIe550ECjznDXpPIXn67cxWZlp9bgQ+uvVr5Fa0n41TCGy+ZLTPRPJ2sre6Z084
afqW6kIu1NokE2rvgot6BorgtUE2OLFgK+0QiLWjiSgS/EOiFhhq6aRpgdP3p9sz
GD8d7Rf1sSR1Qq3BU3FNovSyUx2sUJ1M39Co3EzPhNOeFX/WFZtLok6UXkRJ0dra
W0HietRduH/COXfz9uV7DhLpk8CX1V8CfrF9VZTcGPNEKzTL4vi0RBeUfShAsC48
tWCJkd8gJ0sZevMfSCVlkUFlvHeegRrRALbSX6twKhPwetChd0eolfiQu1jsU66R
juPKwYcYL5iHomqoJtuxr7vOgdHvVmTQSc9PI03SaWsY6dUecHu3feSgQXF03Ss9
/foGr8Z99WwizQBuRMo3KqsHj+7ykxgDSHNsD1PcIQYztgMvmrfriGsUIC2NwWiU
zI7BOUiZGBrLzyEZBDXqrObZsv4UYCxbp+rHtywnamfHJiTvEndVbxsLaMZXrNRO
fLHMX9C4XYchzGyPfqCjbPgT3zx2ZX9420YU+VNzmf7cHXvs1IcB23vpt3C53Jdx
LaoUBpXgxHzt4W3Y2mlrdLqMmMmlJEG2Jx4RdaiQodjEmxSA2Y5gV7JYwU5i9ngf
7PD+guIS9A8CQsv7AbJUoLWevm0b+yPN2Q7v51kpNetmit7wOp5P8lnfQR+vxWhb
aeVzvjG39b1OTXzS5aZvOIEwsbyuICUZLcVYLiJhvG89OKBdc1C5wONZAQ/6Yr1s
9GKJn6E06ckvhqBwVXgguMxVtQC23PxsCFQesUcx6AAn9ln1TsCS9ty50kCnpcVa
6e9T98SfE6xQefDsQzodjeD3LOXnEiTYIRX2aSOzmAuJameumHEfmfrB7//r6uHJ
KFjtfSzjoqTFtw8n8brGeK4gPA2WHB7Vc3Yyy26UaCTKMhP8io/At0+EiGmrAxOX
PPctpzKhDWAloQ2MIfvBfNNgcVzcjUoW7+QK5EMLvjuCa89OrqUkw1Gimihf5do6
ZWu97dVvqmTksm6DVGrNZjluEJ5xe1AN95vmiCKxeIAyhYgw6pxpHd16pl6MlCXZ
Kc3WPpIt+HrAB/leAi6Majm8O/DfGsOE4s6gae1Vv9+2phMjtCdUNai9EKKNPlaP
IQObZSrdh3uTM7Gm9Fe9Wzh81QCqdDV9VtE1518GV2HRQW5gukDTqDpqDqLUg3oE
+aM6JWTGW0e+1iTeuHB8ddqu1/69sp6PldYMeW2wcsLHgaE7vpgc2sXRFvY2HMAI
+pb+kuxhJ/3hPGCzalCYT709th0tqreR+ZJ+QoBUFXSnYtb9idDY+FhTIPfZh3y5
dcLusInFuppP+dYBFm7Ne1ZS7DXGyFvARTeX1ZtUdXAclSFH9/RObY9BTr9+enTE
vvt3tW8INsXpn/HZCOlvQ93LD5hTV6jkUEVugYPkOaLVsfihzbbh31Wt9m9sO8TN
4qS4fpT55JCwey07gKcEWp6Ek04JvcZUHF03nCh4a1/+2+rs1BZxmPEWdGJFRKSH
ur3pUQlYdcJ5890f1QAV1rnCWH2Id2wGW+M8cgpjMVh94m1oqg9YfhwxcuVE5WJM
Qj7P3YA5/l8mFOk2wkTspZJZE9P355DTmQVVwWmyb2+jTm4RuL9K5BFlLrbGXrXW
eI/n2FGJhjf+7H1UtMDmRn8/P7hrbQalvSYmYGXLzoVCne98hfHRtsbzYrghX95f
SglmkxQ6EYjPwuvijCLFvjkqSuR8aaSM+B6xoQoHy9GRleZaHFios6zZw5SGKlp2
quXk2DjeX3V9eY205RZtltdpZxuILhNZro9I+tV6C2s2Er88VKyLCPqpOaUz2ElE
tzg9ao3dSN1Pmx+0iBcMhJlcepa7rHjnBygXBZEEWK1n6c82ax8HmMWVtwVwQjRz
HojaR+iHH85uWoAgO2PKWjK8Tpaf/NZ+HrZ/ekZ4XPG6bbdPE63Blv+KlGh922Ck
a7zaPpJfxo7stcE2leDiBeNjXhQ9DKZG4C0mSeKS6qqRAGKsaqMY+PtDx3oOxXUq
v0J35mnFkiUlM+cw+9n0xVqdTrbUP5BIfdb7POA5ilLMN/tXqyA/lFeidMpVglzX
VDq2TLUWY1OkSzbwpZsJITxWvSAujnPfBNYupe/O/ttBnT4LI0c7rroQ2rSttJak
1YhfI10odpQJYhdbUA3h9b3qXCJAQP3S2HL01pPU0aHrjkNYQWIDJLB+Z2RWQcIj
KVLGxSG2W+ncTCAyLMHnV7jtBwh7JsDvhiTtg+8b7ZMyF9itkcjUBMPRO4k+VRSo
pPXc4mrxT6WY+A7+lSr5fNe4YbvVq/0KI1z8gxjVNF2AEYpoBRsfRSiWMJbKW+z+
/rjxTrugb7Dhmdo0+B8HMLiNP1gW4xpKoQzT412aINRcsj/VYkvzlfaaR6Qm5h6C
0BZB+JN6WyuXhlaJFttvpUkIHXhqHtqHczR3H2P7M+fVkRXY7HobLEZsae/NXXXE
KTs23wIR7alLHLYJ6/7xEzag9bpUrABKxjtPqv6YVwbmC5bX4/xxhixVNWjB5rFY
SobV2sbbwNIeQStboJ2utiRIuucDad6XKZWzFv1bojqQ+4s6wA2PhtiQbP0Hsgyf
2w+8Gz6PaIS5Q7vOD7rEjImg6H1zMyPgbibXZZMiQf9/unHWScPWH0jX1njUE7AP
F2qgBrltG4pKI07hQL9IZ5cPbdEziI51jxMr2GzlQXhi/xMErQXqE3XvjY9KO2Jh
+i6k5K6/Y2mBAo+CxtqtDh5aWqEGu5zy0Zac4twmniKY9BRhtoIFNfw6g6EpBMek
5G+InZt5RF2f3vS9QkUTc8eLdvH1uHEiVGAS+oPmLKZWObJdzYrCs9n6d3UJVUvw
SimL4sl1kmeMKtq7381/ifiRDXFclBS5JZwh/YU+4A1Ks4z7ecVDWLrU0iULdoc/
5gLsaReNC9PnH/zis49YNdF/5NaPsFeHMC4O3b1I9u1XJ8nRuO7LMRbtNtQFIvJt
c2aTDruHfm8OfpGrmcRcAXJczW2evYMhzyTXkJ30nkPzebcMuk5gFDwoW3AeRZVE
zW5Ynj1mFJmJHEmMbKgMO0QDbhiEYr61ek80hyjfo3ZtNoZK1LSgjJ2FVnsCpMjc
MnEsirw2BfR/n9/N9SJLmRyB7WJLUktjoUwP6At3lbkcOarMdtbMB2nQ2TG+Fp7c
GlIpXK1JYBDzjhnezXoE3IszHYiTheWfteVQNUmzcGlgOpi6jzFV7bjambTa7UuJ
kdRivmAThTblDAPp5nlmnTm6MDyM8eg1CVm0os+ZIQs8TTXzQjvCmPTIMEUXWYQA
YMIn7CPWrc3Ff4m5B9v59WODAGLwQdbBhgv8RwzU0f8PHbAFtbBklWlsCh4cAp3g
UZqMd39y7cZlMpT+0wEewGybQjU+tike/ndYVAe+CfdPwUpfyvh3SnIMNdiybqCc
6kQAr6pjSl8up0CFWsBIPACT44S93mDCp/wyxDA/84dxGWfGM5tcqxprOUvXEfOX
Hxa4sf07lv07F0NttSI5P/KhgDODtg2WXTEMLDalKyDJ9mcFTnoXlkQwH0gg1UGC
afkMFCMO9262v1LS5s/gumbZBgZ5HAE/QfSePm4WwR6Ef8WRS8hPlYpR1LVALYmy
eWiz3XexBDYqXDtZf0Og4UR0GJihriso3Mej/7IA3HxUUvWpwmNhKDNu4dw7udCB
ajMawh7hsb2J9bveV36+ZrVcTLJLaTuvrSAkfgow4BH55Lpdylb7GLazuOt5KRLW
rBr+DXEifsWkUrf3oeT5L2vXF39OeAiVR42Jgy99RVPwDIG30HYRA/mofFDb5uGz
VYW1MFZXvy9GRDgL/MvD0D9GQlGpTIw67MUjq8YfLHMdtTlkeDFF0y3Ut7kR7Uxh
1P4C8FDV5I+nxby2THsNroM+noKyoKin89nyJ46NXagNe/4gVC7L7qUCSI4clB8O
HXi6lBMdFZlF0dS9aCDaMMPoybLFXNry12Jlz+GS0Af/14y+CI5ijomKuvcTVc/K
2phQG/RLPUBxi6SL01FJuGhsJQliYK2PxJbOaW78bEbVYncGuGicYk5F/6HSanGY
OdiuE1JWbhcThkSrJlIRJCP5KMWN5zfMoFvdT9W6LqgXAKYZJ0nVO3Lu/dHfKDOr
6VJxjO63X95W1MfcKoRUU0HQDtx0g47/7+ilY+yaL26Vm7Fv9In6UQy1HyH2QmAR
HnVu5b8WMdlX+GlvvncFdoS0Zm22JFuDFdoZh2ZpuQSJW6UuwVMjYmAT9pm80O1m
jEgxXV8TF7B6sjoAm7jRp80nsZFpH5lqsI9tB408tAMbt6/g1CtuER9rmdZSZobU
GeGLzLZT5IdrByvpcVUT1CNMmtFF/ahY6p7Yx+rW8kPsiYQqRsCOincMLdn9D2UY
nzm2CI/kzV6x08TV0P7k134JFDfbJ18JGe2lDwvM4KhBGAkWgJZ0i1vz6rNcREtg
i3Xq6Kgjsk62uW+SWzkInfxMCJKNiOtSCx3O1/CVyQnnlEWijj6YeO5/G6lmiapM
6jDRmSSCtEvqi1AhNITXgLV+92OJwPiMQEPWSbzFO7OSDp7ll1kg4hQn4Hbe9ziq
PQ14KR0aOMN8fOaURk93pQ9srnkb92WcPemLq3Iyp464TqO/H5bzVvk0qtw9uoye
dJdynNMRcQ1swBVbqoiLllNlSUnVOjwGMqRClibOiqX0AxdjhcTVR/qNan74S8sr
BPPCz5l9PpZM6YRt3UO4kD5TTFQS6C7m8cZAmn35GXMno7sOA7LH49K3u0rilg1R
0tI8midJ5oFpR+4leamaYUcYizn77n+Hx9oG1UIWONvoJasVElUmIIv3ngE5WwUY
S8MShbOrB77vw7OogB2fG+rQqabMMQLfps4EbkPwZoAe8WZCjMXItD9DCxrFKfrM
WFoJnv5RLqJdQ0n6t3BtG/YbKVXtUxA0xunfqqjfYlRtF0VttmUFNdXzshrICaCF
oaiGUPTMxA/aZc6l2RwdevK4cf7YE/H9ULMCUqCj6uihRGUdzS16wtiRt4lTFWbv
5huaov2ORavK7u+HoWFR8ixuNd2qzoOaQGm4uNgiHVttfDP0nV4/0lWTrMBLNyF0
Zj34KETxHDRm2BFEYftIUva4MVb4mFjeId1yFPgwMBVLGxvLOSNRqhBaw8v/yONk
+/Jw3Lh+/bMQ8KK4FjSMpFokdvS0D8Yr62cknkacBHFVMvc9VGRTxczt3TDJ+wHc
85CsU5OCOOxZ6kGYgzELf6t1wDHPOVhon+y5ptUtXtlytVeplyuF0XXfCr29sjbN
kX2ZU6CJmynAUKBXUHowLBeq6yuQzsELJnYgEQCrQNa0PDAsRHcalDtMNmbqhVfc
51/edmnskzwXHcaeP3vwjfMwkFuMtGvIHKxW736lXQDDAjPlFqrf4UF+yQZ6Gn2R
adiPOHmllrHtf6FacNYOyXWITJR1booNcJEHzPM8Kguk9OcXT3L51RLNIH5pSp4d
b57bKHsOpX74Kad05libJaQkso6dqXYGmYkY2aOK0Czksm+BO2XnILBv8IU90PeV
Nsm1jkSd0ovX0HJ9i6g6t6dDIhb7P1XxCyXufDs/0geLN4ff0PczYoVF7FqUChqT
`protect END_PROTECTED
