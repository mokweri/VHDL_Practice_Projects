`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RCpPH7652139iRBPMz4AxS6XOVSWH6Q5ndBAdN3CKFG51eGecF4wP3f0uRaDEIYy
EeEm/4mKD5klB3dJAPUDUK+vlTljAVUm07ARyDYIChfVGKFJaShX0fmymWuLLfWL
dXjorcxrlC9lrIFPBrTq990YOzRJdCPMhVvX/DkVLCrHYMgNBNjg/XyuKY5wVnoq
lF/+LBlwBBAZwLQyAG+i3YWvFlBuGuIvJfFMgQJ8tb5kG0uRNnooIUfxJRutNBAu
PcIkq3OKhZNf0+8gkGVPXiNZKSuQ2QAC0MaKFQMIr6MAj2F8AVBdWrrp0Ho78MOe
dVmijGRiXN410nGAjvcJ9kKD/D+z9RdXCa/Yufc6ux2KErROAYgXSJL80N2GptHe
lGiJ+opE2FoNCfAO22B9zfjjXbE+aQfT1QfxThWbHD+nRU8lTJnLZomX5YzWtTo7
9AP6ViW29O0NjGaXyw7gK4lGccPQ5V1uGvvvTQkrXkbDroR/u/x2npzhK1s7sJC4
4tCC0cCesq8AGqwQy87mYsYu11t7JuXTNgqb6XSEQGsyC6KC/RK6tIHwAwhgNk7Y
sAKm4FikX1hPOHho/82pTE/ikVOthid+YzMCAaEb+eVumnOTYX/okxuHfbvYGoUz
QE5nWIHINg6vi3C20XSWiiZ6Gr4NKIEH7Rr6KbyZKAg=
`protect END_PROTECTED
