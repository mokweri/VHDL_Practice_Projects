`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6pgnJaTTFJwVN6yDsb7lzIcTHsclrp5SEMgsHIR/aWgBHWpneXnQEsHj3jcU29E
qmlo21ALHSrcyttLhYdqphWJJxX/ADd7M3P/F3jam3W+2JYv73CgN3/I7eBYfwKR
wcSxZN60DjTtC6wSKsQ3paYmsNJv7YZMVabN4pZszgFLmAfwGafyS/mNYeIkvBrc
o0lfvUryShVvqZ2g2YMSczpO14yfeH0MkxAGjA8bY3v2sk/iFL21MUz+qF3oojJM
npQwzMpY5OYoGEwTG8w5CVD0Xpu2jWLPYEedhbBWfAaEBShBXNgPi6TyKWBUtefI
7KCpdbIJ6ikwvevDfUDc0yHlzOLEBsqgFQJZ8xyLHXMBqR8bREvWaBo5cCKg7mZE
3Xgz79sx0R+cTSCVQOr9ho4QE9ySdhN3IGvMSlDewdEkPdZF9KzywVYYwZwRQrRy
vEh/81OYjnwpnJOnNB3mGvSftnj7N224qcHkKvutaUafZxD9oxtcsG1O5RXpP7Kg
KFhRr2qzO87z7KSy5Njz//wZadoQGaA/+qRPjS3HvCSAjMVu6QLTwvIvcJfSp1kW
BDNGX7ifpxCp7jUEyLXjwoFG++48eeU57xaRkD5gZxAXhqhKq5Y6OOLQ1TrP14e/
oHnTGHPeQhwSk3KFXIMi/9/9lyxGpgAqMzNGJxc0OQD/i1vSD4WE8cIwbTpwzE+I
qjG77d1OAog15Tim9qO3suerug9ina1m1ccL6TaqFszaAnKozK61EtpHneSChO2/
sUAlHOQ7cGxEixUy2oNJOhhVP+fkDUYOJ3dJNDADHvj3pQh2W6yHHmMzw8hhfsoy
7Yi+lbMCX+mbvkgXdMBj3keRSTI3CUlQT5TKKI9nQt320ry1U4pB6n8BXcTjO/6Q
z+nlpOsw3GrYQukmNUR2E17il8VxYpYS2WOBTvJGY10aOkAwac316qilNr8yx0Wb
qhECh5C1ChoP20jTSMO1MY3AvoJ5LkFQFURlVufbJAH1jkZSqhLDVbT9AqgP6Meq
Sdby5dIBb2ez8CYxGFgbw3/1QdKbdxTzo4vpl+UZ10YfJb9Y3v3ZicLMjdZ5TwMa
yt7RC2iK0zO7GXnLT5KaiDQybqAKFZF4bKsZ1QYpRCNEI86g7OPQ9gDWvKjE+fpL
R0qvmwe5h1eu6gwTkb66FaLuJqjFu1JkyBvrz9O0K0e/mJmNkRHi1t/9OWLqiIVZ
ae9/8juo2jXkAyTvlufm9t0OudPtEpsc1Vxs+rGLuvYqf3jZ9lo1ptJrNlAKuGRG
fEq7Exntc0+pBVLLBbXF3cFsvYxbJaAdtdJ+/LeVga41iz/BnqRTenTk6EVO56VM
6NizHnr1bLHHzbGFxe0RLWXDJ0W+UOuHH4jy/RC1whV0OSZ2JY/otp4gh65QerEt
aJhO73XXFpUzq8DoiiOGycrqEDPpfkjVtESSUaBBFysD9MIKNuW8F8E6khSBpL1W
n072O/oTG/0k/9TBKG1IyqBicyd1QFr/ZHop7UpO/sV+9h3DkcnWVdrdm73D9Kzq
+vJ8KfopCE+14fc7qmimNpXgM6eP1zNq1H0xvuBJpMRJ+P6bX43vhAAc6tFrPLKi
2JeAXW3wy+IArS11+Sz0urYnK/rEAm85flAw3idq8wVRe7jjRaqkHeN9284w7TNV
eq5ey+KenffX5kBqRS4LKcFG9pjMkDBjhlKyUz8iFxXhjrF1B1t70jJex2Jm1FXw
QfZ5DGe+v7tAu1hkjd/Vxu6HwPDAUAg815hCowsN2FhGv8HDXxqhWA03XEtKcUSA
biViZqHvxt7+y0oal7GjnWk76UGQGwlf+TJ7fU4pnVCeKom8aAZj48arUEw6M4az
LUKK5uaDnvgqViYHZtKGyMHqyjNebtae0YoBfOelOvr2pOERFqgLRHm8x69ALrVK
+t56ls2ZYz1ZqNXB4DHb0JNlO26l5jYVXYUa6xqTM9MYYE6EnossXYmUR/bZQeAv
0EeAw75sbbjDG9HjLwMmWCGNLgOcDQpncGddMTbqShgOIw2irZSXr3LlqCxGVpUq
Nb/ZtD+QJqirylHkwz0o9N3Z9c7d3ikJbpuqLBKWpORAmEqmv/5MDb+64kUns9pZ
m907yzyQjtWHZhZijqhRt7qcK1wEdvSOtbQO4LssnJMiYMrZjKt0eawh1zkC+yOl
hxDPdiRwIW3QpJeqnkleoi5O5Aqy4ButBZGmTNH+hzOsDtcmak8qkIQ8hSjhW7KR
k0Z0mPxFkjs6nEfGH4dXTS74Be92WWwwJ6RR3JlNvxjDgpSuBgxjMfp9s0mEiu21
REdmlB0kkT0mIcAgTetXxVFF2GFuuwNM+EMNO3JmNfRNeBXnw8z2db8rbQT7XJp1
`protect END_PROTECTED
