`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMtfp4OezLARjQDLal5TlorFmRCdDPJpWV3OutyFl8dqMbwPB5bs/9WtBk7CwJb1
QDvfwdlh9CvPa6PUIzdGkQojrUe490J9+FVQUKelTndZNNRRwnihYLIViWE6FDMn
Rkv8aL+rwxcfEjFaoWoeTSZeWrcL8u3kQZm8s/McJPpgZR6mI4cmGyHL5vBTX0Mx
XihewqYJKpBzcJu2F7PyZIlLBgKhiLPK0fjeYjlL3Xk73Yobnr5tXTAkiUcz3Fc8
LvO12RUnv/l1tAvnX4rQ4B0rvDNSHDmaI3paUlo26FWIrUr/mUAfb2FtlbXma6D3
m5mIGCtt/kK1KvWJO9y0CI6yMRP5PNJAecBiy1KT8FW+uQDDuNPG9R+dqZrYrnQF
Gs4G2jDh10LTut02R1aIoq/dqgZaS9S1/XmrBBhG/LmEdBd3243byq4N2Gi+3Ftp
jfcixzsiIVpqG69oNRB4kWmaE11sEssddh+fmCvGYMYhcwenmggR5QdUQRm6vG8G
nJKPvcCWYtt4+1S/BSuvewnPZWIyZeqZ5dR4KjejiVEhvpDS+TdnYfTBzKhY/gbx
xX5/K58H0yY8BT2AlEDqEfVn8RtZ2M6Vg22iKlRURfaukFMseOWZaRESYrJ6Nd3Y
5OfFMSgOdM5hXs/+Udwt+xxIfqJi/sEIC3rEt+Dmk9GTjsv4ren1QJ5cIo3DMZzi
jZRSPt/qRkyVSAsDHScA47wOlQ0XJgIQ6cqTtDe03pCGanw1N7BYqngC4ITQ43/J
S3yMPAW23AavffvcGbxMObS34cZj78rwigWLBbQJDkCanM+jcJvg1f3E+J+LaP/5
vZMp0tUUueROj9esdN3FIhpjl538zqa8iFxooa8gFI42XU+5cwVzydNqgXXHqI9g
JIeHJ6fT95VRx3JAxteRogSZSkAeAupDTmUYpkmi3axUfBAi6OxutF9zRpV8NRJr
4ksBHQRxPQRlo5egHdrWgQm6JuAEjODlTzJZWFcZt/QwGRg4yO5i9pWDn4Qmm6lS
e9X2NAOKeIT1KtCHLlY3IqJuTvM7QRupb1i53ZPibomx+MV39AcedwKURspH2YJ/
6V+AXqqTuwC+uxbC6OwOII2OMgWvAeKkLKe4zm/8NRAAoNDPhwtFqPVXgAVoEZac
l9zqy1uBMxFUJZ7iSXsjmaGfjvCQjgJcDgfYUgtyYfqvbt1EeEtjXyxKoZi22aW2
1pc1Xygu+a26taq2K811mJf+ls0n8mdEgGCdnlhpDXmb5Zqwkx3vR+r0HZB6MtbI
mmaobG3Jmjh/3oOFGBp0UivxLCdoomvDvYM9w5a0nQx5DU3O8TOEcGOfv6m8U7YE
5Ya1NIOaYpOzOO+jBDlwQHdlV86PDFxqW17bSeKmC0CK12m0v+SvozA76yDx6U64
DThUmFpTa7K0GlJi2AYHfUhwQzW4/mKjjBTFBRk42xc9FMKqAsGMjjEK/Tkc+FSW
ii8RJw7Qloso5D+aididwhVKGXlRZDKHw1F+rDRhcedWN51FcMflSG8qM/MD8hDR
0lAd3qE11j41wvEub41Km4Rxe4I+dJPtBtDChKDaP00y6dkK2yuHnuBsZgGtG6fk
U3mBhFpuspQPais+Bwa0Ek0/8WPIYl5Dv7aQtP96UkryFZM5o9J1hSEL/exN4764
KKjU16A2UCbxCP7qRnR0jXF+rqA7gRRDoyGO4NSNKNJmFbCWViMRYilVmLb6QxSp
vmKf+/Q5raH9ti59sTBUVRs5ZN3yxto060NsyKZTSfIjIgz54oILeXtqY7GzTPzY
wE3Jb8wtr+aZX1p37TZt9QYtCoHQkvj/BpLkTuxobhOhP8ZFbHV/6o9HGM/Jb1/s
qG2m8sHSkss/BmHsEhmnXqUFwPIpCJKdjwj3EiJkebhlNr8Uq+Ln3l/5PTPqrT2o
bNzgQoxNKeyWjGevpsaG9+bVCVuZzgGKR+PDb2d/e80h++9kNsxIxVJ3swiTRChY
2uDOLoWJzXses6Dj/AL4/JmNQUmW+v5CmCpd7cBD/WviTJBiyx9/2MMfvDDBu54L
BSTzl8YCBuve3tJ2AgrUhrKfhURoge4YOWwrFYuDuKZSDZci1g88gvng6soPivVz
wabqLMo+J6G7Ti9kDhHUAtn/VkKB1FF69s7csCgKVV3mLRRONCXkTeb9888z/a3K
gUN2a871dDAduZJQohwVf58rhNdEWjroDTQ6ybHpEgD7OCQ2fPqCH/a73bHxI0f4
NW1p3Kzf0LAuv8RNhHMzY/AN/Z49Pz8dzJYE3a83k8NNRSTtT76Vrvfv5W2qdwuW
K+F66IWxAbRe3HUKSKy1vkO0HM8XA4cEfE4Tp6BbJY3vnguyc/ky19UgTCnCiED8
bpX+Q/v7c0ZT6VCe3nJpxpdKsTkMm8DbBHxJ1NvBJCFvk0ZgR+OBtGZlkCTUDwye
Jqe1lvouORCtbg/Kmn8KooWegOstWeF285BB/HxF09SLb7YbA8iCEUGFvz8DnGWj
v+X0jKr1VHzO96QWKt8XhT9sgDo/w03Y3efsopoeIStadVCoI+eKlLuEYcc54Giu
mvwVzxPxIXjiKYIVKHhFl9vQEtw3vQTe4O72OeAb+Heid/Q58PvWx7V8OlN7cFqG
OI+grpe8+kgDE7xWq+tnhr3bD2UtfyTBlPey/RVB/Z+EG4ywpmMA9KbD6HFcthF5
+3n7Ctp8ABXVwGA2utM848PZ2/OwdnZKbV8C0g9NFKx/O//71yqw5IKYO1gzKgqi
Au549mHkN6IWvb70SPsu8aArMk4J8R9J2fJXi12NQUIMibh/GbPemvdrY7REXAur
8obFWC0lESEeXIHhJaYGGEU/UktnIHZwPEG2nclPYFJs7bSN0dhEHviwotDSUobp
w6OGkZgvzYtCbOVjs4Py/+0uQt0McDLNG5Lk2broSjvSpCbRlJ+dHflPtKiWLU6n
dxgDI3eu6QqICFD+16duCvTcAM7GIdz9iHeC80N8bREMIF7xui3ytsP8otcSR+qQ
rcIOsd6qd/JHjZojZbfzAuRtrkXGphC9UASqvXmYhOwgs2KQXeHSfHauQEfRTDZX
rXkRaor7GjBKMu00hLlvCuGgfTrZqly2M1LHjj5Xbbm1bIPcz3D5bnarFA5XsHWQ
4ERwLeqAM+RjTOQrywH4PcDeg3jWHqPVsitZ/AJD9PfzBTzD4UZnepcqOO1EQZdM
BnH4yxv0HjiWbV9VQ/JXC9Lv+mBItqIXzHypJTAuMsCHltvEN4OBgN2Wl5mKyACp
YUClZFpWfhUjw6c6dBVl8TKIJnQ8XiyOG5HI+U9E1Knnu6miHRrPN6DNs9yfP9D4
0MJwVUbT+nHyipWXncc6jrrQ8nF3HUb1ps9dG+iLLG1yaeb8+P4QFSEulsxOmLX4
Q9qzdn6myiuOATpNqt1UpbhreOBQKrLR9PL+4Mk2QYgNBIOjeinQUu/+WPSVEBvv
NkofQXa5qQuDU61bohUPwZjcY9Bfz2J3GuMN/KhKEeWo96ij2lUa6AllKaRxe4Gi
jM6WdSJNeUA4A20HLIFD/W6vqHqqo5OPJX7qnp86Us8bn17U6yNB5rT7MExGHfIg
rnjn51zkwS1UfBn1jBD7KSEtltiAmDhClCoKZg7BPs3Ttx9vjnmXl3Yzx+JX4NL4
f1+H47d9KXzVyJvcIRe+ZSDlIeBIaQ8P1S1KeqwEGwC8fE30EzErNyzlUmGFX210
fGxc7yctGidq3JDeyuB9VxxzJkpJJsp+G+XIODGKGp+2ySRUVg70B4xhnSuWJ/FL
orabmdltnqeglxlVQBaiRyXjRKJHpF/Xwjq0ANZmWFOqvleWz1IyfM9d8fB5P5a6
gecJeXYf+RX/CioBHg9dTHT3aygKLib7sO0RM7a/MgpXYEjLgeU9LAy3laBHHUHm
Utted7F2Y+Ou1fTkGgYhGUnxM/qmQUb3QVsbyIYO/O7oUOwOWRuJGjRB/Vmtcj3J
uYNLih898bxd2H03Clxmq2b9BQA4F/gydVy9JPnMzwpTMNhy4pR5TUobuNhDipB4
yfbJQYJD59CTHNp1pCnpJf+JJJPFMlFm+tNgA4FPxVO0kAAuoKayp6FTo4XmU6Uk
USw4PRzT51MvBRSBAdFr3yG/lAA4/e7xweOUEayulHQ1xhsecUjzUUJo19+J30V2
pUND1AaXse83FFh9jbl8Ne2F4YLTxfj/MTv1qQ5lcSITLXmmYWBflIEsVaf0SZPC
XnTV6vT19RHRyF3fY4Bphv6aurufrTUEigqh2UM0Zw7DqjTQAvIHELCeAaE4iyOi
6EijwRFGZWxomikuaqsVDnFf9A0byP48lYn9MYxnbXr4S+faniGJ0QmdPUIA8F+u
UJRldKEPfeB1PokXSRmiJBkzz0mSM3S6hN+hkPiPtPi4RuG2baGYugppYN3BXz1k
ygfPAJIHrs7RtbCmobH3HOWWz8/KM+/n1YfvIpkYfqsLZ4/olw1djb0OKaa7dA1W
YNtbY5CewEEFVkErVm9f3+uNbZHId6s307fB4GEzG4dphRVDk1mzyxVHFw6Oe1Sx
UlPMU6JtFgA4/Yy9tUXS4bZcggAAL1jIDyoTtr2BoTze6vmqbJMPv4a1zn2qhPqx
UMmWPbmYcE0eYk3zwPk9ooAsJWjv6k/Sw4T/LZSD+6AynKHwTeuFhUKhfo1C171J
JgiWum4qqqNsEriH4Tg7zlW8hKv8M7dN2QVmF+cOK0zxTkzndzsL9G9vqxMeoXU7
BYpU2sjVcF6F17zPV7lL04f/f277tV4UdRmI3+JNl4aTJSI+dJGqsw/xN0p4seI4
j2e+43B1aR0e5NuHuG6HxQaIrCy/+5ShVx63DiyA3ngJlRuQjnxr8oGNNE0tT2OK
5WBLsIuJP8xeRZfdxu3KXv08s/mk2qYHtWKBZL05gX/iTiex8Laiy7AwuU1Anjcd
3toqktlH97w7IHFw9p3XnfegE64noiAwRN3trDukjWpW+JHECaRxBPP1e1eymlt7
7xT3T8ysQCfj9PjaDmvJdo1WuyW8ledXuyBDx7myQ8yo+kivo8Y1es1aC9dbaZKC
oaCnEzXEOdXH6zOSp++OHiaAuFqmdku+NkeM7dnS92FkbLJwFHLOzRBu2WhL/EIH
wPLfLO2yzzGTiEQjxqSUrKPG8XmkD1ucsHmZ/z49SknbfcUAyre+D5erfkllcxdi
B4/k3ai1Wf+t0bb8OYVxtH4ubfGwf4iFhuvYWeeX5HVYcAx0J8LuZ2YbF42vjK6J
dQZkYIC14chny9UbiyCSqeJTeYBka6GuOqHwui61bhdaImjsug7IRhcze61R59ZT
XTo12idAo5crP0O6KYLX0K0x+8wEiboB4vY1Ov1M21kZ9QoYyQs6J9UmiIn5OhiC
km6EJhjfbuA3mff1bP7T3CN7c6m27SvZF3sr18eur2UjhapcZeTyYIRLvkirrMuO
fxmWVSAWHl457wLWuqcI1kYYNfoP24eW1iOaSZ6yV+IHZ0gm7oTi7zfNEfz39rI1
0iwGD5mye2xuOxAFkS8rSFqUoIB9/ZoduatSbJvKR/8+jL7AAh7FWk+qiOhI3ehu
VGcR5B2FWNo8fCAWbaej7tQe/L4wt/j+W0XOzZpTDiCIFuK0JbZHsDITxJSNt9hx
4bjtilC5O0e99dRGx4b8HG0n0m7ErRHFzXpSISMrJs8GB33W9GzAytcSU2FCsshR
7aKvZfYVGtTzp3vGjsEkbajVrF5Cyqt4aSdbEH74cViNkMAT2tuR3wizTugJq2AH
fohwTMmlrTte6pPa/Tw9ZqJdiNeTpztpFJ/f5Nsjp59Bx203ne+NhWfVm5xjwsqe
bhJsmbJfG1dDmOTexRTC3nOKXXod8Qrir9G6L7KCkAqpIpr+41ikN/+LnWxyXm7m
FkUY5BXoAGmh/J6Qtdgxbj4tnnRmQ/A2iFtR1PDufMrE3nS3JJlA4nkFrONHdFR3
3WT23nHiC5AvRsoWwd1o9/e/r9WzrJSjVav7H6ondaLljk7AobxTguskLkxE6UFy
Wfv7YZ3ePwgcxGL8qgf70iGMXfxysyfhA4r7pNmRxHx1FZFW0ullQ3qR+EyJdt8M
88AfL+h5tocRgbwnt6aEeSCKGe1TYlVrO+BPWwxvz0jrZvhdaPoWaveubKBR1zco
woZj6qh3z2nRRz+MA1fPToW5yDcl+2zYC/lOA/gOArreViHa/pHOrRIo7Vt9ZpeN
1LC1gU5TmdmEMoUC2X4G8wyQLHOOTaatzZAjua9VjdEOle5zV4f0bQLRImh6fBxT
yG5/cpchOnHmzl/kjpaEH7pE9PQaexZQrtNZhHD6o6sxITLhl/3f1G+gR0wAC4wG
emcCWay/6WqSyUgY2byV+XQK4t4Rm3sy5Aiygj8zA772iruf5ffPvOCxMTlkUzQ8
yDolBGgVayXRE5uK9gsIITSUuXzGO0AB1VBBW91U9tIJoPbuNpWma+w5XJGlzG50
ldU+WBugBoEh664Y26mh/8bKh/JysI/+C4H5HIb84EVbz6FNj1CzLkISnXOmSBBc
8ormKwmm37j1We/RpXhxLJmVDM2liWvzbaGnMR/3itMKWdc4ztreKc9+ZWH4MZ6N
JYevSyD2g94jo+hKnJqGQk9LyAIfYrhptSqAH+Dx9M3wKqGPNDjgD/r0jVMlSwFW
ziTtUQWLhuxrZPEYCD8SEt9oSz1YBzEETG0SnuEupfHW7Dy2Lcph+4oTQTR8HycC
X5mq8X+FUsheDwBxWPIxbEZoO54CqADIhufAttYB+uQSgp456RxQaTpgCYfTAgc1
nAdhlA+KSOA98mGbMlgRgacnwcA6Q9HBxNFEd/H+p875yvTbl0mxFmGjv5qf/EEC
5JyKeQAXK5CISfDzhWCBf2Edae+j/kSmuAKMt4RIWBDJraAfuiPtYu2SJ9ed/Kl7
3KjgfcHRY1Dhkt/G08F4O1P8BL9HKMcjhQdizfjNgeXeLGCFJ/PQdrl2jc/Zyjg6
BeW1Ra/PGrRhhkdqWFb6eZgrvD4xBcMnwh5K6aAsrtKqxa52zu5uGYMwO9pOEJ96
eoqteIuFPqcPSdI9WX9e5sJe3JcYr+R6AIsvDQdGHaWJt4zBzFa3Y9Niq+0pBw4c
M3WoMMFzhCwCibn4crDFO/3KcD4h7hu0MlLwx2Mqg81mhQgpaSQpTerrBdo99E4X
MsirQLjHYNGbp2IFOXevx7OE+B5NldeqxsQln6OFAWhWwIX3tuh4Pg60boYmQaKp
jgh0us/EJjqwzywW86ID520qVZ/Bq0bivnzVlg0I3DtB4qyyPYj2IrL/jzXH4q7A
/b43KD4Yu2gq4p8Avy6LEa2Z0+pLggaswWXmqlnvE4ND+4rQmGXcHI2XnD+Lq/iY
HZkF1kJjM1qfTTYTuRMZ16Ll5WBTFaNTBekfMAb2PLZiNBGgZ8A7Z9HC/z25HBof
3dNOW0TQ9c2RgyUy00VGy2WDUnRscbdVJSB7WasmSCypR6Dh8tqIw7gom1H1w+3W
UnSbxCTaDTt0K1+4aW9XYQxwnQQHcaQPN404Sy21lox9D6pQ72p/r6ocfT49bRWI
YIuubpmK1I2fXmCdzETe4jED3spy8xDXlu58QcwTs2L1V0qATWhtGkSaao8hUvPN
Hhmtm/CrM0XLxIHABrGSjWFhAX+gY7DtDP1mBq6kOE3noF+BI4MzhHR5lqo3l+Zv
+Ssq18JVANLW4kMSUC2muRoz4TP6SM94fb+afz2M8V7FGyAmhrQidtcue1GZrUdM
lywWH7pf2W/wDy2QEE0uhQIJcp8dd+ODHxLESVG/aW9qnL5vhTRehPRAvtnORSIX
1A68qIw1t0MVTV7x6lTKcPTs+cx/lW47LMBOUu1iwDI2YSNaJtHb3Pij6Tc4EX14
nrp3gcNyoMVUzLJC1HatVgkljY7KUfkTrog/QAKs8GTUK25U1Mq0MYSQHdd4y/ws
eqyNyF5uNZpbqyWWvNsT5nkEwfKF41iVvjNgC9TI8Xdmw+8rY6FTOnUyQFMLMVPL
AZ/MDqzm96YbKUdK1wMIMntAcGpP6cn3m4Bo3PG/eDmqo9JhkJuWfqDEASwstSrS
KSgtb0xyxrsHYQN+mOhf08Gsak8ToJnpsFqL6a9iRwthXk2d1MYLC86moa3D4ygs
yrJPlMVhhRuJ6iwxBH5+xqk7+4iBJ084uxlzX+qsOJx5ETt+UxOxw9tKQ7kQvR37
bYleDJa8u4VnDSpfAuh8wBPLlhBc2BLP+gxdkDqtD5EyYH1i7hIugI5IGjgE0LQJ
L0cvGlq9LNtDSEMHRo4+6LsMmq4ZtBnIZDZI2PhgJXs40m+3fRWSHgEZ7zsz54F+
sHSl5chl7uv9sFjHRECe2AuL5SM+clFMbjYpp1avxkN34x25wL51Tj7y29nNJQ63
BpaIVo94GOVG++3xEIj/DJb+SnhdxAkJPAyj95upubX4geG28ljEqSLtfA1HyCnk
pr10NvTMnhEVvkltgNLe1DrDtkp72UUU+Kb8VyYu5HPaH0mFNLCWX9v9+BkW7mLr
tz4b9e8DhSZFJE5AKixwM5aO9ChsoZOdLCsCfCNxTfBH/f9Zd4YEXfYuWuQffNwT
CKmFeqRAdegXUbQk4FAsVAxePkDBbk+CmQfE0YQTbFcCxmQ/HgZO5drw9zPaoXku
bKHozqP5iu5RC2LJBWi4u5OHoNMA9fJw6gzK63/qaKyW+M2skVF76JEDSvDEpl59
5NapYPGfeqNY+CyD64H1qBIcYcTFXR0ZDnoBAzmaZQAgqpqALutfpxcbgIWkDLU+
aVKyPf6JJzcgvWwwUD1BunZJVigMPYHdDM3U4dcYIBwtvoAwC5raJ7utLCGtDUM4
LSHO4Dd/UavTBjHLkOTDTc1kEtm/23O6mcWWAzlNhc6UgXrRDmiOBOIE2mYHefl1
nrY8z0TQ1efnq9AhaRarVIFesHGghORwO7wRiXMInhSyP7zY6TS8BzYREFsj2ahj
tRUboTkJ8xQ0d8WBPJdOh8Up/rDRPYLM+ncWiQYUKIP2ziOHJTdoegoJAR4ESntf
xn57gdncd89kUyVyhiHVDwiqHYJINuVapRekjGD1ezt5AsqozmhadJ/wOWZDWngw
so1dCZCufZQip06Pz+Eljb3GK0xrR3rfpNuupfOdg1V55hmyphtoWul4RKolSJjC
dhPYvdYdqREVvS+qyTgFxj/j8RTUe+FfImjbgh9khHhLc4KMGhCEQTkb7qTH2LlH
3eHzyKL8Kqjk1dLpFWfXV7oP4S3/OPeMQNIV53YqFB1gOS6ZhGSsETGbbgz74o6N
UX1/yhlHybau9SjkfBBebwFjhjnKA9r1F6Kwo2Qns5ytsSunV14g2fYuAuePDujS
riY9f3CQmTw8XOm9+pPUM/CJ5aryaGfGEnRPha9XV7b1BgaaICv1uNxojMjrOjgR
`protect END_PROTECTED
