`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khKbY75OW/yvqFFkjgDhNrZWlXzYs+h7zMC3t/0UEjFYgu4vnS8z3gAR7Teg9bOh
Vl5nCQIol26Q3nUlm06n2+Tt+IItJhbiihgzXWPxsa1aeOxCR/DnjLEg9qQC8BkN
Sz4itMT8Jfwi/2twVao007xrk1uP76d2Rmb2670vPmC9GVtMIlGz2P81dimeR1f9
WuGke04vpKkAS7zwLhhfiUBg53rViIxBVUyOAo9sdggtpELde6qiUZJQ5Yh+oZsf
K7XnHvUuTA6fP6Ywrctkuci7W1CoS04vNQrB5Qm48VbL8D/P13jPknQevBiKoY0P
lan23oB7oFgW0jTsnrFIvZYxjdnBVJMnJT93WzFmIj2xny7FXXDAGEpVQExUc7XV
vh4EEc55b2jDa47xX36/pM8cB9z3P4WsmlRCOP83tb6GirZWTXXDpykuAbQxCmoO
rNBGDxuNjPucnLHUepUe4Lr0pA40/d7dVlzveBO5bpB4Hz2lfh2lGArG+owRJK14
L52X31D76AKTu2tG/EReC0VYShQ0dU/+m1ljZ2KH0O37UzBMIa8s3BWHAMnWr9gz
S4maqqGSAqv/L8lNX2KInIEPL+B4J1s4r99VQSbxZjzZaRINgVIBiBoEjF/TF79s
IF8jhL8SGS7YjZSKgiq1yUssuVoUlm1eM2duHK+hX9Hjzm8ubKJRBl8S3qTROo9G
KPzc7sCYKDgVAElbAbltg5HH0WDuPZyIGVEQThk3j5Zu1kbBIOFyHkkvY1FARon/
9LHbEZgEqp8UuVynzkNW5017+OXgmxvXH0oKPgSXZu/bBuP2nT7WtXnwfIQkHYjc
UAb9L3GY60upWoAmZXC46ldgHvkV14QuKHmK/Ex1erQ4AgxbrejThJbuWG1tPyj/
L+Yv56lOZhFNutaI8c9hzLVj6TMM4Gccpki3Hgjl0C+yIPS21ZtstR6iLiIY1nyM
tu9ieI92k3qTF74KVTN9mz51UtvDBiGQNzx9vYr2O7SKFJO56Eo26Y8hAOoAfw4H
23BUp4jMQv0MgY3YwQT79xiov+2zr5snviWsrDNgtcVW8xJzibkZrVhk5Ydvr7Bb
Umz4ycWsgZb4rvIkNcoaF5tJZIS0WX/klqL5ig12XUZhvWLcAwsuqnnY1nZuQsP0
WB6WufFhjAqRpSbOCP/3nRYwyrBsF5K4Yo+D5iHr83y70MwMg+lYxxDOeXAc+2r+
GGiwuEbcQSNtvKNpnKer/x8GkzCxe0FBG2Iv45QM2gwA7GU0VXKeY/qGhKohNHBA
XqJbbZoT01xSD2Bq3pL+LTKOGP3jcGVti1yeZ5CQdSaBUWxUTe4nmiMiBoaD6rZr
kmHmgoYAQnN/eD5HiczGTFxmLJfsOKxpT68/cLG+x5yMgUSi9E0UwQu4W2+7V8HI
OkseSYTOhesFDhp+4rb513UGDZJ2b+LaTNSWc0nVxMbrauC1r26r/YjfMdmgbm6u
wgQP88vCfjLekWK59pa8UPcx21T11yOKjK8ly6vkhJ7Ce/CPJU+shRToWAJR7GNU
mqnWgiYG2nmTTKxa8AUbc7EEok9T3pJ3EYv80FzjZQoOz9lAy1UlXIhny6zhLZee
KcUdlldVXGODFeDgkIIxr8JiXVQX0p3M5tjgBVq5OxKqUCFpdh9BLiw0zPlSGLhy
TFucdn+cB2LQ/8wBWPbI2G3FbJrrbO32zTic5BnHCsshyhmmFbY7aeVJsLThh5K8
C/Oco0Bpb9gO/KmQTX2HiHUGZbDPs7VFyzpLtTRf+4KGwcAIHv9jXfj7s1Kbm7Yw
M51Yl/3vUSHSCwlSX78i/fqAFQdIV4zGby+nrPEyQpJ/RJtTQHOPN4ja2zUlaKn6
iLko3oavLot74yUztvB0h9VLTB8SnvF2oYXp721bTsLwqrT1WAoddIK11EvRJymY
tdayISs+ra9ERFnRqCnRC3pnNJEUGCZCpMy85124EEQ8huDmM7ESufbnR9VSxXGH
8aMGWqwnWR5hwTrlrHGYsOMbpwBH3OXoWNsNZOBwNaDORZgMlZBpr8OVYQSXbPcr
yYfxl0CUQa3GjtdR+ziuqsdRyLmcKKNe7mCBF7gXz5PDgwLe6H6GjdthcBWT8tTE
poCqgR4Bc39WOJLsMI/mQD6wHHtF4RpubW3K6iV4kexe0+PuqFfH982lLsOhBn23
wChXAEt439La/rEcosWMiJf+TNgEMEu9TiSagCef2oPVAjJMGM9nEgZzRSllY5gK
chQk3odSZyHWC/J2aqtfeSD3yY3VJFuodPVccei3KhdoRYkKqWRTLyhyNZukj1BR
RAG9+2z6FkiNIz9BWnFYW75go6P+UMMnu8FrP2YSBeJky8DvKC/sprOx2bk/qdnc
0yaoTWRc45ZfKCya5V9WHPbcpkBp1snbHyPPXmCU58SQg2jrUbfdysMsMKE3Unk/
LNO6f9HBk8qrLi46ixnzEzYRDcewgVX4hfAnjNQujIbWVKP2HhUDx3aLyAe8qA6f
ASOV+im9AvFQ64ydZdmDBm/ur7YHFTQE7NjFVTV2WfQDbmf2S3qOSko/j05XRM/m
3JGGhYRdAxKrf4/Gs3Ko9PiQkIy1ROLySNoqGUJHkAi8BRkiXMIs5gSV07ZJrG6i
qTfms2HFM/7yjTjHdQrvIcElWeip44wQpv/bnStdB9rhfaAW9S1+rQT3IW0SKxkN
7/yrIATVNnR2moS0u3wuFk80ELMM8BUhZpc0QY/l5WMU1zp4S2TW2xHQmhF9tJao
KT0bsMeOW7xr3cNmgglvbpqr31aCaTqNBQ2wviy79nRLs3Jh5v3DBc62xLtkp8aM
1NmkU6L3/dvzvZoezL1IbUqtKEm5PxX9maBY9X9wPeNycP6h4bDAnhfsGA3DR113
WZE5u5C3SAEx/gYdKrnULgVSOwXr/T5V+glwtmXoIfzS+IaI51LCPnenpnbDcyD6
racpQQjJweTJUSobAF4TPQMhEk+K3sRt2uEvvChj8wpH8ewaNPoG06yel9jsSs0v
`protect END_PROTECTED
