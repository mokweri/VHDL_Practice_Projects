`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1MZexvFsVtpMSgodqjg5JGRn8LL1cnvq8Q03r1rgvM7LzlS7v1ize7mcsthNeZ+
qmG4aqbEx7yvbsdZF7qVBdqCU3hHvayKfP7AhuhdI3QsI6aTHDsYw5/zWXf3HYm3
2KBPS6xmcNBVqsKdDfUQj8mnIxE59gF8qzmGsbfhlRMwnMPgJvF8ul9tcp6dwXEt
zYbmDeXRFMCtAi08P/fGBvTwoyXCecLP9WsEjpTVrcTFwe3SMNix2yXKI4Y6B6Xe
MduP1L2fuuVOQnw0jm0TxbCTMLaqhlLJKnUwPshNvjIFkA4A4O/lT9JqdzDiBfDO
7LGaqvgSvSYVb18tsSqu8scwYDuUIw/zaBZv6cWfXJYKSv4duft0z2fzsTJNBe4z
l2YXKj+SwaibDnysIxKHPBboBqoR9A77sq+qp2ioiA+6vNuTBT/RHdzr4Lqc4HAm
3UnY+FvbU9kaG8OqhOba4c4EXzbloWJ+3GrUdlSC+oqDXEThDBKM/u+u529DqaR0
XOGyRtW4+fWlR+wQc9urfjvYicTg4wFl0NdIFUPChs8=
`protect END_PROTECTED
