`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DOidtcYfOpDp7YbTBmN+WucLaEU7j/N0suDh8ZuzhPhetkKq6CwjfgYmO7NxigF9
5wdSX1JtVcLIsDxKlWrN50tGEDxDBBOgK+bhO+C8/2SHNhlQhu56udrI3+shgmez
KUGujdx1PB63w3w54wTZA2tfaXlRdbzu7e1/Ac/vEnIczLUnZcuetA65AumHSwgA
BQ0uBZQfsQu7XpYSWiBhrqI2UZH4NH28gVoi8MAfLCPQchKYL3isydwfngU7OJwg
iSDuk5eqTymqDe0JDPx98rJnvXoIPDukO5/AWLdyLTQQUmXEjJQxy0oBvKoYbUFs
+GLihwYuYRwOSqwDyqauL8kY7ETKMRe0Ti5UtJBOzbMAV+COriGWQs/k5HRVPZKJ
ATQnLhJuovtSIk9RdysMK0gvEd+hpCD8Z7WG/1rONppxEWuBDCKdjAVnbUjpEVqA
eRVJsjKbLojNGz9wAjdBNw==
`protect END_PROTECTED
