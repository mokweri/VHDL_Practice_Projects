`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWR33cwPGJJ0ShOjtC0vXOtPZdKi1NpPjbZPk/NeegZ4HA4Rk1tXuO8KsksshXh2
duQlDjzRIYgB6wNOeXLAYlJwQ+7ivdtbSp2GhXfMKCokYVTUwgk8FxziqaldnoC1
RuZSs0KkVIzkcsur2ah3mXGX7LmR/c4kpNlzx7J5fii8oBRoVOT1oR21jWeMYOJu
2CTvQEONp28G8JQxsDENyxldPrf2gOixnzITR6DC9/HHzAh6/c5A6WufhG7yDvwc
NrfHxgADVJRlcepDwkBroPscz8PZ4f9as6/NIbQqxpLt9zHvkAQSGFFSzFpSPX4L
iqLReu1slGcbaI+JroZAG2eR/EKGAFyvcrGdz79Ej0CTgjQLvbju2FSkoHeZ23/t
Kwjqosw6v9OCqgdMRJblZEU4bb/4yXybTjiPMR6Ok2o7QcsnOwEBo3/yAVfJF/BF
1+dU5eBT2ODavr4Eo0cRRx2I//rf+KE8eUDt4D2p+DZfCchv+XL3BJHeiDUjlgT6
`protect END_PROTECTED
