`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSPLipwNfyyjb99KbtVIc0P39iyjteOUPPnM49p80E9E2PjJlDsst/FsPswr6fep
r672G/3q12wy6Gi5Palkz8TdoxOQ9OXvhsArKUIBjUZkfpGcJU7KH0rKsUxLAQds
sgzjfzdc6i8UBWIxp6An65n+eFUn6pYolawy2n7Df5tAjXONYk7qHL2NGXFyJwQp
DBAzwen7WdRaxzBYX4dJD1SHTyO29L1G+QctSans65WTdhTQ9kDNFO1xOtfW3FXJ
ucqVtAJJ1e0Ufktvrp/QUZ06crgn2sHT0RIUvM+unDXexJUuprZQ0gEbTFBql7pS
81f2eZBuzMfSSZ4Fdj+MURoJIZnhDDYeX9/ROSHxJtTjVd5uMkObNlZ5/fHPKbrV
78Kpm+E5mrVvSV0NaWOfClNgNt5Rla3xSVfXvL8AjKzyLAtuOl1nDRGtv23lTdar
qovhI+cTODO+qyESuieKW61W0+JRYq6tPHm1zmZUWoHsiioq4gDYZP8zy/wirF67
epPMdtB7DzL6YrRmQYgkB82BkTaRslq+0UTWP9F2R2qQpJSNEl7jVUXrWwJuK6VL
t84qjD1GOA//m5asEVLpVNYFZcIx0ZyvjcLHn8WO+8wqxo/gVMNHXAiMfrjZO8ap
MA283+WfX/M3V4aIE9X4VmBIB3VukfJwm0Fb/skbF3n6YOo+yIxPipecn1X+xYnM
nHAk3HS6vzgUvst0kIv9W+WMWNeeqU4u/v2+c+JUnNy0r6w7ru1jzX80zxTWFtFY
qEjdlN34B2DK6BzxjtDtFOiUl0NA2wqSUOEFNfJytCk4gDLQZF6fnPIXk8XnHRu9
/FBr4Sd6BM5YWoA4vMGBp2fWTDaaBeAaTSMf5g/pk7gJEIG0GGfIB9lClx7gjaOX
F4cZDL9ehV5qj9ARF65bkch/bkVDhjQGRQiMjNsXnmSy3YzTzHtrTrgz5g8XRKTK
G0V3746FApb2N7lrulWRmKk3/YLLLsB50/rg2qukL1F6eVH2MbKSwG2AfMW6van9
DaTRdjRwGrVkI1Lbt3mB/6oiC0zxBVyeY4KEKNgMlHbFPX2Wvzt8GJbTTU533Yol
`protect END_PROTECTED
