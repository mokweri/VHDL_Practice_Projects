`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ea4EfglIEYe0AaPkMI/0RuuKqIndwTfVCdlSlxFB9LY6OhswYaz4F8j/xBvZDYFk
AMbkwaaOjv0xia03kywyf0MicrK6iwRs3P+hEf8Vs+S8JfGi6trDBSIs7lMSmUJl
6Zu7uQNlWeiiVxGE5JzEPZV10qxKL6lHvQuS8MMN3+c6RQp5n1NQ4RUTSLRWfxpT
20vbWvJ5HAx4u/My1YO4RzLD0272w/gUpcor8mjfyLVltuEXfF4dAStAPc5aJll7
IpDwifk8pLxZpydMcjOpki+SDjmWBsoSBSShcJTofBNhHVbRVxBUfBKqEdYgjGx1
QjgMiN34PHFPPfQdYw7/HtZgSp4SGwkXmYs0sky5vx1TvTRv/i3P0ppSGv6vXy8J
DsST6PP9qtJgok/cDAllmLGuYoBspl9/KtQa6uH95MS52/+Hx13odbggMTUAPtf4
jHmLi/gwXmAgv3rondwvDRDmxsLSOlzs5OoieSkj/ae/YvxlDxqW4ENE/hJ8387u
21kmS+lYSZwi1UecDbT3PEqhtD73Rqom3wu65nEM47zVUS++vogpDp3PRVpxLCO/
rGg/iQjzDCBC1KO3zc6GWhhcFp3cP7BYFLgbG8Vz4MSDHbByHnZ9l8AdrvFYCrCG
nj8TaFJbpOOhxT2GBsR4usvSWcNmHw8/UOHIQnCLg55Gsbmw8ON3PTy5qzuWrnLy
BzAg6xup8jw6RmSVghc18A6izlb1v6WILkwu5r8HAXRejg34u2pmvvHbS+ruR8JW
nfN4oQYLht78XjsF4HoM2agr2L1HjsuSMoUGFduHJ1pc/YQF5khiLUetfV2Fb1En
`protect END_PROTECTED
