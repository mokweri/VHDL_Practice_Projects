`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ju4nkQsZ1rNVEMkpFAReevo3/8GYS+cSpIG0+cYhLZt75BK8ZHu8nT3XgH5om9Q3
1RzHh6wQ4mldxPw5PVa5oGxko7PaoEel9Z5wTnlVR5xQ2N5vpyU/Q5ixW9I9467h
okNv+7eneQ4Nt3LbH2TLm5GhsE2eeLxSBTlrJ8Hu3ICSvYT51F3AbQbSPEQat5DG
fHxwt7Qm20++jdg0PTqfqqOjvViCpp5KyU9FvkjQ1+FI9jcS6xBOCTEXt4hSTxVG
OxN7oh8B6IwAD0dXnOdyIro0N2zqDlJhOLWkd+q5Si+sSfAiXGuTq/xopi9ho4nX
rQ+iOsNYdpHa3OM2TQwfw0kM+D9dtWp6HPj2t99UZcnquldVnQJs7QYOp9MSBZjY
NMNL3lP856u+uNa8oIMUO2G/1DdKglPJttEPfSOX4yFHhupwG9fa5kot15GyRcJQ
n8ROhHp2onm+gRtDn/HxqeFy9RMgH7jzuWw1cDfePEjiI5E4Q7tzEYiB3/gk7XzB
RAamB3NVFpIqsJ0GkUwIHmSsLuYC2L/OwuIDQIEzCUEXjPa8Iy6Q5eStWeY4pyCo
heXNxK8m+zuMf+no0RYKzSgCjstrQSffx0xbgULwtpbSuV2fBBZJsQ0/bmiDCwYg
BmCN0xBu4AS7d1lHDIrMq1PmAa/6nn5I/ASi/nMcT5so1RwjGZ4vz87pObifgPCv
oQHToSJG5orTQ/eDka7mlqeNvkFgzEvfvMwz2B/oah51GawGm3xAuQe2P5bBz1fI
aWzhjxBJHijPgajyfO8EdpBgROeycIcaxkDVJY8Q9p2zG6zCNfXuN0M7QTS2fahg
5RQE+Dy43CcIK1RCbFOSgIFCcPEWLYcqBFPcnZOqpaBCd+Ssthz7SWhGbFPCwHBe
R0BFzQjVgcQOf8m98tzBfvm0N2/l3br0urbAD54f00uw7GMa2LyvlhgpnMsAbjGy
ME3gjWO58wA/zxxhaxYSZBdwKebwJA2glxL/YoVUF3Ig/ptJNdgwlX2pdddvTOUH
Km+PJZBo9NF+8/bAkT1zKszQF4ofNqIOXBR57GdUkW7x2AsBxnYjE8qzqRLyeNT9
sVpxCUTYc14fbaEadxG5sRDaXD61I4YoL8nQEnihsVgETFoetySDk+8X33DwGA/8
+AS0LRGtU3TdV4M6vCF0JIPesndKu5iu1AnhYk2v+Ulm1Kl83CEjN4g3wdQ4Aef4
0BKkshn+I7mhli9BHwm710E5ZkGucOWyTPC03+uH1ojdJ4Vk3e2eXXsS5XFzr66A
`protect END_PROTECTED
