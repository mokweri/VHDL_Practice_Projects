`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjnp3h4jKhEAQl+zHJwi+IHGo1Ne2UlAg3Mc+I4VClessyhBx7oZI9dsMyccfRZz
3HbHST+ZM/FnTqCSpT7YxUJH62AW4003HCmfVIRLtpCl8PcVHfXIw9dR9zU+mzec
xeTygnxwbDVCbSeCPLfuQnb3xP0b9K/qJ9h4apCF/ZXCTrGmyKX27ZyORoWKFAv7
PH+I/5r4ZB9je0IX/x/EzzIQ4cEdWAAMQ+3hrlNUO0x+5286p8delMDannRrhSmv
JjOgnjpfmDybxVfqw9onv1O2x5kBEQ4EZ13bhV7Xwiod7VIE+1c+c81ViN656ZS/
eU1hx+VRQt5WAyYIQiSlZr1mdrfstg/og1ik9tYYg8okf8DQdT22hvDPxt9Lc95k
`protect END_PROTECTED
