`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LtZp/yJftWRz1zsKNmswM43lQpI2rkj3v/1rPwbG2zIRcpldXjCg/BJJoEe4M6qJ
jXNOSqQvsbl54Y9G1BalGfLlqfR3wv+Aiws/aRyo0Op8UDpYE+1Ka2SBndsTOpSV
M9vRjZqd8my9NBRa0/5bp7xbMCIcfM9sF4rIjV19p03x872cubRusFI/B2V0SEl7
nSJxOjF0wIat8yycTEfIzPbAdKOXqImKMDmOVbw+/jysFkFLPxK6mwhVNq2/nDZp
2sJOwPqFPpcxai30WFYwx7Ka+kgPYjZaTMs6pedqBhUlCSNaR8e89nk2fgd9AC/U
8lbQh1AM8gml0DL56wkSQDSJ5YPbNrb65xv0JDDVgVzlKOE2bX7Q+1QMt6RvKzQC
bjMpPIuVNi88v1a5qllJB7FFUb4lBbpsVQWmlMe6aBCvT73PMUndVYdfGsa6rgZr
MJLlN+HmSLn9Msvg9h6jdlHkPnw8pP25aM0KxbhqqvhsDPUn9lvpWetJ6+vZ2fRY
J48gTLMS9LfVKN3V1n9Eeg==
`protect END_PROTECTED
