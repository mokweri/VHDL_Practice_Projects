`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kC3vg24GZ4zXMov2rmVDr3jXQ731RBpswvnkeYToSSYLrHYqwqYeAzsqUCKMFFeO
r0+XYg8JxBJ0OX5x/wOIK8Dhj/vxkloY8YAS/1ZVpwYP5d5d6M6RetEP3rbmyiXt
o/mk3kQF+Xhlm3+43d4UILI7ELdWWzesh+AKAGrhsbBZWD5OSROFLsVGSYCAM2vC
a5dHIqB12xkV04A0fltnMJQ7p/IDyv5Rw64ENSF7RIbPL7jk2uWYQSoEubiEpKO8
8rtzsezpVa+ok4GiRwYg8AguxLqsO91oZmXsBXb2qWHiWZRv0FYmxPnNNJp8CuAg
MAmQCOAYMROWkyKSLITUzKils2cOgQItulm+5evqpv86ieEWXqDXrNGCXdsjlq+F
4C2kdxPqnFjBbN3NAzC1ovl/o+4k/Ryply1II0VcjUrUFcH2787w0a6Z0vMpa11s
h3mys/L+emLm6yLP92fLyOSJev7SAxKIU9nDZEhNfe/kOgkcqM2qZftP/lB5E+h/
9TKAZXCK1tnUbA09Gs3pJfE/zjvM9pFKHCCaWp1MSeOX5ZXpJR2MzRm08p2pJ/PC
RDFwASirHwxcL9YiLFARd0NyRf5SRU/y/YSzJs7u3M7p1tau3k4+h5Mwl14DmWO3
GDb5oXfhjSBn14PmXLZHxRbKKqhHs+po+rkEV7dVw6YHzIVKitap8+Wxgj8rpcne
nrLaRezDs+FSlwNu+EmNSN1e/qUsOT9dBK1bsTbbqqPPEJDfKrNwktidSwEZn5EU
fqAtWW4bjqBIxdompAFaYWziEvsFAQY6khaWQFzU2kgfzoON8hONvP3q/miFU7nO
3dtPJHWNSy7G4Pt54va7hSpIrq00bnHOubAsXHx6+EKl7rNcbRzf08zzHmSrPwwj
HWzZW1zKyTBTJGId6k+A+awS+L8b+78BKNNtY4d/Aj6S1JiIQC0YQlQkZnbgfWxh
tq6PFzzSAs+HGHPqs26GeRT4IcijOQiK+CskX/TLPr9Gc8m4NJtnvkGpuDxAeSf0
3G0mg/6oO6YhIebbvOuNdBsmXoZx6EY0kSq9/+ylBT2ehLGod+8/yYxbqn6GHtRn
1ejUZMOjXPHHHGSsRkkurPpEI2Ae1+9RP9VN/fLNlwoYqHkgTmQ7JRGf4qs3Scs8
W9pAgwsJl1FqqkLpO9FkKSTtb0BSjA4bZr7Wa03jXRu05sJB8AfJgaWcj3AF79KR
drU9EGdh+LqsrxHNP4sLmqc7SYa2mJ2akhZjwfhoiaC5RMSntMpBccpRKlTm8AZo
QwW3AltGGSqZJq87ziVhBhpkXfxFWaKfwJqca1exjXO05rFL3+d8GXKDfadlVCxp
nA/t6Ljt/wp2LuduztyegeGJjFofHepFnOjXfKhwxaHZGEQJ55iZBbP31ncHaVMn
t6QKkmdDtXiH0oJZM8h0TUz2iFD433wS9BuaWRNt4Fg5TpiI89AuuEoz8ULr58Is
3V1vCOQXfY4ATcJXkARn+J0hHvWNEYpGrYuMU6uKESdcX5MgXqO7flAPV0/RYNqK
+mY2aUPraP00UBdv6a3161y5Lwhenep6AA1rsclTa+CkE5Nlk/eb08UOew6DJJfv
aSUunhmlJKcpj4IeM+a8PvlKN9uGCYGxfJP4KrZoLtdBRxFtYtMnzbpvwLrMi9CJ
KCNVhJp0adXE2tEP4dvFc9zJ/ESvNim46MOxDaeWTBRZMtplCkV7pzUnpKWnZkdo
63koyN5qyHrx34g4oricTbRD9jVYNYa18nTUSlCF8i5EwILwqsgBouA4qz8+62yv
p0CwKUUroysMbMPjpyQb09F/87jVTV/qfG39tLTIY+dZetoT5sqFAaMSYVdwBK4y
oWeaLt5c5JP+kwozMv6d18+AZmXk2cCeN7+rUbAwSTht600Iz6zdRm+75eN74+Bo
ngfGHAIliTsU4zT9CzVzIt9Svbxm9KZPTsW3SNfFUEG+IJsALRpCayoPB0rd1zue
xmdJYyiY8D5VaUifNHIZa8pfXxJMc/WrwHC8tPxFe1/M8RCJP5VXGx8WwMOqQo3E
CJYix9JGhvkQ8tByNiWKLasG+KFj8clnIljJHuOZ8mrPWibej7lwIsXySaNpjPE+
rVfRqks3Wdf/86D1ZUrXVB/VBAnNGcB5sV8urS5QsYTsxxMWonwui00IpfvmJ/t5
MosDrxS7LN3m9mMxiNxsg6dQjzf+XKQSiFAmTxU+wDt7Z0FWasM94qFA+Eb5ZpnE
kzHIn2BtIAx2hG9JH7WSpStx9NJDdGipNO/079SeNo8jSJMtc5u4ooSxB1pW9BC8
GQ0NfqGObEKE293uFMFUiSeEBXJ4PVy2BjM73X1qPTLhZt7UBM/b7xopXPUSHqZG
lf9KI3rwANjmgNkUhFm+2Cv4MCLzVtUVppFJPskuQf/hwOBkQbqE9SWuTR6gkZcT
Nmy64op5O07qh8PtaQipbBhh6Jqt4N8Ok4ysldpO/hhR2K1LG+8HCF3JukvoL9mC
2924O6j3/F/W9UAYE/lD0JYtRPirTp90zNYoklBQjtk6DU5zFoj9kk7WS+s8OI3f
IOvwo50yB2HyDlsZahEttGLOWvpY1CO6VV5kMd4hl1kpmLAXc/7aOwuYG8gLqQYw
kd698MXqoRMbozYxs/IUCt+vD5aAAdCa5MD+qVgr97zBtQPPA2/byOyZGt7QR9aK
GIMoH2mXC3ewi7Pn3+RvD4KYygwSo+ZjGr5a9TsqI8BIzU8iSDwL5WUdeFypRbMQ
UZn9d2D6reOCC1Dp5Lv1tW2OQNBPevpGQVp6yDnfXhQLsxd5eWEaZFooHIaBJ5Bn
FlYBdMgoroiUSQ0H+sUfy60S1w29+Xj02zURB7v6E5fqcfU7fSYx5uNyyaaS2WXQ
qLT094vUIsW/RZPaIll2/O7wlfaQP2GDz5fLap32s/6Q38t7xwsqfQwM/UGcxsIP
UKUx/W96L9QtMEYUMSSVnkVUsBhLCcCr5goVWGEebvr/AxzSi15iR+tCdpZTiCuB
Hvxem4AcKbQw/ghNgYGVMcE3j07SMQJ/W+vK4G75iKi0kgICFaxVbk0vhjAeuOcc
UtWT+MxI4NE2DV5HS5VHP6wZJ0srMq2LBPK1qj86T2Jk0WcdJR5qaxxIZzKh/FHS
MOuK4jbxWaj7gm8ZxuX1VNvh4dI/sHJAOKjxp/AcUwJIjSlwyQ2SMXJ5q8HZcwjo
PyqziBGuQPv4QnS2ry5qa9ijdxv12Qec19yLbZ7I1K8aIgN8tYw1vTTFHx6Dh3u7
kKMuxYxWvKatgwCYoy9ulM+rgHdSiwWiCf74gPLZDRNY5wrwcLdj8JJT9nfinKIE
2XsbPKiiws9xYPRBSEUvwjVR5uXwQwnoqv+tttI8hzvBu1X3Sgyk7pvWzBah4UtD
GhL2tTzr6MyvGUKDdZng1jZQrUQKrbjsas3kZKw7r3p6AbSXFtDZ6ghY3HQ3vLbX
09TU2l7v2L5NvDEYMMZmKS2m3aOazGnFh5IzdyiIHZoBYQeo34jBboEDhSe0b5ah
y6ntsLOI2LQYiFBN950yRJQgYoK/ug4WCT4lVuwmt9yvnWOIv4rflOQtzO3QpxPT
gpu9g1d39d0Vzzalaqn9bn8TCdoVzGqxUV7KUkUcHu80ioots+Aw8XIojNNF99un
ZLstEooFgNv5j1LvQ4ZMPkHt4zfJ51zezZc0jlnazO/UbhjATdRA5qZAkFIQsEsl
AFJ3bqlMJTOrB0nTQNLrXzBGuz8+pAFvBKApclwarWycmV/rGBHzVcsT5i7+UqLo
srMRSsnXCX/OSFYlALJp9/sSPaYLK/bk4Q+SZf12PHW4ycPayCIOE+tyF1UktslQ
VVk0hQLTATkZHfMeRTjbcOogTwf9TC/TF3BkQTtkd/zbwz99zX2SmhfhhbanPnQk
Q9UJrZMSO/yfzU0dnS+gnPexq8AspmyzMttC3RCshPKFlC7ZqRr1KuV57hSRZiat
PI8gfhY1jmESCT0+UVYy1Xbodayhnv2Qk1zo13AZ4rL3HxSSmXGBRgAEDKNDHc4D
gaKDwm/+Mos2aKSA76dQFDnXBWjrLoMUtW/gulq839SibkS0wRPT3q5tnXoMsWbf
QQ5aCSK1hrbzCbJaivMieuUuWSI8Fu4ucQ93ZPnLw1wFF+ASXlcaNGQ5IwFKA+ya
oXAJjBNe+sSaBxiBz4UldRNW72Srho2e6V97DPvVIO3gbqDMuoXk5dSNXs1g1QcD
5u8kWlFG2wJmqBF+Uzk0ou8F2zeWdbeN3BsFYHvRIINDXUMQ580/XB485zD7+eqa
E5d4SiKFKqv25WphkOQp7Xjn5urA9SK6h/yBj3d2GkWPOizmNWGZDcpBBY6G5rqI
AneQmdRFZHXBNw2557oM6Nrc62EMxrNg+xXdZoQUnzLAAimEy1ggTFDx21Brh10I
rH095mjxni4Guh/kaFoIbl441dHdZXU5uJU7G7/kOPIo6Rh9eKDRK+c7KoTDmZF8
b7m4N8ssi5Euv2zLw10tWK73+RBB4NWHzmY2KyrTkyHw4EkPCCVNC5wY577BWdFR
EsH21/c71MxqShKSw2ZmPRsLuJAspKmIf1PCQyJmY7kuaT4hbg2acd+Rp0vAtDQB
yctLtxwcHazfmXG8IZsebQI/n+HIMeP2V/djSvtqbLgaBHG0larHCweIklAiqVFk
bv++3mhBruMpU2UBj/yiHAqFxmmAS35YWPUqOxiW7olc/8BYTTE5ZsEjaYUhYZyK
uhA6Itkn681DWJOfjxTQajfMGhMlpexgess9Nb6WO0+xbmQrVcy51pqfG5DkFfp3
miKalRHGm4PtJGcJaR8aXrMiq1ZVlsFZxwqbURy2aQBHS3RfQiBmms9EcPA2Zapg
f8wA+bAsMHYZUVTQ6BV3QfdCRGaCfSuNMvqyWugN8Y56KYWb8kzrLVui31Td57ny
vm48MJtmYhTKzaAYDNUM6XIQk+n8YD1AnmKZe0MvjG1lhxdEZodnuEzP2tpZ03Ga
KAaHqfx7h3BAQfayhcvF8CQjqWJyXB9yyLj3X/a6QvtSfEbsQeOcNvDRiy+Fqb7r
9nEehAshVcfCeJt52jHgUKP3Znu9yTgUzcYX21Skxb/NXq8ba62iJBjE+ADnozoF
6dBbtTtxAHKQjtXtQAAeRxIROj07RnOrNJw244Oc1kgBg/Iga37qIyuWqy6s3PmL
VIEjNnhRNmwQZqPllNRYCVTgFDM3sGQglkzoJ/jchFToPPmKZgCT+6OzXY91Bui+
PvLjbb1nq222FWIqeRMHFPBm+i4GJh04NMv2ZKTea6if7amN9kukytDv58zHoglu
AebFw4p4gW4yL2rLiYEADZtTnHLnqa2rTRCFB4FxtgoJIT34OY1PHVshb0G7v5Q1
SWS5AxM75lKkwiXx5qo6oNQWYlUjVvTkgBefnjegiDY+diWK2IRwDpQpPDlVkmqm
8mvoxH4/qj2Gc77SuyqTBLON3fEu+XC7S0IIAa3Q5sD9RSxSmNB5IcbsHrg44Rg5
Zg5qHxnzMKB7NsYFj66ewUxNkgtkSaO9xD5MbgHYjmGUalN+q8Y3lf5hGV82nbYF
Ipss0UP2myt0PiVUNpV0Mt7KUpHjyW9L42DbMKj5kQ6OqiH++/5dFzUcgV81nu4x
KutrCXgKkUc6P/H/QrLD0wpkjAgl07w/+HfMAJrHDsXaqkfw+IWrSVPbcKlL67Ca
ylkCjID08mTpIDqob8f/lLAB55D3Dlsz90nzTX5XJNJYhHuiZcoWGnNJrNRRfYy8
Jt4CMo3jT+UtPGIFK3DCdtGDW6Fy6o7sWY70Oh3heT2hKx2JcL1MobAz6pmV4dlP
b/yiOK+tQZeTJd0opmFkdcySurWdgnFadxmrE+TtrlCQ7NKChMxUG4fkbhfPhFFI
a1jrYtEFsVD9DJ0hmT68Io6cKTYh3A1NIX7jlcyrtdQM8qwHVwtyGdnQQECFB/ai
g5czxSXTBr0XJKF5sUUID/LlQJMDTimad/uFbq1f5UJkuR03kbFeHtKUrrgW9tEp
fOSNs8LEFIBJ3Z9PA0aznT4WawTsllQ9Y5TXt+sHZ7/WrFESnuT4iMBnJKccOyWd
eVf8FZN6RZ4p1qIPUCwUVnxnoj/6Jq2o6ZfSKNN6EDGC6TO13bJwvf0PumJ/tfm1
we1Rf4jiekqPQd8Q+Bqlp4I2hFtdpDxLqbouio4SHqK/N9i3/kdIKayP0WrFeLzq
9RfYo9H6Y43REfayu71YawM+gvP4qmb39udn4MWhZqPe+xeckjBDkcOARA4GNkZu
AeH7zRLsGIHgmktlm3UxHktlOi6x2QLVmyv2S9FAVJGGVg3wXPNmHqRPZ86tpMAz
v1AUjHRJALuaPwYjqSJ6Wo26xk8Xgp3A7jNfQNhRW07ABvLYiejza3qaIevuAypm
VsGW2y7X90hg+o4sGywIa3WQG6gTz3WE31LUj0Fl368QNuNxBvxn4U8zH9g/LLHm
cbykDXIYLl2X7iilpBO2ZV9+jfoL5U8P6KJsrned5uRCR2bJJ2VKnoOSFLF5BkkN
ba2b0C3nu5jdmNFg77ComBSjVS9rus3q1WvbCmYBcjqJ42rF/R81uMtDszevEgBx
p4peC1pC49die6oSMtioS/Qt8GIM14A9m46yTaTNqt8d+qlxDYq69KaK3GKkYoOW
TF+e4mfV1p1/BymscI5X1glpq+0IcWKpPmSyk2lwcqIupyz3X/NK5umrSaxoAp0w
PckndIzJe6+1tTwk2APOmONIi5m6fFWsHBXAED/yMlBLjuOO3wyUHXAtofNyRpFo
rfFhZEgach0A1IawD5Nqmkw43PEJZBZrF54ME03uSoI6UzNPlEPAh8aG73n+/Umc
ym6CxC/ss7runbNGAwUvdmeW5GAg5a0DpfGV0+MZ6b912EfV/UoAPqcAp5FGH5zh
pXFgmY4Zc/k7654Phh5vomyMHWrmjJ6gB7JnWfLdf2/NS4LoyiLdxZhyXOhMdZu3
m2sOdHL8f8xEp5gfjrcPAWca0TlQHjsaf8AlYtolr3rRTSztLh6hQZlNQHLTfJFn
mLNHwtqdcw44glgBoEY8crajJZ00UZVWE9XVAgj+/5fRyON0uO53XbuvJA/0KVRm
QXpiWnoc8cKhCLsAWofct/eAFv+zSKgnL5DM1h80eevnM8P0UgAocHmkZnwAqpMq
uu/zUFzMPBQg9+qasV4dUmCmw6KISYiViVVRAwIay1LlMmrdVa5kMS25aMhewr8w
gtzVe100QvYMh+Xf1eOsF1KHaWmKy00iJ5Gtcq9CJvavMsQJLA+MXwgxb5kBZeOY
TuJEe6MduOGs1R3s04PRuCbUN+8du7/N6jp7NCykK7zvYJAcNjg638QQRE98elqu
hWxJIwxOi88wa7zHCjuWMiZL2voXtG1TllYEzzkKF8xzagC8qopkL1/Dfz7aeiNB
Hab18HkpQvUiVHycQQ+yjV0wVl7iM4wAeeOia4D/uYfTyv5XZVN+w6J0xOBqsPpW
220a3Yca/7Z4t8zZe3mDfDWNZAc/8jV+un6+SJaPqhUtcsBJMGeIo8Gd6PrGyVK3
9U214aoWEO7XXktif6OdNJ6IaHI/K068VH3nMBjvMoSrlD86BhIj7quCQLhQdn+O
w3OtB3/PuZud9N0nwxg6G/I2vykw1ks8M93lg+0miIe3Fx4HpqfmWRHGxFOz6oLu
y6XVkOEm2YnZceKkgUcyiJTCz62f+pZH/FZUotRoAreKXttVrcPX8fX/OxbKbx/r
zENGql5dUVeJX+rZQxz2Y9wzj9M0vS3DvY4kVjVv2JrfjK7Zltce0hJnBHNyIgqr
rnZGxMjKrI0YS3GKy3SBW1X9yHlAULqF1931EBcTc2uWG5+j4bayXx67X4xW69Oa
lDGiY/pCGMYdjAQLwUcbMXMhC6KtJQ4nQcupRiOQFZrViaBLZgUJZrq4U5fLH3vD
hHNhCx3uBnkSJMXkTsMHHAhFpuoGU9IDvevTvgJyPr38rN8zNX+fKNZxlmagaWkt
b7484sVaV2Pv9ZKIG30rXsphEFatQJaDq6+7IYs1UGr+xSA7woSIlofy2zJItFLH
DpJ11LJZdeRwEr9E5CuUlRhBa5RJYw3KQTUiU1A4ObdI4iokJVoMq02a1JLWTVaa
Xo+2LT3/epgQee/z+iImC7zOWqw3UVywPYa73pJJe0xYEJnCA+8o8fUaelnh2bYz
Zt0ZWaWia7R4CH2vM89Mo95kJVD52PNgRqosBijMZaCvwYvQbtiRd43n1nCFzSFo
qt3NoCiL0auON+sRgGIqZYRJ4CkJnBs4bDAr4L1xT81Hj4h9gSGk2j9W2mbdlN4Z
v7axBWsNRSOsX/RzLFWGmAw+tameJLiW5Hs/XZNxeOMzIAPEr4cBnOH25KsIzYr9
hTyurj3RiP2Whh38rfR4PCxTc3Fke2NZbQrzsaklAB5ufuH+QFwQoYPm1ygcECTP
0GyBse6ymO425dwpg7e2cr/RcYzpLTe9dfjQzPNkW2grX9LPtOZQnD36R3IKgkwH
bmT4JzdnavikxLamu0E4NAUaz8LwdOnrSVhVnqvKE1pquZoQ3sd9kPbC47VOHQMc
26f33MT7jsPQZOstsjP9qe83LnAJHftuDyURxLKJCukITrIP4m8N/ACHXEgHo63I
2PshQvDiAT/yqRBHFxZ9YwGCWi4R+RvpRPTyv6A3zxd0j9osOteNUz61EQ1li/0a
NevWb+AErU7ckPPfUHdZ1sGNZ87LoDurjhDOjGTQYEButNHHA4Y4mM1YfPGLumfL
OuoODhIGR41ra/YD25LdGnsg0xXbQpZK/5VOZ19Dxl9qesIUYAwuudZxBmXs1M8l
Pn217eEqKY0r5kfvIzoMdNIss2ZRsstcm/VxqxbdHrtgQTmznHF2fbvvZ6hPuLeT
I510tBiSijSexZgCKs5G49jvclwYDao3Z+yV0T3rdaGmUVa15yTFwir7lcP2Mjo3
FhYxl5+URvwWZTgUbt++8NMMf1YmjIisV4bqyplJN9bufTaZX7cj0sfMXR2O2e4A
VCX9Gh2sxKFuWSG6NWblJGC6pRsCNVTI49n8A3I6ogcgxzmgyv4elAmnjFVIuaHo
MItUKWymb8qek9OfyFn9vGt1vZhEzBe3MOUIJTg33KeYifiVDCGTdfkDhniJtHu/
bnYQ/DjErLrEKKZUfyI5eAQ0rhxkPu46VMd87DsURZY/tRRmw3ld8U6ClISxdnTI
rBpvy0Fh2xx92v+DKY1URRC9KUlrqM7yAnS0GENq5J0PLm8Bqwix0v+Q/MJV7aAb
bFH8/lQo6UpSFsbwulIWb2Cd75xEJDR4pedmSHKR9sJ3kxDZaOnhKq9Fpb9EkdiG
x/ySa0Aov96gHyM/lcbshfplINFa9+K+av91w06kAu7E4zRUlrfKeO/jYhSpadiG
yagsR6m+ig8U8oZvawGvaa9m8PM0GGls4ZMy1uQY1TvnHQjKSYJVsWFVoA7SEqUP
NuLIrbgEMTjC4Iw4+UjbSFFnvbaHcZ8hQgdrv8SXvhOcUfENhyfnpPeLtrh/IMHC
c8Y0vcUxCXy9ZFWd16D6Nb5OHF3MbEaFb73rLYLnLpPHo13bvYRd4aUaE7SqErMP
kaRiOua+aIQJ3SJLaQc7nJfNbIlpkMDqGvvYizzG3cvU3fh0sNsyT1aqTnqIAEoD
piIt+yhlmbQp0KsxZMWY3nxGepX4U1FuBSrWr1zHvJdBR8/U1e80quMmrf7eYYBy
AisiH6m1uwjhcC6FuEqLkpv6KX+kHZxr2A7PB04EKs3jtw1DkqOPWSg8Yl+p593S
eU9T6jgAqmS5eysGxrWLEzGJXzJhpEGjm8v3XsRpSPTPf8Y1VNrG1q62mxUR7AI6
9k/+1zoESm7aMnK1FvLmxePCxZgoqQOpTPu2U4s9T0vxuu+in54c/3fhUShsT3c7
H4zPZCGMdynpK8SscU2kvlJdX4spjKn/Hbyv7upkBUz3AE1ZRi579Rm/ReWr6rHJ
VcPNDzqiW6XwXkZo2glzdOaGYl+tFHNRnrgSbDeZxHsWOsEqri2ZowlhUGjM9K2g
0LmmdR5oT9scynDrmiviP7hxpsn7EGJH4wqwT0pIOcmzzIUGK+4IqQx3gIOAgCnk
cWA1izsj5jk8Bf6/525Ry/OhHzdwQICUWWpvi7NepnVrvTepHbqbn8rF7i5jeAgJ
dTANQ+7b+PAsNZibD3BAGW8Ff8Q3nGJCPpsFcL3QFvbr3DGGZPdryrw4qoSQU8QV
MhwcHVwyXKUsv9OEDR4HXFH+2yCYsT/24ZaWUV21FX2mXfOzAIhNYSg69S3u4eKi
4z+pds6ktFzl0WUfyUEax1uPb+Z1ny67Seqp2TwFsK5T0OUpRqaJqs1nzT3iPlPR
JOqOZl/u0vYZT9XjsTnltvfMNvWfZ24OQxg9xWQ29LocHYB8fV4bOt66wa4sIigk
t8Owzorkvg0/c2+TZWyy1cs/mgYvmG5dbTWItA1nafKEgYMSANg82t3JUNFxORwZ
35Y7xZFS/qRypyV52iuAsoem5avoPNo5PSQSHo7sks5HTFjydGvGKuJDXKB2azmQ
6x5Hxgpaky88fZJaENKBnc5m7XVIYXKnHtX4KoGPuaqYEImwG8izcH8S4/McdiWa
/gCvqu96rEg7O8O9253AJAzTt1EXxEawD3FPFHdDPBTEyYEXZ2paTv4IkNur8if3
bRvaZ7i8iJ5nBDm+siC/UeRhNpLTyxWYbCHi7pRgBNC0lHLMBu+nOQ57h/n9zEHG
WtYmHtV8NFpCiuxmYSImbbamnUKPFBsQUFq1iX74ikC0evpUsscT/y0+kZYmgI6D
FWueyXszwt4FE3vsh1txKqgoEDxW52AGCi7U3Ej214GXDXf1YrDJ5QXXdMdNbmBc
j3pPW3VP3jwXIOHGCrGMCWhWriH4KaunDNMMrlwgVMdU34VPshZjdqMq5o1d9VDD
9Q4BzOF7E7reo5MQPim1c71z84Ab3rC7R/v35ySuDtsRt2uWE+P1XsfJ9sWQRjty
SPwiRVgwitIQtoWaffPmuRR9lC5adxHqTy5cr9cPDatYjktL2R37v4TvhrErGjxL
Eji8+2fzniFtN6GcT0+3XzDMBmseIOAZ6r88KWOGONR5SbvO/fCttBJ6W8GnDKda
2t9CzuoVHKi3NA2P2eAZGp+IwKe4Nb+8njAPHkr3JMOnp1NMuNYBj7Oh2phGo5jP
ech+zKZ67ULGMhIUby+80bn1E3u3v+x2T3VwPMeoboFBSWPNMRTE/nDvk6rhF8Fb
Nlv3QL14cEyKUzo1zVkQcKM5Z4+AvCfsjzuzHCpu8nXRv3WBobGWfjE6XyeoOXaV
GqQOeF99icJv+T77uBWGWj8YQ5neIC2pyLD3WDVYQ08bC1LEhZhRv6BwBYNT+A7s
yTYY9YoXs96L79lSzZhTZHAI30LZFKmYJou+LQszytj4bAvaceGoKZgUGGn15ZZh
QA5hms8NaqfA3EEn5mDaN+KOYlgQeekyoQHUb/R5EXS7+jyfwCO9IXLi1NOS45+4
dlUe+VEwxRO1J7Wd7oqCLu46eNF2PaCex552CWQlWFoRFjGZOKfaH8CPtlZCt6uh
q9YrFKguIA4hmQaSkG5M0889lIroQ3s72AnHAKHARjuGX7N0WkyxW0cO7tdBbaWj
4ecnWbIlFe7l+U66gNt95y42PDPlP0UGUZrd8UtP/kFuuLsZ4QUVpukZQ26QAW5C
XpPvw6stL5hGPAagMZrCdaw+GWj40pPddig5WnyqNmvjAnZOLGdoFmInRu+kTlzg
MsMAvHZMMPfY4/HHI69narBVql5J8Chs5VKwvG4hksy/aYrPmLlqkhya2yk7ujMz
ZDuJC+9nbi4ND9zQcJpFWqfdR2YUouDYhp+jHcpxTtQA9Sewb+zablEFWvoxLOuG
HwAKkTPXGaT8kUcodKRPOeIaEZ/bFt4EoZ1qUZIhtSaMJShWrDtwnJrakEA3etVP
tHsFi82n3Z7ff538KQgxgNIqhPdqH1GZkjgPy0nWB4S5FgRS64FWbY6SCupfjAt/
/wT/m3MjiIOXKN7gQWYRAyIrMQYHiJ8JP3XFr68Y/9NriNOFbCxla9b9bALKOynf
Xih/6HPNVPFipYtZUypLzxDo6uqkgjahFkRAg90dprLqzvLA9hI1HRSHcb4ct00C
rqxmvaxiEzLjxDCN33Efp9zpGSXWp+kT5whs9VLaY8Z0/6ZhVelKyqpwQGoSPfwX
NbIYWpFdQPbqVCP6Cpisc6Rl7S+T1xabGlormvuTGu3NV3ZdnpN0rEz8h2f0wGdn
RPYv5y0B5VYxijKM9mNmt2cPaX3CI0AJheg+FwGyKSYkTJ9sPg7yD9MwIQ0DVEzX
aLbMT6K5EkHpFaYxCPhxvxqEZH8Qxtb3EVH6pEI2K4oxMoTpwnWf2oRxefJjvqrg
wtmtmGu6ex0nR6vA+WgnMBtk8+xoPozgaclmL0zawooN6K7NDsuZZWpTshtPYPq/
2ZTqlxESn67CCkbq0bETKEboQcnYDOmt2YXZ8wkbSFc8RlNm4Em17bBVWQnnnbHk
MzhwyDXoV0+CvGY3xdtoWt5jEDg99Fkc3U9dse7u3BSLGcMCExbFezVaE0t2ctJo
JR6mzxT5uI7qwj0jrwARX4melHmIDtN+94Cu3oFiieVbCWeY5l/hamuBiZBh+Sz2
IQmSVrYg/UhDXORSgkrOy6XIgB55fUMcBhg4Uc4SbDI/R1rMndPjFCxmimu8XA79
hi+bxHkQ0kVn3AyslAGJwUTUXtT1R92UMYgUfLUhy4+TonnUlbPjofP704hvQExW
vQWWKF06LRgqVswtjI8C0nYyrkYBBK2hu+HZg0mEkbV2bijXooKVMrjePYIo+TY5
dhP3B3Yu+PUvX7o9NnWDCfjs8copwcTSvqVrTHxLksna7bNAN3jjt5gXcVWRFyUg
BwUJfNGRHo/mt/9EpPUbX9QCCVI2R7F0/wrCWGs5nY9zxihKwwql0/JH8O+tVCYj
ijXkyrFd5EUso2n6fn7YKRHC/44hFpUJmn4GcxDMOfIubDxRN1ZLC1DCTkN2Ui1X
Tk0XwTj8ptZgyIY5coYH2OL5JXbvivDJCulCaxQ0PK3qhNQyOSqrolvaFWjOWiY2
2SDCHxxhcvYw/ncMIbQ9/79r90nteHPdWC4Ic52JFqWwec8FoLcOBLrGYqt4bHnZ
CsXfa3t1oiguNfIc3gqXFCYxSJjchgfQ80KK1texBoCuRqdLuXUxw8dSJy/K4GlP
5bjP1xS8kQcg+9cRJZ4g+YibM0BQoFUxS5f0tB2kED7j/l9l9ti2uS/Q/7wegxmu
6tEwms1w06Ta89HSrWG00w==
`protect END_PROTECTED
