`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
is4y+hAwHtuw09ELmzLOw9RI4UFQ5FGM0Z1shmO12dgPe1lkbum+thZdB1lCLqmI
pNN/VOkCVjS28encvhylmyysFxdKx7BOIi0qzBEXV7gOBSMLroMk/3ZCdReZoO2h
HMJAqygHCbo7C/y0x6W4+bP9m/IcaGzHtnmeakfQ+ueXGffPYLJjRD0/Ihcgo3dC
/ZsjjbnafB+eK+a+ut9ZgvNJl05Y3qL7IaTiWf0/UoOkqvHM/UfRtXUx9ZAKBDF1
FkJ1Avor2j2tAhlwcwZ299y9GRmToZ2xL5aEcrPIXL3OdSYuJxri/Il/CQL/m/ZD
sUHWNhPgmyAdt6hBWRfBFeUfYUsbMVI+k26M/V2Pq+T6qmLhMufT+6BEuFV5Xqix
o6i4oucYmZ8UH7Cv7WDY1tlo0Ew4qxgd2lnuVDZdvhNoPXchcTKVRzXSOg+1PORk
e5QOaHPm97W+K5unZMPsHji5eFCXBvFPopaqzMvqnNS4EYyT7HrOwL3GbGGP0mvX
8tNtRm8rZJxKb8YxlDd7ZxBranNzIrBDGiXPSoOfd0tnVMZjvtCRb8q3xS2z1g6h
HFIUGOUxC5olkaS1SmhjJ+qw64XQiNhfL0FZFpynp4igm6O6jZ6ZbcvaqOTEc+Jh
hkhhMO6ozy9h8y3GkYsKusWDLJ2ecwnhhNkDUWhf1FMGmTJ2crT7kJ8kzc2oK1AX
dNLbMLJ94WNWIhQSrMYSYqfeioe3P4mRn5vmXIuDwWRGqk8Bq/0OTU3TEpajdAFh
jStcicYErOJokeE15WWE+KSJvzxWVuPYgIct3ULjELrLG0WZ1pw6dp49Y35l+1/u
ODjpBgPtGDGyPKSmthz/pzE2Ka2fvOPxctdbLqAblnRFBwlRjYNKCNlQTpBqQ1Oo
TkNNnOc3JIT9ZD2m3kM9N+/4ZR4ikGzRd9VQGVAJRw566GM6InTIlCr1yN3v2pyc
AbUAP0uWABepE4V3IDzAjUsWRfh2EvO2iMtaC4nz6FWIGhCH+PvJW+QdCU+tpLKA
tLgvWhSLtzJjlNr0tuUaj3t7xQb2r4NbO6eKOBR4KCO9t4A/1B9wOl2+A9deeNyc
+HwIVr0eFsGsz66bSa6eUaw97ElMhMAnWKZdDVt4KmjO1mxkpfI39LCwoOTGFG8/
fstQpYovGXG7TqCSuTnPr2ICpWM6HRuPDqBF+PskWPDivdEO18fAi/aBw2smuO5T
Qn4nmvsXOM3qUiM+T0BpNogrRSMkeLl46f8lPmEDJmUx4vKFf8DJ/o6e27FdmhE8
9Tz68gIZ3MDC8SHwDllDMseREWDYDpWph6I/LOJkQVXmFk174OtTXG4Y4FAqbRhk
nuULGzNZFxsPbJvcB8kkkAIROzakrVX47NXYDGixGbcPOsWyUBWxBC6Q/4s3+1DV
1LV+po9MfCR0Tnvqjw8cicrH6vcrestVsDq6w0EtT5+q85/aSR+Fdr4si6QSgSyz
eULkHd+2wJB24qdoyph6lFwu3CU2EaPfygOSvZ61Ax8kALPNutXRH1V22nG9QIr4
29vFfwAMlg21hZ190tNacLR8GwvVrnryc5A1IMOM7YQimicyzpSThXvDtZcusGWK
kT/cJ70RvgZE+1YDeHSUY593gLLZSGnDhUqpddimoSARtHtgpUligr1Rkn2xnn+J
E6UsnzNq3lsjafJNkRcHvAawag8oUIlNDEN49KKSaL+7jA3PrRi6e0bdPnGXULLh
jYDz6kkG0FG0dqZHBly4dLXbUTK2+/VnVqpa2U4LIeDOye9IHJ5x8vZINXLDPvyC
3E/P9v6nG4I1UKTFyNNnoCVOM5K6X1dvzlMdgx7XgWwTaZQIWNJT7wxeaLtyHqsv
VYgpe16/ka2fi+3GxltcmhP6bOULHvXjbTtV7S3rVO82YIFi/7dYCFf1wDzDS+Jt
g68m0M8j45XvEFqdbvdSBwLilbLdjMfzotaoeu+eHP4xQcebZ/xP4GfVannoSOqi
dUpiQcnavnuDpY54Jcd8QFd2JwNo14+lMHLnPCjPdo34LS+0CGv0wA1QfjF7UnIy
c4tYq9Fbp/pgiSq5uJNgMYhMifQFe1tUQXGzg5GnErf/J5nWrQmzqnFqRbRodcbB
eFgylnEH7SSHig7Ay6Oy80X43Utnbt115F72/jfJoMzIIx/B9Uc5mOPZ/yuZawe6
6fyeCbdwIeFqW9aMB9DCgIPIEblMVeFBoOpSWsX90FTFqW/u08P2oQ41/nfz8WVc
MRGPhB9n5KVxFz1ClBzUPbuwvdzlZ3YfPvQNNMUHWtNzecFLs0PJbGf/l5j2PHDV
tHTPCyg8In4hL8DwctbRque0Es9SINbZx67hDRxD3GpKtDAkvNog8QBlj8VxFDWS
qiz+PFb0EixmJQOZz3wlcnxg2N10C/pHpZkm4mJxbre1YZkPExc7JWP3aG8mrizE
C+reHmOoreTfIFAItRGR3q9bdS4/3aggQJ3egcIaVt3t5LmOW/Z3iL/niYtCbJAN
1Jkzzlpp7nQfphYa5fdrCx9zj84LR9NRLnOhjb+JX0yVouYQRCQQv1v1/INdPUlF
NQg/8S/24aUQBO+dR4L+YnwP4AJxU/wYDes5K9PF/7XwPPXXpi7FjPgDvWTDYWFn
9N6p+wYnlR1qRwamhiumky+DNRWUkvD2/bIm6vnFZ4sOG/H+G/X42m2Pv3f6Gycq
QxFC62sB9vqLdnObiEpHi6WY63FMsbCgK3j+N/8hPQIElJ+AmqQYiBiDH2fctcgn
J+fdhJYsjPkyaOeA0yuCI+EwDo4yPqqm7cr1Jsao1dUI+sB/hP/MmjqbrX3q+ZPI
AENtLcsydhVJ+A97KuP0D9MgDIvnIzahF9Ya0t6ABu4=
`protect END_PROTECTED
