`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pe4nYZVkkAlzgo49co1IftB1aqXI4Ak4nA1AnTEwe5Sjc0TwZwR0qmE5Wr24ZY5I
3hx+gS5Xnchu44wNYQQ4d/1wvoBsnphTU8mrTeeJzQz5w62OjCgYZxeGMbJ50012
o1E8uGTdfD0m7rjxPV2q1wkN4Qhy0qgI9wuUtlvhK7lXzOX6w5ucFvjLfnNLySwA
19JVTkNcDrOTGt9ovZ1+8GzAoBDSva40PLd1fP18dH4MSdh6gk4wzGwTlTnLJ3dL
dz0BuqZy+D2aHidT7pit3CTTnyYthxC/IzKggfMtLa+fly2dO66lZcEr6iTT/TNW
Fp29CQwOLUmdCeey5G84hF6canLXJNpgzZ0gULBrNicxPhyecF/xC37QgTJWjyEQ
heRh0Pn0c/CCAwP8xEGAvBHOk8pJnXtDPVWqRpKrwqaxYiZl/0n4wVC621btb5tw
S7xaKCb38NDJMB4QqIvhU7ie8pUTEMr29p7TqmGRfau7yJmU8PzVKTILDLW/gVoi
2+PtlFqwCs1yCWeDgxfyfi+XthaZYt9FRp+YKSwEyvHOlwOp8X9KXY9tEX3/REPW
BPDYKN0In4B98fJSsFs5/iUX1kgwE5zR6stmfqpWVWRozsUa6hHJQqxWC3XNMmg7
fr2iH3Me6plATp8n7UwVHTmjZ3xvX4hF/ArlMIhxdDP9Gk77prO6Lt0AhL1mYpC8
Ztx/c7J9Ev/tdKxS0s4tCpLpeoJim7/rN/p5FMd8XDbXGKXfc/SRhmUYzNEmYEK+
+jxWmPwMwdZxkF9oj2IaOEByO+KVo6wf5DprnJc6GbHo7PPb3h8C9jz3keML0DXi
/EwW35tgSWRICzhXCGpaBAOjwjAbtene1Q1Lk86/YrGcQ7IpmSVcoF4aY/TGlhQn
aCxjAHXgunxbuRKbfSQ6uitcVkfuXA2rBiVDzWPXU44exJiRznrq87BH04r3q2nc
wP/y9UHotUZo1s85dYNw5A1qJnJ5PTn43TZieoI8apV5xjhFJe7VjAQu7sVghLd0
2u94wyQHUyDtrKYGEotqvqyCz8hv6+dBhkWCLoHA4EALc0a1ITZkxUAxkjoFyIG7
EuNQpcVZVMasr4TdZWHIfr8fdjLQi3Iou8sbGYRKc+DiEyXITQbKJqSg/es6iK/G
2/ruYR5CNLsBjgf3NHa4Gfc3WpdRmfIeTzbTOQ0TE8JII2Vgn2+POZmt6EwMviou
+mWXTrJHX87co1u+aRPRoKFmZcYJQKFGdebfo3GpGQy2wJvPpwJOD3/U3WT2+vUF
/jiYL1U9wZmEGlMVT4hAnX6bJ2a80bEPppilTNXbOXXXxMAigZIkB0Gsm7k3Pk6M
krXlFn02cXRgY+jh0x87bqZrMf7dmr/IXL9+2Yj4wKhlm8JWjSiwEqOmhRG2UmPS
mFvP+XFamS9fcQp+jYAflRHEi235ozEBnj5RrJ9Xhr3Lf8dK4pRau+iNwPXC1b7I
`protect END_PROTECTED
