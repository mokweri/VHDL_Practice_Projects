`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zhydVFrh4M4IGiKAkKARem19BdpSNeNN1vSVKtNBtVzzxW4dSRUPC8yCgnmk6Q9s
wF0qByoCHHkFrtJNTOgM/krbuZupjPNS1MvQo++cWpEdOAMAuihBFae5SI4UQYxX
0fHzRthcg6IYa+DKDtmBQjwx0MeE4BB9yjowqv0fWTKONJzo+9Bo/aYCZ1vLQnMl
lz6pr8mIQt4NlthMBUvYvSepjT/No9o/nvH5R06iYUS2iomrT8SQt64TS0RTpO5k
UNI0KiuMr3BBk0gAZIS58C81v3q+G/w5C1/JjqpWJy8qXmi9Vl1knuSah48+YgUm
lOnrDpX47jjYIbs9a0ZTjunSKcVUp9ETtTqA4N6rJvztFeiYDeMlKzJAlmp08Sdk
D/cr/8rji20aMYP2i24NK3Y314aS9/Y/FQyHupC/xj2pWobExYrz7jYmJTt7KqFi
Juunqowk/wlufNEucVzOwCVNTvwbUdWuRLvlb9ItuiaGx6TN1s+MF0WM6rdMaxTY
QkXFyDGoNJaPGpURdeL7Fz2Y/l/MiwCuiL9jGbPeug3OiJxNvZKHasAtam2H8NqT
NZj6/YOA1n9l12s59+PMFP883EJMAfb6G8bdVHAwQozjCoOPKmrKrC/SbPoUBL4Y
7r3TG+epqYnAfb2wUPOHu1wwPYjZkTo+FTnQuqrwg0XhMEP7dsNVTr/x98Wibj9s
sNkf9Smsa8zJGVYx6cfDbu7OJpp2hGTdq36suLnGxTs6PS35skrqy0tKKyjwFNAf
21Adk1zaOzZzzajlLOujcZXomzKI/Hm7stDrXH2O+CMfIvrZBzoaUHDltO+wJ/Oc
L1Z25cKA9w8l6aLFYD1vwFHVZygcbysO65MrMAiBt5QIw/H3j3YA5tlQXMuzz8Gr
d6BhQPVN8RDEJ9Ne/mvfoiJ9l7wIzKvi23FAgHEY5JHeX5IsP4K09iVveRWBcixn
NCseTgwrepWY64f4u7clNujxTupYSWHfyBE8E9Nds9yrn9huBHaSw2BAXzVp3cc4
CJhMHxEhQilWUtSq9Y2zST1HIQe8/XEebOnNNzTqy4Hfl+NLKdDQKTLsqVFU+o+i
TMFYg+SDeRxmsGpEKJyeeXiQQKztDmz5p22VAEJoyQN7mTXgZr68Cy+1BVhvc7qZ
9wy5f7nDrRt2Kf1wpkksvd6FygLozN5D/CpNUra7KDpwVqrtgo2uANjGIZNJH8HR
eApFw3r9W9Gw2Ap129keB+W2vgds/0ZUVpjQqlUrTHH6St3N2QSzOectNGZqcLs+
wsoh2E94qK24So96VuAl1y5we223XKnWgqCtMd4G3usObKWiJ1kJFIewK2jY9MsE
OeySzoe2rj4sCcUJ2/g3P1qw+JvIsm7d7K2iDIXD0i+A9T6gzYVhWa7rUaAyQBya
0+bJPi1sZr1awdKeKGGCqRrtxHF/ndIpJ5M5koBCd1ZDVIBTkGyclr0Qd8c32k6Q
K0NgmLSiSp0swSirItUWyglZS5dkxsC6jpee1HM9CDJ3tZPeOmpkTBHkolH/5lWo
4Ii+ygYAj/KmH7BIXNUqBacoL8unpA39TMNlX2RVKsFgz/p9CavGxhY5kw+PsqHx
aPgEn0n3YmGdYs3fKSPh/mj0Zxr5FySGikDqEQXgeDXkxbLf8YXLWs7UuYVdqS20
/2BGqqMJ8Oe9c5ma9LmqyiAqFL5kX/pIr5gFlvLjN3NSdlvHVJ6ZWwlHNz96PSQ5
rPz4wTqDtGWDhk3C0hDJfa6aomus6UcyujqWC8lpzmhv/9U7o+ntut+2ZRuzeSZV
oFOs9Fryhu71KdzjVOpeGVQKyZvFD9tirJxIXcq7PYCLgImojbVRb8UOvnSI/mqt
zWFza6BO+vq5BrYRI4xCoxdqLNJXMFYHvhk/NqaTmTOy384cL1wzblPRDXMwjDOb
BUN9NAdwHMN7gSxovDIfuCoburxXOx4Cl5kCsgvX83OtY/ZmaDkI6O87XOvsYbjb
jbQH2uhZFR9T5E6UO+7MkYUx19O+VWkRdarnxd7ux2joSNAn3WMboKbC+QEOofwX
GCn44Id7v63FpdAKuaVuZhHSeaTebHMSbjnJJEATVsXZcgKuEEnA8zekfvSFWAiF
RRs6/QMtxdOwt+/zhEnfg0s3mZnajM1q/gj1pU4pL6Tac6l918E3TpikmsDjsa7h
+FpUlv58UDi+F3n7JfnR4Ap6ISLahUX9npaBzBNp/kgpq4+27qkpNbYCPWFRv5lS
nDO1f7gPg1X6REDt/qy8fZ07TMsSxrrknd/8b0pJJBWhMyDATpw2Uc4Po1g2l/aR
s4O4Sdy4WmqUmBp6s/CEd/8A8yjR0gITx0k8vNCI+odHM0SmpzrwWZdpB0g2AJmg
HlxIBJ4MbAEwFpxAHdzCUNUgN2KZGEz1BewBrATdiZe+YUC5HA6TZR84Dn+AgH5Y
FFTVV7JWa+tLjV0CrZrEmd+iTLEIffWnKs54E0UxgccxKlBZCNSiG0STW7gjGQMB
lIueWkjKlpdkuMh7DMMb+jYmthorRtUqD6JDVc7bkNfzPUpoVbL0LjnusB3UD5gx
+d+DIH7YvnwB/3sLA49pMkA6TD/6R6bTPfxM57mZGhYzF0EURW396hr0u9aRqDq5
PUXsV3xlEAdLBZbYN2vvT8BM6h/2p2E2zXGakgiSaqjOYDqt16BKV79xfD5alM6X
9xXqBDvU1DdeIlVTnfMAuyygDFjqbQ9ocjobtqAzL6qPE+85o5Jq+khwMF5zjJ9f
dri+W5p4QGTFYM9fMEXfn1OO33W9ah9DXjpwYFbGALUJyXOe/QDJUboLE4HIwuTE
CyN1njhHwLSZ/kL8eAzgODVT7W4aXWuZ8Y0PTVucMzo0GKyv22hE60KBD4uo4XOQ
FB5FBnnUE7IXfPR/d1lm0dhF1f2ac0KFc1J/BSLPWMzp0AK1sa2wvQT49DR4LmHc
iv1W39ZfPF2ZDvmxrTwA7j9FKLLZ+tXIzD2h5Duk7KzXudS0rYFJyOPvtVj1mwII
nzaDNDUJt+9QrUE2RYodYBNBYdkSsQbGnbnOPpg0chvrvLuZAu9wHsqGnurv13tk
AQSxZxhcXWUcGfAZN6OMvI7N0s12ewHPAmObGyDfi0O6tSGzq35qoF65jrWwFxOy
eGBFxkCdvtnZWYbIsIHWF34lGEXCs66Lbx4PhHTVRh7rt2WIQfYToGCDOFkb4bCO
B4xvVAuEm7T56Upv++QKHG61QbEZcn/DrgtclOQKoIh0zNrdikhzCWk9129ZyIay
7ZqOUj6G3QgRCBOYwRZIcbm1cLEfkVsBI4P7yefOWWKOyUS3C5VMOcrt9dkYrFZs
tY0Eypzq14H8pHigEDWA5VeyTBd5CqNMuFFBliFP8V9sVTnFqCXPgfX4NvVW73F3
H/9nPe0yHsDS19+PoDjshlYuf3flazqmUN8YVv57z+BrXQFYdm4m9z+1ht+YCkf7
fvZ8Oz9lGT4hiJnGI+Pi9lWLgb0xiUZ3RGgmp2OTcxcF9zkkLF9Wvtrwzr9QwXnG
FVI/6QAY1G4lJ4dJCp+8AIYdV7sY8WMk+9y6QnnjVrSNmFA7qVyI4cJEHkEDv8SN
OaVdtUG0pOinMeyxh0Fh2rejjGkE1m4fIlrZYHo8o3I9JyhhKpprSUdsb3cc1x/Z
QY9Wd3Qrg5MgWJODHP1PzLaPLHPpO0Sok9Lc71uHdJoBzLNL8YMV5rB1uGF/PJg5
cxQMHX7s17m/BbE4nfdW7ZcLlEhd6KCDM25Fv6751BP4W2KqjYTz0OIzVBXBiA6t
BWezXFijq/vF+A9vwRsZslXufg4doaHAej1niMOIlkKN2WmVqlnKHDMcyB0LtWFc
BRgepYDqsmDcFq8Tv/YcMD78dTFi9r9LtijN/Z/1W2LMdePvTplpOZQG4YhIittT
vayO8DVhDjUSJsAM1pdtIaAxpnSGz6lsfhK1xAAk9FIfIKqtY1L5UdXGuRBcg+3b
QKvvT2PSQzOqVpr8zzmy9pcj2rkx/yrsXtNSVquFCwZrWbcnDtoBR+wiNkn7YLuz
NPKQOP+JKYiSNpM41pgJgFOfFKNIIxBALDFo/TIVTaiw7LesMzZBt6SUuE/xcq/N
dgMUCuOy6NWYUllTFq8WQ+7H9/iHcCYdAmFyMR3NJWg+axHNOdD0hOz7E4wMkeF6
gYnW9DuYPiwfTqG7Td09MinEVS9sV9DxIAAu/6C4ifuupwgb6Diu+uhXw8rItF/b
hiavOCv3yCRt6veQyrH+uVkX/G7loz/NCUARcTuxLhjuhhtQ0cclF09W0xIuu+X8
FJo+y2BAzSJqToH+ULEveFik0KHTkFQA8/qQkqNzbEy8CuGyIVNcoQR2Vvt542Ud
sRvmaaXq+JcrAShJs5zgxz0QyX9JAIkzbyJS7ttq0EIqpqkvErLt50evFLafQb98
xNZlPiz7rDUrVdwu87RvKPWAfZHrdN5D01tL87ZZ1tpOcaTr0fkMq42V/HMxrssW
icvH39X8c8WAomdnE7kQSAE0Tyt8m+z3FR0AUkuTIgz1aR0uHBD5Z41S2tPrKJgF
fdXkDHIYM0DeOLK1/xwCoBWX3/DCPReNktX/h1phq7dQuHsFEkITPIRhlef0Ebn+
aHke3BdNh8mzyZe8X4r7WOwj9DPMhN7yUoqogyCg8wA4m76OGIOCzuo6NaBDRn7y
9zKtxGBUsLdhaRKdo7xxHJUGqvVq/I7h+eue7rIPrMgaOo92jBIw+Uy4dVPvo1W4
X0NV2bwL8hWxukSnbUMdC4NNXsp806NMAaZiang49hB7rm+V1ZW1+u2M3NP1O+xe
`protect END_PROTECTED
