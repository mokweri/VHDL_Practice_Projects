`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4E8jCW27/APyVFzjFyS+UzDkQ2ur6YBswjEYiu7nGubGgkLnrYJ+WoRVbIxV2U2i
mTEGHbf9haJmGWo+3En+Nd2HxpzZBcS/trh1gzMgvm8xqOSz2CCjblLbBNQEOuJ0
kOMtFZpr8eprPdhEoTKyhw5B+coxBmdru+DCFkY/XEoLAxL8tCD3Qdg9IfIP7J3g
UpdjGRK7pVmOElBaM8exJN5AbhcjvdVzbmnFxXXe8294q6K/KSPqaByP0SXo5e/r
X7/VaKIG3MgA/ZFK+azktBkcbHgfScs6XDn6WKb1VdKK/IFTLL/htsE3mk4reYRp
1E4THkQmCZNqWXOQFZhmBTfxkPeR9+zF30ld295PXtJyunh4xGBZuhFsiX0LmJmx
m5BfluEixsnKCM4a42SDbpdIC6Mc5qx/WJMuM5KBVNVxRN/zGIoFwLIECkuscn7X
xLGmGDklWkW3+eMGzk+tuzkefE+qK2S/ZUxXrsS4mqbKMaopTOSWlsaLNQsbExqS
tK73FluSnfHKx5w2bQ9XuY7JpnpjTcwmtoCMLCkXZTWul3jxCNuTVl2+pa4qKfjb
lL6mRSkbQ5DhcTlNe9mM6yK4skKouKHw9inJVmeP2zDUEOqMlxxgKHEAL+r11PDf
pRtEo/eBU8LZgz8scxoJGD1285a4ZKRS0uUqUWMhNUgAaRBYecZKSfYHAaTcUMSl
y3Nn3raDXtGdPSPZ6Yk0SQ9VhwXybhnirgBiqimz8Ys1k7Fl1DLLE0hOXs+BqG3V
M8PtOywYB/w/IZonLBikUgSJtWtHfx2EnUzmLK4AWfA0Jef2YprH7YOjvW3GUj4t
KJhis2KrlQjK7BYfj6h/VQRv2ZoGLbnUyNtIu7lKtsKW+vW/6iRdSY2mp4XM6a6P
/a1KeD2mu8iE9KOz8TdcdBWvOBg/OOKJdMNXuUNw0Ak+WeFNqXWWXx48UAKmOqto
inq6iQF02FyH/TtDsFKILUGz1pqeyG9XBa7m9VT1wf79xVUTrYWvLLZbA4VkfXdw
KGL2M8jSK6NUHqyUIec1raLHf4EqNgyXyhkYP64v8XtPioeUumAGjPzAXljuIzlQ
GF8izUiNCia+mrPgR7PGAHuHNlTVnmL5URqsoXcpdtxlRrzTcVDC+y7gT94xttqG
IXXhyAARD1y0CEKU7gy//zwv6oByvcZaY9xg05T7GBh+aB1LMlncF2//h9DqemqQ
nvmVG9PFSAV2bpV29kqQwODdWTSDLLSuxZoPqhcEyVk6rWZDNlZydXbHT77fSNYH
3SMYceNFiHZtJ8bRNtrdGyAkWNRbmBoR0Wsb+7nh2DBIVHdEQ6QqO3r3eag5oiFJ
LnklBuxbcd2DbWap8QntTiUcPHQx5gjgfdW4Hz+nP70ECZdsVXYIk6Ls/iWqL9K9
xUD0VLHsKYjvPzuUyHmHTKDfML7zzt1u2QatitNckYs=
`protect END_PROTECTED
