`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+OAyuJQnbVlMn1QziE3IoUaM6+I/IeGlulR3/zs9a8u35S/Dtc5+G00Bxmf77YL
uytDDkFs4ws9NKnxG2FfKG0Rqowo9iUOS/vhbDDXv9MjYitHuvTz1W7oTXqjkk6x
l2tigg2cj5N2lI/yfJzYPFHRBr5bDssguRxk2uyw9DFgU32fYENxMejqiMxhH48z
7eZLQnu5Ps/aAuuVMU4K569ZvccARkWbI2PPgNfA4g1kPAskCLclBQ0ppeArqOPJ
91IbWbwBCKLicspVRfKVOh5qHWs8fVs6BQiQQREr5RLVyktVUSc3fhFXHo9zPGig
qH3IJ8jWE/FIfNHbxWhwC74owAiL5IU6SrajHUhDNO6yz/CF68ICagsX6PQ1EGYi
zBfGNRdIunBWJKhlksHGTdE3vzEVwaAnmjQ5p4dbNNJpvUtKMJ+cLNTFZKQJI3Bj
G/LpczB6asoyV0jw40uooL6hY1mXIO7XoQQuVBHbzU4BbIE267r2u/MwYvITW2rv
mdeOcTF/Un70OMDy6xwERAEdZE5qnb6tXS7qvTbyQrYjj+zm/LSR2Fwu4JSaHN+2
5ByDLoSeWOZgvwWo8NSvMS8aYXAXm2EDKeXw1E1ALPQvaF3p+pWW4IgDm2G+EhE7
VKnPGRitYBNasnBkMlLghdLGubdTtX1/C+c+iz0JhvBHEFZMlkqB8CT5/91b5API
lsHi50r1+j2joqcnrX5hm6p18Vl/4sjtrOHLToqwhmobvp8/v1qbZbMLWbOVFKMU
GG5y1Y3ZCAM8sBTofdYbGZkFBgZC/UEhfo8SqryWxbgy5BGL5SXWVzFBJH7rWijo
FjZ95Sou5N8k2EHdkBADcJ4oAH8SwHSxTySoooUmQNWCk2cjL77DLS1pWKrzMtqE
dwUchCTCf1gD2dX7rP1Xg8y2DjgoefU6TjgmGC+bfGmurpWr5M5aiC98/mlA0qwF
GnBKPoFnwk6gY/LBt5SgZ94a2AHfKXyDe2DqRQ8Xwp1F4TgCtipxfQVTZqo/OKuE
iesoCRS1DRsm16TVMNsPm4+s5cTIF19lXQxhanAHTMJ3+92OCx0d6+Bv+ZVp1B6m
3SUjTe9cFUj+ttA+lCyWXA4SG9sBJNLzaXpbJwnE9jV87XAhLke8Sw8sxN5eFMld
1/gK8997b6eXHhZiyeIn71it5/hjvKbmuec9P1zt8aBCYq1MWMRgj/nrLZTqo3+X
1vAlQFT4MQmeyIUklci3slzXmnQh2+uEoY1T8EulzC/tYxdc/mbuAldi6GuCgCL8
M2I7/sAxGNmeTtFB78jJWyN9gMIqG2yTHzIaOvDe/IlVK+jqh8TeRPj3+UA+JoS7
3VysGepfVt64lN3051381KX6LlGW+7ZWcfjYQ2d5qgxmkOQKwKKwxaRRdVSGyBvA
E1MC01KsUf3m8RoORnpZRcghChIbox1EdvXe1EPncTM=
`protect END_PROTECTED
