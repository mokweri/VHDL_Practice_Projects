`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMdcbR8qOPq9sy7TUrR7La5lHWxQycON0/p8ytCfUtXL4gU/Y3YkoNJkcj6mzyWH
Q+vYZgV615bMLpem3LZx7OhbuQDGuk6TA7G0wQ8YcMQYKxCjO2QZVrNtSpdiFOzb
3yMGlhVr7Xbu85Eoy24/hmNfig8hiSJzO17zXQwaxl8Vda4fBtwTALEOvsHNFfXu
b9LFIP9SOs2bNsng4Z4GY1jEafXsRdI0jN4Ea3ZI3xHr2aVbwA8pONRKW3AzzbEe
3Rz69o9Bw+jB+eumebunUHSnELFDPQMcGUuGRTVCQVqbYiqOq8o9De0WiFBDSOHN
Fkg3T+2N3H2CEwqRDCCld5Pe97dKeiVrpJiuxkSq8PP1+zP29QYXqL7zKhS1XV8N
RscF1Me9KNpr6VmqEH2RYZVLhCeeNG7e1Pv7dSIuILqZ2bqqB/29y2+ISnvHlDq7
mhJKeWX6GC2jFpldI9aQU750KI3+IzRoqqSXjX9D9RSi5ly+ptlDSpBObklWClEZ
7p5wQsNojON9sAUY8HNBTEttO40iFvkL4cjd1RAgNn1moM+GzzOmBmNrvH2nsfFm
c9baTsFYD71xBTO47s6Bwl1OnpIeCUCqkahmEGiWO0xwxcI5Smc5g1r+G6WsTZAH
`protect END_PROTECTED
