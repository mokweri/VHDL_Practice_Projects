`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83Uj6ojGN+59LQwA7eZIvWWZEnLXngaIoyIvtycsv6MEzjrrDTxFwH0r5AYd/uav
edK+n61+netd0H5F9Zf0sTvzFAaHYkmFc015vty2YSj75ozzPn/fiISRNrJfFDcD
fbGu4KVOAlq/fL0R3CnwEohcemtf+v/Gfms9jmdPTvOWE+kPyvEzMqK3ATDkavRS
Ma6o45bGqRvpk2wUiFqqT4bJfqMoPNPUb1t23eNaig7EDcfZSDaQdwm5LuyddwpX
TnwvqjY7F6y+lHvx8WcPzgas4/PuPXx+iDWhr4xVV2ZYMR4xDUgw0AaEvzDt1gxn
+3yyrKeWNxFQ+NHbpuG9bVigxEutsyplv3UFOlHoZM7IVpfa/VdtXxiEFLmsqrUo
oqDDQU+yhi+KOauCLExY7e2WIK2+lwVN1SMbJKwXY3WZvgcxbV9L6u65zujgi4fC
FFclMZCi33vBkzbUQ5zM1e0dmnxBGBMvinw3nSVuC0Sl2nVnaUVfgVEDhgE/oPvH
f0mirPCByzL67TidUYKTOxAkwcy4AMdhXWp93bS1H4Zpmz3CDPFycha2iukImMEl
LYVxsK99Fp2ja8OWVR3sP26VDVhUe/dCNKUjeICaIYKKrC4KEyohOaYwGJtiWjpq
bM5Freyk/cxYBq3ctaMTp7Q2tIoVYpmKhdDYLz3+wHDfLwa8MXyPHScqgfk74HYz
pDijdAm2wdfD3BL9NxuUENXxwnIHYU+dA35vpktmGd775gsQvMbSNiVnPweoTj3H
YIU/GBwPBA//Y4ErTVxDUThOGvmilLJLcFtMimUAEQcVIJioFx08tJWLz5mwl5c7
Wtme8Kv0qxop/5DJu8WkkwWL1leI0WBMazVHTU0hBefpAuo0IpsQNIBUSCQsHfm8
rrNP+XLUB2z2hKMq2XiuY/u0iAM2PP7i1uSpP4JYfuwXm9EEtrGd7y7Qfo3D9n3k
erLR15swYoxQ41j7Q434X5ZD4ycSEeeiuFO1ioM4aHFMkljkbH1PYBBG/tdquKWx
A+fnhWpMpaU/jaGgc1ZMx7udMS8ZGutFqTGOerMvuCMcJuHKBz1YN8iFj08Exn4N
kHb1dlZWEruOB+NqkXapTs3MEmtWrkjUqQ3bQBEMex7sKE5wTWf99TVjQqq3L2EK
yK7F77Zlkk1CLiDzBszZXJXfiFBt0+dO5DKk+DusLoD4/rUskcYygN09b9XrXhVK
74C7XSaKbFPov5WgrdnmoYgNi9zNMbQJ76iuj5WMqvyreglgovr19sdWlMi7aVCH
iXzyj1jL2Ms7R/eugpaWEws2TII5iGN53pIZVfQY0KL98vix2PALNHaazHyyMxyf
FZRjq3/U3jeDCVNwxai4a97y/9YMxSgbx4CohUXngehETbLAm1RErZ1kqHNiyhNT
sBAw0gIWj2jWQw0mYhSkGl7iVt0Eto2CwifQUkWvJvpBobaGksunEyIifAeh9/Kc
1Yx1SRIMwxMX6lRoC+kS2VuPb2Y6htXxx5TeMUEukERk/ikNIYarkEnADFNAzila
NyBcuEZOC/ADY6Z20ZI4asrDxT/tNEDUQbGzMmLo4c527JtS6t64xkE9q4OHh3hZ
LTZAaqcj+YKqFr+ipJIkWbdxK03xRGLiC2NEERNXQeziVmVJxk98tdWlLJKXIJ9w
mXOgWkM2fc13eDvwAitl1B7IPYYvB27QK0WAZ7qS4K2W0DLkhuXwL72bNmZhivCX
`protect END_PROTECTED
