`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wSGL7/pvvs2uzIM3FGk8X/K6GvJwUtrv30P1Dmwj+pxtUd1brJyQzT/r15HGoLI3
c6lOWr4ZRtyY8Il5p5FVvQC7byB9xTRcOWXi5JI/15DlIgPn/v+CtVpBLQs6FjYf
397ybTKe1aiID4rcZZcZsYReF0g20LRSDdo3+3b4OE1cW9puxTGZfOJy9uvYQLnl
YJ1OED9ObvKA7Nlc6OJV0SDLAfDAnhrVWpqZLoqd/vl6WAQCiNxtYSAm0KFg5730
uZc99vHakQSFyPMUInt+haLYWbAY88gXUM4YiuqTt9GSO6GA7RnjXemAOCYi6huE
39bjUl4MXMY9hC8YsiR0tilB67P4eiZmTDA1HfebdchUO7o0f8GbTHAPXVKVnu0L
O7QIVxmu0GqRC0jWmP+AtDTuhGRXyet9MrnpenMzUllcWbS2NM41+OmVaL+YXIZ8
qRSrkR9L9KLUlSXo/Dg2FF8ab/pWLqJa672mVw83DOVS+eOvoO83C1s6HPxYtG+Z
ztZbaIfRy/ORW4Rl4bt8jdgSaO2PERxBiqVJQs5iZclN+GfyZCRsNfjixSX1D65t
CGGCre1VzCktuTeXQJU3QrSBZNklPSnXXHQxab1WUOyhTO5Hyxwdi9omLwZqGNZ/
jAYw+hCxG19RwfJjQIq/UUGBI+lCdC5MELYfDNdz172MUgIcg89L1fbiLjRaAsoi
jb/L8dwBEk5Et5MtwVCM2vO6WvAfi0HbWYQlDosZANF6Isaqxvd+g1cZqXihF/pX
F1Sv7Qjn5XsyxUb4CWdNIQ==
`protect END_PROTECTED
