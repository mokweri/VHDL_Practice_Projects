`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g1ogQFwfmFWL07Ojl934yQ2K9wp7SfUvkjoPDXuWcZA5KsWUP3ZV3XXYOeBE1u/N
sytNb6Aop/zsx2cJNHm6U0DWpiTNg9gy9sEdElS+EFN9Aj+XVugSyBliZQX3CxNK
zQaOZv0MjVHjKC19l+A8rehVl7nv6hrARjmFkjWN8r+1Sod+KSw4dC0hBmmSQoTK
ejC2ohk8j7iZH9hOnHX9jMVvCiN2TRqBvqQNlGF3NgODGe8DKhK7xzNFeP2oBfLg
y+ZjA3cdOUWt+j2yvVHW6S33BT1Ic4TZ3DKMqUjqpurmVDLv8Ve90fkp/RJpZQyj
bSlEPujtBVrqJRf+ebvwgS1wz+wzyZKbH0tHxrDv46QC9x5LhIh4YVcKpJcyHKXk
kDxOfLVLLe3ZmAQRE8hXrC/d93pWytFphKXufNFC5AaCpxXuRVUxucmHoiQ/2Dhp
QZjUiY899R/Bu3UgiXXibvGJBNIJUHEPuRwAdiS9HjG28IBu/yQ/CG2ZG6mvT1op
bb9Nf7WdqTfXrWqK5SRHUtDpPLTRZ4D04DwPnF3VF6ti/jXM3SY04VjBVGdO3ya9
DAHV+H6GbTr6nCCAraxs3XAm3WsO8xKH4PwlOWa8K6v6vWwL+bXRgtJFhDLfwLaD
hCUDgTMZHYRN5BfU6adODbP7jSCNpTFSiClDU5Tn3qLPAbXjyMTXys8rF3NvZJfU
GCUGVvuu2hAR9QdRDdd7HflOmaFmUwXysGe8JHuWE/iEm4BFzs4ybw9BcMKRzmND
E+pty2Psw9j2AjpQb9BIDMa/Mwhd0Z8rbpF6oRWqbi50DhbNW8XmhzaCCRcys4WQ
Qec7t6bqhIIZNEW0tAqjpcb48RBpO2iEoC/S0c7y9oZwKcmGqRIBP89OUYZ8g9R3
gFw9kDuFSBiFSExbG1p8HI4QUjTzGBW0zeKkLR5W+lnM+sYQt0JYk0pj4sPeLEid
7lAToIgaQRNDlMMOAyz1ijklxh0gcdXUp0M2316SxvGsiGyjtAR8VZEYKfYxlYxc
wU4agPhNgQqLJaUw6PC6i/orvGwD7+5jYfFffAzdk+zzGHTBTDZndPqi8iYCvEig
K+1D3pP2dKEj8HYNpBEke2jMgPlozJ0KBAarEm0HlxoKZudrhhb81AEEd277Jp3R
mZw4fbW/PcJnrmqOjVSp43pyJAMywUaTGpEFsMsNWLLYZ6nh9bdECDolNoUqfEi8
dUfRzVgfFqRJLvTvl2mqLCGRRuWjwwf04dGM2l5nXUbL6vRfQd/y8vLPmm2w7vMw
jzSjCZBpVNgvMWhqq/08Dyc4/c1xFVS4vhF638YzCiu9/eAOkWL3dvd6m0+bNOpz
Tm4vjfEDozszd5SnKnyuwRncwZzzBoJHBIx+ZHlrndn+J9XFsmOtbvTV5trRr0+I
eDinj5Hmrtlo3Lbyia4xWGbwETBXJj/L9D+NfX3EEyEbHB4QT6Ot8tCxSUTX9CEw
ovn3AWUWQv3veimRZ4NlBcWxLD+w9UXOs+SWc4rL66HQ0Y0ryeuGpp1aSlVwrsLU
W/CI5gG6+gCdqA7/SRH0M1vZTAg+9PxiK6iwqFSwiTsroT6GmunWk3fG5MnBbOQR
ckXpNmcKHIA+TcgWuh2h7c2YSf1Gqm3Ny7wmAa91d3AlMZ/WsJbQvUGv1IVlr8Hz
j/KXqE8eWIF94zBzEPPRyCsceVfp3WSrq7P0qCst96efYNIJnAIlRBtdd0Ae6/9O
Q0ytFHWAIpxwr8YtGigQcQHs74QJ2MCobv7avmPqIZ/D0C3WukBfHr0ZCINuey5L
`protect END_PROTECTED
