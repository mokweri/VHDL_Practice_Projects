`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEJ3JMH7URyZyE7zVk+H6izGZ/wyo4rhavh82I5T1SIaJgPNLhPrxjVZTyzzmC5h
KTDA9J9yjMhl4shevo9OnocbdwISSYV6yHoMkpsza73KvvWoZRztlUAU6GZBvTWt
U+5dcAHyV0TeyVLIVVaOez0iPbxAxLzZOdWyMjaUuxEQKbpIY6wKTolisCleoEU3
z80w7Z063Fw/mh0gp/J2XfNb9yynZg/+3c593jSbwrqfQVfkLF9/mdivhUB61MvM
8pzThPTn4x0i7iqU8lsG3WZDTdRMtJRuboA6Q+U1cHz/HgIn2GhJYaGpngOs6KGW
kIzk3JgNC/RnOoQ5UZNpx9kAqfKvFtxJ4d42847x5DOFha3L/f8ylSKrPaKJ5gav
3PNFE3xIZAoJSQGjJfg4dcT3qTU6i+1JObYIYdp6Fq2KqTToTnr9mWttB6y7n1do
7//p2Q/+flnFoG0mpHfIZOxeqGYM2pnJ4v7YaMZUa4fJRlsuGcbxbWW/32V/ki0f
5pSFDysN7fnmRIvOicxPOrANgu1IspsoMKuN3YeNsGbTvv4PVHnOqBtktZ8DVSdh
tyhJVl0LLNpT+c7SJSd1qM9xnLlMRRpBVpcGb+khbC55PLbKbDeGcurGbE16b5T5
3AJ1hj8oC6MchtEWDe/8HaEK7/sq46adVZvPJQwEIReK3LBjBFOai0NseCKq13IC
OjFJtk5HGWITOUzRSatQTnBlGZN2YjBbYcEojzmySjBQsIWar/+x/HU50FiHre4L
ni7NbRaZiY8bDvOeNo4t6lLwC6nlVO9Ouu2ib7/QWCn9s3xXLssoPHEuUlOu07oO
h2Zu5a9usBh7YNXskxMnGqC2J/xdczuuKKGjyHR/dZLv0zy0yAjy3BmlTYgytsnK
D+FZgv2jn3ZaOtCSwE9TORSJaVRk1n395ZdvmiA11OVTSvfNRp9dW8o035AyAJ8h
/PZ92n0IndhIh3etjqFl0EI999281MrPZu1L31Xi/bgxNvhu53b74VBNkJm9/bq5
7kms/djQRD+iw4mG13ncBE+uoQ+GWDkrx4f7FgbsDNtafbdlRXif0rFn99+cvMLr
IA6vtGuSowh0cBIYH5BIsxd598k9dXDWFjnNycUpWoPJkCO31eIT5cnkqMxoGm2Q
/DJX6LfRB/13mJVkfuPa4E/+7zrOlp7m7bSPy258SMabsBN9q2/zppDBRokz7hWJ
oKlR+/M5IFXbReCvaqlTKJDs+v9bddHHOmTw18kFdugKfbjnR/aG520fPypgPur0
cSHF82X4JTQJAIbHlZ04YMr13aZB1QmqUXBvtPGv8RyQR92rY89hZh2+smu7qhoP
w4otUC8QaSQ1FPcZh8x6bowI5La0nrNcQq+3ntePi0vr8o0axj1AuEXqU6X1fECo
HQokqfOqw3p1yFNwfPvqIf6yDqzocYhdsR0KnDNvchA3np5abnb97eWmAwQY+gLs
tJgG/3ip4UWSIQ2D9EUqekuXf7k/k0aLK1wF/ZYpgch1zMz5pR1oR5qEWF4rfquS
u0O6y7Jy9qxxvAW3hrmPdK2ZovzB/hsIvGXeMD14tAxcwma6Sq5knPwG7FFy0Huc
ul2kXOZseX/76Ee8ESCyzQYQsvrmUCABmicfchKZi+8i9sKLhsCSM/o3eSg6sOwj
scjNeeNw1L10+Hiz7rBb2BgvYe3wd9HXrLMl3ha7y01Bg77P7gQuCn4PBCeVbA+k
LM4M0icIqOWbMwRg5s3KnJY7wMDFzyHVmepWzfRmyP+5Lz2DzmS8zo1bq3qziFS/
v70F3Ct9bd3XJQFca6WWJ2k8kVNRGm2c9PqK+K++HXKui5BBTjMlBNSy5+WFdETW
VWWupETCKULzpBpM6dfJGiOGInx7gTPT0PnZ/1RbeZLPgJFmrozepD+FEsnHIx8l
X13kj6CFgSkMJgAqsczODckYWmjYjDKTaduHgeMS0fQNbWPUujllJ3UB83wVr8l0
rM9psvdQiLIMw2bEaqIEvOpRcRH0I4nT6U++LYRsTK7ajRYqYrEN+wxB38ePm7mY
9VRSh9Q743ikeUHuy15AhE+dmtgnnRbaOlLCuDR0V+Q6pws7UeheQLJ7XzI5Lr4v
MVAqsmqS0T8rlCF3Je2gZiT8wb0mHQTJYURR7MEkQw49WOBt1jb2Mnpv8xFqsKBS
9jjeVJfV3/QwUGCMJp6EFxIfBjaxF3UA32kHmdMBzZQdByR55DlJYqEv+TIg+nPX
yOBXHgNTvchQ21cemth64OiopNC8obt88fzh0Uwy2FhjbtrrVptAiDbK1iDdFknd
QchhERZAU6zdGkAhnLDQzPpG4egI0VgfZJqmaVGtF8woBM5GCDfkEuO5Dm28TegB
tIKG87zLX9U6LgdsXyglO7SbvpHMAk5h9K8P4beuQNX7MfEJWLCW3aez60op4SdJ
KH2asm8w42hEY/GbXlMLwjX6C2iP5Yrer9dmYdAjWjJ+5ZjRZGPPGVyr8K+nsyi9
HebG1E9BndsKLINte3jtO7UfMuDAzyVag0ndSbBcO3acGBJfUrqMbCEZIB/0uSlq
gN/BCXXjhU8euhONdw0SB6ml6BLHUXLN/IeZXPLyG7oJ6NzjzCk/vjJCcsJLh9vm
6syYWiEeQvrPeGZ1h5wgs/dXB4qa1Ktdxwyh5ByhHvIH4GlptpeQpZbAP5N2fT6N
6RqMR5nEpRbdO0ndvDMCjdzI6vvnqDI/R/v0ZPkEalB65p/lfU7ylclW+eFs3bn7
ljAIKQTO1ka5BwsNeFGLqDw/FomBcOwUbgoQw1lMdn9HHPcVHcbvOCTb5h6Q6Aj2
eWYqBBUuqJvI4bh6xSK4UHMVEmVqWe9++bj44WgKedsGTLjw1160bgcePGqVY3eB
IZ72y3f2kxg05lXmZ8YL5mY2FNKUCQa0//ZhaLRbnsridPBXksCuyyCwhIOPzBtS
NT8YnkTq2xk6cpW9Ua14OszLzOGhvLrPst1a7K2GHxJknPuB+Yu6WFEg6HZzCsxH
vyk95ralVEUHgsA31hCYkolr/bHKoPohyFWTbs+9Rf9/mUpz0VA/aQlRSqSYOqoL
LmEE3xCxygdcYnORWl9vIVOLvo7FC00hwS6nqVurxSpvYhSJtCL5uKrM+UPj5Vg9
sdOk0BQgVOXIBGdZWm+YDRhTX9sDv4+XtXvBX22n2134bOxWvLrneELTPWqWFK51
H8FYO9xRP+rHje2pt4r1EUqPMEmS7IMBOOn6E8yX7ep6aW+WXf3i78JOIjvM1QAS
VS4j69OIaK3Gyz3+/LE4B7fV6eD9n65gVu80vZ33PnKnZPYQxc9xYnO6YjDuWH08
JRcBIP4tqAbaSVnCnskHHctcbPFyDcOIbuYkG49iz8D4++CGHppCBMWmHlONknXt
bA0VDJsfI7v5h4Q0vTsYVavAmzXy45cYD2ZOgZotA4lb6IhQfrWB5MQW1he8fmPt
mj+4JfrRBt22zzQQM58JViWsjAqAaDk0uzBxgJPp2LNIuxtT7tKagYnRM6E/Rjmp
keMkk5YVDxAYULN0xMsRthjzAU496yozv+Ef82dB+E3jPISEWfgm+tzm+FS14/Ai
r8kUP5VWgKovmE5tgGXt/T5vRD5osgV/fOJe8yWJYh5/V8YJwviVepAodye5ZgYp
X9CEcRbyrkuCW8JyvSPMB7Vvvd3xtW05BsqakZeDfBYPvTr9XRjWuNtt8oJpuQ1N
LvpA72JP9n9B/Mbv6RdoGi8+hOQK8QM0VVH3zJc8DLl0NOPWpo7RURhvM1Fm+0BG
p6AUDgoFMI0HnN6PHpm3sYO6OaAwojXm6Df0INsBqVw3zgW0NubuejFuCr+ENGM4
rwHK1e4oye+s/4g6dehyxIujzkAEUS8x9wK0HNzmPK+Rx8lUL6x4bWxJGqJo+rFK
c/CFjJB4F3ZoUyIOyF4rBUmw/1yRiBs1lGIJHYBSXlarKE8E99C+7tZGsJ8LvzOT
n6m8z+WnOFy6r5D8fnODaldX3MD1rMs5yzhPgJrWTmvXEXaauI74DKcJmISvbVGw
nRhtgp9kA4DS6nulSmWG2gx8VmaFvbs95iiQpuClEWGBp3CdrRctC46zosnEfFiR
LKnNAs+0d1F+D1MHAjMs9gTvlPWFmYL3qPnn/EoJI7eqHKE7irmWCKBOqxoRwEp5
a5FDqoVb307cqX/rdAXZ9dxj1MhW6EjcZ2dqw8Xf98ULGFSt7lwv8qWA/S/N6QFG
11Fw7v8kTBKmnU5bwfseAYjF2/c01BSRofEei3YxdG9n65ah9ANv7eCIVJUL1kRY
ZbK8k3wqnsYlcfGGbDY9GVzs3SaX3n7Wc5chxaHrWVUgIarx43bck5YvLQ2zKl+q
t8+upvWz1gMSSkYq+F4TgdSAwhbiWBrA/6iZOhG8Vq13MvXX8G8BwJ56edJBg5RS
aCPu7QFb9ScUsnlEPLHRYPuw4QGu5LvBN0iAcelPhqg5xBFTaullUCuF+7XAE0pP
ixSfJYLPM9oq12VuhT12czD7hwvVs6gDYooS7N5KGGBLmnK1CxlPwkdsmNfPrYad
BUaEHMB8wE4j3maly7MWXpWXzt9r5W81L00nG0bJwWYNMJq0fL/vNYI9R6WvwEnA
LCmlhT/qv9N+9QRfBO+bdIwLnHr87JGqkvEjq9IhuxFfYkVsnJ9Wte3Eo40vR3yh
q9s6MeuPUItggLJEimU/LNelCSbIkzWC+bHfjc2hcq3EhOhhoQpCcT3UaEFppblI
/UBWNgL+0VvQu6WuNUrMl788Q70ZSdhrPne2HHC+c4sXLo1ypBpr0DOo7pR0+H+r
rBu2KXNNH/hpNM8u4YV/b34dyqEiwG0nkAgtcLVAqaD2cnxdC32isKjxvovrpVnu
HYuTNxUhBGt4cuIuOzwZtbcUytfwDjLT2I+ILmp7f1tXH9ISXT0XMwnDxPaYk6fa
PyR0HYeX33Y9QY/foCRWaH3vuqiMXP3sAIqBYkAWcxfs9fRpW2VxPOIKFglKHT/+
+foQmHpuKYDVhILNBuDa7lZLIp4lExrDEtnDEmiKDRlPphQWQgfVTAFipTYb/Ffx
eDh4P189bD4lTVvUTHOSbrFzT3Hfk9R/DrcTzwwuIt5UVpsU+3ONCHDZFesJnUc4
lKsly33QFwOr3039eaSvG5ue8JYd/LJmDwKXD9XYomEfMjwY+gy+WiaSXElYo1W8
TFTdGtVQpRkjx0+SrU/PLpNAL75BRNGL6R71/ekcDJxQpd3HKyrvnRO4d62dxzdf
GMzWZB98amwmjDYWADXKJHua+DbLz8/o+xOZm6sBgQRBq/C8OvXoD+dGdMTh10YB
+Svnnjov1XhZ+UfchvmfYYERjlmssG3U2gM0SZN66vFN3rEBAP8pcWrg6xYniZ2G
aYPDXvgMSouxQluybjDnPOvYp9Xb5QjLhF+IvJ67+7rDKGqHKlTw2Cd+FXdp/xMk
J+6FwGo2GOFmFpj7q11wmrcVI3MXviFARMDJg7uT1F+fDefX1uXzdCvBdBe75PGo
58mj6CU+3jzJXVwPaFmYc3Imj/sCbbX6zrILWET2w2ibTADQxXDUC5ZllA3T8+Wq
udwj/df8pkC9ZhNKXH1WnTmCnTdheCAzaLKCmIbnX/EgMwcss4aNvMrPLhUWuKhW
pakzOueWHV0jzNIP3JOsD1DRC0UbTzSPdlk+Db+fJgPs+4uGL8kaDECmOk1rCKqV
0kZbpsuqBy1XGvytH38PWiicY6MYDbZuPb56QozN0iNGEO0iOihJTGgBxTXMlBNw
rllkN5ALysaGAneuP0Ca44HXDgyQsoxe9Y48m+kgkb4x8XvlogEEHzTJ1qgLaf4V
NU/34pGik2R5mHdCpi3siyc/t/GWgOGTwAvuxcY+CWVryo0L4wiwxZGB+fK3/2K5
y3x1kPlETt0FZWu227TcKrPHs5v9xDzzDXe1VtWULB51Ipec0JsJrM90cII5dd2n
BHfi5BKMNOurVfixEbeArs+UMYdwnwGHTlv37s31oyrJgsyEy1thAFWVJ0+rjK5L
Ba9PcYN68htxDIj0iZxuW95pFHQPcj6be/XP8rtzJDRR2wxHZNiFpKRa2OHXcFJs
DhVwGHBbujVliM592us4Ehmg3EDheSHxKiL8IuiE1FSriu/VjOXOVVn80BpIABBZ
Yd0cmT2KyKSakIjHVhGF3Z6Outl9sISK6qJE7Nj6EZ4/psBxTj0QZjnTSj29JIgs
vOWpo0hv3oAUbSnld/D5vDlkogbOm/FBjyfEvOyn41DN+Q0mQ/piOh0w2IV8zDb+
P1e/hnA4ivGY054zA28e/n9+llNVECGdpEzqXa8SKJw0w91QenwwXGnds82Wu+R2
JaP1HTXyrXehTZm5QPsh0fUEb7fco4dhv4CUSfV5d68i0+O4ATPsR79Qlj/GGpyB
BNJRRkGWqYswqt5xaSov6NteXl3xq+Zp0Bg9Zav2kW+hrAqf07w4YoV9BwItUO8f
AiT3St7azLkeFBGWQtDkbrEXmY4H33lHXdQlFn4YEAxiDqK1s0NBcFXGgOliSfO1
V3Xh8dJMf+2OUmHIzAuUqurtxH+aoJB8VOZMPwegrqrRtCfEIX29FBLXjjgDSl4Q
gpcKk9KZ7Yu/RI0FmOgrq4/1zJRP2L4ejdTqUG9FIpFicjy1PaZQt2aS8rl0v3NU
16cBAAWqpyNe0/NAnRxFwCNZAuRW9Uiw/iGTYhpFyThNv/k9d5Fp12PCj8CQ5HfY
NQQ4uThlRtB3uy1qY9MmGAteORkRkWZHyZ9fOVqBT8cwTb0nB0gmAZVI4OXx0O/y
DwWRZAuu2jjSZnpeXjUHgvlWF61vU5la7hgg+XujQHiPlrCDUTvAjonlrH3N+FH8
paRER1HAW30xrUq0Yzqqvk2dEIKhKas+5s2PvgSF7IbpvHSDopggTi/hw1h8o8zX
CjrxyRvBLPYarv9tkNxQz2g08V6xvWF4U++hSrbzJMpNob3v7IMcC51XpG+xIObc
XTx3rZhJHq9+kgskuRNh41IAEpjWKARDoKsgSl+IxT/fXlXF2sHKChv1tkMn09Ge
ZtAt20+4qFxDfLOSgiCtv1MLsN5MvX1kG8qujloO4fraL7ftDq+jHB88IKRe73+D
bSi6TmhoRxR+skvdkvVovbOdf+36osFYzOs8zItZLaxPHA1Wh7GGBD/9ya8fuFku
Z1k93PeO8qXq9XDlguiet2FDJO9WX5lTnYg24Vax1bLw2XO785smgo3u5Xz8A1Gp
wsSkbjYXUygDmSDF2uE8xCtwo0wcSvdd2eI2QukUv91HR6QmMVUKywK8CC6M00D7
u3m8vQDJuMl7BnQgc5yVmMXKqpsU4Upr69fgVhH6b7bdWh8s+PZbYckOoxolKRLc
XWQyy5n0XlMzu1frRxnzG+wMYGlUHW7VbvYOcZXawcjFjRt5Nby5ykvrgssl31wJ
7vhpZS8Q3jSd3lD0hLmZ9GqeAXmzkMmrgypPp/LEX5jMnr1///nU6tbSna7+CpM9
UOpOa0tnpsqtSXQ/glRjaqBg5TlK31o3Rub1QJgPSHCE8DEzAkiZadUjUTcwcO5H
xriu0sKppS9eTnHvBxIeQA38BZNcO0BNb4E6mvbXh/EbrNELtXg6vzKHNIRfL9WM
K2sTe83s7vFZ15YPq0WB1uNNlwDOQf7jhMg+GPRYRWL5UNRjenR76v+B3hwUrtiu
sxUqELLlI9gPd9RdkmqOvwELHZWRV0ov67Kh7MSlZTNu2EbsV4gOW34Nb+6YHgFk
EulBrwoEwCUz0cVTzzn6TkmhtvfHJqF3C4laT59iQBqizNr80lbUO76qVBmkcfZx
lDv3OaY9eN6GFx64IEr+hpwvm9hhbNVzpS9zG4Vk8D3kL/vfu49aJYcMPIVOT6LK
7xj3wwZ4l8g0shBrSkaNGRkzvgck2rA4yhvOsGvl4705TXQZ2jOYPxyI0lcE/dDS
WUQlA2HDaLRhYHjTMHo0PpSHyojqoKeYjpz+NinmF1SbWu4gZwU6+TX18F/4z+n8
JbqSxb6JCSVFYVIJjc9R4zgWQhamtuSUx8jZtA48vh6wQsiEdJ2wxo8dQGetRGxP
j4SiR4FAqagfx3joCOkU5/86sKS4hANnL9dBorxxSLQd50MDYkJ/8GI24SwzXzu1
7ESawJJDqEqQ64e7+vuqdMWGP+a89tbS9OMBtLTEi6+5jAY8qeRGIZeNxxPaH1gf
e51m3X5j4+vVjSuQdD7HcagJaYYvNgnSnW0AehD7slOgXBj/vTy7jIe0zKm6AIig
nHdvxAMTvlDjU7SuL4662Jj0DNW0ZqYTuw1kIXO0GKHuFHDAXJI9GYJ6vQhfsHjv
15OASd1GIGT827nnQ0nJAR3QSkS6M1fhmdTqk48PJy8OeVnJTNdrO6ii9x0x4gm4
BZft7qTjQGgJu6WENO+KfGynWGyWlMaJobczI5k7jI1Qs+59e0sOUV17fa73KGUn
poP/Fr+0BP2yeiah4pr/CyIr0yF7clVyp7cVMiUijBOt7akY1uNZniCZJncRyZ5Z
BpP7oIoEJXqi4zfU+xd6FjKRuMJVPEmeC3NG7zz5trBMG4Zoc4WdkONcnC0Zq1pX
CeoB0cutKHNhBrdiyYuYkYArOG6tfuQF5l4aPEU6+TmfG2cIKeFekewUdrHAiUEL
8Iz24hTvp6K0kPH88Fq+Su0ffNDjsSHpZWhyl71WjmagptmU5hVXy05lZBKi07Mj
a6evzLDxOBiBsaHt/wiMjVSJvTj9dN6TbTcsftCTGn9kOAcOaULWo1mVyHJVAuTo
boFV/y2DyHp62m9Vodh97MyJDf9ZFt/jdqumOG0Rf1YSC8RSuImDdIl2X1X81Y1r
PEPXraW26C16kGw13LlokBprBpDZ/EVryGAK9tfjEDTyODw+Qs7Zlpy97vbXD9l6
Op0UFmQOvmCWk8wBGmnB1OK4H1AcWl3ot9lC7hTPZs8AMk5QlH3fHh0RvbBxN91q
cJsTcYqePOntZDci1o4m2SfUme5/9f+TP1ReWfK+7nhMboDB6U5tRT+SV3IOoW65
KCGT4vWfd/Bw9nBHTSBAS14vMBWmEnJaYZ3M6aWlf0hg9Hqtb9DZukdawLKVGnzU
eVzBxZZAO/d4x1x5LZTW9Z+U2rW/Rkn8ghpj8CDPc3Nxgdfdl7OuFJFpJrUrwpb7
L5gvPFdrg+hRmepF0xASUVKCR6/C9CoF9g3V0wyLHvj8MivoCXHc3zPoEg+Qn8ud
QZfd4Fx+Kf3bBI7NXmXNlMl9ujZuRdfBXbntGjDLwDZrygfZ3QWEHYT43TBLQENf
+BR9AE2lVtc8/lTMHjRwZ+xuB7sVevlX5Bz1JgT/CFtv20lI7NF2e20wkhGq/eiC
qUBdITYdbmWjznyoRLMC9fjEjLHiQW6ash79WKvdINLo7TpoNpqbYf6C0EgY639u
QCjZuulJwEplIVKHdVybkdMMaemg3Y+8cYM1LEcFMWc1xg/Fa16CrFnIuLsoiJrI
dM1YIH2eWn1vpIsLeQS4Ya+BWt7Gj4UzDuyTqVcfO8iI8yIY6LmDPy2YdXfCv5nY
Avy4dcdUrsIm3MGPVaKdBBiWE+RqFkwZkcYCOSJfKMyW5AajIoX6GRIgxDl6kyRV
r2N2lH6nnDPWjP1/bhdf2CiD5AU/Q2w5W7VuVK038L9SfumumnVtulQp8OYMbfsk
eCQM904CJHBzamE13QD93W/5ubbxzFkN6JvatcKu2l6smXZLjVoDQgOxKlMggy/e
f1bmEchqE9tceJjLuGBESnePGQfAgUsyylTNIubZ5YHHMIiCnjbhotJx3grdG8m1
2TogtoRVbv4SkLXYbld2DZu/+cgxp5HU6/nQdr7KY0p6eG/FNCR7XXXnx5Iqpczw
FKmWjYz3umqrtbB2NJtNfya+eBGUlPlUPlDhcv2x8FFbPFQlbnQSHahMMlJpPcqs
0rrOjqEnQP8Aq8SCrnagklxxrDvoWut2Zq23qLax9vnT9xCRt+iX122tfX+jGM0b
cnONaRPj8FClUR1IX6TbYov0pyi8249p65I0F0GaAxk0nMDUbnPN71wQjX+s/Rrb
Krd9C8CGDVNHHcKeN3MdGoQhQ0g5xAczxRUGKNyBJV39cMWenxCXj56LglgXbqV6
3Ztb+e4WRhYhWcFznX51w1qehz7YnR0ZH9PFRp34NLTL6UiHyMFC/2/RaWEUlbXw
5amW3rN6EazLf0Bc9M7KTBRSD3YnO8RByqX7+zid1ODKdmJLspQZDgv7I1B28qFE
1o9w04plNgLUsx851cKBQucPZWCfdLvkZJuffKHP0YJvENuwfvX9Zxj3dp5j0IB9
TTocKcS83eecvb8i2NyHhPgqDhjPFiB0VXgFTwVS8x1isH86lebv4qg6Gw9pd4vm
5mtxGTKRu6xAaoDOOFsdZxBzqlougYNTN3+rT7fjFwUZUVBA+QIwyo/d//q4yOU9
5gZSlwz+2zDbfP8YD/fmky5IsIhZe6j6HZfneR0IeEBmApjXJSiXQ1t3/Cakz/k7
33u7afKzZafQyCU8FChbZrPjHzAFVQXVM4P9msJNqYN72NHJ1h54lvDvHfT8Gxm2
oiIzIPcRUxGKV/ZC2u2DEFR8qDfPbG6APjWeVB5t6Lj+yk5GA1wRVSzaJXR1hrXg
sS7cgVWZr+tqQkdE6UXLKHsNeCNVmF1QXhKZ0uirQF4hzkD35QmuCvSWhxHHC9bQ
59Kw6eYzBplgj2JK+xdGkW1OcdVuti7zhFga80/TetBmXLe4hU/Ju9hcYn2eEkHN
uiQAc0J+fk1so/A677+y0/QdsQP+rAsbpl+u+teAexLN1dy/T86/Ls6s8kEA45Gz
uvwEJZ0Biw2fuO9w/V73NK6KtcWCVWF0mLHP+PxhU2gFogfCqppxHrt1skxOhcCt
9GwlPPiOlR/lbIPMrjW5HFxRQijXfuZVZvcpps4WT6TysZKmtRRYaLYeyceEwRr3
zeyO9QQUnE3H7YjBqjBFsATdQJ0ZFJEyv60dXsPT2bPgFX4hCVXlFSGYc6AYltiD
Pma6J2Sh2zR0p1+Nj0zJnTD6gHUNHS83KRvN27irHlhp/3W/DVBFb1BtFa/eQLyh
29nTqiPrqKvHTWzl99NURtbzGmAZoXxB9kkh77WWSBwn6q4Ha0Lf8wJhoy4i48wb
DccUAlf0mr68B3E1hHwCdsw78ceh+VThdJ4cdYxjynTgJgtdcICfe2M0g5y73/5+
rRhS6erj98Lb5c80J77DLZoF10HBO03ga2fckoA5KPI0gcF82d33B/BDb9I9vaN8
FGNTq0/2YH5hTGAKLMzk4CR9N5gj6p538ujIgb0ym884BMfGkqpcUo11j2/14d52
o3KC4gZP1YR1WVPqXDSORmtIkRZhcTu3bFE4gjvZFL6iMtmEzCRXMqqB+Mp9jcMY
trfLSo+hG/UfjNYnqrAgFpc3JfRC1N2z4hkSlFq0FvFfJqJzEMDVU3uiIqAAdIe2
36+wTguW7DAbwMlXcAv6/kJX4vQQj/aniooNpfddQ/ldz1+qyn/fLlNkeqjdC8bL
XbP6Bta0muOsYEZYStivlMRQ+gtruob8pQj03YuP2ZyAXsJJQMTrhsPPNZitIQNN
NcZzys7yPJJWzAqYm30C5hUzrC3f4azkUOICUtD+qaRUwVyhnrlFTGBYgktngVWu
TVfz5FL4EcJk7YGNOR9qmfVgttuu69EYMvAx5lUEOPEra4WSl8YEjq4Rzv1Ge68p
4yOeh/5dejAg4KOg/BGbWYofTCJDX7lNkbfrIMG0c5QxyFSXZNiWt3+C9iLbCHkl
+VckMMwlQQVhfdxkURYttYkiZg96+sIZEUxKVp1gRE2C3TXHu6lu+jVX7r44buD0
+luco1lVDoV3cjPSsOgyb2pVps/uJ+6PnzwOoQzgS7lspAm+ovvIiMBVRpMc3JRU
vmpRfPUkJg96pmvLdBVi/WIDjX93h24LeKld2lPn++aX6MVbnYBLx3pM8/q6qK26
c09CvbJ+lW3pwbwMYgAtRoenrcxk9RIfibtLuguq3NHynNPGsqVH2VINK8XKc/xm
4+/zuNMdkIKG+M8eQruUIiE/1tq+JOX7lK16yF+WozOkGFRlpZytrS0gfOZB/Ac3
6EK7jCPmRaA+VSLFiaZeBGbVWIkLImZOOUnb2i//apXlpPz04cCPFePvDHDBQXOT
6OO9X/NlgHuJ+0gqbF3p0CppPAn2lt+SoLsbAYLKvHe2qRBEAMYnVbtgmitdYI8G
Hk3qpV5kTHVnyiV/wC9flkd3LIbz2DyhJp6y2Q1vd/T5hSk57GTXa3EUNmF92jW7
rU4vjgRL9Fl0g8dDlhsNPOVsU2PZrsiWfzO2FL9mDJLbr91RGXIY5P5RLmd8iq1F
qrSU7W5G0JSjIbR58GV0asD66f9ur8W2yXPK/l5Xzm+byPziRU7e8IVg774Wzvpd
1xEYApQtiQM/hFtpfeAHEj5+rgMfYdfYSPuLf800AHQeIShi3A4aD1XHkFGpXWIB
VWv4NWEnxkWVc0ZR5/TkfRVi4XZ2s9WS4KGiw7q76XMni+L5qBzs9lNjffLQDwle
zsTbqYwX1fdEJ7wr1trqMoy3HgxLN9d0O/cqa4erfKbPBGQuqL2Qwd4//kPwOtAY
OWzEl2hF1fMWE0g/FaT7lH2Vmtp1Pe3MonYBU5kg4IoB4uuVaf8WKn/XaIBTDx9C
xuKyouj0KBp3kR3l/4VDSse2vfqPshPtWYjCTiMMRM+DYlU/BIjFBM6Ubc8dO9xH
0FCkxWtEvvxc40oWHdzziJ7+8lGxPDXaw4Uh1iTHdTcXKiR16+9hz0lRY21ut0pq
A01XBrdH/mgj/eYE1lF6xU1xLBYwrK2cAFsQzygKWEfyLnVJmJ/wm3ZVmFY/bsRO
As7C2qLhzYQFaQFSr0zK97dv6NBXL4GYHRX9CsRSjIVVky4FMe0VgH1MoeQ62ZrO
Hqrjs+ZoaUR4A9VpdddFT7bhcy1RnE1S4drreO2k15k8n41OPg1VAs7XdeAr6DMG
AMdNTg5BV6mAr8cLc8kuo/guDiM6Ul0LEi0uKmsAiKU197gNJMRYkYVxdHmkUwvS
+epYbQ8l/eg6fShC0YiCG+h/ZoBE9W0y8ApTAu3U1mxEj5CHnbQ7LDAY6OGamW0G
VoyJfqdHmo7D320AT+aD3x8CJxPwyp/My1p4HCSOWIpI6c7IffnSX74IHs+bY4p/
N+REZDDSD2Pih8OkGRRz/bgaYTB8ZAADUNxbxzz2xtUZAP8vSbRj1rZFiTiy1uD8
2dvrcr3fSfiopEDzDRcxqL26YHXG35iUKiKvpcoUq06w+3IJBKeYyYU73WAnqFPI
85BJoMI2MdO6nvLSOptRNa32QKxcmckiis4mI/i0h3bFlCxVzIuo8uxvVrdjeXBy
WrYMUfEzmp9nt52CxYdTN6DMi0faGNwDv3tUBiQ+w1NBnH2RAh9wrucerMKqkH+s
k1Ltf/zMOxTYwu26bWDemJMcK09rE1u7J7zaeHF6nhKAb0Dj9n6TulxxRz4eyFxK
9ddn+A20WtdQILLl+QRayHCD6E60pLaMDXzTEKoYmxbnEJTicl+uQH2IBVAtj1Kw
YrSMjTszR4TCGF/dk5EPc414v0tZxpK5y/KEkNVYxgeVKURB5JPG34Z5YMr9LhZ0
7ky3clbjf5oThpULA9l+pnFNjG0Q+VQvcQcPt7j07f5Nrd5Re+7u+7+K0wb8hzsf
A92ycX6NeLoam3DuyqGlfJrwxWnADAHS9MzJ7LYaAqH3T8e7qKGcAOhtw/qAaeHr
aoZWE8MK9GtT/UUnYpDay3RUDzr2ZDJWXr0vSeQMYe85aQ+i11YyJDe3wiOdXLJZ
dzLlwB3uTyMEX5moyyJIOLlydYw+8rTvpqZl8oCNBO4HVYoHsAliJcm1lBD4uaJn
EHaztYjmghMnQ0aN2SbBlRxgr6llVLQZbx2V0BpkQ7btBwOg/iEkUTRuQlFuk6wo
+g94Seu8nWeR48uqiW4CAFzRczUwWvGBByLXkNb9n7VjzSXDBPUodKqgSs7RXJ7B
ujI6zsHjW6sipKOBA/UtZCnKFLmZbThje0DnwczRckLYheqarbIESKs3Ew0ITjIX
dZVnNoaM8bginAxhuNZ4gAwlQ8yY+8lmEyzZMyjMocHqAuBmAPlBseXVm8e8q7Uf
BiAvRV09EJQMfxaY3QYQBj6Fq0YzayunaSjby/9Lvyj8KU8L7/eHsm3ylmRPyiRe
DELpWSt+kuqzy5E2JENZ6w7YYJnAed1gLSqsq0kYe58st0QwyJ5Hvul2wPyIBWCP
YB1FLCSAWcvx2WN9VPlLp2SNX79e/xwqzheGj3FcNghkEU6507IE0P8tdLrMzJP0
fDV+eFuP4VqOuFNR/QI7cfMNdHvloWyNH0NYopbwGY5z47ejNGdHLEvmfnIfCYPC
94msYUB8dX3XA+4Iu7EwrVy9hL3zd4ZFaecADEL/66kXChrD0GSzBJUwFM7gapt1
yDILqxmZkgR0GZClKS2as3DSKXtIejOCZL/XUOy+CqsAO/Z9jy+X84ATLMFFbT9I
I/HbhPFxY1aygnGhcTDjkZQVF9DOpMgdpE9GgpFGNmqLMR5Y7PdKpxpgJG8dFzwP
95hk8HSf3mlHOG7DMpGSSWaFDZmcXVdCV9NHSomWlsPZ3xPoJGq04kzVzz9aVGnW
21A+x4d7ArVDdnz8svCYiqIf9V4M7yxiOokq38fztF9CmKCMF3CIznkw7Bt47Kq6
C7Kkq74nqMWTMlmhb5ZCRxLC/R9Yo805YqmTEkwpD6vLYnNdlryRXTrwI6YTtU3u
Q4513qGPSA1AP04agAJrx+lMEr3LtpxFwJSKs9AzZCGPGHCJJO6VqFezl2loMwvA
VAZnjVm0FyOvlnpJ6jYQu3kN72geNJJ6kOZA8XAQ0mcELIjRiuv7Dv9svaF+hls1
xuRh/bDjaViBXIUT7OVeyRxA7Rm+NfmkgH+sUVjC19km5WGEZ3p+WsHfIaTOls0A
+8P/kj35cWGnu9YhfirojPm0JQPHl1DlUw5AC43HdcOIW059lZvkg/9rQIY2ekmk
Kc9YieBdU0oliNttstYx1beYJhYrLdPJvDoIAcaGzeqRBvqsvBEpzPS/VJSsXf/Y
0CdITm4Y9a+YEH7tObSbPnnJVkbgO2uoB7CKHdc8RSqa0q7xvTYKO5Mu106ehm/L
KJvkW5+Q1VV1YrjHw8stY8WqJmQZNdsgWjUTO5rV3WBHEWuLsdBM4Eu4UCg3mqxK
XuoXQpEoPWJKysCbtPx+HM69jEmywtGQWwM2COSkOxKizdIS+DStSmhP/IZqGyID
yCUogFk8d/CEiuS5Ge5b3OykPxmjAYdWg0kFe2Jr4zHJfqne875/Khkgbi8HchZW
cLhudC/4b9TrCcni2qLx6W6s7RU3y86bk5BTmNQ+YSYPSBOnyuixrhmf13mza2Eb
kmR20olaEAIHeVZH8nzPAy3RvQr6BFxh8lwAGbEwCkdd9SlJWu3b8swyjruMJ5LP
aLTRxTTwdukmHNRCQorHPnKCJBr/WxLuIeh9iHW1LM9l5QYTzJwfgFGmG1+6XS5r
kutVX27dPV/T6k5W0eBk3T9i3FTbtSpO/m+64S0eAKnTflsLixqKqJ1FZvTlTsW9
wlZfrKyUwxB1mmrkR4jEVxLzrPzWleXbIl0duC3qbBTCJOxdWrv4BSGqv1N5s2qK
qNejuQ56BgTG/I1x86aaNvmGy24PMgyqF+UyQOSh+UWKcdsdll19oMiD2NiKlfpV
snE1aHkBlJVJP9DCL6WabxHfdnL2vG2IvFP6Rmzc7WgEadoQG+akUNLuxcS2+Vid
d5jnZE3kybBsJwsJbsfD6BbTm0mrov9qM4qsu3eSVUAL1T80XLKxsFHxXQgiZeUx
QO7F2Wup40UeYjHw6zH5gkl95qClOuVQEYttxwIBrK8Ro8UQDYPq66eR/2PQ8fI8
SIRpXfYuaCuWthTxONZfSLMLnJ5wiJgnRJfjeNE4J+ROYwYeKF0pbAfXdEXL4vb0
J6ankQitnSC4emisFvHLsR6FunTW29IwQxpHgZAujfDSW9KVeV5yKwgsnHVlINyM
iBwpnhs+4P10sBLM/b8hW6UTAZIvZVtC7qsPCxyycwW/9fLa3j0xYVxDAfFeVf/3
Ua3S+GTyrfNVA0Vn++CtxKFC2UG9veYg/T9lc171ewlxsH+SeOnLtC5QN54/XRxY
3VXGXWwwPUhq0hfkdMn+Tnx5MTzq6v7CmSpVQfPsr8g7eL56j+Scm2JbHCigWbG9
8EtznEVo6g0yX8LB+lS2ryJ9M7uaN8BuirjykRTrPJvEeZKJGiW0n4JartfmkABJ
I+iV9mmguvtuEr4bJ2e/csvaaeE/zNjhClW8S9jvSExxsHAhYI98FD11hHmhkLEm
qc1Fb1HQofxmDPBEt01XwcdnGrb4TD9Y5gqtwa4q2YkYsMBYLeGXseDW0oJsyHwV
iZ+x7SvMcvRWmdspGQ65dm2KsJZycLTsLOpPjmaus1B15YUBbMa36WqACmTOjtAD
EqQZecoos4B7Yj1dUVfSldVEUhPW9bd5ydSMhlbW+rRQSG3iFNo3eb66e45Wrn98
q6vkrd4QWVMoWXaTiMRKf1N8j84a0Jew0scKTqZc6hdxNV7CXFXoOC4iD7mwedQj
ZuYj/eWXAwhZnRzKothpW6kIPRBErU7nKiaWCeq+zDsaI+88Pz6w9GcvVeVkzEsn
AQHJ/P0GdVh8q3uOeXNiqVJpcnUEXlN41Ybnjmwaj9Thm4weydtz/g4B/FTFpdiC
MyE5iXX3+s8wXWv5oopUyLgunIvs5yYh0AheWIyuA83aL0q8X5Bo/E/AKo5agltc
D0MnGNhIoOKRJUGdRkzhfW2Z2xmxKwFZYyAdQWKctTSxvBaG8wfryfoqPOZPlVUe
t6DXLY0LoO7JGCFbIbs8jlk/Zv2Yalpb72VXzlLMUOdc+m9ujSXjvX9S6Df7BjoK
Q1Pa+NNAEJecl5lDm/RcvZDMPmjJB2uMjeVDLtblUk4s5rRj3Hl4yAGVFXdg+fVV
5FngCI7hxwEzvxFcBSe4nE3HbupIXylBFbwU+Z+tT2ZScLIWOX///JJ04HEp3RPz
i9MyhlDjbPTqso6dCYMRbcb3rE4E491O8mb0mn8GxyNxQcGEa1C0aIAdJM6M3tXe
Q9SysP1CyqJh8RU21duMjIjw2jgOcGTMeLe52WdDOOwOua/JoPHB/NiAZAjt5ihs
yted4ZO8A5mBvupUZLM8AVJjnCcvc7O3Igw+5eXmdje4kHha7SlX66pGXJWdoxl3
/AB0bT8E3XfbNsqXr1xvjUGQHovRnNyxfvzT5ltd9uu3CDimDe60VEIueOpaLF/J
LtP1r5+QlPzJeqkqA2+f1rHn/dTD1VmdjCNoUq5UNzz9bs/cxoCYg0F/qoGbM7qu
WcgzBZK7LQUpOT1ELRjfigdQkkMO+HjIkUnUZ/PjAvIZYXIpB8kTbC9zymd2+4MY
LbR44dFqBKi0MSZcoKNBRFoGRYPYuh0i8c7fSjLD1HOr8zkOqTXs+9isb02czKtN
RVRyZWT+9D0Gn+wDzjX5LvDeEQ9PelS1B/KWxGMFBGEurS+1lezDXlEYRxIR5HCg
3vOKYw25RhcTy6/oQbxE8XpXq4j7NqwpIP5Ge6oYDFjxQMsRbG62aNwmxfmR0PKa
ib7J5smm/5Jyf4yM5eB0OIconqvhRGaxk6P9d4H2amXMOl/uf+Yi3SbKVrd6bgpE
qdlFJ1Vv9DRl7HRvd5rL/ErJidTiU2ANpgHAmv7yhS/qhxTozcrojuRIcaIygxa2
/tPrloKBec6sFutwUFxUowuWluaSWCtpt1nsDrBMAy3+QPGSI8VELMYrT8+lLzRt
kqYGFj7SnAYCy0PKWB34BYRKiTzF07eidYylRwkTx/x1iOQ4CiUA/ydMFt8Ab/OO
oE4RFfCOu2+qeLaBOSMuil0Y7hQ7jnc8VmNKXauALV08SLFrjtwns+eTwuP1S2di
em8Gdd3vTOw1YjZbIdkFV50kiMC8TZqAbtAXn2qddJSzmjI4cP0+hejhISi8el35
IVaDI/kVAYuY+Xq3L3jomo3QWC+b14LddqZ6t5hCFhzWHsDKSvFmeQfDvh/YB7dO
Y1o8+SifAC+TLj8f+DogW/4gbuzwgeqaLedXWfmvBt57ysklCzqQc/DKngViT/vO
nch1ktV0gOHAsoZcnRRJQf29qVPmEoIetrdAT2+h9qvoHsgyIJBptiIor22aEBGw
8JF1i3t1ulThqUWCE2E0Y0AveRAuP8YI3YrZXA8ZxjXMYrR6dTlcwxCPhBsAxoxB
8a560c/oU1kcMjfH/RYzQQQKJgi8LTkOTaCTff3RN/UbUUx6uKjuLIvhXrFHB3iX
f3KhNE94zbdRuR3x3p1hbpOgSlib+x1GUkmWxiD5+sCnOhAdRcVodS0CqrX01NdL
npcQ7KNSEP4gOh5eo6G0CenMkANppQNp6yRGJGGYpDBAiMnZcGgvVF9bKNyMlv2P
sG5pd/cirbxio4xNDimZmPcKY0II1WoSeiwZpfqSn0KF5BGoLavwFma+T43Xdnzd
mz5miAtaypfFJGaIvQQvb9tocjWdH/SnzAu0h6yVylvUy+fB215NERP2yOWmQVfY
QPHUnr7BVj840l7q/q+Koth121ygyi+di8HBc+l60DFQDHjcUsQb//0w3ndBsTE6
A+m0Ax5eI7oxB497+Cf+SiHcIefo7Fk96tYEAM+M2zHMTyohkNL9GouH6NOYfgmH
RWpK1JNk2Iv5SAF0nKLy3NSlKxPoaXzEyQeARG9Pi0I9Ulhk6p3+Tv9fdenWACkV
p4inzqBajWPPKdlbozWs9FQukNodjWm9bv2LMJvTrPKzUjdXw9xPfPf7AYKUa1XU
NXg2+qQC1TjH5bMkWTc1GrsPrM34S5QkXjhjGZwq4QRh8H4G9JbuYy8dKBzb3ZoJ
cAu1D3TdQxmdcoBSEC5xTivE5ra0Y20FIACPBIEXy0LzdnMvPWqlWKVQQMlzdpyq
dRxExkXrouBECT/c5y41QhlVenznGUibJSwnIBbH1YbyKiE9jnvNalg0AJ+/61qU
I04j/OKQbl75N4MJ721f/JplrzqkrQYNpBNYhdvM1X4rH8vM2dXSHFtBuycaZqT/
pvtSupATQk7pGzcxeMyeIUiixOdNHS5+k4Zk72mVBNSPfAjKN4tbgQTWJnUaCQ3U
PL81he0bHWypDnxPXyqyKPgw6DVE/MlnBRs1WehGnjJVAZET20fZJlmg4wZkNvMH
uAfYDtByI6O9IY2XbCmEP2oPzrhIiJtKBv72qb+Qz1RhIoL/4Cjkqd5V2SmD0KKz
gDgQxYWfiEq1N3ThARfUBZkGbU5VUY2k5h6gAQwaWPJk924AGOCiL8gF28JM+c1N
Iod4t202uCIpcVa3aW0xuGbj/gAuMHRhz4XVygMmYIn0mS2W2y5DrcvIq0Zn3Z5Z
2MvGazhK/+/fpLKUOGjH9vpCDpUjPiLFTyPhNitJjlqKC4SEYVMsx3HIzrH++epk
6sGLJODxOt8nUHA40Oug7c8DEnw4Rw0IkNHLTXkrgUz7I6BMt/mvuABrdZelvo8R
YzfAL2WUi1bfP5C+WnmdPyU/X9zaFWJPPAZEnEfGTnKZ2ZPzc5mViCM8dkA8VnBM
+RYdvwDIwZR2EMHRBxIb9+ICiCDBVPtbjmaLndjgkwXBlfBRiKUak36bBl4qiFAd
7c/oRD/OXVzwMNABLeGvJ3s1Q6QzcJtHdMUarPSXEYBgUG5/7aWMWwPDVGL3/H48
to4IG7lE07ZUgXshlr6C4tDZAp4QVhcNym1MpCf6bkycedeALs5yBLORzgqmJFoQ
zJH8wXmMBEjta6XLOs0va6Ts7YEc10SjJXoC5fEvU93sOxzXgEwx1lhocUNf9eEo
K/DzpD6ldGDXKdfH9kAO6sSApz9VsVcBTY7Vg9WSwDVwR6t3Ak9F4diJS2hGvLht
PdSYlFQFkOk3Jm/bGFna8WrYb3vfQh04+Nz5Wbn25GqyLwj8Txx/UcFZthj2IZW6
cJuYicK573a0pXVS3RnhKpU7AXvEDZyahlCRrlL9DnUDMsBnrzP/0LokomiWHii/
ROYw13/nH/ChnZZ+Jt/5HygPYPnEzgAmLZ6d4B66zgHz5DgekqW/1lB3b180lgWF
bVRGbjf4D/9Q3HJ9j3qK0OnaBAKZp31kyV3pzYGJ6F5We7scudB3VoMWbktKWjgW
Pya+M/MCAWNWa7DskV82P2onb/jnbAKOXpuvsTAzTCOzugtAF+bfjWjo+sNedhDp
3izBJRFOe5NL3hwOVnQV1Lhq2l55XX6JoCOnzJpddNV6cJlLh5JCdhwIXrRtvuXY
kFsjBu0seHrEQUcmc5tSuvDFs5WhwrLyUfgbmYxRxxnGjcXnLgrJ7ZpTRZuDnhYc
UVzAKkThS19PJr4V/mIN3n6W2uPzEJoZrMMMWZoVOCbcnw+MlfNJQ8egbmYvv3ct
mefCRubO8WtT903TNjstTOrxucsmUgJ2+c6KAxNk/0HbtqXwh0T5Xz8NHpot8PbH
dIXiWFzFB+TpBQIEFrZQ47RbQgqiIgW1+F17Kf5lHHUU6etC3Oo3ctMaRbgPDAAl
asuQHHJE9Y58PaUIoy1Q93lMrQMYhh0euc8faYuOHoYbIT0Df2NBtX7P8Jng7i/q
kdkBajxvWR6rrUDxxXNWq1Tz96DH+0XM4/6d1EMGbjRjecYGcYACiaPX14N+FyeL
DTFsd4TqsqP4eJ2Ri2zk2bvS76uhZjcMmlWfPZST9+96DBysB2FrU17wxcDdohtT
6fUE6p0li33eJQJFgh298WzaJLdKgWVEh4Pr+6Cl5tfytWJD0uvHhJLOrgpD0EhZ
SsvwQxDk4iOwznV7aEVZ/FeQEy56YP/q/T0qFiFaZlGu7mXwnwbFTUM5dNuRL7nS
ovMD+rW9ruKBwz6TaMQpAzdOoccy4ReB+/NqpSQPWv0i5i7nzwN7VW0u682D7YgU
3f48O6WUNfB63BbZVSR6aZPQIxElnvUNMcQdP/JTlou3v/suwr11bImClK/gsqRl
5AMQhiiVqLhtCJQqlcuo4nOHEK70BQ9XnMeyNhkjdok1yull188Sb3E0VYXZS4dM
dOZ++aNQ5bZOdicIz2aTxnrvPx1MFFFfVJJs6JVIaWxzqveRvXbZ7iF5Sm7Mrp20
w54oG5FhiiITX5UE2cBeTpPrzDEYPxbQMY39Io6YelSIJDInPDaHjfK+84+1ikIN
YX6QFaHLglnXtK6AfMJy4pl6yMlk7NkMINdcuyg9C1u1HCH4XqmCkT1o9fv7G+Gw
jQplPOiSiSmso4kYhTn1G/1TuGxD6Oc5YnR2Q1OghWZXxO1NHd3h97MiWVcBHlkC
D9vzfol4E5f2MdqWHsGnX0YqxK3ALzInPOI5+3Wzp04K8Bt8I5lr3wZeGQ91nAI1
HqGymM8tpmQWZo+BHJwcR2AlBTLl2a2hC6l5xCZ3oZBE7vsiULU3uQUhhodkxgGZ
DjPQauUAELVXwHkn21swmYOUqqN8wZ3yEtfzJkXyND5xfwVirr/+87d9ydPz6r4o
PcyrmMG2ISf+ZWXV3P798AnK6AeGFYOaSDUREq9f9xm0Vx4TgkCZhHLKKDTHo7FA
o4PTuY2c1elvUJ9otZ16em24BB4QqV7vJyDa8so8Jqiy/xVtPOEZmiBYcOKeQ00U
fjexZxBl4Qa+z6v/GJUgp+2p79r9RPVCfB9/Po5PLynTnUqg0uHWY5ELUWXPAkMX
4Xwf6X5Q0wa/nUkbpp1T/VzXM/JrGVGj49JsPx58QSlqFhgFM13Ey0IcaFXSgohT
NQA6fBJcaXhtM6Zdl0xX9O4VCuRZ61E/+Qirn0tIGn61GndM3c+Bc66eNG5USSbq
+a/P8Pn2R4pDvhGomuLKsB0HGG5QzTeddk0yQxXyJ9uMXP1Kzrt+vC8CAssnOd5Y
Io63nqYlbNif8Vh6HOEIvbyvqubuADK6b0eLJ7NN93uH9e689PHe4OBDdPvnrYGE
WAWVG11WgbIia1FyUAioZi5bSWCSX68sLngltcJQucfR7mkfg9Qhwl6s39I3chxN
3AAx+6RBpSoNgJtMaNibhhZWdwDO5BN4NCzUg9jb5Vz+jqS6C2zv60Mz+R8aqJug
pU4iSpZyKosyZWytrdF0oY1vZ6W0ATyTRbQwS2ODdAyvHqyrtifCxGX6EMEWGRaB
sV1C1wTPWfEW3g/0/dWc6mKTc/G1NoAsQBE+wcDLcuqFOU2Pfi+7XAo2FjxHhdRA
EPzJ/TjMPs/wEV9A1jQ+kit3LbuMwHePPiDz7KX7a5CCD5tJ9pdOrTAygGpWRPm3
aAMlMjwBugQL3a7DNjwWSQDQmsidRmC5NdG/wCj73lhLiSzyetOYZNXYXY2rgEi9
Ah4oU153K/2BtqvOyQh/WPrt7HCsY/Td7X1deZxa5MBHYhT7rdECarjA2xN0erbf
Ir6XtqkksySdrIqNfHDg6If0v2gEpSUCUSbpMR53lVM2KifXe8rIJI6PedAMmwPq
r98Q5bylpiHQyg0prjz6+1mzVNLHrxL7Gf+xsp5jf4+r2EOnruVZAUuyjlEvq6eP
QByn8biGfGc+o2iSXdvIbcYKErTkJiAivm62mlQVGOudAyTu6lKQZXAdFkR4uNRi
4aDFU/JCSPkif78i/0l5NE6uTAjP+NPUigLzY6V93PuGnZlaJr7XIrsD7KyCc9Sk
pHV8i0j6KvzsGQpNQkxYbmEhyTNR/ERU4hyPMoQSGR4QGb0mlhjEVcmQ4KrNRaCL
1YseELlphReLhQt5QVr8CuWMIOCbPdm0JUwMc8Sz/5XOvK72tlKloxrt9u95JhS4
DnqLl4/quGmpLzDh+U4KaummCga3Gfl0F22xWh4U9twBLjKwREovN1WkxgqobE7G
16dklj08oRfLInWmV3ae/7Xgi4h1dr3t7lLZLgStgtZhL9ziFBvIJ4jH/yfVkBnA
MpknM1yBiHfbGffnRo1nb64YHVKPB80rk6xGxZjCdhU6k6r+MM0MSlKHJ0tm0uJI
DmCfnpawd18xvD1JljNZSllck1bHC3jXhYbtYAahT/rj5PehyEACXgtJNf52yusW
wLBqSVclvDpuk7ZD6No6tYb+lVkaggxslj+eZ/DtYkdaz7cnBcBBuNqRi+y+NmaO
gMmi7VgvYfnA8GsBYWhMAgpT0gs23Z627sdtkhjGkA2nb1q++zL06noWmobOE86G
XF/DO/iLp6rBCSUkkSB+kwcmBsMZd3VnMVlEWmN2eAGd0QoXynassBiXtRhGGS2K
PYPcgCW/B3Vv1qKpZoPBylTnbzv69kNuSX+D3eh11jS7wsqodabtLmkMW/oSpfgF
fZawJmxjG6sk1JKFlatCBZRKhzZ1srSzDn5HWMY1inaAa17JYqdOxTdv8OSAJ9Ex
v5M0NNSe6xRbl5453ID3MjpZAyZzb3YTrQKnzS2zNByWV8lSq5repBxLlyetX2U3
ubBjEkd1OVha7SSRIHoipKoYjGjIQ/imQosQZWpZfgTp6w1VrKA91G58Fc8KRrOL
5rT8hx1AVZEgqddxSU5OjywuSE43ghehW3Zzf59aydSWygO7VOAjzzn/TZw7aPcw
vbl+iqeb96GAz7dIltyoYip28YMLXle0smjJH7QZqsw1VGWx7lEXYepBF4VP9xPQ
A5Sr2/5XbQKoOkp81s4U1yq/onYu0O6HycaTxr9RK8YGnc9Go1k9SUC4eqolL/ih
f8H4GQWhhMCpZxauNibUZXOPw0Orl1AQPO8fi3q7HwqnqpqoZBS+0Rumi43F7b8T
0kO68WwcqiVO0C5hqA/A0mrdifoYoTCHJqPvKs6u7VVHJ6ufqJjlvmRdXcs6bXkW
y+uS0WZT6WcF+FQQyEL6o9ToWb0mqOhtR1yfqF3yz+vU7+N4NcycaiYTs7sykc6w
caJi9vi4UTy/NEnNN7LBAJaA4baHu6vqX12rfxKHYGRuRd7O7Sd1V4EFVQfDctsd
L9LPEOylqYhyhBTGjS9Vb+ihyCSPjMw651BN9w7iRAtkPhu7/XfE/ZTiehjbrEaG
gDLyqEJpehPE+GRIhKu0BT2OmC3DsyDC17nwZfh6vkmZRq4/8ayC5i5TXChGIz4P
aTUv5Vbb32ikIlMxyVJRz/k5i+w5cSWDxO5FfQ+GhhIUYtewsT5OzzrIqw9C/mO9
7fWBJv7ajyGNzI5oeefNlSf1+DVZVdtuPAGYVMI43GAMbFgOo5ZkocBcLqriLqIn
EHwaQ0tJwHwqXANKLZfwcHwUrOChz06o5nX9vDeK6eAKGvSoZd4jKMvAW1lDbdZh
jW0UGr/8pKoYOe0TzAzdTO7BbMvM66GDzljGoK9rMva5S9lVnLMcnaSQRJsHk3+Q
oKhSiV72GDWBXNj5pu0doVXX9MOlZr0W31T5N6dtk7MNZiwA0Uc9RZeCU+xGUcG6
H678zElaMWujL8JXAt0BCMYkJOGtO94Qwdn7UWbqPC8j+rEB09LL571O98tM7UQg
MshZvnSelRw7nNVSyH5VUzqfNZ5eXkn72ylynUK2KdRHP5S2V7EX21PmyKbvXKTN
MJScstHp3yIFAfi4W5q5/jSMQuQYztJ01//EnmC/dJLoqHDYxH9CsWJ8NzeMXJAM
6Vhvb58rdo5rtc9s5ZbWJwGR0YzLJSLIqMUGj3KNew27Yzc+mvdfmu0aoRkj6u8i
K4i8KrcQK/Dg9TonT1MQHMsAAXkRi13DlPJXAoHNTlHvVMulhD5Zr546spuUowZB
SAUUGwGGUNxuQs7euRQH64h3XOEIUdwRT/rUQ6zRYFiM+ZACZ+3E7/8ArmcNwV/n
Qs6h4He6F5WyHtvFq63YYIhf8mjDFPnAjUb9LOPNKea3s61sQEd7tc495v94ndvt
CBOBPMIFnpu8exbYDoGv2YmB3BJNmjgW80J5sx9lVVBINJfrcOC9Lz8AJMdxuHV8
ZXUlvwaTpF3Ayl5olLOXgQ72u1Q39BZOJo590zAgCZf9w3SsWUTRxM/s8dDYXwjF
QAsSJE6i1A/iGSmNn/pEG2ygZqnvRvsYTionnIcO7N0aM0ssIGVfBHymQej0Pkvh
y7wmrT5pXPuFjd2eXOAdooIK3vWjXipZm1LgeiJbim99ECAQfgLVf74OvhUYahcX
VJ1Ii3QlvTTc9rMB5xSFG2FEAQG0rHojMwuS6kSZL2ET+SxdxeVzNyovnecNSxxu
hAAI0q55w1jpMsGg0LnRiCgK/0xl7cTuoSOqHDUNlX2QYjoahmxymp7vA1O/8o4D
le1Kp+ffT0Qnf9YcOXDxqlI+vAiGGv0tVV5kCS6gPfKSfqAZfnupN5P7BkCGBu+d
Zmv3qnCoaBQW58Is1zuhwbIr6xmVDMkeR89LVpxfjX+VaMgAFFjqF02S33YbbxHD
Ys2v+i7O1HAOF69PZkZMm2gR6JXNsNYSoIybFGs021yFqMf2/+b6rasHEwZ6fmu7
wLyAbb0kmFYEE+sfhaW4ob2rUHREAwYakm4LpylyhlAL/aPXBmFJi42/A9Io9hal
a/n4et+6qmvryH4kd+4ivvasdL8rKL/CggtzZmECaPAgKicmpYP9/ORKYJ+9Zahe
r2hNctBnvpSczOVOmc6/QWeG/UBbVvSinapBkMF0hCGZrDflHpIVjkEN2l0nWxu7
APmq1oo/CSDnUYw8RGk+Z909d0Km3Xhas5dEYi0YTpliGR/QwJzzrN4E4Dr7l7aC
80+B4S/znKXHhkUuXCXPaZMSVPUUi7LHgYQFZs3cmu38hhb+Rokl8i79CDKQv8QD
w8cZqy7ApEk+A7iD0VmDw2AfDfgBb8e/RzaQNfeTktDCL5pWhxSu1iBiAoFbHBOv
8YLPmsmoWcQRvKsj1fD7XNbnpg5lg3bKKNDvAUY9GMg3aeXz4hlE/hAuvbaIgZlN
zBllsqDgwNNI/yvBNZopySERsfW+D/qGIdQTxT/+8PT7+3ItiVfWJyRomR1ZtnCW
I1MJaIaH1k0BkCmBIK6mv9PaK5o437jYvPKD/d5/dVeiOPPGFdyOlKQgWOBYzJDd
Yz09C2Q97wH07Z5nwwg6hhGx0RYVuLvGml94F78b9LIE53oDaaw6hqdRI0TQ60+B
J5419BWRGvlTt0S42/8yIsj/yZXPAUX7LPrsuJop3By+uPF4GiJVY7uWty1NN0bJ
uC9dRK/KGG9aIdXZXC6mPFuuMDfh8ykVPmRKKfc/1BriRFEIHUYXhCuxXbnEsSb8
ixcPqQVsf12Jcn1VzRGMmWuXyzrbHfXHzZWwTGec9u/vifL1+L1MsEJ1olrv1dUn
IHomldwendejso6iVxq/ZkIT+ffAIE2a8bpPbUn22NMZFwAv+ig1K5xFMeFcDJb3
Hq605pk/VtirpDFs6kRvh9yjaJ1SifEpAZENs5ySzfnd7T+2k+nbriePLMSvhxt3
kSWkZlj9sSS/gAQza3l115BZz/FosTTnIUCd9bepXoAUllrV3X0ASRgSNwycIbBb
JX1ERiP/BXPLc4CcXBRmYhcPpb9C7kzyMxCvdvQu2tC8oaPh1MPKyawpx0G2Llwz
W8sLqkUreLHsnhT7Pl0M2sdKRluT5vnfZKRpEcifuAYNiAiri34V19qK4CvQvojd
E8THsbA57wHjQNQH/XHt4rY9bvCjZYI/+BUAYpzfJMpvUWml5Ea9aOlYZxlq7HPd
16EEWac79Hy14ku1Rb0NPpBSExRGTReE8GaUP33e2Dfat1MbW+vFWpflr2YN+Sr5
yMRudgiUssKPDDqj02AZAkcA2u1gkIaP1hyZo1GonO555JwgW50JFrLhiAPkyYHi
VEJsYWKmKn42iCnWJcJEkvnCNE/90+ozqjGsGjc871NTScwXChaycAP5cNKSehxr
gytUthy23kBwaOCMTro0fNMxV7sphBTRhofUgEbhxmpPjNcAXMndq6+3RlbXPjT7
+Z2x15qeygupY5xbf/BAALwkTsObasObl/66UPuMaPF1AjE2jg7qmtcR+ZSleIlL
DoiLwrQ7AWuYyOPKc2zdEtGWzJswJmVOe+966c32iZNzZ2kn6xU1DKHRX5bPoRpE
a4PM2Zx2dTx5DGM8FuuRYKu+dA+Y6JU3hTRC4QpURPOvGQooH+2WQoIMhiUT9FXd
AxBW5PEcigyKZj1Q3ph4A7G+exc2/G9o4xUlTrTSmZE+jgrcDPC475F93kJ3KCYy
CfZMHgk5v+9LhfRzawlTkKqlsA7O2V1QRPySDBpn3JeJrvm6mofLNkw9AmzUaqdV
wzrfl2g0gsSDCLlIxyBtfOLji8YsT0tyUzaW0+qj7OArReRP2wZ2Z/tRWmCyJH6B
LPRxvYsWFfCQWqOzbT1spNKftC7IswzBf4uySNZNEYi43sAekT1PaH9X6o2xBF9A
lEgU+XUADTK+30KogdGMMHDVSSEAwPi8VWvrujoEcHVjTE4SE5ldHZhrU9uKWx/W
wwTnHKTxQUSzsFzZc/1SIgNQAdoJKVnBI16lCokYhg1AiFIyiuQ/Jw2sXxVvrxnX
L1xbIxBB8bPI2PSQT6y6ZX6qnx3Lbj9O6uwupCxV0nJnc64msNgLEU3Q1u8TZduE
CUOVxMyhGS9imyzUj9ywEnHepPodzmTt99rl0l0BsLJchxiPEUuBze+DNFu7X8MD
Laeb6T0a8ETDDgUCH7Cd4ioR1sU70bP6+Tw2L2jn+i/eI8Iti5OxIDLS1MHvHZYD
YATEAPo1owvN9z4oYSRqd0aXJi3lgV5BDoOsnaqj8Y72+h+Bjy3KwOsytqhlUK7F
50jF2vUZ/QS3SN65/eTbZKX2eF3eZggfGaxPPSSv+dQL/evmWRrlkJtRk+jYwIWm
saaQ3VWyV/vk/79k/s3USubqWzk/l05a3Hdk3bk9kPTyIhkuu/rU/dy4FxNP2G1i
nAZ3acjUu9h/yN2tzSX7QlI+djYPfcDMCCo3sgs6hsXEY5SORv4hUOAoLO9YBSYy
hIdvF2kyUISVxTwzT7WYJNIUOekzkcX/FocHWnbZVbqGFws+HYSeAL1x/I8qEl75
vcQE6G8PIcSRh+JMYljr3Pj18Kvx48pvh3F48RcLJz56VUvtl5bOD+e4w6wpxzsQ
snUAyHCBx52Nrg51EcF/KnSKW9cXJwjFXUOMjqSc/k/DubbxKct6TtwsUFAMMAyg
zB9BbHbeV0MnQ5chuGi63Sr3MIdSQjLVA1oPrtECSmurBdFQAiXIvs9n0HmF7gLo
oSnpfnIBt6c6LlyYypEFctK2md++nhhFpGN6j9ZDVeCkFIfxyA2Yy/d9PKZhYnkK
/ygobvmItUjthmzG04jwg46vEIPwSw7xFxxG3mOm4JmQW2I0Jah3WzczQgrg60jb
vo4B6YxAreF096QX9I366csXn2Fm9h1ws88lqmZ3hWvL7EpqUWzudBsxcu2QlAMw
boSzhbGxf9IO6hDW23m3gbSslc7XeA/m/vxII/KaMz1sXnpQF8Q+v7Sx6lbfn0EY
UEPAWzEj91AfNE0seti/Gyd3t2w0z+bZSuAAEJLewZtb+6RqFNwRO0WyyOwHFmq4
1P4Dp8w49NFCO9TRXOfyCuqhFQt1Ig7gxvpAq+niD/23SOn4l4BywS+xlfgBetTv
VmL55yVY3FPOs+tIeMGL2yC1BEkzOAQ9Xjvrk2Fwe3/sXfH6M1NleNKeKMVGJghD
/MQ7cSXmlUN3FFbJAWRRrM7yB5adTek3GsDe7znS+9ED459WkFqlulFpfJygr+rR
2KgMMkxOuGTCg5Y1CjhvtTWFCeXGrUxrx17yN+BRLcFyuEka9bN3Kg319KEButx5
GsoZ3dvZZzjoc58QH0hhJTTobjVNh0lVDxN0gDy1uzAcKY51ZXv+98/7BvnIoVbs
8Kaz/vAmjr0X/PUGBPHKRNvlEB4OXPBXGLgyaXmH3vuQtFHgz/xi/FLNhRtmIdux
GC5/YeIHAKoOx9lMdDo9JF/aCXfUmTE76FFdZd8+7F8OHxGCU+eV749hN0hSFEZA
FJbSPoVH6mHHimG/KSgjNYFc+jkFNPBfIOi6qfKqn50DwnhRhew4xWMaxKnnHblw
IgVac07ZtUWmyWMsRCpcUMQZ0W144MrB8OxK9I2GXo+KCUfsHcb7QhfDLKQ+Dw6J
+SYoCQ9VQraQS2PZL6rOmDs6feJpf2oHWIHNo1qd1B08daN0Ys6XsIvrBYjUfU+n
0SxDwBZmHgqRlo9xPzXLkK5hIr9WsccN7rMPrlaClJCe4yWN26IYx7jZwBZa2Zlj
VxBLCraqzJuyNAuDvdvcnJKcRxbcAyd6fvD3x5E6osDL6iw3ygglQna8YQ++YGZ9
srV2FrScEkInKeGBUdEYTNb9N0GDGwn/D1DpVBQVLGpsf9Q6M661CPj1cHzsU8A7
LrPXGv35fS+VRLzruEieYMfGRBuWMo5iqRpervpt2gH/yxlH/8RDdMSLUI1wSGDU
F/w5rQCgf9OFdfWRVic++hKRSv0JLFloUfQxpKebRnI+ed1TTikA5VrLI17l9EW9
DeUnC2dDsT6R6vVovAlrVYbxoiZqDU1W3mJTqE3Z6XWQUg1R+eNIsJfcdTM2HMpq
t0MQ4g5iaHZNbPjaI6kJNJgeiqNqfINXS5JHrPSo6z3FScxS3+jJE26vEsI3dLC5
AB7DOYel3jG9MuLnArenuJMZU7oWMYGW62Ud/F+rmaAGzt9VvmQ4Nm8npBpD8MFy
CzSL0l/ZYMxxEaU+76yX2KTyZOqa+kltqGZ0dKz+kV2bRdFtTW0t2e9GKcKYXs7w
S94dyJZWB7BsSvEYWEywFme2yO097T3sNtDMnhC1m2vUMNJr1qw3CWadpVkz5sLy
/eniLKbxV7TLSsJ9frgyi7WSiMCQQTjdPTiEdOF15sbwj+FZD1hjtBQpdORMLBhG
GTPdA8pCwuw4Ne5AotmiFAIKIZ2KgSAnw/V1kzgWh/WE0qPkyZggckYFshYDEZ01
cMyovDW0AiR8smZCm4dI/P/b6x5KtqNJBjHuPUyl3agPn00UX3XdtqxESdbf8DDi
yGZopul3/ZHvimMFbn9uKi8oxwUcY2G4BNZ2nj0tRIpTlRZtBh4BOKQx+Aci3Gx0
y7ZNeA7IZZ6SdclmPBkuv0YLXu8rS4BBNln1avJ0b+0Ve39OO1UWcZOwGSSQrs8m
fxBDakozXrWl/1+ODpth/ofk0HCb3w5E6ILoeYS+olMYjQ/0qZ9soc48PCvh/2xk
ExflM2hcBoiLsjJTrZyB8kcagG9G95SVrA1RKNJhHrELHwrNJByEbsTMfKT4WVTb
s4EEo0Cmbx46lWZjah9hfUvvPwpDLdErMHBcY87S0d7U8I7hMbVIyZIt9ujbDEXO
BwqUNVf/8/1DkkgJljFiZSiJK+xDU1qTyrxb4E0+YPNVv7aRtVJ2MxNZwZPRgThF
VcoVWOCLqJ5mcYIX6CwXh8fXbH+Lj8zFsFQSqz3AYOvY+mCqPTVu/Eb+SwgLIkdG
L4nfwYG0DY3ZzL3WM0Wyzg3ntcPblry85P+MypgntfUUh62DcSlqjD/g+E8VF1OA
06/9T2nnUk4scuFk9TBNktRg1qwO5rKlxJs373I2xjQx8zCcxPjJi22sHzx5wFUt
WlkT+Z/KhpGIFrwtA+R67tX8tMqMQ9N1xNMb/rqi5C2g+VIiDt8jpGDU/ceqT3LT
kdhh1/TFPwRiuAwfBXXt8I7BHsVzTKCPCnYKLISgnZtY3T8wzbwHauTOMXaFL3CB
/ehmixIeVhI2g3m5Kfo21FvfomDYCmrReD4gNP3dGNF8XRSaRFjJrLLT8iH7ZutR
NikizZf/C9+NwXkaDGfDtYNbSrth/uF6TGY3tIpa7i1V2reWihmdeQ1Z4RueonAK
KPUDMBEHEB6kb/5O+EKv9fUvPiQWNXnxoH38QUqMLGKY099sIfvqz8V8e3u10i4H
T2uSspmI2KWIWEIw3tJPYlyaV5WC8FXDr410o5pJorZ0/HfvLJC3IVItXuAOIWjn
oxFJptpLOunYprCXilPvqpKXxQH1z5yN9Gx10c4KUWZCyNHb9ExCeXUd/on8GGG6
Sk75hmA9UqEflKyZNxMvDlukpjkQjR5Vz1Dv5AZ+Pd4ixh0AQfClEQGEWxRWhAgW
udJg87LpAjdTuDMOp+wNf4Pn0JDtKxiWflCGwhOXHfeneI3oUufeS9If1s95feF/
4V2hWhdWCugtzE2aqGF2qyKOlPDRXFDhDpQZQP4Gr1W0/ufLKHGAhTLTHY+7/qYQ
vwRA0cNO30A49UVZ/Vj2K+/dLf+DD1JobQr4kvptOq7CoSV6cvIvRjyFfjIHzOyF
li+T7PiKeiTZ/wClnUoCwZLfZji7xzBtL+31F9pxog8WNoHyf0PhTVakeVkhMSG8
3XZFptr5qBj17vcoj/jK6GlrPVNXZzgTcvwYYje60XD1RVmnQ2AalF8Hy8IiN9ZM
pgmU4sm59abkvKksXm309VfK3tLA0qqdAQf42++/TCQ14hgbfr4cwCzNeq4PVeEf
OGpApjUQYhbYXxe3eXyaux1JLXjOEAwt407pa3LShDmqd6BWj198LY9cEG0H5vPW
2h8WN0nKjiSkA3dLzAGQCh77+wWvyyexkx/HeXt0ZBzPpgoe86o5RDJK9Hq9jtc1
87lwMJo+RNA6M3QmzcPw0Oa/HLJ/DipFUT7hBEDokqKXQaT05bR1tCCGhMS9B6ED
L/Yl7S82Tj/jFHe6wFTgceaBGSXN8+cCXhArwx4B1ApwCaIp3E1jNINEI5+Ti28L
Id1z6LSBxHHG+c4WV3fLQZp+OnLo1AHQ4f9jQIgo07g/vu+aTZDULcqs8Zz4eV+9
qwOt4fTuvjTMjPXobPysb8CQ4MAJeXJ9N/5EP83bFcF66Tw32vpdCz8KXdIAq8o3
ffxt7qQXJqVT98eJJIEE/TlaXsHe77ymSDu0wffoS/aUS1nBWebgpZgbGhE0Z25T
ez8nq0aHKjITh5Va/SVHN/Z4UvjBcAuozkm+d7mYae4mJit6GW6BK1K0LfdLV4mM
Zcbk2PT+AN3hSsfQn/jhModU9ftOYGUv8xsMAN1corNoDuLainqQ0hhtyNwrlGHn
pVsXPf6OfXUVnJ3h2Cyid3GXGIv7jiqoFsPbTarT+Org2+2ArriR38g5E3IkFc96
HAPcY+NkJ6VfCkw5QYKWuDXLUBCuUcXjplimsURtrKmPUDsoRcmZp3lzHlsJSzdD
da0a3J5y7xqftPTMfrbZOdwuMKCFF7sWihsQ2a8uSej02nOQG97niH4oUgNQov2N
FDAV3ITxBztDeBl2O8BAiR5WkJ6XORpbQmkk0VxXwdW31ai5Zl0UrjS/2Hw58TIl
H7ybnEATaWjvI+RvjdFLyCyngWy0abKMU6/D9hv3ZjFHPJbM/PFOo8tW/RgskY9O
6KzVIdsENL+9gg2Gka66g2/ccAZvI/GF7TNbhXy5mIkesnV+MKY1hJgrwOZycEhu
Dzrxi2ltnWMdRos5m+nhoj9ea1roIdyWPDxdSLim+9axdSKi9PvRe0EG/xlqja6a
4J8ZHBnPsgsw/SXLOQFS96zqaWlOgToemXa8Iq2ECRKP1gYwZ2ifkN3spxa7aAox
9D6+zkAiJ5D6aJEbJULoNDubp0FgPxY8FIbPPwkK6hJWZ0k1BdjlaEmye/aNW+oD
oofQkGjhOhtYhAPp0uJbMKSREsJak0CF5REuwbcR/XWYG0IJ79EY/Tk1X1yO8Ljm
snjscTO7BJt3s7h7XstgG85eUyQL+3/9i69a4OgAOmsZOjI7tQqYYXO0OIricUfX
Z3K9yrROlfNg6WLipEtiVfirY9HOyO5zJDBxiFlS6z3vm+7lEK/Tr7u9oYmdTttM
OLCjhb7C6lAJct8o4ToQTuElHcQUM6Y0sPJ73aHdZ6HN5SQJ8xyu6GP3LWhc5juj
Xum+IG9udb+vp7MPcflSUa9w5DZXxwSz+BEQQJKZRaC+qvEBVwdLfaw8DjK6ndLp
y0lSeQyjzwQm+YM0E5mY960OvUhjt/bo6/kuyPZD88/rVaqe8XKsgWx312lx6IyT
zpLRim7X2HdDXo/NpveoojWi3CS3DuDQalR2QCvdvGwBfg1XK42uJYBukI771YAL
6JC08a067rFnPWGrqa6UYcVQk7IgSYRexKy86pV8n3zrtXA70xQNpgmwYW4mmVKP
QyGk4npouIUDwcKpKHt5re+7mDdBWxjrH/+8aXY/45h96IYREi96oGLNp/jDR0UR
1m0oUNzSp+FEbOvO5bLLP1/NCATCvVZvH5lEnPPCtlk8zMKMGOZnXqWQduRoKO1N
IFakHLYHdLVOtTHL6yy/Wr5zcXWL/sWCbSgESE1OOJqRy/ZOgTj3lUjx4ZGmshGg
a+AnuKT6LOspTV9p6qm6E6EKbesJCwzBA2aGOQmLnbVdnEi0apok2yziy5dGM3Tc
FHhL41Bed4E31WO6qRDcWvkk3ZU7Bm2l1bqs1/xCSBeSLcSjcDdJdF6JiD9cGZtD
b2iLVS8bMNAYWsP9J4iHVVzXGUQadxSBrtAkv09R4rosgMzk0leG5TYQJpnHR/FC
/lojFmPXUc4QUrVUdPJZdSTbH8FbY8VhZqn2Aa25Q9kZrIxwC/Q/dKxCVFfhdXYg
5ygAeY7vFrqTs6ST7ucxkw1QPQStxk99E7tTcdib0JRq2kVtIA2I0QPA+kjOH0HH
DrKQavHpgrxsdNwewTTR7wNH5wDN8hrtLqUsSi/e3GBycw7ehXa2gS6J2Pxv+3PJ
FW92planA83oT2giA0y36nPbCB1L1kLEoQoihe6dvklrRFfGxcD24nnCSzwYkiWy
8dWlHuXT5/IIYAWYt6a92Keh/3o87pkEpOoysOW4CsqDKC7JRaCH1sV2/7cSIN27
T0L+E+6m+MWPzAp1KmHdgA0zgnFXOudHPuQUK2AVhKr1Wup5GYvft17zcRTB8y9d
tdxk12T4MXEg4KjU0IF84+CS3CelolYwDoCwqVsl1tUVAi6Pdeaqg9CfmUbtBYGT
3aom910LiH+DppJLw45y+iG7ft3lIWskvBczuowX5hSmsSYHfM169zN4B7bjQJwd
N4Nwg2DIWA02/xPK6xJzMMlRGvlxPEnAmCWN318L6lfaW841ngvsaODZJtryiQle
UJrs8NLgTdnHj7G+UUMjOvVQQ3jR0O5KhqDBf5btX8KwMeBgrqs9feKSUws59uXH
rPpuimp2pTeYsiDuKFMcIBKcr86C2H87XHEH1++ihc6B2rDFpWmwkClSQV/++fPe
asAoTRqedEUSdhpAN9W0NBxm2E7r3KB1TR3yZeKNQFGv56zosE3KEGmbL83A/z+V
sOJX3oRsw8tQFJuvY/OX/zfbXy5drLC8zF+12xbld53qm31MlLWkxymcSj/QTIOq
rSsrcvyWosNadAUr/pnaHrNILSQo8F4vwlK7LzRX+dbSzmi+WnVdkajxl/3Vi9G8
oIjMol30SrgI+YpWrQS/n/6WQ0IHfKMqh4Ha8e5LHiknTb6+59dTpAKfVwvm2nLm
CEDv2IDOp0agCz0eazTx4qDZgD30njNAOB1TP0l8wD0F6lcAhzmZuyD5JtxD6x4x
5+Y+JVEN/x5pbx6L8wwGNr0UWMYmYav+oENQLkOWn+xnE8HVyB8V9ZivWL+j+ono
9qxeYT9YGHUYSNCMuBsE4xUcb2QEPJsNsHFHkNYJys6Gd/8g/ibo9+Q++rJ6NpHr
Am0aWoUcNRRoqozncTtRlpRvn3H8SBn5R4vSQw+pKQLAF1QexeuJjuijINyOYU37
20zW3q/MX51qgH1aGskjLYimwhfSBIOT9y/RrK/+NHiTsfSTXTlfX1yFcKMtQ4kB
FniEhXte8a+XV67vf3Y2xiWiGz7ZWtJSVH++LliskIpRnCl8aC+RgwZD2GNcELbo
z508U2HDMkAi109dij00144kPNigjhaZMtNFmn5ggATBIq2udjRmMrKB7mDMidcL
fsWWiA/V5HfE0KbunnlBau7R8cboftbRK2W/9ZDlWHjORa9t8lR/OmsDTgwT8Ewc
OIwibxXAuU80ORFKn+kD3pG2UAUZmpiH0XCMIaQEGFspFWB3NM19RzVz/Hkqnykr
AEm561/NTVYtNKg7mLcm8ix45Suf8qyS1MNp3l0SoaN51gEURXl86Knpec+jxt0f
W0LPkLFTqc/iV6u/qdOrfVTdgzs6Ty/zxeZRhTxclnGTjzLKgF/mCX9CFzQBt4Fg
+1R+8q/lyyzXB+GRtvs8/Kym7d8pIh7bmbTXIA8gYSeJlX9yqUcP+evIbMr9EBgc
wN2NDjka7wE48na/GNZl0I9IQBS++cuYfMVu9REAAn/rCwOIjl6oImTR512qZeUY
87DB0lVPdJB8ttIyEMfgMztkmBfPKqjNi/kiesee3zyeyYb7c9r7qGQ1RjraV8dy
6/4j8mgvAN/w0YCNdHhFMwWqDqRvpiWVO0FrshthelM9bzIXXybtYLr/WpixBELI
ykBqnh1JPzW0/IHBoYXhkYp6jC/vcblEO9mUj10qyHkwy75NZJRspwXwggyVeQIp
XyfNmK6JXiR2oB6rtxZM8ZWI/Ppt1fv5Kf01KZGQ6eh/UXTGf6VFy6IP5oGohM9D
lswco8qjoq5bUdKjhCiA+COSzwqYJFpJCKKhjCA34cHoNcPrWd2CC8pdGNyCy/V4
czo/i+yuNTZysOSKonG1Tzq5wZtvrZPYCvASm/qB4rYNrTgPdbLvMeyMocaBtUOJ
U7FFK3l893hTjzxWL5VsqTlrnO+eoSfdQoruFKo7u523e3Eu9igAnKYaUx1Py+k2
lvEG3mkugxKVF3qMSCDu88lbXmkEDEIoqtNeDCyEumzOlQSLQeoOmcVIcxoUo1PX
KZ4Saje3NR8KEOcfDpMJKDkrDblg++lzIRYP4mLF1OQqiM362vS6J7mb1pakSBq+
GwJaX2hz4hX2fCspUhM5oCpMW2s++dDzSS2P1lyFRuiBZ0Y53SFRJsQVT+XCIRWl
9RCFr902nTb6IyaQN1UmGXun+1v/wDqlFpYJCs4OZ/7aXtU2ixsV2ixue85unOJi
sPyDD0NDNxnMo54N3CUAfC6Zr/RN+DCIaLgems7BD5y9JLQa2ZCiFbMkW2IsKung
gsDS/uS/CQV1e+t9uqWmkjaACLt5/JDruUh/VUY0ERuhdYcfiUvTOahYqfslL1It
xoiLZPNiLJEaEF0vdt0d1q38AaYw57yiRpPv0ptb/on2oBNWaXm6W9Mbnu9Wiip8
xziD+mlrYx3y/fC/TGNxznT8pwsq7Zwa9Xblm6W/fKgCVcRA+2DIqwhKrcRyy+bx
nSymKImx1kpvbsXtCLB4af4dIFC5wnzpkcNZpzlPW/aQWbH9NXjOJZvlo3t/jpgb
qPuGki0nMliNaGDG1//pJvfCxO97YbFK8TsnKO9hP9EWcSR8Tfo1lhA4xYJk+ubF
zfxKnWTFXEci2NjJVBu0FlXT0Pg2kzLOgv4SaQ/13vTPE8xuhDmS6sn308YzYpbQ
1U1RfKLdM4AIXq+4WAJv1k2X8Y0U/s665oOj1h8/6Mo7KasJCUB6pqfJ5K9dzUZl
Hj9HEtc7rPAEfN2n3CjHG8jd0Pa3/S1q/8tuVD7dbpNDcEnDd8nh4f6/nCOGeNOH
na6ctfehM3iZJzGCEGbvrS/N6syZD8U/e7nL6CTwBdNvHyFwtARgqySCHd7s6wyu
BlFauKS2GK5Ztpljj4tNkSdm1L7ScshdUt7RjyX3UM/wXX2t8MfH/bNqw2TT6Sr6
NRTr/+vHF9f8iwraOaTybgA9w3cNyGRAiVrMaTFexlsnxnrmKT0ZIXnbkKeBDy9h
aER3kHvXvSxxFfo+q+/PcH8KH8hL5z7JsYp+Z4OV2VFnvIKCfQtAAznwVR9eb13w
EGa3OO9g6iTVHApwDcPwo0Zgoa8tG4Q1qIYFHcVN2p29HrfxWltUPezjyvnImX0N
y4geid9MjhbFOc2bj1UubGbDfGDdjljIN5jonhKlx081PIa0uvPbRwnJwnr0XCGm
NwtIyD1+a8gbZS2UboZa28MjnVh/lSIPH+rvfOpWRnfLFnOHD716uNS+Avdey5RK
ZTBJvOJkb4Mei1ILS7vWsHX77FNAMD+Cq7mqGtu6GuhwPht3oCWxCAKd9yoZPjgs
tZManVITJwrga1aaV4FHov8MLUvA0Qto0Zp2knqa1LfqOPyuWvCAujiDEA9wvmlx
2GYw5bTaXUSaRxvVJuirv8AYjwkJ/GI0J/yIdPCrJ1Bp3o5+SPq+q/QYk/gTtPE7
eZpt743aExF7oHiErVJJfKBU4AsA+nD/tjMFpdf1Chjax8z/SoLTh2XQhIsmnYTQ
lFYUSDGIaDy2iRm4aYcBA2jVFy4ksFdchpmCh8+oOKWsqaL96rXEb8/W0SXH1Ggr
W/lEjRK6hzOtKIrcCSufmVhmnJDtjexocJsH61+KwPHkEA/d6aEJF1aNc9QITjlO
q6NtyWZwQcBYn8tPPrv1CJcOce2qz07eGSbB8a+lM6+XBrUCqqMGiRiYNnUzcoEh
qH3aR4nroiUyC2eNXrWoS2jmWy2OB3jXK7CSVuVB3HKOw7G9Ql3B7KgtxgYO6H8p
x5LxamUV1keuO90mPWFxuDRSNG2MjI0TqmB2+9TxJ0szdg6HB3lwSi7FJp8gDFkM
iVce1+qKTrjDFlLwwBBlGCzP2Z96Vv3NImLyIkvG58Mt3CjRpPcLmzVRyyTdH+Gi
9ChYefgN5Ko/ScbJ4zYu1gnUzfEpPKdBnAhDQcvuTByo2R66im9xypVzaMAsWpi3
fA9UfTRHKjxsyKpXZi/1wHL8mQbO6UiwpOUNNPjtxSIiecUhvnSH/frkv/pByKj0
/kZkVRhS6FSVAo2p4GdJms18pVwFK/W5d5jwdMAiel4gReXPMl1IE90Uhra1b0Oa
b62USjCCT4xRyfUdUHL8kZCmrxxzpMRPj17I2NpfGX6Vo53OqkfsFNNsRB0Xt5jo
gX/3y6N6zeHklZvpl0d1P1y7D2lekhRxOUw2kK1+oK4q4nMkRvcZcB4WIJB6t3kw
fsFFZ1MT5InmezHu/spDu0KPPh7baFX472x4IGrRuxYt2Twnbww6kHWkDwKVH4FU
ZJwcOJDxpbzHOuC/AvyqOKYLkEfBAEfmU478iKKG1RNuEu2VZwkEWnI1g31jcv2P
Uj1mr883kN5Aq3obOOwOXYDorLYZgnBmmGLIUBbfEMx6qglDazkZm5z1y266PXwD
/BBYArn7xe5eJ4olXQz3aTJTs8uPJK5jdtcT2XuzDNRpcJkiJbvCSCQ7Rx77yXEB
tbi+JzbQApV5edQtVY3kfRJKxd9IiSiIUJJinA9jyZ9xq9JIVZuanFLypn1ZYHwV
yCpcvuBgxsStM1Fyshy6AJfIoFeC2shZENXV7CNz8RXerMwTZRI1HsHcFThBkNX5
8/CbTGgeilOzUGtV/WAmxarc0J89oPrR/Adw1m2Ya43dq+MUWZkVOpNfsJ8cR0Q9
6PLSKO+dqsDebF+BviKdrMmpswJDxf+X8+mKvxFz0x2ootG6leHFdUo17B0dZFqx
UcrTRGyzRUsDzyprR6xFou3lnhT1L/qnF99EILjBVw2j5wZTdk21oT1pL7YrBk/l
M+fiM2AmbfHyOLBS2yNBDM5WAk0TDQ4GkiUO2hlI7fdX5MvqG/SgYHFOCggGdLzQ
b4RW9ALPqgXVYLM7Kxj83vDJxTVW49axMNi9PbkfTS/748m/NcBIPm0fFY6Vtqa0
ZLhiC9VqH/+iq5ThYCEliJIPlzcSKRmRExGCiqLm9RPK4KYUL8+5KmWg3jfOdfrW
aC7uwDseBatzIYTNDVyg58yNpmI776SGxRWsBdTMQa/DoSzWnI88T/0j8MryBWLi
U/rAio5JQs7SttV3NLY9GZKeCjczcA/ulZEg6bD2/zd5WlQOE5ZXdhuctk9bMexi
HTnIMzuIlboCtj4y60KKl4vEYNT2YrPSDvs2LQ44y5ql7BkZZCAuulgzLksejnSt
fCtbM/Ayora/tVEwoNQx83u45yhyB0ciNwZfnNAJDddc6UZThkcjQTe1xGaWlm2d
swhDg3mK0P4lFAYybKO6JqksbwMWmxRD0uFlejCMW9ccAouAEc+LKQyCmyZNSeVy
+YGDTgKlmvyCFoUwaGTsXng7Z/V2t6z4okdhmbXIvlZpg39smsLqhTjf/2dMwN2A
sHnf2Qds4HKLNcj6PRtvm4ttOw/ObTciKSPKjj4y32onaI7zT/mYlo4U1M6+47hl
yXbKnKvAcW0O44CGdMWTIv4/gE8VlWGTVS6kMwA5zfgDLZ0sjsvG02oUqIu4SF2m
iSaQAO4+S7yvoPyC5ONvJswndOh8zPcILBYauTSieKUHAWriJ0iPNlkcGALHqrx1
nMVuDTDYkV6NdLzBlbUSM0HJZWxTV1F+lyl9i0rvm5beRFfkQnbYqwjNmk6miOmu
/MOkU6mLUZhIo0ojJ0RjqcD62XWI8meS2SgxPhLa5zM4dOOcazjwjCc2Xr+AJwPS
DukIK+SOOzX7cw+Q/9hHb+9ld+2xlhkx9y7X7BRTSpmk66A1V/VoiJuxmwPDaSgt
tw7+tTmCriBexQUxgI6q8ySPqF2usXj2W2m5inI8Vyx8GygMF5HDmX6FlRYTpnbU
Lv//xwPTy36UAHlxTm1bxpVdIIsXOOYyatPLz28YsgriGgppTLNM+YLLViO6+E/k
89rEGjwKFUZe0flrHG3JWUgGyRcJRa4gFTU+3QUvdih5W9Wk84qNUVm0/GiewyuK
HC0QKAL6gmw4ZxxdDN/6L5iNYyW3f2RUWlPekY7B15Q0/ibaLfZ5kIF1+wvC1iqF
7pEO7uEDo2wEbwm4zWTchgAVcE2Z5zY37QZwh99miuUN1G0O9gui3h3H5Fr0fTM7
o1+LQ/9hy+Uvtraq+4qRi7l+i+/SCr6oRiQhbuEMMkZJ+EWBAEF9CA/NB7BxGZ75
0JG15LexkmqcVP1zyan1GxePKBf89Eagm9idCjQRGVHkkXaVCxrD/OZeHI+fJH1/
xhgsYliRSIM9yH2n+485f9LiejLVh4sp6ZCAbm2ObdjEhT5XbhV8ZK0YoFhyzcne
+66gkltps+lh8yCG4Q4foYqQZ5M55CMD6e3qPXxpKwqhWILFAwOCSWWCkxyAwAPH
TqKOkHfJDzk/A5c458TvFGij2L/HjHVULdCsWrpYFCm/20p1/OVrsS3J0NSeoKAd
ZDYnZ5KdBP8kXH7wf2VnJf7rFdfu5tEHsUq249WqyJ5LIeAYXRZ2e0gJFi4w5RXS
YrHooiwscylacz6GWsq7IKEvBPNHB21NN2KuUeR6PqXMfsGzAuiEyqIDdjlpG8bM
4hvY2T3q5qJF7iMO0qZO2Qm2pT1cFkaHaM5Fj17ccHy3/uy3FSFTI4mLZv+dq8Dk
o965wFa6Pw06F2yUAdGT03GL1ikHfSmLtkfIGNC2spr85/LkCZlBABtAe6Vldc9V
bKuQS3CCyEFY1hjk8CRN8ZfgkpkTKLyB9XyVGegn5YfRlqhoRYSuQyvjOGrTDuWF
ajypX6bEKzLq8mMjgqhcYUvf6IMrwCy4pye+NYs4+CYGLeUDpVEypLM/YVbVLbXW
E4H4OvUaYtFM/c6VSsLWGQGw4TH0p6bBLPQxgGRTDfDbmPqdPm5FXyM4FvM8nd0L
IMCfVRPT5jZiBmjSwbDGAoyZfb8BVxI+FxEOVr9jRzUEluezf6N6YRTp4Q9ZgV8A
Je8Fg5vCwiH9COGgQqiiqwGZ0qarH8220UTcjFp3lvVOc5idr7Hm+DiRxxs8WSSq
DzNEgMGtV8ubJA+U7Wf0KuNon4IcMx0ykC2iQnIso0WeVjZD3qGNZk4nBcxTMUDX
DEb2NL/VEEVKF6Df3tj9FQ0WISUo2kYq/A3yKKxQvI8mqXLpOrDEz5kwfZc4f6uX
0HZ3RLDjV1BlL1VN+BZINa+0LbWi/U6rRb+tzfzm5XOBf5MMOMWRk6Kmh1U6QuSg
HjTqWYVwPWiJgH9bSeTZKDI5rpu9/uF7QS93tJl4oytMnVWKeQ6s3a5KTfEICusx
z0LStmwf7N0mEsGu2OVOZSs3wEmO06NDjgRhwyxb2Fvx1tTshC/7tqg437KlScsl
Kob3OTxBVMkAe/5117VKGr6CDBvQz6t/boZvnnv+fmoJNLiDf6Jd4bTg4ZS/p5wt
23/Pj8U+xQAb1xFUt0xZov8MtsljQ5UzrWCcgad5gLkhx4l2h7t3k0btbveU9QeH
O7/0D5hGYrW0atJuWTF/VvXFt6pcpBsHBcBu2u911ff0V0ugMHcY/6kHQOom90Y1
Gznin1RyzWo+xsP8PBwVcumR9odDhARauoPrrC9eDrqzpX59FPW5faObiBxwfnyu
lZevgWWqIlWXxVaG+CwScBkQv2lME1ffy4avwRkKn9gaOKmXU8xjNMlfWHciLxUN
kaaNt2iQzW1SR6w+ST5Q4wazCjCAfj/VYfTf+L2OD8X5KwF0HF3xaHl40BQ5OTHV
HYXhLZNRR73Hd/ijVS9qtCLMBP+L7hTwgkI2SZx0nzpHT7Pfuarq3Tb4h37tU4tm
fbhqTlK7hLZA27UN6/jR/rSIeYLPaXC05tUjWu6SpI6Kzv1JR7PlNgwqjOzpR6zD
b3CAuX8Esn7ZCbvE05p3eSM88WAz8hae0/Eu3mEaYEr4LXWL/g7ORdxGogAyNT2B
cblhiXUO0nFV8qLR5ZCogKVzc5IIqRGtyE6LSMVYsSCrvra2WSGeavg4ioGuT/Ga
zOomirXqnJubWDcwfm2oLHlKb4V2Dp7VtsWcKHPwt7qDf362XjGs/BzR/gvK6qPG
UGSnj1v3kKuYlqTPgNbMHLEAgVMTJ09NuRIWCNlogYpIkOg0h1lrUXlooeaDJGPW
mt4ZgfU3W3EPLXMbbCVjneBOIzMDXEnDu2ywVDpf0Bif1P58Hs/TwFheKXNsiaH4
7zriHHhx6D1mpWxViDBiwCBhMm1f2zpiJ+PCd1NFcEc3kJdSAgOLVjoMx+Wbzr72
OLAv2BhRDrmFER5HwSa/kUsE9jpqdtTA6sTnRynNeZdmA0/CQ/lX6gqxDsoWrF+Y
FLHQ1j/b0cxkmuiFCMDfa5HbDPgpoliMsKPuc/HWeprNFX/s8RKjjzNMfdLZxAuM
wIpPiIXfq2SH5H8GKBs+Ug6G/skcbDpKF48OpODHEVT5aCvNwZv5rJgBPwLm4LQ0
uClnT2GlTP2MdY4B2vS1eLruqvszkp251n4lY2/vvZ0c6tdWgWynbE1wZYceHuvn
TPGxXJFgqD2pJ/FYTzrQsJuJHwiNWQa5VNABQr58tQfNU8uROF5N8Ymg6dlbngVN
9/+ziZeSomx0C4aA5eNVZ+Qa2sLs/kFxRWbjBZFBQr/OBpsrrN6WQJaKHpej7nZf
RqRUYtowv5IsX1xdIk74xZJi9x7255U+ClRWE9jduXjiTBo9K3o8wbD+b2sC4OPS
ISJCQhi3yj8Vx/w9yEIDVctWHcdrAQI/7F5i4y4uI9qzossVZYsSfF3KfTLfFVCm
lE4itbAf/nkVj8fJXjIh6qOAzDOFbhdVHzpNYOsaBE7T2C+podMJQHGRwShtzT59
5cXZeiGf+PjaejrGeOJjc36DBel9VMOUcb21l5a1y+yBBfw7VV1VwjxNXjqstDZC
lRFOm5dQYXdCcdRsjQDnSonDsClk07YvdiD/wUbsSQevHAUsQtBFccB8XaADu85w
S2FPh8P1N9RHPenWL67JcnOYbAgXXAuNDwYnCB2pW52qSi7geZ3PCOnzITnmtlLc
osJe57L5a5blz0tXfABM4IqRd/ZoySxZvosNPjy/I8QzCqBaF0VTqbOc34YBB/59
E2/S8Gsfn6ktFgALoiqH6eExxcS55j+DpbcTFy2+0icD1MOgySWr0nGxJ9Ml1vp9
AfpnDXTslf4ufxKwNmceP+uLuKYyJl/cGF8gIEAR5TjRWljYj2IszaFePljPMV2M
+17kWswBIs0rEu+oqrbQfnjm146SoRG2+zJZ6AgmlkHs6GppE6d2d28vUKgarKj/
60B63sys1GwSAMhDQtZY5ueEYbMbT1dWeO+x4CKlCOH+b1kYXt8jbT8+Numh7jsz
8bYjJCUYNrYoN9zA4h5Fj6OvrZV01d/pmfMllFelt+xKxhRCEO7SZTQWqxHYqTzC
59p9nj6rc8v6hNlSxoYfRdGpMspGjIwjBTFZvr07XkaaauQ860+FjTt1aXVorLZq
TO2xX7b0F1FImF5woktYnWvFr6Ch74GseE70pUmq7TGZkgeUT0oXARO/S1TsxmOu
hQnezQPHeilKBtKj43HC2cua3oaB9cr5p6CxXtekP2CvOUiwhUrN7gXUPnmr7zhQ
e8N6xfDBGwociitWuyuTPwGHss80dXF5fJ3NDoOLs62A7XZmT/fJz6bVaxByZeNu
xi0PdMf+mshK40Or5ROTRTQRocQ2ANNJdndX8/iAB/fW5nPWvXFM+ytGpysCoP61
3mQP5BraHXrG2HNbHnzaeh+EKliHPNG38gAsHg/Th1EbMIKiwFbpXrVZcgT/sX3L
6mUUI7HaDJ6H5zDdDFxRXO/0OY/RJfVBH82r2Tyns6dv5FrAmSfIMKLU23oKGSjR
/o5imbN/96HxJvRmWn2S6XCuAM0xNAp0kaUaoM8Xl5dyk7Bjrd/k8Lfa0OXgWLTf
BhvAiaOIrRSddUL7YclBsfgVvcoQ54v5U3+HSx32ZITLsMMBu0bdbIN2FGTFaepy
jfSnt5/WEgh6Wxq7idBaL3dprTdwGvg5tU3tvtkLByE4Z2yeg+x/2yNKO52ql7wk
beiIkYx0wjFbsdz9cjhgi94H+Zf3zmuRf349m90Hk97raOaTZCY2wWo9rzCtYI9d
LtqVYzv4V6x13n/ywTNdleVBpGH3EvVEKIjRA0CBX98FD17LCQ+YwzMP/Fgv9dzS
eXHyXl6igtqiNN6tL8l/Y72JZ2KAFz2ZkPLeFq+MRxdoY8yiSx6nhLQrZMSKLWrP
tWogGr0151JV52yesDiMdXSb71ogQOKoiHpxaJAbFRiLQbxRvQFajRKke1Z03Yth
xShsvrwy14AcB+FhQ2FF2zN6Nr+Z3cLHCD2e2nfNUJZzRFjOoK0ayUB0f2fm8hsf
m67pPtaJOpjpBA0LQ8H6P3clZhpOTbtbIgF4iJInXoS//8+HVL2DUDGifFwp6X0y
bqcoaIyhzzsXGr6L8Mhc/3UOQoLVY+ZWXkc1dtPB/dCSxDseM/nGrd58K3EIwf/H
CCBhJupRA6vHy5wJBmR9RxqZDAUw50tlnyynAt3HXKzlU+FIM+JA4cw0yurxfBSz
nUgMeVQG6L2svaPY/e2TjDLh7s/UzN8pBZJgs3yeWoYRpM+CvSDbHb+s07+z2OxQ
ys2VC0tKt0bul+mOcdfNWmVw3R9JII8OtAxS+vPjNQd9BkqpkeVzbdi5bJenR/sW
Tk4fyrP85aI/ELG/psv2Q2/yuTWP2gajjjiM+ZFByF6QyKNWAOVQsfQuFVSxNhTR
TNRxjjXrjn+heWAKoUhI+eIXRoqnhdKG6vtzHNB385wEX6f3dUau+dpx77HNKXiB
V42VXCuVrvV3n32yl3IsaWVvHCyjch42yXiupvImSMo1RC5zt3kC42l1/kLvP9Kn
mRhsUMW79qdWgq3zh6pRteIc7ae3jw87KTinmdb6MBlaCPIyKT+tHszeJB2bzk2y
coBa/9UBIR+3UEnQOZbQckt8+uwttWKFI59iNZ7NTYehoRVu1FHEV0ZDxmNxJArT
8Xyh+ZsLLkkEhIkIrUhwHTD/wpQyy5DAkhODXp/8191EOmC8IsKCwbmAT6r4wvBz
djNCZFjn21nBtTuJ2iu3X2Wgq5mIT7AGMybxVc82DNWdBLaqbTsbyunlU0F/VL/0
tdGePgyvtobTJly6XWemRuCJHCEmBPbczv56Yd6ChufQV7ZazO7f8aY5/aK9ntSC
cy38sUsO2+y2XkddY6QwNj7kffRcH4Rfz/tnAQGKPYr4SoY4iCZv0gmFHFd64VfM
RN1nZupJ6mW3Iv+x2f7hJ08FxACahB6HcLUVjyajpJUVvlU0W8heQsFHDgtGkzU0
bFfC1OWHe+CONSykYZNIGYLiXGRLcZCZn1QH7uMvGLawg7g1Zzq+dZSBCIWKsBZ1
VEId+mErZLR9Fe5AsFymcWhblXHwOnxrdFxmDMgZ+7ofvfhCmF2mW9a9WLq08k5J
g+sA1gHDSm0XylA+V7beDKO6KiymATrFbUZ4EHHisDZ/osvpoZdHzUNHdsBvhYOv
sA8LnPfLaJUgoVg0dC/FRwNffal7fQ70JeFQ8hc8aFcKAOFzzyTYanvWoaqD4zZ/
yhYd3NN8zXctwwGDK+xHnVTQuWPm+UFn6mO956mQVA0DtEGd0Kpue8BScmnF8Z66
xPsG5J28aZ9Zs/X+3799XUvI4+nuyjwXLo/w9SimOneO+9qML1zrmbSyrsljMJ/4
IDOPqBQqhAJ9y4w6tu+PHVz6M0B0uJG/ap4ltFi524KXuidr0BfWwiIAUhyHUqG5
xYQvmkZvKuuZq7PyKoBueWhkgaZVu73PyXxzlVuQnxU9xcaguS2tlzSs+/AbXiyx
ClSc6curPtG4UToNMa5RTJW0Eizho0HUzjqXje1S3Ytuzoy0pXl6I/Bsz6RiPvo6
PLb6bf6qbWDzG7WVwQ5u4qezPf0QvqnphNlvioKOBrds7W1zVvC9WlaZne001XCv
kpzZxYPGbdghDa0fthiYg04y1KNvjb6soBGw/l7OAgpJbZCmYuwKPvCIGktlVVm+
qvxtvwuaC28Bv0QTm38XeVvUE3QF2nQsmVVkjHXPxl/41tl4LJIVC/SaQolAzMLa
kwWHBmEahsIWvtD7yi+bElFIHYSZqRJXkmBcQojLlCSxxVN+J88CzqF1uZF9HOr3
FUzqIyFzuiBJw+HzGlZB6qpX1pB1oVqIISlTWM0D01Ov4E57Tp/g6F6ypi9icAIh
i8yEN1m+bM6I9ngthJn3GzDouWodaIBFEt4BpHS/AIaYXCzO2X3FNEqNwIZSFhHJ
LGdjdtp1byV7yhMRZDOQz7XyV0SP4RCMlKWYAB4zDp5yjLwYuz40pmcAYA6f0+LA
sPNtQhl3lLSx7/mNGdWNflJJ5rza5CQrbeFssuhQcXoD9QDgTVd2mK1g8C6MigsY
6Xj5ZPCepWW9GPN7zJ16yc0VBVpaCYViaCbF0QXoMLitj00oKzAQbSAY00frUCCZ
iAUNnxF/HDTN6bZwjyKUJG43CUcND6y6IjBu68vk3WHRK8/mv7wELUr8NfaT0U6x
ag6aX91qtPPtGwZXn4Rf2cwWWAEbyu0r/IP03xAB+OLlYUrsWXSut/iMU1mU+HCF
wNvxyAb4QbLlcmoqS20YIbenHY0X5N5jKUr6wQpves30m60vtcqsIEIc7K7WZeNP
Vaf7UtNYovtYs12Jg+4lTER5JAQ5NdrolpQ7GDGunK3lc0ZDcemOrypWE62s9gbe
Eeln/Oqb1gPUFAXHC2u5LD9fb7MW1YvMQqrQYdxMpq1KCokdFi6lF8fJNdAozoBT
YsuWImBC060xxj1GbU5pGSrbNFn1QI+GQg5Qp+atx733zpSIcItb+M/VAbYpe3Ns
/XgvIQIHur7JUxndnFT3aWOfLFWPohIzdeG62SVIoFbTK75VOcdxQRayErXD/rIg
EHU/KEatdrwMQpvUCZWfhe3U+ucG+n3NliojgsjQ2aiLsvYMqYGNmH/OvM/Hhenr
o/lZE6AT1T2lb1UK+qmwoNsEmyy5K7zSgxTMzPwTbFsZRCDuO4gNGxdu6NbHm/BV
+ULlF3xALXfFo8jyuwEO5jt7IshRcIibCnFVdQTG0YpA3p2c4EUBRlGiPVrQcodx
ge3MzswZsdUMR0ykXiCpXEwhAxp3M4qaA/V419MPWj37tcwHHjlmQ/4Pl+/DKJxK
9pu7ktsfZojH1OCijunL+VLajtw7IAsawpKCc/iXhTXeQKB5m+ZZgc5FrFmr3yCh
idiKpm+eHhGzNLiEa24ynqBWtFWEC7SwKSmucycSv0DavO4SYQui7TcM/xfFuz6W
+opzbUN5L9ZCTDEuYr2iBxImParpf/PMV5v/XhXoGWY6fN5LyVfqK5ydDTr/Tmjm
CprcZXamQ0IWYarKPL+GTNXLGH1X+Awhwfxiv60afgDCYbYKKnFApU9e7wHjQTGA
g8NJ5yS1Bprz7HIBzaBp4NyaSwRRzgiKxS0fEIcA3tAY9jeIIL5POtEtd9sbQDYk
9y10Bj8aP78OuXQYTY+Rl/72GmPHPNY3iEHsjOQ9arOr/9Njp0WokTRg6/z2eucT
UueOVISTx1p/l/UCgQPK784hDAYW6+N2AJUx939Dj2CLSeoLTLIokP33hxy8B3mG
Zza7+/pyZEzZIA3n5Run7JHPp3JXrdqpax2pzjYHkGnzL0sZvxZCI/znpdpUFR8F
Pt8cASqMpXd+Iq74YqbzX/xwFul8DUN/n1THK9wZrXgLkQrLg4pX+8Mz0BZkMt3h
pUZdsmWnmsuIC0EBN3/xTippR89cSzludkvaipDp8qL/XaftmHoaWgj0NAVUI3yB
wzWwAIqCSDyQXY9w3vFpgpRLjYRCSlwmuO9zB0hSITxjapPphQaXCydaPGO6xmNd
i3Cb2xk+EhmGVm+diBwoOTo0/vEv7KQdfsabK6fz52vf3OcyCDyEmiZEqIwfO+Fz
nnX5srMfU9eMeh/qsUxCmdwdv77iZ5nvPVPBCWZSUaqt6cLn146WsZ564d2a8CGN
Rnyw+7/BLcMy7cVuTTSk5CXE+RyZCccN/A4xhkOHxU90+Sxx40RkNqIp8DdyfyKO
KS4V7qr63hRy4LlS6RIRsDYRJ+fMt3AF0nKR2Hb3exkMUqYLkLST3H6VQP87C0mJ
taNoN/dkIvpD8ufPFyE6RQbel4LzsWR2F6fNr/lUme8tEZ/AUuuOxaEhJeDYzUDX
+KY1b9gb4up2XnVmdJ5gVMlcCDsKurVlJGJa2a47QZB3/pgo567uTYrBSOQdJTG/
XD2OYY/3mTrAtb4HWQt2VhzLVvaXN4o0ZNdT/mXqVxqBlLHoJfqUlatd+9PahZur
v44AVr+SWBJTGEykCsWeEjgbgWlKFZ9MItLv2is1aKch/dOT4hUFjdtrmOgW3U8m
puy4prE460RYHvsgX5KfpESTrEA2/qVzKQSXpgV70otxQYY4hugk3qvUgq5snIqO
uY7fBeKXDcFbWuLecF1lUAMYmt0JyylDHr6l3eNaleCKSe0vDLJEURZLN2u9mYJ7
/dpH5d4mcf0AF9g1s6GZIARYAlIbIvfFIFWAcnnqpCV0y4ZfG72e8vqZGOkQTvnb
yXInnNtd8MeQOH94mRJ5ylHtzLVdJKO+BSL6pUTbAs4VOhi6cOTE7o0AjVglVSRg
hDIWArfY2sgFSu7skZ4xG5wSUbsY9QivTQfGzREwKtBvm6LGha/JKaUYnRsqw4ja
B84Zfc2ClnMLYZk21adsFVyKmmHjdf5W0VQtKdPZb3pUe+ij/rFS02ECn3Z8n6qe
pmWlXhYq3ROKeqKJt4xNeuUoVvG/FsYrJhh1sTIU151S94+1tiRUuHO4PWuq0k42
4ealPB7mywnmE34uMeWHLzwfFVxzCvDs1yoUXiTy/Hb+sQbdxRDgBZid9nlP5DGM
fn4sfz2vda2RRy7kI7Bi2FXDaMufEpN0WuzQTM9HejQRpXCVMpcWwQcAyIYAExV/
CmZS/LTGgoqv3k27REtAflX99zG3G6Y9kH3B1o5gKLsCbVkjJGsO5QfQHi+mqVKp
BCJmheqwq/qOl2Lja0f4V860QEdWA6d6lvpGyYnuFlWgP3t4rR7j5ptOmY2KPr56
ThFdaUjP/bAmEDEkevivXEnfWJR1mCNrsl1mIF31VOmVJVeO7DrLUamRzCOAu5wZ
eDwpMzigiSS1kyY48q/Mi+5EAV6ngHKqkp6roH0/gsFt8occ2DZYW/wNT1MiAoi0
/FrMfOGUv2bNbW7K0KfLcCCiMPk+T+4/VkG1qKKLiSTo5NKRYClkdfZK5CAz8rZV
USnaBN1ltByTdH+Hgk7YC68JIj8aemA38tBxCJ+Qerq0tZC1WOJKO0fFzAJ4niyN
8hnaVo94akTn7edC49Qr4vR6IDhZU0beoWTtuCXkXjC8SKw803bGeLdFYYcmq78E
ShaBr1yPvPUjMYhZARTRd4dJ2Iinx6ExNo7OD5HXz385QwK4W5ZZC7bVwiiXDxRO
YBZGYZevwT2yMMo83QSxTmeIDI5PA//vcwCpy6XDVuA3rq+2SQNSX2am73gQvich
HEyfEYw5LQFvauSG4m8sIWmVENHBwqYI0cMGxe6W+dMhY1waTJULf8YfGgz4dRqX
blXsGZymfhvbUbwGHJY02GTwm/lJL0r5ie1+AS2E9nUW3BlfZ7XOhgxRM5so3d0a
C5PSf2Ygo7pvZNhU3p2DTrgBpP/9lyOsA6op8Qm3F2KKAPg5bl8kLGtY93fem+x+
fL8RS0f/q3KKR9BuNF5BA9iJNSvljyYrVRvLdPFSQ1Ks4Wr6zyZx1JqGCEtmbhDZ
GPHSU9ij8jGv8LD7ZQKkJtaHXt+LmhBywhacbVc677IPLxxnh/uhir7/m7c5S4EQ
68BK9NDouy5q8SJ1kDxOZcoyadHkxTem0ERa4HehaCF19DCyqnSMThQiQZk/ffCi
XB8jzQfVs++0BeRhNLAeaPQbKveDNSUyqY/DZK2Aua0O7uU5awOTC1H4S/hId2mC
C5xOftTfeKD4m4kFP4VG7e/fyVad6sD16R99MvnwGjH5PAv9eMJbnWbCorytrm5N
Ct1rauxNt70uAz9sGV4lh3N2N0TzcRPSBRtjMoSe8T21bb7+f8gwkaxcldW/DXJn
mgs6lUFuR0ng0AMLdpMn5St4BfQHIq1zAapBKTaASLm13mZQkQkRQQ/DLkt3VO0u
q92aPctjh33vQfZnwyz3n+/mD5LTATYk9flovjMyulu1445RjfVzayPfYw2cLZms
7ZI5E1wx2LypP+EZSQRdRf0RLWY03MdL2V1cpzrcE3JGjqR3BfKHHp7GvL6O+RVL
ZPW1T+AYj4D/0j/Z87+LiQLLHqBLFPHtSXGEl7bxlz6uNwWkDFbcu4xs1+MZqXz/
vKsHtfBWo34GT9eqvjm9TaIaIizGxRZglZMV/NQ+eQ2cGMIjFwqIkmmjecRKeZiy
AfVjp/MLLwM2SwdvMUSj2IN+Eg4cNPY3lvhGlKIoOEOoQUNQG68CeFrJCmxyU7EY
grr5VFga+NN4gVvO3q529oPpryRjKSX9zYcIjnOd4Glx65M1u/D0LHnwsLRsKKxt
xyVpsJ5TI04nMtElin14D9RUumw//gwG5UngNs6nGMbY/xkiehpEx5ZzuNFmiC4a
2h962qxjH4mwwYOQO4g81fCPgXIWMi6+KKUl31hbv8xIjkouo5lPGPm7YtrOmzZR
s58191JoawOECUGH3AAEIoAwql/L/VaTzNeDNb0lO7dkrIsw640OEhKp3Dl7B8E4
xRq9PEa8Lj/VoYhVh0L5IlduiH7WLNEaSZqMydPUc1wUpfIGI6txCvWBfwIt9z/L
eq9rvP+hEVUh87Snsu69JXm4bYwSiF+IM9gPyW59CR10C+BLuRP2Q3+cRiEeKfU7
o0OQyvp+I8Xoq6+dhTobmcM7hYjSevyMcRRopZArZaqFSNYPAn4rhb+VudCo0/VL
RmGbiTPwuoh5XrI84UikaWk806XqX23I3SQfmtnAdvC/sSp4bTAdhU+BqnupBvXd
KFwjH/v6W2KqSbHB5Bl+q5yPMWq80Xir7L4bnSJG2ZgBT4tyJOeBZslgIMCdMHHp
fxRkiuODwQM3GNi02oWWn3Wun6LT+CcAVyTP9tS/BABvXGGJ7iLkLoohiS9i0fDB
8R0z5zK01tmu3eg6k36MtaevMtopnGjSj+5yxlMmufxvks4VyO4e1jdjBWdeIAce
8AxQ08XC11h9Khqwh85oDRhV8YG0lbGCG4jyOu0+Zjh3NgMI58WkJYQacrY3c/LV
q9Gh2B995EqXqxf+e6PWQ1/tHxOqrnXU7hbmm5G5SgL71uo3NEdyJINdPExXO5na
fuxNJSH/3uG1NpWBsXO3VhqisZ3pCSgbbNOzOrZJbF//hbybdlQmDPuTIutf0Qzz
sGCB64zNwOYSRKAhVb6Yoc9rWMTmpzasEH3pto3kwIlwkucnIVRS2fUjyigSOrxf
3jsoc9vIuzzMCPKsEgf5hGv+fueUbo1XR/Gz4KBc7MrFZgz61xAvFmuXPlJMdyPl
KpM3BdVUdzX8s3Ub1SbV6ufkkCPGxV0QLQISVf+l60671RzyRjV6aNDDIqo05zLf
V6lLsfm0PQqCEqWwq8/APJGs062dcRD24jaAw59uBhwjndTVUoLofjzVHfpna2Xp
/KVceOA5D8Ku3axZVGtEoSUW012mlq84ONqot+9pemiNUM8c5Re2z4HkqzvHg11t
5fqGvSEEI/m5Ya+fiy4L/ZqdfVa5jmiFRczfV6sj/1p1Y1YZ7y/tHBtcRqgMaFBU
Nm9sgXD58cD46nNWdhMOpKC1oNkyyS+0Zu6MlyMOtMiydgj4oCGjUeNeop2uIMPF
Jc2uKwHUFGsTdZNv2a5PeuozFLZHzjikZ9aycS7jLe3vAMT7Xc1Br8JmeYDE99pl
0cYcgjlksN94Ib9lOU5uYsOJ1Yix8TbM75scH+DJf10Y98z42KiX3srEPM2Hnbg1
v+VbO8c9MgyangPjYy3a7CbDhJEuBC5vyh+2Y2wfPNESpHA5V+kTnGzg2T30xNud
kbqpwJ+jM6gqdOFJmrCXw1/E3zOOgRQLZGLkpNnUQ8VXu2wWgzXyKfQ3+tqhXo5S
VCooXhGH/P+Hqfq5fYOI/Qi25TB1k3aTwXtOEk3/J0YvW6eI/nqmiuh3ZW7nsWgK
E6f3k46ZEPPdiuFSDKTD9HQ8cDManjZaiiZzjxq3RQtnFVlRBOCSgdxJhr+QZ/Uy
fIgPfSt43lCtIR6L5cR/m6xA6TcWZFHvJv7/Td6AyB8PquvbCGTmrvwmOmTi0xBH
43tpvlIRYhVmT/yKxsKfBzscMXtdUwYDIJLD1jEw/Od0C3Y07PlqK2LdGoRjh7Qi
W3ENPtN9xFWUy640VWS87+83geEzhmEBacoLNJ1MaLlcB7S3LqXrpQe7d7NoEwLz
5BlNsnxl8612LjwT+/4XoQu7nvDLAE6Ej42qDHNMBqqy55OWfDVKshofo30CThyJ
U7bftTIce/MklDMf3NfM9EGKSYpJVekAZZVYztCu9OIPVeT/LRUYrSJiuZ6fESI4
SnCe2SfiYXiAAM55IACnI6eC0T6Pn4ZLpJDt1SPJP17TfP3XSVebVgxUIl5lfnFF
Iw7s6ykuvfg8mNfCqROeiFaY89ICZ3Rwb0ro3SFrntHtlazdIm7Lj7R3cdy2GI4m
EoYDxIEUnvNnU0GmfBonHVnFNZrtgZe71ZHbKD75KQCGMBXdQcEhik26vJmIP/zR
KyUof0wtdqmulHGBk5SVbEt9zx3h7cTILAn1kIPm8A+QtQjk3j9ipKIQaNUt8xsY
aZOSeX+XBKBjQKbsWn7cf1S4NwL4iFsjhI6hOPLd6eW5Ktg63u3mFE735aB41e3n
HU9e25D9bEildnzk3BBLxcS909I8USIlu8DWIFEgof1OZLPfwcW+FLoMUZZamxRb
8tyyKPvkCylyikLwBKAlLKuMYEVxBsd1yJLfqBUFb+aSB79e5+1oXRIyRPn3/PXn
B9TMxpFsm47CvhQ3LlzFAQsGXwlBy1fwnGjpqAQgoh4FnIBVfyU9/jNpXxa8L5Ei
jK2I9YPXsQI1SUnRidcrxueUvULKIivHsdhZhH9t1ipnHoD8jX86u89fBUhUCCqu
7IuCTYUZODTwXGehL091YjJDYS2OkZxcmA+8A+gDogj5yZOVZJk2k0dY/W2pZKII
Sy7TiR5pnuUpYbzyJ2KyvsTSVI8fX+j0qU0GqVWtaRD18QNfeYl/CMQOZyq37e4b
r+Kq6bZBDItz2PyTgy2Cx8qQMtxg5auoWZfEszZLosYsE/fcU/h9n1aR3kGPl7Ok
efL8Mff0tCYgw/+2bbsJ6+gWqxKHs/nT6pENEe9xgPIunwkCdnecp7UiUEa0kliy
OEjIwVk4ytwXQ+FKLvmIAkHHZESwzM6dhdtBiuHaOkguvhiSI8zU9zckl9OdCw4e
cVrFx5DTf20IorQSN8hWqiGGwaRQg7MkhDtLpJeZXzTwYb4jcNGAPKXlw41jkdTH
JVrVuJZADoJA/0npL6OGVokKWEFuFJLoP5yfXVUN6y7uWnQDMnNScDrLO9QQtPaQ
+1G97YmKJlWtSV+bsqXUcZSdt0mxPWc+N/thfsNPMlin00xV7xEdRK2AQ46+l9O5
CySJUifxJi6TZJv3DXjWAibPB/Bmerfw2MlvZPO0CPhjiCTrNh05gIwdLbNrnvtB
JvaRR4FOaC8ZpNU+QAU2X3WhW1u2xRU76slK0QaRicli49WZccs7SsaW0ai9NEzY
mGZ9I7s3h2oFU3uO6s5eVmf30nqGcRLkagUeOxesMPgOnFAzzMN/yX9ZMa7C5VhR
JDDdFH0uw6qsbeUQGImiREdFJCgSOu2dLGyvnHWbuDjyxTjUgr4L3hzrUs/nhqlB
NXbs4Ga3DYVFlXlYTxe7oYsY2mlTvsQn9V0kf6YQwX4MAN+JIrQzfOvtzpqInm1l
uQ1eRP27Fgo3xcRZIcvtpJDNLrxS3gBLazQadaKsOOltiikVvFetY6JP3JxzCuQz
0utF3g7LgCxhL2od4vV51fNidauf5NXQqwkvJqGaLaoJZWWwHQ03D5DltOcGw5kG
FtlpnAXPrf4NTtPlk9aOMHxbU/F1ZKqivl3p5AlOrB5vmvAI1Da0JYusN0IQfMeu
ofUOvf+ZT4mi2ubcza38yroghuxfAlfv7/TZwPTSw9dsXqvYa0rXAM3X7LCQXtMh
vEBszkVlZ2TePyLrZLPNIvLZi6UJ/AIHg3ufN0aR4cz1lzBP3dv4UCypaMtr4ZsD
rp/1GPvvj1D4OTqyvyuYM1NYM7GsIXIaMtBTE9jWxrQme/QrEgoVtdpkRP82vznV
F+4g96ERhY+GHFvmJIMSKoGWGsv3NTG0x30XQ2Dtytz/6kRiiH8CBibI7kHcVWw9
hMQZNZVD3jVFK3XLeRoxkGaQ+brfeQPJ9w99pqkRQI9D5BMo6aYJC1TJf7PcXpQ9
xUwoFvakzk+OO6qmF4MrsnisWGnoyG9WVD/ZaHa3xBUFXk7CYmNmOIc9a+lAZiYR
WVDLAm1kwDYPRywxIfcI5Xpe+f0BFzeckGAWN3Tq0h72HXC+fFh04OfOEILdBpEE
H8dnLo6ymKDVdm7JqmNOnphMdQ5puVS5Ea/P1aotCEwiBTYsH1+erLB1tKW5hi7t
lyHzcLuL3NEOnHDDZzGXqsQMncT9XXwEIaGpTkqkkTx9gMEnIu2AR0jyVZrUmbGt
RyqkniG9wUHGLBonATmxLctwqm07uDVcnz3peIJE2aX8qdjqCEO4ldV4+Q97kgBg
KdwTH03o0hvoQIQ2Dm/p2nQ5tu42djeLBLlHZs+gdtvJ/OomKdP8VMu0uHUkLhmf
Uh5g2KoYXg1FD4YhT+uJ3uXqkjy6fBe50O+gwAxx9WvisWlwJDRZNGXdhKEcSWFe
vVtVnetyiAC+pTsR83wta93wy+uYU3Gbys5dvuFL7rFjNPhndLUBcCBxoD+1Xa/K
OEmCWS9QFJWmkmS6Zc6PCM9s133gosFfOPfK5soMHI2aienaYmG8kOvAv1Zmi7/G
gfv8JZ8XmZAicP45MYyik+QuAzLH0sJ8hq9X+Z+iBYWJewaMOO3PIISdqjXlkoOu
AYF4oTRadLDdCFMSmxKifWr+Tj5+USaFFgRm3CnXfqEmqNwtwaN2SE8fAs4+JREq
bMHJZmmXedH+82+DRHOPIRUJAPeSLgAqor2ZPAAh1z0M8PurfYZ3WZXYVHcvsTm6
4zqJnZ+Z7XSsVPYRu+VAnC/ReUtVgt0WtP23fq9Nds4VV0igFMdNqmqs/SpBegIM
LArIM/OdLcRagZ6OX68+75p1RXLeVWlWSvoGYhAga+xxfbzTW3N5c8OI8UKKuL79
8WnqHeaxtvsh0xi6/ZnYKPHBZA0qzstG4E4PlcB97/Ij2x/aET0q0YJi2R90VfII
OCAe+XDMMyze+rDCiVaWMvO3FvxRcrWmky5teY8FZ3rd0AN5mFRDTOwVlOevT6FY
v2VOW2S8m4K0t8UvFJ/xPVxkz6vAW0iDbzhe2tbziT7EDAG9m8kX46oC+a8VZlFE
wJHlL3Gi5fpSWn/p0i235CC+3g/2QrM0nG+0jR5OMHzhBcFVpWZLuNAoG+fLc3jg
XVhZaDbh+eiQYT8usGoy2xuI3uw8vauU/kZ8cy1kG/DFBsFoGAL+ndmObwjjOueG
Id4dAfGrm4TowXp8Zc7l/SXozgQvM/tbjjlvxXOW00urAi+X3LnGajizSygT+2uG
KZaiWGByLelA2vOF4uHpaUrJpF201rrrA3sT+WmRIIPH/wcuVqfhgIdS1drNJTS2
4M51/pAB6i1EaCB5h0DQbBSefUVR838RPVKQbmAv4jhn2W+BSDrQ2U2e9JBqM0KO
EqQmxQU9NhZWiwNj9ykcAg6piNxYt9jLQkswL2rl0RmsWajvtLNqpayk154edLXQ
1AKuLUyzLUCPPPVrF0PTh08YIBFnparffJga85RcVZZ+02xt/13eBoTYKn5Ubjy7
KsYRcRt0L/Xyd7gt0/LByQ/TIYQANd5pjQkyd20jHvVR0Hpxcxbnv/2Y7pM1SZu6
MTWexgRDwehMkG1arFjVkCaXdpZjAjzWvTZxQxEIzfuTB8OL88OvU1Y0rayhtESg
z8W82RzzVFstgh6Bl7eCnF448HwV9QPxn7PO0UJ2aWuTkkQA3nzGzQoG429/6+ic
C2/JDd6R24NdwAqiHprk8NKknqNdFIcqrnmSClVpdbusA7kTvxnEqiDbP5JntREx
DbHRAjJYxlC2swmsVTc7DV6qJ5BwWoKqh9hpLsuyjT/a5oMIJU+e09nDuoegDdn0
3Myq+AU5XECHENTNLK2GyZev1SqbLUP++HJuVIZXzkEDemVF1o3CX4i02m2TU4m3
+AWDnmhdQQveSejIIJrqtot7IvKIVhwNsE7XkoXzrxoiZ4cHAjo2/ybKgy7hNUs/
vADL/Ozy4KmnoB1Zqg19MVHryzPDJiaRllzwvK2EQEnmnT9JaQ72LclNjnPlkhoe
I3TG3PTOFz7hmLdlBrEB6jyP+Mma+WxirxDh6dspb1YAznNfQqyC0nPaoCOZHhxA
AVua8KTt7X5X3g7WxhBQattUh7vlnGRglZntenh56y84ZHVKnlQiedIxE1MGW7YZ
rZ2w7CGgI+YkMY+tJpXQR0kUo5kZiNAnng2/Swtog9PGoQWqYOsMl5CtT/2eC7ly
KT4RrS1iWh3+aWtn1KCxZyr7wxSI/YLTBzbWBNQ+lnIZiJCzAWbBM0QR4PmwApOv
v+PcpVf9Gor4sxGroZFQEZDUIAbdkL3XhMUzGhcfjtmdHIoGwJoI5HGbrVR0OvD/
4xktbVTJkyqNYbVE4uCLJcQF6DEJi+RKxrm/I/ZtbMxvvKo6ctMFTdioKIxu2JWs
viMCsMe4zYQyeoci+CmZlb9vfhgTYqj2N2jrtWW2ZMKJ64EAiTcjSBZYHYOngmGW
VJZvcHoKd99Pnu1NQ84RxPosU9yBdmHvEAiTveOyRZpBhV/Lmx0mVESgVmMjqxon
8cfethKzdnCiwDOoFFzDMflxBBj8hA10b+iesEwdeFMC3t4lj77/Vwxwar817j8t
Bnjhz9TAlCT7e4k4mp73CvU293uhp35pzvqyUce94az6H4xdmqcnQYWStzgTcEO7
vvfNoia8d4oyPqHtDiPFmh/800kGDVDhPKBmFkkDIM1WQgAJnMBnJCe8jK4Yyo13
WxoCQofmBjLmUEiaGPmqNmUSuYsItBzE/wGXODORMlLNuUoz0CQxEOXpR47cgPsV
4PxB5Xz39nScOjgHKXWGQxWZt2/+c2h+rLUUIIUdEUFHzIHCz8eRbqeRqwc0cTAv
Lj7DS8M6DpTR5Ce17SLM1Swzxs2+IbFI1Z+JIw5YqC5YRK64f0NIgcohOH08w1Gc
+YqEYfm+SKPQ+vqi7hUd+cI6IeXI5kFXHdyBc32/x3wqf21hTCD7uVL6HuJWCF5u
wtKPn/qm7KFUR0c7ge0+t6cPMAhQrIhJ1p4hXQVvH8E/A5WFTAVfySwfryZ1pbjG
vLa7V+G35Uh4e3Q0BBijTXKgWwI8wSiM5aEWTQCuiuX8PWP2qG6+vJevxGMtziHy
s0Pr21e9uyi+RK0wbUzRzH3lT5CDpAvKkkmV/5KtTSGDrv0HvowIXW70Hi+BwXaV
2c/hXCwsGT/tVt0pr8Lc34keI3kL0GL7UrRVJCTypEhbJLG56B2eXZCPoEyn4/Sk
NgQ8SJWmve3ost0fT5fbUJhP3W0R39fW/PlPIu6CcvZciA2qWdNajKhyyMw3zSn6
C9iU1vmpgW7kqfYJzGiUUPSpKd9wc3coO3mrQJHwotZjvUiEr44mrpfo8c/dKq9q
ykaWPqusMCrmMYRJyg9NCA8OOjOT5K1i5VZiRNpXzNr96M0T6KMJkE3Kl7GEvftx
s8rvPqF+jM0Yxqzc890xdBlUaxGj4nYhYtAIQQtfSYLvJgmxw3u6fB7CpXgktS+I
4vWp2cWVJuYnbpW7D9pFE1RrPMJPxhAJ/ClAX8snHG0JIHTV7qJX2zDXV8SDB373
tMGugnTSrG4iYCIwb6pTTwVrFbGbzbJB//Kqasj5QfiigDHmHIBqJMrr132iXRpt
O2TE45hu3n3fC5n3eN4QkFn+1O8CBCTDCUc+mku9lf16cY2nAsvccfCaehoS0LDO
Eom3oQxnnQmxQ834OdbI27gXn5+2iSWcU4zRyDgGvcp7zAA49bo2Pqq0yF3MCHiH
7i+FjmzqXX6P+SVq3c04gUI9z+EDlXf9MKvBHH2ZccaWQ6mh7gJ+zxNLPu2andAh
AZ158WDJXSRX+aF1bMnCZdY3SZRy+fFA+HcBdaIyQ6jWsFVlgQ062JXKBvbmlEhi
8jn4cTbw0cVtgZFzImcyVMpvmstd4PN0zzzRruJzj7KgJwY1639hBhuP02BEO0hF
a5QJkb9V7fgic/fPbqQJtf+JWGyLcmgzW4uNflFincLVVvbRiefxFggrlr+HNhNU
h7e0ZfIFmTozDxV/3rhvW/zj78yDP9qrT0038Pd+mQ9zAy1v+mBTRLdnkIEObCia
1MgSNP8lxFXzWrft5FpdW+HZlUvxoNfiRjB+GH9dNA7/HPyYLLkMIPAE8ylsHBt8
b1QDWNHqh8gX78XCH8K8xE1R+acd/pk555P/+cJnm8QlpSjq7Ij1yv50EDt6DWRe
/4hnsKKNbjWp9FNvqLiQByn8GJYaDuEZQgGRdIGiJFbx7jLVPiyCzEop44cMNiq6
d+nrGhWxhw2G16yD+TqMJPJQCXRwo6kixb4RbsIahHNEzYMr3jm2p4r51PahTmV2
NTufTA7SddwECr0g71i1OLvU+fnelF0nDkuBY0Cd96JOhFYinfwhOj0+Nokktro+
KNJG6JzzKyXCRMWSMXIjiZoKmSvw5WAn+GODTWRJhVQCRDgul4tyQthIhN6O8tvK
w/BdsiZTrJvzayY6vaSSXcLA3DgOBUCtL2IArlAdjK5XZ6H2xtc+XTA+jAUkqYdh
prS/nFLiz28MVNwoxhMQmlsBe/J542GjUXR02tYjxjlbrDFRyT9JWEOLTooKxyo9
cRrZPHMrWJCTmkSyVPkJwtVLGHgVwVL3eTn8YpgTikrNernBl2BDhG7W9Pq0g84S
R/2a0vR9rzVQDOyrsgwOOu7eqz1iPZqCIrd66gvKItXtlPTm+c26X/pEQiFRunqT
sKcoTepRsABJhuu/FScMi420DperxtoujeI00DDocMV/6vCfHgSw3tCeKPXzwFpi
sdE7oIkZbMG1Q3Rbzw/8vPqcx+tHve0fXNOQEHn+3mggzNsu2HKIVNybVbsiN2vB
vPTXOCi9pRyLYnmjKQrvYwwEDEtofdSQDm3VivurDHFUkvnIkhzC+/Y6wYI2bLZU
rzENFavSggzPflcUSeX11HMN+hMc3D5FVkp0Rky5pca6Es9KvA5xO8xjtk0RQ9QZ
9l2dCwP+vG6YXuGlcozU7gNi7ghoLrLPnTITCyZr14vvGBP+XBCzlCBBCvEvrwS1
V/nCRbmk/96Bqb982j/TBePHEF8CTASswy3z+Pj/H3/KjI/Syr6OmMHY7WlfYHbu
wz/mL5dXVtWoqNhEzsVJMp8p6ZI2WZDRtbGQQlds3w8sScqGThzP9P5meQ5B7ZSF
0WNqxyvxVwl7tyKHhoVCbVVKnvg2N5ACdke6RUIrKR4hw1reeSUx8RkaoRNguhxS
j65xLXfyzEwjpvpcJTQmOxJo/2/zXLFl5c4ddlx2TuvxdWpMH7OefhpxkuLVXLky
WArsklxQxWTLVj+Yuqyq7qUFJC9D19sbkHYW5JNems7P5u3VXjBO6JvSXIt4FPmr
FoTM6WYr6zTiLVSxHOO6NCn9S7Zd2VINnhSAMM12i4quVdm6pzqNZfjZi4b1IR+c
eeiR0FnF1Qn7PSYT12ld13X8ne65OumHdqqnc2AHZUOEYmKBILRLjrah7Kfz0nBB
SSYiK0YzPJ5xhOGZBnlL3lyfVyAe/iUKtPoc7R2fFxCuUreA4NiXOJxA7iJfWjGb
rFF+vNmpF3iiJT6T3f50Fc5hPcVLq7rg92iEoNlrIuoKwcTZFORZasplUJgCwwFK
Rd43xjQ0VfwmyDYjBiNjfjitWbvKh2PhWSNmofm/vzyx8GF3yaur2FILY92RhpcO
agQ+w1sMbUjj24AoBvEKPWiRCzCeB+tZOkNbrcE8V7CoP9Be0OqrGMmnqAeZqr2t
z1tFoC7rmzGDdRJYiFtROZZy40InRLk7PYY7p7xeDmiMvelxW1sFSdQPrGVSTHm8
gCgdhoMKPw2W+UusdxXd+4rIkxby/5NSzXAvJ6UAl9CBPQmTtpqXtzSNtiVxbDXB
ka+WpEguXzofKeQzUuZBniFFJup+Ch2EpHwWHP5WhsKbE84On1fKlWeblc1KPJ6I
c8eI632Hjgg6MfTyGb+M6cuNStHC3cLNxCz1gshwTi0L3iwzLXU7bBVKsN+iD83C
cSeG9bcFZzFMiMa7iaS8ZBmW10XmQUSSizyx7AidP1MEoD5Bh5z3V3isOvR5ryXt
4mHh0l9ttS6slesa+CBT0j+K5KfTD39A52cte/MAwzJ9B9Nfa7e3zzg/wGmpqbfi
QfbmHZp7bjEkN7MFsEmqBAlQ5K6/5O+zfu4/26uwguhEATVAwZd80/FJI6h8QK6P
50Ce73oRxMqiYosT7JEkiaqDcbglPer+SCMZSGjE9Rzn5EkUu7TYxouYqiTAJ/HO
KBkbGOqZbUbnxoxgf7fY9aznycvSbk1d1sqetFVtQketexLDojt9qzM1NScv8gFX
8hBdIimyRD0guEyZ+bObjDFw4dunUDeZ4YQGVLbtbA7jGWcD92cwym0yLyQ1bgbX
05hdp9JbSlh1F6tCPn7ZESkM+ateRZ0PDNtmhETEId1R2RGyTvFoNiprplQRAU3L
lzw6CjR1MH0PF/m7MmfhzEWpU2P2FzRZM/gh2SXbAzNmmi71jOjWGYCWGBOV1iS2
8doA5jqIxORQ+VrOAPUkBwdGGdAbEVupqZM2RKvmejFvbU1GcBr6AanVc2n3Qb7I
TPOyfc6EdWsVj2uzqTfgEWsAoTiWqNg37FNtOPKAHeQQVA78Re0MQl2jD6RSdsV2
uc8db2AYrsjkA2oRAWrRqMm8wKIUquRdWVl3rOIr7xt6faEYSF702BGbnvHh/WE9
dw+HO7qoSJQ3kaOSVGb/GzhaHl8iJ49RZKqtxow5blS9K91p5XaYqfenFLrX6d/T
sWunB7+FdGmZ/OLTOr4+qfEPsXhlkLGvMfcO8bJr6+aR5XTIODYt5USa1tMheeHZ
gXL6rm7Ko2t/e5sIiaca4hyPqEZ5Ho5/qd2o2cpyA65V4XD3iSvr3lDbZ2xCivHM
VWhdAMNArdLYmYWQRRu4VZPeRueLBRmSlUSpDxBVHld+Nvq8FYxJYLB2iv8Orcp3
49cY0bzsiSevLTKEUqagFj4sXzs8c40/0miwZyzxGzsuCWA37gwh/in+ouhq7jpf
t4bRba4uMlpjnhiSBS5LnIFljhs9dmC2RoJAWcUVMOg9/u40PU8gyBdmc6xPVYoL
K3zQkAOzPhlN7BX/PlFDJYNXUrGdu8Uv9zm+y+yIKYABXph3c4Q0LFyN/dtITX2Q
szy0FQYbzCKDj7ELGpUmzdeoEIjk09aN+dpIrZ1GWFlBK1GMHNAlXGm8Mrkins26
Mt3amlXwmyeji6r+T1/044vYWg74b6EGU+v9ThqHMvbKgNDPSaAJMXY3uRIBmUdi
/rPzZzzTAvxqzPIN8VCiPTF/ewiIX3apjxqxJxryxjJJFOEZSwn4KWJ+3HJRCdB3
PJrj0Jq7+cTbWj0cGBjSbBFLsa9xOadEb+r9AvScmgHE8vBZWavEybYhyugKDDRf
yZKcDJhrpBljNc/yhSF1qdavKxpgKNZz8+cIOao+QhGMcmOxJhoXHAMdg1FNdSdw
DknYrVR2JKaM2P6ropxnq8f90OeGLqJvHBelufzeh1cQVUIC72gf+hvI05PJU9Tc
kc9qXb+gwikfegwRM2c4DCQelYe5B2u5YzMQwXaL+BEBICPnJOBlyeKqvKEwShmM
EcX1ooUEMlL1GaixUFmpbNcSJFdCVthDUruME4Eleuiko9SxRxinmpv6czHWKww1
/r61sfGm15QbTqB+22WGOwMe8AXloUvmDy/Xu4aobJ1hq6LQ528u4YPL1AvHOw1R
AutCj4+WDEFQTSI81zARwcxtZRevh/hTWGhoDid4aK3dpk+68pFD9wBmefU49ElO
yDpRq8HaP5GKHreqE5UMcjS4To9BLjZEokl4e0TVRDNQptLEwunbgJybhXpZyzfI
itTD2QdD6EsZEfytE8NSKZLAAIj6pHGnUI5OADSkZICL3rjPIJOn19VhRS9hB6yf
ziHzNuEo2luVJdDQMHOiuB+brKPFIAHqfudVwOxHCR0ev30JOAKxmBb+qH7uhPOH
7SdKtifNCBwn9VyoU2nJ8TMUAy9w8xUIYT6RoAueMlmPKDWkMMHFtlJ4Bi4nVGEM
ICTk1n81hjCqBTL2NqmJm2o9uzH4O0zWt64fQ5D/KR5MyMgaD0ANZuvvJlJCxAnJ
72tVRu0cQsklhiwazIAGHofH4a1ku9/a0y8AebHM/Waza01uTI9acrehQA7ctARZ
25EZEL/7VN209iZVyplCQ6K1qfAY7SK/2+8I01YHecHd3Vumg9Wos+oDPE+3kAmj
ZmPkM/rfzqKQq7NouJHSmqq6kv3oIwddi6aCG5nxmCn5fMGQ35aV+Fd4lXHYu2Oq
wpsUzOnwj+6Slkfyz3VK4BX/H7s264rgriB2yO4im+mabDI6KAxCEP5nZzsg5qlu
dRs4ZT87ftafd4AlsB7hmKEm1IHprV6bGQIe/Dc/jcMbI1Ao0/9fUUsCZUcYzfSy
+QjkkXd1UOb1ZrV0vT9UNDAWJKvOM4egURnAXVRpj8x+xH3/PEx4wS442HLLALPM
Y6692Moe7IbPmQuBztIRdeYYg3eI7m6gTHgaucuOA7S6OvtWmn7yvHn1s+I1gacJ
4ncTCk+r31aqp71un+L0HoyqiWZQasGoHMxhJtaqvumCEsvKnPVm+njRNXMWDGLS
CO42AL/VoWfVjeOxdlWFPmVo7cEC21F371FWqjMyyHMrXG+j0MEsSaU6ZdXxPuG9
za3XTwi7J58eq67rUACKO0knkH8JpLyhLqSeLKq3/M9WGmdH1yvf3qWRC+2FLToI
GHiq0dQxc+vvopSlL5J0+RXkawEkeJmhRp8j3wL/lFAkagdEwgAZTNFC16ccuZSi
+ZfoxDKUl0iVGclTATWfnUzf0IBoZxVZBdxSPEjBCrbkEGsBBh0ePnKF8SlOvUyO
fWQQmuw1h/3ep/cD0EWZ0JQjDLWcRTrJ9EX6wk218v0opFsFvqqSE++cl65Fp53R
l8dbEknP7bUonKJK1Rs+sleuGHZwAh0oGohnsLxSxnOKmqhA3rFOf6+GvLhPUyBm
HbK2CrTNSh3zXQwcJ8sNZXNKhTbr0fGJY11OAEbn5uARWukI/p58iELOqmnkY3tR
RaoHN8mb3LcJwt8JdyU2xlIUsj5xLFWXl3RCWmukRGwI0m36Dr1uneQxZwK3waMn
MLODpdD9MK09D9+e7ZK9dDW2TSEX27ns1SOwZ5ap3XpLNKfsSU1WdIQJrq1T04sm
O9QLHtFSpgBUsLK/Ttr6Em9U16OR7+odeCUYlyrygAYF7aWAE0bXPmm0zDFDvH0A
027m9ymHrdc3FPkM8xuhfe2+ONzZIAsPJnA2Z3lqbNf2Frm8YZmOLrsedEUGvKs3
RhL7nJoZc3hLE49UNG73Z7Os9f71yzoEQm49LEdjIsNfoGilFZJNy5z3HrSy3myT
kDOE/n2prdUvURXtruzLISCNR6g4lIg3fjATfsSud7G4xFw5f/k9hrZ0Ei6TAChb
CFVFR1MacKiqlcwHy0rtajSgc6/AUpdXY7+E0QMX4cFUsl0mkz9EK23luOeqVcz4
N15DBBjs/GOnxaPwG1kSd2dIBzqq1wvDzGZc+Nap4Db8efwrfyK2Kz+hzHp3+fAU
ACtpIOjRpvMCPiYTy7t3uyhhsghl8dMdBH48xLmZk0pyl2NiGPmF/GnIECAJ1x0R
XcuulviW+6vTE3wET9oWETWhStXxxqicfHyIFjfxSeYf7VK7Vkk/Ve8AVOKbkez2
yWtQRWnvpwrjmGZf/C2IMb5Xo80FK/8uwCEON0nu7KtxqRQgxFD8OY55mWxsU2KX
mBpK3gzzeyrRU4cwcVGDJI+ogeZwX0EFmFAmzLb+jz4jkJgLsXEoFHPqfx30D8Yt
on9KuRr0uYpmgpA0UCB6Rv6bvtbYpQDO40tKH9aOR/Rd1FpFKRT9edPBMO8fJglV
F6HSL+kzRZDujMInm/8i8LVkiZVdLLJVzZLM3V76Tajdns5UhKebpw22xEe0B/86
3O7RpbFy20kcFVMU8tFkRw7jz+B8iCabdN5TEB80Qyd5+ojWPp7HGEDjZIEBl7tR
r0NVMVQmY1fJmG6IeKKj5w7ZLtyR5Sxtehb9/ImVIkpq5pD0yJufZOtUts9DSEP0
TGUqSkR7GTqG8s2oQhjN1KhGtFfxxcQioSOc6tDLz6hh12ZCnsWonxNcK9xFo7g4
akT62FeV/YoeegGIVXTXHfYZvOQuLpvYl39vfaxU+PGeMP5l2wNSvdyfn/xs2t7g
TuIGH9/Pzlw9qknuWWXf9eT2MNfdXjFcvfIPm88ytGZ5Gg6wcJam4lVXYNsc2lro
aYpYF3xbUVI7x1zimYVwKEZnVMXlv3EDEQvJaE5usNC23+5NIy3RAa7ud3dU9RGi
jR1c8UVhhYZ6pQ/MmKktfd6eJ58pImBuYY0Yc8rLGvnMM3B8u6lGwgUE0BLcQnaD
cpOHH2xcO2IGnSRzXpOJieqAu6wiPv3GzIUqxIeXMiV/rDGIczyMVFoEIXJBsSOj
fS7H3k6q19PWZ4Y2kv9u0bvrIu9wRQ1a48GZW4nE6mJczsyvLVUyvPfDe94y4tnP
7/92oYJxc4EbZrKGmXVemn5JDLQhWs34K9SeFPeaeirEkej4tJYpVgJYRCz7BY7M
NAcV66mHQJ5YhxYFagk2SL47DifRLQuh3TCj4Kdqivyjx1hPJb0SF1j/8QlEWfHP
dJcxagneFPacSL53LzzIvdKJ19sd4UYZCjhR5hcOEdMOQFRCRxGcMmfOPySCkmSQ
XhQ+PAIwJPukw9D1HFxMYUFE3qx+s144XHPeOwngLee3oFP+0xmDP/oRnkqs/VWS
rBD9rHtFgJmPDukOJvTqhBn4bRWDB4rKO0quSUXu8OMHL4gJVfSAnlQeZaLIN4ij
uoL6XZeq+dF11wGB0eBmuS+KqZ4G3clz3Yd20/6kRwcmGyf1z0dxff7jQrEz8xW8
hse0viBnGQ+8ZtIWSQyDCr8VpOsSr4XM76w2A9gl/HtYPxBYs4UnLTned6PyevCT
Ezwdf/FqMgqOValLwZ2nnvGISjFWUtgpXte1ZSlo8CHCjpcCzT2yI5lNN2Tw+kaT
5U5v946FMHF6xZXEgFx+wfEGNSrv3qiBcwQpZAsmoP0h6nbVcNWzsgf3b6A9KDvs
F8+vRywohazXnCUnd3xfWZ/zCDa5iP26TPNPxrNjdKpXYs2Rgsq6t3kwfiFnAaEn
hoZGam82nl1+K+gCT5sbq/IkZA5uUhWYkDR3EhgyalhXVmTNwmyuGt2hE/jLOSWU
rgiptvEEmDNc6NTPyBaNxURpRVlUr+7ajL7c+vR4c/VF34sXCyJD7YJ7J1U5OzGH
Z3uWLoOS8OgsRduM8fJzALzVILHeqOFEjE47r5kq+dP1GtLCOkItcDRI6jWwByQt
8/X7sGZ9pgved272hYEYyC/pH6LEJ7kpgzZcbMQe5teEC7jxm3nUKQ1CJbGIQAGJ
Ulh8SAmfJiGWMfTw2+rAVk8GFTSIR31KD65pQEOrRTmxtF2DoeuqcDpwARl7ymH7
UU4D/0gKgRtiNyVyQ0HBbuy2eutHK3NONyi6izithwV/a0FF+P8JHoGVztPZ52w0
2hRdXQiEITmjQHsr3/XXokqco1j56aPcYRNeGLBaMlXrg0ScvchJEAo0G0YfKskH
kXv/my4qB0PKo6dIwcaMPPx37kbK//jpTBDpsfVxNsa+o9ciTbiBm/5OZ+riG9wF
1trPsCYn3kmm+k7TcMjVxQsGafj+fQuoJ8DJTS6h029FAfiKFLzPIBJDbz3BuxPz
yIfjanGYILkqzMWZIrGqGZNrwdaHS6JCybibmjIB1wl5Q/OasYDCfSMUPXILJyWU
w0+1NUrmejTeMg2hu/4yU99wznLmcqsZ3VO4cUgTzp5TP2qL8FCoasSZt85VIwt/
Z7qqqK3lhi0OEnlWTUzZ5zCj9IpLa1mfCmtjR/HXGaLLp5ZzkbtlbAGF3nJCYZ4r
xo+Ffi06cedIJkAflY0uURUCI6zaovX8jcl1J62D5PF+k1oFqFIlLjEMlHwxgQJJ
ARsU3+kQanbJ7COZHcidcelDG6+xV/CTjnXNz+kdCguRoPXdZbFO95Dv7XKCdsea
8cg5bQNYsOFgyXLFaV0vAk6T8kirgbM98p+vlMwBMgIWwXPpAVd1mIwdJvW27f8E
lhpxOw6nwfzfw649EtKfPcF2zVuBAkSJCp76et42EbZxno9GW1YA/b3gFc3DggG/
ePVvD/Zy0HlIm+07Eys7t9fEhMu+ho9vOFduaIndEjwi6nNRFhK5FwbGgsAoSwMw
IliLpP6yiBA/8AwTuJKA9jTLTu3XEyKs56o0heVTbkrEW+Kvx3FunyYho/svO60N
LU5NMUSbIZCKylOzsVQUQ/h9jmFOA77KjF7VEvXeNzfqrsCDFOfFdIqqQ13191tL
8rxK2Sa52xRLwiiww9Aij0Q7////awMwqsxC8z7E1vll1V/zTuOCjDkC9TYQPuLE
UOGsEoUqDgx7xTnyet9T9VxKY6oRw5ISQwG+yvAMCH5SL1L/g82CUXNtpDzzg1ee
EeVkQ0z6AnFoHGi9VuT0nTHlBg9bbNZXRnTMgjirdaM1b2e0+Sq22JJlr8HMkpxR
eCWhdgWJ3BD+OV8mnDEBiymPwqmj3NtIEbvJwWId7RPRaEpPW8w8G+XnUpVMmHfE
2PIV09cztavFFX9S/cd82kS0WQWmo5LM4eWOYj8eIUVKDK3xT32Fw5odbMXW+You
h1Tr70fjlsa0dcvbwCHHggER/vGwisuQrHK5EwwrMDnOL6/SNzpoDpgQ9xunYNwz
h7rsEvqdqXsmDpQfgGMEC0AvtyMFB4vAU9ictc5aNxbO5LOZTW/uWbtiXxbFBHcc
7ls/gG+n7QBwT19KLmh/AoA28QJzLZ+aGX2NN2dGguoBgSWihKY1VRjwjiT50VMF
jgsZ6UBdOA1Ma2dnJJMJ7WaNLPiJx7K7B57SUsUaciyGNOUfof+60a8EyXy915rb
ZoPgyijuDrrxsunTWkJTR9scTVi1QAO4c1N8b5Zf4SqUDo6z2fmah1/aPOy+11O0
YNTlKp0TwidQdWC+JOjiEYg8f35IKbTN6Pi2sDTCcE3ASo9GFULiCtYGN8shqTNn
q/V+LfYs/y8PY5fvCetck4i2sjTSaVJCPi/QeDtF8lS1ku96o9VIiUplPhPIS/Nf
vLva3jeGiEjdtKtpJE7YtAG50pDKIsXZMmMVL1LDPeitr+jERR4FTy5NTovyu79S
sXhLiMA7C8QoncGVPr+ZddYys0NGSPuvePnMtgSUKpGWNzVVXEqLv6t9B7u6GGMd
2iAbzxgRe6er3uKMhPiDztaTfBFUbYN4G74k/yOy1Ua2NyRkMRV3QVE9udjLdpFo
xj42vGIPvC1bzTE4Hx5WZd3HxEWPxxXm9RC8/sqP5ZGitBL/ZIitESz7C34BosUV
m92onZUH82J5XMuXWHC/Bkz2ILuUQGFL8/a8B5LaUqsLh+cYrZz42ZcFDA50h5Ya
wJjNb9Bu+oFqNwxZkqCLCZE3Oi2FGeim4Is4Aegy5QU5R4AnCEBqFegZNPkjgGFF
hzrjVPTkKyRQushk/kdv9FzYHy9j6BoqSIrmEtMqQA4ZKAhLUSSUEw0MvLhQpYqg
Z21JvLefdga6GWRtv1Zm+z6d2bgvh43pHeR5lyRvTH0WIUcibBb8Z7FwtqmMdk+0
GMGIrXBTmhvjKDKs7L4Ra6fbYWyxEc4yoyqkGN4TqrrLS21Z2MILwupNejxZFhUY
1+uvcXhMFkt6mkm5D/SM+jTAcUKTA+PvkE0VyZHRlDfjwBB6hofKfgYeXLkyKKAr
JcKw80kpTUvEMLH7/BrRsjcKi+FfayUyzDoNkjf1hdjo0wFbmjZ3aLt5Gj6/v5Oc
CbNOhC/+pLAYqcw+1HN9uKypc47Nnc55d70lt2TvMSAY/yrxYYwooAZV/ebD8GF4
lVj3OKJPHB+oU5MdFwoPz2JB5HYCQeQYbsqoe96GF8SeyTmBfpVFqr7gEg+sum2a
peGTBrMmkuWxMjTzhjAMYxrc5B2nB6dX7sNYs/KoJpA6elBvDGGa/jzHvVe8w/zf
QwVuXQZvfB/GN+UxO/3eHXnMKWrB86gsAfCuBl8n8iqERe/EyaAaby6xUrdLMSWY
8DeAPoeOda5kFMYTqRFb1uAdpEOxngUfaztTGru8locAeyp2+c6gVm1S12r7GwiK
MZmBZfNDhY0W2fV4mhTWW/ts0pqGPbAKlW5KoczCUzLA4Y6w8lWCxXByNSN3REU1
plbDtbYRnqsWeE98Iv3DvgnCRwcRaXVI/rEnix5j7L9fRuakeXGIt+cCqvr8hBQj
GsaGecT8V0axw9TqhJh9hcCJIbf/2zqYGEdi+DpfGJGpRtvQ3V8bCUCsW7NKrvSl
0F72rYm7QVglk3wuNPWdTShKDwdyDGYRbWm/EuxEYfZGJ+BQ39QCiBP0uW4Kv+2n
orCnxZfmmRHzJeprkKK6Ct4qHr1t3ihvvNauuMoPYm2xCf8xRMUf6HF8gdFY8tbb
0HfS3JaYXY1DwFYv9W3UKzobeePhBcUVZPJzswE5ZAxCq7VYMwJ2B+l/TwOjLOz4
AaCwf8cydyuhk020gaRHrjtWFZg8HtJkikuO1yp4G8BqPGCGCJRXxwgN+0+XfZui
rjiRwddrMlMfRU4rPnVnSd0WW5aO8RAFPSMSCTBlC8U3CYxVJys1ZwxQ7CNI9kPj
xXNfXnUZ28a9mVhK2L3/3MB15BticsQDvEBL0Ocnw13OYVna6mfwjw04fk9tZlI2
m3zop/6iB4MZFZZxy2HvWrQ+aEhlBNW2AXxppijZqiKrCbsn2F4oMQ2Cih4i//Ji
eCV8R9L1ubIyTJyDb1WWpNkcNqDulX8tO3yzLQ1vTBoX//1PxUTqedXeweYu80d7
q2FHaCJkYyHzsfurCXBw/JGU526Xy80WEvWdgOzH2zzAZHmwgYkj0gL79cguZSFK
oXqaX0/cjwqa8URYvNQ3qT5z6+rAMY2soGqq9BUCY4ON9T60k4hHcKMCOcSp7ozL
2IUqAp2ViWcZhT2TQVWt3G4EWA4hpM9aNjE2fHnTJn88hT8IfSYgKd4aYZoIsNRa
aMCdmeElnF1h18dADiM5KQ+LVhfZKFVjahfxyfomdM3/Wfq9oNsjQNihnY4sovgj
+++A76zpHUXUc9T2b+o61AKcSwM73KDVInbOd1lDYS29h/veloXMR4vuAlEjxdXd
u3GzDgfTXcCFHJtaC7hhjPE6TJqD2A5BNvl/5QCDtEyf7QJoXGQmFsG40AOuNkZq
LDSkOnWdX3gX4+ews6q8dah4WNNbT8ewmG3nT53j9Ums3G65MPpxTbdrm60ldltb
kzvM2QMR2Csgmy3QwV+2ZPafTic6QgvkmNy1tFnSO/xfL4jRdV8lrgUWjmSSupPn
JCfjABvn9pTwLt/uZhWE0TB/DYBKN6417K2hQPSQpRoClBYEWKMjjMcwH6NByHA+
CK6bTiqo8xWDSfLbLYwKOn8FrKS1JT5T1gnfNFcUIOw+I6AhOnsAz6+s8VfJwIhR
ha//qVx31i+iWCNuu5O1/X6Q1r1Y6liFAH7DEbn/FoHnd4ZynTosL9VFmLtsakkv
RV8A4K9dG6i0aNy3AkxAO63RRFD6mSfjApDjHRAUQuUjF83zOHYWA9P3qseVFHen
VH4M/f2xn1bmpm8qB7liEucetjCjoOeOq07ag1mmVXFfY+If5Ncvypkg8n5jNU2X
fRxqIgLjT7E+3A4kI3rGd7+8fYHC7a3jAMDW1zuAx1TyasuchP+Ed1HnZnBumBmu
59a4M29QShSJ7bSkFj2Yq414apYboJJNSmPnpR/8eeOwksXFrEk2nHo+b1+HgawY
o1ZNkLcpk4pGy+B0R0Mi8gtd0Xgn3k+bTbHoCCKFpHuI3OmAP+uWpVxDR/4/9Ryu
VjlZLUQSAhzW5BHgrIZJYTo7tcE9c3wMN3Fc3At3ui5UJMy3TikcssGkBplx8nLr
sYO22JtrCCTUMg9liBDayddbxuwqBVtQbKje1L11ou1GqulvrVudXS3K7F8PBLNf
Zd7KbSSGo2ZhnBrfE+6bcDx7oIJSNQDWjBZzHzuegrjbiRKvL1BMHNhPwkrOF0XC
3PqFOKCgVHdl0ekXnSnYR49QeIc13HoG44RyzBPMWLJy/odrnDdE0PnP3wdfXwd4
VxACbcjHQ8A26hOEtCBE1DC9q9MNXahk5bNMImzCHVgRcamKjH1ktXHi67XQnAvt
z3kFSHRmBU89GJrsg98TPCGRgW5OX0rb59BZYSgXmz/sxVjdez5Ym3MGCU29NfOH
cCWKUPnx9KVmGL7XsavMmrf5Tgt+DQkDOjXZXlJ4GYpf4n4fni9LJw+ywSr/PTUp
Y+nl3oYgre0Cr9LpwGH0FnvN3VTO/hJvgyvxEcmHk3EV7UZ/MI95NG7NmO6GRUHg
D9P996VYTr78wFMWuCW47DeIh0Uv/2khElEVcmFtoRl+8p/8eDxf1Z3toDOHITB/
vuomNshhZeQhX/moT//SBIojjMNJ7iWhYpxbMZ7jm5pZd26U97KNgjxLT3CnHRQY
JfTokGYW2VfdQQ7GAy3I3Swv5Fg9uwDO6EyjZpQ2zGt/BrHtPDbIzL98724UXVpu
9FPGrctHm0iiVV3IdGR6O+1hVsstRsKHWFWZT1NrK2iHs4kByjqEgxB5FxZC1cmQ
LMefE2uHdurh46uVzaAD90Bg3+vkmzveUpIxqQNL2HOw+7HNMgkVOsXodV3ciIlt
7eW9RDlHpB2TbP0zZaiZLTlHIF85rjcJesWxfaPNiepEELatsTHA5a78FEwC8gb+
/ldmZclx695tznx3M81LXB9ajnE04EudUJxQxhzpSBqzlykOQne1UR6+MzX6YUQr
7LmKprycltjqqm57KscwgjkuLyuEOQyI5tniNyui057XLB9W31CVdyL3BR8zlCPw
MABxevP2EB+iC/ve2Vv6e9QdDLTfeQJFgQqNwEN8Nd9zqt/FDa7nU8lft2uBrQi0
JreRYaTG7ao8id9FFhjxeHkHAju/2dRjrrq7C+fSv2qAKMQibVACBrUV37sJ4q9T
P/leRF7KTjqyKz0ryVHHh1udwPb/b05OU7b42YJypIE2TPwFYuBKtqLLFMDPV+py
18Cb14VnwsZlvRUo0e+Hq1C6SvnnMqZj3QMNzsSED5DDT4m5f4jnnJrhUC1jCwJG
eRnawmvvWk+6aXAhrRg9w6VcPrJ2Y+uIxDJ4Zb7u8krnoLUOccYq6I6VQd5AZa3L
X3eXCRosoVDo8jH7GON8KuE4hOJw7yde0CmYy+/Uv9cHnbzb0STJagGZ4ORUo5qY
9HHzS+rYza3KCK/Ddh+q//EnDkC8oaVOZlnLrL/aL6ju67AxMXmFOFwljgiV1zle
VM2czXn9Xj8EZXYcmnxc6dxslQvUfimZ3VmZXo2teMsVgrq9tc80pNCF5wUiiStt
Rt2D3Y/9jcSsT1qor6nYYpqDSqWwBqiurlCpROkaoNmAohPRYKR1cd6n7aUKgCyg
yN/l0FFD3BLrJCZOALDG/7mE2O5rHjkxwjVMcOQEMianBW5oOc0uYJ9CVVOeHIa9
/1reNk4e5+zB92Bn57PMpFs62SU6FCAlku1vcPpUT8io45rD2yfS+/VAlr2JHIRr
/wzTRz7lGN9h+4OEbn3G/eantiLegYhyhGKt8AjplLJhuUXI499nACmk+yxYB58q
syWd6mAKiG9BRGkXSEuRyprPV01biVk9qvMWqZxSXN9r+B5W/4oUFFhawPMomGa2
/JcwrvCSSuPndlnm2h2cuNRTbhh3IlDgZIEBaY19sihSqFikrpXsrNfKeKQF7ivg
Oe41lH3d8JdlQQ6TtY+FhyZBnb0Tp/76eHLRnElPTasjw6fzGSKFuQBCm01vzQgH
dO70i/uhHVS8Kffc/BgzKB7sL0gdMHL5VYdRju6/5h7TyVkDHSoV3sJ7NPR43Yoa
+1kcVrH5JOWnHV+XVwHFdU8yYPoHSPqmsAdvQdt9MHSZ2MHvObghHhmHDxjDQX/D
BnFgZ5kVxWkEcjV5stdepYhnG1d1L753i3vZxBv/lcKH2ftgZ0XQJXPUnFOC7mUS
dxPiDno33GR5ikLo1R9rRLtktcyEzzVur5cTOFG88gfFRAi6k9y5vzUsSGVMBeEG
0qrSoxGcgXrzues/x8ifJT/KeEH9pbzGv8qvcxH8NIIKXYDetccOGS3lwAA1UlIx
HMwpEC2hH6SC5h+lXqxVn1WWJo3Pi3yTlr8MjBfnJ+tffj9sPpAr/CYPFloVakjo
QL3Li8ukS4kynWiSRSxeR/Ql/HDN5ACYErThQfot8LXwU+heJEDJ5uOLgTNwPJbq
vZlzEf510Hoi/hpERZwImXt7if/UUywXhQPSefDxg/NZAIta/tC4g7YIsOnz7P+2
crKjXWZBnfgwan5mXImlVbIyD9jFLOA3uQLumQBOEErgXwkO7Y+6AaB1WbgnIryL
qjQgNPEBk9QI/v2FFKRlqfh4DHv9KIDtmqirq7I43dFu4VncvTQnq8947T8eXosl
BC1yEGLCNoU9mWrhzwFhVLOSzbunzVSFwv/Q0pOhZjTQjH4Leu2cYSBpSI7e+8nZ
rgBVFErFqzhhMQTuJxTufYZFRylf6ZmurfgYZ0L9tSdoCre+j3z57SvFthULHjaQ
Np3FfVjNbjbV7sCFe3hEEgCq1hCmCgtjErTt073QZSBLFGWB4rXgRcwO8fHD3aDA
vJBbwkxUkaEtMPNLf/641kXt72WekDwGzED1+qPm/cpGKzju7wZI4Lq8+XG8r/fu
zf6wKxoLKXfmQiU4FJTmiHN+a2qrzKVInvN44P63ZCSVRl8MaDx58llxUk4vpUIK
F5NyhzDHcDtrHge3Cf7hN05rRldInB/npaOTBEhONaIMawmFwyHfvpv7VKbeTXO6
RksFzvmghIiJgb+yrCWXeMp8p7GuGS4ydgwkEetVD/y0DINleh79JxNPO5LfoznW
sl7mbUVMdMRGc9h91tLQFxXJhC5+sNp2//zhed32JK9E6cJmhlWoDCoX9VB3tqXH
aQvfLWZ0lEWKgb6k9bDDHksGvch1UhPJZO1VBnXGDL2kj7LFNYwJHFmeFkQN9t+/
jpCJIaV65WV0O6+c2muxOebrGozkUG+Rkntbr6koE9Jb4LI9FrFV4aGYUa2Iyqs1
vqYtEacKsznOhYQCtER7pL/+z+OT/U6ytZGXcJQAuc0IxxKpV4FUMPgF8pY33TVM
ekAwWwq1BofnXHqWelH9XUNUTmgp5VG29/1HxIkdrAFbtYR9RkqK/wQKiJH9W/L+
S3c6dBMJKHvYFCfc8W7/bkn0WBaH6EJF6yuHYkxKfW838Fzswi7TcRPLvul5KMQ8
S3/djqQguKSMo6zKeB3mVNBrrZqS2D63GGm+Y1J6oKkPp1h3NksKxyY3YW6aXYWA
28jPmqHrOYKzztQvA+TAAz+YytBU7Oex4mBg/8uSfropPmGlRmyTQRHGYuyjWQkT
YDT1TggYuTE2Q3xhqEZYdoil9Ru+V11vsz6hEwvdK24L7E+sxqC/PnHnxIConIQu
Ubov0DxrGWmcxIJ9jd7W9Gsxj65nu9ay3JAPTEd92m1/ooCDaOm+Mhb7WYz6JDpK
WXkV4TvnBsHh/dbCeHkRAmjB8lUci2oPDg5ikNW58f36aZXhEknOJ8vzeGKTM7Ug
oGHIKRZWjRrPGZtOo/LEn4MzRwqwZT/HF7MjTEDHSOZPqcu2nsEpR5+tcl1RLyrg
btMzyP4JKSx/uXtQghqOcF+l+oIsVjM3udavZnjR2pvKnw5e8l+8GT0YjaiPGZwQ
S+gCpP4N2vznsQEFIWZBykzP4qSxKWwZvdblAR2mmwQY5yRtamD2xI9BKwf21gZm
82A2JyCAUe9F1CKAB76hmK6nxRm/ZOBWRuplAQm84/e+ty3t/jTrEw9tvcQm/PFD
sevx8997HEtjLMwAi7ffGRUMEtyngYfSyPx++M2vXQhvS4QR79rNC7akKQyPveO4
Drm1t8ZY+HD4s7m+cGz326x9qM4cB+BTr7ui0t0R2/TGi0n4hkOTpDDliHSzew3v
Cjn8+TE1fysquSXfIs32PnKPsu3O6uojQnVYMOiqbLbEUT5KrylBomuc6R/2JhWO
hS2gGKbQ0CnO3WA/XtU0QnsjUpKODiL4HwWnv//6eviUN5fTZYhgHCPQ0CxpoUDY
iLOHDaEQIin5P1VAw7xo/z+lXJMVkhFawVW3I2xYA8OPMq9msOlb1mkpwPZ3zTJs
lQLsmFkDpg/k79BCf2MH8McdrisihQOApmYgolDUGoOQFgj6j7FBK9I42Dt3xWhz
6IltfAV7BznKOrSbvduNrGNk8ZafWGXliKtEvjNMav1BBTaq6nQHODX5+TZZGonO
qgiUVok9Hy8x0oxPKVHkdNvK6+5F+zlec6eire4I1EaM4cZ1azL48GansGWJ+gLI
cxzL1oLdBCcQSCBvYdmlzBXDwX9EoH+aDBykeGtvB3apnJTPxKY1DkD4DUxhv8kA
xCPJqSBLyA0FLgdOOeC/zLA4th7YbIG86ZY/R/do9r4vJJNlePaNd12dIWYA+IFr
B/9XOBKrGJisUYgzDe7q0Frtcn+q41MYRCiT7qCRrIWmHVXNz/153hZN7ptwcO0K
0xsEUngi/4eQtGKIIIKKV4UUIjOduOqA86r16a85nlShSavQJzDAedwZ2E2H2eWR
IIGLjx2CqA6VJocXSQbIFoqOJIwrY/nWl1t5fxwKLbmzMg0vY8jlAdD2V+BN+C05
8sG46nSsZIZnFJJZ8EYjuKXMhiVsxGkAdBCmFhml1baYKx04Wt2kgKcg0xVzQrga
yJqrS3vY2bPV08xwWOl04GrbTaph2t9XB+XQtN20ar1+Eo0OFaEYWd6l3/dUkFDM
JwNtv6tyVj7Z2PHLE2Gh4lXskt10gEMrvNvf7Uos3MCAZnPi+kfFEhvzp8WJCxgd
GruxEBZXel8JQVb+OU15EMTkYJpNvIuw5OSluz6lVzyQTPpqfcADMhzK45P49g4T
YI6v0qi8Boqxwv8zHQogaM+X056dUu91atK6Wg4wkZoYSdZEl+LpOUH1RUfwHlql
XlMosg3YL/4HhDOmhM2djORAKYA1f1HVV54BsKdvqmwZXEqmbtq3FZ46IaWiUJw7
R2CmPcvR/j3TSemB1lWo1qdBXIOFGXAX3u5gKjOcQi0czeCw7K5wkeI3pwRtfnk4
6GZ7ZdG/UGjmTrm8WCSaMIh3bd1FzkGNjWSplxHPXwaxlvuPILpZWAt9pBjy6M3A
2MsMiYgFvewlRb8LUotbYkq4UNr552IR9zJnMrEXs5VFO/2y3V0ib1ESkVuTqgkc
gLpdNm7KuY4Ua/oYj5l7fXYAPbJMSAFZuKW2ixysH9evWxTW/adNAzdSSiWD4WRo
PLlmW+alIsp78NJNB/gelN0H6Nfi/zLGnfv5BpC5HFHHa3X742Ytk0KQP8e8r8bb
owTMWdcPs+t6jtcs39urimw/1+zKUmldY2kqsDhiJTdNkT2sFutgLeToYKlwEKUh
hbSrMozd5ebe/9btdQ/wKgHYn5Owb0UiX8bfMz6dp4GLMa3VZ/Cm2ZEp1QMWmjsF
7ltyvsy0hRkYaesd1G/1KRYzccC5HoaOnKAE1tCA+KYrsjqQHAOp48tKqrMqlfA4
0irkQ4wY2pbPLhnhifG8zxULlcNh6GRHGHtmNB5bEM7Ai1rSZk5HVWDXqK0T6Qe9
Nfpoa0peMU5RaTcQKKm3CAyutwQZXnB/Jn/Ff/xasN7mga4+YsY6eZUM8+1NXABe
UwZD74ZkXR8sBhIh68YrBDbNLw0zHSokdirzRqXKgei+DicRSOTUPp0sbQFalQs/
7z24JXa/Lw8orZXVWcsB9I6tiJ4wwPeYMO8FSnX0S9o93Pt0osLboguUZ7mvLsSn
L4BT++GKC+xvYPYzGFMj53zbdtVJXk2UsGKyjegPycWOslj8CsUKOSfzImbvCBCJ
obVYgxQtx+3nCcOrgXPZxRs7rZmtdjaa5LC+HhOeDj14O6DjYgGEc3OiTvrahuFw
Q0eaKaTdQFJ6wTCHhcxwipL61UCt9LO6rLWbAVP+4jn9exM728p0m00zXoec4w2F
f6ILGE1j9tvEWDrL+iLR92CtCWhIVtqKWM1AQwJT1+3oT/XTXwRnxtTifkFcve25
nwjg2gPCMqbD8J8g9GAnulbIQQZqA+Q6zsZO8f+GMw0TKA0pCF4PeJputlfMFie2
90VmFaSW3gf0DyrnQZmI3hnOV/AcBQl0vOh4uP3LtzNwcDsW1idied/1vKeDHKWj
hYyQYQgG+6wdA2XONwAY0pvidHJLK5XBKYGwmlE2YE4jPN8/xME2wvIN6h5jkt1I
UzxU5ApUiMok/gFHqn8u8FK5Y/Ebj81WgnnWmUdWWQK3XACLEam4aIdtgQc+EqA+
VaQys2QyYKrWXy2CHlKqiAmii2jwJ2NahB6zfAz7f9//mhElAsAawIjnGA6r8OZy
HGpQaYD3nXo66ICZBZT436OFFlcaYBy+qkXg8M5YugMzuXVnAT50SQ2A2eIWLxoJ
+pW58Dr5yf2wfCYkFosfxnYZHAyYFjFgVe04IgCeH8rHqSaIo1RCBK5KPTtiicJJ
rsYj/BI9Jhw3T6k+z/AqvG72iyImxRg6ku4RzPe2OETrBBZzuZqIhRvmTEs2/gwQ
+2CmM52XvfC02IORbvvj+fmcG+zYexkU2P84VSm3m1vwMzKqp1+UlVSfddoXnITw
7H0CgdSZ+6f6BEtd7PNa0XzzK670Zf8xJ01WGKChLu5XAyQt9XnjjvCfDGnn7X3N
s+akKSEnvrD2Z1HVHS8k6XlZOJwrIsa/OjR8P3L7qTOCXPe2oTiGfPnUxFK8dkIy
lKwISEpWl1EpePq1x8t9ClQKgLXMNBpbw0QDLigfOdUlN5c+N7zPnXXLhpUD/0II
bKptgCR0aV6hJlMc1kOz81bs/uIR8ap3UtENaCVD1zCerdWVbSOF5ULXb2O1Y1f+
iJ12RPAAX8Q3oTBS2lzt6fgRF0gZVaniOMQ5Ve/E4nQqfr0KtLMacpQynoTl2lux
txE1Sz/XOH3gcVcnCE8blCgAx6Z2PSDHu+4fpwGBXXpiXhmp4WuPXp1fc+k5dD34
xlcgNtUD1TRJNH5tXzK32FWo1syw+Npakms29Cqy8F08dXJtkoxoGTqqNYlK4q/H
FfqosUDfyOtwiL9/Uc8iLafby8Q5hW8dtPOJQCTEzlTgegw8Z66xaZNdxDoQE6UF
ctNEsZDJeg4lTFdgI+wsXbg5H67oznrE2QupBsnCQZFWI9X5NjW7y/c5R7fttD30
NZ+bQMDFEqHbaUe4Ry5ghk3eYhtt3woTDqo0VJZygbVErwdXtnHZGPFF+oUj4Lqq
OGR3mmcL1pWKrjy9DV3BuNRhC1bvv/4+PyRapGBwCvuvgl4SLtLWbqF6Z8jw589b
4bxyzPqv1fE5lifkeOEJGrsNIpPy0ZMeTZKzBXk5P8JATSBL4VMZtYr+2eIvpgOo
KnTWtgDI38C+SkAgzlqXxxvEsGWnenkrNdICHUxhApM43t0Tq+CMsmduZXTMqrJB
WkgQVULqmOP13RpnmyZxCf41C08Cf/lld9JdZHNubtPvwKbBiaVSo3AHIp3yHU1N
U4VZBicXGy4K4Lee4XQF9EaxLLuSqHZEvHj3RvtAcVWq9bmslPFOhKCFZxiKQn20
D6kGkCQbF6cey1VB2MqTJW6BBQvktDbDGgZ7QRfsqxp5htDk5kKuIWJPf+m8wMWy
PgwPhVWhBdmf4LWNUawcumG4wLfK6AYxJ26eSotqOVaDOnDSAilFG4WKluXAVENI
yCWthXOznkqM3G/VxemTYflJ4Kf/qODcellZB4QQEnrgS/zwU6zdpxqq/hWcfmcX
NP5J6axJhlfE+wlobkgGmnAvDOQezP0TpUGyGcc0E6xpAH2TUbfw2uoA8iBNn4nK
w2by2fVmTGj5QGRa5ffiqF8vCGEVyuinFG1uJnJ+UsiJdgnmUvlqlGZrtmGGWOG/
ZCz7NAEH8PNXmPO5QFJ/+uwxg4a5SCKziarsTnXT33NwAB/n1ouwOYOS2hc44gV4
pG9MLDw7oAQ0wa8dacQza/43eht11U0EtfgvO9YMQrWrbFL2P6CZxefvzKC54Sk1
pAiT6u4h2C3u511Z/y+Gn0qjGpf2BoShU10KE+DGaWkvxgHN1/axuDaCEZ4Ndlsr
oqXAQ6eoNaGdAL1Xc/YdNp2LoLE13bAl4Y1jasLWP96JOweoC5ThY/SBSdOfrs1K
KeL+1ftDbvcdY/sawyaYsAa0NVT4UT4zo1jG8owm1+VNGFAcBiH2dZFngexLOrhw
UlygHugkv40sMWq82yRFfdEfXqUUD4QlWwLSqUH0nMq+lMH5DsoJP8muOrsJ1LzV
/OHidIwRFGZathSk9eoTfR851009D0xjrMMjAEXuKl6rEQxZk1FQPJ8hgAOscaiD
L3v3JByJQjJQhHL74TsXfBohzS1eZt1IhpbypAV3lqtcn0Jr729bIoGlf/c+LVGm
7mB8qZ+twxdwixMaglZKXliWqCvzNZbW+yuzuK9MF0uzsHCGBjS+Xjvrg1nTi6UG
nWk/AqspDB07SkyDQyxHi0NfQhpvrmf6WKniy97T3CCc6PyiqNEzXIXyar2u0XZc
DlXrnhgdpFYROKMIE8KCCBCexvfjtuVyFcQRopY/vPJJhNvg0+meNpS15XN8lpZy
116D/YvM2Y+iWuckG0AHGAOtzh0C3XMR0AUxvjauOw4XuCck2ET6dcxnbVe9iabb
vyHznbWQ4ckcGx64sRgIIg5G5A4yS7Ds6S8jJzDThUqugDXOY6cvwlGlhPBFmGyT
jJJd1CI74R5H8fZx01n2ULmmD2DBkp6xiIeenXkBQqoLdRMSK/R8/oDkfl2NLjia
A1GsrPHoDJpUrJ8Z2OCrM1cKXAY7y0i3q1lwxFxuSGDrGln92oWwKe4aBqOYq+Mf
zFpZ0FpM4qZ6OhhbbCp/O4/9OtvdL8GrUAbdL+9mDiHTsK5P/pgML52T2HQvxGlk
FGCPHxsnAD1HCaRUpiTk7nGVmW8F8Syg5bIhCjnDaT0ZaQIPiqarURIQ2veqUJse
NrgfQjKcpg+ex8XOMFG5IhfxSgeKcSI3/O9+wfw8iuaCE/zPGrQmvosfyG6dLs1Q
gW5aZRg96yF60U9po7p2zHoUgtMl9UduAFraFXo1op2zxowTHQ6XdTBjeDv+yuHz
pwK5k3UcaprNHkaswHoZZh22oYjW5RbNiUp7gTjNgfS5y04D+TUYv4dty6NrCV2j
zFdtf0gO5gzK1QpQC0JG3FF2s8WnyKyfH9XXjfPl6088BRwVnx9gig/BaWxPIKs4
WDAxtPDepLP0qzxddkgGODscueaULkNm+XRAekc6k2kOu6cdDEYf54Rr3XRfgjCK
UUxh4iTiabrT9yxVWpSlmg3tMJxuOGWS+SZNp+YlUPNjl2//4P1+D3tWjXTRGiil
6BgrQ/4QDZbth7/lnQNTsBSuZBRq4TUKdgJQuvVXVOh0b3Cxwd4SBfc7gnxitjAY
EOzuhHJ/qJ2iM5o8rbM7UVkKmqmjty5OqigL4DB14+E2giWTzV7bfI8/Hn1+ixLP
msempjSbmnl2bh1HDW3FMYBViWFhqUgAfSRlrGmo6wwJGzqrf1WDeLmAtUNwHDQb
PD89De4nX9kOtgz2BmEr7xJ2a+p1Pm+FI754VMCZpjXDusB5q+kYAMCKQBtxOKQA
5aG59oLlEqF/YEVXm73KkgDPs4JJyhjyDJBxirH24ZCR/fZQkMkZ1lc/cN9NZA1P
5G4unJJG0zqFnaiW79BseX7F1rw7LzdZymKpAJaW8cZEcJhtyQsFp/FUD9mM3mOr
VEI/Eu8F5bHO9cII6gTxHEUdgvWB3229ALFjmrwsu25rSVRqLHvMSFC8rxMeLAKo
4DW2jOU8/sRm5myGsroRCzPnqzv3zxElH57Dy2x/Ezhw9MC31Y/Aq1xecbJxEzrC
uHMsaHyfb+gPKvvRx4x3OS0QFy4RvfyTmfmNUTO2cX+h+bEuCkIsMbAXDGxcqtvv
cmfk6hnQPIGlbtRJ9szdPLTjelAu+qAvNvZlHv73u3kc3wUtU5+QcwTzzZ3vSfXt
JKXqdF0iHwjYTbAl5G1FTkfG+FYcJZDJLFet23q4mpGF011s2xsVJv5vrsNFUlaH
XYHxSF9Bwsq1us/F1uPooWUHfiB0VLKMNuft3IJ1BlXTFqBlE9i/8D4EA/Tiqp1G
VYD+dsIR+/x8dPF2rv8/fuVor5PxcJILlJyqSDAS3rd07GPZ7l4Vf9Jr0I2Fu91c
SofboGvLy00YHHa3cYmJghhnaF6sGAYZUp8qdbno1v44hv157fRywD3RJ+g3yvVD
mvKKAOt10ZKlNRNkF6NBdslQ6WX2b6bPgaiiZPNQtku1VORfwlUey6G2YYtyzKfh
WYCH/1KXYRJ0ek3hLqlIwX6gJLGWUgBabkOkIHuvgIz3N3YSap1hoo6UtzInPf1+
KqF0hN1C1PBdPv4wyvuivu/E9BgXivobGcHrz4BvyJ9/gtsIEA19yY21jEi3BQ/9
NGt6DTegyNsNRZnEK7BAb+PxzAiTSFjosOUeeQo50V+YwUJBCUuV+SQWowJv7+I/
0ttP/YlvXuMkyUIk4eHWYvCsDFmJYNiP6al4ezMmlVEfki1jOeYd3vNtaby2BVaA
EQYuM6mNaCyON4L171jTcZ6hX50S7cB5VUBpZmcwaUY+vhzVP0jb/H9Rgu3pdF1/
CeR5GYKOGOkkgtItyBBpKHXofC/lcoSMxP+28ySFSJhggCTTvPVYlM5NDCHH/ms3
vhnRtZG1G8iGPPQrLyt5xVP986FOZC7lgpEeiepWel3JxxtFY5yj93QsS87aZLoT
VBTUd9BrO9+cIG6tE8B1K97TtXvBXQRn+bqrzG5vEpwYTysFmB301XjS4QN62UI5
vetAwXyyXPGhUGOzpqWQPzukbwiaFNBvWuIKKlLzGwhSr/QtfVsQeXyPpXENMSsg
mPHnX/wYZGThhQb9vEF/eYAq4wSvmm2tiRrAggHYil+XljmrYgRoTue+xxZ87EZ8
GRUrSE/nUpNl1SOMheoloFqaLY3R4XCm8VACJ/0A/i5FWaqO3SZAYiZ3u3wMs5V0
XiqqvRBOd1WIaUGi/YcuSEYeCGcw02r3+y7XIT4+5vWksrFiNih2a0ahQOQiqQIQ
Va6IkcV4N7C24SImJ9rZqqo3UF6a8DTcQjR4F0Mou/KPOKuGJVusHj+Tn+yJO+PQ
4NeySVN7Z1mIPWE3Lv2Kc0rPV9/jKkC9oH8XCM3wn2HG9TMKTUHkvk9be3cbFJGr
Ak0WlxXohb/dMruvbNXuD8KHHM37TMeEVeGcZjIVaYuLyt9xEYiSmaIp1iYwLVNc
dIj6owEFWeFl2cjdrxntpMmiusu8QeDMqW7B1QdIAfWVUVPZIWsRuohrjRGiCJPk
1YsKQsNrrMu1flz6tfqA6oM4qhAAMrMze4ex96kFtAZ40hbqEe+gN6kIovLtnRlA
QuRKd37W2syZz6gdj5txE/7ghh15VufnnZB95ZtlIphjYnJwG59ZMFuTR7A0XxcA
uXNp/NecrrakxqA9W6g3Y9/kZWMTDvvXR4t87gTItneP4Mf5kHj0tWo1joazi9YB
21LHYiunuXQSvoYB1Mh78vj+5zGzlAz31yxgipb4WoVG0IQLGyqkau2bc/BWtxi8
zIPoHRYBY0h5Nss0NuBny4iqocQGh/lS/CWW1zBrIRsSp9G/XjfWxItKznjxJ74l
xsMqRO/x13Mi3chNMXVtKrn7sYp0RUiJwfPmqJBaYnZB2f+OCBGiFj1iTo+tHY83
sIR0z91GbwpK4RI6VvOGlJge7LIZbq7L+2bZga7KkVRRHXrhDEpSCRwmDAbHi0xF
FXL5RFR2x5/V+Q4lFipZiKpO7bUoLmpgtSfHgQ8ZLo0E21VwqsyGHdVcISQBof9Q
U9h5YHGekrrcukeQLf7AfGzkHhwZm0tDwV7khhhsFOhu8nmYipQob8mYxojrO3gT
cmU64iH+IEH3mmLJjeE8wDAMIgS8HkZ+mPH19bTv2ooKBzfyUx508LJdNJh6tzwU
YDFrdE+ju95aEQvd68dI4+pJ8LSqcsrlImQQqvxsKMo+NC+AzAAQbqwFs1w6VD7a
A7MElLdIWKCvgHgBY2kDmDMdc2cfH4Vz7p6dJMrIQsmVWkuB/fV4ObpMAajyzr2T
GFg2m8teuOFhPIRYrmfg7QWsOzRicjQsRSNmIK5ucBxBFDaQFMetLl2eDWjwXhGW
sniWtNvxjWL9yFNiFQhIoC+zp4I15HgQVLMXYK5fUjAhtOT/ObUA75g6yCOgjl9E
xidoO5SBDFHygKry6nzQEEuZlaPnC4QQ7AYNXfbJrLO8GQ0rIOFxGGWIvucS9bBj
ZdWN4qk7704nEup1u6jkgVH3P8bZdzjYk9DBt30fo8bb3x/o+9avr5UWPfUVlrDw
uaBmCHGN8GrRlhZ2kinImwn/M07k615rkn7l05jwsaudnpGGutHPxhCQZy3hXjP0
JS6NCd0slPu5xn3YOzGNJRBLp3uBchBJKMthC/1w/c7e+950wPlIst9wiuND3W4y
EGipJcjITw4FIB+OKa+P3aMRJaTq9ee6F3smgETcuqgc6VBIkN6EqlPVX5Ll89QD
6kAJUdlKBO+sFpxvr2dbwNY0tonahozUK2QrspFtYsYB/ZtQOvzG1vyEjflIm8ag
aP0G3YNZlOqLo6anxy5N5PgTumk4dJhrdLTvicMTm7pKgv3izROBysziPwLSEqCA
bJzeYpWDwmQ+18UkOzC70STgqZg9T2v4a6qGPzioiZ9pOEerVHJi2TeV6TsKdi9K
CJlRCIrGVdejBPLJTaGpdbsaBdhZ7gaE9BeUVU8jz6KM3GBWqWQwOoUC8aOx1vrT
GbLt2Fn+AN6HnaECfIIYKWN5Gr59+WuZ559cFw38Qr6KTO2nd/ch17bcHcdh4Fv6
0K5d3sBXwZ3jQscBygzfcbjxljyAX5RukpO75zcvUYcUf5wOgZ70o19eg+lbCIOb
7cnsy6JNbKTscpE9YCeiAsanXgHoRWmqC9eQTuryOKLxxTd6rtnpAWs2IMSieFmt
sIo81p4AfTf4me1jkzZBqXK2CnJ2XXARae569qsVv6uYwiIc/bqPVGlsKuofMOnF
H5eZ30KuHGfbz9iwaJs/XuOAkXy/RG/ENit1mZUChhSxkL2W2Xu2zD2muF4BXeYL
+k0XbGycdLoRBrjN6A/uPS+g9cG7B244Q/Ri/1RVpnMm4F4BbjKZCGDvXvHcVv65
sAQV04eo+uTl8+3iW6StajaePtQuxSjWO3o9z2DvBkwdqqcnS3s3UE1ICwDxj9Bd
NVdvVUTcsfF7LbAeVnLx/g0Xt6W5HUK9UY3lSOfZGiJcw6PmDjD2Zf+lSP6IQsmc
ehOCcNhmD5QSKymwEGXlbsHIsiMiQERC7iqzLscb7XnLlvm4U+ArpXXnKwOJirJS
wTY/0FRz0aRAQbPlkzGpcNwhw1VSTZOtsFvMtGB1r6emE3lZIWIb80h4/q9V+dIc
bOwNdJrxBkcLL/lte6Swsx9NiaxK9g7L5sX1hNg9nnK5YU79RCZTbljhxRjeLp+1
vx7AviUg2z0PDs5cVlHEMl8voIIGOHo64zH6JR8qrlCpu5nuT5HWc7Bbmpbc7GO9
iORnwDcVakRM49PbsvBZjh2V7vddc5JP9/wHNdWCtpnUZN4PkvJRqxbbTvVFgBip
9Y8AQvQNsH1EDWBvL+Pm0iFmuJ9cIhWlT4iDFRQ+1XR+TJAbejBq9MzkztVbUA6G
rWGB/sSz8u8qyd6NcUUlTT+Z7wVBXzDIMTi/EZQIDnmTzlrIVqE2lA2ie3UHGfbG
FngYv1ZoGvFnUKKE5Vb9kAsmKVlfa+wQ4K39Gz4OSK3GhOjEWkN2iahGXiang2zP
BU8TdosaZVEwod0XLWJMNRYUALMPZB+N608twGCtKQ6U4olGW9qMPl7sgp7cA84M
NEMxMvTLrOx0RcWFo5rlmzm/foM8HR3t1YxGY5IDhQNujVv0cGuQhjHb1l5huZsj
5KDGDb1W0IWjx6Y8K3IpRIluIQ/3YTWqL9rSXtG7R+ullkdfSH8c06ZRfbdin91R
prgT30tiq8PudZcBsnmZGhNnhPcc7qVxg6SSnnXutwFHf435RAM6eyZUeARyx6gs
c5kicF/yR0YTIetOSlsnkSCd5vchFsHdYQWMm5HbErn3EogFDZXg/ZRKd2+iwUXJ
XUTdoaq6cP1u5At9n7lkPdB5aZidmoUWBqHA6x93yuA0hNCwc80PLP0//mqt3em6
ZK9p7D7gyZljAxuD2DU20g0BLw4PQZsQfPL+zPSktgZVJf1Qau+jbck+4v1dkNOk
vDbEIL2jIDdhaxTiT/JrRXkY+rljsiOaswezXZJfkb5WW243LJA3IEys3qfOjXrl
GCH0IAvkAhCqQs6nZy+G53VhtW3Au8gSbSQmFsYVnd6qVelmaymah+mfiZ8Vvr3d
lRzQZzQnBtw/1GCW33dBsXfRvYoQIY1IYKQlQGh5P5e3BVAHDCVUg+jBvqeePhkC
ADLGN9HwKNt4SeMGIQWsw+VkmOPzHpIsEvsrCQmm1DVSHAvPxDcI2CLq0Zq32eF3
RKYl3DrNPNAlxVUB1ZRzD0E3kT22gJKd3u+xuBP3OfpfgeQLBWqtF6whA2kONpn3
NG6dgP3D3h3ansXOcMNSih2rjM3gnpd5HJepyV4fPBEqqb7hf1052rwT6PPhCf3R
1q6pkft3FgTwRK5ChvsPbYGaa7617v9Sr58Nkf/7QaqPokTKShUB4v1QUhPY0wXE
PKLBoumggLVgIoQon2bS3SgabuDOgXjcT2/7P2VaCpIU64Q07RLzUs+gyEsCIiul
88NjQ+AdhMswRwr9Cp8KTQHEspoSOVPP0LLmEHRr1PbGqM0TUPaMQ5Ai1QkkXAoS
ZNHx8UEsMwMgG2scnyE5sLr1u0EkjZlgud22CI2fi3UEpQjiz1U7iL5Qy/8vFaY+
XpQk7mvhAk07MSml7FeCeZtGr148YawkWY3P8neu28j9GKvdGw2PAWeLy/5N4PSY
DZhuZk0QIAqS/uvZWxofQjnIE7xwnKhXV3drqucBA/6XCbeXii+F58OX10rdnD0M
hYwHwMudfZ7UTo3PbTIYkfLFCf/LIDHL9Oq8fWcDyUDcE5lVC2CqT222qTcIIxPx
0b6ul9ZHIJRCgUIFhH/PYUthbhbrHmwiuos1T9GNOMM4kxy7ZOQdSDok+yrybrYq
TWSQjCv8ueWVB1Uat2oz18YN5oHOnlf9HPilCGsdfYt/6PoKPLomc9I9FuYCbyFo
k1rz94W+Z7smxzHNBZhAOwNn8u84rjhtn8GpqMgY0rcKKdg/SCSQlBYZ9ADiqdiS
EgxJjHISH19hqcEdqfqfN7DjTn+iW6PyqQ0AD9PVPZ3/gYYmXhCNLWJBmJCcs1ar
FGX6TUwdhqhBz7ROeWc96nmhCWjKaTk/jwY15b3PCIu390/WloFCH8fKOVc9jvMa
V5zN33HYIEqDmvGjLljtyvPonk5K/wp+cb/BeXYuBoGUguV/bjgOUVL5TB5aL+K4
2Zoo8ZWyYFEbh8vT3iT6iKFjw0NH9ZazLkTiBy1GO+8CZf7O0sLnizLHC8yTUSV/
Zou9F/xeDddBUR1gcJZSmGc8rU4+Bgmd2kVK76GmpJxqLw0wRH3lXMzyPesarGx7
Wl3bIMrSVMr1kIb2pLnE2KXll8E5vQPCfgmcP0hYl1aCq/EnXX7hrhFH9MCtCubX
mE8WgZ2FeRqCf2TrMzNKuMzZhXWpH0xLMkQ4BvHcNuuycEB0OWpqZ0LDQA3FTX3a
whhk9EDc2UWrXPhSF8FvtBEdHnA3BHCVGtTKqJLp8i3HExWWLW09+0NhiE+LYEWh
REXJu/GeG9dnIh4KdTlq0KQJ9u9fzYRvz1IGWyT3Q6af7Cb8kU3ekN+CKkaPX8Qt
MnPAxvC93UapICLfrIadiYAzph4l1gCgqj6AnaEIkt9LHYfNKxaChEVQGmAABfdq
xOUp+ltpp2O3B8q/WNcfz/6dx14JoV4kKyCH5GyeaJNo9pu1b4qD0id8GWpmCmI+
s7Fsds6nBqJdBT0oU+PONRnMlVjlMV6KD7xs1K6sXDCSMasvrHFPBKg/ZjxkNYfk
g39nncVAEY5s4h9VvGeCCFgAmGFyLQWniSfC3RsFLYcTlxVaNp9tY6MfhBg13Oab
6O1aWBO4VqHq9WcVAc4cSdGhm9RnmAwSzE+SYQWMlIQ5f5Lrn6yiTa1fuVdI/Ey+
Uz2Em72cXAGnmUkfFvWXUUxN7qMHZKaQVNDDETT9S+ShFiqcn+lCpBscC0kHSst8
O3TSIiiR+SgX0BxE68jpWHdDA56DAv/WdGUwJApzroeLKMIdMjdSUNpQ1Z3JePNv
s32HU0wmVpK3PIO0+cVwG9AIrnoyf0qXF6ke7fZClIuBAa6L+/0LBV/aNQDh2h/v
pILUNcp2wYM0iCmKbHxHpYTvJC67AYjsYGsSiRoGIRZX5y33E39VxpSfWaaq54yI
P0j9efjU/A5wrmJbmMpivch1OjqUOS8aWQqSSkRhGsajyToQDA9DnxQgO57S6v37
q+7ucPvOYt1ZJB54lO2kiac6v35SYCxvH3BuYWgV2saMyU/DHfxFatLcp3FERAHH
pmHDDQxDiRiic9hz/tvk5U9rwe7GF1br2/KNJ2qYeUzHZcQ1J3ps64sy+JKb+a8j
FYZHFukdK6HO25KwF5pkW0F4dgTYC06JmSMKRN/awyTBbNXIbwU2xeJoFxPL/xOp
ZCS/pM/q5ErqxuJWO4c/p7DEJ+RWCd3Qe/x3PQsz35hCsiUAH1DPmlqGQaehl8sq
DebAzur6NaMlFHiVPCGkzbA1zyekfJZ1k/ULy6S2BUEPkDM9e+lqHGQXY6sDtqfk
WPioXhVrDaJeP8oKdx+Tc2IShDPHNpWe+FCM+VHGpv9YdI5B3d4g/LTxIDIHQb3X
X7eEIGB6ukq6QBXFu/FnHFSKf9xg9QSHBzs1CVT6pWhEDeIHryMTdODalYi1X2QM
Go8v03tYgy/VthwdjVPvysmt0O5w9QvpJ2ijGKo/m+gj2LCjAzIxVnt3NWJ4XmeI
ol9ZxrMWt3ACtO+9sp3eO1kA2d50NkKzj8o+q19FbcE0Pe1bXzrykSkBAaWshYKb
FFaKXItfiETPQvgtJs0LYE9jle4C/I9CsXF3jsmQJZTwVe9vo9r+c8tYjoRwT7k3
PUW4rxuYDMWOyN3VSz+6FdQpAU4BpsgeyEsKV2qMMYjG36PTVUMFTinxMedGn24m
FUiQBqB1HC+5bFZTf34c2CGUyvuV8ChLhiyUmQGde7q8CUfMunjO3k1IHk9BjjlJ
gvYjmDTnfTAwGfxS699piWik/5foEsKIs/4NWIsXmq1Pzfwvil2y7WH3ZcKxO6dd
2CRwzNtvbl/cC9chrArTtbSLWpbT+851jxLcAxXhiAW8/GsD8i4jInZz1UyBlUVP
NV+9jufx5+ip8TP5Dk0R4JTFcJnviy8BzfbWOoIg5hHI1j5wHizN9prfMRRegjZ0
sHdk9wOoKCgnIvEPygrvtca6eUes3+quKb/pWmOi7ox5rbhYQvLUvRsbBVxY2Kd5
5fg7GLVjv9ZUOlg6CYuWTeIoojtwE8uRhrGqPbI070743yAX2orX14Mniu88qRF4
VRBsgoQ5fupjKq+Pj6CvVZ++kjiLjM8I/XgOeZ5R5opN4ZrULRikxLZaMG9kdV1v
kKUMY1xb+p+WnQqLSP12VnZddB9ef0H73o/6Q6UMuWEhOz9PHNVkwVAAHlIrPAkf
uss8M/MF8bKnDrmvP/yLHl75hv4hIDZu8C4LYA1x4XBrTILe991vT7IDbGoXyLD3
DO8OaTrBURfkGsf0YG4ftU6ZCOlMp/jJD6YesgYHZ+W/bbFcJeSAtGvTGrAbdJ+i
opEnGVsviSpyxuA5vZRot6og88R803IyAyazbK0Pu2/PXNgOQuACij0x3dEgDJUF
T63F7YKj5eJKUz1qNUSoZNIplhGgY04Z3Uux6Cu8KUX4gV/nA+zbQnzBLAAmIOOO
hBajnl1Jiwq4cNR7mrQ5BoRyOvWE+zzaM0Jw8lJ7plq6e6Kdkqf2/FrRmQwXe4Wt
dqXnW/XmhCUb6Z4twY9Gud70T3z+TuNqy0T4QIe8CIhxekgFH0hFjrb/+0WDqIBw
PAgaUA0/SP3bAcr+mbV17/whOqZSpSIWFSVMVQs1308WMFTfRzd5zB0tFOytwfZb
XesRsZLM9Pj/5MGX/gpd/XH6sGRZV5iGq/bAxD5WpmIdC8/TF2XK8nxRmIYBlcym
onFZ5gX+DIPHvLCJSHAmGc1CRy8WaRzwTliJngJnq817oB5ni6WboPdVYjp+RLeC
V34YaUYYP4IsYgAcSlQdnzgZJphPgw1rfj9d5h3tJp4GCVydgKqvV+T/sHORXjZy
nQIC/iwmPWn0kPDbxpyHHFtkkiRGt3gpV1DPdyCQjy4oh5u5VogPopP5AMhou478
Iv26BOKAMJTPFfbK/cBGZAlqUYZPUW5gL0aeCgUhCrjtaw9O+SoNn0BxCh0fP8s8
tTafIhfSfRgqKeS+HbidRD5bYmOAyg8tVgUs/AleBzotkYFJ2amifxZwkWaMJ5hL
VCNAiw4lZ1bXhL0TtxsKabXqVIhcVoUVRo+eg/wp0jnJyUZ0hKJNetnMnnbd9xzL
CCgwmSPBlPYRHSK+vP1WS8SUOBAQYLP+Agx6y1aV0auUzSfwrPEMrhyt/52M1oHd
88PoaFuRBbLHgchOOFObqLROIm69k4hnnrr6i2jctTJID9v5OyRoXm/JDYS3AoV7
ipmyNt6+xQRai9dw2UntZ0C3RzP7fvtwlpLyKqjLP+uIKj6ApUuRjTWHnzw7jlRE
s3vtTu18YH7yYFsXbscc/f92RHJ+vueReAq0tvi+qlp8Fcy6aXKK3phhPiFcdTCr
vURfF7D/YvI1xLsZb+wycP8PZ2QW8kVb1JuyyGu/wuoc1btzumIEOoMdK8K1rhaL
xCDEO0LhYt6W+n92PFA1Ja3wOE1zw/FrZZSk5+xkeY6iMrGGGKCvnLxpcn194OI6
Nb+cBO7zhJg++A20y54vZFEgCtt+kORM8nJsixrKR8OFRPXEzsFHBbvQnzTHSoTo
RUbkEC35HLIdIeo+Dn1cNevLaR8qFWLWJebp5iStBQQaxfGcGSsLgyS2if+Wpsio
F7CvRnITTGUsgjuFEA0WmyfMsUktjuZ1YgW1O8lqBw7eXLIilKW9mw9f9IN/p7Mk
DZnvucU+10/MfsBjVTNziFvoFNzpWnfJbO9GGEa5wZezWBxYIzpaZPCTGCOHBy9S
PzC7jtOvtjW3E6xbFHnxRwG+9AiSYUGhYCxoaOEoiET4lVO5UDwbc6Cthg862NP1
pFm/87H6LYGzm4uEn5LqDuZDTZvJgFqQCfxHuctFRdnmy72ex4WZhmFyBj+nJGwi
oTO348FKaUqBcJl348CChItTc/wgA9JgdPKC8ViP9uOQc91km5DaAXes6/eyKnYf
9eYezcf2vN9n9m4yzZTpJsceferCKcqj1tR6I+QdIY0BK2oSJF5S6KqwPXMEc24p
kKysIpvRLm0CZcSt+ySSXPbQeGI3k7LOpTSN10yiPfhhksPk+qlOo86xwM2Rh0yK
HVFkTMhqAd3UvOtO9m6m5NICh+ri0NTygvmSLZolCfhXODqtTixf14ORmn5B/Ovq
FzjKsyQ3b2fMxwojrMgqAe292QtBUUYN4Wq72loTgsIe2LXs/cvqOZeqMi/KpTBt
xx2nph4WJZhn7PSx6nl6GnnrRN3mjlqSWkUs2w4W0uXc2zT5dcQA6/o6MnTn8tVB
OeZAgUVlAyBvV8dHgFdtLK2pt6aI1Ui1Uo0nzqc1VV4cqtc/AnK02+B4yfvaPusS
32CLww+esCd49uEaweoCZMAuPY4/govPq1DbDnMfFh9wEYX9AnJ5ic6WFsIJa2SZ
eQy0eQj9ptiS+vGiOG3aR6r/Ug4TNiR6+StGUKpE+CGH4ZhulIkxgqtZIy8ZYxxE
2I7G7ZFgUNlTvuF3XBCTrufcyziLlg0nVkK+z3DCkNNWCEtqn8EezsCUEemag1SK
UuOzaUY8t29gUeqY7xGA3rjapvIYlBMbMG4PCa7jOh92Onl8TbDx1BGH6nnEHdxh
DEiKiD7dG2cNGgghAKWoFIF9EIrFqS5XE30ncrPexNiWUniUb+l08ba0h2uOLgj1
B2TdnkOPmxLq5VXhrbG8ZTGotjIapezhmdxJnySueET6NdtQ2W2BzanCQ3ItyCEj
ZOEgZ3KaFTeTfCh5FCOI9y5OLJSA2ud/k7HtvTtedYLNl86dtsxTJWp9CwzdzP4a
vIeqXw7U7HDC9CGtgSXk/KjfPQ4GdOldZwhUe1YW1BLpoD/7O7aFovYJTcsexppk
Gd+UJpR+Q190DEoLu4U155tznod+KVCharwhALwaHuni1vg5Q2aJfMBgYAgq6IBE
ljDXO4jYSW8ukg6AWHP+A1y0rGXr5XXDxten4YdQ6GFlabbqtE/z0nO8EPOoRLy/
vYSfmENUIYRFMBA64Q7OBtvtlnSsMSsDqwX89bRrlDpxqLavRZyEdA4kydBujxld
Cxqsmm6Huh9KHnoCp8Y+FQ4l/56rP5PMKvJzed1+R5s8d0Kb6pIR1S2pA1nSeeY9
aDF33LISC1wMoWS/su0QhULXmHe/APUaGFtpYh2Lho5pmYHsJnMDEx3SvOu+7MKp
Cf7vCQ447idyUKfpJL2ApqXGDYZy8x6DV5hNUNiol8/8eU4OFmxSR5UrTeUlYg/t
Cuad8ABmuk7dDzNYbBH8h3JPw3PG8a/2Xf+Ih4XUgbJjbh27OkoWDUnG1IUpxobs
LhkhNzgTHfrC9qDpxZv350PfDLQGNKWRrRY7OMExgCTwQIe9SD0Ng5/zRcA/8P1j
32M1HMqA2OvwqswkHuuis1mljw2AWVTyzQ7Qke77SBKGDPQkpt4o7oM8B1HJzIyg
iz2Bo6RR1D+XHia+Ggy1qJKxYsywBlWi1wRHUBDAdSUv0yoWjCa9KtfFCwfWn7oc
abTykDBGIMX0DIERu1+S5Ll5OGCbplGoymDWFpk7kyYp5IoyJNsrxAH/So2ATrJj
z6vuTVKBa4Zi1uvN71NyrurTMTkEeSHMIz5IyO+0UTrMKW8hV+Y4xmCGy+aqAbE4
r8hjxehCF7We88cfFKiBGqbAOBrsm55B7hKwNMuBkHoc9gDvbFGviuOtZmjRWVjI
1VqvWTMRvqmowKav8zYoKnVyMrX7mzt7mHC6dGIqUDnyer3rzAi9uYJjzLaEbAB+
j/mEuN+a/X/R4ZZ4/U1A4AfsgxNMf6ncbTwxNDxXjezDTPNUSM6VGdGW3RsUTi3+
JDh3C76S+REkru3GqQfqIfqIJ8wZEtV2Z0fqTYJxd1by+Jjl+/IWkljLLDrcbzJR
3GxtYOfk8xaT62vLF2XR731gsQR0oR34HbcMGEWSkEpLEKIHfbaes23Gz01f0/di
ku743ZwcJ2khIPeSlvEPsqcgFRgfyul2iObJvS6oGXZMsuDM1HDM1jGXcaUBvq4s
yzSjbxUdz5spoI2fWQPe23vPndz+VSPWRPyuNbic7Wu/e5AzoT6Trb4QZtysEibk
TlBXw3PxOI0yBgdtWZq6UAhuuLAedLkcjbxeOG7XQN0qsXxKUNn06Hv9i1dFcHno
3rDCOXq1U9i9vphwBIjJa4qY3Ki7Em8Y1naQF39N4ReaPEklEFQbTTCdZsv0NofD
ZVv6yq1J6kEaIkqJf3JjgaZA7rqUZUmcPsAfllW431E5ua7gqwmJsyZV87ZQXiW1
mVwM6uGKvDr5NG1taVK9kP+da4h6dxXkYXj3gkx7odu7SAL29jCNTGMqcSLQhHqw
asvNrFYtOEtDLU+qgAikelsNbfE0ZRccgR/dwUCkIiupOaVfjnA0oOm6ZZtosKNX
JlnLo6ByM6UzaOvIHjwdkFBpaVi0N/L4hd7ljXk5e14Th0R+wkyA52OLQNWp1BHI
161bBG18ayJKxGNRzfLx+3G1d5sA3lcYcWZKHyE0Tg+pTYElh1lrfh6A9hR5888b
JVG/VnOgZVQy6KfX7qlJSAeBnLJtrjpgTVYkZUq75/Q+u+McqyqQhXFpPAuST9Pe
6/CGVM5fxNZFsR9RmoaVGCNagW5ZWr+UmKndKycdQSGl0Qr/vwTCHvUhN+xce4Yl
vQOBw/8WQK5tKoT6QPoTe/RME3Kv+s5BZ5YC39jdzpVRSXm8N4xBK3w3KeFU+F3R
fPbDj8pt95n8k36NXHeR3MCo6CLWNMtVLLuq4PLBla+HIhF6Q7O1D8rX8CFeBJT7
seFLzqQSVZtpo23VJfQ37Sf9VuGZVmVaaox4X6/iQCl2lvip5dbAjBM/ANRNMsUJ
OO5mIt1ydndz3VFS0yf5DcgbIGSXMznj9wyhpfmXtWaR5poCUsS9E2usirbtN5Ox
ALovgxiVhoiF9rtf/nKRWRf9QzNJJXzlNrfSZ9yf+ez+fLiJNEp2N4gSxGp1fvXF
KnfvV+4hYkgBjLg9rzjA8tRRjniA7S0N6RmIvhxt9EsBV+3qfoVikXXae4ehAkQF
zXxi6BkzZovqTT0Hp3TFF4EnzA1V1mCn+P9sHS9K6r0adEAIZbsbnPmD9xZFlvUd
f151WnWKbfA8K5j+HGQSFn22WeXOKgOueOiR4Q7cGoslJE2ivi2SKjF8ZreG7jje
qC2hMz4MkvE7o1oN3V0ro4WvK8vf+rTj2+GbIxin/Zo0TbRk7f2rtjD5oc5dZmBA
1unP3HHzdoWtMZOUoxZs1sIZmlQ5Uls1QaO9scDbKL1kPUTheFTNrXFsPoUfqn8t
ve3Zy3UpHvv+oJGIhMHL+LeoEeQ3K7tX7mZxUGvSbQ2WIsjMTS2e9/xd4uAAsQtf
68TkMpD2wK8rzVaDLxa6LzTxcoqkix70d6VzcsFQ01/2gdoJOzlS4D0T3P7ImDI4
iAFuoTyA1uHG8TRKyUt1VlmXq+hL+Tm3knb1Ajanmw1mCBfJZ+UQyBTSAdr5c3vF
aXq8lRlSrAz4bkpE9LZ2mCp5bXz2bpElmxyj/0Q7qAsjLpWQQ8G/nPndrwws4AKF
1LKGUa16XwBc3Vwt53HugmM5Sl1c8pl4CBaW9jf9HcwJzypvZQkrteQ0ZzKh4x0n
YT/KgfbwV16QxpkHtlUEsn8Uz6iatkH7IkncOJH1siit/lEtqG5qfGLmbCQdo7xS
T8/TpZqP0ygCfvuL0Jq8Xz86vmtjNN+ajk4UDEUko37roazt5KoySr70K+g0ql9a
ZfdUIRUaBUQQga9owfK8ASoUSScnAEKueAkFcSfG9afTlUUx5hJIkNna7TYTADcu
oPT92IBL7Qa7W07W6yX2rEXyUr9KvnAopf+N+PyZoh6d+w4TymgNaCNUYM8hEdwG
pCy9kU+1tMPh2nEPDgr5S0ilTqEDuj5uD6dR3iZIKynkg32Zf6GN4CUi98nUwqFd
9MGvioDGVZhSefblAwBE/YRKP7d1nS5f7QI+p1WkPZJCnHvGwv75ie00/0qs62Rl
Vvdm8JmkARa4dtzjc27hjsJCeA7n49+CZ0R3W02+YE1H4CJY3b3Sy5A+VDREGs/n
CSpuQX9MdD9de70FprLMzzClqpsPk1UgtpP0silQft6HOwH8xvxIP2Mm6GByDvcW
N9s9T1xoXgwkmYMqyI32XD1f4btXtaJAzMVDQYGs1f/dHaV2AXt/TxbTAF4TST+W
NqHFItrtsoy0Iqnv4cj+jZguDbxjoAxtP/OG1TxHuyMGJnxL+L6FN4Oeq6ETFeDN
EiGghf1xMs9t7NcxG92btmRRfiichJ8yhS5ufRsscIZgY+SyYROda7YE7G+udI7L
QRF+CNCNzCS2BRMUY0UcblTIcCc0DKvSbcDWD/yOdszI8kTu7/utienLIYBCQDzx
xXBND2+kf+RBK0EndLGdg8MiS27v4BH1Te3LiRBtGFiBBH8QMTRZP5eISnHSOkNz
KoD2myy15tB9qtn9AubF5KzKxgEdlQ/L6J8CFNNZ/qi1Ac3U3UkR+zqYRDXEXrcP
ZkvlzGXi+UDq/+gk0dPLMVa9ncf9LSD7ypDSO9niWxsx0BTVVBSjqqHIcbIgWqST
ZiQsTaVoRiU9eTNUcEdpqUxOQTiXeC15AByJPdhYYSQJ4XNG38dUzVMTa0ieI35h
ibneLFw6wiMWH22loQTJhpv+3yxRdYhwVfFMRpGf7FaBY7ZynjG6udyxD+EgynJK
Eo9iPvofPAjs44UBAJCZtQfEZavFw5m55vz9RRnABLQmCuULbUk714CtNtzaqxRO
Q6NsccJC2eN79jr4SWo/qrD/PsgkWggyNvUJ7GB6GNyPBUxFLlbV6o12c6iD32os
VV6cY1onW8ct1Cb0qDbQTykIdcU3c75kEqSbvv6XRHFARCUZttan29jYQajv04Mp
6xxKDnl+LicM5A4YEQLgUfaUDAqK61HeS3dEIezwIiqMbRiDQA+3NeIWcBnFlb4v
eHWqk7cSMLrd0U4ZtvPYl++I11SbSq39IBDQAyMN5KKk/y8y/16gTs62nSIgMPq1
4Lrk5ZCaGU6M8qJPOHGCZ7y9GC5GLGzWfBzEF/dkPa7WUVW7rGNEi8OLz7wbaB64
x6ffZ/q10akvxINFDtMDQlo8bSbsZ1xCILWmFgg1ERq1d8guvYNayoGrTXkW53ob
wbo3fuxz8tFBvGKMTPRDZW8cN1chPuTV/zZAABFR7bkB+h6vRHQEaZzxOLLzqANt
xXk5OutfZJxgmlAwzoMEdDHJEy/JE6EjIa5Y4v7vtsrMyV4FjNfdnkUURbzkzIwx
IWjXWWtTG1L5RBVo3+AjNzVv2A9Ibl1q5bD9ziFYhoiFMu6CNYTeuYUHb4ybRJrL
IjmTRMvaFxHHfE551jdXOBw4PQ25CREuc4bvYS4RULvD9Dx1sOpkVOlCLM//GXZj
n3wKj7uHjbzhCmxaBjsGnjPKnWYPPAn2lOeYOzrctdKOId1V/kI7r5LtLn1LahAN
R7R85zeRy1J2U+uhEvNw0bjk/TR+DD+XNSbhcaWBqzqBJIP4MiPxsiHVFK6HdWh+
ICsJiKQ1O6qTleoepoWCmzf3YornOutu8hhSi9onKc3T8smrZjf9Aw+eZJpmFkDk
SKZQS9hMRUyIqFY70QYy6x/XETVIFM40J76AvmtJnXshJRFxbH+hOOK09EPUOC9j
tiBo3Mg3fMpb2aj14QolU414nZ4BRQU5d+wpGenXSNQIXfTO60h0OaddzKBFBgVr
uz9hFjcE8GaEcPIaxLXT1LxnKx6Ke6iij8IlZ//+3q9Enn2Xxp6IKE+BDWynBCe/
xL1kt3ZMRAHl/N4/T2AA24n8UB/IUP7XRXjiz0RNYMjLwbS75tSMfcWSgdanaBY6
QoJZaCxnImjscF7yqPDhPVkSXBgdkwBVUBNeAzOBVxCJ2uZHSHZ30hvBGAWvJZge
uO1K6yma8W0jZ/jXf+rqAexF7EOZBdiSbyzW2FR/irmunM1XEyA1tmDzYLB92kZo
hfWyhyliLZfz4F/rfmYh6EGAthnPAJOOkJmaEHr/a5sP3A1i3Gqu0brjrmlFwyMe
3ygEPma1tk55x9GRVK+W51XUBU6/ho4I4bhgR3dYjMSgH96ed6bEBAIrMv5RRkb1
XuUEb48tuzW1VdkEjhFl1XLhW29nYJL3KgZcgfzmOQye6L0RSuB0CL4woT/JiFqN
Lgvnk18SnZRJSjOlL2fQV4Diuc07O/EpxmSpfGXK9YGuqZEX60Q+ZjB2aFMg/fTS
9ZTYYPwK/S71tIax+XcSzL3iaw6Bc3KxcFBcTFpmEe++rUEj2HrDVM4UtZxSynlb
+/Jj5TWmusypvLmpo17rxBzLK2ndwifErzq2Z7mtB+k/MrPaP4kI/oZMLVVtukpd
NCwUSu2F5qPkoM6f5sDGIpOnjyjl9iILE9Yl+a4s4kKN95VzzU/1LnUfUpJojPT7
TLI0THg+0HurYQJGyLZorwBrSDqLwPJ+UEtmhF+/YcTyZHvMK91DFO7yGVmmM63m
EnQltfFeUiRY8mxxHPgmtNUEwaPv+0y30XrzyLsEa2awokiV8DQpBi3wQ3hpW/Kk
vffx4Psoy19vu1wXi95PAHjcOipBGAWtkRARufOH/qFM6p+KUmCHyryYB0IP/QP2
/IRTPC6/HXOQh2lhd7jJ0YLN61ZUoaBIMnv3tHgwgo72Z1i/KSzDjYeDOTZOFX12
mL6xw6gpOo+utzzBpV9SUOfyzG95OTba3vu9yykEhl8P4Mk59VnK9iWDYV1g+B/E
Ueds5ZZCwJcKbZo9QgaomvK8yvhd46Sf6tJqlqGQJGn73y4MtY/qs8rRcVih6FAI
ycboPLgIyRJx6XRDrdCokcm8kac2PLvsDy1XfP0pzzkSgeGiH0KHanHN+z/278aP
FqqO4JjDp/9xO0WMsp0NJXdKdGX8zphgle7RYr1V4DWv5hqQtxUJHrBAtDs/TG/g
1/Xqa5gC+3wPqKUthvR6TuctL5LQqyTcDOqERDT8WGEpVVOcpRJwUQbwHXdX9B1c
Y7GlB3g0aRlU0D0u+CJvA16VvOEk1dnldsBFQcfSY6xpJrH4w9ieUCxzrhczYDWP
F7uzCU/SnMpwLcerjiFE4QCSoEKVBlddyCDJ9j75HCwMo6a1OAeVDWnhxRu4Cqxl
TMQXKmm3ITb5XQtel99EMl4laMcCxtLGgcOm5C5hbka47EWx9bG6YL/WNUJFnV10
Zy+kcou6ldHrlASJ+LpgRVnUgUHcenKemfrNfsfmRLWO+NWNENzbo9Blpyqhgnvx
Z7yWYR+W0Eb2s4ZUPrr/XgdWYPXCDQRm4cIx4Oyy0J2twyMUc8VfBtlfnPkbPIDc
l6YPFGqGdcdH+RcPwRZXZVgTz1vXBiWW29J2JNd4QQBpoz3xJGTz2ChhxlduxQ9t
LFuzQXGe3M91q08wXP0EQyDFFs2XOSJGjPXcniMs7qlvUJxmSZkavJqzJ2FJ9VSL
Lo2FM6UnislrMDGb5ZftvUULybBqefsWXFeoN3pKTpZK8YhVffp8VG/DIE8h6KxM
f8ZmoiKNSrPx9/QbTXuLFyDzLxcOaUVjxeDLaUS2Ns+N86QWYGrYRYrNfwSXE+CM
bAoyj9Y0yL3kFk/x9yRheMV8eCAploe3wdN/2IDhunJluI6v8zQiNPa7Twt2Ccaq
P1/Y70JjmyBE7gZenkcp1O6GqHPmBaMt/akwYu77QvzsxMHCGgr1ALyf5DD62jab
uLgq/nDX15qb2YzniveBFNAnzm3MbKe/rrhlpf9KA15g/fvpiKJxi/53F15Hz2NO
g7aMhSwlwpTfz0RlO2ZySH6ZPOSQSBJZ4ZeDJebXITnUxu+h97AtNTPEYLrTTJWx
Izy4fcP1/SG/isAOBjEmAKe11JLae61WMl60G6UUOVGp3lLUWIYcq2gPRYAoiWlp
5uKPO2tEuExFLE1n9aUQsecrMeTscz4o1DBHgHGC298xNGS5s8+g7H+3SFQ4EuKk
vXNJ2zRYOFcG/dT+zPXaWvZqRvIl4CcY7XCyR0pKFWdh+lECQ8YyXyVlisp/WriR
L472Om181CApPQ4rRo1ilHG4KyuqYL+8CvPP/VNQJ3WussZYD08eKiTXQ7c1Kk8T
Zzr0EBYjvHfLoGM+eCyVpNMxnfeeb38wL3CT8+IgivSSc25wJRLaxOq0DfWyRWCH
2XkzLIJBV2qsc5/IBShtZ6MaVMrJRdgCqh9zDHBZaAMpQzZGbUVwX+09ucEQtQmZ
XKuuw1hAIZvyayPSO8bv+zl6uhV8CvrX5RFDdEKLjjav5UwVZaETDuWb51LSZW9X
Hx4caMhOrVNplAkMsBPKxRQDUNgtLRSKipZqbK/5xXAfhc1hgvtsrDcTJyFV0yCO
UgvM/haP7iD4fCYfzYloRKzaD+bhHg7SBWlXSXVtv/l7UA6mCgx8G2F2yxF3T/gZ
YAx+ZuoKmw4aDX2NGxow+9mRrkNeHb4RipU6V1e/QzLLU9K3Xxc0kuWJkuyk/mNV
y7S8SvvF5YtLhepKOqrITArUjzugFqhD/G28osHqH+VX7dgV2BTIZyNWekrzy27e
d4sht47pFDokqG2Jioh8nIZlMRAR4LyiiSI1fm5IORXYfx9dkHKpTpDH9mo5YWFO
KnYettnONrnzH+LVhePGsX9V/gI2CZFyrm/o+4+PV2rlagcM2Ln4S1Kl9/danCgP
9Jakh81d3OFOt5HOyqJWrWge7HZoiuQEex9lTjcumPo4yfxXidQRCBb1Y1t/9LtC
tmvnWWIh5g+4xDVE0sz5hdKQtS5axbg3iBcdVcgunA1kT9js/E2X8qH7I/578gnc
43u6tBVkLqPGsCuz4D2fCiR62Dyn845B/LckqQnlCv3IHKCvNlSlP8HSVfPHzJC9
0525/mhtbx4i7KmZz2FLSZr61s0FltMjjjfj+VFyEWGAqnwkfe+72ZgRcl4T4nTT
PRAk8gswY76nN+dOc/4LJabJeUw3j2RVqMue0wncrQVAwtr/Uy9or4uhWUvA3mfG
zi6Ib4RSadrj5J+URHzY3quHZ5O0whB900w1E9vjiqfrJlTnY7xB+Dtop2muxDfO
KPrvtx5CYGsHDp9bXHtivNzolnNgG7t8wV6TPoWFFoYaPNSQ13gkwy18EmHr1Ob/
L/0WuiFt3fuF/F6cHlDOu8zYtzRCa3CcTPZV02PRAebWhoSF75ppHCCodLjjanvh
H55Z0ddBAxG6n5CUYnX9r90I8BpTOtD+ZCfLTQtUveOP1+PbOQt39WpqllEtzT/9
MNpWgXr14uIbyQJCfqv6Oap/3TacDFT2cR5uC+4CgAoZZHK46+bvRcC1qMIKMnUE
86kECeSYm6UQeXQBYE0GBuIFTHXPHFS2rxnStS61rt7WwcLRAESoQy5GEEj1nmH/
z3exictnl4LdvdKlA84ooqGUfsS4d53BrMjAKASQsRBWXeuX/eBrN1stOJWDrCfi
7ncqh4EKfNJLu1PZKBR0IyU++87heddKizxBkC4Hdf73MeP9oLkDKonUVRi9aygE
/xLbZCLIzqDqx+yHbDe5OvPhS7rQA1NA82KPfDs0d//1S38D7ZgWjxYHeuM0pHWW
t0MpGMYa059yIqoYmEV0DsM6eMQDXY80pugsr7zilrDTlmwk9KlkknCXnuVL4Roa
Iejjtc/hHomWpF+NK2YiEte+yCOm1MxqmDv2G0gunF+0e/CB4OhOwtM5G9s3t0Bd
JfXHNh3S57DXu5h7TGXXumt7cg4kETKvbQLfYC4AQ9PhWqquzOq77qGMaYxfFnGS
fMlKXPeZdHiTN2xSjGIMPN+oZQamb8Bhh29rVAF85cCdGwBKmbVixwgQosXVOeZN
CQXB+DuQTMb0ZWXsssfsQibJ4PsIDhlFNHjWrnvo0x8bHlMM3Piqq3OQ21p4lscK
QhEGANm/NPpIhbc6o3bxt3Oh8v0jLXN7k/QZ0/gEQg+zwrkl3LBbUBr/P1uj6mO+
P5DYUSqurx6lPg7ORt9cL1/dl9sILuRo4hA92VrOozEwh4pVkjnt/6atFFmv4L6e
guQ35Cd7rZlV5nUdruBKIrj+DO4MHxsoPamtdZsLzjJ95G9Ch6uZoCsThGkPpkKt
dFZum8pueIFXioHlsJ+tQ4NMdQDOh+tNKT0DTXk3KX7U+eXLl85USIvkMmIQMG/w
ipbopVUmuD55C58pl96Lp44HZnnfrvLHu27gyK7h9SNXVxho79AGC8TseO+0VOrV
WNoillul9R50oXN1P9MfCpxB/6coRKB7uLdhrziQNNuexjfFrnj+1KiyjzXtVU8N
Ub/UHh52Khy7prCF8ayjqefF93TObqsTUMsp3BkhC7Sgjpif01ff8q6EZL44WUB9
shwKX0MRU00skz1/S6tpgCqbkuM7UkDfGtadC4Bycj3j3bZ9uSPPTv+YdRfAbEhn
5WV1RJ50jiGTnf/Q/GxID5+rZOpoWVErdRbSa/E+7QXMoe3HmcGNxsboBi3YdJF6
DrrRbEcFT6m2kTwVYUQuorW9PES5yIRBoxYtln3jCo4Ae8ETWqjHLl6otd1QSLxq
gFR1xn2RQseGlTQDmsBpmxsT6aBvDJoU6WmBNvJrupoYQg8gUjn+F7At+Nd0Gs7A
QlD55RylK0LJo03/My9743LOsoU42upsPDXLP4ZTSrf18tqL/d1cDAaieKFa+m2Z
Qy3EuSCribuC3wyVXXzcs837I/mGBBi3xGuFArhnFlhy40yIFyO+A3GDBwnmLhL6
xvSSxVfRTxmu0wlhHPu4Mo6Nr7MtJMNgbsRwocwnIzJSfVejc2vSBMZD8YEKlCKA
cZABAAXYP8f+CLocINnqr+udQUmNVuSehuAHxP0t5SQ8jLssO9ucaQ1qqQOVuC1u
EmqZ1CFy5MjSlwjx2zTm9UPrjV8fpNl+BZAOQX5cxQXdLUkYM2RwPDpe7LpqHheu
i6Mmh/KTbdh2R+LDLI7JLXupVlen0a/ITkOv+ASUBNJhZBmnQPeJbSdWhpuZLPns
UoTXxoRUWYqffe18LwalZeCF48bl2chcG/HElpZGiXx3jlwLvl+BsjbF8uTpBCK5
8GVx7oTNsaelzTEBlpte5xw1hpZ8jZjGRVglR+FwawMuCWlz5bI+4W9HyQSL4MeC
06FSf1l0Op+AGZuSgx/C2Qn8Q/OKsoikYzIkRKJ4MeIwwDRv0NnmQsI8AjSw3BIH
a5t6MV7Ot6zAXUfmOnsfqBGS9GmhoV97VtlzAWvfNa1V/Tlor64Wed6O8wiORV9S
i2vKt7pMbUXeHdIytcLs8mwYYQLRrFZXoKiD+hjqPXz938CyZr1kpKuxZx1cI8eq
TXuVf1jN2gnwTT97QvVrRZlyrGBUvw7a6rYhdotTJOZpSmxDgf+K7t+/K0SZjb0e
BZhIVftmhSB5d7sfN+Flamjs2aOrhwkyLHn8kDyhjW3WhRvEHsdwigKXl2NdCAIg
AtDyFEN3lk60gsidjgnJ35vckZUKLQ3qLWLVPAO1CoJJiObqARU5/V70NhuDgULL
thdwOU+IeAhElc/uRrwxxR4Djh74KXZMES2a5eQH+aPWUMT8LZy1lyvXVVGLy/AA
+ZEuoDlvkG8ngSEhljYue4I4l46+JdiE/IFmw2it4tVij79fjgazOZbf5gOfnmwF
xqhguE+lTzHV/hwLeVrNRhgCD2Ub1r4Jyx4u0tGAX83WDTHNbJG7usgHJB0D/UHy
PBklQQHC3DQhQnfO5n0Eh+C8WuD7CRdgPBbPdfyPjvZH0jsGjZe5P0882gA6sdn3
8fypuWNhc8or61JwE/LIF630OWnRFkNj1rc1dkfBWMztPgBU6FmwKhklds1Atzjr
PtZ9CYhPuoVhEadPRu9hQTq8OfkmL18oC5bTSWZ2pPEPdG6uQVeJz9Pzg4Oe8m+s
Z+B6nHyfdlGp74eYBTYwdr2fcx0zWjNDY0FCachNxfZ/p3iuzOJIUW75dnqeSTHH
8JvZqBqQB3RIsOHo+yW5MsVil7Wt13Hqe9LvfGGsiQmuJYhBoiCEQMIiIhpm3ZP3
dFuAFzmuQIIzCT31qJw5LNFucVNKQcGMU2RBcJszYz/D78JSHFAJ4TwWX0kygZR0
UVeHpqDJ8xAUFZYyv50opDEwpFkE9bRU29WzcJNhwRYvzRQaK+GFNpbsKi+DrGAs
L8BiBMVERHH9vN8H5CboJAqaIMHNp5VSsxauSDmpBFAW+jP7SLCKyfhC3qttT01J
NI+iB/sxc60XSgPkHjPXVYSCQ9TQoRNJDVadQ2xpRf2p0aS+4gDynB8oC0BxkitZ
xLeoNSsxnDuvJQh5Dp2i7Nd+74Nt1qQw29Sw4Ch8WaQL/RnnobPlaMzZfM3HIDLD
zrXjjrsP7LbS1y3iqx93I0ur221sDoXMZedkrvSxaYF7HC/CxuSxmcjN9wPa3YTK
yHygxL9esgEJVMuT1uOHSE0yK3TSEF/pKqpff4oJCZHkIJkVgI+mUHn68TaosnUm
u3jHMfbyBDyPJB98whVj6gAq/78RxtnWqNRfUnNXBjen3kE0vVWiPi2qWvxqRLUo
vEkZiyGc6I18YM+2FGlhLOEZV+w7DzESFCQ40CiZR4J9EFzH4eHOR2yhHbkm4Emv
ThIABb9vpWJbILQh34xadl109lHUvbRgcvmB+l6uHyCNz3825OmPr+YqiAZdE066
RKPKs5OSqvcst7M+SAWP9lmqxWRET+/GYTGFKrgaE7AQaZpyaIPOIS2bibZl17vP
C1EdDdWGRgMMl5/oUdYb3rYDk2V1tZaAMwBTDO9A7ZgpFCPQClXun9H9/5/jV4bN
OSY0fRT+qATZeDDSoIm8w3FqJvOaQB6xyxHq6wNj+4aHhmk9Fjjv54juGNOpnrV9
k2UT5bEZb7wPrFont++OB0hCF+GRoVcjEgEHoIXniF+9nJLkR0z9RaBTiGqbF1n5
RRdcohknfbGAD1s5qh+fwYrBUoR7hVOJzerw7tUcWRaAt219Jm1BHjEPVRtcwjnz
1fAV52B2hdkgEmOSYB1uGDeQuEd4/tzvty8OGWtx1FYUlikHPDxLI4uIcyD6H0b4
jYwY1an2C2LpcwdV2MI4PnWRXBaRQVOFx4j8adU/KIOYPhg1k9D+4Zrgk/0Fyodh
jgWjhnI+o+mfRU6slcrG8gKyzpj2IPukwgF+P9rwGZFVnX56DrjgHuqqKF9DE3ef
Wn2cRkf8jzPUWM/TytO6YHhZmSQopCv3BkbOHj7LpAg76uNjIZDpXwGZEEw23Kwp
1Ge031elO5EElsg9ONMw+K7doDAfjZhdalWvRzcKZkF32+2aytBTPZqFWv4dtUZF
5rre1tSMxoOw6A7zVbqV3HqN6oQ3wJ7FmXZ4rnbmZX+EdFMyYuyBIw/CaEMsU89x
sqUeiWRmo8V0pVT85VjfjajBTodqvw37U+Dmb+BxXXy6F5f3uVoNr51u6C865mUT
OssuLtlBr0CBzhqdNIk7NotzET7zfldL+7ocHSnvMgRbwRuXK/s6HxyY0DrmJjYA
X90qTBQFwV40fcmoza+5qmv9EiCwy/+LNcZH7Mn3CChNq77jnLtDPFfIXtNwcXnR
98Fu+g5e/ttPe4mvfSzVRVy9W3EILItSR5IQpRu/OdiUxWp0Jh6cHz4xFpJgMbrI
/rLIVJSskiKojYFLuyjsPgDkjcbDP4qsaClMmWuRULLJlgrLJ3vPdo0WnJxziRVJ
nncULyAc0oT6glrD2J/4jlpWWMYByIVWlxkM3Iq1J3hrSlmeILRozKhiAMRvkA8Z
BnBp3UTeATOAnUcZcwkRHsy8+NkTZcEmNQsTTawjqUr5KLxNdqwliC+DzzEQ2Ryq
I25fx7BeQwvxqzkT8PC0+EbqyOyLr4toT/41RZJ+i6U1NHWxaCSIP5gJsAgHQ+QN
52WZyQYectZilJkdFnZk57jm8kvAt9qd8TkKodO58kY0VQrk/Nrmmg6GpbzimJ9x
r747Rh/PXgox8HnR9ep/EtHjiztlZ4SbB6cwuB1SHjqYmUY89P60ZONFLiIIjXk7
ySbfGOBAoKSIYPQVCgMdca39F5tDm+GWHkqEKj5/XqVq6qwLXKvJUV5stKbwx6BF
1jKEP9runZnF5dkEgo5h4/kJFPt2HehjSoYzQPNBK3wFyc4lEvWgPqAkOO0cZUny
85/JVrlfCf7kN/g9QehGNOCZWiEbns/v3gBZSwOYtZWwJkmKZAWzdXuXz+tiXJ/g
87qBYRxY6Z8PmVdGkNBMfKRS1WqcfVUI1105k+SRkTI+eP7tMW4fdvOF5x4Vafia
63XVqT+w9kyPxQpAsW/3A8DBKGbJzlPF01X0jmYe98e7dJ3mpkSg7Pe6qMA0uWwS
sN5ihOwwP/dAYLtatlztSo+tvbDmJ7gNdiGb52vX6e5O5onWgnfiemxfwQorHWya
tmchH7Hz8krjiglOKzGvqugYFBO14yqjK8b7DMsrNVcYI4XeR/UzkdCfoz8QSEjJ
DqkMtyLpmjy3TMDe/ricTWU58WnDBXszvcn3hjsTTsW28+H2GD+ysQKR41xu6x9G
pqiC3SrN/TJmh8Pv8Nfttue9etltpX6/vnbyqMYszyuMtMOsiGtadpc+r6DkD3XD
0nm+u6wKHkgTSzw/bhx6K8eknVZHWunzycgIulr1foBsXtWEu66ZC+EDQrKYtPTD
c7f+GZKnx75yNV1w8U8Hd2lzuOPHGhkeff1dyNeygl4exZYQOKNVbWn8veYXDhCH
n0RxG1yg33JVqUrsOjA/iumDosPmnUne0jcr0DuVP1EPZtIXv/rrSnMWYKc8E48W
wVQNF/ovH0Boc6Gi29fLbiqhe0TWKh2ZN8SHzM7CpkwGxmxiX92Gc+zhILO4q3i3
lTUDfCtIRlKu7lB9ai9hRpA6+yGvZmaVfnKpW6a7sjRE/6auqGZWcNW+K6R+zoPW
Z225PEf3oCIQkIYAYNntk/94YpGUzooueD5CgNj8JjFQpvw7ijU5V+68IC8/v+f+
TQ+gsKXdzd5nE+oZYnGaIFrxVbSR5qCEqH4ftTM/71l8W3HCOZMQnIUiDmgvWQDb
2Rm5HBUjzJecVDrh47w2n4IJSYqgHKJqSu+OObZg/GDGziVG7vBumijFrOiMdden
C21ivJ744cYbG2h7foAk464+uc1WMYXrHLrd95iKEBPH0lgt0UHbXq7KLmANPjx/
xLLaNkTUnlSWXa81n/OonPpZaDXM23aoaCutZtdbu2MTSUu6b7o5qC+VX/DQ9EcL
qYlfcSmezp7I3d+lozOGoJX6EWxPFXVVnDg5hxn08xphlIXoTxrshdjbkBnqX01R
5ziBuFuQpmMxwYhU+Km0LsXiCg2X9zIeDxM0PTqx8K5LbQgZ1WaloFM+mvx49QL8
Ywm+6kLGBccGceyZ/8ZsFwuR7XL3h8llSXEk3knpyI988i7FQolAEsL05MlIBCYB
3W9+HfhJxoJ21rQ5K8cfcaeM505sQ0yp6ASc+QG0iTgEC2/ag6iJLFWTWR+G1xZ6
tcWWkWum7ZXputDvSHt0P4ROxyCOFtjHBbjK7vql0mIX0XMLx13sg4Y2Xl7gFbYI
pgV7bDSHd+Ra0qUWu9bMDXAtKhX/FKbK5iyKScLxV5sU4q1oI4UNaC4WyL10g8i3
1hYcX1QbDoOFJGOUEaf4tRGr8IGck7sVRR/i9PSLRs0j0CFW4seVS/ucvlwTMCW2
SaRHJhiJHVEqGJNgtviewB6sGpMcwyq6dcTqyOwhDwnxQoUIbEQDE1suyWBORrFk
TbqAbnHa8BlDoQeJaUqOYmHcAIWw+N4QD+wX/5+zUJoUqcneaCTftnsAvwDCxF1T
6+fKFKqjO9X3xYH5TO9viwyTFtcLHwqo8rXLhi/2ChMr6eGpHQU9czTGb0ggv5C6
3ZRFeHhCIApRsGEwY/sMnPGrmwSoIkBSuX9+Unuiz6Ln/SQf/edzP4T/SU/yxbnU
ZMev5yfVaK1J8vO9HTjqjXuUT4y0DU7y1d9WVlIx+LT3SD8L35CGIFfAo6uq996T
6nnAf2huOtbvQqvD5eQypo0LDlGPPhpvaS5dRG6c3be2uBIIdUxLjBrmn7WgAu9l
cPb4GAjG76erbGaIt7SZnfvf881KWV0lAnKWWLclZzgRLaCsr4H3R4vIaCGAgv4W
KwxU7qd1eCw5yiTY8JGpjUTnlkl2i21RvyzIb9IpJGIByhRMz3EiZFpZAk9Vw5ya
QS/3/HkBDLkA90eGrmzYayBmlD2O0RUW1En9GuSUEmgQbBkcshkl/WGCmuk5Hbj7
W/OJyIeUJaT+KMAlI0HJDKKgbUPsrzeKY6qeSURDpRlypurEsKCukLep6Sbjtukd
VRen19W89BHT8+O5pib+B+Eza39Dq0P+X/Ni65w3fdvHQElc2uwvvriiJXRIaDeq
3h00UPRKUr1fbjuHzMlHjrbk4PD2YGHlySP8X9pXO4iO9o/XHbXji05mg/L7DUIh
YbABG9Gz98MBKZPfIZSpBwouOGiZmJGAsfdWydkLPu/JN8f13+utKmSt3g6ciddX
BXg7ruEOCcqF+7oaEQbkQfUc7ljVV4GUJJT1kz5iwk+RuWI5o6Dmpcl+jyqizDBo
PgKmEIaePKxrnxkB47JUDDYio9LRQKbWWYSKwy2WJXm/vcuDUaZugeKL/hpfgp7u
BCfUu04Oi7DBIPP2jtT4NsnT9YQXEKJtPCXKHtrlugAu6hkGlmk58xj0caNp2z92
XwEkAv9+hWanbRi25sHd1Tze+6AXJYrwKFbJ8P+aZgBumWfl+5jGp5hih3gIyrzn
Ubk+gNsMCPQu0WqgUMnmLEXNyL8EOdgXYPVlh3+1SFq1wj71kRVjGePIAiQb2+RX
JCeWsCwxnAPwQ20hAIb8cKLc87h8dmLuOLfQcy24ZLRDbFokKVFo3ZK2h0MeOzWF
N+J5eVr3cYI8WG0ew/0lE3WgkzWDLKkFF6h0ScvU+U4/94MzHDrF7vzo95jyNMNQ
MSh4l2rSrKS+ThckXEVinfHHhHY4E1lc7pVLPLRmBaw5xp5XjvhPSeCZ2wA7aaDg
mcPQR8IxSaI5pPMEolTIwomWfRt/VZu9eRv72jUmN1ItRoqTVmuZ0QOvO4ipGqfY
aFCsTAVNBWXpB6O+GdHJjuhzmJ8I7/1fZvofH9D7aoHSiypS8FE/hgCDjMokv+Gn
3PkdX6xQz3vos1F5NQk0em2DT8QxzJ1V9mRpB27EcduIvKqhfJjqyLoasw4m2N5i
AeRblckLwqCOW8sMyCfQl9fufrbhl1m1sF2WczwfuEFmot2ArIfjNUJQV1M04BLq
qwcei+3mqHMDC959qXE4CGX4xsL+wTiXzsa0zV07UW7OeSICoLfdqmCufTz5by5A
/w8KaLaqp1FUT0fSXn/9hJUdxVUgOmFNhNH4dUObfn0jCbAO0c+gvzKRrG2qYuxx
/3JZGdbNlqL8vys+A/xcXz7NXiLAWkK4J28RS38VbMmVqAJGUNABZ3M+1pTb4vyK
F1oaVzemIdWVr+AU33EsGNQE9++J38AOQyUgYEtT/AL6VoHWskMUhOJjF2zfOQfF
XWMVuLHM/EnpAkyrrEfSu4K+z52Jn4kmo95zVz2lphOcoJZ4n1YD+GVp0DxHkImy
BydKTAIfKCsQTkbcLLvECpq6racKQ9OtzqJG6/oZUbvQYOtY9OsrhEavlk0x7/Ez
qLIOtoTcdad98wR05EixG3Dlryn9d6aQtqZdbgerwbfFMzlCuynUK54/bSSYgrzb
1SoeMjYV9oJ62ICafoYsfMkv03Erzta0CjsYGNZryAM15X3xv+iRXSPGsPH86SK7
oEWD3yrLHFHLfOLP8OeBDbk/YjBupEDCcZLzCTITAUQ7RzXw0oTGCu8cIAs0+D+j
7g3s00uCYtwMb7kkQp58+qBBYZqqbBDWx/hfutgxr5dmT/Qgu1zSzfG8T/Ae/0kP
/YcO3RvgTX/WPMSpq/y3HXDKnR9fmacEzFtOqq9pF7fXnJnJMzaqhmAriC3sKr2L
C4PML5VVAKxt7r7gp4XbKCVLv+LnUWsDKg5bd1BtXMWV1Qcdz9lwszHS5ZXXfZhs
a0n7j1JqI/B7vTk+6/tKRt9EbXytJ50dISuXbvQG1tajQhbRr/k/VxkUpcCEHDL3
ndnvl/mnci5GyHXLjbpQ8LytJkeOU4GE9VSDhiAFp4bqbM0ww4aoUb2Bx40riDqN
/GtNLYZjP46vk8ezEdZ+TNcPVKcjnkCixUEFVnojnQVzo1nrhQO+qKtIuwkuI74F
cTzNt7n+HNtzFtzryTeZAYtU5f/BJBiwWPDa3cskEeryVH2HFPIhR2NBdwXLVIqG
vzGYyxCZ89hb9LD6QoHDxZHccsw87cUa0oyJbY4rYIbt8WwW+frsw/JLwrSoh0Vh
lzh28wFdelKDtbScNuJq5VMFC+Y38uRm3vlJgpXhWx2IZT29twXpHSs1Qb0vBVcX
I2ttcKQg7dAY1O+k3qj8wT2Cedt283bJo2QqUa4r5Cua9HDCftU4777tm3hyAls1
8D4FlCV91onb/JfbcmflrmfpwUKTWHAkFJ1OdH/SE2HqMrL1oDerDxmp/v1eMeyN
qRXxEFtXFjyo9+Hbs4SxmBNCmLUPhrjJMpUydr6zU/NlDCvnlxBchfLoNxgod//I
djZSAO+RVWbhTpC9jkLETAXpMAy0LVGtqRlOcjEjGA3643W8L7RolixIZVl8Aspe
0171dFr+yI3/1BVy1FuXz/TMxh4Gv2B/o0wW9JZRThmjKOwDiO0u1V6ypaQ8Yqd7
ssg3xQkm1lOwzzF7CJ93DJRQUD7BTgfz3R5gDS/P8AGM+feFsq+7xkNT6oD9Mibg
ngW/qG9JzatlnNQlejW7qzLNit0aWCgQ+OJx8YVtagQ+L0gNAl84KHeoOX/S7Oe5
z1O0cyhdhIRa4SVyjxG9wyKVM45KQH+CsIiSAeyc8kAp6yV+g24l/ZPWxbxoH1Dc
VOrgt0TE/IunCbyVf06wpovrohfMQ49JYDjGW8dHkpbMbUtFVNiUZfrTKs0m3yVa
xNEwJqCSwDFF0DrZzZCobxtC0SkDk14akDFQvkdXLNkjfvmSMZQjBezYkpmRL8O4
dkj7FpuP6U/oQ3KDvFi7RtoxTQ/9vInKDJm4SoTCVvyUdHJt11qhHVax7lIKEpKu
9KL8sC38iJYuDy11kNRvNSzNOWSe3ABJVnUxZFR4sAPNwjyYmAUs0NjtonXaoJzm
1CS14cTW0ZfHUI+/G+Bf2Br7Z9+E9KNoKbj9SPto8r3hl3JE/hRaV438iBttWLib
GmrC0wPqtqZmbMQsLwbEk82HF5vzhO4UqFN+pVnQj+VQWUYQ2iDZU4BZb1+qYq6J
RKw1O7cjQRnAS6JtFmcYscL+/uI1vYL7EJfPhADiLSOAANtvjbFVrDMt0oJoYEA8
S1hmtKlXPJECz1N4rV0Uprqppq1ghAikmTKfkKG+ALTu9CTj4mWIGqm9AgFjP+CU
kIfhvx41eNsjMlD4wQurlCiQFm9f/1bqQgk8JIvy86CgtnOKlV8kyI3dlPtlTrZN
RFmGeDevj6ISKNXFuVPB7xy2LD/UvW+2Q56Gioj0/s1gRJPyWgMlsZMih9W36KrK
JfnNKWVwW4HIhlCY+ieeTzXScx4YFbZb8o64TWSEhj0=
`protect END_PROTECTED
