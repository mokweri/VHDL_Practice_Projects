`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PXTexYFAcIPUtQPlNoIkTGUtDMPJPiw5B9LElFwGDyduYHDiADLsYmv0kYWQe95T
adniyChGHC2v/VU8jovN3QwUC1kh3NENPRdwCYZW5kZrKOkU8rrYoHY9kUHtYa2x
+6pmh0vwySaOPM+dzg+E+G+NGGejDOu8UlDkEOM7vQC5wvzSwMV1/0niRtsgnirr
JxCiXnxEv8k26NmAwa9A7X/s0iVkSRXxO9fwpNkFdIh1UOyk47er+Xc6ZwvhsG8y
Jv/Jf8XdjctmeFWMDHw28eVE69VL8kRa4A/n8XWCTsCIFHH9/QeH+UwkRztyDTD6
yRLljhjWfu3PEXZdH0QqDSBFU4s4FzW1wwBNxrhPVlCshr4p6Fo9JOIjBDJFyjn6
y7sAFzdzl8HuSsN0Mkq2J8sz1FC2Doi/itJX2c1uRM8wpPZBFF6GGUq+Sh29qRQI
DzCkeuO/sWUks+u2CpZ8+5NaWxjn4qXaEHAj2BikBsNdW1sIpcP0dX5KR//0QRGD
TCrUXXTpzmOEuE8jEzm3I7qoYbiBOZOyK8CfxAYalyXJS2mz9q/PmpzV3bVbhftQ
o+/899UcTPBrTF6GH/II37kj/leXaa/5tOY3DBi8HFy5OTR79dC2qGeVHsmptynq
EmhzbuSeweq6oIdBxTQetpfToatQTyIOBsDmexQreJBK9jN3+l93xAOgF+ix+VxL
BKhECCuCHXQvrqeJaUMzTFwa98JvjJvUN/TAXJM9GTcQPrSbdM0lirdTs+WJyQfK
4EEaR6FirwwdRVuSVbejJvPwpk3cyuab15FRNGs8FT0s+h/XS9DRCNWP0lXunHus
S8MJOz0841gIuO4c1qnx/n6LYJHhrrqSDbESmb0Qv6gIXPC8t8f5lklars5BEWxk
AvLq8xUqBE0pc2felwz+IWMjzoyGPvlHrzJZcFzL9snVBpWTiwjZTYexy+0Ua2qy
e5ImOHcvhM5QgMd8pfkXBB7E2Exox1/L+jLXYABAjMBnZiiXkaBt6lyZtyNJkS1a
M9P4e0lJSukN+5MPCOELOubUVlzahcmoplazUa9sFLjKftkMlyHvgxM2WC75c0TG
qtkti3ljSTi18yX9i3Z8eIf8XTgrX0336fQF5FjljcTeIv4EPg+9T/ZUE9v3qYJ8
Aqmv9GCcO0Jlcs/9xiJhFAATUSmYOVIdsm0p6C0i0ZlGq/ZIasNzkI+XsaVOHRWs
IEdsZBTSDyMzLAgArp7sdOBPlNs/w+QEa0AvFwavXwGw7yrm8Iu7NeHFCs094Y7C
2flFm934hUv7tZLuwSmGCNjobIwum/a0alKip2q1RruQn7aZ/Gr+cAS/B9wLm9T6
rITPrdTLG8Z3DpH12wovv1dqnbAtQFtwaGzzy0/rLlxOauxMB4usRkRGMHghabtB
VoYdAcdLi119ZpOmCVM62mRpB5EAfZ8MgrlcgZdmIn8ivqogWXd5TZ1t2D61C7lS
/bzowJIrtj1/iqhVrrb4voqM6nbd7J+FRcU7hrMv90aiZapuln8KyVW7vSE+Konv
YFwj9lr1zb7Ag1gAdQNJ1mPZ+M1ylymzq6nQjLSDsIc9n1DjJ+sqdZoS0vlQbjMq
Cz7BkSK+QIKv9gyaKa/th0jLHNTJ6OQcYUvFYbiErOAcjtaO/hqOx/ol5hJDsfoe
jMH6HSQOBaINXWk4Is5rhVcYzTFajGSlg+DFHZE7YUSAwn8cvY5tjHu5wHCqESvc
m841mgbWLe9YYA5L1/EcRltfaThk3px/NGt4EGWkuIORB4emsQRts2kmYcFGd0nV
c4S8jy5qKIsXKqZ7BOTt/JmVAbMZGu+a0ijMI7F7T7gvWCTOhTLugFLy3Zw8hKue
rJWZXWeSYgmE1yNkqKZQsBgjFMCDCQ8ws6EDeGogsCQ6ePy2NzUEoOkKq1eOedne
/EwoZVBcMC6iRVzK8pCjLZMhWqjTxvCQfns73A+g648SpWS1+p8G6bbxvLYS2GgN
ps91UM1u+aKnqNrOdmoA0Ij4bUjQdTcw4hJvhNEkC6Qu8nAGRY2VKKMlqTwUOcPB
fwd6nJLBY7jypTHbyiZTboZz7p/3VC184tlFa7Z/gqvPpvpGBgIikkA6ifnS3KdZ
ky7+hFK/2azajk/wu3wGEfYdbvyE86kWdOjnjL1Mv3SxBoaR6WOuF5iLkrX2CBj2
sDgOifBDCgw2e/v99O1+xCPhU1KqAh6THRpQeFlGk2FSmzB6oJv+j8+j8fngluMo
O3RE92XNvBdoJEnELJkYX2yeemlRuLEhd/x1lQDpmJxJOVZj/5c9nTGhYMWxQqeO
rn6hr2eGpD9GMIdpoQH6fyv2pKqKEWGEHci7hO1JAuQY+Sd53BneJ7i1V9Fk19P3
KQAZWuNVzTYNJfB/GoaKD5tPij8apWLq1ThiCsZf2A8WXc7G++Bm/zlbDBsQVQoH
czevzbcALBdaYcLGv1yaiPBNg0RWTNIQb+ujSNuYf9q09kI+IgI+uKsfaYHrWDtE
fy9Gp47GljPVBzXrzM6K++XAqJZnriGSyvYS1nXeY19YMbiMChcjOgXaYgT8qyRM
Fb6Jl/RK1WxUV6ZEObX8PVj8ED9fGNpfTGnfm4f0jOaDtCXLJav0KowEuIbaC+Du
ltp0tFyMW7HnKaTEMycquo1h3Ieb65Qtm01oyxulTJEG2xLu0P0lFzuMGEwR96C1
rePvJ26yH/dFNGxAMGB6euVjY3WO4VQrrHCAtFv6l/Jaku24SQCxDRru+O60ySFq
x7Djjc/PlWsUuJP1vVcZKIGxGMZFABp+bnZ9J2sgbdLsxR2dsgsELI8jcXqIzpX2
9OQrbc8nlK1qjdTept+vP8yaWKaEt9vIFpmKdRPkJyv+Hjvn34uhBLR4COrwY/ok
tAERwypcoNH5j1PEnbq/K+NqVs+JuggVTh2KwuMqLy1tMhboqQ3bacI50tUWFXd3
Db1OkK84dtoAjxP63uKBuLlRccvkB4T+VQQCIoVf+cj//XO8QWJ8oR+MqIpZ0pYx
IZeeUEOqjW369PWQDO22B2uePI6V3fKEFk8j8sz2SPcGsvC4RWpc5R8y0XSNqK/t
70HkImb34A6Vayb1AqiDLkmzCbvcOEO637QRPDnrZqtHT+tvCVaJKADjk6AZnkA1
c0c3f3bQVY7TlC+X2AyDaKY5fnrIBrDjKM4nOH4gdxqd39b9SznVBy1tVYbzoI2l
4cHvf0WYuRqLxwub+Z7tsPLvL4ptQAMx7vX8RxwjcZbGLLG2j4c1gdyS/TvRbY2V
7HUeOu42G4VBtClqGjhlOqzpQBsiIFsMt++T+wbTVoe+TfaAyJVcIoBVAXDzdHbs
py6+eJkfP0Co5buIccSuBBFLeoDg/7kWmEaVrKJAwVLx7vCJaTqmWcheAjZ3PsyV
Fb6jwW8Ziz9eQyuC4sUG2ybWPJx/AKImk4tVFORIesfUbrvEJhEIYF/fDQcfGQnG
HkLrkVqz8YGHdJVugkHGxoV+IuhPi0fpXFKUWrTxBsZQyR2dN671jYvE/KqRgEyo
/4ljkMlkMVTtfZ5G9vONlPTSak0LkFUv2Ynn6/S2TXjwIS56R/qNMjMScRnAN+sR
9A2pFiFJtcNhM3M2aX4PZVb50O6mf/c1ThyBEKXIEGtXgagMZv/xCJ9aBGHLjSOY
isSNGWUThLt4g2v/V0nutlYrD8ArOR5VRWAx7NRWlC6bLyK+JriSJxNxUT1u1LhE
lVfT4Nc9EOMgn4LBp8ynI4lLR9oe9AVAXlos0gXkmSwK4nokh281becmtZlD4Hy2
RG9fok9wgq0an3DxV93ZTEY332WNviA1TdFrfRsmnv898cwHX9xghoYnVBe5DGJW
M+Bu5Q4AExzVVK7Qc1dRS+8c0+aDp/LBpe3irz12wUbidcGYT12afTC2JTuSWEI3
U6z3nq4Ws4Pkiw8Kjo7NW/13QAWB1gdx/WvyW6NjAnph804qALb5hSLQCUVjfLnI
/gqdlQhkzR75vrPESgkfxckD34ELVIYbpNcr7azeTbJARWndhhJWU9Zs17lRYrAF
D8E8zXmXoUe9PKPsn/33b7Jk0PIr//d9Yo2aFty9MR8/jf0JcVvtzaiW558pF1SA
j5HDXj/WqRi9BgKeOPwX28l91fUp9sT2DdBSdlo8qFKov3yDUK5P4t1IGNylL5jJ
NfdL15kdUnFqjzBD5htz/E24uxcuPmFHA0TCLK79ZsfMUnkAFYoPr1DiqmLOQjGp
70JtGOjbGIEQBbXaByNcr31/2KXacjzKfiU9PmEnhWwGHuK8TfZW6MzE3bQIT6u/
kTMf2tLGJHGBRHe4rfVnHtL589Rg/+e70zfAFLbiRO0nCDaDjomsXQs6EhypvkjW
iqF4uZaXuonQ9NgsD2Fh5+dp4wCY9MRuMD0JjaXKy05YS4ThiZHyDOZMyRcC8C7v
HZNNlM0lbd6v2702e81BZ8RyuPZkFnp/HnKXButaFT+x26FmTJSALERjq4nPQ/Ak
4Jz6pHTN4oRI02WvOX4w3o2rcLYOjC9m+enZ9ZYhV1tUplTi5LpZ21dTtHq+WoJl
uqa/yVQk99n/WAwNmoVWN0a3pJTVc8R74WPEL2GfRiRp7eJTFiAuRGiKTc9kTrCc
u3W57M8vNSi7vs0mXadUCVep1tB0mK3oVf2KGmfXCCZkAzYwBTX3GIzAHHN5SckT
cPsJga/Jy2R1il6KOt6fYhljakJbRNH3t3gdBh0EJDHwETdhEgeWtin3HTRbwT3S
aIeXoHOFYhHOUoSJX/BIncElpQIVbAox0NMRoBYVrNCPfkGMPsyYl3r3r9xnvqB9
A7UkcUpVk3tupKiPR5YXnjOWF3rEbkwptIUilKh8p8wR7C5TYwXa4MSstfuI+Z8b
+vlih51x04nokA4w6A2itu5+/zSEJwfeapgO+Y9JKWOtAZcSK/M8qxNMrz8zZZ8O
YGztfcQr85ADJtWHVKzHtPebeGj6ODyTf8Ttid7Zxaf1VLq5xVKxjsnE5X5/F6zw
vM0AqpJNa/gr8BamwaqchqGVqLu+ntKOWP/ilIKf/zd2Jpywc1aztu8UbTTrDrVy
ICZLwUlzJK9aMdPOR0FaZjFRl+GByGoitOuxqn3yTYN/KDU1WAQ+wVhk3EMXSesN
qIu3uMaLKGwsPLVgyoIhNcwGOfKBQ41tKlOtK2JDU1PqSRGdqJsnyHbt2ZhfKG8g
OpTJ3Ec4ayJoF3ATJu58Tv0TD6BHj2PU2uLrSvEVfuZy0MaWPegdJu0JvwxM9Zzq
PjqOnzTvutGQnimahFjErQ==
`protect END_PROTECTED
