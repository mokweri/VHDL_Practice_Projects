`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLNbxOTtze8oqCjCXT3UIJ5AbTIPny97cKHffGRoAe2ojtm5gLBCRuYs42bvu6YD
/h+lyjhNJLp7ezXQmhQYN02aBF6cNwj0P9PDezyYfIEsH9YY4zglg4/hlsyNZdGz
sBtdMedXrMoacvjwngoVT4chY8sv0amLDlE4GrhsKLcVR0+dLDxEE5sJjyCg2/ZM
NwKjSfqH5zGJhlGdgyX41SPaxcqepw2+aAM5lpsCVLxCXIbKq2W2g/SVcSZc1Ji6
DxDYAxBDzaX6YZ2nf48MyiO+o02eLi39d1RS06XcvPFMBpokaIlwYpZGUxvoees2
WDn+ZOZwu+lx61DYpWpV1n5ZEHeFeTEnsFUi/YFX1QdZ1jbnB4jwovkr/+PvofqG
afpgVpbt+GJuJibn3HJYZweN0zPQ+POhXMI8KaC3zAT0GjrgNdUmQjr0IRS+UgsL
ogxMsgJzfEtDklwjL5JwK9UmMZ97ey1f9ryqiW+XxWZBpIqYOvyWD6qejk5UuLIi
iNkJMhjd//AvnNMetcJof6Y3LYoszueKHd4Rcbqs9+quUxnpIJiOIFCmOHEoK3R4
DzyoUA22J5MJn55TWb+FfGoX8monr6n+4ANsrzje4sA+k6M2D4nUaG2M00CE+rOV
BKSMOe8CRqjeo+Hg6H07UGmpuoCP9aBwqk1pcpzUQiRKHbQYfqiU6L6hWMQf9Ia9
vxFO3u8BvG392FyTWqQT3Wbqepl0S7WYD2boGhSe4QE6oDFaXH1kBAWU+0KfCdAU
KaCKL4CrQSXGnJqyIQj0QjmQ9YqHccLoTVOiqd9Z6RdFZOS2A1b7AFe4YgDn/U5x
xZsI5de2E2C9K+WypuTC6fD2XtMqGsrCtsfRHUrmknNr8kjLpv2aZD+H9VVgB7Kl
Nu2Q+FGsp0+oadOXmSWltwks9Q8g3xztV8ZZXMnDquPpI1mLpfrrBIW0ETTEtzpW
kWEfZbQLqrCo7JkoJ2sOrquv8c2Dh3I/0kBd5XpLCX+rQiK7yOHR26Fy7o5kRWl1
OzRx3qSxJx+f+OunJ1VQzsuh+oj9akp3HYDX08a7e4rHXFiWiwOe+tU5vXrwMoRI
`protect END_PROTECTED
