`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/RvLLkRn3swicjfi8zO9vwWkhNWPjaYpLfRbHn2Dh1ReK4bofQyvwKGkZ+DRSKP
gQunOt8SrQ2h+kP3a0CwHrWYS1twOavTN8J0fcwwEHG2g1NTb5rdArSAt+tQ09j+
pKozFDDLcSHC0K06+CQWWc86+k4T9qBybZ0kGdZ1kM9f+wR+g/8neeGTlGJvBhV0
Ox8MgOiIImRZLbkvR6b2zcqxSmJI44YNnTZVtSdThrEc0u7BwjKe1DoBSt2UfY1z
eCR+C83hTk8sxRwbAf8ebL1QDsK6rLdRkaZQgq6O6S9RRTampi4V37NXzOfgI8F1
AffdtRumKMer5isYy7gY9+5xtQwpbiynArJatLcRd7hZC4HVlKy5O+OiPX/Tpu4w
hjsYVT7/a0tH4nEJ73ooceC3UTS4qApGypBfRjlaUgzE9vneSUawZTXI6aw/HY4T
H8IrSLHWzp2CEGOix77XRbicUVNVs3SoDRNfXjbscTmYJ//veC2ajSzd/t2zLR+F
CPg5lyfvItYWPmzkOX7Ld5ocvqY85GEbbo/CPHeZcXVGSJKIxkQkoC83dDFjZXMf
7UYI94Hz7ca3zx1m6B1/UBdVmF4ewR28k6SYWXfxZgpSeIZghHE07DzljF/Kn1uN
42WmUTGoJ480JuNCrSS5mwFqyWIXJmno3qu/ijTq6OFJ5YAsWovehUgeXiLhuXQB
IUrFfPrf1snHEZLcctyXNFXq/d8qZemNYZreIachBZOQ3VBIj9yO0sS+X/fHW1kd
1CJFQevxVITxAeveKGJsd+jVjWod4CFJi6uCfEqhnDiymn1molEIeLTdYeKHKRks
nL0wFYsz6NEgalUD+4PIcbTGOFreQ+6VUCU59nILX5OMD/eIXEdh6nLixEp8HyCi
LVKbNUhxc39Kb8saXrXznoRBg9YQDVq7SP0qo6p9OhNP93C9XtwHZeSL/I4YGKrO
nZ2zhOOpWde9jjIG3EarM3syuLwrO851N4etPf/ltWc3NNdOKMmZGsW6ARxWo4CL
7049OGHu05eCmrjyr9msQH0v16GR0pTSUf3qgbEMEIG4g4mz3KsA6vdLouKkUgpe
BIZ3A0xf1bwAOXrCfKRde5Wxj8o3LiJO/f+HsxbLHKZG9CEbbmHWdJ5tJbDv5g/L
Gci5e+wXvHVEjaEs9W20iLXRyzl2xgsVB20ebaYjDzbKpLYacCgwiLjQeKmke53l
xunfkgwC11+QdsAkCHijoaw+Bk5JMvGJh/sX9mTYSpSppDqoR3Z36SKFKK4plWry
hFuR+E9d/nxAnUa/UTdWfh5Tfqt7ZUCaIfImwV3VmrG03BK0WvL2Ookiva+0p9zd
rzSes0xaYOKwBGSOsAcrCxVojzaxs0/hiIZnazeaQQ4rFgtjsw2wtABJivdj38td
Uienxf17n5G5zSzJWYfi71vU0VPYUOD74xeDj3TuziOl8NoGIi2NxCdhQGCodTKV
46jSyUTptQtqhnHV9+lRCdNWjNcecyRIA6B0+FHAE2ZLoC7QwX3VPRW7led+9AaB
HIKEA5r55IT5YUmOd8laNilIBzkKTbJ0peytHA/57lhs7udRSe2aCuoNQUZjTCL6
N5fjDi/e1GYDudDN/PrF875omRHL9I+/Wr6NAozwbkT93cc/0tv1RbbnBIQB6Ile
R169SzBS4VKBTUPihE8XjXMc8+housjIfmrhw9Rq9/ZdncirSzbs5kRlfxsVGztm
P4eiEQqNNpF6Gm+xaLYCnzzqKMT4XPOt06fMQVpvqTmr8uvoIJNfQ9jtGjjHBHwM
XtnFRVV1dFGPgX4eb1g8aFpgB+FVP9rLVgL9KzRL04KA47fHILfZqLfJoCWAPrcx
K7SkxTQSDdbjNmu7k5XZKCO1cFMh1mvaBULPx2nVhVZxgjH0AM8a6dL+5XmMeFqZ
90rzcuwHUUcd+JOEOIOfqQQiullb84jMIK0uTzwaQgKbBIYxCze+O32nKcWTr3Jz
fUOIMfTkEjAB+NJGFqWzCfbi5PJRAN7ncQl8CROHjJm6m5o0WZ+Mi37lywYkwITF
SFd9WKq33/QFx4IBn+jKpH9PyiaCnfcHjr4YPQ7gwcKnpEPfxXuJ3RDcXIrcisbv
ZD4QV9LIthyDkOFrkIeU4X++hsJ5dPgdOHkUSf4/QtC+/yfmNYCcKDTke/ZEGG1n
AjHKqMbwv3oH+nIJRO3JD2rK0P28VhqEgbcGa2ahX5hzNAWlL3kPmHLFl4wkMTRZ
AQdkteq4DKbWR/m5ejn4x/SKGSbn8ES0CVd9Pi0M0FQ0gYme/QoLZ3n7onAZOzrj
+WhqGQ3XZnnwAEEIdBVAo2ejFQ/pXUq7x2rcxJTo2CxMTCw1yTkv09+6cj0dhoy9
gBzsUMw2XCEuUHYqZk0z96HxZB6/7774qwwWg6mJW8G8nCVUMV4fMJpUqVbMl2RS
KOzfTZdSXHSZHpH5bZecX2EtELY2CHuWyRvzgFVGyNbXJCDxJjL4reLsAzqpj06M
HPFgS3QNijEX565WDhkVKcsDFfyNEx04vnVX6U+72QTdKre4Hs989BQKG2c7hSAV
El5BWzLWIScr+Nr8TFrRkP8sRAzq5PulBR+RiUL043T/g1t/lkg4IbODE3j8f1ei
BrGTcbcNuOBbliWyNTew5/0ttTb+CKDxEhuX7a8GJvP9KUdjEwVnxW9Nvn3I/25R
DK9mTeXHOusMtDjHHr74Rw7540fn5uBm+N9BtLFkvZJCclAX6fM/Za+79E4LXA0b
CoB6E+PFlEi8dwvIk+24HA==
`protect END_PROTECTED
