`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwCQaoLwbdD4aCUcOYDn1zFdfhma4Yv/wj5lmr0oGsX4UHh4WV1ymvUNPaNp8pIc
Ln5hKCQxUWvic0dCEu5YlllgQ1wE/QxnjB5s3uQmjv/2H6I2J9yUtltjbsXiWg1R
yJboRrLNhzy+duwKA+OJL5VZdXAmIPPGuTbSiRrm2RZ3Nv003uvoYbjq/9aB/5lY
1OSvv1XO99FkyvFmM5pcuIvpKZBwg4wbWddQOlgAj8F3kpp8zz/xInJgsCe66Rln
V5Lrksvw7gVy3cT8vRrnKd1pKh91MRNefEE+R6v2wIB4i2nqHHjmIjJnLsfBlQKw
l6PiiC+GSCz3TeQQAM2npOk5IfoNZGsA6S6FMUx6y8cPfJRHJS2cKlfKtYlouM8F
/R3HADj46+ZHEOLQD60pG9jFHgZL9+cUuAds8c7O1KL+/7X9Y9+GZjsfmZ7fXBSB
NeRmqi0m6mIkvPUezfZOEfwp9UQDmyHStih+/5VRN+bYWp1ZAtmvMsUCmFKVR7nO
Y/q7AY+rjroFepOr82Zym+xCeOAM8I8gpYs9gbdR/f9L37dlbi9VALVCHR8QIiMW
j+tRcI15aqK8zfKrZLq9CYeOrQdRQpqwkbcqTwDe0+7ZpV8i7shfIgJ+68FkUJes
x4b5x1bVmwY2xGEsVvQldDAJyWJcJigVA07Nz5tfUIcV7vq5uulFG2W+CrOTPid6
4T63/Vai+rYVHgNJ5RymkAJBqna5w72Lem0rDH9yCsRl6sq2kq+SweKcOqb9+UcB
YUlKK9Y5d+biFupoHuYS70ZCOvxUoe/r14UkqY83TFuGMihkOPfaIZ/D6HoAwAMo
3oY3SfHB4ELxz47hWjjcKWeOId5CcQ1wW9eolxz8268qmEF2NhzQR71dAkMhff8g
eA6sg338KiAAMhOL3v+ei7ftdFht6dGoobqTDx6dC5qROkgy20gCcPuR6aJCV+/I
ePCZqeZwsVohFbJlKE2YBoukWQRBTh7VOd8VI0y6iadItBBp+cCBXKV4EU2BZf30
RaaoE3ehmxcUlQisVnt6Ag+6YbjV76qp4IoNvXGucBFrP2HHOENg3zkedF2gLp5o
9XAf7V4W6sCnC3XICMo5htNt0ko/QA2onddzVRXfnu0h3dwV4JqVXs2Wqz/3aidT
Jwe52bqGBrjZJN0fPhtdIVum9erzFqLNPYJH6H/JHz936Zd/RJCZYZWGxbOqZs+I
CIOR3XFZeYASqGV0MpBvZ6MgXIpF6a5FAd/AMHYj+d0T/Nm1lpPQ8wyXnKQHzvY0
EpCE1JUZxICydwRaoiJfQnthoiDd6aS3g57NeTUXoCb68S2EHONRH06tbVetbYCi
4JQcbHXFPIp9Y2pZQNuk5R0tTNe5c7UGASwZi0sgfIIrFwtMZpa6cw91Ipz3eEjn
3I1uzUvlcn5DA5s4tVof2idYvExbTB5yBiX6wOKwxEvy0qB7XUzztjlbef9T4QV0
Rr4nBYFPvDSOBKwvNaYGbAECWymcag4UAsTZ76rfa4MM7TxTixfNyWM9awNLaztD
mhYPlZR4KMeZxYkla3knJkilFjUKos/P8QFY+poNiMQ5L1Qh1CpALGsSz33dGAvt
fTxJNfgPOf0cWjCtblxRL3Khk/DlZkap22pehMVkYSwj6DKR0CAyUiimNReHdpQ/
G5aEtgQyEqptEXfVKT/rmISyY1mJLGT4nLOhysCiaNMCy9bMZ6t6bV7Y+gwabGoQ
xXKVPymsvlAgh5PpNgpcIMG7EG/o9BARawO97YQ1RSC4ulgxoD23zJgtuFnu2tl4
+VKEoOc8Kj/o35xVQp+AVIabl9zMeGV7wbHfa4oAW+M8AwYvxl2JpxHlbRrxSSuA
Eei+1b7g8FOHvYknS5MqG4CxVteIde9ZTW5bIKYmb8JUzAFUytK9cURSaEfTIC3U
IyI/cCLKo1s/ZKuiofBo8RpiLvK+CcrQld37+e69IxoccmdWAGgLVk2/LhghFftV
esNSMU0BsQbJNef9KVTGKhvVJmArWJauhdSWeta0cAEYqAdhj19hTk5RwAM2hc1k
W6y4qRBgouZcKx5okFkzPg8FW6HvHYqmlc4ntJ6N2lfipoGOIqBCgBi/pM4y7kqs
DxldYCLmfj4L85siOd76JXyEbDK8VeaUEen+RMUD7LIFoQfQOrbDbc6SHHYAQOjo
2b4KBD+yhwvgwNuuV90L7EGJnsfUB9bQdQs9gE+vNuh4sTgyAU36Ks8ySexRHB1J
FBN9Ze6FU+KOYpbv4YfzzKm+GfqjUQO6oR72b92yHi55wrUfFuHjIGwp4ICbjrnj
fVwaeP9PSTVt3fBvPUKQWL67CXp8IvD5ZJOPex9pXGtFsEsa8OOu3wsELIhnrv6n
pc1WFX9BkSqkj2/cTr89gykJLqb5OhpoKeEAsrXVGDFlGxvtihV1Uz8yE9Qio1Qp
RWn+b6A9wgKDh/iBSnBGvhzsauRblJGu1l9Tq/m/SBJAKcgYRU4dggyQzCNzdN6g
9Z0jtPdNs1a5Jq2n3oEQGXHJe2EpFsSwv2IeHi1bUIJ9Ny9f1HXEXMLPNNWaGZ95
9ElVnMXQ3X1duy7090MwjG3WZB2cJ+yEHkHs7LAxeZxJwEw+g3KdxsybuEWl8+jT
Aob2BitWY5AuXk4CW9pjd7U70KTfBROlqShpyBAYu4+Ol+SVqge4tQ6FQIlybi9s
+wkhOuj3U3G+JXOtd8TSd8mqRzI14sr5rTYMmTJAzYH77iFmYuOyV5td4ToBeuzt
W2bVwrZxnbfZcd73/FL3uQVT0J43kiUJq9xAkQali/Y+p2PVm9mEx8qCF0bdYDc3
vdJd/FkXfTLq4NzC1BW6KzUU7kNiUOx1UsNYnqlZjMRZ+0lU7TAFF4pyGZiS0V89
VLMI3jL8b2cpf4WjVRSL0ot+Uh0m9ePenjO/lNMHr7pCFvygRdQBX4uz3yrKuYRP
toJBSmIsq4Eul97X+BWwpMgxhShsKOjFN2NUGKDntYlYimdy8v/+VodlB1j+eEKT
LkibxzYRw3kzX65Zs/Y04TCjvx/xFEMAwHfDrUwuAqMQTQ7XHjqQhQX3sCxEmYl4
jUCg/A89UU3Gmk3Crjmu7nNlW+aU+0CBG7NPvqs0Zc7uJaIfGnMFCkaBkhdUf65W
AYeFY2vdDCwT8h+Bj4WZTGt/jAEXhhzjsZoj3WRwMJ0aA1I+RYUDZ/vrCLqpJ0hS
fSDaFhl4B0sbUQw2VeTTscoypyP9MAA/CqIbBcb4hjPAMkEPq+3qf9A1zjI34qRI
L4Qvc3VgHyRIV4IhppvpLm1KZuL9O5TcwZRThN5Qc/PUwEorYVq/cYCNxsA4LUaO
tzPiDGZrFKzYYhvpZAX5Wg0qG6PXKBDm99e3VGoDXmJNCzLKTRK2AXIiTjY+r3Lc
2xTS5zUuyXDMlklUv4CWzzFfv0Wicirs5M+j3/8cZC6t9FqZ72nyOV6Ih1Xrwq2k
w9M12aJZt13RBO5XXOHCj5LRpW3+jEJJRgBMri1rqJvTt75v4MxX7hk7RQPtqfLk
i6d4n8y3Myc4ZdM6S/Cn8HiJuCYHaBeqIu77Y0Q/O+KTpW8Gc6rdbDcKz1fF8r6D
U/61g1IjULo3+NzDg5urAwQQYuZj8FIq/8Iw5XnawrF9qUMfYhm81TpXqYUQvQP7
6WfXYcxRjh83MRgLAUtnXQ==
`protect END_PROTECTED
