`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDilU1yRA87L38of9LWp0LuHi7gyi7leoyvmdQiyFUgWIo3QrxhTOhxXqjMD/HoP
FXcME2p+gRujhsl3bnWbPFcBtrINijiOiCSHWD1RFt20jibLZXi1DkSvLvACdgf6
wbw1Uj63TVicTCDePDiGzGgVujI1n7W9lF1gN4gAbziuajnzp4jr/sIntn/AOG8U
vigAUIQ9YBAi+iZalyrq02cxK4u457kdJu8KCZNrvTwqU2aPuZSkcZ17EQ7DBnyB
yaT9sHJpNmuZjcSfuxSluiNbDgg7yVBTpXxwzJrV3dSIajWHI9GCXGbomdZsLGRh
43mH0i8/PKxuBHyc0DQ6F7UzoXrhMmR/WcnhkC0llkef+EKak3MbOkCwfqW3NdHe
iEQvRug50WEuC/1jqKFG2pdLP/06o8F5LUERRuS0wU3wj0PJCnO0QJ9ynutd4qjr
Hb33TXfIMIBqCVZhA94tEXgN5IluaXNeOy+LOozFIUc2hhpSHGWGT4PFXMnZ1bbd
bYBay5rb+3p5tg9CK68V2wGQyo84qPOpIKATyjjAJW2cWUNsyzYVQrm4DsCApqis
2r/lh0Z5FuywJMIOhpuTW/b4EsqY8JhM0LjFXRstlgNTvj7e8pVzCw4Qh28fBbwK
AGlyN50leYKcScu68J28qEieP97FKRyy93otvnYfTyvHZwVLADoZXeG9zmghS8z1
hBAMvylzKVyrR2ahuDsg3pthW/87EcE7K5Pl8HTMra7FO3N/jvymZW1Z9Dg3Caw6
H10l0AZ9Fl7Iwarpm7w6taAYwGIPs0DFduYdkkzW40UBA1PyT/l2aEh/2CQTvmbY
Oosd5m7f+rVU9Yl4BGGm/6mEMSSKl7ifyOFJibOy3y4IKP+F6ybma6cGvQ1+5Av9
MrSh6DxHeHPZ21s0QljdYrjSwY4BvuXlUBMBCwwNav+3/9V++so06877/+rLWymU
gQ04jmm5GtrB38Q0u1Z4F0qlLRLypBJuOtxWIwCGezWAkZMJjcMeugWN4oCJfXOf
8gwDT2g18iEv0e2ZscTX12gQ2Nrc4Fwk73msy8jkfk4feKqAhgZC7Dqo+gmWNDaB
Z58F6l859a1BgJohFNiXJZCq9EjQieJgspKSdbI6lnIINwYDhQ+7MPcw3PD2R9M5
6J9TaYdmiatdelvQbDpuCh33estF1b327SPj3LPPAyAnZw9/FN1dLzx+PjnwHfqI
CyxbtQNf91TN/JthbJs1Xr4tIhnPLgdG9xY5AD1TKdHyVceAOlxEpI5Yr5FpGsIF
R1vOYtr0CIsEPLKo2lpRRnocpK16COendPbZunsgeocLctpYT8YwAMeuQNf4FCk4
MnsAsqPuAA2q8NX2VkeuyN+LTVrLCjRZNoy8fGKUOyqoQj8gL9RVgMdgW+Nm4yeq
Eb0weu7RGUjSVVV51Ets8XWAus2GTLV3fWsJqb6I6AU=
`protect END_PROTECTED
