`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
isDK+kCU3l6wKa+saq510dOw3l3eZ+3lk/ZbMH2LfvQ0dk2OCZGmVHCqvhP25b9G
N0HaFdgd6h3msT5psWjJs03rr9quvZvGXtjXCaUU0Clmi0UJl4qs3PUej7ubIb7/
VqAQSMYhkRnJscNjhjLsgClOh9rONq8CoSXg0KwU6M6FtWaPBSv62BScEbp1jH8F
eS2SlCg4UwWEhQfCIHdkQK+fB/CndeI6lU53YCggR+MuGmeIfvDq5xcNiD6RygrP
cQJHcsXOuZ74VljElvqQuWCp4loShcEUlhKCKj8vBlmBHQWqHTWYxUrK46o3GgF6
oAjmvQ086ddOO3al5slOcGjaxkB5pShCjXgvrmBc8ROWa2PZGXB3EssZgr9dswEL
Z5lCXBAcXibs85K5qN1/1r9lbbM/wuWxT64eGe504AlW+8pggJc8gcGfJubgnavq
z21ol2SxjVLC5sHaajhGuNPOwaxWhv7hHVvXScWlTNe0b6fpmIUg3bD1h9QpRzXZ
TmvEdNf9Ff415NJ8E5SIOtBPXcQtJ8A2Wa/iaMIwUmdfyHVFK00TlQsqHYEUAQtY
JUXtGd/tvv77C3ESdLUkyw/MjRAy4W1QWAzL7RCCLBMOC8TBRSXQN9Bk8Z3m18N0
QAs7neUzWURczxf+7WP5ga70EezVQH8CXLu9OratUMszP2VNtpNN4GIOu/Y3fGu2
t/JJaGr0TpCwphkS0izIxtnjlJgIWIMfb47DZQTSNmlWtOprJIT+edpuFpcz/uxg
V/41FrpxdCNsXmVdSD754qICD/qVtujbGrNmTACE29K9HUQAVglm4+GrRGuUqLw/
Dha3eZtyYHVYPiTk3hLyq/0p35a9Ipriq9qmlaCwxccsKbzo8PsvwaUkTAip40Ta
PUCOJ36yjP+eeY83NeQwjUErj+8Xmzvby5TDjAfjHryGqCfMAxE/zwihYJnJb5o8
HlcMkPik6335OBRBfo483FbTDMZoaz4nJy4UGVdIFxsGPosXrwL4akP1bWc1Oq3a
8DAP2kEdX9XIuwxQRWT9OqJgYZBRMqFlO1DMujYd9IZjV8igH8XnT/DpWnK7ZkLC
xOW20HlfGbe8W6RwTPzRxLkCUJHjbeCYuKiEqKoflXoPAsFwgFyqergIozXy8+5s
fyVXfUPLzl/zTpyObR/GUE8MJJCJauLljd+HXFD5OF3GRgqn/M9cv7EY9aNxkQ9L
2zeObeV1ByMboNisUTv0RDRt7ZF1j3cLcaHREcIBS3viJLeQ82qItKRtdti28R2s
EAe9dfP+gDpGAY8N3JFRV2XG3qQ32XWXmn+YOGbxoCdJk0AtvwhyoZXJALXVTPAu
bh8+E8+zBydwDN359+0cd8NwtQx5F/uNVq2iUsDDBQLtoDxVcUd/WnsxB7xO1qpw
bl77qjCekgKBkAqF6VOBK+faBPdH9Qv6JSYHWB1IOG9nKyUSqtuHat74kNsgY3YS
0AyQiHJj67V6qI8qy3Erb2n66iLSGhEh3vGRu2S7iCZBOXjedm8aAUpqPOF6WzJg
S5dBZ3h20aadrtGa4uokrWCklpCRV8qWqACuVquOWHshvEVubcC5+2/eDryZTvIP
Cudb5tp2TuJXMr9/6zEWE9zjaIcza5W0teA8fVmCab6gTa1CbkIDRCeejheoLtOk
Du8ogiX0J0e8SBGWrZLoRCLUkDS+Ur9l1mflJ3oLGs5cUzAI2vxKA7tVs8TPxEmM
R0m97a2SuMzNwkTPcGpuAq+/HMVJC8aHbkkWrT0ceIuYXZrjFKFa5J+5vx74mxfg
Io92a83hZWVbA4TZ2Upv4GLX4sCEhxd3syCo8avdUZLfQ8VxL84eYZ8momDmWL1e
ja2Ke00qRPmwdfzk7drKY0WWaZLTEdGlhjwuoYVAL3c5/ltsGu6Gos6/obuwXvko
d7a6JgyaAdjSZHtMNR0K071EWersAA+A8RPiIEVjSws08v5ZmWsE6cAekzM6H8Mf
+XOuEbcyKWZBuUPugFyTN/uEjNGe6w0jMaisIJRYx/cMlzEeoPSr+KXwA4GgH2Bg
cAAC5Ewc4dIZBhoUv9MnD7dQvisuZiWyDLvUbQzXA8NNWzITnMHLWck/cyQL8pGt
MyWkP2gm+ndOm/K0EcBEpkjQ3jvmveqORN0YSitup96HBViWBTACKO8ndWXUnQed
u70LAuzX7FZVH1Q94H6RJaHRUcmyht58QZE4xyivzVI=
`protect END_PROTECTED
