`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUcwfJmefjair6OnrU2G2C1PjktLro7n/U0VfNza1wloF2omxDBMTuv3EisSShaX
/rToYkz0EutOhwf3H62OGbhEPbuoLFjGKgf8/P/n1rtgHX6eD7hf79L8Qmtny95p
6jRGFOq2tEm5lkw0Sxh0eFqJE+D761h88fNcPkuQ2GHn+nx4O0mwtsjmc5FFEctt
+kAmSmay3U/WhTlj6wPURM65Gyk8+8MfQ6mfb6VsIc5QDsCX1TMWyJBvwgGjXflC
7dU/VbNcEnbYZiO7L6RspBF0AfCtqG5f+OrNBzbSGReonoHWYzo4qg4ijXF/YodT
DMPagJGmXb5YqZifTyeA0VRplo4R5wl98xu6lKb5ab6OSGRAJMLsoa1erANptMv6
ll+oEgQI+T9ceTJDRIziH84m5FrRofakOwxWAIN8njXCqE3yv5bsgnj/rR9PIzZ3
2sSqce8Bv01tUxbd9WkQtagkhK7R9OTquojSjH1w8S07HZR7JbzfZNjONsl7bwwj
wBiuCafQi2uGQuyJTSE3UsNCpCAqT5F+U2ZN2M4ZhOF6MhhIKAm5CkCVdoPUZ8NS
DdRUPO/NsX42iV9MQ4+StlsVLTse3OfFZyGmN4Bk/cqbN951aIng1WRKdVe743YH
77ros00Ir44niPflf7UaqsqrcroZvtm3LA3GEgrtOC+MJMYB3Qnwf20/7IwuvnC5
9FLZ3ov8g2Y63VRHrKMY/5GBZZgBtlIeM2v2x+9dwxsj37ul6LzMlYjEOQi5zPvp
41b5Ciw/OVXK4T86HSFcC68XwZCzFJbg8337DAr5gTZSyIvJioWIEnkCuaVNV/OE
gtArhd1Am2bx10zG7gT3fSZZG48fxwzBFBI/3wnGr3MaLTMvxCrPVJavaQ436in3
HFGZbnvXwzre16y0fwL3zh9em/yxFCbVmy21Luvq9whtQSMNQrbRtN72Sx7FIrTC
ApZHMWOL5wFP/6Ploa0oQ1Lv6RVH3s6F7NU/r1w5E9c1DGj499mF2jTs0ey+wr/B
AUQJNC1kSbDt0Y5nHa6TJLisxYC8ZLqdt+sYzkmQVakQTCPkUSK9mrQiG0+cLeYm
hewpzPtxkoHOjhWHiJc0X9xGlcXYJnLjem3K1UWrrfnnhzRdfRkkP1rIXyDU1X8p
xf1hn/tVt/MPyrQyzh8cfO8cgSueS1mo+Uk2d46gfW1LIW0RO6en2nHB9EOT0arg
bALVdkcTNaaDvmpkO19UFbJHR6SYk+wqXjDjClvfsi4os1NH6aF/csEuv7ko8mo0
Po3tPk7MFRrOJJvVfH0BadR32XJMzMp8wdioqaAVwyH7AEvHRebhCNiz7eu7tlBY
kdPCE3CXAYQq9MjVbcSDcIvQmbCzLUukGhcY19p5Wa9e7MMwlSB799q+zv4n410b
l4OiBK/aVkoKqfdSlThZzl6Sn7Gntu7WDmjZ5JXN3DEqH+yzf1I9fHvbSZPUkAUM
kS8j3UxaADT36iHd8bFLpLTwvfuHceWQw/+d73/QGsVU11lTgxMZ3ucDCAQ0jL2R
IsSddDtFc25A1GOJQRZXAj2nQnRaGTXFU6UCYXZHXAxU5vue96a9rNG6Eee9B17y
FH2d4zAgyF5l4s+Ixp8TnaKd9E1eRc5fPgYmGp0c7r4SOnoV1uTToYJNhb/lgq60
TY1UYWw5CqvA1lPoMr0JT+eSUetReeSR5sMO2VSrM4DWK3fJ1vhTWSnRo116S4in
Qg4ALjjVnSIThZd3ySjkh4VHDmRvLEEnH4zGJttjo/h4qbjkXRQhu7IXd5gFKn63
tlxbGdNlwMRzAYiPblxwZr0V7rWG/hkpJcNcN4UNbLyKFKJSEyViLlB9AWOallk3
6xzU9YMLh232PoymKVl8KgyZCSb2FOJmOlsRrxfdUXo5hJEnR2sNFYw/ZtOyGu/d
WaN0Ym7Pz8S1WvCJOUQvpn61UlCiRBq03M8XynqPYmZO0aSvBfToXC53uPfHwSEI
Bge0aikWkWmTxXOafkqMVFCwaC9KG+UHOoj8Hsu7ulgzXDvdmVs67dkMEbvgfb9+
auNRVNOkyt/dBiPjEWNft9tQFRrFewrV6f9QkE7ELAqMiUNVoAyJREvUz8OYnvX/
UzX5TvwbBtCOcfp/xQbXEG7dVB7xB4VgTGxInoObMe2usr3bsIcALEVVtnpaTp+W
nVu1Sk+8PHAkHFGmp2ZTGu2T6Wf6oG3MUQ1wRjYt0edEGnEYex+6AQQtu733vbYr
Cy50o5EGq3UQRg4pw656B8fTBOTB5hAYwfKoc5Pvy3AnvVNKcoxENoTfNvlArDYA
/bROudHil8b7etDoQKoyT6Om1zKESG3e1MWLSwaDDLQE/skOUflrew+0kHK6C7e4
wQjXvFcfY+97gsDM5F2Y3gx2VM/3Kgd8P/E35OtfnEuiIWnrYvmqSp3c/VsJbRrn
`protect END_PROTECTED
