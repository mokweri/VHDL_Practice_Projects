`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUxuJTuUaWMVyAoCC/JQSe7yLkOA6/2lxoXKqKzqDRarsWeHVmXOw5scV/L5gCWw
+n2YcvAPQuNDTMDZEEqGU9v3641cU2ZitZOTqHS5GY65iuWgtUOoNmvexGZHJlQy
0iKvS/xNPs1WhO/l+ly5kqIiX9MYmFt4jhXxE0Kk4f7lrufz0OW+PF2CXL/WPisq
cEDJnkhBqvXgGuOnSL5HJiULMfSWm14gHkW1PlDEFrnxHhQ8rmVfM666tw66sbYI
jvcgKBMXcyh9rk9SJYZB0t2MS3P6EGnExVh3+F8Na47t7vfS/N4lWHoRPLiVfhKB
3klj2GcDQBOdrCERellYwrNtVSVb3QmS6if47NlJyFNLhc7RdRVYbgZOR+UuIaGP
c+vOP7n3LqFiC74Tanxb3vhTm0lJZWlhxrpJg2kTWji+BSsX0DhbzATYPHB7pMFC
5RswqMzwTswd/6WqnLTuwBhc3/xBygCIuLAfk3gmQO21bdzwaoWVGOuOEKteJ3Jv
QUrvMXF0DAGJ0RFCiZ0YfJXR862ZTkK71ME7niRrTPmb1ciK7TaPiI+bWGo070xt
pdSDzo1HIHc40QmpQCj6dKgGswAbZPw/aePxWQ8VPIWTtmSQpwtdEcEK1WZvLmyF
crdcNOYb0/SkZJWF2ONzrsQbYUpkK1JRTrYBao628yGQdl+95XU1Qr6mIwprNmAq
+ZL10FgRnN3NcD8oEuV4iF+hTnirOgI0AutgBAtIx33nOeLSsr1eGzPB45nn3+A5
bhOUWSCGyyEZ1kbLQYG6kGJUBoXcU/DWvFW4Hp3S3554Mvt40Jx0N4jxA8Ljmaxt
BJpBODrATm1srEioNqF/W0zhUv5EohsntIVY2RJjMYvEuN4upjxOZgsCyRoMDdJe
uDE3Y5OnNZqljKr1eCQPxYjNnd+FTUbkjbH5YPbbTiEU4s/ksnp/ydFkilut3rw/
HfK11Kp5+EpRZQHvtK1JxL6dkoPycaZWeu7ymdD8Y/orlRtxjvbhnpn3s9EaWq97
uzazcukMq3wAMWpAc/WVzt/SY/nsaRdEz6yJVblyfmjcGbHs/eenR11NK+HwC0FA
ryvpPHEG+qljnt0ThqdI5H9T98ccmP/FJlVKz7nNSQsTTfLCrQOfYB+IoOvIeLRw
9XVjTKHCJKf7AwB5gYGNxcpz9jf0cQxuoPGLEb9gk+jwwHXNxOv7NmrSRtSL3gwp
j/k9DYpq3rraGhZLYsMfvFinhv9Ch2jM+ESl2+yQG9ewAdrQ+HumlLjGAcDuUw5i
1G6N0qWU8ZaULWBL3MPkw6mmu9vkYz22GFErFnq+oS01Nhpti2LIkX5Ndcnzo4X1
x+BNStB/vZZ9KP6/TbX1/6TFaNZjKYOt3MXOxW95ba7ZDTQNzwxVBaWbbcYAtlLY
HkK0JuWvhudZZKCtjMJkLBAk+5URsAcnXu9aZDO8ixhBiZLYT1EnQos1nKxN6NFO
1SxY8sR4ovl4IbZVQ3G1R3mHAQFe3fCzCLVVMjubiLYdNiOd21XJVs2vDcXqwGLX
xW0ry2Qou1X/7IEmEgqVHnbIc5W2Ly77S0NOmEyEXVzMdC7m0o1R4hFxcPgOkgQU
zzrxBnAUsJfTSRwdMVatn8Jg4kdDMpkrtD6iEE8zQe8Z8EVf7zIaN//EKpNJSA+k
w/Ih6Xak7jLb4IuzsNnVS23SOMEdtuCP+MmKRHno3lbwu4T8gmSsY28nCg/z4ymP
tcYM2cUxveA0G6myvpkelkmFE/zgyHY4YvhL8DYVsfBQq5G/cBw3FHnAKxEVgDdA
SfyM+8qWpPqG6W2MDs5665qnXhYdJltycLPGCxIKitPS6Hc/o3+9tEA+y+uw6hAE
b5DtaVipSKt8jMXJLSUsa+d0i+wYtTfQ0IEdk4gYop2rxzb/t/TywhpdAUxiQ+eH
TImJd4yhFsKoOPlknZjSE9voYiaCV3G8JkKb12jZFp74HV0T4mqvlDI1Jycufu/Q
wKNy8G39ygxvPAs4i92/TRPEuyijmskKy/ieMDp7gu5ulgs6TT8U6Yi3UfdJ3nFq
+2ActrTlp+rM/rbW99P2YJwUicqWo75zdSo4w/enR+ZvFqgCycMJKpt3BafY2y2S
YGlSqxPayI0JLhXCms3J23qhGWF9IA1bDqJFnveHAvwNPwNIw80azPBSYsz+Fbgt
L+el2vPfZwzGzSDBJp4sXSPx5dv/NGCjtNxfH1W1L0VtSJLGMpU66tVQ7tDUArPQ
hFpSZnuQ3khDkNVY2SLmEx9p0duYwE7dyQbs6GXbMuQv8DPhIhnLGq1Ul0JvjB9p
V+VIg00aSvQN6obW7q/eCNCG3XLwZfkKMWs3zzFsMn7bv7/tL+eAMbwIlXOsfWVl
oHpzuqUkdbuj2Qb+IqFG+salW+778MM0koL/Prk0j/Q062WokSk8fMfWTlqCh06N
hQax0wC8OQklkDf1SRmEyoLj4+2WbjRS8IEFqGh4x1XwsgGwbBhrvtT9uD2Iy7ja
8/ghfcbQlOKzp6FvfTUl6oqu/Oy7kw+G+BEJLgIevnqlYz6duc+JohiSfvjzfLXV
SRJKrPkTDdYWS9SJtHht34n61Dw/7RRFhmggImyoNApqOfOmysQeaYPFLMcHaBvQ
G9sBm4WAIMzMny7MASZCHrUgEvI+EVJPIVWdfX1yD9NrGPnAI2KHCUHgEuPCGQPT
kjA2VQ/ag96WKOoRN9LzwQHttNGV4dn6PqncwtFehi1SHnXXzApFB+VL7P0sJLaw
FmneA31QBO+aiZ3KNNLroIcBbjzUY/iF3bAFutFQJRpB6sl74bV+RxJHIL/dp8j1
/VkrvduPCS6fp5dIGA8c2lsmwMMJCTSloI89gOw0h0sqBOW0U3McvQUXHtrC1jty
ozuCRQaRtW/GL6Z/bV5N4I0px7Q/T28jSe15eZsetCoG/UDARVyFahDkPpW8oSzj
sDFmJGJ+Y7BYH3qm8g4BmdA9uBqsyIMDsap9pRj2PrP6GJMa1lBHLwt/UH7hM0pk
OozaosBuz7cRTWAst5xXAoE1htlckfw8xruB42I7zvJFBp7Gt7MQKPcT5Lz1G47p
l7WZr9r4s4opl/tDhbWEeSFNpH7sbJ0mXdlxX9/aYg/XTrDa8MFJSEnunNdYVPgZ
7oOVaUZFcNeYJfSo2HAxro62t5wyr4xx4bG6r9gqrdddwc65y03Ns0ifmLU2CJUz
K4A2UP2DT8dAAvgTgddg4nHbYvanipM0HvoTbhZcObevrHegu/9zeF+x9Wy9zhh6
4LtE42+VKVBxY0Pr6SvtzLxHEetzth8bJVmHW7xD2lcFtU0NAuCZWeRYN1mPPcN/
BTvL75YxUh/zVMQZclj/LTDblA/vCboWV6FEE8f5LDxEhDG2Y5rC4NJEudi/lW3+
LYihM4aufWakbKnXLX+W5n/kph6eZhcwG3/9WqA9ROGRWNN/L5/RXAPiKI2RbmWF
Prvs8WiPgr02ltTO1ol2sFm1YR0Hzz58sZ++3gQeh1UHKFBPr9Oq5MrdauF7aU2G
hEa9DFeCEXUWXsH6igvzKytefwZ9sGX6gtO/zu3RonMl/bKREpRvhleWiC3ZR7ui
F8lFKeWz8aKL0xRu11PpzkAUT8LRjucHDex3+RnHMC8OErn+L1iU/2SWgYTyEWuZ
KxCMRYjnT8bLYq455iIq8eJ9LUX3CdY7F7jMzdFgg05+faAZpL5dpe+wkthv8d8M
3JGaESHE0K9TvI4YRb86QndtTSfjD6+haFt1541gaP0hjo0zE1tGKYyKKUqol2R+
YMjxwDwR1/eKOqaSMp63Nc8Rb858sxnIpJIkEW5zOFACb75N2eoOJXUHwYHeUo12
HmP+yFRq3ZwgcigkVTp66a5ZKS808W1JiIEpRV8uW8wea4BCkWSGDfZTjOr9h24+
YlrwumwQYHVxOQJY2iSt2zne/Y0Qg8N5e17Urr5qAH/28CZuMsKFlTTQakgY9AAX
3uMQ/4zYHBxlesDuKqyl7iM/NrBLdBW1uPm21A5X1/ZR7d1pFGdayGCj9cof95CG
EOJFkBvWYBAcbuANC6jn0/SQHVtcOPMua6X01LJRwLsFJT9y43ZP3+/yD7bwDoo1
HFrszdIbhEPA9uefNH+VMS9JWBtsaLO3oCKz9rVdFLSiDzJOZH6naeH7vxqWSzEh
e6UpE/xWKRtSkTGxPqGmV6Tc7T+Ta7rfAtV7jUWsxxbyj4ZyC9pnEES+XvAqB4T9
UfMtXqq2BzN61kuXWRa494zWkyg5oYkajKYbxfl0u2cO8Zemmk2UMw8w4SjHi/U/
lgGtCdpmVMWM4/oHkQ2jWAchItO3IiIblEmY45znUpI8rwbFTSdsp/FyNPwtPKs1
YZOKLssS6tRwiNkBB/bpJRsAiPGy12mAbGE3hNFT2nim0tZshw5s+7y/SUkX3XWB
uQsn/MwgbT5GIu46pzieOPuKWIRZ0g2C3rBL5p87VuTZpv2noCe3BkZJLl087ppJ
w54T0EGvX8DmbrSvKc5jZbr7SPcgXsbAyrnXe3uLsJlU9GTCNnORcRWEhg23G5Hr
bf68chH2MgdaS4YzU4TJ8N5xIkI4pbBVeshnzlKpmrR4xOmvhFgWsdy4DeLwPMwl
ZjcVPaPnXeOR3fMkDez46ugXC2697H/kybsP4AzZk/bPb6fqZ9uf1vQs+marGbYC
xDI5f7SuGV8dfcKG8tY1Ty61iZF8ZWcqQHCn85xFKNeFkQgYKKeVgtmW5upkotbs
oPxn0KjnIiSEp+PBg4mTyLDUeVDjqkXiLZFr4JvPIviLP45nu0stBEnn5ScfHgXj
I9OkrzR/knjHbh6A40aU810ezSrwubQTiW7H6NgesKun/MDxb9UO0HWG+NtqMJhR
cDcPDfaBYqxxcbUTC6fEumrXCBhDzbOpqaHk7qyuynICduUpc1pV2uhMq9mA9YBY
9yc5sTArdajOaijtrXR7tYvr8kveWznWej/qfxb/oVlP4FGHA9zqWxZs4+67JFj5
/C3Ap0ir2icuESdB4fWbedJOu+PnVjL11kIMN8XHSpihTbzvMY+Wc1ZnZuNeQFWa
rVhlOgmLCgz/OxdQlcojmDxmLkd+LHSVmor/LT81DP3lPajstGMoJFUeO3rXAcMT
A9nHz81ClkyHepZX0BToDE9+IFYeARTaSKSCOSCNcxpdHX4J1rnfaWeiQTVUTY5h
CsO4xE/Ro0Q4pWoL59nzzL/RBV0H4o/cPl4F4zI2MFNMH1yEak/m5u1dezJaWAdy
c9krPJ1qIbnMMLHPkZ06dQcNLgluYSxn6iMhxRHY2gun2feoWWp4CBTwySBQwmng
38Trk8a4TLI1BlO9kov1YldvwGKoVsJeRgWzGSEZqmxZNzNdbDQY8XOpBxGqub9W
ULcHsnomRS1vRnmM61ldSa8/seY3AeBFroJMyXXUHPGSm6MM3OL2VPbNzVLRiQ6d
mHdb8Mrzg0mj9Bh1R/NwOXGlhIgbogU8+p62CyzyL9dyOzFfr+z3cOGPpayh6ccl
+E41lHdHiQxYpj5c8J+8qY0wqfRBVu7M9RwwjYgNX093ieoq4OPLtPDzdHhZpyTq
YKFmwa0Jsd3i0UR8plY729GzB9rRiTZzGqCRkDOIQtla8sqBMx5McRTKz8Jn7Ina
Cdbre6aj7idfmoBsioH6Mw==
`protect END_PROTECTED
