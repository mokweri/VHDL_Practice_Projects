`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQcq3E6fnZ1z56yDSD5ARa/H67mLsobVDfuyze5TNUfjO5qEUkYNY9AWC7qAkm6Y
CHEEyw1LkQsNmVPVgPdEOfj7TM9YaExLFXD8sUttB44vVJ04QQULZsZUphHKdSAl
VnOOLdt7eCy2nS/FdGQmr+QsRaYO9/RvKkpoq68S0T9PyrUsOscj/+iXFlSmDRBn
psBZd6HPrdaXO75kY1Tq4GRfpY2TtP4UA2v+qH4TxXarrnwc6sNS3rEUNSQ1Dk3K
7qIrgueWKRWxvbk973Nwwe/PT12o2TJYxvmqLJJIV7Yca/O5o/e44UlVwEvlJcq9
5GH3/mt86myiV7knQLUVLOD7XbAXVmgSbEeVv0C2TtfhOXvtqb5g0T2Lft+XRF+Q
WlWbTG5lL5mgcrGgVAD09Uqjru9wpUuMRy75LexTZgW7hA2Q9KlyHmack3EUkg1c
2KmbTM9pgxsl5Ox/0iaTUqZq5ADAmwPqTaDb+lYxo1RU9xydFpz7p1Wo+BisoRm7
Gxj7roZnK5VMHkznpRNUHf4ch9ZDomC5ZzYSZMPUHDqj/OeB9rRm8AwopHtDQMBN
CI8E1I4Jlafrq7kwvn1OAfrzONdCeUld4IpRh0oR54Xw1FUIHRy1ys7muHLz5m8t
cnhQAgYECKCj51NPErEhoVqJIxFTxoSuizyQphKrfdPHlZO9NmdxzZawp/2cqvyG
W8OGgMb4iLyIl12Z5HQQOAxAcct3Ogg3Z+XKNc91vtnhoEdibU3SBjTPpKcVumbV
2LMh0EhjeakQrqCTx2uvycx9V5kSBRsJuTrmGURih7UlbyoLfY1VPt3qcUMkxY0r
QHHilK1WIakx/D16N+vRH/VJsVP5QuNDmvESgQbqRkvlUEFwRcFnYzUgcP69+xrK
7LpnigPCgbN5xOdlfmXJl6MDryG03lvjtjb4yWFI1luruU9+CCMZlL6Va/cGdCQu
a70NSziZ85wH1SW4ePHBVjLSkBldUDqNcbgJ8h/Ck9g7YbaMPzLowElqOlSl2UKP
aOyMziyPI9f774lYHuPEhXzg0xw60c+Fb71nZXhijcWVulntoob395a+GxOLVScc
tqwibpLzSsDqbmA4Pu7gmgmGMN9R1oPaHkIIEQtFW7EN25nNmJ4lHbw4iteJ5fgr
s4gvfI5B/DHFY49C+/e7+J3BLWhGhAfv042Z41Y5app4BBowukY6p4CAEeN943CK
wpqqDogiYRhjtiyQQ04AjiE5uOpDdAKIpJBmDZGYIY2I2ZK8JF9usmRmnK+xy3QL
MFwfskKq3x3NE76VI78B0JrKzdNzIGcmBd/iztByfS8ePCq0O/W6XZwReG39NfaW
0lfCcnCJ4u3FubCsirxByw8A0memJeutE31OWcBlRdAbMmX+dgD3fYkDA16uZ1Ju
LmTMiFKPkQ7UJDH08mkqne+th2OdIjxi+LbR+x7sM+R2k0NXcE8CN8+nBBgMbI7F
yW4RhjluIRnszZnQmbKqIzdGp/2goNcq1TRgJxjTo9fAPBdTvftDUhIRUnatJpfK
uVIMtU8seN+pXWQgx3Vsv8DyV8C3CR5yD1qPhQQ8jR/LoaC+jKVVAV7siDg1DoCX
q/7Vz1l+W0NM67NPGJm/dgXsCl8RjXgKZivJniZYHTekj4sHXEJuSBZoY18fWfIu
66IfuZethIvco46v1hTalZRFxRIKs/jDqcPdK0Atpi5YaFF8prIpRY+whU3RyJ1w
gliKX1YDd9II8eqiwzpS1NpVOwHATgOZIW2xLk68AKLL4kLhebgosUC/wtM5RDDz
IggWki6bP76GbN11X4p1e/5wC/7bWSLmqQaC1L+ygzUJbF+U4RhP9dLEX2Kjqm9C
NXHnXkHlAu31B7ht4VuKXOebKcbwnhLKRfn3ODncwF8LZ0gkA2cOGde79rv44dJe
OiwZAzW9mAKC9NCPJ8gkA1Wen874JNBkUeHoPP/HtPMTeC2X/1zbiJWQUJtoM8MY
2co5JuP6Wx17AeBtggGKg2K0sSZRxisX54SFxFXGN8e7lY5J/QzEJCHjAww+ABFs
Lv2B/ifo/uS+fR2Z9UAK6Cc8ey9Kb352aVqG3/EMj5mdFY4VUlWYGayONZMX1Baf
EKIDlRmlL5+GCqs7T0IdeZ/9BWwQy9np1x15Xl2XO2H0kwR+XaYOfvuMvKTFmKEn
rAOjbqeu0VSune95bBIocHi3Dx9ywn3w5l5I7SFGbs+bWtStC1P419kdKytUF5wC
dEEnOBqqnTr621u445tkG+q0t540QoLo8HLbmS9cUYzOeicbzeWxCZSPBUjvWsFt
9aF7DC9tou2MFSSXzys8evvS982fH21I2hIWhWHzTsfCtz+qlLT+0QjoykjB+7BI
jYWi5doxgcSxHiTZs6u8UDfQ/0uggCQcMROz4JgcCyFY8oBke7VLraM3IzL8ovMa
fRpUJ4acZH4Lq76rs+vppYkGvaRIvr2up/Ndw4RhJnrskjhyjjWYF/Zp3BMbBy8U
3nqAFgR3WNJU2/tXr8Q49nV0OY6ywWeEIyr1yl1unTcH+WYgp7SgIPXFWZjI9Wng
7lHWGoXqVo7a7JAZ9BdY1k1JBMGUI525F+GBmUKoPk1wTtL5EW3acMFeX8i6Opmb
gx5TmpruCvLch93Um0zROQ2VH8Od3DhnlLGHdcepC3mPsd+u1zzzP1Vzd5RN/15B
v1gsEE0nkK/5YvFhK2FnyIDBwHyzMBE+vRdNzSNZC/tKOwemoXyMDHAE304eD2Fn
I12O9Nno6NjrAagtY/TAcYtiR9Re1dq7GXNdWRpJ7504uftgSWTZaFJ/4rZzfEuD
4VlrqtopngQZ/DL9DwjOHxgcDAoDjy4TqQtTH9xq1jD41R7vvY7Mz4J8vCJYd2wn
EpIahbzxFuXc3DZ6aGaXtXl/RGXgciMlIY/3O8pQ95D8hZjY2I4+i5ONfq5joE/Q
Eg68FD5L4CqjiaGJraTaPRgplpES7TGe4YcKhVopnqWljmgZ3msV41gIQj2/YGj0
+++z15mBUuEdVQQ5OWIOpxlrewJ52ZrqDnzQTCDxXmG6LyXslWrFKLTbpXw3XoFp
upQeWjh8CjVRK4QZruMK+8YV6FrNE7J4Y6jKJRaEiDlK8lJ8YHD4hbboUrszy+dA
k+ww0egKoYEnMrhd/WFSCgPh39E5vaIINDVMGa5aATLV4x9gSGW6Amjrr50lD4F+
UiAW2DLpGvV7rceE1yYlOROeNcpIyZExowFuycrlWmZY0GH9Kylqh6anwRauHGI6
0Ojv+4c5Qm9kATeqYVVMewaXUuowijeVlUhdTPtyvXzLg/BkHfWvtYu+kyGbGDV8
hyqDjqEU9ojZ+fIsLVKP9hgl+uaKvIp2QCB4M6kbdN5O51cKEF9usWvYES2VzjIq
TrodJBgguavf9MrlH0tIOVI9TTrFEmMk8KSHzFbrGA4o2x0mgLh4IyqK59Arx74k
fd4ghKwVCIJ/Zglw9p0m3K97UjNeSpuvRlVG9Hi5TqQ=
`protect END_PROTECTED
