`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kt61VANxVxsVhN1+aIpN2bmEIXPjVwq8p7fYtem5YKOyPJlCzDwu8nOPPk0FPfRJ
O/mcio3AJCJHA35lXPaAe6jHbLVXUBMZJEeOl8EdBsJ07n0SdwooJostBRTlHjYV
7SU8N8MQ4rurqvnY122f2Hj1flaACni+5HdeiXtCM9KLIdF2RwRqJ/QJPnI7ItWA
1S+psqXooep9ijkY/B605UDrjFb94oDZ0y6O0w3+VKuMp8nJ/tcNb0VD7QkREECh
lXkBmoz9kpXgcDEYzndazaMCupnINbrSjowBr6Bg+hw17hAovMOE0GztnKh2vrvt
hcjTQRk//Z1Vg60eFgyfjb4/JnyC9/R9/2pGpfGuZn+8Km4r8chLTESTxwwzFn+i
fNLc487tMyCMr2qKgT70HOGfslCfJypsSio0vK0geKg02p/MkxUvc4OvHONjsOB4
npk1SHkrwPywn8tE49VaYqKapkarRvkFywnXLnFxrQLSNYENp8imoKDcGKQhg/r+
KZryla3BAphnjnso6fgUj1IX8SZKMi3dwT5e86Cu5j0SJBzUJdZ6ft2ErvGFnPBV
nj+NU+f7JEqK+UdykR4EKod9azlzO1NK5EeB/z2FR5ZdxsKZoL61THkRTWE+Hd0s
gUp6wQdr/YYLBOGs8vGMTzwxYTSOVW3xpiioE6FtKNkIE7+3gSoh0k9wH+oGJeOe
bX+SqcxiTTPS6uZl+F5sxmOO9O9KCPp+rO3vsgJPHNHAvfapN4FrenXy6M6CLvg7
tlqK+NPVzys7t/LCdb1bhXxiq7+gNLuVtg008qnc6znyBD9QrXrQtRvHRu1+gszN
v9pX6OkqC7G9hU/mM1K0Hlov/I0OGtTlf0CGMMFRZQQJApIDLjToa22xnUVwdhxJ
oqN0BzPNH7GiEjLZC+tDb5b/9ROn4N/wxL9FbM4fIkNTWflXR/eCVFKkanYufAz+
HYnhQDcEjt/C9WeEde1jAVn+eLMIBMgo2WpM4JRxjFuAEK8kgaN9Dpp8/fDDum0s
zrH6K4eQp+sVQTFC+WL/hWrwQATEJZ6nZPCkzivnuPl4RTahuYF8QbmM9lCxtHSP
WXpAeqOz4hpCXOAGxJ8xlANBtUjNh3F3tuFeE8sopVLcc+CFSbAHZqIxDKrBRgy5
P10/4uo6KEY5jTbB/oV/WXmQXDJ91sUyTJKWSK6MSlWpbfDOuEKTWQIY8CV35hSq
EF+5LmJ3CYY88m2cRoUuUr2yOrbzzdBrBukcPSVVoA0P6s0FRH81V7T2i+l3R3NA
a4abHE5AsVBMIH2fxwGCg/fFrNDI7Zf6+ebZ7U0q2qmarjKHR8PGuxAHDwg/RN3/
oxLaYYJ0Hlf1phcqw0SFK4582/m3DQpg+1E0Ip1TIiFMEvwi4M/fyy8q/o1sjmHf
zA6PwGGqfb2AxjKvu6hajUyF2MTODmbf/30s181zQklaqi/0Qok/VaWVmvfjE0+i
MjPFaWwg9Uo41ZAkANEDmqMcodp9+VXBQqhJll+yIxgoFtDNe93UB3mBeHBEoMom
GtEo0T+yncDrpVHZMn8wd/QKl78bvUjXuXpowi8a2c0sLc4eGLKCCu11lu7rmvhv
R0VHImna+YSSyZ/eRCbKWiTsug0UgFf8l/spFJJZRmWj24oowM76EW42MOauH2wD
YmCloVJpULVbd3+X55QiWKcBgXLNI/on4chRCxtrDi07/U8aSga/Yy5RnpPubj1s
psS5an13jrOi1ISqtlwh7BMOJyTG+dIHjl2jxzIGaD4FK4SOOZwM6dbBe4bWuvWB
aGkLllfdOQ1II01LyIg9xA==
`protect END_PROTECTED
