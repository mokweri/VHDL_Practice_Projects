`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBTxnbucw9yFnI087aaPWrCWJB55RjUI/nxjOi7dHf+/fyJYv6T6SWgB0MdP2SgA
STNRisF/sjX41OWaf+PbbegzupQ8Po/JeRCe1nPsMYHZiEeUG4Qi2mkPev05domJ
QjLRn+WffFZSwFo78tWpFSBEuv5yYSFgfsOZfbJEoR61ieSEzSmRBbKgX8z9Dhj+
76z3USr6tDRSsV3Jz52X91f8nVlZihTl/XNRCXaalCfbVx138Sswr4fUFhpBkbVF
00yQ7pL+N/4JIBBKAmmQQPDGNAjIfWEjzf+jNwGV7/BskmZ7c+oTEoL1FYf0cvaB
1DY5TEEBnrTvJrc+ow/uoUe5qB8gS1PysH7tT/jgCTueJnVzXs/UVoHLuW1wQlBd
Sn68JoOCuDt+ZRpDpLioUq1jOrW4Tx7QSji8AaBtlMOFbM8PqT6SahCxO2ks449g
ozmI2I7ubpCqXhPPYXLeQG9TrVCLzL/LenqtJjJ2S4zKHcOdkeyd+APGKjbZbYkL
GxeZgTHxMzOnRHYR5hhQxmsezH43no49asVEZLhCnflyqUCaG7TGYdIMtrolI08z
rxW10/0akWEsOoYWGN2fxNCee6+f3Eb+ZJ0aZnSWqLRk7bGliLU6JDRpGpDzzasv
3DyDKeh1m40xA0J0qpVf3OZgfAR/N7mKf3z0ZNzc4xFdmAlWgZU2b8VCct7gjLoX
f7JEsZTJlHQpROVVXeIaGcTAOw3CGMU6x03kb8vY9Av5No7Eb7Q7aPOhbd859GJ2
nmeZ/whuudSBvD/UOCblSI/pR1POX6Pl7endI1j6jR+G4SuHiH1h+tQzsPeVrfVb
zArRYh6ERtL1pOMVZL4EPajai4sT+GAenueCXW4IEDLpd+7QMe/VU2RCRLBs/aDz
S+oEcq+21P5sF1oRj9eSVtXYUFPTZ5ouItfbAlpfXoTqUEN+e11WeUu2GxK4TNql
`protect END_PROTECTED
