`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yc2eJd7xjQm8/7AeDTjtZKar7ok3gJJAanFRC/pZ9Qyz5abDIPWy/htWUzyg94r7
rJeI5FEKMIVsFYo8TUYFtwmbHsEaIEu2X0GMbBGhZsdVIr9m4dFvSUvRxDESI9+3
2+qxp4OxthLGxoevpjyZYZrWYUqCDCDZZbo8a9RW9SblZ9FvA3/ZTylIVuWBjlf6
qlmSSYWIgJxY2PEKzzUft45GXQwfIZ7nO9AjUu0m4ROlYVUUXOPoG89G6ZljPO1T
9LoCIn2IqF/qOg3+7DnXDsFvwTMGH+Vj0XEHvX/FfAfjb50rz3UHDoWIa/1YFFJh
6ofvyBH3NXOVrgDz87UUDEPIOYMzaJ6Mt8NF2A8QKBF1ZwP0GCl8DLAV2JUUnHxh
kR4++zfynxLt9+6rdHHGBp9ZVxA6ntQhj7vMLozoyWKjP9VB5WUpFXhDlTUHTdSM
lclPrLjQ+1hdWQkY4Tpw4G1a2SgiML1EEOpS9xXGstmoz+XS8wBF9wtwdT1x3qnm
dTZuR3PZyHsLzlhT0qbkLZ8SRXZujQefFWrKJ4V4E54=
`protect END_PROTECTED
