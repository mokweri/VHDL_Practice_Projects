`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QUwW2OprKH2TWaMDF7icsh2U0NZ1c+FwPkk3Rliq9gdDqJlzT8KzQLzQKSyI5PR+
mqfYbONaJ0YXscDYqy+7uVEQsOYY+4aS99EuIdX6uIEqxBF3GTOSTISVekflrwzd
9rQrL/8QshYBwgNJmO08KwSQR/A5ZQaJgBEoPk3xeLeQypKl/98sj6fKPBpso4PW
Z58szaoVJ6CFl333NfjXQCLShhRUkr5+nCtGi4rGistV5fu4K6HhepBQBEwxv0+4
TodhaX+OaE66Z8dbUdGfTl44JYOycescGxhovYoWIWeUDNfcxdWsI0zUAj8GJ/w1
yOrf3m8SYcVDBgEFjuLb2ZPxMCQQgXBjfU6xTmx0wOYEzdbdtHtZpIkBQOXbZAQs
NrUsXr4CW2DUfBZYN4Nx6Ut8BJafBi8BtWAiS7BzN8WofRpRGoB6IMNysjbxMnkj
qkpWfFxAxxLIMgKr0VfA/LcZUjnvjuROeqkutfB/uJHPR97DBut05YYzJdHvy1D7
a6uI3OkjtXVzqexpkdFuMUonTTy498YijwcKSxGk0bjdbz9GxcsP70gevbXvXNxK
Ud7FvzrvKKnW40XSi+JF/dkG/4S2LUEzc7LzESL8p9pBBqe2V+CoNId0GGl9Sa8X
7xqvgtGgZYxSFiv6iIhp/4TgknctL4i6r1Fcgs1BuTDNzpTEzMeI3+5arHPJuy0h
B2wEtrdd1kGIlRSi45t+NgzE9DYvIB7BckdaVSS+1XDAAf9NWXwmLulbMKMgyktV
9yBjUG9nqSUgpHjvNT4KCgtU2YJecvE7fptHnA3s3ZR3oyEYFxVdD5eDnUHpNK3W
lcLekr559k2fzLS7PNzG4wyv7RRwR7ahYW+UwjZKzEsU7Q2Nzo5ISSU9FCn6DM6I
`protect END_PROTECTED
