`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6MzBTaRbpmYoZ7crULAZOyKTOW9x+iXQedR/MXud5Z6glPFaArKWDE7zYzIaEty7
w3RiH1aTwRZ7jTHW/WBMeF72EE3F0uJAIC24Rw06LSHNiN6kfBjklJsaQG3SDQdG
t+9zGAkHAlH1N8M+P2WcFObpFfpN7eKm4u15XPpAPp19Nz3Ug8TUeM+WZP0VC6zb
pddGJeq4KbSlJ4S6MXLTQDEMp8Dyt9o6SgWfpip5gekuAs//jwndwiQqwNB1tNtA
EspefDuwJBjldeTIpgeQMUfgQUYX6TvYhAy6sMQD+Q6w3RmPytSJZo6xWxFditbf
9agq4wNrhqKUumtHpZ3czaocVN7YHgbQnMeXw9i5PeV2ojviypP3prlleDjTclKS
qTuuDuOitpqVXsA/wOVRby6etWvk34BSgp83VJ+n4gdcKwFWy3AJbnHdbCUpi6BL
JQ6xShaYbfGcDKLxIV+nC+dDnvK+rEGeh4eZyxB55WjlHLrowK90mk7iy1jJtZio
iFYe8hfWg7/sqD2MMZuhNx10+e/NpzXWTljeVPnVOVs2wdzZpeEgxzN+cVLBslYp
hD5N+wQWPQ83Qh+3v0JJcxfwP55ZXKjxG4nHfWTJ5jN1wFjKTQRFi1uMIET5hUea
AfU+uzLs6rtjgWVP47NsehpPlym6hcRTjhs9u3OPjasvpQzBcFkNoFJRndxwFUNx
OlY2MmHOCXKjrdTwWC7FioZZfrRqkDPRUe0mJkFxDO0ZkyuvYIsdQ6BaeBw4kCDl
PLtcTptVBo05ihuVEcFYCx3TXruxus/sDn3RrwFDgLJzDJ07P4pwjuWejD0a8nY/
65PTAvk+wip60XXosWbZVA==
`protect END_PROTECTED
