`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RZ3qkZMnaQRAGFZr3FA6Io01+ExbZeteF+tvJztQd8fcR0azltuWmvS0nWpZP2A
0GRUEt62l6XTz3cQCZohO0JFVdlzYl5sWiy/Jz4EMC5AxNbedKQT1cxP2//4SZ8t
pxNv2/jLQmL8PmD/2KoRLat1ZjyLfOY0Pj1o0Pp5OfIYSQpBJSYxgFxwGtsEA1Bs
`protect END_PROTECTED
