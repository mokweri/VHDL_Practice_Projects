`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pstMNwhNEHwZEBAvUgkJ1u7vsIaoEFTlC/++lD8QPE5dttqqsQFe0E5nsF95qW3F
nfiuv75rxAkrS6U9esb+TdypAqe50L0FueDR7ZuaCmbcuRa2CeDGZ/3fEej9HbM6
oD8AJdA1uaNz44LCKaJo+xaHQtT78talnte16moAN0vwm++VU7CrPM4bYFDFUKdT
BfAqJ+J2W0MKyIj/xmeGWLbrMCSjYXnGLWY6u5i80tQlIH1mzQ3S2ECDrwBd0r+i
by8tTU+qXbdKP7Mlx651i2EOMWVh+enLh5mGu2f/icJTe3X/ET3Orknnj5AY9+Ml
zFGPFe4ToNDP0f19vlO1skcJade1VEepARTMF3tBZCZNrLoVvQ+Xsgg0aDDGgozy
Kxqv35Ro6Y66Mv1vkS3WtbZILZsoPlO4RYJYuKC1/HvPc9YfPcnQjZ+ArsuB6g2b
G/WlQ70vP3t5PjvDJGAvLBHePO7ZeuX0/oJrZA2uZKAfFtqp6kUWCbcSiNrcRfQp
XnVm1EIzHUPN+Q+b1eh3jKb5vhGsHSo2IacWrSssCwUjLj/mp28bNzSX2dPrKK+C
B1IrnVD+7dmHOtbxHci8nXBjRL1mFA2CijniQ2n3RqBOBJbhAZgoZhK3x+INsAqy
PLEbWO2r8T1Btgc5AWpLoB60whpWIPEHjiN/VEKkGpVCQ3SyqGwBWckALpg7ew22
5rVQUavW2TOtHHGRzDO0rhobJCU/3wIqqjY3VjRspgBBZCAk9tnT7CAwmVUzqQG/
HLpOuU5q5FqX9HlmXor0a6XItyn9uIi2gNuvm3ZMgup4HRN1D+2RVbDvZyct/2v9
TFX4pXE0D+iJW8cXultOTkKPOJwyhtfE4an9O5QvgUdYFR1bgziC5UxkTHzL6PFd
jNk//1Q4yrpgGlV+lppovs8F3IL9xP0W7PfWeZx3aK1JFO4FE5OKaB13+DvrEpun
roDCQqRDl05GUjD2iW5aIZvzK1iiVd3yR9qZsRhsBcrn+hdySHlIjTZo/xeDxkLX
Rsl+JbCi71rM43t2FL4m84up52iltDDHqlJ4Dq5mRdBP72sg7mPRU9nONBnQyBzK
ch1gfyzs10/nFYMvBJCAIG1wp5QgHFdnR/gNspVJv67rCCHkLy6VNs/Ex41nrhgC
yP0EFp2xjivdyE1iJcKx1+HHqocXjEl7tCmqLfE0a90boYWXRQSwQPlVE148l84Q
wP6ec5/zE7O5lCBhPIeo3aOyAOE3Y0i9CXG35IsuWvtDr/Htb5s5nOJaeu3/LZnU
DCDQKLcGIiMP82CIPI0qaDyO0Hl3S4Ar8nVOKPBfWZ3oot2fqTYQ4y5cFK35P8ZQ
bmH39BpRwcrW91YgASC5Rlz3x/cB+jzLrT/Dg2VfwmVmEW9vcdADBhoMpS+v3Wxo
zz7CjLCH2LMG83CKf5Q/jMWLuiy5F2f27dJ62P8zraKEvNsQ9XFqLcuvK14rS0wZ
xm+SZkbbROMNZ06t79bPFaXjpA3kReOJMvMPOSBdQWTV8vPygHinF+tkqNiGHVXo
Cv/5yfLiTSoidnSv6XaUOwT/0NkfOPWdnTdruzEgm38Rw0Z1m9EQXz/GMKnVhvH6
/63bvL5VJHt3jSoEMX9DxB87TQLo5ZGq1BvbZsxyZ7uxWUmVFjHI+GDRg5/5aBsT
RFGdO5whf5jKBPP+Y97RTqv/wGL+zSfJqtoEZG+na20sfV84pioOs+R8GNsoDRHw
l/kD1wYNTLUWv82lI8DPm9LMgzy1y0qa0XBEUFPTeXYDRJ2/PZ6QLprFd7mvzrPH
wycwT90i25/YV9kdF+EKhHrxO6VLG7qf47KW2+RT1I5Hss6CiHZAqnjsphQuBiBD
vxkRuLhczmYF7ctwZgxDqWJu1g2tNjqJB1hQtOk+IOBKY4SPtAEg0/JqPvUZKS25
1Ehjwj0F/TDFhuU7FfRISxJt0JDtjrG35tynvVN5xaA1cbpE+Bu2l32ph4Em4u8R
MJL2V8ENPHvcQHROadRkb8m/fqQ0cd4p8NxThqA3ABCY242TA0nq9DT4nQzvw57b
CoQyPKg7glONc9jl+CmMht6VSOjy3wyjUZ0eePqviq/7dpHXfWY4YJPm//eHUdUi
+yonbw2LlpyRdtNBiewO7iNqQYW4WBDgX57qDXg26+r2wWVmliXOxJ74iwTJDq27
Wp15vQGHXb0bw/JAry8YyvqMOfKtkIc5Rp0lts9znxeJ9YLmElw7eZMEOUJv23MO
rXbfGM+/1IPm2BJRFlzqpkOWa6MbJe3e7nKs+ghtaBwzFWM2CetxWNlDg4VGV6WX
+2E+0F7PoLWyUhrAIn1toosAqNVzGNAk8PA14qoZmyyar4nwo9B5d7f6p28S5Pny
HK1U8ajZrsV5GdYc7m9W6cPMZhdRoBD09tmO2rJIeUHTZzlr2GiA5aEVUFcqzTuq
3MF2Gu71DJAswJUU6kUNSIfgdFXdlzCtngM+7Ej/Xzf0jo7KRlHBqIHd40iTKlYV
M/C2gSXZ8qR9mcTMyz7qnfDUlsjOpxF3sE1xwBddVRn+VUqTGG9o3njlkwor0XJO
jNa87g+tdJ7APXisxHnui2UWjcIaW8jEumIaZZBkaHMthDqmSjW5LoMgKvd2zl8X
PD6BSmAAA6aKM0LyJoICdOMAA922b374v9F57IJqQbM2W2ul0DQKs3JM0AJaSpEG
YM2b75w4GYK+/P/adabRMicDF9ft/ptV5M0m7PYeY/jFizObekMHzzWjCe/rwGKG
CQsGZ/zDKwfM1IPOraBaBFGjE4A6HNg1hYvD7vL52Qd9UJURzBMYUFtlB06AcHzl
p+dtkPjhf+LrEGZAM7/M7I3NoP+liOVdwxCSsCzRqo9SKoSNWGr1vxeNT/Ozw/Kp
pVeWvgL6L4kKdBfWEiWmeKt13qCO2tqGUYQZBWWmpCidgOWV1jDbx2G3MEiwr5/Q
DsHoaDZnVcfSTwHsZ74zGgHAmE9k7d7FlT++ugvQ0pb3vjuOcYLoRX8s5LF+E/Uz
2vSH99LVM6+x5rcY1nvfo+Jgmja41j11KeJaZ3Wyctb/fc1HkZghvWXlGasfAiGu
pKAdPmbg/loU86njkAN+qUiwdNShB7ONPcdoGh/ZoISLAuULyQnYurI8sXhlqogP
UY82qPp6txIq5y4WDcV2OA3tz0qyN8UF++w1olepPWeKX9ufhmQ3RWYjEQ4MmSe4
ryEKM/au1saDgTScqeaYu+lAnLm6EgWvQpG50Hr5UqDr5TETcqP8N6F5br6Kzf6V
S6BLeY4gK+wYlRfaNusMNidyfFTVTctbZe9JY0LiZRaM7HRG6VkoAnJvvjJIvGFv
nDLptYZbeNxrFBgn+hacSrQQJD4DaS2UPrKOaCY5ZJgdFj6nBTRlH1cLNLt8492l
BdW4+Wx2PywvZw+PnBLxDr3Jb0eHFR3eoN0O3ZBUErAZnai/BBczKfVA3dU17QXT
0/iknqrL9GB3b3qE42m8mXEPVpo3fmzjCu6TKcK/X+CG3AiYK92AzrpBAr/g4sjS
Ger8JlTKgpyVsMyWVEEks0HzRSUkxe8iyvu2qxHmhtgcX2gn2uemNguT4uKOoKnZ
sKYzOrZb3Ck+PIpdIW0VXhmMBYVicmCvH9orDnxWUjXxsMsafeUPS/Lb0jPcc//y
w1VVuBinJ8fgo5oBZdxbb7oHWUE8xiKgdDDeK93DIGBFNpvsATdMnvW6WXv/S0hO
vicSzimcQiR2flEpe96mzmz27n2J0xC/zUIxYM4STKqp8m3/M/LXubYvnio+K2ey
MVG1DloprXTQuQQURf6DDpRMRk5fVUWbhI20xCG0xVtB2G+9Oy4oTJvdirqR4346
SxldIoJlDZia5qef/61V8kPvNVB7fe2AliMZxcMq0XzwvNJ1bbYWFV2948LA3N8r
i2KF7D1xARBhWMfhfmYLII9Q3JkQOhl/ZSkUqj46BwiPlUONZ9Piq499QpEo7/aX
YQRLBF18UpGPTDULavK+TS2LP9TFN3H23CZfbadc7x1LEI/W80VuR2lzr1/25+Mm
kcm8mZARGz3gLRCplzfuJ9rQx/xsZ/KI3zBq2YIPH+ywvN1+zaYX3xVchItY7vje
lus1MbjyBo1LXJbajoqk6FoCZJDtWlemfmBNCzeJeBFNxoJfhUnAfPE3HgqknLN8
gtcHqDkErCIkCmew2bz2CTWdBcgIeqk7Vs2iLDwyFcGOn0DhrDCWQYY+qZ3uYlXR
UcZiZE/bMzlIxIjCKo8FyUsF3zojZsR5EnnbJmQj2+vd1ol/LkgygOcpJV27BB27
VstpYMqkbsa0X34vkhQsyAsWrs/NiHukucQKTzq1HwVCfDo99CZ/lu7NUuE9FDxu
pCWEbrmImNuCaSpgBeDJIkMehGn2mu911m/Q5u6zY+rB4r6nMt6oXfXoc1+q1E9d
Nm5+X9JMFNFiaTBuFyg/O0lZqo+FjxKcw89tc6CTRS5aekL9AjcqFRKLs9WIPimI
PEdvJmNrQBfg2Z3daJicXekvsx3SnFWcvrF4ZUILYT3WKGzlRxi0rP+FJSloLWiB
LFzjNw4YPQkHckwZTpV1lDH0hOIUmOhX03oW20V9ToJ/Ty2UDKl0Wt77/RR6r0HH
3T+9Jjx5r7sgJkL1I2iq4JPuB0WrbKKfcNBf7E2IbghDB2qEj8pbx6KnqCGTHGda
QNqTHS1HMUd+X8EaD7nN6XZpLuKXaeWpgvFegrWfZrIP7rSohaiz+GYahqgwZsOm
SUxXCbCaxzhog1IFmytXGeC7rEpCBKn4uAUkqPXN3nk2c0HzCFDn5mwmUx9u+pLx
Q7J/DN+xGJjagDXrSHbLdMTEa0MIRy5nS0bzSV+yRgzw4NDlqIVXuLcP3lqPUR29
A66Xvz+yE8rd/eHuv6pCCZ0jUGI1gDfUYBqJKmi3G3T1Dymud/bwvvV8iZpSiXCL
/bxWHaqfq6nlLmjgylurHeungdqABZ03XCO4GhB/3lYRH6KvegUCDFeNK2UECYlk
dHhhvrslTHm8Vj3LhDCdWX5sgYKa5x+uzdXyXqhZ6lC6K1ilZDrlNda0VXCZL8y6
P7NLeWzTJ2EBwy5xdKR2aghB5SplAj4q5nvksRsCutdpevdGa5GhTwzwYS7Gfdrs
6t5whO8pdjhI1SpWpLHH9XD6LGc4lUovgjalQ76JCg00wbQAtD8V5L/Czr53pR+E
iSXZXmZfdPU93V6AhgeLSzKsLCDutPrBdopjGA0G5z3wCllMpldHFbUUi/KwHfp4
s5cXaAgs2jyNqGoz6rOifqEr32M5R1+aFan1kFBZLmqXMK6fK/dIDl2OoqK58kbp
VhaVgC40Z3z7rdOoZt+YDwByn9Fk8lONJo0t/p/Nl8a1KSPFIRKevcAxxoirm4g3
IP/eigZqUgUEu0WHK8KcJNuba6SDHKDCJ+77M5049vshvoySnoSXbREqTLHxcwDH
fEsMQvzMi2c+4ICWTY04ujDkaX2+XUL1QeBYuQnfnZnspJ2wHPdJtX8YOHKkUsDv
CzUP+0Fj9qPFbPRCupBVtARdDJKUTH6q3mpN+mzhLONLGE4z1vBnVyZNJhXmIlA0
W5HPNjKCEGatcxlvPhpJNXeQ7sGNayjbB3MC2tYDJ9n7RP6d8JxCvzSpc80NFleR
AoWfJF7RfJK6oMCdzYLza9w6VVvvuPIHEsorJi8EhxBY9GfFrWOOhyVxormPF+Rq
3ap5qd4rkuivc2iYspD6oC22f8s1kuc/k/qyl6Vweh3mxsyQ03b2omsXHYGx5q3f
IPBFWrrJM+19WR7c9lhFXeSrhH2wcgd4VwcfKjQOfP98Smce2c/4uVEUqJMgQ1G7
d0OY17PGKuwL3nr/Gth0WPQ/KFLR1vsvrUmL43ga2aUqM36uN0RAf/mhxqDYvDh6
jDECGj9nlffG77byeH/93FMNnZgqLYjbyr1Mt7ntTtx8Av5zpcF7gLxyO2erZ96l
o/qzOc1NLz6uhIL8f/7LJ0YjHnTrN5/bfjfseUKBw/YtVeSOBw94DK/bJ9dL75fk
eVFDf2a4uDlRMekPSYvQB6VIhn7T4gB5+FPWYe4k0dGLvGoEfz1Fvw2ydmKqjI0D
6WoaU79zgUusSRc+eozsUwDHKccaXBLzLIqX/iOovFzFj7G7hTc6D4yFqgCbdWGP
eCHgiImBZgCJf4JbHe6ujOb+/oqwSDkJVrqH/oLm1luG3bYo0nEH5tJtT4msVVnA
y2VZ3ccqsKsSqV0e9oi8RvkhyqPCTpvJ8EGPzm/eYT/fcVhfIFESN62o19Sdx7lI
0CbsKneqnCfpbDvleK5OPs1bab/kOs6tWjlrFRhTnDhLlxS/Sg7S/vA3ssLVL53Y
VuEufVda9kZFXGIbfpAO6eLM80AJ5noBbhwD06ry3SnJE2Lj0SkoTH/241ujwB1k
cdNdVKMvpXjt79UIlnQdaEl15PLhptjhnOHr9KHLBeco/7LFthu78wVGez7K7KZJ
k3tXnkvXxzDQDu8N70RE0JsI5yomD7kUSgS8f13S+mA+HqMgxsdv9UMfzLgeFDws
Grq3jp/lwtvHYmBsPptSseetILo1ehz1xzh8WGCWXwpK/jpu4NZ5pXrZ/kc+C7Dt
kMv29zrdUjiVMgrTrEXAMhxEQA0ylp2SQ5H8x3EkF4DFczekA7tKrRq5vf3sQ/5Q
MiADsQeiXvfJdl7KyADQTeypOaWp0rw4Zx5ejycSXC86bt27YuDrDFVqFRZYy9Bw
6QXDdKjuBjJOtdsDbD+ZWJR0rIbl1uWMRrNwCUH2ItC/YWj9png22FCPqLxRW/JT
viJ7WWB+YlkhyriC4Qil5NQRENRmzhqFjhZ5f47P7FNkOlDUBJczpCrpAicv1aMd
ILZMixtfYnoVR2lgVbZ8KJ5yh3kxO5Vu7RUr3jq8RW7s09cQNt35IJ6uW83AZyXz
KF2wBAZHaeUjegu8HwVr+BPFm2FsybcJzxSxyxIIdjmFldw1qOpitqok6VlMwDB0
tg+NEjzQIRMZtj4VQGqFcNU4WMIYKJW/xM88RmKG//h+d8ePEbSSd/2SO8qXaRSx
mqpL000iFGHBbaLhu6tvFkbpUWD60TRwkyIu1UuhG1jJg9Xkpl0fSdFxI1ooSccQ
ddH4Pgk13YQYKEkioMZRpDVOlbFrdwdVOuaRa7wLbRkGrLUq4cQvfx9kvf5+eMgB
hzmHFiZnxy7gPkCyEmX75U+IkHdPkqe2E5H3b3G1+fXC86KpnuBEOS36zeNDiNHs
AJf2ioP3kAheDrKF2A7iK3C5SzZtNFIGr5yOZ06Vq9Iq/TH+6xZ2lPg0TBWVYw5D
aO/S9Oz75qJjFITv//SiA3YuOCIQorFSMXTd3HT+7i3Pm5gHSLCo1dq84NUjGdFC
qo+q4NTMT7x5Y/amxyc8eaaXtDUeoE/nzPq2Co6kYpEBTwbGtvzN27nZAMIE8Pa4
3pIj13YJ2Jk/eDZVEaI0IeR1RlBKZDPvDuidRwXmMb8HG4ZkCI7T81C81SmAVt0y
bpAGTQFkB1jRGQg+0ztOlL3Gbo+TYrjEzzGRaBIjcVvEk73b+IdqPJQqPEpYe9Pj
E0Wov5X+GTQxwOAcykAsOT3CX0mmIAMaLPosJYLjT4XBrBS4lDe1NeSqY9ZmJlwg
fDZCiFAv98MHfSB8Kt5gRMEL5fet5rifJ2FyPhu12tUV3aA5SonzZimBd6wTZGTB
jg87RA7aaG9aLrgkD5g5wohgbMAN/o3+BBGVk0V4P62y8+tpkApuhZcM47l8zrp9
nav4Hr5efRKVWzlipUNcm0fDBu4UD8GW77OVBPAEuM3imd9GEMtZa4w5qslXeAVd
n1ojPPc9t4I6nuSpo1s1SU0LiH1R4pD0F/QlqCQxFdqlPCBvL5uLRZUA1K3h2Asp
k2RjwCYciFMKDvfQi1RIJPVAV6+nHTplNctX4vXf6mSulbcS7p2m5qDicGmrdTTu
vfGJCnQ40rAb8EICqB5mP64JvkRQ24OQ8V76Wu/+eYKEDfUJ/RgSNGmdot9Px1qd
Pux5Ifb0rbPJKFi9HAfeCfWH71/vxCRmNWkmBZlihZDJmrvQ2shQId3cGoDj+iqr
xncYK0a/ZI/VbmM39L3JXZ8XwPxkjM4fPUxf+o1SlGbeq8yfejkodOkdOdQh36lP
zM38V23XpmpNuGPNrrdCBDjUjzbGIVjEPjYw+gu6fx1hVfgi93lhGTUXqiOe/e54
9YuUAypxHBahDtE+3F4HZ3G8Cj3u/5pvP+lZh1Y9BfRmsxRxjZhgvrqdx6vX1nAw
ylZd2G1xVKSVfFsxkDtydO5xC/weZGHnnnCiBy5acVvhCS/DDBWbTNmoj1lWFLAA
UoWNxzkhHERIG76SU8QFTJLLPymemVx8vMsK6dzZZMPBIOgA5eJ7PRXpt85HJi6/
MGgP2+nIKzRBlKzC1jByFOB88wNDSuSu3mOW2fPNYyqATp/jJXDOrN3k+mNjDHBi
v1jF8rdPZrNY/ywFugIyrFRIMAehv8a+MFT9cU+W9oTmLU7KFXNFd7HQy0C/urEt
c07T3gOO8IRa/HjGIQFdpA6OaP1zTQvOwpR/gVdXTtnUjIk7cqAhJvMglEy0eLH5
o9lgv8VJYlwdHAc+IL/MnR4b+pMhZ3p3n1TknbMXx79M52rh3/v/0S2cNz0EqNaO
5Mr6K0xuYOQeDdczASUsnY9gjw93x+PNcK/eBnNrzi41I+pamOw0v8DEvYar0h/T
gayIx6Zs33lUdhH+D1qVTps6WT7kwjAG6sjrfJcH0p3OB9IsWPNISn/G9EaoWc2R
aRqR5u0845tVAlqV0Pblnkhxj6UeJa+pTV006+Rqr9wAfw4afBUqUSkfd6BgyKON
tS+To1d63I3Y2FtT0HeT3GIqFJhL0Lo5ylX+1OKP2FhvATOSAFukJdJEOfh7J0qq
xoC33RUkw/+M02lcLESanZT0OTDDdczrB5LG4OWxAYOMif3BKAVEGe4lI5rQkg0n
v/mYSlHDvXQPkklS2bi6vPw8Bg0E1eDFu6QtD34BNA/FatZuhvZKYGGMkV29Pzj1
ZxMWKdjfC4cSPAoAWTOmEuCatxuHqzx+R3ZR+K0KnVxurkfx2O+3UPhW6XvyCx4m
JWaPli7Gh0RXS+yNNQi1zrKhKubYFwdD+szX7ZjLQfwW62sNM5FOsT5O46L01wlv
KD0ES6NSBXqvpIPbtTHWUMEPAirKzAhHZDbzbaQpg1f0dVrU8DFUP2OyESsekOcV
jRKUFA6RFrwt2d20wAY+FxT1dQ9o9u2EbQ7BWqVl0Ll54SHt8lXLEblDbRAxc5UR
1L27695r7aEBF/tCzO6NdQLpTr2zXuYkEi0IkWIxHkcZ12ZyAxvZKOO827Rk3eKH
wHyE8a5UbXE0LhlYShGXLAybXwhdybo/Ixwan8gtQI9tLTfXd47bJaI1RDuZcncg
mQn+ju0osEyZ1ztye6Y3GuBtJw1TG7EyKIsvgFFc3cslywOhUKi7CWnAdwbkNAAJ
YvzkJtAas17U7kSL37enoaKLOqAw7+X506cHtcIF5tVIdyVPNNVw4VCHTtRKCnu8
47JUM30Pekv5IA6/Udnsn3/kgOB2ZCVyrvJAh+9ZizPjdjAzdeogzEFS6iB2YfwC
TzR4BsBDWGp5CzqmOjK5wleJAbSQw2S+v6+XmPxpMagx6uENov/Ti7Bh7MhZfsyz
l1J/k7fhAL3GCeR72nPKf/Sla2vi8S11M2UdeCIBGGJSBFLEx78Sg8CDN4J3sZqg
wukSqFmPO4MM2beWpL8fF1vFlAehfQz0+UJQh3fW5Ls6qGT8fPVD+OL55WD6kB9H
GrFAMAeUTLXZ3rOSjAB7T8MXLFijT/TJbPOHhygtBux+EYbaAEqNiouijFYX/Icd
oivUnJyro5WlHJ2Hpet2kY+ZJw2NiVFNFdA4R00NsPSZqAs/pPY7BuHnjx9VoZ7A
AbsEqBt5BO8+2KQC/VhydBbTXVDg93q1x2gzf4j570OaK+FfngFHreoVUCnuaQJM
pI95tEeXOVZ0pmrDUyJkVnsa2oDlgX4egz16cTlk5nMwFk3sIO5w1orDGTCs+ovA
kDDIjoiWIz1iQEG2xeadUkdY5qokWIT+rjUUkuhOkcUyMUX5I0kTWlQvKdy3Av9y
HN0uzpqQXpeZK3LtOWWsB+0eWnhM9R/nnbYga2m/RKViHro/ZnLHGA6U/HrMOxXp
w4lnEMi46TmYjcAcPMGi6pgjce0kSLQpSRecTy9MxTF1JKqSR6iznqCWTnCB8RPb
vgsGcGLvU8WwmHsoFKc7bvzyEr1ugMMT2ooYg9VoDGAxfrTcJnLUAh/5Sa1kbHXT
MCjWrhr076jHZLfcHcs/vSCvbZn9MkGo94rfHRsAL9BE9z+ssvhGZIHPB/TEGIOJ
JuDyetNlzVC6Zp+pU92CuG8Nzlx8zmBwfm5gWqxjQWICPFHx/TsVjNhIoaQ0CA3N
L+tL2fjtmox8rddMsoRT3prSCGpmEiW5jCJepcs7x/qM/YkVCg+6p6eCVwZNXRNk
20PuW5meZAszHF6Lsazs2RR+9FO8KRuvDF9vLJGvRHktjqIRKSXAS5G6hq1d4p+9
NSpkf5fghzH47BrkTT3W1HPJSlIjlKqYX6csDn1w2AAhD5s2CU9SryjNE1O5LuU1
am4cjwn5Snx8bOtLPuPmCPaYaenDv+l1hSQET9MBIK9+E/IX/ezQLxMGWwHJcETr
prokbY+OaEEaS6vvRu9h2dAmOI1cSfYbb80dn2pkWBmJwVKl0FNd4o/Z6+45+1dY
1JvESOPANfTVD9JQpaPwpJptqwNwJyzxJKpGM41+lmA23WF9SzRwDGVjMxxnsVYc
WQ47Fpg+tdn9d04OGDB2+SgpSycyMcUQFDH08fq9KWS8K9VXo3GgWDP+HKhcjttu
ZJbdWxBuvV7xtJtK/qMwj3y8tCCrFSql/X/w1N8PZyMUEUJFeOWOInmF4VFfd0HQ
epX8yjnAA5VPj/6+i+3iIw62YYnrUNsSrS0Fq3KvVvHSXDDpeEtyGOKwwj0aFOEv
yoRw+u3AHcoOjIsueGkGIpCgug5QBW3oQLOYs9NpUktEZwFr7iS+VnjYIu6e1xOu
+HGThmHe34q6VVfkAA7eEw35KHTy+M/zLucNWRufApw2D21wvdIwzQLsj+XyZDik
ZtPhFNOKuUzHbDrmOPEGoBZHGFVxRhaOUX1tXduQf3q4ob/RlxsJEHdz+PKvnLCD
wXpGC8/YkEt8tvf9tvTQ3a6UOuplhJo1B8ygsiL8TSievOTG4CtjY7MI25oSQk9V
GrWMTSvHygFqSlUCLabdIkqb3E1w+pNSVG+tarOEookJCIMi+euapv+qtXjK+K3E
P0i3G23XcC5fq+R7PNLE4YAWv+7o9Y7nPdio/UED/zMSOaxN4cDf3Gntpw9wYrct
9H7TYAnublEyUmKZW2m1sFVTU0R19lJw0u3u0JeTZpQBATON14F2iOJT5qCIBswr
0i7jTuiBpUvY6bskaXagcDLVCe1FSJHMbSMfGMOBxQxXMAPAYuLfHHVgfhj+FEJp
ly+SYPDlYiK5zNGXouuOX9rZtJN/BhCOd6idS3NnrujrdHpmk4ACjs1tiuFYc+9a
vGu2e3990E0hr2RS2A7PlkRUaHx17cHb1j/Gxr28TVyiHx54P53tZwOvUYtEVncT
RxcapJYryi147XDQQr6UGgR+7vJ1pemUcSPwkKiQdvl6IqM4+fO6SUEji/M5A/AW
gQ4A3bdJBqX3CC+7kTYInALS3J0s7fVtu26wklWKxfQMGF3L5e1CNv1NT26DbI+2
XQ/c3fpKRka08f50tQ7Y3IpXhhjhcBQhS6A/WZSZug6Wh5qCabtPHF0LIzkAtjnC
E60qAFPRXm2UOKd2LzLBtzQPqj/1eX+YCtnXu9WW1EC1Hcb0aBFha0XBx5l0+uPm
eocwPLH1zRvektdO8zLYgQHw6OxyHbDoCAngaxrCqhh9XBfCFuFfLVnUdsOGahJ4
XhecTHwhm2b1hIRyHRg6Ui4xiGOyg7UT2n4KhBhcNhnQUR0VZVXnX8Q87s6Tg+3I
EQoKaWeGroQQ6eYg9SJDGFBPd3QWciLFkrdbxns1PU7SBzLvre8vgi2a/EXEMTUQ
WJBe+SQWaFasR0Pj6aJw3jysDEmOfdRsg61XWRy1k30yAMyzMNB/FSAjUcMgmVhq
wT55dOzKqNDdzjjdymWE+kKYm4sltvrtrs0PDwsaMIQZYnryRYmb7crzSnRMadFj
9oYwrVVSSiEebwAxQUQTvRB7Du02ll4/hcoSQ50vO5Jv1Lb8x9rC2uiuO5ue00fc
2MMQtGi+PcRCun7gi8mByH+xyomoW7t2c45s/K0MzOrryFRwt7D9z3mrtXtGngZo
wyOwBo2mF4e6c4k2GL5OqTq7DkjUlTg63rshuRXbyRAKPkXniDno9yv2ynZQk+NJ
/TfXqbYjkP0w4cflgbSj1blOiPBU6DN2uo+xo0FWnUnVtzW6dexzDhRMLLLwnpeI
RWO9O8wCnH8DwcJBuA48+2bD59VGTl+4Dt3w2Ne62iTNJQUCv6X2x1GPkC6OsU/3
6VqBvXk7bD+g7SwqFntA48DvFjqFEgEZyhpvPnDUr12m4BRsKMVPkC4tVl5Y8YH4
dzYuYWgRkcVXManfoxfpj9LT8gk5uaszwq7GjNU3JwzJSJaq4RR4O/t3JkcQblmf
N3vsb9K3CmYeGGWNvf+ez3BfhgBt3i9mpXCsAY1bP1XG9CCfebzZppoBD2tYcJfI
oyjhKxUoKaAytRrER09iy4zSC1cfe/L/4I/2DYKeinf7OBguenFj36ZU+Qjhz0AN
6/NN7lRHQPSaUdW4S3mXEFu2G/QRbqHiUQGivA5X3bsM8e0mpij9UwMUlFW4JCv7
fDEGpfCbqeof8pdMuEWgZxHLRxSkd9wfJxZTCAFsfzHTU5Sba/eJMS2WxMAUdCg2
5mBXbas1UsZanvoTutPxenV6B6akuhFIn7T3QX50dMDFZqOLw1HYrX5PEvdO2D93
6D5047mpZaStiR0FPdTJoCS3Aybgirf+k3XyBG73P/pVqSG69pNEKlejabvFUyY5
1vb664tc4XxVhrnhIKwnljxG1eH0CayEeOqE7TP3Kni0olrqFfAFsmMzD3VpegIX
QWdae1AxbujoOvVT1xQcVimV6d/Z5YU2sKOtwFcSKx4VE7J8+TiMc3R2LmDvQmTf
nTL02Eaa7o4IuogYCwN7u5AXYJit6jZll+qAR5h2Nzpcp3WX4eU8KGo2lp2wvcs0
l9tbsd/DhS+CAMoOX7K4oV3h4g+M62Pyd0rj133gm0pw9sewoE5qM6wgswh0HBHD
WklyKj++FaRibxDpCNjjwH8Ys9FHOoexAHZSoAf6NTgwRtmmk2rK6c99Cm87gJ6D
9ghX4IPp7SIsfxUpLKyYMfeohubg7v6syFyiJDRrT9jGyZ9NE5XYtf+7i7fJ4UDV
8JCYCWxA6l/3ZTaIZSGgFmdoCw+LyOpwWzI5JSzVG+1AGR61FnM2Gp/bkRnMOqVr
nN2onxYMrmxDjWj1Pg9XgXtOOVzNmy5AYLJ6HAiXzCG1TUz8BgzVhpGMC3bxMxJa
vdqh14nwNAj0s2radv51JVoqWxsMWQSAI/CEz/VQC75LVN3kCDCXV3PLUzjto4rx
QgoT9hk7FR3FOHebKsNJki2ZrdrTrjuj1hGxt+ptTdMZ+RRO8DjPL/hpypM6AwL9
3ZDqENbdRPZKQLui6YRtYeieRJEeKmv9NUajboYmwieK0ZZRR7omkqdqsQv4fgpi
Hdr533nQn4GqgRc42Egx/h/7v2Yg4ucML2so/i7aPzkNSuEfRlobQs7KLPPjTn3m
ScGMRfwZ9AJkJiFkZQgYh7xpydnNshFV35nKqoS4cGdfzreOBsHzNh9ZB9aa14RS
L5e1w09K9P6ifyPQanXXf3ye9m5fnCVKQfmZypUqGTzYN9N8fZzBpdKMPXu1g3el
hBcyL1/7haP/ANwJLCck4my+yzLsHveJemYfxYiclMowgPZjEUEfVY0hd5nirN2i
BenV7EutAp0TPC9NyFykRJ+yHtHdl6DUcGP+WsdjD+OEvMGsmgVRmVPfDySvKI96
urPh5oxoCD7ykJucMnWBCUngnuhdDGrysaRPYRD33mLun6Z3glcAZ5Q2+2s2CcNI
s9a5IieR5zz4TiTEJSfkCogNsPbLGl0lV1JFd1EJydAEvkLZMbbs/5dr64wo/2t5
uiW5BvGXz/NWWx7uFKgDTi6aukLOWmyHH18puEmrlVCtk9nnkVqu60smuUHxC8Gf
Rgavnul4sndw9bmPcOVKl7rAt0iixCBy6tE1pbQ6idEYaTWWvKQ4fmUdYcE8hBHG
3ID8fLeovo2becHfwA/8mwr43WcWQ00rlAK8oJdyUVohgb528Wv7pcGhXaDipQtn
mIIOvlUguaGRxi87EwYWYsPud2/L7oTAWpHI3PWJMcVcjwOFdDC75gyMO9+1WDgm
IWt4iNz5tvm33uDHA8ItWhjYGaCtfdECb3zDr35q/dNgX09b9Fdit9IKaf8qsArE
buCTyYYX9LobQipqj2LKH3GgHBH4yhgWP1NAPn3FJMDB8MjEPJye3z/7SSg32mMj
dwxsfD465J1OK3s1IRM/l8QjVnjqcUg2CsGcV7XguEvROmmqLUYHCrw68knxGJQF
zpOn1pApWdNXOmQ5/MmCPypvrNrym8J5djt4cMKksbZbRb3/7GDtS/aDPsTwli9Y
FN/U9FiyBSsVMlnGbYkL03QzGXsmaDxVAvQmfwMM1sYKx4jEe5z3zKtmxHFnMjxV
L6l97RxFkcHN6yS9U9QTKxkjQjsDVBod3R3CMxxILP6EYKbYW+v5nNdmZ+4XGhDz
2a3XjFdIZbgo887GPudnVhFz8/dEZz+mq8VnHVbjFkDuduGWVTtCcGF5ayNunbkM
f4H6NTU5d6CgU7X/3unok/YbNEMVeoLLRahqqBL7QrEXRYL7lJ7NtFN4wkGYfCAa
L8yuG39uwK/SAAwfVjtfbIi5yGxS4wiZmBnYq8Wuz2XEeziT2Q7uHIMrM8sGC1VI
vqoHP9WkjyAEMYff/oE9xIymMh0BRxxlHf1KVsVn4RnhRKp5BiHnFdfYhNtAagAH
7H8xWp1UYzMnoxF8QnVGzbL7V5vZ7ALOyfseJJRznJn3biV7OVJPUrwKCFPsEODS
o9XcYPsCmScrfk5MKkOES++7ZYYbohSya96AxT2YKuoRMVgfxYSTx5/yDLsBQZWk
8Hbl+dxBDV6Gn4BxN+PG7rvu9+JenSZw3oJql5iLj8ftKPbqepdfsChJOBk7L/Lp
EJFHM3iWUIUftVEX/D8QZaj1JvzLS2LwiGZPs6ps6pwMcSF3slynSEbwCVGLahb2
pHY08DXuP1Pw6e195sNYkf68I/tXCNdlG7yy4ZMuhfy4PJgPv2KpoAi/H8YoHXIN
xRN/nUBsR9cpdQlYOrkQ20Y20+UOvSNYJgyWZkXGkFKrZcm/mju9oqreLQF2bi7r
TJo26Q1G0x6S3paXCa57+FqaH4vhH9DIy4YicFqDs+S8oSdXOfmPF3UKZQNjs5df
AP7SzCZELbk6RyZB3Q7xwXkaDcH14DlqACqhy9sEbSD2q5DPq21j9ZMzqEYAFi/R
O/clOdUm5Ff/HJSeMCc5GrZ6YGThTMxLRORPcMAhmLJXi376hWbN+je2XZ83O5h7
bV4MIo8praZMlmrUsvfSav5Yc7Oq4o+nr7SGBnOtS0TVFJfbe5nSAiPdNo9s6DwM
oSzN0XZdoGY2THMoag6oKalxzwX+Se7x2U0jgmro3VAHKiLx7G1kKOylAp4A+R3G
YGEFM3/2lvbzawzIfE0nMAK7eE+Xz1e8t+GXcvj+akdMo/TBFe/EdCfFd4w3jwKj
CTrshN1mW63XX+HvbbFfyUFmqPK68C4/X2ywv/aMD/rYOOoOrG7OYRTRo7tsPosq
EdMQsAwW/wbxE8LjnfKj7RrHEr0OzDHoKEAPy1W0wIwre0zRR/WzICPvCcY2zNT2
nWVsGthYR5cILwsFMzoeJqyqBdsLyvPQNhNgpIJ9bVhMV0MrvDReIeZIsrBou9lF
GNODlUURDX0MtzkQnyoPLnHsbklP+Mmk4Xp43rPhAGqmyKCifwLxitSVD2wfPmdO
496C+p4ZPFQKnPd1JNPq5JUnSe+obOZWqBIaMYCpUCLEU2YNDyWTAHojiVPvYGKF
fnNzsKFT4MkkEfS5BNwsofLCN9/MaXbepYGwyPWvQAFtGnkWgRqAAH4dJnkMKOFx
iq7w3FM5/nMMEyCeFlvii/qrfyvkLWOYPLuFcPBzJhcaRHIAl9Igm5G45zo/3iOr
g8wILwthx+JD7EtZAd5keiZstzMoJIBf5/Lls+Wg7cpfJdvrHEalS+BJHBhODN5O
53yoETtebiJchzQSqbRgdgbtuUb8IrB7BrfL0M9SbtXXNsk/kQELNML59+FjbaS3
uWq0sqjqwcStn0z9EM8apeN9wQMhxTf6yA7piIYVsTX8O8XblfY16O933LaAQ27X
s4QYG+fPItl2UxIEYw1YaY539JwkgWsRZe0j6u70W6cZO1xXYU9BDY+yiWrntdED
CapbdxUisRlnbqbqpGMdrI8cXj83ZVuWPdBpq9jh8pUg2lwr5oFaNjJb7UDrvYa9
lJo6Vdd+TfhH5vvBt4HISHpOMPBMlhTkLJArYJOPP/u0GHH90P5cHkj5Q72VsmcY
eKXi/+hlhbReYC/z3nZwY+SmOLvM/yFw9Df6+tekFk0VmZNlWNHq2HHjGf3oCaZ2
jLcpZFRw83KDrZ5TgLag/LleaggNl5T8khVFqtxEt8bEKoXRgDAFc3SGKWQB2jLU
mUXj0ozIUU5lzVPfz5D8eytAYKva4kvFQpI9rhNCeioGP4DaOEVKAe09NB2kZgqa
ZMHhLdSpVBgzUEx9gv8haBcvskyw526Z27FCJJy3A+f5oCmz7joYUaqKdtpgnrrk
OmdLqyIHc8otms+vO9rN6weL83BxLBq06Nq7CK5uI5U/gYp8kkTuHKC9m37ZHBLF
YT/HlSdNfn6SmdsEKxKe8XPNQnoKWOt/zodeAmO55NbNzPyX4RGJVlVEPdSTc9nB
Nm06sUb+Tl8VcmI6LkGklwc8ldblTeK0qr2tBacaEYri7WHEpyq2hwCKqK+w068X
3vTiqq5De/FEL+xD3pIqxictNpTE0e5H0V5BBnyVw2he5UmDm/jl+t/XA6lScuQs
j5ZSyK719dxv5URkRKf8eA/5k71yiGATXUzeEi/PZqP9qASD4Ag5A9oM6k0iSBrh
r4RplN5SPBCphyD+pvrf/XGCOAsROHgmW2mn4xur6pqntOnd+44Mwo1IfGqlmtuS
QobB7JdW7/CIJGNGrLGubUu0XT0lHWtjy8I1cwcJ8NA1CNNqKkQxcHLghVmUaoTR
25ckPKRfV6R/HIjPC6ftjB0lZKTQzsf1DRB9qjQK0k8O7QW348/DXf1iX8d26UH3
WsIHaBvWHwtHSlF4dNL6WajqBpNuzkvEKRNgePpS3xWbJjzloEG7DsipTg/NH/Sp
zKQEVAxG5d6PBj9Em447SaDSYzZblHE6iwXEP7YCRhgbBrJ9Kl4yj0m76MnEkasu
lFwJR94onn7ySqMu0TaAVnHd/mihTDWCSshwdDYhk3AZOzoB2vNexI27CqIrOGI1
x7WvCley5tje8LPPe8IZiyFs/+9lGUdWmMpwyK4BQ+SCd+NC9pgrcoYVXjEIreFT
nKkD/3Wc9NGI0i0nueWoBRAAOXf53Vzvu9+PNgMiKo8KwENvW915myY+2/nrNuXL
zQbF/beUgZp8pi1/wXmuoyEqhraYFb7886y0wCZEkZ2VdOsVUjy2NDEBeyGAjsGs
ZgGJz5uBhTRmcNoYkakvvJBSd6ciBVvnSn3/Z51lzZrSe3OhNYnpM+RZnNd4os4V
a9HM4p9irQFP6m21/L+JkhdCJTBZ9qaHiAy7HBjTk/uYKoCre2jpye76xOGuIHPb
LhdEiqUNayazPksyrYbyt+NAHEzUsNZDfnIICRmbyfRfUFebTu1UNn2w5pMhnybR
cdAACDvaLSsXjRg6G28DSn5nDxIx8qSX/wNJ+KnoN2cHLvcP8VgfpFOSv3KSVsen
drN2AEQ1Grn8ZdLTAdXKsFbbUArX2C4MFMwhcvdSHiE/ecFrQKwhZhEIePdQE0cq
KDMmJrWmqbzLJaLYmzqRmO9P36YSR0AsGOCmp5zEBc3FPzXoPzS9EPJfTLuuSB5U
exKCtxigoFvPOJsc9VtNlFv/7t5FtbOffgJKeP5Q6PHib9Yvn2khww29N/AP4FiX
93O/2+OPa0KGD6hAMVzU0mN/LO6jlRRbb9aKA2lifXwX1wM2qvQcrvXjrBN8RztY
Vu9HPjfhAGifbUzNBCT0OecCaytG0syaORaWnfgbYhIoyEMEYtw+TlWvMMGwm3oh
m0WreW/xbWh2tVK/K/f8yqQ0t9p3YQoRx7VkBXyvoTlZ5tc/TycujJoEqzFFb24E
Pk4wpGlSE4IGs+QSNklAoeOa1nvkYKI13B9fDz3wOFrPRnlL+GfPV7qtAbA4iVFM
nUh2K+xeE+NmL48YbbOJeZ5KchRr1nA7nCvGY/5qgxD/wuBYc9ob9Mu0SitMIHxk
aZtZ8w7NeDBUkVmmdppZdMiB8ChYa3Ee0uOpRw24OcFTvXF9MGb9z6FMNHbGGFIU
gkC2GCCmL6dSIeAZ3TynKe5coWyEfuw4aflrwHwD0b6ubhFwwwR6Bsa41GgZJV28
UBp+gBFIWh9xGeVxx8ZTVgKRcra+wqpbZVuZ7s4f7FAONEQJWIQA56mZmecu3rrk
cnOb72r5Ek5VWZetfXLu+s3Ugq1N21OzJ3LKK8hyUf/FweQ+83v7NzFTVRmFHW3A
yFSM+tfmeUnhe51eHS5WuIq5QUBz0ANtCGyiy/UZTd+X9dgfoLrsEP4ozGQJkdqF
vk8TTDotDQ8JvtkwH4vRRgj7qkA9nGO5TzfOGUjhieW2o0HPziZbaApu+wejrIDQ
IRGbj7pxdqu5fx64O5+9Cz0FT611qIFGKQd0anCYv5k/Jt8R+5FxBUjjRbsEFamG
FkHrRYRCvDWtk21R2w1ZjNPZPhpj7cDyHX8uIVtoLMezQGSTsJKRu6kxgVLYtGgT
Zu84EjshEQAEkC4EgCNNlnTEJhYPjb2e3k9s4fKF9ovbA/h+A9K4HcoIaIpUlFz7
akj1s27UUVNmwrIE3S9+0kKAYw7HiEW9u7wxP5+AWeD2a6S2LzW4BucqxDmSBZWw
tsxoR3w7aNEdftXgMMA3iJmS/t6+pXJJdEVY5JoTKjD+NeDglK50vpEIlQMNE12w
3OUfV/EFASXFa5tJtOujUhtIS8cc+IPTN65zPMTurHrV5p4h97spO8oQB8EuWixl
X8/fWbvZPuOMscq+5Vd22xDaL5sNH17MZgNJJhWGQxoyDfo+/3mSZsQ4OUjRVb+0
hOS8blohqvS0pA4mlaCadAEjjRcm3NicGHK0BgZm65UnjSoy8jEJ8dhRV7ZImZGa
BgzcKfeaKQj62eHO6HqZKdpmTMyV5lKsiPiqSDGxBY0OoKadNa/BYEHgRQ2RMCWO
HovCwZ+3MU5n7kPZ2nboWDOCYk4a9dbiMUtBjOR0Z0VWKEHchrqDc6sPBEPhM7Jo
fezhdOG27fZeR19T0e1wVb71OEfeCJ9JsDVUzUD7BPrtA7tPUB3xadRYBdqgfy1g
Bce2A6Ca+ZjF/VIFNm91C5X+QS1PXvZ0EFTVS4OcizsEVFxTD+VYR0VKregzZdNj
LQMRSiZ+ez/vW2SyUu+zJroNdJ+tVSVuZB+mCeiXzco5cs/kI2/Lbzmhb/qexDTJ
YKTHLAWx+zS5rwUnKQbKCmOW/2QlzjU3UCY5qc27Avf8dZEstJjE2yD2vHoydeGn
Efl9DoUgf8VbLuySiPJZ4tX5mOkytVZZJrXpyjsLT6KraXrsEjwD1nZRYvHfH3jT
TG7DRkWvLtajBTWvmp4toT7QLQ9Cm8tmfs2c3a42Q6v/F2i5NaCFD54KnJkgVYYY
elfSTKNjYFoNwluUgzqy3n9eOo7xhRHwCSfc0bE/z4uhc/9MshzL5lj6XcHJNQKC
aPwEnrF456SKaVID8MH5TJny9JkuUjuJTqpFdEj3o8ZVQb2s7X5JASSnsks5wrYb
7rmpXESSX6koG9VVMBHnCcQ/NbBTeGN5BK9C0ccA7eiNFI760vcwmLIkKkC1Z/TX
M85oyQjxQF66ih8sseWpGT0tUdBdK2FKjZ+YJolR6QhfLGL1lxI5UO2InjW2H6q0
P3r6vgaxkiF71wJXPOCYOoKNzTh8liMkf+e1rE0UTYrv0VvQmCVxlveqVaUI64LA
KAH315ltt0iSpB+dyrm+L9Xt+hoKXlWPtPv+TwVQ0Glm6Jjf5q3NMeiSnQUuwCtA
m+K73B7J7Ird5dJkAFSY3W7KzTCR2JquDGh6k5s5QjVcC4qa05r0Ms+0b5Twn1Fa
U9wl3q1vE67D5i10qHVeETTmxRFX6dlRf+64r0hhqBQMKr9h0ancoXljSiupcmxv
WfDuMW9LT+ly5dYMCJ2HhOoQIG4qtPIP/XlqsGwd+Wcp0wKQeMY5Ud8xfdkMbAfa
eRBBytPJgU/rmIz29yrHpDK6Y52M6xqLA6NDqdmXUgfcCzFgT79yTtNm2tzElh49
EDHzshmwSRVmjmJYVeEOsQ9iL9seTz2rjGBlGfQRW8Q77olA8KVfHJTZKIpw1YL+
F35BYgByoJsvJxMeJtp4MGff/z+hW/6zXlZvfVIkQUZw4Vtx40DlQ0chSvCaVFNU
xUNm7WRDpCCuZimMqP92t6cZi/041o4Igaf4ajCL63yNAIvT8bK/lSqKqyjPruBE
l8W4Qptl9ZOE4ETScjfNTOZmZcnIggxDDCAhtde3GgGsOpXooQJ2LF5BNEKjd9F3
HW+viPKmqMbwmvCXioC5sRS/i18eFyF7TnwW6rDBEZmNB+WFVkN6RL4f95pOcYkw
J1D8mT5PBtFkKgSb+Y18bHMm6S39oFUuVmkO7kUvZzUAgvNtLzvf54rWAVWMvWcx
+qTDzZOhbOQUpiI3zeyALlKOce5+ECiKhiN/ebLKSfBwX6Pc6Jw1/i3Q752QSS+C
D5knnhotLeA2kmxGDen7jWWb+SlSGBwZKB2o7R2ZCm4b6GFxEWZKDqOFb5vlF1Gu
ehxq7MDaIRdc6iyGlzaAlKM+kIYZtZV1QMehL22zyzwKlN148tDKoTI810MANvnG
J/lytJ+TUovoS4i9irDzQ6NFzVE+n5BVJvmNXAvq8/BPUGcGscqQH+ZC9YWeMEtO
9qY8vRQnNtypcQEdQjGLsBCB+nTCqD1uShy6m4LsOWo3JCAf6sKe3V3duNJ7bdO4
fWrVEHcYzgYRUsKgSGLwtC8Sgi9TtoXYHvZF2anEKCDOcYiLtql+CA8gn1UQnlaP
wKvLhTA+eXw4E3DAjYUYUntO26tp6fn3zduHXE3j+hq/NvK7PWYAoBOZtfz38K5I
ZtOwECZSdx4It7ApnbmaI8X4/b/rjxICHouWvGplHzLIYOFId9eInFL9qSx1cbzM
60mH6NGHcufdw+XD2mDTzejPVJUgwlY3kj4+SY4GQv1eLo71uSMBzBESRj+rcVqz
t3ZeOqphJbX7+o551QeqC3KkFRvgSX461z021biTiRBzhOCVB97NEOs9J9DMWrfD
wQF5YKWAWsL6lfydcV6CzFD6sU37dv9SuE0M2qf6k4z0/LvexWEaNPlkr9tYNXBE
DIuliu6HDnuyX4i0M7TLxBG5hnRfblH15y/Fy1UentahEfBxjFFjSGMRv2vVKxq5
w+MIjS9mYngGvpIf1zsXz4ePU2OD98YJ25YUCjJ8osLTF+5yHOm+WGCbQuZrJEc0
rltA2nogfpRJFrZ65yAd4jWURY64Gg1xDysWiu4gjrz1mJ3BFqqcE89GVqxp7LEq
o858Egr+UsdX/ccGP2U1jiaSYWrJYcq+uaQ0SMJhjtpSDwR2l1a2egUixYyytM5A
V9sAEcCqySMhMGzLEP0zT+K0zWeF3ctBeS4u/cEsPMBc52rU6S1tquWcyErbkcf7
XkWcwcd6EqapuYKPBgIU4o0qfVfLKxePH7/G5dDOAeo0iTzq7eNLwhXAWrbVlwJH
x3IgjAWHIgA7lQfZz9EBAZnzfe8DdTRlnXJhoERoCyT0Nt5iVhRq+hILb+CDcTtg
x+CjvKzDINFqPt4i07U9D81C32sVmuIU6pDtZ5WV3F9nO6o61QdSx2BicEFkZh72
QNyLCZyFg+/70+yqSPzlUwVN02lkh8ubl/Kqav17HPQm/jvkKd5uj3zp+C+FFa7n
cXNG1PdoME+ZeENUhXFhg7fAcMv++WPpYrrjFywuRep1M/NxtUAeLYdiwOxvqpdW
7ShMIkMFpx8BMcGA3258Bl7LORdDqqtl+fNtrnXhoeodESu23kVGKMCjRytMsJ2y
40lPFa5j3kYM0SPhJwaLPFsgqfh2Ygt6KGJ5ojNa3g2hNIcxFKdzIl1d0gAbTJO6
CDtpaBmu3oMGibyTIvuK5osGYPTip5K1KOdRvWUalpeG04l0w9tlsHbzAeXu+I+V
XXi1VZDxCGR2UtOiYfs9yEbj5+ZEeNjhxiqbNjGlVD1ZxrPsoec/7IIpQFICnaR0
wLmSOwED3D37BnRZatnsamsLq6o3YM19MIEqeZd7n3nbmmuWKqgZxueSmk1nKj25
QMztSzcaxWuBzPIVOzmHJ+/F2037at9VYdBq287jMVtwKc0cFOdpALkYUHst0EHC
JcmSSAuuYY/U7+J+dVD+BNk4pbXk621TE+2YARXLFDNDx6BGcjsNJOn0CY8GJuUg
w7Tku43dAmpws0TVodSYgkaQqP2TZ0rHFOWA6OkEHqU0HJioB2GPrVMbY/nq3FiP
R5R6AgZmmsntejtX5NIYSntPNUZMCFEZh3Cd/kgv64R0K54ucaQBrF7qs+c2sWAS
gl+Z3rlMBd7lgT6yeEOUfE9NplVsTkLfv74JNOLjuryzovZoJw4LsI+epaglXaaT
R7MKNaBxT3ORRru5VO7/E/e2/HzjPYmTKqT4uRlzpg9zZAnXu0JvpquTNtMPLB4H
SpjslOnm7vU92rVyHlJkAPoI+LSxxBUo3Z2C/nBYhzWTBhOKaovy8aNuSbT80ljT
wvqbS5I/9hjW4Oat5nHJHerZIKLvIeBoHow0srhhvrDAdrkeBUpwQQtuPnCQWDWd
S4LmBd9/r/Z6AWoNxtcGlvrVEE4v6eY+hm+sMxLBNH30TRcZHsaFVFmJjTLq+b1R
nw+YHkqJt23kGgpG481bR75uX5IrWVY/RIsu89Zx94A1UwU1uRthqEwxIBooEcj5
ByANFveRHBgjMo5LSS+qKQckHF0BIGT/GLwZUC9UPmbHFS4DeUyk2+SBHZIX+uTR
yiv/+g8Acd1Oyt+NAhKgppvpciwjjWiqRTfN1T/Onn5DbBAnmkf05ZS4B+kCiKpl
1KWtMZoNAMxbQ1SS9RTVr+s+oNIvJYSVumg7wHcJpkxLEl9DfVF5HwsE16fi/Chh
LMii0TOV6X4ZJf/RVDSKcEM5IDzkpzW26tV+g9ovxnfKyDwd+s1gK5FUVGAmglqh
RQWW0sJFl8xnnQRKLq6VywWERlPdkWf5WbMjrn28dAC+1FGDOTWVx5LUC4uG9PfU
vzEVKgo9R8pcVU5ZnM9jScE4PNTUPccK0GN+FsBSnysNPue3RjL6e91FGfbq0D78
M3XIb6Z7pWZwfM8NMyRZkby9cKw35SnkM7Rq4SnsH5MCt8EFu5GdaAHHt7ZDlp1a
oBiaTdIJCMvSetMJhd7J/yqRRaCagOXhR/zrEa+hzbSKXu7si0n1CfiUspqA8MoK
nrFGbE1gl3rMfZPR9Mv6CanLOpmm6nYFWHcQEnxfYO6PVYbk3XchujwgQgueubwg
uJw5FA23QOTYFJCifPAMJCjgA3limI24Lsks9j8/64Ls1w5EONV1cxS0/hB/TEOD
C079pXyyIbNLB9r0fyJEmOHG+Q3b3N1QEg/ohpTN+gcOw/x+efi6vt6jrFNpT9mR
C3Ke6im/1hKUQary7l7+Efc7Pz1biC7XoQUc6jPIWV16o255u3PSdKbIE2snCDz6
N7XafqhDiaBZPmct4BSidCEIrXY7ey7cv/03fzZL3xo3gWCvXn12ayotnx2cqNMK
vT5xat/sVJ7NB76pJ3/YxuaiOvTdD9xl0paVDCImhlaUXOQlOAkNjAsUWFdNyLJw
bWo+qOtQSJ1+hfYKb2TqtdqGpELqlEbUrLMkq7TIpXDlAkOIDekkWsjLUtffir5T
Y3Mh5MzzTC/x970Y+3DBvQoTJmBCE2j6MLKHzxzZ7AUxzxf07/1FxwPSF4MzjqO7
94jF04bpLLeBpPwz+J5QinFS3Q72ZLGxBpBb+D+g9673xx3KgtDLzrmz63sBV5Ra
8rh87GX3ApvWOnTSfVKtvXk7/K375kT9sJOmC7XysMMFd/m+TEuGM42aD/1nx7uy
qF0kgSMglRgY3s0TUkU19ZSRWq6wirP5t48wwdgtphyee2gnJ8HE2pfDGj/10pOh
73Rg8OKIPUi0q+HtNglzPIiNgXcH0ca0JFjXKXYG6nvyaifVplQpeENNVrwEo2DG
OSkBG7RlBFMyxne2HaEL7mQyvle2y5edD7hpNVePka41ljx+lWcoq6nnQLp8k58W
V10+vkQ0s733t05R/gZn+iRsbD5A/l+fphGAY63TUJYVVjQ5BNUXFqrZWaZctG5q
6naAxFtxwkP7oRkOPmC5wFo1gE6ULAB7Kqv6x0U0xyAuw25jc/KJFkOIdq5ofV1L
LIrBc5XT2oqjzVKEkZ5rlU9wpMx00f1CGWcMCLWnygohvC0XCqu1a1c1hAJJrEZ/
lNlY78DF9CmNye3Vj8JdejrzuC+0HkTlTJnM/jF5x3wSdXLi3U+4Ai2kLw9PQGuI
Uer5YN5iTyTmY26jzikbFrFKKwnXXSS61BdkjIQaoqcU9w9iFQLFDRbX+7zP+3Sf
zZO1TQxufhKo2Tc80quWFdSQWvQruyELFZg5VZwYHgcRWsUhYNQndyVomwR3hKuP
ca775TLRn/g/VOTUPrh7Ok6Yjt/7PthMnS/OiryvCsTqEICpN/OEqz5r+L6qlbaj
SB1u6rRLn9QbVHjcdlK0/4MMOWT3Z4/hUocvQ3jIxoYDRQ5OdcUIo+QXbXBnp1/a
DMqypa54h9o9fdK+6aytPb9ZRmKTMcv79DxlsSs1G2wpbKeZSGRe36HBRp2JALpj
vCvqD2bgUv1SmVSpUCIF7NBUcKsl3WwGNO1JFWyuzQwWHrsVDZ7osbHaZAB6XCfx
LP9SeJeetc2kZB4wdvces/cpju9jU84JVaK206h+RZtoBtUqFJsHlJDcnze986mC
RNx06Q8gZdIG87CgLWhBU0wH+eB3eZbVVlvIORQRArZ6AOzRmM70JMK+q4PT9Uy1
QLK01fHneQ7R7NjswGRiU0tYZIm2MQ6cF7bAeaofR7KpbD6rKb0BDIeaCDpU1+Xf
4buAjqzgPju5snhYpuarcbCC+BPSNZvPLPQcUqYQ08vV11gxPF35c6QoMRGTAXAH
v4GAnhnWJv5ccCURd1qlCQAm5nTT1v85OGhhtKQsjuvk933CIk5XAa5t8scEpZwp
FBVFLmQsvDT/V907XutZnNRYPUYGyhRJBjQkXtwMEVLNQ05QyJctlPxVi59slnL2
qKe69oOdI/lzir4CHXsSML15Gq60w5mz0qN8iiQC0stU6z8L88NdtXh5pV5MaKFP
ZJ1Nrca7wsIOe+B4olVCk8ucX6DYU8rthHvZR1b6UCN8PrU+8hse7Z60v2xmTVhD
dvgXKWWz9l1ViDKX74dZCqfhprG9r8PS6bUNLhfogNJwCYCBI2L84f4k5OKdlFDe
8xpUv7epK6lKsUdcVfKNv1REiHfM2zC5FpwKQ+Lb4gM/ouFGCflgEqLuIt1jvIqN
UvQ3HdLDoqwbhPk8wYGh+VpmiURlqXhA5a/h8GSaVqzE00y2D4SQt4C6EsXWH/SV
Gpbe2GblDbqymP+L3hUTBKg+wytE0R9ZhIvv0DSqlKQ7dpv9OIHdKA5cOJCOwwXo
WwIicuFEkAtQ1lzBQvDhxTaXXUCDGoYTQfMzmaKv+00VAmUUTEPcVw6RwzghhwvV
YxsoogVtRCuU3I5IzKHF+NO4FGCpI7Xjy3ZR2vbds/bhbZbZSH4DJVzxyxZZoitL
1HDiAZL1O+PyGlO12dZgXiC4vKW5va3QPabVBJG5YUhq/pXlwU+aIgE3xt5peqHg
9WY+o6PTdz9RGRUy0qMdxxs4dazfvxusvZ5eoUtZVl1cZXpsAN/5ADrtS5xF+ZFU
sBFHBEmhpYe53+b9hVv7fPsPOYC87/6YY5/KKNezsNzRwsKqoyl2KVTdCWXP+Srt
p6tHd41KgFx8xN5ZRQu7PKIm0Gqa6Uln0fm2DSbKSX99YtLt7Uwws2JktMZ15oGc
PwyLaCpCQlhnhFpKS6wNvWMeLT6Tx4hX0oOw4+x/bRU3hm/r4ZUBywI5KhLijBvg
mem3jl3j95P/4POwpQG/pNkt3w8C32q3OXySE1swn2+L+9XUN1AMBz5qwuA865wb
1HllGsTyVm2Z/e98QMmYYAAjt/SFVTkBmXRX8vKf6nq/Q33RV1gHDyX+djjLiYKd
wBgShfI3HT6HZQpR7UkkjjXDH7x3coa/dCCObeXv+9H8Z2a9+ITw5Rjwv07RpkjU
PgQCmPBO3tkwoth/M5x3TFlEHBxOsoEAukCnfwEz2V0D1FdtKvBRen6DABb5adKq
nykr2toGU3cViZRPvd7E3lsnfh+VUm3npPwUdBtL0NlFi7yx6kNTPq1s4+wTUrav
/MCWNCmipTWVB9t/2IY5lP8XLk+jGv7eJt9JroU4iQRpy6/7MU0ew9+XLbFQjIWu
hI/sx9em5+2kZTFZyNMjuwtE4vKuu9Heku4r/cAIrzJKHPNW4TLiniTzGHHquWAx
6n4Ie1t+UfKKSuuHnE8pcpfdk4Nd6AyN/fAWZRs0eUZg/lzCnEReBmFKPEUNQDre
vATfrSc+xSr+SXZhlfX3/8UBia4606wFhUqBZ1wTYDw1eepwVgh9OqhY2TYqoxU0
cffDinbH9gibnEahQAolvxTBDi2hjB9EPWexJP+ya4xTtlJWxrex/2ZWUnlRoCY+
gJK6n/WmVxjWIUiCmVe5F2SqX6KEwvnH1UJNorN3s9UzGgkzq4gsb5MsLfeQYcAj
QehjNSZKwMv0HurQnMGxwzu4Vx7kGVZ0QxN/S96RmAsTk8sXdKQh4V0RyrlCqYPK
qqqOvdJuHXiUNYDuKFOedaSPcq9jKPaw5CKiMP82VWxqqB3DC85egJ0I+4E5s+1M
R/b6+dqaKIqp0P8cjgqUBxvFYfjud+vO+k/oYr03ZuedvxJurr5SQEKvNDGVvCte
L8esZ987dSXEHcU76tB0Y3ZhVOy7C9fwduKQM+dPqtxDT1Hq0SZ5lOaAwkfDF/Z9
OPrd1bN7C+1GH/Uu4JDUiG6TDCkkyRNU1zMbzzke5S+fGxuw19CCs0mECO9a5TDR
4G5k9p3Li83J/iuF+UXHnIgDeiC/k0r8azI6dC9Alx63IIU25YJ2t27FlTPlD+eE
v53G/UIWIc0ZxPEYljfWGcZwJUbffAQYmmMpciUQHX5FngONyRe4z7VWu4ZVPQii
i5l/AQlLlmF+fr4lQa0eK/ljJyGht64nO08SuaAjHZrWN5jnXggWISUvkntVyXuc
WZAQPhpcjCDXzxiQg4vBbcrtLyJ05IViCQRNH8CuLKuv8zbRxwjLjJEzJUloYoaK
LhYvWJuRUc0vt5J8Z0OJJwRXfW8wHqIpi8+5uAwFi+DD5ZSEuKYMPLJIFafTfwem
FGYaAk0A1c5bv282DwhQCedZuNwr5pFeWyQ3LJQ+CoDz/TpPQ5iMqEGJt4Hn65wd
zU9/LH4lWJG/suD55+AYJf58AlHcIu+4usSclSgx+reI2CvIUpOO7T6Cd0aic/t6
RXUGaaW46/8Gej1qIG9lNKw/1zLAk5dtTRKHVykK0mmtuYxOsGLc/jcm8BpqPpU8
PJx7H8jIPJxz0CE3wAcl3kw2niAIfp/sRjk0RXZDTi5DcZhesy7y7uT4hVnNm/s1
N516GYK9iEbBdi6hJVkAjndLB6ncOluE9tcdxBFu6AjUWVHEIHmdqUZEgN4pZEz7
iIVVTLKqxr6KLgkpnex4sg5tTv/PJGcs1Hz3wd6J6MhIacIJY7AqZHAhbSed/TLy
j+b0P1xJynvC52bTFtOdRts/fFOWk+ESVvZWjr2ugw+B92QTqjoiekrXknh46A8O
+FsL54DxTDL6E1ZaOIGDLea62DgsbTtDFXtLG+JgCo4g9V8IkwPuBX8s7qkpcu8L
sE1hHcDKG5eOouXygX3lfm1zPtcJOU8VTT7rDiXfugb1nOBn3nKxJgVR1AK6TgwS
4dHjL3kyiFCkG/JmEvj+TOq0dXhjwT8jqxDKstWYTzEqRzYhDZCWBaFQ3iqP7uVW
51jALHxKvb365ypdeFljSGWFbmSCo+IwcavaWJOhOkZVMQGuYZgJqsegcj76B7Qv
WO+mjRoSocxJ+t7UdI3KtKGs3g1G32vEjuf0mopjJhYnxIc0lZHOem2sx2pqc70A
i29h+no890BqrlZdo2Y+HlNruqjtBa7HUgynsu9MrwE1hlRhx+0aNRHX+LgWjBO7
uRpwemRN+RFQm89zeUJWBujSShsr/xl9uLdlsce9fybjaWrQrGGiXbBFSu17Hxcg
lltAI1RwFwIeAs++QbJ3A9dJ0J46da6rhAlVdoSSnr6+Uv2q0XbsI+fXL7lPHW2K
sUaixVZrvOuZBYI0Yrvi+sdAq3WwnRDAjJsrwbWCLe3XQjPD3KaNSzf/+f99Tqsp
4GYWoqBSm6yffIpjEvqdnMwuH4iIgZcYFDr9xLPs+l28JGB3Mlm9MU9ANRiHUve3
iyWwrcjcI8R2dR49bQ9G1sSTIRlN9Y8Mq+2BYIhCgCUxqsx00agI4Z4AQqH5NhCK
Iyo144mJC/1dQ/8SyjCgfnZhOYDREtU5vuPD3Tj/086t42ESSYQOgqYJx8EmUL81
sQfyVmW2QJ+ifiZhdp0cQiaA7kTyyq7sS73e/+YPD/aJOhilY4tg7KBlm6nP0kGC
FTYbkrj0sq9spQnqS3YQKcOp+ayMuOMZmPdYYG5jKzEC4mrlYjueWslLQv6LpChe
SNOljPRRnLdumxqxNwTS5cPUju9FqFJQfVCXozZEc9ACMB/u4fVq2YbZ0NVsbLoK
xscGMt39x9zqWjV3gJcVos2UUWktWqNYNGYwB1GlMAzYbE5mcISLHfolQf52wg/d
y7IFqlqMWZXZZ6qGgRVJ3jFRJh6CyiYck00tR/u6CGqCNtXuMUkRkXuP3B9lcm2l
qo8VhUsuvsZx71NeOWC+rKr3Pg7bgJHEYZI36Mcv1OX04vF/0o46Kk9QibmEty26
ZslHTSs0Ss5M8dMzGj+1A0SBy06lDGFycjWZipd0zDvgcgK/dIxEbVa/vt9qLvyK
Z3idpBc4fyImnS0Se/KK2gSQsUkA6b8fmKDcjM9dQv+SLw5+/pWSLWrqz5vCsP0o
w6yJj7Y7apuWUkXX746xBYHkCU/9SxPCgwoWZAqI50TP04QF6McPFJhm2xfspIzV
SC2TommBh9EiiwjJJwvmIAeRNBwQGyfoIXhf66FUwa6GzXM2AZlj0fLBr7UnTPRe
xmyZWiLHG6lKOan0W8dGzK5fSuLtcRSQB+sne/PxkPcmqCCxqG4A+70ApnBUiLPZ
9qZErJ2GUnQqrKC06r+9XsHjja6lCJ00c2Wwmhe2SYdmA7f6SPcDTFlZXgNR8ZS0
OIRpXBwEIahova8T+pqgs9ime4Aq81n6MtJU5tnn8qxgbfG6DWLYOA4TX6RYpgxS
gKjPFo4uoSuvzGS/eEUS6XGfScVmdSGYSVJRAW9p03VqreGDfPFjg7crmlta9iPc
M9olr6eBCSPLCKyIdgfX6bl829OD1BG+hoRRuRevJrbUbvmuJ0V7u2PmNbg27ZSX
TGZhgib9hl5OhEJJS3LzuC46ctFctSunzJM80cKfe3t2lCnigKXJyiMjcmjI5mRa
9E0yIlpNUUA4FS0hNBpeEvknEEUaYba5X3dQdOQMAqrBqlDB5jrHIPA8QeRZYkYw
SgOQ+snusjeWLzmUqpALeRWrxee8EXy65noxAenloUv1UfCN8XEJ5cQTBp3imhEE
ASSFJ6BrFjGVAg7LFSjSZogQUTq+O73h06m+Qd40xkYPAFAiNwoax9LE85QlDLUI
HpUKF0YGNwClHP/azO1c4JD61ejQc+DKTW3gETt176s1VciSTZS+wIukDJthbAe7
haqa3/QyBzloOh32OJXhzKZcdpzehQEHh/5aZY8aRzuNcZ7IuVoDeuJM1LqZ2QME
3K9QMFz/KqSosgGvYLSbcAQxDZb2m2Th67qto/JDyOp3/m1A2afRRUeQSmvZkORo
kAQ8jH4tQrRna85WrSXD4+Y5vrg2NFaJgvixLFwzXYbibkpjfe33KAtRAuCUoXMw
GcrQUZGRvkQiI5w2Syq5SstLJvaMh73HpwaenTecezd0cOgOdMS0eWK/CkuXEbxA
ZmVMBRm8we+RxVML/UO0+8k6Nx5ad8BKouqMLn9UbeiP+fxli//uHi38l54Vk4zK
bpnqb7qIzeTr4LZTKph7pzfo38aL1/3VJKu7m5DsziyqknWVKqmS/Mce0bvlgs9L
+kfRABEvpaaeWxbnnPm+gC6flEI3jtt9Xpf7pQGsCq6dGqBCwjFeOzXvCAfRGrta
wjS1G9WS6idsMzIf3jTKXagSI4dxo3BVHXaYNDM9T8CaY32ocxKEB0nj7GbR1XT9
Z40H1NKKk/pRC/CcwilgzsXuqb+1KrVwvxHVBvk1MdRNbaekqsK0X0meYnaOocI2
r+afVVOdYKJVCwSBcCcnozkzmDqE9CfFqc3MClgjSNrAYwVEo3GsqPaIyj5n8g3+
YrmvMPZs3uaBDbUdaX9dh3EYlSqd8u4h2m1DKoetqgm/oZptr90j7FBmXwFBXHNN
343kAdYSYGHwkk4IUGM2kitMwVtkSrxGqBv0hJK5JKdbNjfaeVr/Z8XrDm9MbzsL
Qkug5qUMbbf/MkJMrjgdJwVVFdoln3gjszmbjLceZA2lu0ntAsXZ2icN/7CFXy4c
oBVf+0+s6UYI1dTYIYlAzTvWRFsUsaeR/f7zu3J3OD9zmoiUaokw9YtCOECxJBc/
V9W/EELuq9nrmabr7A4DF8M5YKEMLj5i9iBVW7JS+k8yq8kGvdf1sk7USX+Zi+tL
LVpyqIRW1umJIC+7GX232A6lnQJPzkHKahV3AVbOACMA+hqr7F/9drVQ6QJ6i1Ju
D5cRjJuGigMqJiR63rAm8+IukCShXVsje8IGzrT5PN2UoPPZSPQ99Hh2N18uaubP
A6lkEplaDJn+bPftTMDcqww2yNpe7Cil7wwo9nTJYcqMtSPkDvQiJ3Jj72D++JhI
qQKFOUNJ2kURQ9dtLYkEb4+yAqqqgGMDl4uB0GK+ClvREq0dJD0uVanuNORo05e1
DX5unGfTT0zARnrO74uptRCQ6sOwsXNHKrsV2uwPg2wse7trEXsZTJfYvisjwGjJ
e3aI5IsWFF2qZUy840WKNn9frJbzfLu1ko1aRBI0JTxzQKpLywhw/muUpSM0J2o5
X9rxOOF7z7PRXg3iOMGqwagvy4k2NQ7pBQzk09UvqlNDdcKr2vD8X8ipI9h58QvM
Zz+hEfjAtqdO5GSbDWi3cBlKL2D0MmQmnwvvNpq0uYDqD5EEDIXTgT3UCeUeaTVs
DnXWaIvkylFU/MuFDJViiNZF9Rlt2uSKpKuBDDjPDAxInLj8OjFJObH27wD+cUuk
GAAQN1oS+NxRIl0VgSDfZBI3/kizLfbD17UpX958uUTF5HvDNZ0eTJq4ULc7A86R
7u1bJCiEOmU8yVC51LFLoFV6Kpx+Fzp3+D2V1FhWHOZI6nmnjk33K+1+EtLJ5rUx
g7O9QMYZobk78+vinuX5POoA65sp2T2UVFYbk27wnQcftzhCScMvqxPSV2o5hrEx
rHFI/xotqeDGmJ4I1YTWt9kbPBHTYjgO5hqqEPooQylLHZatuuprRWhJxhpNyQs+
k7pNYpV3d0aTKShfXKTp+VmK37sJOsyGYGmYrKg+Qk9zpuz/NO3edYMxqq8w37a/
oqiayLyBc9j9L60thtkTH/UXMp9qXVYF2tjMvbPkMdDW0AhnI9Le+5hoaCYkFpBB
ERN/LIKBxz+C3erhBBZQ+DnIt2E2VaA7Qc82W+fGnUWGS3rlrXLK/R+DnlZvYg0M
roTLoUoyu/l7iajwp+Xp9qsvvVCBjdAKIPptOtBz/cUHK0zsTZB5efYPouskUkBl
PxwiaFRrYgP1VIXDFyWI/eA1HX/Avic1Bat3olC8vY6yV+rsZmi2Aq0wWHWsczqA
CgWvKl5oPpNlVny6HfwqtjK3FyxwPkLRol8hq7b2/DbjNQTccjdZNytWmamzCxRh
hhhDsWPROeRop0YtGFqXhEa58gJpWsn7Cu0nJnJL8oAMAalEhr88VctEH/xBr/45
YE97GX5K/UWZgSIsXdG86QafP9DaCGEcs7EATl+yeUrk9FeJNxXJsh41u3PE7lWe
t20efftF5uqwTSWOo7sFNzpZmm0k7uzizlvw4TnveWV2zOeRZvFCr6gmXQJLOmTp
C5Rj/5BhSEk6X8jf/2gB1SW2Uua8vRmWmGkbq2CCUxZRWqbvWgHzT1CnEbaZuCix
rG81CPC05W7QMHJ5NT5Cm6k7o6J4zyjP0e7VRZ7Bh1iVTj1Ge6Q3I4u66xiiqjhK
DzKvZWgLzi8QfT5CfrCZ91PueQjbHdK45dalUZi0FlZEvu/Iv7rZGQPKbFfcgm+j
Xk7GFcXxB1fLzheRyikRL1rEW9dDoVZ44u3OzLu7ut+vNE/GCWGHVQaQLuuQ+Ux4
FaJsEyRkeoVqiqW4ttLX0aVIPGFpvDe8JHqvLEyIn3HAVj/F5DpOfk7ajNBKxv2j
qxZy7X+rh9lptexnE+6p9ZTcVGdKSXQrilT0xLkVfeurdDzMTwny2A2U1VXSHxQ7
rFSIhlVgCQz4y4YjjmxNm+W6xqZgvevLKe0EHmbSc2LUjz5DxSGDtpWObqzB87QE
ca5ORl1ldzyhRGEp0NBQ3RO+x4obbSnnq7exMTjiXsjGsQOn3hwsY08DV5818tcb
hoAMDg6eWmnU/0Kohr7pQXuwCi08+VlRAyipgqfTUTq2yqp2nsJkFGh6eI4bA5Yc
WX5ymqakFcvVglFVorsCa4Sz5VIpSDFuB8LUOEep4f7BtAJJfDwGt1V30hx+xKKZ
34r+0KzjOzdizESX6iHK50yiycLKdlm1FYWGxx8/EhsEa8QxNGxMU+5dWq153Abv
4oo6WKwKO+tvc1mL2FoPu0HEApcaiKK0MYF+ieIbJ5+OlPwFuxbSQFgUqYmhXn+F
LR6eimbm/NefdJ4LSNd7OggJidFNuVjJCeitKjzqxXGJgTUs7lzm37jklvCy8jkr
LnGjluWF5VcsUzi6EfikxXpaxGA0yePoqVRbXby2TrXNYQ5uNH2+Hvpq3FJ23aVS
icQ9ZQ1fCiGDR9RDhzkgMwzKpcz2OnTPk9a9NQCVR5jub5zEjAIAxkg4mHEcLmmW
/pqEtphJJcHAX7qvZkXV7qri4mAuOQNt+eJwEDj+tOGjMXFz+uBv8E1M2HT+lShQ
mIpJsH20j6yLY9UzMqPDvZRpGbk5UgyW5AvckVjVU22t41DhFYICN1AfoBH1jBwH
3W4A9bxTJayb0ZWhPaaMKJ4l7f+41CmK6yuMYSYv5PVwRKb+3uChTJgkvhX9lNc0
ygykxGHb0GOcdNUGoZ8Ye+ruP/s85xij2kbmRaVJEGZqfXL7aQU8b6le00Jlvovb
E05b0YoCWxJ5CWC3B9kWz2lnBOe+hdMusbhgpdvkm5J2OY6pZBgGyU16+A9TGI2L
L19qECJ/b5sWvVOczXIgqY/Zy28FtJFel9BIDzJsRx4FKzX2BCg12soYYI+tExYl
MuJrQRcG/2PDX53O0wEhuS+tAZUbnMIBkoxLgmik0G0gI3wxlhRrpg4wUWp2/z86
yUaQuY6IF3kQ5xtRNITXuSfSWqWwGIQ5JZHZ3RdI+ni6sgZwAX0I3ypeIiPSWx6X
fR4FHhnnObOyZU4UFqiugD406eNOuaUIIo22BqedVWo6Yr96Bdza05LmUGcVnSs9
rEIBDCcq1+ZgGt7fjKckQq+KkzE9HDNW8dgCqjyaHAsLqoT6vcFbVGLzz6GPZCLb
LjGwvxZGCh/vDeFk7XSGNayd+K5jM+QM/Kj4GzbTHyHAA00lgrBp1TdGJCIyXXsi
06HjQXtmuq5SG0Qk7KTZM3+UhRSnWOTYHiOc/TJks58fLOd+2SDQbJEP0P+I5RCE
fOtk4cbPkGss9pqNkCLDdpFBpPr7yWAh1Vmu/xp6zXZTylCieL20VFGLDfoGHZZS
IethQ3lzBfnOdnznyiq3c1NDyVv0R0qcEr013xYN4GFp59416e8CgBdbLdck4S1r
6alyuaVnWAvBkQC5lCOeE8GshgGU49z6MeUb+H7YPQoGLxS3skIfZV5DCnygcnEj
a5KTCOHI58o4NZvD6g/m+PiW5kLx/7wNQcFVd5UW8c+qt0KxnEjao7NsRn7xcW4V
ThdnV20UixXtEV7IRyZpNu7Y7EZr0ybFmKvq9HfwS4o1zsuBZfM8QQ2j5CSLxWk4
MD8/USBlZgYlhyqmj/K4w5ptfxatmc0iXYLQWJKPtmxcsAez9pNX9dpOFgp3EuWB
7wyrBrly6mQOc0veLJuDN0K3Ee5DFJYFcM/yJ+stUE00YX2cfHpPJAIKuhxZO9CH
GLfqSOHuiUBEsW2fGKtvPk1sgsyXH1GhAuEldhMPSowxXRXNSq610TwFb497JeqS
HJu3v9XAedLxbJ/i9oIl+8u2wZCv8qAaA7YcFwhAUCXCcz+4E7f79rHtLQlTy14A
dPOrKRS2WP8hZsZSkvQwdir+Yr2MZ4Bwxw89qS/8kV82bKC4KZ0LnVewE8qPwFWH
GSXOHRSH5vBlhDBH7WX0X0ikwx7tdFWr5HhFD6iDenF8a7Afl/b9Zgmu2thL0FsC
nmrxq4of03oaQRy9u0NpJI6a+wb455ppLQWS0Eepo8gxR3bvFv7TbmZh9j5qItd+
QtJnc0KUfcYFV+06sIoQON7mGxOT0WRHt7bfo3DWR1haopjn0vkbwe8xeEFPYspb
26qFEq4yhwURL5V0yg3XecbuzBZRX9eIM4ynuRSDDMGyQilg60dYwBulTfLpDJVg
fopQXFpFs970EE0+Sbj7Zn7Vcr+Ur3SxDoH41LAYb8+dF713tknYtzeyTVC5P8+g
4Jteb9usMsMMvyDamaxUhP+14DQT+Mot7+c5hFrA68yAA5O8wQx/uEmbx4oIxVms
sHoLmlY67Br5Cr5ewBqq8LoQ/pfooQ6cH//RFhmVNhRkd66PKS/LG3vVPVVny8k+
QKgA0DM/RCiWbOmjcpEkf7NUA5lwigQINWA66XqRXLwMsHUsMW1U+kjTHWE6kmed
8J+26To6e1uRAlo8FlSdQw290+wb6sDnLCC3OtqpOOo3JCDUOvEDDw6tYww37vQ4
5mhARX0Ji4TAsdzmB1IGws98TG0179a0543mjeJBFLYgd8YZlXMxojQsBhukJgpN
UMXoow2Zo3NXjkx7NYf4oS3A3FPBuaAJ5OmjkEahsoyj1SDk4a2TVUNsH1JqmlGI
SooLepaDjQyO9iXPsLRUyt9smQC3G+ZcXCeOX78LkA52LlLhKL/R02CibXzWhL4v
QoVafmBqVMidPIoWJ0UH7+5DtIM31PXSSkIK/+We1paxf1Z6J8mz3o9nujJhnsZ6
/9HS8CS6xVst4E1cSZ2XRlpW7JckQ4S5NSuQZNndbl4N46X5UsHHLUJ5jvYEPJt5
DfQKDtSMdANy4AauG9jrNUgFWU47cd/9V7YzVLbR7TKewT+l4nnsfJFcRXCiEwhy
jUhaCiszbUh1JXII6wKZ006oxkop4Ma03DvJvm9uef/NQKc1e1AcJlMw0dpTr2p3
O4aMEsgipfBGt81bVv+yxuCWMCW0LaZPCmsr1o12iGb+gRAt1Ed7O6Ev2lgVMl+n
1sfVQ9eB6JNylGqheCzkdkw2bkhE2wDFQl9fOoec7jBANst7scNnZEkxXoD8GcE2
kI+FzEZ8A/v86BXVT0R9gcRrXhOHfOoXenWx8pCuG0p8u7ePKZWJZXeysFv/zfY+
1D0t7g8hnD7Go7GBo2vmFKslbrfSsO9wgiI6/wvUUbQc5ASS7jgRjBBIUtBoFJmT
eCFf0LYGmmhRzP7xbNhXT19W6qzpNILO19xTDNUttUHWQIT1032NMEZGVSt0cOle
zsmZsIhpyo2M6k/DWN1ggTC4ec4k1cUtRlIuE/dkv6Uhc+px0oos1P5VNpKfPZUP
/zBhZ8SVljDDBTwYWsVp0m1Y18OBdfxjxpHU5ZuA2QPo/IJqfgh4ymGV3os9OPp7
gEnoM9l2KTHzEb8NmDdPtJrTPq2ja+C14ukU1wp48yjlTtFjj2oChO5qqfo4CPT8
KpxbWQVu7hja/J3PwdrRtE1y8mLIWYqIjD6F5KXTZELFH9gLR6wV8C/Rnvkd+aLB
ygQV/S78pMHabRpSYWD4dZuqUjF2JM8mNmLuNpSaSeewMMFLEFZ8yxisfygVYCLg
nqAzApvGYunJNPnrMUQWXPJnv3HMt8afaa6O+8cbRtL4UCpSaaFMSLx7wYvhCYkd
e3Tt7/Z5XTa7xRbrxmvSubg+Q5URfq3T5KpeYHNHC3lUhczxPyYBQ84WjBb/evuw
ldFgFxtEYZXuCX3skLWHGyxfwxDLwS7kWrlrhFdRkqBx8INTC4osjrya4JOkHGEB
iWIkK+cn4UkLEmDsV3828AOFOEqG4QaTfGJDRer3jaebnu/9FfYXpxhnDauL1SGE
SNRh3nCqBuhnH5FnyhLE3Bdvx/h6c3BYTkOz7hnGsIxMOUpi+nkgJhKX7TvzmzN5
6aDTUnbqBx6nzYBG2lm6yzDh2KApLxlI7QCgsVYIx7IKki+dFve0nywbrWCNazIR
weQ8pmTHSD8ar4wqMw3XOOqwB0452hhBBc38rC1xwPSdMKmvwysGjvLeXQHd+BCG
BZyn8ljqbEOF097SXqq/++gnDqq6nJMTIQGjD3mmZqi1grmf+4ocAv5VC46eWMDD
2VvNrQWIih94ss+wB8bLSmU0RL++/3QgwrHFlHmctpuVaTsSsk0s1kJWzeuETsDv
Ef7M/407uSy4Z9/cBW4ckToCkTlBBsoWAAKFwiodnou+JjrEKZoVVzOCG37BLsmA
kHLeCrep5qPKX0P7VJj4a7z1UaRE0fdn+/Y4asZm+C1ynoXEnSpVlqO0MKcbzh4h
fPI0VY1cjcr9YiTVQk2A7O6bZsZxI52ht5MOdGoFW44mP63MbOi/euXDbQ4jmqdh
FHNAkPuY3Adflo8ncczTolQEbje4PwnuZZM10ErIKZPckMR1nKsXvKqpOYGDGAlB
XN8Q9HATdrhSagew34V1bq4As9Pu2fBuanvZfIbKgXmYVK6bhpl3zCJ8gn5RaTgM
1Hhd5l+s43vQIed6IB+OHJG/4H5mst+ruF7C9sTPmF1uMCgP3QR3ke8fOIuu0ex4
QJqWADtMdl6SzXNfEpJmvPn3ZgSK936wXNXL+QB5W7MsTNPxrKMX0TnrYCzslxDx
TNNrTDzmWUMm1Ec5ufIhnCYQYUTSXBShxkTCGGObokMGvj9+sy8uhbihpNj586Pg
vXi1f6BfEpFxt/G2JHa516L8Q8LLJZEnywKVNfdcUxaWuoENIGqqCqESs4j/j7CE
+UXdLs2uNnGrWs/LYi2rtp30B8Ns03K074C8jRsdQ2YhjLkQMYUxH0JMBu3nn65T
0tNyZx9HNTT+8LIXDFLOwikR6veS3cyp+1R6Q+S1V3L/JAJAfu2ZY8tdeyeM8Ucn
OCOFsOgFlwhcmkQrHwQHtQij9NtLbLPplYRBSnihA7/dzWWCeYzE9c3mht7F5eTY
tTHeAMKNTfmUbdQWZE9Io6UQHiMTjPgbd1geYvr5Dl3NbtohfSa1ZKbfM4ulL+FP
8Jm0oczCjmZqaxAS1kjsUgdok5bEcly7MYohmle5UwRzTW3TUwCj5ZnyCe1WLQHz
6dR7yDJwHX0XPIUSJ1JEsCt0Bi7YpNVRFhESvPT5Tvg6OylYCduc+bI67seBLo9J
dAZUQP9uC6xAxqnldHDyNJjq16Mc99aIeTpIj4vM57FTDhrhfoJhfqgHqpccAwzG
UxjckcpsnftHdOfyEc0FGljjv2dHYzV6zfQG+aJChlL0YK69utClTBuzGvGiqVwL
zf3ziEpRc6xjzH9XULONH9fRZapd46jGpls1DiLhiMGW5rj0J43RyU6EyeJtLxEu
VxD2rfoVojq4til9k/UZGqCjTxgRhPcpAAQ3ZKlRRS50dJB6cVX3g2f1TI7sKVyX
kumuzfieBsluOSx7QWvPpxMnSM9oao4arJOz4fY+PwfaJif3UUL3+7U/22kLWGE1
3Mm3HO4RoEhPAKj+7axpqHpvuswciRbLj93PAoFxAKNlwyqjm7Hc5W0jdqPC4PI8
TRRWfzTirpW4B6wXRZ6guGV+wj7k3FDIoL+hng/+m1jISKiMwgge1X99njOVvODK
9KS58bYyeWvXsyTtvf3WsZ80N0xtUkFn73xXt/foz3lZiNVLbwl1IrLCMfc1JSwR
OLqqq/uHJJbzXwxJvZdR6FGjBjPwK7J0fE01Ra+PM2lEb/5zRNkZeW2K7fGMkiuH
bSfSQos22qGoQPcUBE4PFo/OWfGvUdB968yHGyBhsI1Wm2JvDua1bNzRpR1TZHtL
xMH9Is8uFmZsNX2SE8NBfvi06T1Kbn2E9BO1vTkAhn0nlhkCzVD1+eHveLqI2UdJ
aKfD+sYxTkkL9b6lGwiUggq6Vcgr18IoDv7dTYxflraIVxbUrq5Ya2EYvR2GZXRl
tp1X5CJV+yaYXvKIMa8kEskrMq30mUM0TTJYDbBDP1FphFQrPxiNEZVSu/F5L00H
cNWtqPUkspUYk67mqmgutCNrkERThHBcGgebWce0tz25mMiMspkBX0ISkLlEIcDM
k8AetCu3/JdlkG9lvC+B/BQw9bV1QJHDDHsARN1EwI9GNpMRSmUZ/W371P/Yg5g0
dfi9PFbrgVtbH/FIdxY3vseRGZIYJ54mBKRWGG1AOcJ2kPpjQYSiqAoA5maAm3hj
BV0u4CbQOs4A+mXif1GmVb9jnV4A7Mr0l1v79PUmrlAPkbAl08xHZns9IyGiYIdD
84aQr8Fd9cvVAC5dvwBIUpatPLLhh5wY3582sQAJHiSnHUGXCnE9XfBFW2qTibW1
ODtjnasDtZodR0JLZU8ZwMVmZEKbuDQT5b5yAlIneLs3ENKa2bSccAAJfaIAaeYP
+WhgexjDnsIGjYLDhHjP7cUw53YSWlR8iUz/euxO2T2z4HV92jwTDtUwNY5a571r
AO5AxQA49KhsZ8GSi90y3MI5FtdOCkEUIYQWk0pp8OfeDKJSrDSGRCZ/BX/Ox2MP
y1s5Ou2VTJYiEh1Qe6pig5VeDWpmIhMcnTdjaarijRQqv6m6fzPV3NVDuOP+TRMb
lF187igbwiK629ZRNkwslN0rSMKohqOXcTMNFj7lzMUh9reRLr4RWxf7pHTfflqs
QsiQXAEhdTRfM+bf4MlspbpPTUMbgje3mDGQqu7817MrUhNb3c5b3ZJIOlZIbRNV
STHHjsH9uNlOF/sPJDtbijWh9tGmwNWmnz2B/0qU4IgIv3JGt5KEaIOkrjZJSPhp
7U1B8AzgnY/ErxUGfKr2wRmEnsZ0COaaX+C5JpHJg0s3blwc+31qmte1V3oZRBWn
cNzLac5HcGDBpGq4dw4s2+LXWyHT1+c0xHvEojnI31SFHhaPDrE5g45Pbhg6JXq3
ECYssj2wxHhKEfFyQtyMAGpo9CWtjZMvVa+/8aud2Y4vRxEdAMEG3akaDzsRvJRC
ivn8Mugcab0ezzsDq5uNyZbmfpwT7FTInRsLacXYjBUHA4FXEpeSyWiMpxoMEwzc
nWDlEbNi02bxun74AlN8IelNXXkQxcQ70zlQLbscHVkwh0Unr9/zT+iEMwab+kk7
4ST2Vl6P/uzira2lBRn8zzlj3AljIx7/FUpriJtX3rxCbGRum6lq8GBfv2Jp/+Zk
aap6qa4L03/dXO/UmDCFgHiZRiG1m2V5MTQw3rCRRH4hf2wvbQneUf4ktlVvJGhL
/i/9ttN1MZjmuZQZHAmxQBGmqDXc+Ck1L5nSxW8rVEFls/u2+IOA4gnrR/kJBNbQ
W9lBnfoG4vWOU+SV8UBnRuNGDxwc3zr+I/HGzh/JSDHYffIDcRJinnTcLN6OKpQz
rtXAIXq0puamy7TTY3vWsK8PSCyQoJO0M/EOPxc71qFO3Db4PWWkcSU3kygCj4L3
AXQFrpCwhUbAJiXYZNgMII9kdj/3uLrQSB8QARt92NeOuToXZ+2FBWL5SiUREsij
xl2bG8VqAUxSZ0/0dmIiiVqm9kuDm+RkXV8MpTQjQPuZlTX2nc2uKDX6aXXHipTU
ruBKPu5oAkOXpPts0RHy+OYUy770rMdneWqT9SktSu8JA1CzCnYIdhuh692pBSEx
nCgH1OVdJfcFNH/WRb6Zsj+DV9kbnQwoPSh4swL6c5MmuoCylUbSZyj4u/TzEa95
VFxDEzQ2ccKXeMGdxhzFTFLIOnjFKEigxpOFJGvlnMvBNEQva2BdtEZrHAWPvtDs
SSzK4KiLFX8rueqqg+QF9fnCIKjivrO3aXUNyr0tzsJbfALRWbPnfprZLtYfLf+Z
nU3QYvAvBpsnaqU/L3HSJ/rZNoxd2P1CRiQkdMBf3sYZR9oRTV8I5hjDIFAbov2v
tRA3CrmsxUbXBPAjwfnjmHRSMPKo0oZm8RPl6yIi0GrknCo/lHigcXsIT/v24XsP
G9nyt7oa3tgXdU1jZP76dvUuKgN5coPnxtfwTTnTGOaT4sk5mzUnAvllFShFS7OJ
286E48Tdvq7RSNltMTc7tq/AkeWxRRRqfCBVUZqnNj3sEy3Vp6ye50zqswzsIsKA
s98Dz1t4uCqoz8/4R7DAgQiRLUqRpwx+ps/RcJ02AV0If4YzbYHmXvB4VvvZBqu+
7Trw5X9Fg9EaFiN9qd80DGz03VL8y1O8btCLqgc58dEXDQu3E5L67Seuu29IXwbS
pdpg5Y8P/0PvcfEXXJQUYMqCdAwQtxb54d5LVkxLZIHNBRvBZ3JlYXejAzu8of8j
sKz5CS5YsY/c/cc9tlQ6J7d0K4EN26jl+COuh4nvOc/RPggT7Qrz15PHRfOW3VJZ
l6dtJxJ6ii9AxMT0tgO5MjeYGd/Q8qacwGYf4txgORAeuE/IRxIEQlDH5fv2n2JY
co68mmBiqSa6reS+OjKbqWtwsgOCvAzQrYFChlMukEdwYBQh7tSHQC3+gB/Mqh9G
UxozYPXaBBNiMMZlyJoPjeoQw+XmGOl1RPjOeB07fpJQ/1iWPiV057KpZqOVa36F
qw1ryXv88u3u/7CPDoBLCyW6TAtH1HkGtxaQboidRoBN3cKPhxse9ulcocutIis8
+klFFx6Pz3UnY4VoP56ra1lHMY07OKwm0HF27cQogbcnSGVmPLZegMz5TohmNVJu
FnW4UwmYGiPXDUvnBo3pC/zkiQGskGQQIXbxMeE4iEa3eMNREK5Mhr5LdfiQl3ou
GBz4q9KqF9bE2aeh0KVV/wT0e82tUp2CP+X32uH+ETEMhVH2M6ZM+3b7C5em3VLZ
SDhsJ0VRB6xI2mlHdFwOC0R9MmP/v8C/2pUtFCvKJJiR/a6YJj/Ku228bQCe8jen
qAOi7Ef+kj9Xyy1ZDUjUv8A25VrnDfQ9LYBTzLClE3qCUh6uXOHUEUE5Yf8Za020
ExbbEkcJwOrKOFjU0iP4R7u4tTJ8ltrkR5laRvLwVgzCJTjBGcAcfCDN/IiMJocB
BDnP6oES6xt0lvAHtfxu/8xhX4TrUJSCWdck01D9x/OeCdRXwdUOCmbYvzb5d9dD
7aOcHB5oBKrdHZBYRiHne0GMPXMfAtHuSzku4RMOAPZf8lF/NNFM8MgUOvNaS4Ww
y2eN1AxBGaMIaXEsZUu4ePLphltdfZquwfyjZLJ4WR08nhCj3IdJSeN0kn4nMHKA
ydVU10FQetIZkxDn8btPrkZrLdeSQtAPZRr4ZSDyeeYqXJUW6ogYgL9sIhi7r8Uf
9z9erzisxzQrXliayufuJt2GUXLkxDmtc53n+paDmv7mAdvWcntXt5D0yr7ueNie
CkN5iq+rw3GvOY7cMycKTWF6T+3TJwWP+8GAuUp63rfA0nb5/Koovv2Ou75/wJBs
KhNpkRMYR93/nlWQcR5oKeuhKEcDitFp691kn1vNNkDBEaxa8VzYrDxIktqZn7jq
8IUvmdPl8XlpNWSMLXN/Bx06L0OqROzImmXTLm2i1ZSyJoBytvH1NZrha2ze2rf5
ZQwJuJMsrBEI2P6Q+W9qsCjjbsJA9S0bY2/cB4U3iEBKUuVK2vvD3MW3FB5yWmUT
Of/OQdtqolPO8vE32vpzmJXyjrEAxHwxkl2Xp00cLR8dgb0YyuEb/HORZPR1VPRl
akZhebj1cRQzRHxblOQUXcHiXFY2f3FRfb2wXYj0rA1DkVrgLdUTX/6w4sVH3UoI
ROMdkzcOKHO07GEVIIYRYDA8LZvFZ6kk6mAZKQ8PgGeHEhR2gLaKdZQ9KnusZszK
fIi+Vi0Tfq/7vvQag219cBajFb57r9eAMUWKxGAShUMSDGbgVzd3S+7KIhK8+hRi
nKi6AV0UZaQImxAkcrNUfCVgkiBaRRZEBafEjEdZUEClUkoBaNDdW67AIYm7wEWw
fB3X9Wg98FZNUXzlN0HhAqT4Jb3fxySJoUkquAmVzo6H0RdqPSECTQKOBt47yPte
qJ9qwTvxnZZ0XD8+wDY1BYlW1AmergR7hQbKBs81Kc5LXELOr1kmSnhF0nA7lC6U
n4Pn7zBcYXVvcnFca4qQuyhN7BmHGZAhrJd9XD6EqJMFWseorTG8bGbUxqJnxeqZ
Rnuj7XJrUIy0bjmlJ4FvyDjn0eNPtE8U+ZbOCgMJRrIQPOuLB3nJoUJO4Q0p5ZKl
gjv/FjYKkjAvkIjqpxv3pEEdYejQeE5FhP9i53pCEoF3zNCZ7JbXFEZqT/DQ4k7n
ga8sOtcJzFWYKseth0hrCYziDVPkeVvW4xCQ1GnXlEFXfmun0eobemLHfKtJImKW
0+uURL/W6VTp6Mas/U7PIjBkBE6Tjs2irP3f8ILixfluN5JCAIe0wB8QbH/9jzom
0A2IwfYj4dYnVJ6MKjz0k0BOGQcppQCDwIAuoM87OFbJDbgDg4vBfMz+s7nl+Y9G
SVXEiGImSeoT/TzWYo8sfcgHd26XgPGHPz3cdJRatuPVzd8Tb+QCJCGdPr4rYza7
ddROCOpnmQTpCiRa8aZmI//M1MYNw14HL5EFnsRF3kKEnX7DvFCmgYn6L47A/cjh
6yT2e7fFJHKuSqQjDDViy9/DD4PmfZEq4Y5qIXbaopSPwpwoojUU7YCIM3vkwUwa
rVjSmvD6B79LoR2MTdGFxWbdTuIhpT1KYkJpAFAQn+V998dq8B7rGpx14zhHeJd/
Ow1lILY7tnbKTWW9sKyxaDoljxzm0ZWWtGFiJmYVJFjmMjRSz9kxn7Qy2YNhLNWM
h8M0QPdBlJfJ1+ThlsShbg82whDB2Rc38cJoSpiqs2RqCFLYOswBn0+H/PBpj4eM
oxWGyw5EpcKnddgu6ddzp7BcsM2rznyyjYHQ70ZQRSm5Qb020ohwlbjAhG6n2ELW
WvTOj3wezRDR1LQFS5n8Fz8PhdACFWZ1bRbq/tpbr/+zu8wXV7jFtiPyorxFXZib
FwnoWH8xmuwW004XMK+vEgmJxVX/rwNmisCKiIzvTDwRtNzrNa38aCWUzqOD7h7F
K5AV9s7GVrHEQoU8nbfAgADr9uUL1uuaHWPFJApFFKvd8EQ1rrd5GWxBFuJ3dVpD
xl/Od3bZNk+RCNBlu8cdpWB6QC27hKaMK9zDJ8F4B/i3dDdIM5d8vQC3uSufk5Do
GhSfOP038djfJF+fZJbBVTcKr4l6jPsRdlJgW/mOfXKXYgelj4Wp8sJc7hbrxfX3
pcCUzDOh041tpIVSR1crWZfTh2n3AcgptJsQKOPsL0xza2UznvabU20Jv7/hFHyw
x+Vqp/Hn6LllUAK1CdF7d4g5y03PYVKtAphwVUOcSSA72tNx4l7Df3xplX3Le7Gz
GC46vic8yyy8MDjw/LdZpeEiiy0FXNi/eUzHwHciqiLaC47u/KciWVRS4JulCeIt
moWZ3hLWtCpYr2EIOco97Ay6Fldowa4jzzQgdQMzljWpq5FfB+kQDiy/wIt8NqB6
NNTlpnrFQjadMwxiBYHCBHZ5BAJh4QiBMdrDzZRG9fIweuk+VNtvVxnHAGPlsovD
lNhqzVQ9uXqq24a125l3w7a3QiRwM60HLDSFktJMtC0K2rsd9aq6YDPAET91U03I
/1pgxnNMT3GV+3vVQxO2JyuRu6YZ8Bp87pvTUCbQGNttVdPrFaoMMoFlth54OHQt
CQVd3TdBieDRxT8yGChC76F6aqV3m2j4fzo8QL9RdQYa53cKam3CN14tPPAemCeT
IclEZR7iOgxJS7wyU5RIi/2tzoD1LhEA8ZDoAJa6Bm2SAkfaDP1DLijyTrWTbeDV
1cpzVI2epWPRINehZAZAhkd5aAqgLIke2CxpzSYz1IsVfe14KqlxqvupC2KDPNpa
qb12crtCvyEaIVl3/3a4oM8ft/Dd9wm+cXqS1vbPx84aVI37ooCliuLgPONion77
xC2WVjy8/wYWMa//9NJ51a3UJWUhgtrNno9yvswwJL2a0wC0QJ79VuQ9zeJQyiwJ
Ue03EEkJq5RduwxgnScfEf+88NuWcQMvc4qV+7yUZtQvMzTTFKzL9zNho/UvnZnE
6CQbNEXNXbU58/YFlWwnpoRLSYTOZPMwr/i2423TktqcfDQ2KfeGckdCAiv5pYdG
Qal1hb7ScU8D8K7/JNsb+QA+jj4t2io2XVbsYAIeNgeZnIqVtWOaCdSK2VnyJv5x
c6vBZ1q50951sn8mf0Fl3OMBIUO2KMjUjA/O24iSzBuz0Op4wilxaYR0sLBzisZe
uzqBQKZv5ERFD3pavVYciPI5x33UcGfPsIdFNnTqShe8EB6CcMzg1c+xuP8cpsZu
Szn97NxZso5/ROKQSEL6rrJEgJ4cwSmblZaJrmNwY4d5jsLRUal80UKj280opVu8
c92rvUwiOpzw1UpjqjKc7AKv+Q5px0SHnHc10gPn65DWYWaHTOLYT+ahjzGVhdKO
tnACqsqimxHyASB007hQHA3OutSCPecINSAV8eYt57PtWcV6lUlb6TPBWOznl0dp
GlymOtq+StUgr/o8PZBSrfkmU588aL/pMcCH1jeEOiM28bjhiC/puGwoGie/NjUO
LHDJBxnSD06Vs2B0vvnoavrZnL2iCHsDgQMNfEN3K30l84t10OlYmqafaKhRtGuc
aG8Jgk9lL48H1GPVWm6GqA+Ev2KugNQY4m90TMd+Pvz+VH1b14swEe3xbWP6Emef
SK1Jq9L0MxFQ2gjhk4KYEJc+QIfhOYKp4/dWxRhMwljW3Nxjbe5V6JwltRZbXEY4
oR3FyUiCOMiGfmX1+lNul7dpZcNP0lvJ7EdkbJYhMnUD7jbZ44iISiFFnlPZ3ovr
xtbwxl+vL0BT2LfUyIoO2gsd4k4RODsdTL78aHQFIm9yLD8W5s64Ifaa/kXWICYb
FBAZC6K3KIC74UG0qqji4PdVCblTZZMhmh6smFP+HKG+Xj0h5SXutpZgWO2/limy
6ly5kpSFxdvse2XA89xYKQaHgpeCTMFE5WP5l1fEWYfEFN/ko6vtQMapBALRUz9Q
GbSAke/NYGxsdZgmvZFwQNC0K2E76yKj+tCLrJwoe/UJobLuPeT8cB2GW2wkz1SE
SjdG+f/GqridvGhsfFIZVADnzN6raXeCoPViEc/pRnJOsbGsJiCHaAmqIf+gnk2p
gh3dFThP1q0/u+ylH2pzBvU7boSLSAPGhhZ/graYY7X41OCdRWb3Vjcx/9Qp34Pl
evPMbVJ5zVTkMV6zNaKC5Kmls8z+cBvurW/xb+GLyJuskN2Lf5EwynoNBLvdjo25
XA4pWqQgd18/QHvhUHCHg2DY8qm473zLlvvui7CL7oY=
`protect END_PROTECTED
