`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2spsmwN6jR+cMTnvRCA0YelAak6ZSFP3AYV/Rpa7+ImfcwqJ/TsUK5JxlBslAo+I
dBklw//5vypltn6sbESMI57htt/Aglpb/yiyMpWGbWdDw8Xrculgaoj+vhK5aboa
lo03Bz8u0rZU9Mf/z42dijSrc1I3Bw0sDfqsQw+L6VZo4QZdHJ2fIf1wlyEPh8Mb
R68Ra33rboSqmTIURFdQ1ufzCF1UBV9SLTB2vki/cGVjcMKgrjDNQ33Ei9H5k1X1
IswJHjW0fAPSfYIzVtHc0iFCiZGuNa3mPDJOj1nrEAE1jC2x7WoQyGdIhG1yel4Q
Qf5Curf1+tWG2Tyw2b/XKKGHXhrCkaRac0DwznzW1RESA4AROs+tfW2lgAMqrqJh
VBRJbj0mBJ/dHwHxD2crmje/QIDrMKs5VVDLzn/xY23Xq/bCevlmEEK6rhlYjqtA
gUP55mISncUbzsWUGxm67pw5szjC8kEOmGRVnLe40/HIYA7IhUF0Vo+WOwU+rKRC
AOSANuO7/UcgczTFbhm/mrqTCbejYCMwLNqsHjBVHUXWUqlfJIoozoJZQnLLKioX
sYOn93vDLeVOm8ZseJlDBPWSFK2k3ryICzYQnTHPBB+tOMZQI3AKoBAmpGMTryn/
wrZTT5iAEO0TuxnBN7tf+LVWlRwvKgmCYpwocUWD9UF3HFl7MuQ1GYlo675/gV79
vsqp4JsroZBZ8yqLufJYJeriV57xcZhfqC7eJ+t+r6ITRgHtelWKxFa7Yr75svZ0
FQ3s9xS/Db4Dx78HIlY/eOudii8o2c0kHfACKiE7Gj5kD7C7ZkkPzLchSIuZ7vly
`protect END_PROTECTED
