`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74byCa5sNOlHhfNVuGX/i1sSK8hweHKXqBbmiwQ71j/aaCOzbSN/MJ/SMAPND08K
nxA1R8nrwaK/OV8F+RkvMyAjhuVR9X/AcLv8GvvtFR+1Y5akx8TdBhrmFuDHmxRl
FnSYJZpVh/Bh5al0vV+oyA3yXqQeAOngLZVrhwdBWGPR2Rs1TrlPmoBqVNLwG5/H
K2gLUQ8iB7UC6ieQ+Y4tDwqXw1FABvlDpxzWyNPjpFCSvWgm3yu+UZxFN8H7Kig2
TsV/MFIRYszPebTgIHLdYCsslV37732N423+ueu66Y1Dk+1TpBsBpbq+mx7Imh2b
WxnCVPnZo4wto+Lme7VuGqpNY80PoM5Tfr0LZ+zO3uMrJYE1rFYb4oCUWRXVnK7O
tG0PGP4QwqF7nUxl0OWb2tOpH7jck0SXu8TUDMS/VYihKTkWBMgVkyrPE+80oIeG
s+gF0T/I1eylnE9OCyieMDXFGhkmnIQxU0IJA3il/uP2l9MILW+ohDH7//CUfW1T
OsqkLP9yTEHxza7DHNLx/lWqrXm6od6HLfSsaVA1oKCiFZ4M3lTLksAwMICLDqEQ
/RzkHTYQDkp/wQqSQONxPShBySrjzL9hELpxnaDVfSyKyUhf2LIB85Joj4K8YqNY
iVEc6Ok3G2j3qTw4ULbyaZYlHyzY+lD88tg8ifyhZGf54m+6BHtCPLgE4QLD2UW1
PHRaJ6nimgM8ILyKF71MX6b1MDftyIS3Vpe/sbicIstyTcTsgBijn9Jny1ZzzM1L
UGyQQ0tJXTBIbvfg97JOrQ==
`protect END_PROTECTED
