`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rW/OJu/zSblVWB2BkiPkMNYpWFU1mBotQdEGCIR7Bqdt+UOLaPsCJeW20ICAKKxZ
+U2cszyHI1+xupSoeK6ENlBsW2QPOqZqUDmfwGHbCMRvkLlsDowBN05YvyxjCE4m
tGSLXDTBU/nM0jRdHoNns18cGOpXBlnJaL/OZtK4JEPczpr3OqHaQbSLtMgoFZnu
H/WJVFHYPyTaBcp596KcK+JiYusIQKJzumNKpPZqcDZSSSEzQ2RVrhY1fQG9/oVh
e6Sr/iB1sW0HVA9/HmcbKi7pgjRRssuwa6GWMmIUCaZaHyXNIDscTI+eaXyloI9T
LmIfbJFuCQJ8cKCNU89qSz1HHHoRTy19AzPqtcXuKjmrFwOuUxEZe7QK2Fd79/KY
h3cf640hbHdKi8ki5hUat2rr43m1iFYowPHP7oxIOVnrYuFLjAIuZgHEB5COt+lL
uH8ZsuJc9THZGIx2Rmp+QWt+Ie1qiQiSO9/NV+QklNTx3UD1B/snkKq6MNeqc04t
ItluXRUtEEB+F6idqfythBsQ7iUzf3iy05i3N2+3SBb6Zb2zNHUgi4/v9xwQuiBf
tF9bk45dugZeEwk5K8dXY0aphJtYTF5lre/TQ9GaY3NoDqbJQ5cZQLS+zbNStpva
6AUPk7k7pLTGt3JEmXXCPXov1ACPwMeJU8Iox8KpyGvfiMhaxjhPQjPX8ka/27O5
b/vgFFqKZgLKFoT77fE24w+8Ao7uH1pHv6ySbE0htvgRFeD3sPwQ1Z6rLijAFzS1
mQsIhbSl1O98oAdrt2Xg/yX9I//4YugjHXOv5cDvmbhl6QS5SG6DZWltPHZPXPch
jbnmEL57ypmlKWyR6MuEWCR+IDiKK5NHWS/BZ8eQ7cpUAP/PUVgg1greyzcDyYyC
a+Y5yFo/uFKUMLrOdR/n3nOsM6Tchsx4GlbM5pgnVRjD7mi9+gvSvZ27ep3sN0Lc
48klB2CbNfVYm3B7wI5wfEVlS4TFBl2XkD6VutmfPW0opRNxctmzmdmZBm+ngi1I
f3YBROr+B1x+1B4qVDTcyFTczYa5TU33vAgwzNB2Ns5g0JfPdnf6hcRQW2zuUpS1
kroy/OOzbG5icdjGyV+Fi1LKnpAtXo0ndmhKYlACc2SBW68F20FxPI4FwGpu/Eag
TwF9OVyTpxtQCR+ETfSrxoMHgB9dKFqDI+Yuac4HiD2baIx8rLfyrb4BoUjL33KE
lTri88z9y3GOqwTEzxbXxlyV0O2Ax6oh5BsCvb3CqS5wulDoa9cicXlsLVjF4qcO
GfadW11EpkCyrzK4XB8u2kpGSAtLn+h+zzbgDR6MpfAaFBEhfHUCld6qOeHBQnmV
S74yQeUDvIM0oEgNfobRrnnt9oxzkJn/qrzA5wN7N2Ekildp7T4YG/GsufaFNU+j
bkLysekEnd0K+VJQZ14XDbiC6/cxoVpgiQc3zcjsgPT8Y5iwkb450eoynwTDPmk2
`protect END_PROTECTED
