`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sTDfcvbNiNo54ejlI2+Q/wNSDmGqHFixI2aC7Zof/syR9sgs9wuctgX7DrnLN/wt
OFDUicTnWHF6RreDjb8ZflCHaI+d+WLMTvowszliRzwOieCEXj2cXafzLS125HBV
Dgk61bqbKfvIO9XEXYYfDnccCnaE8Atp7Y9/VP4e2zX4PUCiiLYx+U2ZSspHO12P
uUcM6X7Ieejtw01WOG5qRZ9O4F2V4omP9YLw2GmX7kBAuoWG8BeeobxjsZppg+El
aasjHl+MoPtH2fBBxOnehwpJWgJqvuaGCqtifp4+E6/2EeApwHtAjNz7GgisDZCG
PEVlMhGWxhsI3+v4kV4RRWm+ABftQTdoE2hAswB0CaKFooxtmPWJ7uJo97dLLlSV
RqfwOohZuB5FenTYi+48Ek6cvs3ylD2tE7jmW3VjlZU55Izlnyo7fkbwjIjsToaZ
ZL8DepP7s4f4QHCiVheGh5s1BHVBxLem57jkAFJfAa758rV9hBuFDcE+CskoEGe8
kaXHaFIttLiD3m3zpcEcqQiM9vys5QACXNhgqswhlgm3p6+lAUEF1ahH+YYkaSj7
wCuqX0ss4UuIXyVQ9JNhMBqfJIBxqS6AmrXoQN2LVvKyDDj+pWFHQ+4BkPmVSC+Y
lzWDwDehtPZr979Oepg/mOEKx4mgadbwQeoTN+8Byz0d1wMK47nuecqm1us8lLtf
E7nn4KU1eaGFwvyrJTjdwogUIngAYEDwFP6Dmf9slBeIgiQm9mkmoLClrTEMFtJm
/f2Yt0z5hG/ZLogjYCGbTt4FRQ8Xi9C6GbI3WMYNbZkLSaeT42Je+ZMdhoOuLFJY
pePfOSSKgfxLPqLLdtXEUKd9+QUxmI1WSV8gECdKVlvbCvK0noXiwc4AVUlrtjIK
p2/XP7JrG+eRgMpCa6qJI2zJeV7J+ZQxn/ay/U3Zox0Gtm6Zvy930X+D3Byw8kWp
dt2K71hODQRUGdZM/2vIL7bUyeM4Bn/VNmBgWOb2wm8svKSnqRG1FK/WnsdNKkPZ
aMfowl42LBIOYlBlXEY5EjpkCQT3pdeiaPv+ER0R46Pl0yzmZGguw0T3caDy8tJc
khnVdOrkgxXbHFHwMA/cD9PMAHA2MeEikfcwm5cgkM/y1ACfVeHQQRCTCeOtRzkb
yFs/5qL/2bRVN8cidK8VNN9mXSpNZgXGwHGom/JA7ErUjgjQMf6o0F5waviOYnVd
yhNvg4/aH+tTqZqeLRa39dij8QM9cdu3uCcSTLwBwa/3X4qRzK+vkoZCc0QzDyiv
EsmIALGljHV6ASaW5FuoZrnDt7zhq9JJX0Imycn7QFyDezvwCyqpgvVkBx80G0Qk
gE6P8oiNSZtUsgjpLe5gwBL2kfNEmjp89sIZ3GKjobYhN6czv/TiRNOYfUeT8Uql
N6pT03LhIHFYZQkAxsPp/l83N9jyOzhCDQK6Y61xnACcGAiySSmfcPuUTtlm/0Co
dKtBk0rByqIxZBFAykrMyr8nfWwszLYhmnAAmRfBFuuRWIvHuuZdlTdmR19VQiMH
j1drs2asB6tc3V6/1Pg09lD51VedR7oFEzPgFFWyyq2vR53U5kRN1xi+6cDlbTvO
YAp9pu8kU72u5jIWxJROLv4ZjX7/yzYQf0sl/t3F+xTkX0sQe/b/dqoWqUkoclkB
hqSNWZ50cj3G84F5nMpOMc6SpubHOYIGaAAZJ9xjgNPJCjp+mG/u8cZtfB1INUN2
7TP4218ktqDltSzqzlxdlFf2gEMLU290p3zB35CJ74ASGkAASjlnc1sP8+8wLLNq
bLGOVmwoEoeE5c8SnSQ5vipbA/0kdJUIaLVrgtZI7Pk1QFtR1oHHBKifQpZtF3Rz
1xPk+WGMhi7vWX0eF7IXL5Ge5UNn1f1rvxEcmRTbcZ8aPkg70nMmvgBln4LDkmuy
mrvDN8tiPjAOKz70+8BBlTkWgRbIPC8g/VHikdHNebAMdb6WuvvTVyMZuXEMFQ3m
rPXoh2zn0FaKZHJnyvSQuC2FhMGoUGxGoH1p0mFjCtUdCElyNI5U055asIdZjK7l
pnZ2OzyVAfDBCrnT7vBsZow0J9awcr7U5YRKNDc/tMYcrlqztKeXA13UUbAK2UFv
UfaEOX2I6dvzJPITc7+EFO9ybSwgci7aP+WeMEiho6MNvFTqC/pTYnoIYyvU5Dek
LQVt8r5XJPEro8cPnvcKwh2VWAWAdXjgn9/DAWzA2YjLJpA1QguNU1SDIVhueEdO
o/swF+JGwTIlpe2NCjzjTHmBjRLfy2fuf3Nw0Qa8focKVt0ViRVnpQveJdlhfLZt
e/vbqlCrXmuzbUvI3JgdUMnkmtvv3K7ThbcJ7Tu5F7EAng+K/p8859n6FeBwUPg9
wqsUzKVS/DX8JG2xK44/s9d3+eswA8FCLG/1EA5YvilaUIMDci0fWMDkAqaS9BLe
5eo2wV6F979fso4XM94czLbPMgKRBfwM7pp8VTBWm0XMTROJc81+Fpj3YcvedYw6
lM5uOhkVPdloPYvWFbpISCPaP1KY9Sf+4mSEfsyeyp3dOBLXkMcFAVmUNpsATjgz
POa1/ahqJDz8Q33GA0I2RqtM+lDxAcLqVpCRmiBOJSxdpRjWUX0d5XIXsauTXn7q
3KeCeQL2p1jRF95dpH/FW9GiD64q/Y8qum7Vx5h0QUu1jMtUJzMmHLmFqGHfMwNl
P/G0o/7PpRAOOeeZnzrFqJ4iVftDNgxFX4MlMgWuF5EoUpjip8EvgGCjjQPgM0dz
wDCUakCWWCgE1v5yjlsKTcfo5pptIsmunjzOskuxsJ0bBXNa1heRwImmzfBI01LK
xZrJQCFTp0IDE+fQLziGE6XjM0cLv2FlTAam6LFGK2DWzfIV7gx+j0rC8fUIkQw4
1iAHbevS4mQ+kEZGEO5cGZMDtVpvQC99WvzFl4/HFDJJFXFt/cYf8STyJfvA7Xyk
gTaToNPtqSRTlXlkLtx8HVILujutuhGtckwyL5Xaecqjylk5Isix1lfhiFXxQqMR
9pK2JqVEgXoS+DdTTuVD7MU6f2zPPPmgiRfTvYGtSJ3ohI1f7MPe93ULK7fp+IxE
DFFH178Jlff92rh+m60aP5yuTuCu5B8dtyN93o9w6RET3UcnRpDv3A7+O/sfVdkC
qfKyamfzyQDTuv5HVu8ZnIspilOEV7rYaE97lGhKTGAmgkk7Y0xzKHCEXmwbp3ol
A8fFf0tXYq9m3vjIrZLJUYX9cdcnE/AlO/e71vc5DVhorUIT2mq0aw3aRdg98OVg
k9CCIi1Y++fPLoKV4zQliLCCJmmeYxaFN8tvGcYrBgNozMHiBYOohni4SlcLvhbL
e4KDQd9eRDliZfI409Mo1QfnSLCA0I9SWZiQiNOGgwH9Qe9uuBvZy4iuiDa3VUux
qdsY+MdG6aF4TQIelMzDsdh7w4AwdTeVxdF8XYcnXAPYsk71AWvMB4rnb0JOWjz1
Wkm+wmZ1U0aKQanY73hk0ip9x7pMkvhJHPhdOzm5ifT5oVc2qZd7gJus/N4tt1H3
CkDLqs7RLJQZz33TRePkUY4EZ5IHl+Kd9paMT2s47ufdMx/nRRfUDY+oBKAhGZJx
yWjQe9GgZCWMBAHYBAPjQDXiIC8RIPDv0V1mNgxsAgPyjv1QD22oD4DCUUZCCbXh
18RhCjQPwfhwfvl9Kx0LYEqCN5GpdyzjAYM2uPnFmOL2rYAL52vS8fNE2zWrtSDH
SfcQfj5zVOk8WXFbSBTEG1pxgJiQgxOa/oe0PnbPRWK8ekDw9qBgGUytE9AeUKlW
B+hOZW5VqFTJlY0IVzWtHgQ+NHzx9mKO64M5hXUNICF2WAJXnJisywjgbUFb+35U
MQrOFzBJUvumHC0y5Ie5pHTexMA/BmWLOtXOpG4nj8h/q3HPdQcgQFSUOyGrSDt6
w/7yHYjB0YarT+2+ORJRDuT9STjZzwUpLIPr6q3DpxtKKlgUn02exUMom7qhBE3i
gh/KzRPbuK2One83lSmSvh4a3toPL+vsFj5dJwNGi9Sm8sHxsh/OTdg4jda5Qi3A
LbjITCdEyXhnMGeCWB//jxkgf3fUntXtwdBJYzp7/HJ0wpmpYUH3Arss4wVoN3wz
sstc6X6hbh3JnXwoKYiVGY6nqWUIkOZWigX3t+VFME01/qUFwcLhTKGDJZo1hdGQ
+2nvzWVQTyVJlHFady+1ndMx2wnCbgB6p3kvXbAJLi/BoYgktzuXznuQ/sNy3m3M
5RptIpNXTCUYqZPPg8L8IP5QnHP0/BWpYaCf2PrMGCg9q2viNe/YNDR999MjSKLp
hsqwekjtTLP6VQZPN48MQWeypdgk5w39gqTP2PdHXhy4uALStgLtsb6c+DAOFo5l
iPBG7OdunDKjrl7ThfzcNPt0suo1cVNSHxna47JzRDd7sd7xXgePPd/z8Ps2R/2W
56KmjTXhgajd6i9xUAPOyiFfyfIFeR15/9yPkTjNGKzawoSzG6BUvWEbcjrDnoKU
5aBCADYK7i6LBmY6rQZ1s9zu92tB5AWkoy98Vv/SMlmxu9H5uUavdFyMiT6J+NsD
81klaxMwnWjmUvwvqg/+clS7WLEzP7jvLhjCq4H0Ir6VsHmqyPFTgc1MLST/4kUr
Z5GPUxKB81pQuMVOQX2+qpyM1Ni3Dr263gAyfVPKtnrg7TKc6J8w5tp3sWq1JnD4
5EcSMTRlwlhZeXNFD8bzvNeqLR//2RXvSLBEmah/TvFur8Lu42FasF1PrZEzEpEw
QpJRQq/lmjO1CW0tn2+PgrnvpkVtwahex/vO8d/uWEc2cgsUwWQff9wlmo1OJLew
tIbNMUJRR3T7PWDWqejBb0vBO0APhX8P9+0uWT90F5rTiSIfKMDDN0CEFIrj6QFL
Jlu20uB67pNiu1AQnXOJqfxxuwT/P1eFI/2D5VqiTaHhts+pKwSXwr9eqoNLb2M8
KLZb5Fm8e6GG9De9UvXHiFkGMyCMmWRCX2O1/ebCKlVUG3hYO44FkamvSHHxMqzM
gefQnZAsfdTZKcnGxk9H0VPC0zGnvqVEBkXTbCToB1VSTb6+7MOcXg/zBsMZvnQk
qZUZmuaaXn4qXd8CFClrjpk/Ds+SY3sgELmUu9R1KeMuAi+UEE0pBh68Z3509Of0
aGE2YEdAlODpdhxgtHhHH52qPBbtkdO6P5L9C1F5jb5wUd0O6whDP3VnYa8dgjHA
PYntS5BnFavbkY0BjnXL/5OR14FVYPNLD2Mt6uuSJgz9e4NavlJTQq0aWkvn2Map
rBkbJ071XQTKSr6DkfLGbuVtnPqRfnCNykj704ve8nzGfBYY0bNl6WH3Mc1/g4Us
B7+2ZXkB+dQ1hsRUifcj0m7v/AMPmJ5MmARf6Zsb7V9Ozc0D3MZP8l2+mx1IqHnQ
b/mazapE4KH9qJ4BcCtP14NaUeSbKTKCXObFem1nt2kXvV6e6cBBcIsikr1e/TLC
7FLkuxqh5vbr/naTI5+5QqnANGDJTfFg2GE204YxDsWLn1yFqCkCzcT7iSBXpk3W
VnlGZNnsx26VptfYncXkH9XulxuVvsrAmtAyK51YnSqcIAHByHYNrmyeaeWlMgbm
na6ZjHbAFgkdpSG3NRCS1Ej6HLT7obFGyjGBRZwtgyfeJ5vLRGNRmplhZpW36b8N
FD2d95kx9Q/QaB8DgWBfbAHQgwQ3JlZNdBuuLiZZa7eAa9NgjdPZ6B/50nTpfv9C
Oc+Z6vMKewteTrQr3dq+XL6lh9ZxxemnaOwKX8rLaic8kJg6oZTqSAItWlKrchiz
jwgc5mzo4ICgyHwdHT6jw0pNzHXH+7evobnXLC1JI0H2hGMT5wb82kVt+KMDdAPr
B1q10F379gkoESLeq+Ls5MDnW/7MWtpLFA/LiV++LD9pozsPU4DB3qAJym/68SMn
oGFWzqD6RxagYLIaDSF2bsVzVM1D5rdrs+CF0/gzBSsduS7lbRQ2OiuNBx+tbYHd
Og8GsBipJTHFLSzA4F5AZPjUHOxV/Lo0gJ/PxW1o9AXCHN4P/PrV5l9Av0YAZ7hK
yQxNaIsbJHNnmEqPAYjb8kKADc7TmcGsKXFDaYp7f8lyq7uV6paP63tM6bxvqZ7m
5D8jUHPQyVrJvHyY2ubstbvnvTdneOUe2jgDHJ15EYLn1Sy47yb+NmIRWDA8H31d
ecQcQqYWXj0JXym3aAVfP38SbxkV4epnDTa6J8jT+9hdlSVozHOQy5vyaQSdWyGT
TFuYvzZsd1hjdQD7uQkbvUfQoI1bo+qKzqow3qYKu8VPrxYDRNCHTVDtGib9+gQJ
yHILJdQES53GoHlmkMKoHhhkF0AM03qsql+7MyCsCqr0O4FdH9+RgtLtwnRPT4/D
G2d8QZkRsjFpuHLwMiAQ4nIyq6276rHXrtTeJd6K9h8fvV+AttJavatdaFt3GfJD
eBgm/48+obuvtT+ZJRWZA+LwBQbliOsuZNcVBs/IOovmkpE2kEkAgjwHnqFDlvM8
0CrJKySOlcPG3aINFfXRVm6VOTqsKWTliacyh/eWBe/bz3qsmcbgz1t0CGeVTX8M
F/bXAcYqE/sukR9pcg/Je4tUuzRQQZVMLUxklbkngOXTMe8FdEO/A6bwEhrv2yPe
3COAHbxOqmoGB4v+52yZwF7ert2MiYl4bZZ4f0xkHxSIpqlU6t/6grnG7049GcDD
XhCJ+C5TEabaUzRQyxHDRpnpTD1HGOngkKe4m+1qnO/kQrTLcmI28NsNIaDo8hZZ
AD1HesuyUt1RXEc5p1K1u42r28DIasA6heuNEcPLvH8QvgVEanFC7tnIzasJrfrX
R8m2IVnn1itTSSbydyFdYS/zsb1bU+kxuFPVcOGoyRR2GvYBS/Kixe5u44DAALxr
A8MQXvKLvb6oYbea9qDjUO9huArgmmRIFjxMTmgb3cOpzhnm5UEz5Vr0tS99otSb
lmPPgAXVS08vIKG0DGfqJLkMpYl+ML1KQZMbVCxjDao0c/cColFm+8RS6FP2ki/B
0BPnAb1NgSF6PPDffUrudc5hRise/dzNMv2in9Af31CLQC6WyEvBiPHQ67KqdAwe
PWXbE/GSvdYW9vtdKLorDAq0pmg6Zcx7kPSvCdDIPOcSczzhkC5zBHdR7E8dQ/84
nlJLv30APxFik/OvnmfLBwHa7RjFR/QAZSsDg+FAulkYGoAF3z840e0QYnKBfO32
6ZKuUJ5a58ToM7NGHE6bD2umaWqRJJaKjfSNdr2B4ux1VriVJf1Y8i6UcmIPzpKo
WJ+oM77YmFA/EQfgj32T9cKepmeWavygeSKpSi76uUoQ7v18a58QAwl6WNpR3Ojj
oov1VeqKdoe/2qJizGgp9ThENvk95OI/qkil7nuBz0ejv8bVtKyzC33qAQRNyc+z
LA3YNRCNJAtOcwL/uDcVVZ7dMLz99+1Bi8iD3KOkkTS+4RlancHUHIA0f+AtOBDP
FCEDZtbVwqZRaSxwo6RgZtef5/Mt3oFwP1BygQ9A55/ErBj234dN85uszDii5HbG
eK5BVM8sJMHlK3E477xS6XT+0tHN/SFJ7kIP+TJCg5v93P5v8xQSRzOyGE7wFter
invdmVM3LXY8qrs12vZSEFCWJ+YDMo0bSIA+sQwgtHEHysaFaH9cWAESm5604RN5
V3eIWX1Viq//38pJgs3uHOCAf6+pZSZSuntDvzWDVV2g7PJ9/MtX3g9grA8dqv+M
oOatJutlMcbt54wkRKnx4ONRUcitckweggk49j9O5+NaN9ZT9bsNvUWLNlm1sXEo
RBIjZP0lY/+zsyYNGPIAoKY4gfvMH1pTFSuMa3VJbuPsJLuCjmhU8aCR8FoQqbnB
wd8cBeBjaOnhC8KzBXnpD5B4bS1es+KDtTc44MD47S8JaH1lCt0mfkbUd70KVUgT
V02y8sVHNvwm7n4yaY5yP4c0XdtB0jvc8/tKmOLiYPPip1VdmXXcbNN8OfF2qFKg
HCN6VJMjuNvEWqIvh0KfEzD+2hWRc07aU7hREAGb8s9t8ZeExsInEvdUvm5seCvm
J2p6i4c/cMM4dfOYrjCGnSjtS7bww3Ki3tJF+FPEZCBBY2E3HMo3oAqFS757aKr3
KWUwSRaHffnCGK7oD80xGqzkuBY1b5hIH00NySWUHIqne+hS81unubNIyZ2MxzhX
LFFxEgZtekJiuLzmuIlZ8obIqUvPCOuJbZyOJ4uwHR+u0P+Un7QpEJY8OmRCPeJ3
t6nRS4sdQDH1QMN6bOdFAO6cNe25t4e6KYpo8sdCWgad4pLlwLwafCpT+kUgn2cr
MqMWsFbQtka34zr4WE19/sdWFn7zaLRe+1fvu9qCrYlX6lsvwqfB4vXJqhHDuB/z
VIoplFq6OzW0UJsScdqoaydK+1rMxirUjoUMkWfpPDS2YqmlYppRJrzqYJCMtsuf
EVU0KfmQDRgo7mDxdVqnkY+e6wD2scjxuHqEKb56IIBSolFo5OnSFqodd6UNXrwO
D/hueBL7IV6RihNNtXfgc+/D9CWbv4BzsjEMJh2T2fe2WldmYSBe0v/IJNrha9x6
w9D922aDccfIvQg7Eay3sraqAa9kTKyk+wscfQiBkMwI5wF0OS1qKCWKVpH76Unk
lD6l2VoQjQcFd6M3yWEbhmW4c18wE0Pbbcl1NBUSpUdI1bQznrW69F4dsCsBTNQ+
SQ8S3FlhqnNAxQyviZHMlCQj3vK0w3XFA50YMrfcl497y0l0zOvu7hVjVH2uEXSh
0abktpxFa8N9bNKfTRCzR0j4fRAUjJrTSVoGA4ROL+2ZglvQh4DDRIyp39WRj7iB
rdFDZJe/8pZ5PzpY+4k9Bj9qU/Fy5lUg+UbU+10/RraQTHIeQF336/do+5Uy/Nw3
rks+jDvsPWwL4AQ0kx+H3rTRX03UBxSAKzGWTVcAQ77AcsjvjHM1je4X6jk+r0xl
cBGFDNm2ppRzzz554YQWOyHQK9qrwZZwJh1/UtKvbZkR0+8o/eyjJ3S4Momsp4vy
Q0N6O5Isp1c9tzUChClRAZbaAh52HsdUzV8FySqtZnPiAtdZnaFuzrHGvAXifErb
oVLzikLOkM5ncJxRUDQ1B6l69L/L9ywVuSBqUPNymrCmR9xpuJ3MMvJIsGP+OOWa
+zsx1cGuzjObTFMaYFqufC9r6gfBy2/90hkMPkDkc5RHplezIWSURLUWqbLnyNVy
+/KkKBu1vpGXYYAtOxY1Vd75OeUncMUW4RGSNzo4EtYCpteXDB3n0Ugceas0Szue
PQ7Ft7cjF2ckb3SKwltGYdrrqh6yVFlBsHQFknePa9X46sjIUt3IA0HPR1yLPGJT
vrR+6hIhy2QcHHS532EjEIlGbpHW60i/+9bv3uygYDciFe3o6p9MZHw422v9ea3A
pjnyOz/4WAsje18ObUnXVJF6RoPAWkS54rn8tWhpFM6sqlla5fixG20feBBACXTk
XfDkDN+GnDyuZgA32/RKv6/7YHnGHONoyK02VEcyAhvns+3ID7/JI7tfQ0ybngEq
wBWrBJm8S9Zjb4Bji6xTwwkpaZBZpUWGEGGH0JuCybaDldA3AUxKuhqv03uyXddd
5tqL5m/+Etkf08og7oC82uGTyvdfIfzAaPI9z3ZJNalNFBondnDdmoRWHBMGY8FW
AQVPYTJSJ9jFHAQe8ArjQruICTXXHoUd/CT1uk0kjrazXUvSz/vvp7OCxvn/3VKl
bXQH5jutu+RVWA8/nEpu9huW4OOA7/onHWUz0xxnJLrSMtyf3G6DFkSttgrrZwF9
LVETHvYRb7biyk2NLpglsnf3uV1HOI9RUx2/odJMqQ9QBAxe7TQarROc9wN4hc9L
q88mDHR6xi0Fx8LVWe9daFuXXpiXRY6GekJpBvZG0/ITzCz4oxdsYozLcaIgCO5e
I3nlCuDO6duhH9V3S7UodR78X4Nq1hY2OuhXJ8yJ8/grvKBpbuZOxtyopXZ2dQzH
tiTOvxmmidPWHtJPRcKqFUPOmkMkpbgsdgpnasvJEdf13Zg8vqA9zDfPSpQ+yZWF
wFkuu5scUlZH5Vv6zQQVHRSvNGxtoDhhq2MJeXOm8wGulMleJaMu7uXY1KVUg351
slEmKIf39opMhQxPD2HU/6+d9/o3g2tRP4pKhbLKYR2WjSYFYtqfJqTO95Grk+uP
e4uvwBC0egaxx/0lMfw31gRzQGizKuLtKd7EfrsCLLWCP/bb4KycP2TJly5sa8/B
liYHeOYQzqVBMY92mfoDDj908D+N1T96s3Ol+bC1MDlx7+aj4SkCpuFBOA5/er4K
ycrV/vBlhnQoxg80D6eQDy4nKf/AwTh3zIUmka8w1L345NPBIYNzTj3HJVwzdSmP
Md7MSB1JCdSqfAdLFfphheaGeN0AT6HQLtPRbWa89avBqhxW8XlbUxtcDQrvQy7h
hhOKzvMtG9/NDgwHKbmT5rRk1YnzgKcvDjBS10yGp7ovlhowWJLbdc8B2rO6WP4S
Rb/7Va85m3FnOgjpXAtbpnTr5rjuluEeh88R3TaAH5ibJ+2kS2D7H5V4hX49y363
70bTDucxL8g87fagCzdBrAcK6UXVS9oPLOrnUZc1RFn/D9oR8Zp1vSv5J4+zhbzd
lsZaUOe+QXP4kpRGw4KF2NObnLrskY8415EnePai81XrVM8AykvWaGPpIsorrQOR
EgjKdiTWfyZNn2abKitCkxV2XIAUHPnV0TtM8ITriZe7wYXbbbklNMxZV+JdkrAr
ZlgmVI83o8OAOw3KmJ7oPPOJxXooG2U/RkN1SjcEuFbCBWOKDRlXSWhDPpHehvL4
J2lhr2CfygWwhS2KsxHUMblnLCaIJkNaJ9AoTlI5R5rg1A0ZTVJvBvHRdJVQUehB
U9AZad79up4M3dfFhcrph5f1a3jXYyfrvirRlh0Vy0CS027lsApKgHGXU8PWcTqv
w1HuiFIqXLA2ya290z083vcWWEzEmst6TJbI7G7iSpRpkLZxf0msckQPur46aoGs
dUV6J5nkPhrlgscJufcZgZJdBSe+IL9wFYLCdYJHaRUhhWijVhu0+Vg+sbK7GOp1
zkw6yachmBp3K6honl00Kcxd0RCq6sBfOFAgrfKAfhqfmo1GDo4uIecSv2nyKYKR
ERvCfuI2zsWUIdKDlNkb/BwOTH66yQjSBhKwXj/sDmoLT4b/a2LDEyQZCpFEsi8s
i70pfnciCSscVUnm6Hfr2MFs3bJhcfvAyT+7hKMZkGqYWn3Ir3JW1JfIchAyaf4E
+fFclD2vsrzoPvIygosfv2Uz7dAp1N4Kcbw6xZuBU38FQmrFz0DEhI/ulwNWsmdg
NZDAmjXc/AYb3ZBoUo3emZcbXUsmJvx2MohlwCzpCCeleOZYKPc48k2EteBFjwzK
QAzlJUYGKUeeW2SzauzlxuzVcjjGs03OPKRQgnEn2TLlnTOzNkZUXBkxAn4PRQAS
VS+KvyqSMYrlJJeV2RZPw+jPM6LCKIpL8VoW1tm+049v6lHVV2yZoDA+k1Wc+kie
pmyQ41y2JLZIw26OxU8A6jtcXkSXDHg/wgmqShcSACeAZNYTTJm7CxDTK5SMYSqF
BZmtxncMUi4Y35kQ4id4u4wk9DGgCDXO5ZfOVtsWxFWmwgTVYXFch4BVSW7+QgaH
kU/hWh3mWTCjqBCmBpekMrNNFFVPkil/8sNnT+u73R5YCqlyXZkNNtyh6YaBGaTy
d82p5DWKt17HoSl3GShLXtA9A8X1aBSzitwH3Nd0zvGWC2sMqv+gYe9mezZQPeO9
Cvirq+/f61unYeDqm6o+aUgDj4QKKeWqtS/ay875ZIyRZA0LrC9WCXoDbirkEy2M
e9fEF59JDfsqFUs7emQ1sxjK6Ij1XG3z/PM8xE54uCuzrX/G636x7xCWo7OOzmKT
ha0M9yA4B2DJp94qTQwdZjj7wggoFDNE7P054QFi5Ylf2nFHmLPTgUdarqkoZFVU
CBcPPj1I8Z35RppactgoUEKdjYze1BOLAZEJ+PtB9vqAtBJB0pABZIta+qgzb/7Q
EBuhRi9rBdT5/+6+yT21hAOMvXy74GEofSunrj4vuMhCsMghUn6TFyunNfgaDvLW
96Aqb18Wb0IPkoUK2MLd3aeLnF+2QtyNV6sJzQebgsG7JGqNq1kW3BLPDGRDtAaG
M02i8eMPYgI556gD2B3O9/jWj/7pAnigaCT79e2EYfdBLR9DGj6GcxUv1Nez00BQ
EcNg5kerjrwps6OZo73CHwrzZZxwJsyLT2cTv3yS8aD/WxJ5oM/JkvBzlk9oaRl2
q+7f4ip/i34IfGFoDOpbq43caIZ0opzFFKOCaf/SSu/0sxak5e8Cb21u2x9QWMLz
RxOjGC3SFrZ37aIhVtWMBeRx7An3FfzMB/E2VAWRNJQTnoozcdpeqtLQlEM6QlEf
zfaRNfxVqYSaB/QqGSNQJc18vCXZX3hIG98BrQkRqc8EesXz4lV3bR/KKrf/409C
NvrTbdb9WQCMQm131VIhtWVTEjpDFO20iVkQnENOQrCpn/+zXrPZBE6wh4VqZwNA
N6zwFVCEusMuUW9GAvFVD+Eavi9XYH9AHAEy31VZG1w=
`protect END_PROTECTED
