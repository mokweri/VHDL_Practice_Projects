`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqO0NQm/4I9ArXlZseEdwV1VE/SUS9m/zmXKPfsQNhCVizIUWNX+4TrEB9YLufM8
hl7u4vP1aZJreEw4YdXaFXYYwCu1i5atR147bxLjuPghryBBfA0hg/k7MFgXLiqp
TGiT4pN1xHszWa1a3UwTrSkpiAgDThfp/1D/RH+fLLHYnN1tphmQ8RhIv07TbXRi
z5Xr5IDyAthA/uRuUsJbMlBbln6dQYuiWook+mdCUsV8YMkqhzXWCkF0fr47oCe/
n8SKblmMexEggE3zkwVMoKG+kQ7vVvBkM0AmapwEJ9aWO+3t+5V2XuHwg6WjlmLW
+KR6Dt9Pa3tkrNJQh7eVDOUf52FF/oJkdFdldGCB4yJdKNfW9qeuJHpFGcIlb06m
GbK/hinNQIKq3L3qHQxwRF+LZgJjlBaO6rXFsVPNxuHPz6kkEsxC7k4geyuHkxWp
tlxECyFlrtXTPF1t+o5hkpLiObVQoAmStUYf5YwU8Oo2PZ25hNi0nMWOjVGcaJb2
4bVeaWLVA5d65DuELDlOg9IaNg1l/5s36vo2mqzC2hUZiG6D57/M+G1Gg/BuGg40
QSp7ewRN80jY2IkEi45iRR04A7Ben/IcTkU0E2NcsaU=
`protect END_PROTECTED
