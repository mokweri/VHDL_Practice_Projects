`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RlnFyApM/bKCQvzm3N3dkDluh7USc8OVogCuvQPTbooM/lhOx2mm5sRKhZ+BPuu
qWODobv57JjR2wYVEEmAxsFO6IZL4M28xPztc06DWnCkeqRgneJ3UxwzXQaU0lLG
sbW6Yt3mc6aj8R/rtydpPWgEgpGtCuocNP3nH3epplx3+Jlq9yhlPi0MTgEPm78U
8HDR3TVOhxNIKL2deZvEPcnPjWgqtR5qzjmjZT2qAiz/9/YO/QfECOSGPtWdu0qO
sSEbrXwu0pKKovRMAyV9mIQzvEsgQYDdEExAceAThx8j5KhjmVcFTxeGAifPkD4e
a/MaF/0ug93OYaoTM2AnCDQtJrvn/eGtBh7borZBTAa/q658JrX59FG+0jnrfo0G
Sfy/d4sMCMIouP7S/s5e/sUE5/WPdVn9Zhph4oKqBGAl+igV8h2tGS5ffXXBSAU5
0pUYJmaoMsJ7+XTyptJipm/n7ewBOZk5ZOmjNe7CMHaR5Bx7RZBUdiEHNY4ev94N
3PL5za8633qROKUy37C9iFFYg0ZVOzdQMer8dAaipuiPgke/wQc4MwzEKWXAmEbk
fIN9eSLi+SNpplLoQxKr99wMIJpQQ2qzEcDvX7xpvbE6G1UMPVsRgQp1XPgWalLn
L4jtsxirFTr/KBihAuBb/9EZQBJU/2QwO5uiOXYLLt6xxloUn+KR50b3VmZGzIU6
l8S4R4ZvzMX+AKbsIPN/mW/EXV+xjE4+cjpuq3zo1oipqYPJ0vo98uCZTszp3RcD
Q7fGRsxcBwQad80mPB30om+0EekPW12zo0KR4wTfaY8d4Ow1t0ipRB2O9hu0EiJM
xaGjYkzyY/oku8mWRMtMt2ClirYRn7f1UhwstcHbzWX/+sXiBbh0ZgWpUApz5/cq
kdSkQ37Vy1XMqMz8wEFoZkPfKgOAlwcoH+fid88GQSlEaFnWAx9lTFW3nEzBwpUp
5Hkrpe8wpnL7yvjM9En3u+qq4eM/8sDqxhVIc5tt/J0kMxavWnSNyzaMiK8nhSXe
MNEB90ai8da0Pxag8cbMbNUigwMzs0Yo1eL6p97RRAH1hlF93wM1aPl20Z3Tjad5
7I0sH4DJakkqADC3SQewx4LjGS+6o8sxC07qGllEmmnkbaurivMP5QiCnpNi2rX+
e8lda0/jOcUv4F0JhWRi7jUlMQnX7qjBlbHTXnhLHQTxnkzEuWyXpq9OgOUK/38I
A3sQQ+0H9wRQkVwx7CzJF2VsBc9EAMXRKjEeXb7ANEit+dJoultS/Ca7meUSLn8l
3H1lsPXKXLJcl7+0LlfOgmeT3i0+J/kLPM3v8k4kwcqn2QYl2NIIKtZxfVePjiTJ
/9NszWVzUjTxBCN9213h+p/3Q0A02yadZD9RhywLK14ngX7X8eHd4ZiZwrRMz1p8
BNsEuEAE29+6hA6cW/TVDbq7xHGGd6W802otE0P/8hw+H1S90f4CpgZ+gz29z4eK
rkGZ7bMdgj9wXxsJSllSwSBFHBoPtHY1HFtY90/Klg7QbN7kEcCFnS21izMUU/oB
O8kICtIR0EIi3ITsv7AeLA==
`protect END_PROTECTED
