`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QaRIt1Mr1YK9qpa2CGQ0LDiaT38WHJFztf+mtov33ysLNA8YuuJTtjjpJ9t5Elb
TMGbC6MNtKwFMFEyRt8QZQVI+xp8t1cJe402ul4P9DPltyy5Tdbv/BrfRCnGW2Yz
1AVy8QkKbwRmW6MdgigRu9W9m0N5TbAMHls8YdrbkMguFFcAqTC3koaRyb4/lG5X
LUzPtbDTHeoFGbRrqah4UK3qRStfaiQXHVh4D4hr0KUkvvnY6kkkOqRiH1W9uavB
fjx96LqqZtnLIVcOFdQ0dFDAbhug6TpJCS2J0gU5ry5SXQQOVYQ3z8aPlnunAvpP
UYwXGk+BS75NX/BzSDUhN+PzEo4t23V8kbsXoea2/N76oYKS+ammEwlXny7zen2S
iPSVPIqkXsNashZig1v24rvQcVIu28/c07sVmVfA6FTIR9MejD9LtCBnyQT+8ifP
SdoCg3vGWIxUvBiKyEdb5ZB7ifFOLE0Ec4Bw5TdEk3ZKKlrLOFq1Zp2baarK7xBc
9h4khFYkY2juO1VxgnYeovAmcdXRqQwCZoSB2GFz7IlnO0Zt5zP8S4RJPWEEQ6D6
WI5t9Rhjk5PlF8fiB4Wpq2F47eGSuaP9qWYdfhCX/Oni7htqpB47at5SxWQ9Pz7H
/FInbRNkdTomsVKXHY5qLE+4Cv3n3HrY0lJhoI9DCg3suLqxPgO4rVJfpjNMuEYo
03enzFNTKDlEyy9MEF/2c/5pjKKXdKY6zvpqDehUXNaJYmc66hOtGwCIEq5el89v
EJ6x8FmY2vJtQ/o8Mnh90yIifHnBo+GFdNUmCZii9jCwtzTRPJvL+Rh4jGNRe8Qg
v28zFh4PSKW7u4j5AXmDBOgFf4UDxJMhN6Ebr7/yjR9UjHl/dDEJqh6tlDcdM7CM
zHiP72JeAh9eMlpVxlOXRd1z+/C33yA6pDXKKhP5D4ZJ38JA7BYov8Z5XhIEVrvO
ziJt7shIsmJaV+1lQIosJOEAL1ANzyIHAmaIJlIRGimHt+MAPeopamRMwa3dkvZk
UkyUa1AICr4stsAA6jWBm8jkQBP++SMfpzIyjPvFULA4lIS7s0dkX0iUoDM2iI6Q
SbMb9furHnUbKNohSgkUsG9QhO+BYTC1jkGNa2Md+R1Kpq5t5MiGTz2lU4CxJUli
wfpY7gEqc8bEOq2TWob35kFHcMNEGiNPQSu+oC3Yjk6SGWMF1EDEGyiiZd32lNNg
Qp8NiW1mknRFftvWuyRJTy7D2qKRkctEXn8VSX3L5Vq7n90DENu7PDY5/xUAb0RL
ligZZey41PeVAkjrwO5poBsnIv5ghBpQ8vhdkOWDDxdGAXyHFhh6Yf0NSnRufijO
i4dUHuL35ANDGSR7ohYY99hsWu0Aj1SVDck/onR3Cix+ONdRIq/Hd07RNpTKjADo
gnBx9nW5HklTjOcBLP24slkLlEKHo0Jp8fMO9rhpcHqXPo6um7tWv0QuXtKe4waO
MStYaEkvz8+qEBXfmcJtkhVR/vR0wAGVhdqwegKmILkpiUPoa6hQmkX9rd8hop2h
xKPG+AoQVWsbqIww4ceD81kor/Pmymg1VkkDHHM1mOy2t07jX/cnitlvrCtjkTB6
5jfcqx3aufbZZOhphxzctea5KUzpD/HWhRhEsrmRRxox+j/ddspr8kuPCk8KHE7W
vl2QFj+Yha7EAemsmN6MEuq3AtEFXr3aWqcKXiDEGO90T86T2GekXDTYe8eMeuyj
asaW4T68ocaUZvZK4uUTqKV5t98iuNa+qQhj4+m/ChSsaLbOlMuq0qjh8Gdq4XdX
YJktQqLDc+TI7yYCwJn80NQNITl3mmZDu8jbEgrxP6E+890Tzv5yepL/GorUMPZa
1Dp1dJ+AEoeKbNmL2u6UCRUxyx5DskMOKNeo9yBpVyIqMIU0dR50WB2k/V4s0Z4v
+OWgBVjyOfYqXv6tU6iSsNa92m6wCRGlNMC+jYFf92bNWNDXdQu7cmhDqT72hLZh
IA8H2JFTF4jR2RqdGj8GX5ds00icONk9ObDgLjE1yPVVKp9iYOf22weLtY7LxLvu
3HKiBGv9aaU1FGO189xj7AgRTjwJh+yaruF1xCEzgxTDs3nIXiZ3et1hfGUDCYZ5
zIutbOhgYFwsGBoyfr3ZFcRET7uyqVc8dgAG3Nnuwst10GqIcgvN0Dd+awDUcV5D
aXSZQVwfpS/yaB6dRhAHWPCwI66eQTw6VQ/+hcVTxhlBHvJfyxckoQAyq3p9z1WN
d2+R9uTnnAWrTvtAEZ7JgnqXhklLIWgN5/jmzZRvpog1VdBqJFqrj8MVgSx4FRUJ
TMAn9t60F5vV2ZXGEeG070mHeSfEmnjJIXPOCH3R22xVrw6dB91DwALUTP/t68Fg
KTkglzItztks73v3W8kmzOIy6UFviPVlZ2OEsIgn7ZmjqCq5XxlkYuIEQBv0kNd2
JyCGytaxgqVA9KmTarjg74QnR7WmNYCBD0Bs9OPDmWYBeXt/fu3r+TyGgpyTPP7o
8Yvl6vfP6amA5rz+Cb7ZpkUALT90idDT72Kyu1iPH9UNf3me2a3/kXmiAPawjliP
CoiSOa8d00n+9JYfStiYIiFOxPd3vqnv5cZVZT/8vZ+HTyA6IeonzHx0Os2mlDg4
ElJcDPg1TkX/yQ3+cYL5Xy0AEzUmvay+5emHAEdO2ozpISpV3tXGW9c9KH5fyIPI
Ikz+RG7Ho6drDQi4Ky9TH71p2Tyka7xDNEyq++00nw2MYLFJZEJXI7u6GAuO/EEk
vNp6JFkAl8MxUqVqieRPClikkwxm6LnliCuwsgpv8UwQWJo0YU8K9N/z9oiCAxQ/
gh69ctqa4LIxsxtLK6MbhfVEJVCngpyBD9UMI+Y08RVsNsNxw7342kul0a3Kflnc
nmPiABrAwlp4nz1lwZhEd3wSNN/7Q920FkEQXaNtvRBa9AMP9bEhC7/lYkJPFZ6G
A7qbs9lp8F/s/LNhY+DLRWUOVFDox59ActCiIX6XoN1XnQj2ZkM2j9+ArluIHkNC
gS4fhb0/kUeb6JDDwCftyi2lyQhwu7nuyp9DhAZNszflC69lr3uNJ8dKvnxxB3sf
Et4dHLnkudmdmlirtFYz6FOgoD1CGwPrgk6pl24CoBG8BCPu2lGfyzWQF3amR+H9
qw+Opd6MstetPEW9ukcWRpujKgHu1bqgl+1qfy+vjZGu6rjqj/NP1oiAoyINCEM9
dL79RMMZmtk1FcsmhQfac0iEl3o8V+DvDtDuxB2NxIRbrA6QIv5yPJpnKlvk00zb
N/q5C+vdD7uWZb2goXkZ8cGQFKBSBsJNdAg2kdPoFxRbu2dzztBhGiENK81+pUmy
YMmCarTmvoFGmGblIqWY3B70avWA6WRI/CugH3C45Yvvkm2BvkYdp1ueT0jYyz+1
S3lPozfwYeY5ZtsgG/71j/ILNRuqp2f3VDeTzqU7FBpnJ1qB8yvVaM7HmAeGYKxb
GX20N0D3ll7D/5eaEtN9/uwZeAUNcCqIj/+HoRoD43YanMK6GyaMIEswV5tH5qys
QCXY+ExFE0KBwVCdEtGt3tP9wYrl1428tNZqJKB086a0DlvOfAGb3X1kciYg0M6V
we9IdQGDt5snpL8vmwxLDzFHX9Pqm03/sp1wTZimDzVwtd6eKVoZRuJEiSQX4HBo
uQ1dT0Ya9pfO33tUlHtpqGOycvChr1+aPWvs9JiXswn+mkeBtz8IV+lSm/0ZkL5H
3B6+YH9W3/yrKcu7bOCGk01oUe2h4B1Bk4+HEut+Rqr56cJ3R9YS9/LRSOGbwlXS
13RAMR9YQ2fG0dX9wfQzKIYowasllcNiSEvnJ+Hx6XMGgajQgDKAd5bX/7nrWt+x
5Xtf0yQHZM58W8wOiiXnk7aZYd0N69qtEjnEXVf3YSNeRaOngTS49zc3Y2prseil
/IXeRzNluoZRoNe/6x3VNJAdBatJRoGh2tKTY9TPJ7ykaNYEuPuAl8DlNbXQfYRM
cOG/6vsxIXHomOg+8eOJHokFPROvCgQOiyPfpsr+1RH3mHPHZI1o9mnV0v6iPtlK
DttSdgkO/Xo0ZnMqurcV6j2bhE+BHZo8hRvAmJqQ3EPNQQwi++BUT+eTs3BiO6bg
0brh3vgBpWu0xTbe01g3FXXA4DUKrDjO2KNgrEzT4bhhi2s3l0y6vvkYukIyWr1U
WuC2wRkz4n8XM/BccC0eUqiTnE4X5yQfHkwgKpacUpwr6VlojYa5puNZ5D+iOd8E
leKDU2bGjUoj4tqVnf8HuQf2HUNERKaRl9n/rjKPW0ukECX2x1pzY6dTyclCSZl4
rijGaNUjR1/sinwqswOq1IYPzeT7fp9XVacJC9SBZfFe146txUEQZuZyZ2v1rCic
/iNz986ZiU4KYOgJbT3rqAd9QK1sSsxdsiQuBKxggZX4+E0H9cXabkSn2mxpCQNs
waaTGs/Z0+Hy0KVWHfly0kzZI0uwSMaP5rryJtVF2Mw81dUppSzc99SOc0M7EL9F
lGCLq9NL5vC0HpQ8Mh909XU5nvZtoUNibRXMpm0sFHTJw0yNOlD/qz5AXr5pq2nj
Sh0o2NLwQggmR4pqDkbXmiSKxbosctR8WMHpfra/fdWuPajNwFfhg0Q1tz75TTBA
ToBOOeb948f1ObXEdbW0WFydiGK2HS4zod0/qM/wLKbk3zmPI2w+/hHMQdDgKy0I
8scbnYiMYzYLZOIsBSKLb5iDFfDoWgfwtLF51Ke1Bcg+2+TKCP/DNSrE85V8nnsn
bIs2kVm652LpYHg5I5IZ/sKO6kLMpaWyaeNyOtCjeNUm377CfP652vHP6SeoEgfl
UWV7rV/759MLKy3ch/APNQ3Ztn3P33odOFg3FSW4UGqnT0HW3k1kbFX3IJH/p5pF
ahwpZOglM0H+85hLq79762w+6wTDuyQTTRYCuGkOfrZ4QgqDiRwd+Uov1CG03aRn
z8b1I63CCMWyXDXmUn1V692pxSJOyNMKjXqKB71JmgchqJ5zCMaiterHFTBlcQD1
xu+r/HOrebkkMkbmC0OeLgUWgeMp6IzMwTneodbhD8lWvE5x2y0lbWQlmt/515wB
uSTOsOO3gv1df+rYPdqZ4P4Z5v7IesgogZDcO4iZ29sxUUWsOqukeVBQbFdjvQAj
VKpNAitNpU6Om8lSqCu6TmktZO1DMcDoItKeCZHjp2tte8QoTWqeQ/lz1PXIfRhg
XMmfmzKypzjQhdDAoIX5aPiUuPyzzLRDeGN33mHvg4LTE+vOHUWdjFoUpwykA0sV
zeB4QocYJi2GCoRulhFYQ69/oy097A4+R/EFBVRbDzBEeJSeJZdfGWNtFI+igZD4
k+8vh+MGSfQRgITZkJUtyCM1EYBLtMMTiNwu7bwjVhXK/7npiVzRqop4fr6C1AVw
8Hcy31S2fp4slnvx9TsTePAst48GYS53xFVXz9iHc9nyaCFGYSqq+cZY/rCElveM
voPNKg9xvkcVdpZGQT16+CGvRNQgy45iyPSFXlPrzoLbLIeJzqh8e0XqvU7igMAE
ENh37eyo1VK3HNbpodVQxzP5kwEezJ2VSCZofQJzot4oIXTke2Xl5cfucg+0NEpo
kDvySPUfAliwDcry6h7MYsp+VMtaRvnfKy8H0fv1k1U3RZ5DrP1xvWVq9jTaO59Y
qjYbcnMZwg+v9Kz2XQWTaH2AMBbpcU0YCdnIkMCXypq4WXs91yvlrwX/Z2qXBKD+
TA4QX+NNFv6VGT6BWDbaw6hpVwhpnAKy8l6Q4cfETiz+Jvl/KtUYfng/+IYFh8Mw
XehM4bHjsHg174W4LcTf51lxKBEVuhoznT78Qe0N8puVZ4iL2l2+Hr0vu/wHp7gq
mVKAzvHTVkl5jJ3xSxaIxvXVZvQRQT5F1IXQdYb/0TGqMiA0xuwRyooDDyhul0Cb
saG+iVemq13FXxt5ohFGvCNTF0y1MNifjVq3y46NoXIP0apAAa9+vKgj2oo8y5TJ
PRX6vhcsuWmIC+MWrD6llGfIV/uffWpwLnropNmACs8oPGJmg/A+RvrIt33O/HID
jVGGoCIciiYLnpT6ZUzXeLFsJXPVje/tw+HB9Dgju//6ikd/7PGnrjIG2mn7x1Zi
fC7OpJtQ7MbCP7yKt0wfofmBkH95WCq1pRmaXO6xv7d3a4eW7vHnj44OG5roOkRw
6iQ6siYli65duo0xCrWzLOqCd9ONxwAlshar2NnxqEGSdNMb25UGDe5D9DuhC3H5
0fm526IooWhM2j0igVENIFEbUkat5vBPJ3OvbIZInndI1ZLILd46jKU9x9zbSXkW
A6TNBSM/CYp3AxAOIpM3+4QmCscTgJ3vUsRReVec2IzU6eRaNHYasYtnMXY3GafK
eNW4XS/6LRTUehGSuXW+eKCEZo1FbUcOK39YbgKsAp7FRB6yTGduKNlch7RNGqLY
ucglXcet3V7IUcgajwcx1DcbiJ42O10FyH878fmtY35Uivyn1cm08bsehigoMrbT
VDlZ7d5XII6rzDAatCjCpkeTYRKMzzuG4jyuQJ2RLIxcN1IRRpyv5iOHzhP8e+tD
+M0N2ZQ78xSwBDucE3DWv7WmJRIRHKlXA3tmB1Y2Op+TSvBVG9RlFKl/3RDmO5uK
qvduqK/AhBQeMfmwR9c7Jxf2wLFtjFuCOu0EXIto5wwfF36Aa5fGDfztE9XeBAvV
duc7HZBs8f5ukEKi7c/qPDzNgSstZmPsEJhXE/IK/AoqKQcDGTm9bYLtn+/2mDkP
rh3N6ORsx7M10mC+U5+4eVMIKJwMK3B0PBxK97l5W9mxa4rMOhOShdBt/d20uEJP
3ahLNmaYE80MUjjNfjWre846Ludtx7oJ1Todk/y62CQIDF3HwBZXjHolKZOZVtUO
532k4Eq96tCAYA1qFimf3oaOTVlEg7r2+En9QE58JBatCuEqdEN3P4mCurPhGJlt
+RU6hd0ll8g23RxIlv54vsw+FBdQyn5AGCsk9IJAMnY+LBRP686owAW0sWk9/Qbw
nMNo75pawEbNeAJBoICttQcqqLjF7RFWNPBHBI5Jgi5HTlMVn0xxdFRW+XNqkk3N
K1g2CbIuPtkH8nJYakTgBX067UyF3UmhGttCA8ivBiy0CRyRNLwIpKTsSfT1cUrK
Ebak79zg5hCRgjZ4O0Piuy6WATT65wPW3426wrgLYo7OVzeHXiMaZMkawV4NpRwj
bmCz3hkG3+2uvakVDYR69fO/ejGa/M3qyvZVlUqBTsYjIZNuXJV/2e6icqGLXUAJ
DvgsX1A1nWAhETjq7TP1SKK0kaL2BGi/qs44NEK+FiV8+MxR3A5V7Sl8Gp0qdVtI
B7vykfMkqeQlPfX8ctVewjAJASM7oP92EbVN7+oipxqU8d9UIXpqNrotjvE77cqK
NyJvs4DW3ilfzDIL0lHtTp4FBkw5PXKQCINrFkNH7QPiUKFHUPAPFsVneKHwiSe5
tPOx7mqluXNv/ghdnZSH523cIzULHF+Mnwp59NEIZ9fRN0VZepxmWdERxKPl6Fg0
FtoTbg2BT3gWXW6FnvlCoubmHFGaA30FHfgKw+oZeBGQsRGd9Qv5elJwJhh3hvw/
zK0wpvcd3bDRh2u7vcUXYFuFZuyhnbkvGUU61zuHpazju28ejCSTvx76Be77oUFH
+I1j54cW1P7AR3lAILU3BTy6y+uNNOYhiw9sDGgp2NsWbSVns+KF8r4TgXxYWAgS
J75T+pBytnWuEkVHYIkS5kPrxVA3fGgUYwwYtLJ7mE6a7OJIjqgDUHuefFktLFan
KNCNBUgRMDomNgXH2royz1ntNSg/P+mrDgtptfHTbf7+0C1pcZd0OpJr8SHISYtB
Vcr8lRqjQgBCi0cWw7bMfFcdn5LjFWTgZ/c9mTT/SZerw6ZH4Thr9BcQPDjeFSMn
U9h7N9sDgg3ywrjwUPtDaxZAubqgvFzmJi370gzyE5ZqIn/AYoGZtiBVs9wpxT2/
yTs8RKOxUXexB3wnaByCXW0mVU4UdRg2ndq1nXgepB8+7vkk+gyhu9Iwss+eMmvD
Yfz8nn6FnS/nCIWHj1sD+fZof05+209LiXh5PMY9PZ2bwZhUqM+pbvvSH4xvZjEG
HUERsbV0ub5YJam8CdWeOc+qKuVyEX/c3W25d6sQNQapejZStjob35nJgfRlUP+V
8aastlzziD4f8GwtV4rjP/cHrDlcD/uv5XCYJehHRonIzlUPTrOSJ7oiULB/0NeA
5oPbLcPqJ20z18ywcdSiTGVL7JH9xvKFtN9jwpAj9SumahQ8iJCzqaNgBIOedwXK
/rfF1vWwJeBybrcwJ8NxaQsOCcncigi/K4ZVTFrAiluWyL5dNjuRlts15H+mLD/d
Z6ayYRhDWnDTfnN6ukQbgTW21KlygoCFuJAraU/3H/LyVIx9Wq03Q8IpiFO+Oc5p
2Di70OM3+CdKo9Y2/AzxtWcf89hMPKIFROOsWERjdD7BaurH5n0ixu8y0So4lsWQ
zenGi5PhMNyAVcT+utu2xlNfmHnzVFXw08bmst+zAgBAzwf0xyB1hjlscHtKjMv5
V66dXIT7dr6Eb6oIYqrq2+KslpB1wtJG3l0aD7D4bTiefrswuKlcfHCsE/T2TxFT
xiPPbF9VMw3Ns39al7BqwsBa1trtQhmj17DFN94LDlGE0I3mGQD8BBi5H6zD0fde
rPI98kjG1k3pMQ1nD/VKgaLdtnN6znKrU1wAk2rSE+MBROEQeFxAehDw1lKChOCN
UFFvv6I+o9rKu1oUxtLhPb12Lg/NV2gU7Ve3nN9ba7OrIkMvtySymrt6xkzfoat3
0PrwmsjmK4XNx6+541J+u9no/ZNWPx+7ADAQEaZ2Mdf/wYK1i8lz73KeIZBWSDxx
kbFmZyUIo5F1Uft1QkdEZ8Whu/S4OhGojcrLqy0EEv26EGvqWIztoy5A3kZc5c6K
Vu8gscA/QHCzM2+uuIwMW6dEuxhBM4Z51bJZFAwKg3p/QTfYrRPAVlpZ+MC/M0aj
mTDVzlMD3UJP8P0vPb+05P1yslbt+V/77LhaAryJWMGFc5bYIUxwYRC5YPztpV3i
VRTxq+pNG42fHEIukHsFjg4G2VomQfyqRku6l7gaOYgsHdE/tCHPO5nCD6Eno/uZ
2rCk5uyjdSqXOeIc8fLTSguKss3UpMIwJtTHF1H5mxhtqZIT/+EiOrjSI4hqAfEC
Db9ztFXZMx3RqSWkRtz601lgUiH0h4IZnppdJqlnqdNg2L1bdOOamvJPNIICcIM1
HBpwMirZn6KCSpEaZezstZOj0dFrbkCdEmRSqjJc9xi9gVYZrrBOdAGapnpdCmC6
/X+SZMHaeqv6U6Bysce+7VS9+SGfaRSgBaKh/PCdS6wRPXujBWTAnVR5Z1zO5NJc
rZPS+rfdcDTbJuF5Q3ZKoFbCqqnV7rk2sM7LmKB0ndG23zPxtjv0wtgtfqORKW8G
jWCX/qk22V1zV6kcJS8T53ED8RqEzKWp8N8m7A/U8+aQJVIB166Jv4fB8wfO9BKB
kW8tcZvcuuN0IiDlJ0dEpEovju1WutIfwdXNC1WIMbaFDRPzvojfrrNRNwQ6UItZ
JneI55WZS7qThjcXeHVGCGexh/bw7DxSFklnekcSf0h5RVkFlySLOQ/z6lO3KoGV
s9r/C4vv5ev1S6P2oeohJ8zpVE3BEvgvS+NYxGECp+7aY8e4Pc+btv6bSKijW6TA
ofN3nENDp8S64W2/P9dICDC7fSPCoWc15YE6fA/sqfA44f0hLbxWiySkHOq2clSF
cSajIFn/xvFByYGMV3BdVsw9kjnW8X+XOAqmAAmD6RyDscff/wPJ/SMX0hs+Eb7O
OmQYBudV4kvtQuVaNlttJ6Vb2EssLjqx30riQGUzNhL7OMYAFdfKz4d21r7dYU/m
sWXSTNigmP/n0YAQK8Dekh4uePqNdDayc64RI+YbA8WwxNF410qYp+b8bXQVk9Q+
szlJ3Du+NCJtze06c3uxT4J/mmhiN6KoI494sc4fofPJyeuSPw7MQdDGK/xdXTrr
jL1JbHCbUNdY/IBgsoRFrSD0ZeAxPqBzv2vh3vnJ2Wmu0OK/P+jz7BxbVuAAjtPU
PPj9vH981z09QXK2Cq4lo0rxbuRuobVoMSicq/QebEnxYdoFpw50vMjJVxlFN9Jo
2Q42BcfZ109F4VLjjVhfDb7FsM8yZcZW/x1YIOc7wfQa/kDY4Y0nRcF+PAX5ekMm
V9/d/Sn75Hr3hfZitQtCdR0iYUS5NrAIIM9nz3SfGVQ0sRNSPE2vC2WUnVk3XvNe
UlVT9H4HW/ePteU3c3bBbDk4IyIjzpRU2KGvKnA8MI5B+VJo6pwcRn1nGpQgT6+R
D1vnM4keZpatLEy1q4LgBZ9mxl+6pjjDrUcafQ92NLdE7PLPC51bitHMVSXe7+zq
Ls3HBvTfzTvfY0sjItuB6rFZV2HV4lU3kmNDt7eB+qs0PzehSuuKbrVGNad9Tw/n
D4MAIfSkl6WOHfLD+tAFUg7ifz+soZUP5mlSmKxCFkurZ2O+y/tvoKsR7PDK3/0Q
bpVq//WDzIZqJtO4eqxp/k+6FvrjRNdoZrVXEzCPw89/rotoJYgH+4QPcNgkpqAc
lk7Ac/d1eGQhb5fmeQ/ACP/5CiGprxrmUv4vlNmk3B/yqN0WHpnNAJWVFEhJD+3s
F5XfEGaNEsQbQYYkiwSdHT/RTATJ2+mhqNfTlMW0V6NMtyp9hjUeqvEmqZYoiJO6
dzpH4NKPIe8LCxc2A0K4EBhtMZegNC7xdN8AZdrIU8IBMroOIprIIIzNmprYbXcP
7B0eStuQQEIi4saxrLiX/yFjA10gDuwe1cAlkhhrfH8CbfnPJ4cS5Pw7VDVpXt4G
b1ppPoc7n4xbO4NQ/J1vE9smonjS91n+Ofl+/C3gb0BEviDPuiARuMVnONgSBQNn
Z2SUL9GTT+FSGnMAF9qmwyIIbIpEuB2TiO9vX1Hualo=
`protect END_PROTECTED
