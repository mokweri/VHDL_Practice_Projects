`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vk4DT1T6H2GBcILA7v9nZWuc5w7P28/FXEO5aZGH9kFPj/7vd4pQ7dsbVoBCVvV9
OQnMb1LX++x49lAluWXorZT6DyqSmIbxSJ+hSWOEMrw8D9LMoDURMuIILuPcOl+e
KvjpYMe1WEUiEJFKZ2tDFFaWu2tcziKgciNGlfogWmeMLOg1KU1B5XSWskW+TjJM
O2xEeCg52FqGhEio+LBSA+1zbyOWQABHowMXunC1JqlnCsNoP/92ADVGcP2fSdfk
ILVSDBoDOoA1iN9kdGRGj6pLl9cVGMGo1fmZpQOkrqXxEPOuryQ5x42ozp+tg+jQ
TrcJ1QixrEPmfEcy3WY7r+PjybouJuy4LlaYeRCmzbUv4cTDFgRDSwQ8pdkppcK+
6aANmnPbcP0zBuNlyUFSZ8SkWKxhiSodr9vnWQlRsrKzQG703GEXELtYzYGyGLYv
bO1OgwBlFq4/LygVFOliA3fzDLTgPpLhasbS3aUaPzRS9ZF0VujJANRkwXxlVoQp
yfH13m4GCEEbKSwWVWk1sMmOFrreR7PfQ17KrYJW+ZBzZB2imAqoMfdpsH+Jdqhq
fiEFc/dgiKHbN1vxUhsVyil4N4ByciSpAD/WcA9n11zcBAHarjkjIn3tBSSKuiij
bSee/scXe1IFi+qMP7wiKLeVENZqlWLL9ZWoYHgoPzE5fQ4v4MnxednUMboTvTpB
THxseT/sl7BthuaMkhisukHaPK5QV09EkTBgT7ImtAaJ/UwjeMg+sbNir2qL02dG
F+aIFKXetl3v+/DIjgkcLlh6UmHlp91eQ04j0/Nmnzmo/FOCec/IncQkP49HCurl
3kew1oOb8JNVKgEA0n/smlrNuJjjPwT027NsHWXla9/IwIWPtmOxnRJWfcC2t4VF
JoKs1GYthaTAGdUrN2cntPIXiqV1s7QQ4t6ngCLiYfLfBcC/odAe29aWQrC/2QBE
ypnXJHlQYV/yYq93ndaIV3+7pJdMDLgkCGuM2zizFrsevsV8gKk5H3+PhPclvsQK
n55ZMoQaCn3mJBSgzQgOA2ctHFSlkQBpFOSklE6Qwq4//DzwWMQ2lzqKDl7OXX60
jcBu3XWlYfnFzLjBn+NYKiH2PKu2znJ1qYx/8K5GeUhDwsmFhySnsRVp69JrOh/c
wiSlONPUV6QKHpjnQ6DUTGIxgTOc5E3sy4EIgMWxBTlLB0hpTymxrdfgq4z78Ok9
44xAR1aVjz7Dj0sox57BqePPvMfHg/DQN1QXISKnfwx5tBpGKcu2bKhlhrEPkL9/
4mbpDbq7MU0OLzemSRoyq00luJCCYjLc17/MAZ2z05bFG2hqTrghA3n9qJupUHI7
Q8w5ppi+ndT6LDpSw38wQKQoNyF29Vl4yoQ8m4Z8MGDSlDw8NTb2WtYLpkr68ZpZ
V0JTtsX59/fZvywFZbJ3rdMQi+jh2K/kB1DE3VxqaRb0kVYus/4txmZLxbpK6Pto
Z7cpv7H71kQuQ/QZBdIFTLSlVrTspfdgQOjEua6vBcFMxEgD0XDCaHKnhgNLaFQT
ms2/v26LSBjtWmG8BpsxJ20nYR1Qh9xz4lTEM9RhnqG2J285sJJydCGxZ0qbCrnr
NtuGgTtlV/VWu8XYNQ4bMpmk9jKoyhp/yc1BG3aI4IURoPp95rlIQrTXje/Et5m+
pCqgWabsaeV1L6fu1X4eZ3E4wFV+8Thk3HXbicQeTTBJJHYcG79hrAcedesM8KNB
TtvzG7ZwK1KzMVDkhQrLFHj24VTmj6S5+Oikul1PMAKwc7IhgacEd9v1gy2zak61
+69iZLAQYrZ7eh1VlgJWt+Vg4JcCQkh/Kz7u4qhA3gGGDoAatCEp5RZgcAvzFy65
lewQcgmqKJ/T94wX9hGa5u1gaYhY1gQkhUdfGKfdzGYQ8AhPjl2uEdjqkjTfsFui
iP+9Hz/OKV1og/5bOo4xBQ9rx3EUFekkT1tNFyGXauyx3PI8i5ZhTz5Jr6/XVlvY
eOpKBDELXztk+/Uk9A7iQaMKhl4b4bbU1hDyblhKukqqHJMSHdvhGjAULKWzoPif
fNpafLY5zkBKaqpvnTRyC1hlrndrBkOKac5rnLlMN6d6YPq9VSyfGS+mJ8pqCQQW
cd1rTP60lMk2MhqzEVGu0CLmj6/uQ4Z+sZeO0atSzlnQuK5u6uw1z1+U6AEo7kP6
edyEOuecjy8ix5p/OPetAn4n1o3MEDAK1WPH2v6xiSjdE3lBT5c+qbLvc4v8KF9C
N78JwAHvtpBW9qYg40B/kaCovCIcEY2P+3r9JKDiRtR8bsardu4YiD4+DR8GqoiH
kfuxxti+8D9Gnm4C6ZB5aF2UeaL3gh/QusGHQIa4pFXWy9jXmtDY0FxEuP3Aqz8z
19X42xAEqE7e66hZ0gBj9eRBhwwtHIvSx2gveV5MqVQ1n3TCMewCrAxitJn+0Miq
2HuY+wHgpk8XwNPYvieVzGxKQNg9N2MN+yV8dyqnhiE9K+8fzqHeIj6b6OyPVBZE
jaoNWB9sNtcc/yF6zQbr7xiKqSS/Av7hgHQY2vBsxjrIbqnXaEo6OiszRHT8Wef1
8ED0TAUAFawQ5ohYyy8bpJjbm4unqOL37SDkrZjrYSomsSqfDXJ9I4Erko2M7laq
cPksy3EYKqTtUkACUTttp2OWBZb9xgx1vOikONJrpVOB3yA766cdHSZjCEwmzopP
EZis3MyOzs0okyd3uiMobbTEr17UNpYNZrMlXoEBHxQleW+6XsztXRTp3KVziQ1Y
bIFc99czYOyvORJnB35KK5PYueBDznRnMlyH3U8o6tW5sOq0O5o4XmzshMGjRJQf
iPHy8llVZrImYRZAgghDjRR+aHHvWLgbTLKjXifDOk0cbr0fBzkO0UOEXkwQwqp2
9ysKZJuZdGiOirfzz7pXYapMPTNaBK2bVT8FjzOBH8uTyaNgPXMza99fS19prk1e
sErbhhZE++mYgcS310F6zRYf+cBhduXUOXn+WflnLOGJ/QVU0zBaShbDlvjqtFfz
lm5dCmsHA/K4VVWvhZ1Q1JAPbWwxxPDf3M/zIx0cERmnlQuklYBjgP9RqUPyZ/55
1KbcQLlJdWc48HFjiqZywcsqz/LYMoBbNhRSNxxoWqzxLsUO93OSnZOz/lhG41VD
QkE01z45jLzp5tyawQFGVWZ8gXvl3S2XbYDji1Qqh4idcELxJfldaTdeIRmbcrSp
Dbgu9LtO5+oYCrOzGdpKaDblo2v8i5E4LMSIkEg03J0iPtqO5ey6ggeXRHhdjGX4
c1A8RJ4fbioA+h+MCf65j9kshXd6oqAg1NhLwvPhsbWazIJu/XBMgYKaiySeQ4mz
VF6Iekk9oCzDw/cyP+ydyckjjxhgD2hW5xVY3WgbhyAHOeLcvvqKAuHgm5lDfZmj
6naPg6NlAu9cBRYrqAX1IEfZDrexSBQu+4fzzQCxMgxEh8Q9/fGQqjYS076QQrau
KiavItdI4SSmZwk5n0w25Nq8HEE4lyJPVaLeuM29QQNZ0c7//8DjzkLIBG7hlfL6
9ftaNVtetWlE8OFGxEZx8Fk90Wwxwtb+Yv1mznwrwrPTsPmceHd0TZGddsZL45m2
Bt/IgsVIvxhysNm6mSYxEJ35fS682lWviqMGy+8z0yxc1eXsVMJIa0/c28Eq17b7
XTzlJ1sCzEY3XdFgmW4wl/l2Vxt5SqygYAvWN+VE6zXPaDzXSLkC2dMkKIdPDPxh
ZjRG7kxtUeTdvGdmP3rjwf7E9EpB6oC0wvzZeCqAOE1GAu8qqkqjg7Hoh+xfuZIC
vBx+AGNIhdmYOhBY9aWCRpwV3BymPiDBm7eooq0lBwREdHmX+oeDrnH77KJFEYXY
GiAPgI7diVGltsLNYe1p4TUASSZHJd9VU/Q5t1G+2JNxpQCy3fvFIJzj3QAemj6+
hb+CUTNk2z3NE4Zne41AylBW2THYrTE2I8onVEYI/knxgKmrDN0K57y8p2Z96gm6
k2xClj02+huca5pmexwgoPS8Lxawy+H6NYdLyxD0WDBxL+QNrhUOQK1lajOakFCi
SAC3DWbrIetlZXpsncPf96sUJWIrQqQRxlBeOAbnH4no65jU42UdNGq5YfZtTzE0
CoXRtQIaUAVFwvv5NGTVTKoydbd88U7jPRkwIiMCfaMxd46LP2igBAwPSydfLdX0
w1FeidwxzD2PxfnE/Y3dY0TCe13O4IPtu/VERa3X8LrZHEf/Rzxtxq3bi28Xyh+d
th97SBOdTs16icT878k1ErYNg9wOAl+vlKF12r7boc6sCbg3R99eUb/lTgvp6W3e
EMWDwnN1pYUD2qWWoExeVp4oufr36NMWBTjDg/XK2aIGZ9M1kVcYaKW8wKzptzbg
bLNAHAIlCz4WIIuH2lKEIHO+lfhsLV4RUKBme0LsH8w5oSI6uFisKaZExvYpQoxQ
8kkaLD+17uODwnHa3SyJp0Xi8n7kxgVrK9SKjYPAwnDkC8MVK1r685chXsWdjf9C
SsT0No8MxvIThsJt8nNjGOJ8eMBq+Hut5DAmtY9cqhVsIKs4tQIFTRqlPmS8jMzT
niLEZxxs9ioFh0OxPt5n5Z2EqmX882jMqzigZZ6h/gRLoYdlIWxbLW4Fj7fmMUVo
c3gogmdIX1mMLfyr98nx3aZCwZc/VCsbV5yYxNSHuCtXtl9ckIl704acA515xNQb
N4M4tmpQfyZ5lW3Cce8XHYu4x8X94qIP282oykdi7u5CF3R4JB8DnNggJLmKPPBT
OAwQI7i2RMrbgq52kZbrkEut3VXyH68EGC2Ei1gNMNIFyrQsFy3P7IgRI7CDXT7S
`protect END_PROTECTED
