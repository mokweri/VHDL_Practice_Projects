`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XV1yEyAJ0Z7hqOVvpTPk6Gge8AW7oJbl5J29chBK4C2dPU5xr2Cm+kOj9SXiJ7l
qFnU1DwE9N24stRU2eA/Ve2GRoCDfdRqDf1PpW8ddwZY5DgckeNPtlmfi0phzUbm
BBJaSu1isIcNYkOx+1853dDFKR/etYKEAqbSxaObZY5nhawuUnQ//OU2Nk3gZWTv
vvl5One79+sTCQ/LrLR7MwlmG6KlYOXH+6bLMuLzbh1fhfwizaNTtcUKdkj2zvma
+Qziuk03vgQ13I5xmgV+JD7OmuLwHlik3S9/MAsfhPRZAg6+hjTODn2tDzuenvlT
/O8lyKgl3wmin+QsxZB9ZDVR3FvGrASd2VxOqsN2v2j/oISHWt7/6qU6oi8uB9Ac
cJBabVkW6wv2/qc++RH6qw==
`protect END_PROTECTED
