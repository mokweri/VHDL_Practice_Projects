`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p5SXJybCjyvIVpsZsABJFSdaJpIP0NMNFkPVxr5NOHOKywUN1exsDrWpLZvV31dj
T7lFvt0AEXQOVl+36TEvgPIyDIKrJgVC2Mhs3N20QqUCzZbPOsVFkNXeoa+tFFiy
GYAFFcPZCVVpZDbrXXf44QUaeUHxwa5zc4mln06z/iVGpf0P6gJwa9vyKfyLGtYU
zTeHzVb4LDK960Ueouh+aZiehIDB4PZD+ROepX2ii4AnOIUnx1/5eR0HqWJhqac5
nMUoz2JUjrnkCM/yZ2oj3Me1Z4pGqhwOFYdffZCBjb+MctTHsEhIHqguQftAFCQL
VJh0O2LjW6KXGEww6nCIemBzUl/xGrgpw9zXOSpX03tnlfnCcRThPFDpDh8VxCN1
xKcYmrpzEVMDCmLIX6QF1X8q1Nf40EW7VOxI764DnmXDpYoxLiOrP6YIk+TsQRBD
fRT/owvwhKsPJdzhMg2y5VXYF1n+p3TmNGLsf3WBuxP01TGEYWUAYNCgKHxVtt7T
YownFKHBAFswSNj5s1/nVE9jMMV+D7DpjqZ4k4jBsMq1jhJlxJkEB6APdmGZwnNU
NqLAQKiSYyklG6X8YxvjzSYPsa/kRpEqMo7mkjD48whPcM1uDRauaa0KGg1f9sPl
+lj6PQNIFEnt9nO+oqCsNqroo8TPPOyqYHarDCWJ/ipwIcdDdFjSTxWP3MQh87bz
3BHE7fgoIdZcugwESZ7J4mHzYs2PMJkEtlsT/f6Y4LFDgaKBSZ0piC3GFZOxcl8q
LC+fpZ0UFZyoPy5ks1UBi8amu7bQuS1luKwZ2ClIw87OfoUFnfEUxxsm+y8Qw70/
69jTuSnXSL8OJ0+m94eDYn3WEpqMJ5DIrdOcPF72R3A3GZrXo0YAUb6Vt/wIEjpC
KVwT4PFnlxSvuCwPjacj56hULZZ+Mkq33hE6Ne6x6by5EqrwGt8m5f7MA9Rd4ioc
+yj91ev6pHAuShfUrh2EldEhxGh8b4s2Zu1ks2zY2pa+joSx7+i0qyfqK93KkwG0
HqWLaLwhvDpvQZ7fAnLDb5zVJzyDJ23s6kHp850Wgx9GTkDX/HxbfUUb4kYsjZLs
Jo90DXmsICaf5BSc0x6iYpZ8hLmA3pRr4bwhzzwom0LG3eqH7tv/JvGfRQX3eNq3
lNiLPx3Ei2PL5p44En2aR6C4hAHsclQe5oFAlnLEnmVmQZW5mF8Fjm2XNgbtJfbK
oyjrjBQR2CVPrsjghLSEbk81TT1jIylV2osVkhA2hu7nWB7tcZVcVcCcyVErJ8D5
B3dWb/fQy4ooJQlNHQvYMdAkucKel2p+Wi9AD0Ma5XneTpq6HOSWsQH48wFpbsF7
px2VKTqHLO+/aW5ghd6ho6nSL8bawD2Ns8PAf755V6tBZpvIcj2SvSOsxxG//ak4
Mc5QEPnR/GlkX/kxj0mYrDqm+57BlqZ+tqeZ4dZsk8+E9BM/ohfrHgfIxbpP4A9A
Yb3JrDY4/fiHBY4QpBp9iy5aAck3kmQb0tr+NpaQ8yMF/bw7QxGL5qm2jPLVA0/w
x0zerVqMfizmjFxEzwg+eIFSf+Uvtme2PVya4PElWIxyPjgrwUejgg6ZBDtEM6MZ
jHutK+zRI1twfyQHkqQMwVC18fXS4FM7sW+23qu5H1wu49BMWi4EpE0S8Jcehnoe
4+i1QTWgpD/SCrVDzenBo14VkdGVQv9hsPFR2aRElmzWtflPCRk5kmYXOFtZc4UA
5JEDipHHfj1tKdRux2275aqUbkefqIzgBQ591TI9yDRjrIDW98BqI1uNV8Wu/Lu8
I3qyG7PkRNGb8uZLo4lvRLzhLliKJK/bfljMGJhVufc9tcnm7D2aR3LBryz0yUKJ
I9482DJj6rC7X4kw8TJ22poJ5BbAj9AnF8r+SZlPxAmlhEZ78GX8WpXobNuIC0xO
6z3UsjZJUk3rqxVpqeW8kzNM+QruA8J6hlxx7w5ISpzZ3NzoFH/iVt2OGvNZDoQC
xP/r/FjeVhqSliKD3vVIBME76KFd5RYvPEAdl7NfEkUEJIo5wB4HBMD61MvGIUA9
chYnAQNNhVRxL8ojSyMpznOWFR/iJnkM0yMRfRmsg4bBwJuhEf0sRJ/DnBMXdLdn
FDXQ/UG9MqKRu1PPiG8cbxU36RpHYkhaWd1+pSDyOcQ9s1xGOxykuOC736VAwOAR
1vedS/WSrdXTWH9yjqE22D+pdNkjF9INEqqplXH/f8Ffsb90N71n3654+MZXx7GD
ckpQPxV5nTgKiq64PNqmEj/dLNeBIVaNFSIYqemTxwweyTuxwNMD2lt0Wjnkk33p
7t4RRRP5K08cbZIQPsIbFQIcvpbHI1dRNhhmVY3pM+V638Jy6IbFtpKJgQAjwp+a
uKSFWiyX65NEIslXIOoiyWQ6jzFstcfn0nUqZm1VltEKW0wUvuVIljaDvszoaSwa
7lFavska3s2xJ73Abtf3ODz4Q8vqW2AM6VGO8dAdkBVuySbjBuX+jeTIpAsn/wKc
J5D2Ltmx66aP1AGZpGMkhOZhTl4282R9eWx0x4tlQwVgRK/SQJh/tJX88OlcWCHW
2oD+fUGsspmwidZP0sK2h8slCcu6P6Aj9PYHlNB4OzqZkdyWPSly8hoOHnGAI4Tk
l1rWdnZoe6mOeDLtSsM/ImVKzgmoygYybiinLhbUsXWWoQrcuGaWbxv3VjuC62kw
r+447G6gC5rGRc2tu10Neuqyv8nxPsy0b5N+MI+RoteBM3oVMUZ7wEyP724Svrdj
giGONJc8N61KpZBWCjfnNcSkLtpXe9mI7/3l5KZd6Xn1yqeDFcln4OIcK2Tq0VT2
CmLTsXNy+GSd9zdc8z2apGo3zlIlK/8NF6lSZD8pQJu9pP10qM3BE6PQ149WkKSD
mVsYAtnmPKcWrNTCUA3vEE1Zp++6Xyl46Saj4ZAwn/IavQxfvt2oL3MU5XmhOl6i
MSPAdEDOrhZYmmU+hb0BxwQGKAPKIZ1cPdC8VNtjgoY5g9ii3pIJfsYWVVKi0nP0
8Fzwg6aIILGFSFZUNH1J+ktbbb3sUX+4AEyESi6wyIJmgf+GmRhdF8sigT+fUXvC
FlZPRSBH/aX81a0ihjDzJwtEH1UQTwYF3hI1dkyb77oPIKFH+pTgI2tyABTUe5y7
6QdB1eYpAe5M+bGgm1deQdf7QTqmU5EbEZqWvtCzEg0QJZ6HLZTousoaOSITxWvv
RNlR5jxVrDOCGhNJTWLlgU/+p4hyAuKPIVV33JoDpcHfwExR/rKmuA5HtYohr/ft
qdNpDWnZO2pGiWE7zHLY9+4DQZZPwwYBMhEogTYWfnWb4+XwoQSGAZ21mZ2vWBrV
TfonRSQteHVd25oKIDEgrwBVLJPJw1QfPk+wuUY9SdTv173ZjKVvInoHdozxnWTX
QWatmN96UW28cZ+wKCCUpcSlXbhhMqoFjgwpgCRkoRlIIhBys+8EJu8OE/HG95bX
i1kfMxLHzsCkuSldJTSCK4fVhfuWcR6KRZVXaMXG8rqcQV+ZwL03XkLKRVuQrDRa
a2gyH8+6PBaUNzlV8cbPANUz5ltZ5S5q8r3rTx0up6IgP0aEAyOU99cf15J2gYeL
Vxa/42fNZdtHYVx44wwuPRqHf9IMenUmWyUTeFhxSMckxnSST8UCTtc2lzm5uZKy
t2izlvLtLgjO9FgwyeGGRn7NGz7H5T7jFPoLts4txaEwhnHI7qg+99MOOysXS4wb
IVyozE4iDHEBkOgHVAizMLcDv08D0DaNaz+e9mJFV1s2ZAriY9FqCS46gDFYdjny
SICHnKkKe43JVpkm61Kw+hnkr10GyoVX//MPAN9WLgLynqWfOi8x5RDGbGQ8rKXa
NLT0VEYFGXj3JHLgNbBKvB6UIQDvfumNkNY52rW00XNfFOf3lHVbYdHuUDhDkRwC
xmTrHSdLpgrAFxcJl6o8ZB0nuegJ/k25tH8IqNgqy/mHgQZw8BJJVus3qe6FIRL1
QQDuneupr+aLat7Pc/kUNtKDGCD9025TKSGBPzR/BpldDYgw+bR0U2Zl+THmcmJn
0dDw6lOWhkP/IcG1i6P2ka1C5Bqg8u7uLiIIHPXnbUKMbmdxY4DoOwUkVjE2t9gb
0i9dZFg/QELw+mUMLW18GuK1MrBnVBrnavBdrk+wD4/8T9JTBkRwDo4cIMwgCOzp
/4r+1e9dVdKulnirTy6C6L70HEo0F8Cnq9rqoxJMUiR/VIxdTn0/+d2EPsLQdfSr
L4wUYRrRx9blKW1k85u/q0raIA9vHf5xQJ8esYu0fwS/MK+qiRlC3B07M27LtNuZ
yrUl6WqzFHV4iTZqgT35FR37JUBJ5y9j/bkF5CDWS+lWLuNdOJKWEVEBYK9yBx2v
6R3T9oXgc7Vg4a1Ll59etdnwOBHE2d9kQJbfCkzLhZbpIqRLVNXp3U+r4f/mAxZW
nP2djgHjZQnbMPvSOQfBefBu9ivTCF03vuAUWdpwgacoJLi739xp2ZaZ1MvouX5C
ad/oqJdAvJr9fq3b1gdAS8WGpolSOgMnk9Ho7IKpkuWIcYZ87hKQ3bAWkOksmLd7
n0GJD0QGmGO/GbzfdbSeMVVctybkPTPCfBBL9CZIeIqz+1012ziUOSEFxSvIZWbD
I13aOHvUjDqdygXILpYnrQ==
`protect END_PROTECTED
