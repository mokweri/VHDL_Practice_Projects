`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CuoWyC4RzD+ZlKXgZcr1NhoKcwYYl8OwdtLmORu8IMqzgdZ6uJlkARwYU4X4+7Qr
xtDBJqrhfytZs2+Uv8N0s8CeyjjawG6bjIZa8hRiYfXc6iQH0qUx0CwaIx5df7u4
EWb7hG+8CL51QAovXuBXvHvODqsnnl0e9tTsmnDpmK/WFxYxrD1o3dM/NS2eabSz
MwYbylPFrnFlGxP9C1CfVPuBRNiQICQcxum6RqK7jkjMUAxurKyM2s4uFEfrCR69
+NLKLV7Rum4oFbhdzOKeqkeuHAEhsqonoLzzaMrorp4uhn9y8FeSwuK96ELvEnEy
b4ttPUEK+ENGdETBhhgNj2rxq1SnIdD61k0XtavtMYx4UuhXtYLOspD2wn/lEYgN
cV1ym5cAeW7FHThvyK4hg4AGH+AWkx/XyTeXfWUWZxbroVekAcrUp93TLLqHztlP
jjHF4aVa0CYb1d0x9R8WH4RqrfZ7ETQMKaexQV+WIJOUhWDoN5ZwGWQnz3k1qhI8
I7ct27oTtJm52V2TaogMO2uDWe00ZTdiZg0Co0USbLPhpxEObkK602gx582t88iL
uIjw2mzti83NppYc7LhS9aMwpKHEwBtHQmfh01XF4uAACOtuOMp26TJAf2g/PNEY
/+1o1VdcZfEmIa9ekP74nE/1DtgmAL/rTjGIbyuc5FRaTX+J5nEaky7b80oRU79m
uH5+1Cstrc6icoWx+Te1uRgILavAe3NIoYRAXIzO/XQv+/d+Vf3yleQXGn2kfRPX
YbzHMBJ0valT9FJ2rm+hLphKksSx1ejIVQaOxysQR3/UQNsM8iMD41GgLAerVr0R
wakIpG/0AxaQuRbQN+aAiNxFjcoX+n3eMxK5zv1EtP6ZNkMd6QIUugwHgqTcqm1k
oioOQFJpgXnjvFgLhuBG1a2HzDp6D0VyYDRXN0ongpdZmgjHBAECXWZe8qtVMB5M
U4tn4f7iKpR3uPQrMlnpzSGOmL4dPiZhHY48PfCNdyuDkkV1C1geexQ6/fmUjWMP
3i5aaSAEK8MCF5zRYwQRHDvXhC4DWA16w27LrP8Evm1bBhuci+qtPsMtUHpIKIuP
zzYKiNDz/+/Gz8kzbkMwfssL+QV4gBA0ezJnz973NIBgEwmVu5jW5/dK4rb4dbIo
OmIFoiC19bbELBq4YKPH0K8l8JGTCiBK4zN8PLYso5XF8cVsiyZhdK4owhTceT3r
yltkNey+Kjk7cW6QCxNSCwbsYxd6dGL2uR45ru/1xb9NjslFx5x90UDQw3i9xzDM
DiflpupP4Nw2yPqo6VtD9wg4v92mpJ9G7Fby2T0RQMK48iDbwEwBO+dMsMZpYbCl
HjJaqA2rMJNANuicbOCOTgYfYdL5ddIl47ETEGH1MO8FVDpbpPfjCuYa3Jr30Hmk
+hzfg+Lv5ZJpx1NCcVOztb+Z7Qy598CWNSoc6jicEue3f6eeS/ykYpOs64zjI5za
84Lge8Z+ZSa2VY+aXFkteDvMkqwXJiJ5nNyjwjWyXMUS0/C6hF1sNlFheNA5gHDi
/44bBF8YMBfT2QfTfknjZr6c9ugsaBMdaM4I0w/9TCQE125xbP3lLkZcdf2vy58I
pLdf/R1eK1pzJ6h8RRR2wOfmQh0rfXyXV4fbHV/zIXZeC05eHoBgTO5I9XllJKOH
6fO5mSySzPK4eZzumNN6fNsFO7zqfrgG051lVkiYJOg30CFkTy5CyXCvYIG0y5EP
G4naaRZ+Acxr9wp5FSqsyH79T66iQqqUEY38OUExoEEF80zsDxaIkG7cBmS0GIje
ea9v3EWni+5rAJ1L6hBWpLiurzTJ4HUAQgTkDnj/Ken2BCdywXrn1B/7ojUZlmRC
/dBFJ/F7enDhgkA7Uu39WIgNpPVXUQgdn7u/kxpYxFg+/zZb2axpzOzmIENh3HpI
QNa8vtkPAZxC8B5+cG3mLZDBcxzgmlMJkrrm/O7JR/TDv6dNTpfG8TaN6YY8il+/
zEE8Th1OF8e9c/N5+jeXT5QWEpsOQXhQhNPOm6ZLatMPw5jNumHuTcJtdF9XxgIX
Ky1d36mgP8OUFsRtpgIhtzufwE5fW+jBehYPtNzqzAW/Nj+kdBmPspo9UcyRhfYs
4nAnyagt8gzOAobtjWuXlzsLXnj6ysnB//4a3q4fWaF4pRGvQn/c5Q6HJ8EXuzcP
gNrRZqRQsTTUhWEk3sB36dtHbLe7PaZR9klcabrzMNBkRbW2oRpgdYh1cyLv06oP
klT37k4F0zZ8zjOynIOst7ftJrjlzv/L1uj4TBgUpzoPjYN+m/7velhL97uicevf
OWwXgsT1pQD9UtFp14/3rs6whPbr8zG6F/aFy0pa9bSIDD5Zz1329GgRet1JwuAM
xBdPsVbIclebPVDp08r6iflLRXeZ+a6sPaPGQXCrZdE1NMUDxLtTJuEqw/a2xRct
OkElLkoLxCPyf3LcbvtauQhXqvExGePiGhheANwWxmgY7PqxDdG3P0kpVPtrHPRN
Mf40PUFde+qEw1YdSTxiVN6v9MC2fdYc+ojSqeF3+RZaRLHQSdjNmBL4bjOvVETo
tnkKVzPnJx3r0AhaWizi0m9lT+B3DKu51qSOmktWK2FbNorgRMe51jW+q6gsVslR
Ek4hsnTGCPIxDixv5LwfaBggoOjVxGazC0P5eqkPhiw0+iZWpuumPXQ37jylGHYM
r+edUFT1PPNXXKyVAOFOo81Bt6VYIc9kMzY4pPmnYFuwdmAzSoS6gl96WXy/hVT5
ZxOziVRErqypz8B061KYcyWeemLk8Euw/KiyCDoSrJ/+jwsE/NNLPkMJEOC2pmT9
ubvjJ6yR2bSNgoI+H8l5eQq7WupIU7JjPgpQobq/QDRVFC2827FRVuFglZA9YUcs
nrFDFJofoR5DlaDJlu+Lo03UPu1EwUyNHDVBOLJLwQv9TlaTlkWC/O2tBmPf+Gju
01dK2QUD9po3t/6OqWWMHslhkjoVRgoWhgQ8j2gsJ9fV5pItw6pkhuDFsR8TR9LR
WoFTwqhKG9jWJgAv65g3M6tGzlXeC75lp7z2EppVY27DkA/9Vs+ImLBdVlNmoCm9
rl6Kpidpx+FyjJgZpYVyKAZv/cHkwErmVq/6m0hGBCHTMeP+UN/u3Ut8xs3EqDsQ
8kDPwljLHuToWAzIN7Mvz+XOkOHZAaERlRKnyt89efOx6HkdQK04pxoCZWMhyYDQ
pRVs5U1G9K8TITFC7c6wn9ttxY6UJfDiflTE9w1rQPEiIK34bbL+qDhvUT2GNEGT
Y4jQCPmztYj1+gOL8u5jqwTqEIxBEQfbtRRctcuAa9mzjD+T3LHQUHREHsVJJzIl
avy60hYOofQJf2z6XY3h44dcfrhUrk3uo/Vij/kFhmhh3sv65ebQU6zgnIVf8egL
HaVwJvQLpK3YyuG9Ajw0Y3jveviwvTuv73qX0plpMOPWBfwLqouUFKpn+CkRaG06
61DK4hfIzXn393ZuMMir8FFHK6oksJ0MhYO2xvIWlzyYuVxiM+UZJrFPSeSyI+/D
CjlU9xOneydhajQxTH5Hz4uBlq6vsEhKHiOuKNRVmWePiyi7jf/x9xbtxMZJeE3C
Y8A4+tBenvtvuDkwIB4zYDq9ClIBMrCIEma9c7IkFyXXA3kn6jQwGXSC+nrEg7OM
XyqG3wirAD+7eb3kh7uOBRwm+UEo0GZIMTK+fhxH7BuoyINnJkAtMNE8XYOzBT0f
zrROVZjMdYvrPH3Tk1j1cAYaeCCHLBQFh0DtN2aDi0mHOwWMYiGAsRC+/O/9hYBq
tqtrARJBV48vIW7dTkeNtzc76wOgVOttxEcksaS5tZrH4a6L74j+GaZrceImYmyi
k4pgKzRtoGr/PKfjACwqL0iiztCfN+gpVSfXzIW73XHeYFxbieZhXTbApcktl+qI
2GIqeacm2j4GGZzZ64i6A5veHpI+s9YUbMyF2fY4T/+uX/2ZJXocAqMt+1LiZf6i
7wK4RhRWEx0yICUQFTF8TExOOOhQ+BmRBmB7cYfh687j9gocFQ24HnC33eMK0n/W
P2WsaF61KyodHBSOz+l4qBxSeu/byJTILzntNvNgdOyMHHZLy89L6Gtc56NHQ8+e
pOU0dmF9GwJnjvSQqH7CNmmTOHPDbQ8ls3R3YK5JkdaFgVhd9uVDcnQctD0G7I7n
9+J+pSvdtINqP7OhbtwPu1iGyizyFRsXVCpYm7adbOUyVetM7YTV/DyjH+olvxyU
5UBNpx3OVVuRwz85LadsMzl/Njztd+GS1NDOf/sTlEGxvlYi555FQfzcHnWzPQhb
`protect END_PROTECTED
