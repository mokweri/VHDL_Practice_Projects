`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pki4XJ4cVIaCr9lbeyHrAuFEaveGNG6aKXMl3Pj6zo0TisTQbUAq3lDsLkAFQJYx
fQpSlNB3x7ZHjFgxsXaWZ5uVI51yuH3iAZfBVIVGY7Sp8FQSo123vW3cwnmgoQtO
gH1sZ++utn40th954D3/iyzH2psskW6me3IVIDp6ILTUBaThbE6rW9Fiv1ngAc3k
Q4quxWZ+E1t/gxlR7QQHr6DX8EQlXYSHEq0zlnsZqYctPq2dEMdycHgb5iTte2jW
dH0V2pcz7tM+xZIPuJ09o5wDoRrqfOseV1PVWhWbnnEh6l57Ct20zA0cjwgseKvl
SrpZYIatXtr4mUHgnQn6Qt+9TRw7/ZDXTBZCSrfB7bzR7H9iwNPYemnEKbpgEvzc
Ysp6O8wxMr0Err54q3TqypBMLqWwDp+c8V5HFpgYAR+a49a/zhpI2iwSeZ/gq/oa
RwZgrqqUoElzSOSpBizXBrNQH7EhBI6wRla/iUM/OhGW4uD0l6BaVoORz0g/hByo
j+A6s75a82FvhV5omRgXdZYHOaGkDrq28Ad7tV9FMRl6470SUsWoLHnWC9pIbKLT
lNYdT8Fuk1ZNyAcEEjnbTdFr0hZKGCNWvkB41bevDAM=
`protect END_PROTECTED
