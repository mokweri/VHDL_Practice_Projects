`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRPNwCzhFxu6Ov4Qx4/r79pNGAbLwl3ng82Cb0EaqECA5avJM8OrwWPVbEUOY65K
R/lMh217cTrWQbC5k9Rcklnfispj0Is3bqpRe8R2DAcHt48H4QnFLvTLcDC33Q1f
Z1wlGA/T8N+LfNJq8/8xQ1pxui05I33Mi2r0tZIc8a77bdBAXHSikKuXCoZiSCj0
CThqb1REtU8zZVyOMSeXWZU+IV7PgepcY+9lH6gfOc+EJcZgvXQeEGqJq8BuNkWH
cy87jZvc6MLJM5imGizhDb7MeCvbOhRtBpjmwN7alN5W1EwsAcKIEJo9x26Ignyx
Dd236f5xuKLPdwd6b/m10H61Q6/JPoF/9KAw7IM4/uYaomHWkwHwcVJH0CR07Ibx
6QHY5n8l6XH8P2ie+5PxVnOw5a4k4pXEwp1BB6s+LvOLD3Db3QDtdHRdGm4M2Tk+
DCwoSSwsHoRq2pU23H2Ep7RTV7R762Vg3AxDcS+Q8E7S2ZpSAtpVJKHv4WYZnVWq
+2RE6MXYUjjfaC2QVGid/o5cPrChPWF+g6RrM0mMsgeka0oClT76VVn7ResRX6sr
Uo8/gj1ssWe+qGYY9YlDHF59NBIvofQ7WVyPvEy3kYG11+DjKng5vsUWMFQ85nKM
qcysL7NO8W1oeCHNTr2digLTO3Fpl7RMzOak8GUs6wL9EY7zni+H4uzn5MgEyy4d
7rw4lfcQB2WvZllsrjbglrLFCrWrY+jBMWfw0p28nU8KJ+5Viw6zZlCsXu0nAOS0
wKYg8fOtEQLT84WTwxjmdVvXtgUjGOszJ2WaoeH5E/pwZDfGkpmnQzptJkptGkas
jAXOv15HpzkdfSaeXxSw3OfnC2ImJFhfMqrOKV6gHYGna7EcsKDon7Ggrb8tUbqy
ObAriBCMFfpvX5sf5YBY6SwoT3nB7tltpedS0E9Gv5jtdeLOO66YnOAjPcgyPaYT
tptqodamS37dYAPBIyPNjN6czl7Hb35flm4JVs+v/swV02vJs9RPIe1McAYTf3VB
jLrv6uWc8ICXMNkZ+0+R1XfLYUiIjub1MiEVRvXdxlv6898em+EiLTi53tpiyLzG
p/dJZQ3e8HmKy3mxHo5q35xIvYsib3nq67CrrJHbS91lQkkgzg+5KqLSl3AtMW5E
mUS7tt3k3q76PzUxaAdAjFKkM73YsUus3TrfpNMNIJnh3LII5ICQKXzOk9RNyJK1
9asv3+Gb+vZcWgPbkr6bX5j0nKRoFVzwqlOnsg+2xuY3l+mA6CHOY6uodRJYur67
Rzvz3I5us8z3CJHASYeS0DsvN2UCg3wR86HbTLW5s4raStLTwnRXB3W/zXbMZY3J
fCrBgSH7FDpvFoqBlqZg+sjPL7if4AmW7moPZi2KYFuwWOmSX7PnIcZzwruXlXnF
DXxf9e9qfi1zYrv9wzZCUaCZoKGMudmiJI1xaFyOkzB3ats0QWK4YVM6hzTvsYaL
EWzpXCbl2bepLfuvKLiP0D6Q320oJFE9Wxbw9hPc1jd+SJXc8ZKiGyGgpOmrBn/s
o5PSKUKHqh7KP80SHp3w2Ai7SWzChpS37X+6fcLukz7Yp4v7zl6ZCSU2GCXCpaR9
CYgkBkWluIAwDhl7usO6yrDgSqLUdvSs8/ZK4Vh4JeH4R5skudjSroMrxbxeB5c2
Ho+IOUuYrstpJV7Eu0NB05elpYwMFArMxpv2M/iMxx1y1Dcjw2q4FSgaEKgdmddu
sc50frn6FCLLUsjH3WObsztkUHkx3KKrFHV6K3uOdcDVj6oXCsIGUNKNXVRFZt8Y
OSxTF7yJoyM59w2gZRX0N9A4LmNS293jXUVNeD1FOXYngYsVCpigSAH0FM7RtrPM
fsVBGlTRlrwpGTBjD+ozp2vYMihl8rcael/oZ7krXIVjUhK3/4Je/BdJ+ahx1L0R
guYFqkjPiLS1A2mNjwia8jSE31LDdiL7wODFsiivzfQ++sRQo3JqWRbKDNq4QaAm
1nzANspJgsSpAid9QNabu2k1kMEcP1KC/WXNp2Fv+fkfEq3+wv5X/blmJrDYRmWb
Y6l8pbrOAC51pw7iH8znnQ==
`protect END_PROTECTED
