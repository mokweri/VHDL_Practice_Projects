`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CB1l3pS07z1K3zIUtpXoG3bVtuodiOTG6hpWQnsLcC2H3LfhU07JaukviYagO3EH
nacUaD8l0uWaca/Puti7Vl+xg9WI6c/U7rMivL/QHnkazufWkjNDRNWTLsYB7toT
6F08rCp1LNu8t27fL97/n/jf73SsnMZXVIahAzWQVRo6Pw2hX1CwGtdtffuxkl1u
nW1NtQAqwkhkSMnSKhdyHHKzE2yW7UaJhDz24pKp7OfmMTWK1efOoib5QY5LkaqG
qvyW3FGF9Wd90SdnIPJIDpl5gabSdzAoc1tSTHiRHiQjVQsdQ8gsVH0D2K//3bTA
89ORgkyAg4FCxQlE3ensEZ4tIpEkzWvEQ6hoWKCdbIXobbSUeAKmNlnjggsoXMeh
eG17Ko+LnXWOtH3BjjT3IMFZH7n8FTibX28MOzZpSDxInEFqxtLULaBYr5d9LtmS
ehcAfL/wjmYskcQURtC6WddVFZywjkZAbGOgdGr36zmOVobujJI+f+Fvkc1ReQMG
RRBaqqEY1T08a1+rFVVQQ+0hGy27eEIW8yro9H8baoD4AjvoUgDhR8c6Yct6KG9s
nFF5ZLntb1+s2Thw1hqH+wVPcMcdUuMFhN4q1DqEOJFj49FtxKW+WxcqUjfOLx5k
QKE/IMGWXx7urZRHqZ1mkTiDIrbMFni2WCteBUUs15EN43E7+L4qt2QXO37JKpjE
Tzmw+XYO24tXtsqRDEKTvQqLB3h5OX65WCXcfyBN9Zzb3HqjCdfU5u6LLAMqYMTJ
ezPAEQbiyFuYBFSyclm/zGBebp+e9asWFyj1tKhkQ/Dsk9mMrcN0QO1WXK27Dwd1
qMN/35Bci+oCjkO5KKAW5MIdsHPDFdfYjWKSPbMxloVTnXq1E4bIT8sD92DGIY6x
CzT65FEQzMqwWpSgfW1Uxgvz7xD6bKun3AphP/eLVcsYi0ec8PCvXft1z1LKpTEf
3HW7YJS4Quhvse9AEg1Qiloyz7D8BBeFMKDByKlvicNqBQpYdZGajOwdHGuE29zO
xhSI5Sj0yTwhotwoVVXK+ZxA9B+K3D4VUe4lyNWtjO3RNeBNgzMw6IhgqRdM8PfN
Jtog+pW2nM92TbfNSqeXKTaVTXOhn5edIcEciA5yqe4cce0DNCdXY2kPJrsHFTEW
hF5WXwVDeR1MUmnI8DssFuU4YkwJgOCmdOEdMvD96IF4MN2m67dpxtUqb3bwiMVC
Fgs1VrSwndBGqakqfRVCcQWBD3cO/WrwevjXhySDhI5K89eKdNyTjQ0Y6QsqD41P
yCDbBwgSAfLs7Z77g7Ly4TOtUYMED3qyxzWUz69uRkIC4D/aJnf1wHzO5RgBjYoL
qTCMnD1fLn8zeNs3YzeQbdCb9pg88HX0qAJWHfABgLCq9e7H5djchOXIukjC4tCa
mK/ie/2H+T7/H2dhQ58byBnsn4Dyg/57WvrKe/1LMEIQJShiOa2kgJoYe901YmqG
QVx37OuoU/mEq1ztJrPvI0bTar4/vQcu+vxA8c/qJYzL8jkN+DThcUeAANTHl2+i
Z2Dn9MmewGsjnGwWFcNyQR0bYFSeZCEt283cDymGLku4D4eiNdS+7+oL7cwKeWx/
c1L0mGUzIqmjT3nDKfW55enKOuLE3Jke0PDGYk3hHNtXEDzilBlXS64eFNlmoUD4
lo0rIkslstn959qiaWAE4GHQjKOCnvR6P/nU/ZKTQyXKNs8tsnzGc0eKH23k3hjg
SHUh2E2gCFlBc04tHrH8LNUurldceBjH2Jnzdxv03rLgmwQipxXBfrINkjQc8UlY
vLoJ+6evSw9O7+0drpa3+maO1OZyVxD80jaCaktYnGLL0PDK+7eG9lvdkikesegP
U0w9ZvGpqwt5dcV0I93/n/3MW/oSkyObybYonvzvmZ2KyQ1JDmcq/b9rB0xAolb8
Suah9C5x/x8GPEdRzjs8c41NpQWYqYLE5FssGh5ZU9XtlperLr1bt6uT0HAbIegi
2dcK/xI86hNlEYhlE4tttcvesVH9uUocbcAO6PiPSZ4/zw0lo7Cj8TL0zyecQXFe
5LveL/wnQnklG2ZhHap1d1kY/kWPKv8qJgtzAz0nCWjvs9Zlw/6Ig8BsrY6mg0Ei
pvmxR//iVVr3m0QLYGP1DJh412ecarVDiZgneurQ2Pm4tB2VcJ2WbLeBjYTJMdod
GhR2GVkHXRXYCCmWjQBRmz93emZ1lE3F1wRtfBLa3sp6dR4pnc5IOvAj6hgRoBQ7
qcOFidPjZp4+yEQbg0kL8TaAjSO/VNC+jAMwGt8edxszHnu7DYT26ed7c7F2IW02
3+udhEO5Zc6la3hysZaSkBnnEYebVVh/nvNenn3GPJ+CVNH/dxTBG98DrX1WJ3+E
3Nalu4mATbGMrWfd/Jd0xv6fqNidJrx9tjURxoBqcu63hUYWWlK7MkxckcAMhSzz
ZRiZgUDCO2TDCWidXLKcR2Nr1GivwCK5JfpNOfqbxGYSras66foHDQqWbqdtbHgT
AS0SGZ6BKai5Xx6FrFbUKPPuviLQ61rHUbt2JFXwxaYkN7yfGA3oZuUK/4G4EqtG
jgBhs3SX2+IMxVff+11+p91BcO5dwhIs9B+QrYCo1NSb8fTBPBFTU48dHQzsgHGM
9caOFsaSYfSuZMUR2nFIEI14UQ3VwZovJrPBXFoHSabrHoDiC09rQI0qc2Af9PBf
X0DCxdYvhxJpKkOSh4KrGQ==
`protect END_PROTECTED
