`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2gOSHcdMO/lam1sj+rZ+Y72Qxu6oDw4dfXfIWTlmyHCNkx9mJ300uzNZPRVxsmw
kQWQ8cC8JJ9HCc0nghJI6nZqEWWT9zyMQJ/2Wm8UzzzGQAq9Oc2FgzvkSkunztTb
5oNod7gPBamD3J+NBYmK289qPoqYisA76zc+lk1K0mkRE+QfxWwUSyGx4W8YXIxj
mzUWC0kATgs7x5vnwnKpuawdan4OwqEdqCm+GUbXN3x607idOKreCToCvriAqHvz
+M2odt7feRGT21xVU8MNf7E657BpOFeq9o6sD+gcYcWYiPnAvrZOpyxIbqEfEW3u
h2vXIYSnTnw1mmVBb1OJHjla/NsNVLDAde3HvwvQQ0wrrsENVT29/nSyr3pLuId7
mEIDxa5L1e3LVKeNdDRTRUGGUD8OhBj47xodiYD3icHXkqZx+YTohAJtgix3p9W7
3IvYnV2LOqbudCAHLf0nDn/16WVzR0lcvHZEieQMRN8lVA6fLaxJrqsKZeFrNH9A
m/lvliPjnVm8NFSQHTZtX3QwnP4Z1jaQHX/qr/dSk6iukwe4XxNlWzXcKdWlkNSr
sRyD9pwiNuGRMxrmVBU+5pYHfd4O2TUpljpP76Ozj2BIrO6cx5oG9xK5MICQw/gC
hKpoyfgBgK35W7OVMkSu4pwtt2FeLyuPlgRZNM1qJCmYcf7sHWFtBslAfNIc4/gJ
vgq3xV34aueBUvQy+WLc3o1QTz0s5V7j/4jEB9EvacYghQJRxrKgSmt14ohaU1IZ
Yj5DOSyuQtqbNQO4AbETRXPWfJIa6YDBLEOcCvAaXUZsEWv0jqBrYcT7n58u8jYZ
AMoMB5iTowfgKQKkuY/0YfPQS+30pxF/o8Y+1nQfP3cwsrzkuv+d8t03hgYtVk/c
1qj1J/7xPCPTIii0FdqTdoUif8dGZX8Xtm09VmeKaT1v1jKVe/YfmClPSrLK/c1v
rTG7+kly+PC90H7SmbisgE53Op1V3Q0OFLrAaAZ0IbEs3CVhYC++d6IDdLPTdWXn
gXdTktfrtTkCxQYU80p3S1ApUu5fqTrNNtiRmPIaPr6zO49jUX4Oin5GzDdyueh2
eh2n/tJOsOu/i7hbQukrTc2cFjkK8x9POx5VAb/k6/MiIDE9EuBeFQhsOQzmtJKM
MjqRtyJ7yQMfAnSH8UEvttuiraMhU+FLX/7gA+8jBGJgTzRYJ3qc4xqA85CJYrLI
X2ilKlzQ8tfq+5xKo/hINO/TyETNibTrtfVkQ814YHVSNdl7q5yNxUI9Wahprsm6
Jy/8IM/tX4pSfFQ9OWKTnERRpmcvds3A17NkZBXAjpLaT7pw3TPnMVSewWWq1efb
U5q7YRtNpyWTvoj9D0Dp88fP3TNnue0hBDt44hsmgjVMUZUIuCKKTyIXNKDtQtJv
WaR4yFXRVr/mdvqFBJlnc/RoVs9ZC5HIQCflungCrpm7z8uadBuhQ36o0eZXFzCp
Ae6/da1FFy2MHQjI+0X0vJWwWTkDEoBGybzvOrlAy85JyzAeZL5HNPtU9DXj9o3O
zNaanQyjzO27qxvPiP7nn+WfnkJtU6pAosNIbkED+mITh1HOPd8zAFA84bbYju1J
54UAetGX4G3CTskbpaF7+WlFYyR4JMgnIeRwhxjf/T+RptIgXDmg3p2pYmdE/k2W
KluzfxdMKB7BojgFjmxs0Z+W3NZ5qgWeUglsvssiPC4rYeJbw2dHpFMmryiNCmVw
crQfswJy0TooE3envUqumi/O+KwDW7RGrdHj5bmR3OnzaTIqr/6KCOPXL48UolPz
KI26QSBSC2y3c4UWi+Vbdug7IudPf5TiQl2Uh8LOqQMKJ/UAuod5ZO9ANwWqOqr7
7EQsPFDzAM8LIKopZcMzxymytl4JUI2BzXy/JXOe1wLrhWFarFmi93P6FsN4MM6f
GHyyxJxR8zDuDP7hUE8ibg==
`protect END_PROTECTED
