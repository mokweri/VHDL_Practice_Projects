`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GbtSwfgcqhHuXZgjnv+z0/vcnt1dr5OItVGu5C4glU0dOpnBEHsm7Ge+LlBtFVM
Zt50JnOM0BC3w+wL51l9bFZHf+2c2unwTSFAsD3uwjmbe9Q2Kn2wEHjGvoOX2Dxm
ZhHAZO2iOT3J7sp22EPN625C6VVyzoeNyRtF4YbkGh+UckTIzCnMJPJKv2xPy7eQ
KShUJOGS48oAsF9o7Lz2Pv6i0e1BsC9XBlcOyLMD55bU/+S0jVoZroZX6EPapyvd
rW45cIOmkNh7xjI+8vTA3Q8tkUCdg1VPkCCMXUn3+SewlrQglC6MDbzIzKZnorPf
ezZ8PfxdQWG777P9WP9qUl554TwsNhDMnfBDdWeRO2M=
`protect END_PROTECTED
