`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NmC4ppHnMVC6VH6AEv3PoR7gmOqU1njULZHTeAZFpsoIpNVzVNqYvrsbZLdTrOEF
+kYvqzYIa6FVjmJl01W2ttGknSVA7ezyY+yq5yZnjPzc5Q0hkjjpM5PfdbPdMFVU
kgiWgkjIYPOpfIKjxxpdag1kz14ALhv8+vcL0V5kLFdZQETHGLpxl9if473KAVWk
hSptYcMcVmGsStBikRUt83qJ74kI+SCgd4eP434MsqELcuBpheBeccorLUxiQJV/
dw2DE7ppswQT5CzdOuAvzei9CSGlTS2LiuCUqlL/xNbnNC0psp6mQ3jw1FTjwxum
Zgkcf2TDYjrotHKl8lHYeDlXpqA+jzRiWbIT+CPO79pPDLwCGOkaFYII/m63Ey01
Wta8VOQ1mPqJctAa7NYp0hUP+9cRGe82BtSQiNyF/JJc0wZl2xF7dgdTdvDFezrm
b5V4GtT/WJ0kFqpGlRlOYjwqiTSQA7pTvT0u2dBlGGis0r6v/Jt1n+/FINZN7vKT
IgRwzTRhWaOniXJ8BSDSvtD7rHG6W93qn3/3Qbv/U2NpER5vz/e/IRM9Z/h+xyE9
SMlhXMgq5PJSVDHIqhlXexNhN/BTcYxFChvhzfVPbDVX9ocNDauuuxZ6rY+Mlg3J
ds7IkOhyBa0AddN6KB0SKj4MbZ+H2cQX7fWO6ubOPoaJ8g9Wf6RMpdShzdf0EQsz
uhhnlNOqzIiyHFn8fNaP5gEyvsypac9HCbX+A3MH8GTI8zWwDcrtneowkmA/cb+P
js/jwIYWttapO2nz5urjX1U0z3+KuO/XSOSGEprG1iqIdYEn41uQ0a4szxvahoi/
HKJrXlOGjYxzCBQ+TF5N1Onxa+O8NPwC1hA5K0rm//DKyhnDeR6bEUbqor6bFFT1
qANH9vnQEfmcTYCKitFTQLUUrWk+NnLUk/CG0eYsGBzlNtnUgWfza3EXg+txu9pI
/8xqBGPmbxYEKH94vmRZ/vKxV9DO3+SYKLa9tiiq9B2Xk6pdSC8qvgsN885C+3nh
cq6q7MhXtE9lT3KGaxHV/t3TlU/U59VKrwi0iZeXZqJxqlC90XNGzUZpZLPi75aP
olS0e4c6Yg7ae7AFbyWm2oNUIp9nc3nos8iBuKMVzGsvVMf8rcadXODChlR4vpMs
hDd4EPyGLpeYM5uF7lCIpkgbRAElb0Otq9xy4ka9DuCmig3v2z1FOBIQhlxlIlUu
MBzXx11xHUUQSceTSiUSnuMjBvvydou8bppsF/VNu0zxzLk2/ENfOcZC4YBd2Yu/
Kj5rh0zs85yMzmk+gSeUOQCoX3Fiu2eiIUtOtMQwLBiVKifhENe1VwHcou/OlJ4q
s+7BCYn762jq5Om5S5folNr6QLkDsH8+orvRfpwBXWT6oAg59omYvh80LJyB3/fa
9Tp005t5ppEGT1pzeEeNzDFCfoZXEwW+61qvLTP3+k/o+09PhTokaEefoINh0U0P
DkbC87I4A0unAgwjvJpiKFEj26ZyNQftDk8S6Ax/dHElXtukRdeewLYxfTWXw//G
q8WCLpvQfbDQo5GdfGwzXQ==
`protect END_PROTECTED
