`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IJ9Gj6IYKI6CRqew1bjczM/Was9PP1V3kQnyim3smKF8Z6pkpaLqgV6DAOfoVXZ
CstLyPYf3diYQ6Q4HrSOinwJHs926YMc16+QC5k0+ocU6WTrkdAlgNZEdt1tkokf
hgWki/UGNTFZrddsebOo6BXD/QBaQjDHJ+N3VZNIsTKbezfaYF3hTPVzggThIvIW
7KlLI2emcPccWGj6aVS1HXbG4S1rkYzi+4W416M3GRFypEWaMyGHeslwowFCafsW
PnxPgRNjM6u5dJmanjc+ekN7l/hchT5PlWmgkW9IlbibH74ih+dUP259vdzv9tVG
bj8Q0z1UCdkTkPnHVe/Fn9FZRwe0p0zecrOzCy7KnM576KXsnt3SKuZv3reauica
g9Ee6OVZ4dlgGIQ3wHcOkKzo/l580YRZuQXMHpqW85Yv/HLmvhV1FqSRt9YEgPNE
KXSvwV5DWLJfEbuP98Ke0yDDuz02NE6HopdyWNRjdqFG3uBfiZq9jyIb2rwVak/k
LqZGzMgkVerwc9QyoxN023EEArLAWxIIyFdam4qbUy0pHFNEX6GXdGf8jwDyW4R8
IthjGvNCGtFPpODnk5GsdJu620LMUDvbhYRR0mBU6HVFPUpqDMGR7pkBMFxZwf0a
PrQRPuK0wof6h6zjHXtxpjbniY7blaaKBSzGJdmz0IBWACfQgWsl1iOYHXtQ7WX6
geyRNWq/3NpflRkayec08UclVU5J0sJ8JiuKrv4+hvj9nz4T6jfWjcFnY0nwTzZn
`protect END_PROTECTED
