`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkVGqp5y+o6pmDDJpLJ73iQAB2y/tbAcB+FcIVZsCsl+YTSpeJJ0UMOxQqwP3ohb
rWp7P5jCYvolnx7tq/ewT5snfwW6xc+WIL0BtbIliLOvUaDNXpYJSW8rCCSC91fb
hAp1u8fbnVtIghHJxErgYfo2VqBDsD3k+xjlldjArRyPWY2HN7W8Q6FI0X4hjhTz
ewH+Qv46rAh9pmi8idkunC+jO6IC+ad0d/BNy2TDWo0x3wEgkHkANrm7elaWIaIT
9EnZB6+UepbRyh0RSPUeltWX12yBDuv2Idq5hSATS6iodOrcpkKOAsXyTdbApC7j
zMJPFa0S1uMJADE/abGv/3GFDpLSg1G+o76CalyiYkp7SnlQnnQZ7If+Tk/9X4QN
iex3V66u4pz7/DjxtPTbML6moSupAyFQkt+wFhPuPjTdQ+3MHvDIzDY1uxWA0i0a
lg1/jXMjjIXuNBHdsWrg+AEZ2AUJboiQohq0A+Y1jbgEiw/VoFDofBb9zU0xs2g3
dWh8m8cjt6pEafArTc8MKunIJ7MwBJ0niWYjoSzMOObi2go1EiCylK7RXF4irsOY
MlytN+bA61bMA810bZyUvPbIfrObbWopcvPqs94GSeHN+V2gLMhm1NIgE+OUined
Gp71OJ3v1MlcWQ44VO4hW0kLko1pNCgvKSF9EzXVInLKdO9Icny1PiwG8rka/xc5
Bg1kLdneEHms3apfvTqkW2WHI7LehnqWwfPnE5KMuA7HvzaWVXgwNIG8PRub7Ti6
O0QCgRUSIsUSXdR/1qGEci9lPPF0+0mwQkXs37bd2shjrCOje1QuAUVmWmYFaVog
guY7wcAq5QvcIjXDvmU3OtE50Iie6+CFrE92Ipi4FrG7iXLOMfgMrgzeGpXSfFlH
0HNAG1PA6D1uxoMgh34FdD3mSSmGHm4ABGzPEu2ZlWVQkRktfUKiKFS52COTx2JC
nTGDVjyy+8GS9ufFWI/7ImcGd7V01yATMS7MGyb+XxbsdCNsV2bSZb5ZDcNRg68I
4Pa2b1k/sAQlRP0qQUn94YQijlc89OV4+Bn0497NEzioC842x46D+NNBage3MJEg
aUXMAb7EO0TnASDN00Aw9SiK45+NoruLTL13ODGqoK2Gew0hibbfNaFkFbUb/qVK
AOT6tVvUJUk68J9nXRFTGoNbiz5CHmRkCFVCXJDOsAKWekU6wmUoos2krfMXwZ2P
52llG3ojPWFbezKb3kuDKdOac4J+MTGDlwZERQoWINCynkr8SNdBoXAhuKOflUBn
le4Dnew0iGBW+1wcR4sfnwZW2o7uDuIFbLA+f6dQF4NnqbARp6Hgciw9fE0c9u+Q
IbusTfomSbeaDlTqSj3+O9qVppjilh7LE0QW2AFPBzO2NADWbiQRMckrEFsDSRAt
zA6Ac+1iDRJWhXwe+t+Oh+GR25sMvpM08KxOZiSeyBtEt/ynv5u/5nE17O+JeFhV
3DRh6v5vSBZXdJJfvgMl9W8LkorjogF85f7fX49rqvv7pgQ5a5HaRKgNlY3dqn3T
wVeDCxnNh0EoRfNbLIEeopq/tlqzFacC+iXqMOg13yF6TDWynCxauuiO7NsFKd69
FuiQ1ZTQ4aXgPVqKQKOy2kQCx1CpinKhR01AgZ8104iLN29WnKO/0QTIqWAscWdj
NnuGngLHj6L1Kb67823m1U7mL1RbcfM8nhmBlXzLVbJ9gSOeQR+Jsv8ArVrA88Kx
p3E13Odf9iUFr+1qxRe7Rn98timgVQS632DqegsyjHqnyVRtkKTYT6sMu87+XTgv
QGNFrxeaqdPCrxd9Gy9CFgulkes+DrAbKqwOF7cc3ZhZGyGUIW/lk96kFdebxwYU
jjSANe1lOpKxce1ZLIPhgeb4D6lh8WV3c2AEld2LiFGe+YkDJ1Z9vhDFa/7a3BFk
DdugSTUz2f0bW9UwHaoDgODy0upA0ULFFXjOU2/1/YXRu79j/ev+FxL5PwxsimaJ
0dSjnzvtp4+C8UBKOKV5ReP2/Py09HAPAWUl6sR+QIaRzrTZbUDIBNcqm9BjV1LC
ZmyGwyfR4q3iEx69ZrIvgs64DjJKdmN+N3ekyoOdcw9nh70LlG1qVOWrB3MtB6lN
pNHV8QwWSBBailvUt1iRkrOv30pgU1ou2hTB/LNPWeSvUiudvsLSVaoJZAX5Cfrd
EoW90NWF5oCNUnxyk29JKMWF2dJGWfm0Z8DYPMU/XH8vNvAmIUvmlZP6aw77zcCJ
VwTyOZJ2Co6lSHWqg5ShDD0rfH4E64V4XoOvLvwKl7WPZnDBSoXatQO1ChNhZzsb
gDyZcNpYkl5ZGnqylxVBv63Ne+SlPIi8ooEoxRZ5GYfAI+wAvbxDGyR43pTp2sCy
u8b3uhYh6IDfpd7+jQJeg8FRpQ0m2dThWqg6U0OMytShfuE92e/VjV5MdrtLcMgM
s4X5vY2Q8RK+vfu0UYovKoPNqj/EcUKHfzeL/dU9HaHt9qL1I9qB0XCuE1hregFo
Vs956ofugMwBRBT65B5dqdvF/rPjT6ZID5UYn/NTF9FKOA4a7RWHoicdy5kEh+rT
xe2T+xFkSlREBWws+wzKVhtmeZQ9yR4WHLwk9Ne1+iXLERtxqvR3qOn8o/biVitD
YCkuqQYJZjaOVqDN9LvH/S/73eWafUFAd+at4DyL2jk7dmyFTPJ28Rt/Cj/6cbFm
9Z6lxGB/56EXTvzeT7cqaRTWXsOffFi8kl5MmEkp0Et6dmOwELAehh7N6jDcmYVZ
G3Zq4mYqMTA9aU7WqSVeRfqVgMUTDO4AvZPofQ9P4S3pEMPhiOqhVEM9TyGfGnjY
8zk2hCl3S139Rw3PdP85xvqouwfZt83NkSiic0/MyBxzjAGTKlyJWNV5pNLLpoVj
ED0aR0S+UyEqHHOVizTRPBlvDvivOvET3aWw+M4pcgKWvl/fIOnE5CnnMKTpkU9f
+gvxywvwRPEMsLre6tZ75UOervwUyK25/S9gda8UlxzKXialxw9I6HDwDAlNljXF
czOj4BOFjU1UlJNEJbaJuj0xC8R+y1mzLQcOCA1nxy1uc8mb7fKiwGyDfcZ/VE4M
st+X3DdDyaj20VuV06caLvOpH/QUD4RYWtJkI/rMgufTWHiRnrR0mUIkpDrgxCZP
FVtpiwkGItH0TScLcWFzVb/wzBIOyfj6QWbbOIX08uA0kcXfy4M6Eldl2r1OKdit
hGpSTmLydQQZkl486lyRUkQNnJ7+y1L6RsfUMvhJzOiBgUkgvSNoBzz2yJCIzi/s
/V3tehOmgkVgKMMb7UZAi6ytCJFbFWAGtFXWMuBjJjlmwQvwM8VnlU3IIpSGltC9
FCgmdvatWORcfNh6DZawG8ljHfDkthF6HLoaQTv/Q+AiAfeyOdxt84WpoRScR3j8
Tiq8yRn93npM/qon8ya5H9OFdfNKYy5LCc1XQgdw1HA2d1p1oh+sBZeVp+k/t69m
nLmfX0sQuthGgPYQgbz4+95d9dWjUj2dON/Wlf5VM2asGAHJwVDtR/dxwnyGfwlf
mPDNu5AuFk3y5X/SEN+DGwduAENUFQscphiFIIZQX9+lbuANHGDHcPHED5hIOMTY
mOWUda6CDqzCcT39hawD0/FhLR+XldHEaLd9aUnwBVdp3NOyDvAECFKUKeXf3AoU
hkkayG/yG+PuRRbXnkZx7rO08yttq7fkD+1LgMOFQvab2X7U8uef2L7ZlFOenCC9
QYNWfJtz8dkFDiQYECnA3xPcwGRKEyaIb4z/W6OzMCjPdOnMTzQJ1SLOHPJGHyVH
FNDbru9iOBaDfwHw16NW8k5NPQ+skYOrVL8AFKRe2WchVrLVT1kPx2C2QU1/i6Pk
NGCm2DXI0agnz6FSXGsxVAcPonKoNmmLyR+tTg+cKfXaWSRU/8w9qGFETpUqG4KI
E45flQaDmeRnSl70cl/ICBlpO59iyUSNA2ubMVEh04DwbcBHgobMPO28TovZ8+vE
2mQZOCS65EK8FuKF0lkGOXx+Cd8NVCom16MCqyBZhMFJJ8tf+KWlABAvXV4qM9Yq
ItTu5ZKWXB6Hm5xtOJGD0RqGtw7JJa83z2Daz7n3Wi/oXWy3Z3lRAyz2bXuL2wr6
KQgGbuPC/CUhpE2CPAB8Y5jg6hjtZgS7pZ37tVQ/aaG258MB+86rGLqKeeGdLPry
17SZOurqP/IWcD8jT5s2yAjihXFvxjaTEFHpQgjvxa1EzZNQukOVPWARm2DQk2Yv
+uh9fqgIOAkAtCH7eyAJhowkd3HFkYK68Ylo+BI/zFv3SYdJpUOgMuVOFtrxAjJO
sbg7bgFy704JJ4gY1O20wl0Naj30NIBim/LFu++jg22PUWkdDgOtwgAlIk/XjjSt
PnAxkGruADgSBkD0h3aFza57ZLfUs9kF4bFhodkEaRWiSdaUX7cD1/DrjXc4cvFT
pNzK+UvRicOXHyMRY2b9ub0QK/WajtpjLDU6/kqxx9QqB3K6oOypIeSNFpvVDY+l
`protect END_PROTECTED
