`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4IpEDXjUPO4qLSvXDnJQiFIIUU/Aj2+5qc1JWkEaFPfqnDZ/cRSRdGdXT7eXQ/d
OrJodmoUYvSORDwy5Yd95Qa3BS+EFDlkWhNnrWaBfVs5UTrCHx7ZSBNerBzy0Qve
X7zYdaj00oHeQUCYviqyC27kQPKVGMssE0tfrcjlLOkckQG3fRUqCwxf2xzrqkWn
FOS+yNbS7WyEEB2MRK2a3p1bmmgSY5EKkGLpqvdjTcVREf53/cuf8pIegjbD4gZ0
IzqFRqV2jsmncFCt1WzB6DfcyLI6Oj7WIRVI7SnX4LfhV3su+pmu1mPvHD8agAUL
SqmgexrWL6e/aYzmcw1+GOEGOGUBBv9LV7yFz+AHprQzZLqGIuE0QZxBA+QbD5ec
/SRXCNfbCWsCdnux5TDe5cVebK6XhFEszjHEI451ISvgEBfcNq4+lZgrXfA8LJhB
YDHyMwaIJF0qtrIQGXIW2Z1d9/7Cjwcwx6Ue0+1/a6eb1SpnF29IQgp53pm2rAyC
A5joAN6zWQppCNticRUuIRkdjH5uCZnNKHaT8koA5Mx5y65zJYDUxrva0ZBzVfZd
fXQb8Xf0Z7BjmXt9B76S7nc4z54ho/TEO1JUMA2B6x9sml4rKupIgkB4KaOenL14
qieYv8q3I5t6EdVLKFeHXjL3hiwOvFNDXoLxyyG7+ZP0oZVHT/4cWoBiF+PcWVmV
QWF14WrndFTXK8zU/XMgkK9mdKPJpceE1kpB2BQomnWvvUyuBVSQDzArdt14BZHc
B6k32zi4pqYrcwMcQ8AE//mN5AQaeT2lfGLotXTwWiNknwDlANxlRb//FxQfms4b
IExzOqiDNWWYBVYbTh3chSGWDthY5BT+vTekAlSlKoH5i4QhspKIiVEW18oP3Tmv
CmyFE3sCIwlDwAzqR10cD/3wD7AODvK8ef5pjVowZqkIYRO2dvlg9dB3JPppyJ9q
g2BwNgknwas7CxO447VasYW+O5Vn4YlRBfVJGuVTe2On6YLkLQytQMPIIw4jVjuj
tFcHqVMTEJeK4p8LhFRyNee/bs3KVfJ53sgoiuGjPXVTPZY8Orj+m1rJR8frMo+C
GrS0tSwgUQyLh1npUPVZAtz0ENrza0tmfxU0bxOsGnbrDyJnhusmky1vhh64rw8M
D9GM6LYTpn4BW3Z0ITBYGxHj6LDOYPUOfDgd5FIwRGtFrmnLeIhZiN2mKTwqcV9u
BOccVzWgeFyHue3E0zeooq40UaisUk7tHnWydLDQngg3KkBKpHBI+zmUnVBEddlv
`protect END_PROTECTED
