`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/+F1uLxsRXzK4WJVVr8RaKfKyCFUEVDS8lgSS106SbHOSQ0GqWO8U7L9dAKDvii8
Nw1H5RQqzqVDctMBCzokBmDPTGCGj1vtpjc2MdfbMKnYygSe3vByERuEMbN68SCD
XUwPpsZ8iePYS3helaXR3s5hFIX2XNPxInVsNybIaf9syiM2QAtj3mS1uStUS36N
LY6PYVB3EnaD5AOLZlA7cuE4y38QZK629/UdfeO6FnR0Vf0siS1A6v7fTbkD2QrF
CumKa2zKFLfhyT4wx9meAm5C9UylU+LpFWPMQiVYqx9hgDJKPEB+IXjZFv9yU88s
p4r8Fe8h+J6/qmfxUynLZiBk0jurjxN9ySx7eMYUxmgBKDcet9TJ0uung8LMUuum
aRkca4O1CFB7S35IPC+WfvJT4vWjFTBzOG2CK1mLXkAqa15NkcgJ6x3NHkbs/cgN
mh+JvTsG8rnUidO/hkUGcI7isBsJfgdM3jwDji4jACw=
`protect END_PROTECTED
