`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VhGIwFxtmfBXertirO6b3adFnqT+G9SeotZTjBQS6SDirv43uK763Wjv4PE9HE3S
lf+1Ch6gHlajuJkoyF64binJ7aznRkpIk23FfdemK1n6r1hJ0af/4nX4WMXIdXqo
Z/OQlyjoOeUUs0h18VyQRMk2jkhE0n6uuyGIZcxLNRPurLGrLBtMs0RLsTI47hVx
YTnmHqGe+mEJHNd9Uzm5oO0q+3vb4hIJEW03Gy1wXGEPmD9IHePtZDhA9LAuNQAf
5wCUMQln8hq1RNhatfK5XPypRQK5j1MnLTWpZIbJm6yOCUXs+2EwOk9jPfCcCetS
h42r+PxS7AlK2+BOGVFjXDrd5QJujhXLOsTlGOIWS4GiknqTPG7v2C2UR6rfZbVh
aGBXmaF/bL+PsjOr1q9YlNDS9uqrAiEB0na/jbtJRPLvNwAIdvQTs6I4rqXwKRgC
8Zh7I7WZkK/TzyIvXPcOnQHTcpLJUBibxKRwxSdSCR0oBj+CnTpUGsYeh+J5zjNf
UPjXgWLdq4WKBoeghOz+A5tSAFXVzrjBbIgBOvQb0+P/rNIQLbIzphm8VYLvHOyz
OhPL69v6JL86Ku0HtdG8/ALjTu6qo9608WyWLqDm/cd2wfmSpF2uSU6O5YnVpjAO
hTiqJhB8g/J9Vfmj8NbGOBjqP3IkPihL0p5c8SjTLAjo7J3x3k8quWvaxGwHhryL
xbuQ3B/Q7x2e8bvWL5ctGUPa1ON+yWcnl+y8SrjXzT1q3WwmozfcB0zjWI2ytHfS
GSqBvwSMbSnrsG5o6c2Ol4BTuIV1gF2aDwblkClZnFPWawga+H2K5LdqYo1Caw/C
Nsp90HFo/HCzgmuuQgu/L34U95iSb5aptl7txmXyRs1MxpYm2X1YRGuRk/rMbLYO
q1/0CIj5yiC58xJa5nLMoL9J9dF/lDpZ4QrmAJLNL4ro62SjgPFhllvF2G5iKchC
2DQsYwKO5vImlOTOne/G1bfdUkt9+2WEGrWKaT8JdClnjNbntXkXtTDcfA1mNfJy
Yea/ZfBxByQ6LJtYar0VPE4Ssh1nKJMP7kEiZHtVUQzmwOpIyk0BcsgwmTz7g3nO
TB3gb+YDX3os4Q4faoo06oW7Cdw5TUPrXuAcv7oSoLbJsDgrG93OJwfNDSbe+k9r
DL6G9IHMcU84Os0aJqwYCgb+auVP0tYoALhX99b4uABV9smZ8XJptkkIrdMvmEIF
`protect END_PROTECTED
