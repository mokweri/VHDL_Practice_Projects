`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KL/oU35zjtE80xBZ/hG908Idtm21p4GyJ/0KtZnlSmO3qREw3YTKcB0B+WB/uadF
IjhRpUhEXUrjMh6UmjzV13bWkex9U+yJ2fWnqOsIoMVlkkKE/3IMKw2F0FDfX+8G
dzZOX1DZSr1pRolxrzMkhtQTjKu+CmoUaLkV6b0MJuN2Jpzn1hhsq8wlkc6GmkHH
pW8cyuNEeVYicT9W6IeFnp+bq24XMdM6y7ZW6/vV6r281k0tGa4MJYXMvLNir+nZ
7NQpeL+WLPNyj3UKc/Uwt/gfUjQw6lKVTv0pAVETz4TqxCEVP59HRdsSzsAFVDLC
rF0fUgLE4ANhgD285FkEYkw2UpefLqyABoAxUJlcZEWilAiLOdst1FxIBMGT8W4c
klZP/WqIUhorvuUz27PphHMgTItMExS7RabU6UuOa+XZiMFhne/CS8ml9RkDNRlx
k4TpPnvyhyVCoDN6Bpju4suvf3B5BKdfyzcpzmKn7YRTSUw8mGud/aZaskXqaCuA
+xD4GMu7k2Zlu0SKzBVzngyrcIhfe+VHtKE6olbm1RzB3GR9JNB1KgYj2vJKyri1
W5aZB1kkJKA4vD68LxldZGsZ7pu3lv9M8fwqnzXEu4FGQ7CXJWok8c6MR7PqoGEX
Zmw4yuNvuGq/+ORLZOzd2s8PbNhNJcEw/aeVM2sdDgxEcRB8vGzLedtuWwfVnnjF
2yomQ+chEYhXMmLOJXKQsfhWaawNm6focSdalntToc0EoVqTWmLKwliV3FaiD/zm
Jk4HP9dyO7ZeO97JLoMCarQeFBCRvtkomjssqd/3dLJWicJ8HihQc9NDiBYqm8e6
2nvvkfs1lcWZ0E/32n5D6aKRcB3LHu2kw9BHxjc5JtQ=
`protect END_PROTECTED
