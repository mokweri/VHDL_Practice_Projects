`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MMTSSN56gzWbo8iLCr/9PG9+hBkEbDluFW4j/lb8aIinqCk9bpgNYV1FzalUeL8q
EsfmuXs+uivvJV3vJtD9G+HLlZxhNBX/rcEchSJoIBLj1PK1HvtdW+aBo/KfX5++
rtZrkQMLAKrlug5U4l61QPnWsBoz0N1YmU9ca7mQoXb5wD9gEd6rKeBYICqU3QQc
oTo/LG7W9KD58+E7FwPM7b3HsxlYBfzzkK4z7HI2LoXKoSc8gyoADGh2oFs6wdKJ
W1+5KNmYN0cyxl1YtyU+LAvz3uxi8w0MkpVizjciQAgncDJu+yoy/+xzLraTW9PU
aZnD2wStjA5nisAmljX3/POc7YtGV7G5sV663eM2GeaUe/nGSyBQ8SBDwiLjAhLZ
MDpy8qUSjleDWN8vFXLTxFA/S5eGGmaCz4ZAVzOBG1/y3kgsUTDvgqO237r7fVk5
xfj38Y/rOl4BvDUiy3y99UUDEF09p4UMuJ1m6Z3pXqdFalbIlrW38vRxKuFg84MY
bhMcOQ5/HjpyAiW8Sozbv3IIno/5T0wjV1dOZUf7+RYKnwsnZTAqYIXxCWzQ+wMB
34L9tJupzF7NESqeZFs2m2/y063edLDVB6uI51eSxUbZi6TA3akywih9BnwR4xqg
hHGkvAdDIYa6cox3i9enFK+ADvDAZN9dLqW6BkkHmIK7WSN/nCvUFr9KiLS6KBz5
FKUlwbG+3P1zJdXZXuFFGqfA52fX/Xjx4NgcC9mNZ2c8RDfDhO3Fa+QplBApDMsV
/LadcElu4WBBZfjeZmarhSokAEyuhdbbI0FSz+ELxioiizUxI14oZzmlOLyBaUIK
smBqjjnx5t/+/SLrEtMVbFD+H+EqVTDW2DO1YBpXk6aNCII3hj/WQ6f9eTin2wWh
7GkxHnGng1GQwGb3KKph1ai1Hs3akmbUf7EOiaVNCcyjQTe/D3KSaeDXrhyUdWBe
bgHmkT3g+QHfZ6WnuKgyMPPQBwtn2TXfTdBCi28PPTZQsHoW7NV2F9JCY3KAJjvY
wKQmShzPscSqBBMdVUyzO/bbgbf17yixOt/LBNicMKSUhtSsVAlaX9lEHJ/AoX0I
5chKFtIO6WCLhfSq7+IhP8tfgm8FSueIM4lUbykFX4YbwEnjn4j51U3VE6OcaoxF
+Qs0IvFYErrIUeERUCkYEpW1PGSQjwHvsINsMniUEavQdnl8jb3xCUfSjVD3ht+H
++bpOEVid4WPlUgpNoyuFvxX4T+5uqlxT50MOYRw6tU=
`protect END_PROTECTED
