`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bgWSN9JCuvZzVHNtV7mIT6oPcE/QMV/tFkBusHXKBiJaXX7ChZDAC0vtckDYbSj
1XBKJb5O4lh33+OkStjgHXj7NI/x868txnviVTjn/C+TujbLVU0Dh+zj0B61/2jJ
biFwVBXGHLol7PH2CSqDW4v0RZaQQ4A5wtIQxITCllLEaUNkol2ghsA10lIjP5TT
q0VyoESf5Q7Z9cCJ5wiQClgkfzTy6kJ1AVVe/M6sDbqAJhnlK+KfP0i5iG1elXWe
tUB/E4egBLt0BcDQsPdypsXg2QYWMbUc1QNYeTjtN245xgDuUVyk6HXmhzEur738
o6z+tujmYQQ99T7phvDc0Q7IdBknYL3N44g1pIaFnSw21QYav5cX/GQ51RJCE+d1
431S1JPF2gROCJms1/4jQ6XuLeWNcvwA939n8+pzzIZ1pqsFYDfndTRZLKZtmkVK
coLSa+KKMtPs7N8ns2ZqDr6aHdesUh7LoXIkHyZBYZ5MdNmBqu00bmVmVAdf+9s3
+jhPkdUm4lpIIuId7RKJn04XXNp4fRT5WP7NJkOMcNXa9NbZ0clfUlU5ObkWguew
O/xA8ghnFYiP2yxmIuDgKvtFdFDtA04vNx82ohLMzEJjMLIepcasWltNQSQlgPNA
BL1oe+gk2cjtWmjiNOV9tkcyO409c6bi9auRWp0Ite+NoS2sNzPC7JntPc0klB3V
3NEyfldTKPkeYV2aM2ONsSfwBOM/ElwFsfJ8DQiNj3lZkcOMDmvj1vQpyJHaCuUf
atJBac7t07YIwVMfHK4mY/RdEM0iDhbEwGcHn+UVFEZCgCzaxSSpnLwr/ec4mVDD
85VN7hE2e0zXqrtdGYDXgnH28dVoSVrgG67HK+D7zIZvBXQACDuZ2tTCVbT1dDza
B+BK70jPoSd7NSmxu1LX10Ng1gz7NxL5tKWtKCYBZfSjtaXEfMYpycuNDF3VYtFF
T0vUg9mbnT7EHLFhLNGGmmUq7+/Bh9XgwYuLRw92zS4kDtwn20S4AGjPZipztKks
V3N2oEML4tJ5NSJn7qSGYoJq++niWUlh9iNRiNBSg8yXVPmRUC1zbrlN11MazRNM
+4ZgvFXAPfrTxe8zYv60XvNW3pqjTjESDVGvHoHV9TzKxd3bYQW4zBNItLtA1b3i
ncbxKgrZjAKhFj8sRXTjGiL4zUMwvLQL/nB+ceDSrX171Me3X3F3/B7AniEC7rqG
qWbbklm6jEGBujk39XxPLr9hf4/6JqsMBEujPDCdkaNlYnmHXKOrdpkAKRLQBaR7
fTVBWfY7vTjuQncTNxIplj5LKSVlaKT/+AmTFmbebiOsCSMYyrkz9HcjzLxYISv5
jOeWTY839hDWNI1eFn1fOS5w6lYbXG/Oezp9KgxmvZQIPJ/NyI4vC8tf/OrwoTpG
y+epUpXz0Ytp3FXn+TE8x6Df8HKnU3woeBU1cKYinaHwQyg9bF/AfAde/DSe5O8M
ColDsp3KIGhADe2BSocaTdWtEIooFcZBbtDgqyRVWOtjeHRDow1ZL11QXZmw+mSz
SRD2qXUGX/nxKkQfxKxRUnrz1Ie9dAhH0U0sUwEgggTZ/eo5/DwdTf0QOIXTW36A
Q2Q0+amC2HFvwlNPhvDG1yU1QrNTJnhfiKlp5eW8DwGI4VZkxs/BknQ8LoxAljRr
eKOWGpdKc+G4CsXwDFl/x+whFJFGERpIXnkNR7dmBZtrD/Geh3uCgo0cWE5trdU0
0Iffw/gn2TDKPxf4NkOT6GLEkj4VLfId1jfUZn7/Jjw0iPFpcCe4wFI5DSrCtvSl
DdGrBZJFg8g9WgvHuBZPNLqqxg5JVRlygnQnYgbwOaLjfsTikND5pBI4MKq3WrsF
/PlKP0f3e9BvA39J3XA5pfSIjk7cMxOP1Gex0b8my6Sc2hZdyrQBY6wGDlx9LHY/
MNi1dSEYy/+SPEsJoYhN7w==
`protect END_PROTECTED
