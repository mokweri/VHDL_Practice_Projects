`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W6YWYWMzoWAp6AFqutYNEOPcsbtPMTrgadBPd8/1Eqg2puCe+y2/eL5pDQUd0Q1p
AR2KaRUZkxnz+iER6n7L8QRGt9m6P8LO0soN4Skon9FZJUTPCDAjKECNXZ0ZDMrT
FLubGMs8h+cz5u0RgNyIOw401SE7DnlmTixunNKt0R9ry/Gbt5vYGG9P5AOlPx2P
LsBs4R4t2lpAg66flfdEdNb8WtS0Hr/bUAX3SF0mBkVjBlJPWPk/3Nh3gPMB49Xy
gmlCHNUPaDxh/qxjHaFQHUhulebdX9EAqoPy38HZJ9V2ctJlWJB1OW2h6c0sCqgB
2LLy9X4xzqpILPYLufhTxmaAglE4ZGKSpzFRl0NKZbLCM4czLvmSwyryqpfzM/hN
107cv36VAfDfthFRSlK/n8K+Q48ATRO83P+je0Wb4YXyf3OZbeBhgHgs+9Yn+dID
taf+fmEdyjkoaic8aONoAOtBrx5q65/q2qw/cdnq3UhfZhYAw9wXRNIec7ab+cbw
ExZSWuRCncJFGqQRDMs2X4IyU20PH7z88G9x5zSLaS4Bn/3O7JzQoFUZFLa048G4
AVmBRwIO/HkmlIIPBz8YzL03fWw+q/FKGDw7ljGwyB1MNUCxbu7pqD4wfIPQm+4F
Dm/IcwSl8nQTc1flCo43dA==
`protect END_PROTECTED
