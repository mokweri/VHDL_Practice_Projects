`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O8PA1pS/gWQF4UOM9g8sjD624d0wavdG6vyIx/4t0R0bcU4XuB7h77ty0N+DGuin
gWr2n7vvBuCyDl8eRDE/DwZBhRTskQSOBTJlaa85zxDzVW2tG41kW3ySfnMr0o3n
54yWe3T6Ualw5cAJVcIt6eRmHNNT7NQSwaGXsEt0llvmG7GGxZzI+6ze5l/Nj9rf
YTeUWRaHJXUEj0wx86Jtvid2INN7eudodEwlevfRZdDWzdp7zPv726qX05eT6I46
nvmySHYy8dCNsow5o1u2mH3kxFCA1CE86fer9qb5IzvHBPHNE3iefA0qtz+O4OcV
Y1IukNb9qDNi+hk+C8juJS4exoeuTgy/uqs0L4dJqzZMO8idGK59zLHEeRWQw9hT
E4ZgVYFV+Hb9B3XR/1ahBlhQ6d2pVVN7CmTrswrHVAXnc0pwYX9IKLGbSUwLzyNR
Z8gUtFyT7eqTT7zU2Oav0DxqnZl9Uv3fdMtXrXNhz4bpIBoudG06/mq0Co3RLevd
LY42C6OpbjtIVc+Rejd4L3en0lI9hc9fqj3AOc1EPMsHLAisoyhzbnrh6/KEj9K6
+BWCpW7kFRDFFqiuHtjlP2OzstiklnI33spp/5Sw8ZzetEta2D4ye5lWZeQSA7qv
NnPLwJURfr5VDvXqUVNZOkowAMzoFw0TmSf6ezgFIu9dzQvoUL+tEk0raFf7IQtD
gcxRVJvGxfPtHg3SfvHA5z8mHjsjRKlTconOWCqTFY139NWmccBSWauDjs1HyqCi
fnr1WwE2jp4SK8apODNTF4a9ARkv5LVWEr8NLGP/tcDawVGtoUv7F/Bi5T/PtkVD
P80meshMXTfDeUEt0sY5aq8OrWQJXeH5X5WpFWf00HcSy2TcFitztNuQyhnW6/20
bhbSQ2rHiS0Yd0hLe/vK5XmtFgm6Z0Dpy/+Ejeec6+ZKfAFaI8HObJlcbXM5MRkP
7+Wl5LlcQpqEHyipWPSge8GI+06A4sQp/OHfk08g55cFORFWACt+6Nkz45Ixbr+k
mfwbvTwS4gs6RHvWWiergoRMWWxpCsi43xbEVUYCVUIeY9Xmr80L8t1pVIg7bsLI
JYOb3fVEZEC2e/i67P/84x+mC3bQV+vqtG7Ff8Jv1nuMc5n8nmzgQ5IoBw3K9BhD
7xbhBVq0VED/YPyYZDu5vHAtSI5K7g/3rMiZO/7pTc0XuB4CmEWpeHQ5vaUFXAXN
UwKHULx384vnCv9QJ4sJ+lCRfsbH7B9eJZ5K5+77Egt4KYSkSuH96aQ7h2HEVL0R
nlc/qQujm3NLIhkbZ3YGZ3D1UvARbmcyM2CAkSR3FCn5+ntG+nLs528Pq0WZfxG6
ZzLfaV0mLzf37XthnRCJN2l6Wof0tiNE1DbqMGFxYlCxNsNOw2k3hxJjCtntTeRp
jRY5Qa7tAzkRNc3gfwXMYBifcQ0qslF9UrpU33pEwYCoFTQyGqcq6FjgvQrvEoWg
d6liSdNJv0iMYh1+y17GQVejPx0XVqb1T9NO+xWQJPZySsBild1en3fwse/Rp8It
mW6IB0Vmb/skJEHG8MpwI8Z/1v6Hzua9+jv64qkD0kgyywtrzJcaQKkWEvAb1GKb
icY1qWffnfGukWMuMli/IuJ/kFWwD5ttF7mbET3rShUlu2CAYwFsdTruof6ubK1Q
F1YwE/qNY3/XM5BdE1cTcahHy38r5lhmYp/PFaeYLLIFMkQ15LiwlrNFV6h4BIDa
uwIw2OgOn+U7VyzwZ1zzaksUXD/l2moG5XS+8kZo2aKOiKCpF3+NSwCsuMdb9nby
uBrPS+cijP+You5yO3Vdg4HqWWhquhB7d+L8HCbmPmkIAyZiSDlvs54lvoaORNGD
ykiDIdZ+A857AsWRus1r0GlbSw0+3+h1TVj0TI2OV0N0dhhdWIDULmgV0HqQGLZX
JmcJyd+PhMT2Yl6JeBhC1551gPPX0kjai+XsJGgg6R/QX+MkHjiDYfiq6ejFPPSA
Sa1z+sHDhZOlujdhsD8nwbzZZyIlYRUmFlVwt/jPBDwXFdDq5DYBYFJastkSUArM
zQkPv41/NhskgfHD+SPyXSHkx3iV8FKXkGuZtUKR/hH2ORt2omRtOJcZxHVsXddK
d8FmVOoJSyIPPiDpsEJJDkE2trACbihsQMRFmZ4q+0vyr/vK49PvaKOjwOy7Tj+Z
Jfdr+Ez1dNF4OlhmZ2nfCznwiyUkoWd2TMLr3eK22cOJezLN3xfE90J3xDIv8OPe
Zw9w0B8tYZxQHqKGSsjYldKGAdRFJ6Cq1ybajNUHADB77Y4R26xli4MOmMiZC1Wj
UAj0o15pihGPCwCOLsBE1SwpEfhJygFK8m7vpTdGiDujoA8EipZynVcmfWt6ESuK
KzJAtYr9JG0y2Op3+rZRfT0OGRzFlyhaBkKNGYkkZ7AVTodUoSSKl92IsH6fr0cc
GnvatzJ51DF5y28UMTLNAO4C8ennPonGQbteidxFyxdAQEoR6v/SXTv9KzoYutzR
nvD/IfpTNTKe6TqWWrkIvOPfQjd++49uZ3kt+fV+L6mZ6DGxeOqVS4aTv30+37Vu
3vocgT8cnWfiqpf+bn3NcBUOuG95TAlSJQBMXy5DDwbm9FFV7WShQAr0UPpadjW9
QC8x3lYnb0pOV6G+p/ApY1wMqPl0qmFu5FdpfCE9NCIXLoP9qPnmI07awdQyxnMc
juQPzqYo/bQswgnbx2p2ZMqJRxSC7nMGZZHn3i5Bbij/WntVw1MJCEofCmgoKwh5
8HBzDJUYSHkPjxBOGBsYYaFVFNJ6E36N0dYlv8vMGLI/UY31ijrfDOHKAiRvNyhP
vGP4CsBtUQkS0Ts04/aqVsjrmOTROTd9yL+obUweyQmozrZ6uVGgBQAzyzgPZnE8
MdPlQv5BQ5T9ww/Dp1jMJkQbEQt44imv97XENDkJlzeg1zK41Yy+vDoQ0+OQmqRK
SWRwBju+a2ZU1zlTQxOaLaAdr/LMAJbUCfKYFo/EEE4q7axz9QkmMW02Xh6qDZFR
7os3wwGoNoiLv41UnlRYFzDso934v1MGezFeDbWgdKc5jpzbnxt/vOOrTqZd9x0k
atvrNVIuQSveuN3i0kIG8M4bPfmZS+e399KwITjL8ehxnJnmRIIJt/z/BmjBJOXL
V5z4eWFoNBLDVsjm9G6EasgF1yqFYaGFK7emZr/wJJTycw4ItMn3JM1ZJhOw+xJ6
08s5IxnhbjB8FvrRS9qoQbXiLB/7H2OG9f+cmfDzoHIkCnPJGJzq3PAMKyWFfBY6
GWyDrymya6PEOP/tqw2n14aXh6atsBNum+moSeJU2ChMm+GaKdnS+i5QcMLcK7RK
p5yuk5qF6UC2EFIuthd00OkkZDxyP1vcy55LwJT08zBtO1As2LqKkAcd/YN3NEk1
+ka/mYMdiLWGOXHZWz1XFZlxFbSo/SSNtcVZj3tFqd7bemU/mjty0emN4BlpoDPW
FxOG0sMnPK+wXo/2u6mSKXkyn46Vkf0wU8BVMq8HYJVmIMgP89j3xBkgypmBahrI
QYdAov5aHr9auKyahLqS3kYu13QZ68CAWTTip5bu0OZ/JjD5hXsPT57uka+Wv7uE
la7foIhz0GLgU+hdviUahFKb6L4vmvlFeUlcQPkmyYCU3b06cAS4dBPKcw45p3bL
0cTkhNKqnD6GDm982X5CHCWTF1CO7Ph7KT4+xfkaThxPSmkNedksG1nbJW6OKiFb
1Isw1yoa71HTOacNTgecqYVuk6RQZbhWUbsD98p9QKEcFR3Tsxe7F+dbGMZs+RwE
ysotridZZXRz20VbqKKRL8Uz77gb82oP5P+KP7ytqL4OJn5UU7DmzYeAON4ayOef
dUVOjJ6OY3bE9IFUuJ6pJLkF6COn63EQG5ZEanhvUwZOzjIWGkDAFmVJFnx65ASl
ft/F04zGjeBuTON++q+YEoNNteEFfVaFHmWnv0UhvpbCEvukfFZ4UM1wPtVs8D6U
o72ERbDx9jUq2JEJnDyAFrMa0IPGI7Og7EaHreo3B6Eav3XEA77RUah5KgzOR+QL
gjtJ08D5zVwv4ih3dctu01IIDOK34qXtQLJCQwWIQRO7SwkGDxaPqgwyhOV47au4
YhwkxQcWWCTalN6AM/NCxNvSTPx3GBtibNmFeRyRBACv/uZqr2vDflww4sMy/Ebg
UpEjR52vzmGA+N17XCCKS6TtXq8Q6fa2nKQg0KLxPzJ/IE9rI7hhY4dpl+olB95g
5v9rEXjiSpL5Z9GY43A1aDtrYZBNDXYs+wJeIu2BsadmPQnyltsOiZrjL1Ouc5Ak
x8cFDFjGZ5/kjN1L2pa1WkRy89O3bVvHfiCsp67KvWe8wbi3AqsXOYLz9KV2XwwK
ckRYslT9J7hIfH4UyP0nyHG8q68F+Tax9lHfEUh2LUTxPy9Q53uDx+c6nP1Hc1PA
wErYyLuL6aYpxxNTOjhQd1sQZeTRcsMpYiUq0SixdNeDroPt9dWZ65NoKFborsdM
NDPLU6vgNUUc86vJNI1zqUEnMyrqoDb8zLq2QIqZUn3j3PPvApKl0XFzIEpIYky5
vOLpfmKHH+Fdv2L8oOI+Ot/4u/dcG02ie6tWmY5Eg2KH/HTm0pd2qco3kszsjvLV
setPUauSmDlgRTiFNYCfcPX5NgDiHQzkXowlK328maT/Pqkf0atp652v3bW828I9
Y7BlnsZ+Em8XOQ1V3YphWFefL/+r464JF/r/oCDGIMyjSJDXj1XunJ0QuwJM+BC2
q72W5O1j7cYON4Ensuq9w+/QM+6W1YWWq1e07dnsZ9Jf5G+qthJ8x0zo7IhypFGU
MDHUnTnvY4T0jMqyFbgIIwov5NkRTJie4xvp8zy3QxgNO/HeuDwjtiNgNJGWM5W1
5BUqhVoJcrB7uCoaXoR3TVyxnk7mXPO9UmMofpXv6Pfkx9bckN+IJJf5QKy9zcef
S4hnsg/TrwuqHJmssGBctUL9yi1JjByTCs3xFV6S+cJW0CVLTcacsuyCp7La2nNy
48IM/iIkEclPwxLAAcj/nkUg0xOs7PeKt436Tpj9jP9KonMUhYmh7rFNCcqbOsXI
BRNZV0huoazh9em/62hgapIT+A/KStml9fQG+c/W19uZ1XeecjlPmk8VcOnUP6Z8
59zGb0LTH47tfnS88NUMk7fuqeWei/mRYD00WhKJf8Oq3b+mGRKdYnHrcwpMi/RS
EU4fBBZLs0jLfp9PKDsGmXf075YsT8JdvTIar1BksrN07uPQVnwI39peM/4cw7cP
5fQMiCLdFFpulQXtuZyIkYsw/lYpioM1aV038wfqpToSQ+AmVMqejG7wDSWm0AXh
q/4G6xXJxfmpYUyo9VLt5i3seF2c7LnN/F06OR7ncfGruC3MqqqpWohbmtUI1ozp
VMI6FUSK36rgrcumhfBuSIMIzhob2a/VbHiH6jCFJPDFE6dfdN2/iP1TAUvrC3OH
V+4/SDxPMjA0M+nCZG/sEqfhPwsvD4rAB7/kt4D++TJGnhpH01AVr33zQUKyuANn
P8K0s/YUZJ523BY1WD8e7X9aOsSNBg10H650kPYD5efkM+nkbm/GHWBJTuaIjm24
bQ6We0v/0OoH++q0clfmO+/73BQj79D0LczkJvqn0TsezUA+T6CeS79CjKISJsum
msz2joM9D3I0M2iCzZtIDGG85278yGX2Y4YLcanr2ZN+iHcluu6Ng5+oJ89ugBdW
ZtvuiQ2kQa004HfjcfJSpS1Xnm2DOLyVkivFoXF5dDZ+craaSHbVKxh1vFQ6W/kS
+FgpkRKdmdDibJ5WZoJg7MXaLT916F1Cg8xfbgwfkm+VISP4MH6Uit9uQuf3UEQO
1GvZ2HIQuZ2VltA67wq4iq0qchp40XlJxEV/FvhM7Vk+slF9W+LhMNIXqc4kezep
dMVwYZJ/Av5549xMRXsPzZdaMeL2/CprzZ4UzzLOaslplSbTPt5E5M6j7ETSReOg
fShnKb3t2B/N9QpDJYOXZNVv74qcx7NfX9UNLGC3zwccYT0A5+KENImZt6r42RpX
eL6hpEERgnRKT8hS24ER4jVfQ9wJWGjWh2MwP0A/aHPPMpAQWyg/rJW7qVRTIrGO
53nNXiTSQVlDBe/0tF+//su4xRmZgjR1gl17R/9LgfFhD90w4VSFwOGBjG9+v0Yd
lyTxj0EmRRcQK4ff46Lewd0dszASz0UWWRU4TLwjAFbiOsA5ZIVUC/cbJ1fl521f
voeOAW2TJkt85GxRxdarj3W95LXxvjp1j3kQu9P50EcOih/Bhotg1+IgEZgT0pkz
GrBgI9MOP2cKQC8q1bnhCPYnI+51P9M6XoNOKIkAPTEmPIVwKtGlCy3Ib/XcvyU3
QE/ck4b42LKEET+5WU+KEvmTozOD53x4OUyWIXH4qNpyd6QOHQrtEAXRC4xWNiyO
8kyqiWBMZGRUBsHmXF53iSxhRCK8sP2w9xN1zidZbBBGM9o3lSwL9GXS19B8T3uS
W/Ay4A6jNRAU3Y/eqKrSPTDvgWU4QTOp3W8vdo4wtYOSYFt5ZqXEGF/hemcKxcaf
8CHS7NWb8dz/0xFlUpUbFqWMM32VwDyItO95kZL/5EKJWjrlLByYtS9FFrYzGy5k
78XP24dverzBh8tecRR55I7Rdc0Jlzgi09bBtY3AFLGbiBgqVF4GACLV3GV3bf4P
asm2oCup5YEc7QVJDjCsFeg0/FkR7yDR2hXja9GDZOUuOqV4DdrmNmLpr2Ah25IA
06o9ADFJEinA7WCBeGBUig86IRu9aYhB88+S3zOf5U5PgFvxwf7cJoXWOcYzGNOb
AkWUBCFNJCOg44Rp3/vOEccCGBPi4qNkyugJMGhp0WP+3DVMYc/aKPlb/QJTAXqC
sKYFF4z1ilXVIqdhYpXyp8CrUMeVqoiRwQUQCkD6I+7RkpXzcyJZINg/wp/F0D7Q
3KWdNPLrlbLsWo1pBCP/O/9kcT8kHwaHTZSzIxkEXaE/mb4LZcHBvwnimj2VL47q
bTAGeAwoJ6VvleWVYYCZiHcz6DVJWnvgVoBv7DxROAXJCCS6UH6X6eHq7V72Qc3y
966dlfDSuoG/QFuJgnjfvL0FNh2+Z2AsnJ5pMHJbBmn5VH4oRwxYv9TRZRx1AsMz
Ur0ZBltLFwlEJ7B2ERm/GKwk06GWCoOOc1Tejk0Pp7cHhMbvbBhmcJs5SiKJmu4n
8GSbJR/MVIw4vwNKmzPngoYyphJjfDcqn4QXmgi4oWevw3+lTQYtMqV1NqJKR8Ok
ttY45BwEjbEumBWKGAL7sRSZAQf4vr99ozx6KTnsvdqQKeEVI6BoJVFQcewQpNwv
r7/9TyP0t2gu/AuA+Snobb1zbuNXzM9vGIPgH9YgOMI7MjgPGpn1LnD/DVZxASWf
kx9YeNKI5RlXnvCEfzBrgdw3gl1cPoWKD/t2RWtinT2uHxnf/dDh3joP5IMzjKy8
hA16a/pvzYCAVthJR/nlPiM1nNT9ERno60I4KAvC/Uh0zHgK2n06FphPK+Mug5QQ
117CbSstXt+iFDScWx1fPsB/iVJc7/sT2kbOldvlXnzypHmveQR+AK+Hx2CxsuUi
sY/+hJvvYOUxqm3CDfxA9Wc9Hjn9nYwbBd5msOa1GSoxVnlaluUHlVX+BeVtFTiB
1fRk3H2PO17gXYcqZ8zM5Rv4iG4Reh7U+ae1gffXgIWOnwxN//lxtOUpSIbcgGzy
LAccN9skrH9/M6MNYyOAEgihbLuVTiqJJDDHzTaTHzfrW7Mjs8Ix4ODlUb0Cfo2g
2UpQ/ULRx/dQhwvWJH9/8i7X7yMBCJmSTk1US68A8And6m85/KPDQKU2IqAEC+t9
y5BeBROrOvP69XlRCxhR58grmBHUZzeH3lDQ0UbUdi0FemqyQ4VP0mnSQ2L3iwvi
B/cnHmh9NO0JLzwKkq7Wc7QFHqdTTWbACxv2oAvpboKJODb3RFEkPreVGkMQ8kSw
Y/zPG7P+/XNy3Cfr7+AMQND+3yzq/4IYVLoSguxpA/03+sb/Qygsh8EPLebYt759
zK68yg16sapQhSCt17zew9VC0R/vijtYKfrIKSE5jNokuksvI0iy231iOIiEvYK4
PskjkXbm5g7G5lSkyfeTb9INxS3wlMJO2Tau2Zvpjqm4KtLvgtvGx1hHhk4ppZYR
HzpR9gaW7b65nWRkvp+WATe99PtvV3cF45gFx2O1tGnAG5vWpC/nvfoVxRCikSBg
JTGsV7dlExzBKxidonxrLmTpveK4HhFtOO7dMThLTN48FoSfY5QSbFnK0/tqpQHe
ks0JXtTuffhDdsm9Hcoyt52htp6c4HJCHlJdj4OuxT6Zg47HQ+LRybBIwhKFZS2C
1blFL4qc+64cDpjuRYflwrHhwf0Xof4BBFpeFn8pI0tcrTt3RIGBD8appI5DXrri
mPVFKrcKLabMRGcYRY64nwA1jOeTX8VeWBhsv1GkDtYR72K+dyOVo+NTSZzOiYIo
vrpQAMuZ9qbwd9nJlXmAfQqLZr+HvOv6sF0AVdYS6vx7jRZpcSt5H3TP025KLSCs
A/YPTVRgyjIJhIRd+OicxQVukLz2lEq/vySUCz4E1z77fKjg7OO3tl754WLyTFRF
KfcxMk60PaoVxRsNOujKJ30NpXB8Jp8nWiqqls9QkbhC0EJBiJuzwEsX/4tOfZZ5
1diMpYKCIc0dMHQUpw5o2RBSffcKeR6wT43oo27xDOzkSCuW+dn48a3BKKQR7RsT
MhjMS2KnDJdTADgAUtKn3Wb5nD4JUg4TMy3LRiKVr2im6fhrf/lEiv0oT0DI3UqO
sv9y5/iCunjUK1vo2d30oU0JyxTEMnEQIY9dkmvAd78CcYjs0bSnRXSOANlugdya
12d4DbjGwsq6gHJaAK4XuBvRsDfA++pb6V3US4C0QmXtoMsBRfRsQli2dlTOPloZ
gzTfgDCSkAysaOpahB5uPFJ1fZd6hmWcPXfRIHDs0yi43U5RMLd1fzHFpjOFT8xH
CU2An2rj4kBUbVhUVW7IorKZaqyzmjmxDe+fx++dVr9bWvMY9IIqXiAEd0iIC+Mn
8yxpfRKpbDH/8cKtySxcaEVz7Cjjrys2+x2EYhYjRt5UmXzTHcMeN25hEBWLmt2q
yB9ueS4epIONUw1yqLYxJOK0YZEv6cpkz5ou7SdteBvtVn+PBW31lJcaPVJtsj0j
iXTDlmF78/wtpQp3MW6axv8VWaz3/bfGMv+P3kBYbpqNXUmmho6irUafeKM18ThZ
CqcBwI7Q9c1q3NJuSEzLug37OpafS/hJz+Uws91tUZjgFwoTZ1+L+THNcQKJomkA
sppGm7RSXLQbwYQhTrrL0WNzXY0czxxllUcmSSrZt4/VAlalrEJbeQ5ouGQaA+Nd
lO3/YmoSIGxvU738ybefHNTIEkV9bJ/wXIR5gUdKpY5hNfDN/gS39jjvfMMrSYIk
ppoiseQFQpi+n0H81M6I2YeDcR9kYB0rauegETD9t1GLyNyseOiYF4J+4X9BKAQa
tAZnLAfqRZ+gScP57W99n6R8wjzy5wUDPOYSnuCJrJb/vQvMy5zdqKKSwc0/4KjS
6GANFjVM5fpKj807ug6VFVl913qFN0dqwZb2o91GH3lSYpqwkuKmhn7SVxjH+8x6
Sbin/975srfEJ5m8+42DYpYBjXwBSp9OebBM5/55QSE9VcVRTxPAEg9Z1sgVQPmz
h2If14rwuubOH9J+cTBWAQMbtPMy6QFOxogKWgvgMGAm+Co2g7LZfBJWjZJmRL2/
eXa80Rs8mbv3eMKng8Gp2c2byhzqye4R6iB5pYtKe1/1oRhh2ttUwiIBJJH+KpJL
q7PGDClCXE3JCXMPJx0ZLK4ElNp1BcqBlSzQDn2iIAZWQbD9n0xfuYPmz3IkTaTY
MZ2FMJTaC0iE7wfhq+EWtfPDkG0OXPI/0XWrEPkmHIJ/lbxh8DpFXfZX0pf/MytY
CC53kqrZ3ecDws8pCfhxshz8ESQyhfFBEtGMBzesrY+Xw0t4cQ9TRs7nBez2auvb
v3pqkzqO6bwJ5OKtNz2GRLGw9ogZKjQEbWf+fzsKvHsilOO+w4shuQcGZoeMfB9V
HJTgY7dhcUxxfNlFnjOekeR6FIYfZlKct/D/CxtUvKZ6RzQQ51uadur6Jz0oTls4
IDvUOVvzAsYQEgnPkOCyEIpM+UUeeQ6j5znt/yJsmZYAVXhYBbfXB+uBJnmnCbWs
+9Szm2qMF+dlOyDtf2tmbIfbSSsaxMxmWbZPOPzXYsB7CcY3UaDt6QxCTIISz4gg
1I8wsY/JGkDjDqoarnmA1HPgwRyLHLswhNWktjHsISKMFMcLbEHx5SKg8TUDlldA
Pjp5vsBC6tTNwaeEzNbHAfFtIjqnHIuioZmj4XAYxz4vvmvHrqxvfSdCA5jynlSO
zSWaaZk+mtEZeLkA0nGpu6bMRHe+hVXTySlNByWwE2XKPFTRW2JafXKC0D66jSW9
x9yTCkznUeCk8MFP4RCOuWWMz3bP44GULd0UTSXKrsoPka+bb/o2wRvB2mEJsiHe
pBKYLcCBJb9VRcCMDXO+NxpSz1Kyn2uTOrrF5w90XxRsl9fy24CaxVgK1AZwus9a
ty88EYu6p77l8VF2BhDQI6np0tipmvJ6u/sCn0iSaQgIked17IEyrnZD4MfMvwtW
xNws2pJHM29camkvC+1usAaYrM4oL8MsVUIZwpPVPwpTckPKzX+c45bpTQifBvq3
Dlsa1JqCWQSacxAgGItODNbV2FAvaJg21+eXDDDPa/FaEuZZSPNoRz7dDYK6Of7l
fCD/wc3vJ1JdCTicBsxc+1mVb1k9MHnciX04d9Z0IhGWMiUO7FH5DPj47bAFJgYE
vKwQDQK3dT/KyPkct/9sFuCKwj9l90FJKPgWlBog32TxycjpozzE3oYMWdoVFae5
mqqkYhv9xr8GzblAFj/8FGemwdgHXIV7iAGKmLCv0oCTARHepUbAt7mmisq8NsYO
JHYRqGHfW1DVaQIlMXF0nM+xFVCtiNgcIBrM31/RbjnpTk1+1SkalmaUHHx/z35+
8SQORoZl8R3irUB7bO0EuxCYtAzPkyn2KTogcetBmjxl6NXkgx5Al4H7wwthFwKX
Iu98B8lCrrmJ98A4FoYPbOWGz4ZcbGSJFFu+TIKaiyQhmfYGtgVDGMr+rCDD5bZx
2cdY65Z/PNJUh2vgGodNXNGRiV4nLmGDCjecd9fW7iDZyr4RoW8syrmzutIGZDH+
QmjvS0V/aW+l6yGfK9B4vEk7msOxb5ZS6RilLL0dOMOBu9vdNrXEnsaodcrU3t6K
5Sr/HvQGtMSfrJRNruhuV5KVhvd41xvZmJrwhcDXtKwHczUr9x1FZt2QwZHw2/vh
9xaVp58AYqIdWRUHIRstuzZO9WvJK5ymGf0cxdLmRU+apFoYwd4ySV2YwgrRHjbj
1Edh4EWH/5UaGdmxo6zkHcsyYzh1tUFxqGsarFVjtwvdVsZfXVwvkTBwljt+FAgp
R8qyjwlqAOhrd7xbsQJQd15NIMDfGkcAZIza+QKULPutbQOY+44yyz/Qgpc0CyPp
X/x3y8OaIbhVakikwtzsVF3XIwR7mymVqyxgyo+od7Q9U2W9pGBCPBvhq8R77t+K
16b7Jo6kl/JMceBtqvPmW/4S3HxLdk0Gy42LLWv2uu8UHuQoYZ7bGz64i6dColZ+
zM1fnVgcBqG4vif4XAfCQTvo34AGnLKlvVzhjYRBm+DJ3U31W3wPM6tfFRlmeNji
7tztUbkI81pHaP1z+0qLWXJ3rRLfiK/wiiXrZD2Y5aIge2eL1X4wDN+yWNsNEZEW
Uol6zDaRdEccQNWAGC+ZN6irEJ6kvBTRXefWCJZExTfs80+nnNo7XHmfYcN2cxK3
kSY798U0Ag3ifrCMEVkZINC+olRZoVidClQR2V4JJ2/t5GXlXwm76p5qTnisRSUb
wVGgWutX1rgtw8XYYgO4eylSDXH1Mzujxg/qbhZZ2WannvGWJ5gVa+qscc9qi+M/
WR0WdmfXhFl+FwsHzbxw+eqY1pzhRtkd3r/SiP0koCF2d3zPXPHRKaQ42Feiz44Y
2/HCe+/cCjsUkqS0xAwvvnsMAKQ5BayJi/TDitwiH0pAU4zaR1nV9h3vZrfEH46i
jZiwHVUWEWVyCyjzorihi4UAroE0y8Ztj0vUoy2MSZof7SJSW85rXH2gddtmclQw
qJIi5PaT2QacMngu81FvCtUzOaa1VA9Feek7LE+4WNLvzMic9GcQUOC6i97cUaIF
WI3dV81R9dISvWtbSUhMQHMLD44/ZqldMGVfdC5oPOd/WrTAfHl4VSJi1vRpWBsb
NJ0R1QBoxWvguGB7Q6te1yZlNvuQ0CsQE2piP91tn0ubUv0MlI2iA73Czo5eYEsq
FkSC510mm6OfWNg2UypRsVFfUc4YckDi8yuaJNC9Cfk4aenZji9IalcPjrzXuBcN
apJDezHJUxXd6NLoJvSgngQia2hAs+lElFlWsC6UoravspdaJc7mMvBpuy2fkn5g
Awgzbtu2T/JCR/e82FdEn/m8lKTAA36v+d/TIRHe2Q1OgeJpygIn15uPAzJMXNDY
Xe4h+sWu6x9KjjyN//d2C0zqubqwBfMtwz3wmxMDXJagvWVxxQdXQ1YP0Fao5JDh
Qgdvn/BgCB+ZJbcklxQpHm7Kd84UCR2YOdPhhQvev0vH/iJR09zbGuk5eizRoAYK
JCKIipiVsw769jhqKwsH/gqBBsPSzul8ztBUjN81TglMnROtEUNv0xVd5/kP29zi
/uNRX4DbBF1gCN+sgSIhoylvguPAetSbNrOcmPOcBDcDYxLfeJWCKDs8LZEliv2m
8qG4/nUprs+ub3qMM7F2fWUDFBxSeyUX7R3e6VftKzla+7LTp3pxy7byblpNhTli
PIaTAqp8SUxAuMQmHRhOBoQaHUubBtILqD9bNaaASBvqGUz+pujaj+tTNXJtpSzv
C4SjH2PMeNkOzCoyR//uGhN/gYDrLPk8Sxse547l5Dg8CEXsWG3ndoQW5717FDEQ
TH9a3wrMNpPSUwY4btUZEizbi3a94qdMrzioEYz6U3BigW3yJkAjFMHIz7LElgYS
FshSJi78Mnqg2We3kwzg/Ryfoc/wpuoaofewRnQ5ekP0ZhoHm4umlktavtBGnK75
RwXEomj4vyZlbl5CbUCp/hUWZNBiSY7+ldqTEtmgbOHEaHtlqT7+845xVyq+jXSy
oxdqXFog0VzWvV/5MF7XIYLBDZS7V1VuOSOQ29QWOuVy/st54gXoWLWmSVzxmTwn
`protect END_PROTECTED
