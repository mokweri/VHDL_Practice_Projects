`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ApjCkm56g3/k86vrg0vjYk9KWF0l/ac29FfP9aKHZWx1Aem7O4joe7TZ3NTdbuhC
g5hse2vkB4kD/zThAfvR2owzts0WH9BGSOOOZ1TwS7AdRilJQ1rJQbxXIP1XaCka
X6l8V7xkf3hlA48B8m8GH44nJWbX9WBg47VERJWelXyyMqd7Jnj+ql3K4vKSKjvw
FEjk9spr73mlTKWYHd32Qj64BdjYEA2mHsyBWfnL6/wiBBvlIVEghHsMf954HKMc
V7xypUH70aia/4EeYvwxhL2h8qmRaacxwDBygrs0Eqpj9IccNHMgrwZUrHnxeJ89
zTUXTwQqEDXKa11KErNNfZeJqZgRrUbY4K3GUnzxyQGpEtICdzqpB0e4zcEWKMG2
bK0Pk1HWKX80L9OqmYin0wWiHwWOshhZnFp3+riZXKmb2ktAo11ZEV+TNUO4l5i+
sL8ueXkvG2ZS+b/3LDnCAQitVA+Pym7r6m8jM4V0Gmycr7o+krsxDdU6tPu5XZgI
i8R5o+ocRUFOR1d73xHbjX9Okv4KHsoJVD32E0sQDbLDw+lOWxEIzp/0aolsMhxg
hDRCLCSNbxVxLlli0mvZa1iKWP7JUMCd/WaheIkcHkInCDQWrzKlhVH5ZIiVZBzW
x0V0bO4CWaCrbTFAe7WmecgfUcRkzGZ4l+y6Sfozo77QhOCSLDLgKo/zqBAJ75ky
3mvwn1wNse8DwjyH1upMb0SY1iOnOvDGyD2myH/RjDVP6DMSowwQYrodVM9xk333
FRvP/qUPS91ZNNp9pDHp1KLQFsYSx5CgY/3dceJ7vGmm6kqXuuQrfDnpU8LEaprN
CYY5dlRyPivfp75uPVl9RWDPVlZPcUULXRkYLY70h1NQDOWiuiExp041Vn/60Hx6
14XKRbGaDj5AxjwVQLXcV1InvVg03A03tNxS0GCSboU3qJoGJhRJ+pz79pif0O6E
cNJQTrsTfl55qtyxipmnDv8RaWDeEPsOb+kEQhGcRd8iJvv3fXrVhZAWTasHs8DA
P8C2z/C+c7/lVQMRgdjhMtKv/EIPkNBnvaZQ6JbrZmp10D7uJufptMBDv3bY520l
HI5lDcu4A3xYPcwcTTJtxPaBJ9eUT+eAcOE67EIRJE839VeVy8a3wF8k+LHSujsk
luSgaLhHec6a5DrrBzCBe51Xq0U1TT9l21UbUCPWHSUwZjBZQ5OETsZs4ydl/X4t
1xlAfI8gahcvWH4xXJp5/4NhaQdXeAQ84sIkcUlNOO1okgLTIc+zf6/ARx8eCHu1
EK4OyJQ+DFl/EvZHQPirlPAcAOBSg583ALGJUrKvqqxlCtNEs+yvw6KJ0n3jdWIc
G1a1Rphj/x0pGwvsaqWR7Dd4sKm32O+ThFb5TISnXgpFao39CCQytpbxMxr0apwW
gBWcU4jVKNGRIFcl7Q6mAa0y+CwUKkYCbDoGhsjr2D1oQ0sQ66oO7cMfhezhcWsh
AKwD5t/qoESTtPrRi9Nl+bZQdVlzk+Rnpo8l+3rIUdRN9H8Q9RAZExOye15TSyMz
BlgkBHKef0XupnCshskm8ExoN4+JyYwpyBlCNAwuQJmhtokoMUyYwHpLqQPrwLbQ
NJOi/fE7K/PHdaVXKbG+iAYiAVLsV9XICLpE9kMmd0ELHltpouuKWf1L2Gl927CS
nmsVkTgu083e+0EgTAAQpDB3Y1+ry1j0Ub9DQsh9rOuMoJzyu4AL7O2wwQp8BC9H
jQ32TpHuLvO/F4JzwvBfPwQFT1G8A0fo7Zsw6fn68s5v5Zc5en019GvKl94j2tFF
QAkRMvYe8ECoGntK//EzwQJfyeb22gO5rIP1PW2+Tg8c+WEJWnt8R5mG28uTh6RA
Je96Y4tn7iXSTqUTM6eiw9YGCNwOIctI/1LTK1FIoAkkXuRkdZ+I5Ty9E+lHtYhN
i2gHVDGeMfvsxn/1seopwUFAY7JZMS4FlA8+OVlvbabXa6EMxaeQTqfb1Kt9GK9M
qjRHWGzS83GSGrZgNO99LZdCuOYPSfn5ON89Qc8tBnb4Bp5/9+zp8A3MLtGuM5J7
m4tm2Xwfkje8St1YFAb9IESFbzCQJUZ06/QQ4njdq6ENI5M+P4YVgsmWbZiTDq8n
qzT8M1aru2/xwgd/Zew9tOcLKeIyPYT2+a2o2lE96hscNCQKcWrZSqItv96aiwgZ
UpyHKsPqk1v+yU6E+dZ5lJ0hNVCtZoZDvDFF1b8asT9rYDwCs3fPCZex0hEI47u2
i+GAEPU4FDHlKVuEPWxPPr1TcPyYxesSj5s6Fblz0bqALekelfpAlIOQw67L8YKG
N+UQfvGj0HHFXMmRg7ueCrMMiZ3eeuvDJsrFjBNGLNO95u3+vKPV5+qHdaZaJyej
qwI6CzpQDBw8ZMDQDQp0ISFIre90pye/ZMpK/0hGmcMYEvdd8me24hgulSONU72h
ym5kfUF0v7aqgAVETILJlVUpIJT4Ex6W9yFyVTB+YCd7QF3dvQxpXj2TvkHZ7IKa
wRFXRjGClNrXcQYsDmIKW1LgKdMzmjuBVmK3papdzrw2zedHUIJN0WDBvf2hnK1E
GCvKiufPvoDu69toQYJXPQ4H2Drc+ALoUwc0m8UpEU+GtX0jz8ht45aVWdFNNYIh
CkUpAELAMQpCJTJTs77sv74OkNQbFB1e+6/UqpLG3WajnL0tH56DgmN0lsuuQIQl
e7CE4B52GkD8v73Yv7z2Mfw7hjmJuS2a8LpO3OVbI6+qzDfy8Zso9oWBlqCGx4mV
VFg4ze3FfUbCy6Kvvh8yA6KURJhFGf/Em5UO8d5iDeW8EHMePkWoqP7NV/41cBDm
4RgboV/4pRFlRcpESMGiktDreOpKhodlXphvyDvQ0Os=
`protect END_PROTECTED
