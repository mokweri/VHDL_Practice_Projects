`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nvZgGTTDsCLROU9Y/1TcN0IVOmZKiKVRkos/w5WfWshR4V6C+hr0PecgF/DfflYh
FCah0UTKLba5sw+ZJidt1XWCEphtuzu8MzIKakJ5bBoFcxx+AHfn3C9nl9+J6GGS
yCcZCJHWl6rVWvIv4BcnVcgbetTXBi4Xlu3G+t/B5eqpwuMYN+XXKlvgSbAbOp02
qy0LQkz3JqrvoHQNrv3/MWbfXLijqoxMT2GAJq7uCSqAici+eVvP+ROsrnpDMu73
rB53OzlqgdxAlfo5iCIOW30c7iDe1WRlYQiivXS/nvHprxgALfJcUZtlA14KoWT1
bFD6aNogYVhW9soNCCyOFM02g0uObNsQTpPRlXcCWDzq+F2w/7+ZOdAm/E074rKn
XDe0vFB8D341on3fQ2RwAJe9/Fr08ynK+kKi4ZJXTrWxCmOY0ZWohgv6rNMQ2Swh
NXkbOW8rEDgA2bQXgQRa0xCtvoeI4fA1Ep4R35jLQpy+jwO9zf5+aF8kDqihe45/
VjfaUhOmGivJsu28TTj6VaNqrQ8OyKTb/R5O8deK/VUkV8qDRovGDg5EMpbdSLXz
XW3NwdvdGRTAdKlMPs0Drwdnze9PVp4kxU9dwGp07ccNa4tVkQaSdowmOqGvsrS8
Jjqu8Pz8vfvzINkDKcU1bkj/gVsU7btC75mhBVNF60Zn6ZfdRR6ifYok2dYf8qIE
2sqiaJKt9ZKQAtgCiqW6vBjTxeZHMn4wlKlIjo6zpTLhRwFfFt3uiSciqDNWsrXV
W1FPA7K+5hq/xwSKuh6eZI1RWvvkF2Cz22NEq67hIPp+HlEAql67MFLONCFxbiAR
mMClwyRhrYgO0botlH/V3xpNWb74AymP6PDD65sgcLOltoNbwSLhN3RSY9j7sD+6
9sdqlWcfRc6QmUaa6kDjiN3Er79OCwcHCmqmKE+tCoLkpkLWT/VDPk/fZeCQcSMd
x2CoxGfYkfkcDwvmM7dpSeg46r6H9FPUzxC7ZKbQquoKjy2sMZIDaOWM3qIyiTG3
WvyNAia7eWgpMXnabMgLMWQaTbByl3TX/200I4AH1kbhMJwgzbTPt0LhVvnnmTnW
`protect END_PROTECTED
