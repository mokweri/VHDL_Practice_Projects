`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pui6yPimQQfaDeJWunDUwCqIftmTaE0LZXUJcW5dmvTz6YeMmR90K4mc/WtW35GS
Ka18ATkmlZiFVmjzpRuzigx8wp+EAvkrZ5DM372RLqnZothJ/rClxI9V8V9Kb3tH
a+kRVrmNNcF4cijUGWuC29hBZdsCPEafl96J57E4lLKX3SzYsEgW+8GAviLP/UPM
C9qN+Eu/LhHqFjeOQW5XZjbBfyFDK3jOZwh7hp0kTDaCivwgqxjoPxyPSO9oG3zc
tvDEPd6ll0xAn+N6ANbxDoaBFGQKYGRpMnzmzemcgLHNtRsT6/2dxqJw+CHDJvxv
1fFZW3d5//8yZC9xlv6uyKtdXO5CYPP5fsA2y5GE3UtFqbP2/bBJL5CWYQOczBPG
59b4dft5ErEbBGYpL0IDo/snrpu4T2lE+yYmgbFy5hBMqcMRZ+6VOgD3MuTCDfd3
6T8DgtLI8O9E8R3IaiBXCrtZAaL1hodmSLlAKCPIlli7zrFb0dKuXGsLNXVUyBuq
41lmFzo29k4+zIAjT+HQ1Bw1+P5/hliOly6094m5A+132YMf/xVC+5Nt1JRYcLyq
FV6QgfR9jXM+jnCm7D0NCA7FIkGXfmfkoMemFsr4p1/hd+ETXcb1pmBJuWlS/PQ+
LaeeMRwHuRigYfVW4etJJIvGYnlW5rCtOrZy7oMOLsEBQLmGyXT6tOQ3TSV1LHnk
zYQzQ35B62XZHsrI2WmLuot4bW6VaYkGI/LgkqxSmcmaWWGjR+nqLzapz6UToq0A
ju0uhLC5bBVzsH1NML9qDUzKwvCpn4q6i67aCPFkQz8c9YTn47ZHuVeBkNoVW8J7
cs7okLOF4JWsgc+NlcQxynabEnMRZT7Xnvc2St+cbmbnAlzE0YDmmfI0YFstdxxE
G91msH1lu+8OjoyTvpjZfVXIJlw2CQoGeix/5RSt7WFKaceFn+AoMgoaj5N2qXET
9OQ6kSN0JlHZuPcQRzWnIKwrlsWQ4mCWucIQUZcVaY5xdAS/fIvUWGLCHJlFSeIL
RNnAfnar3yS4wsovsOt4SnbPpqV7xg5x5FWs0xGuyRj9HpfVCxxwEnGoG/IEhrqz
SHlxRCFupo+vBRr/2kwf+9neC4hj50o2y0TYyin9qbtVe0E1iXpFwJ8/3aM1Cgiy
zRR6r9ecwenZoEDq1xyZ9Jce0w18RzfD/Mk7pa+YOTu0UL+I45zB/C9yKkYUFYW1
zSXBph5T+H1YUZbE3KjtIT7cPVFliE3g70L0+zZCMm4nukOE+wkbLY4QmmUIJ5Ig
wjhay9niBS+v7xY1o3YriWbeixyz69Pfd6uITwRRPybb/9m5P/zluLEupHOxrb/e
CmxKi2bGWRb7uSoYRboDgfGqfP+lR3HSX7uKlDB1sn0Xm8Nby+4CKIY59Eu8F0RY
XWwSIBTzTalkK3MNzfNuRIv2afkVsvGEyaB6Mp/U2dGQWTHDSNL32Th78eHwoGk7
m3z55n82P6GsYsHQN+NVJ1YKk6X7VeIc8zXvmFdaV7TKxxI9zw6/+qmIsBO5ACck
wf/kMs+ZoeJhZg9FWIrXe//jEraXWakB1rAKZrFnIDfWYqXttqRPQQ4y98Pf6DRr
/dnJyddEroBOGsu5shx5WKG0ypsdt5KSnwAqDiXPaKfCuu8rkrl89LRdQ8KQQqpc
KM3aO+OZREpkYFiRtCaOUIeinPoacu6DdDfu6UiXKKYW4yWAN4CaS+g0iTfrKON3
2KPLHTOGADiaq5+QBzyG0/y29GI3TLgZ/qlvt/qs2EWKT6slfzhgG8VKi/alK/MX
r5ivMDSJrqYNLQcK7cz44TlkyOGUNdjwrPCmPCHTl5qRm6x2AihIO18WhwVEOoyP
XVQKie1mC7olMn/ANiay2pxqUWca0zXPxSRVfONZjVnFlunamirHyW+tBJjg3Az6
ALdSAlbjsmX5C6lNL40OjegN+2IWZXDqd9DFcLz+apaZrNtYNEZILir+BXLMciQa
hyW5VDSA1+qDHShHhYnlj3DBJaN1exKDSzSExK7G/HtbO4DP7G8/m3hi9KyALkvc
QURAPIvwzwYuWNusfwGNQss049UvKz8PmH6d3UL7+3IF8lR1RCg3NzylinllWEyy
K9hMOnqiUryYf+KrvsN24rzzzvfPvd0wp36/RdjmSu8aan6liKsmgCN5ZZ50aL3I
303AIl+w/LUJpT/4Isq9B4sPwbnuM1iCBmMBsTptHIiam+qmk/qaJPqwRhNxKH3s
XA2ZeBzUWiKrNQrbE84WbyAH/KIYxvVQ/hN3br+D4kog1Ob70+tsrfvAhNg9O1Vr
x3BD2Qt5jiaIcmLFnLM4dvLpMqVL5uqrSd6f5XYV0tAslgio8efhHmuRWTXCRHX/
qOQRFXGKyffXafGUEzrh7PNhOlVDB114Hras3HsP+IKITh1WreNgHWxZ6ePDZXDT
ApIuMa22BQ58Y1nNVf1r3hzm6hu+oVw2r9cDoyFxBTQ9Z+XdMMc9iC9WVnaFXHB+
xXwhl2w32zN2LYVAoUSv7UU19cyRt2pxlQiIjmm3Cl5an7yWUficdMNshSbu3RlM
1bREoWqEy1AS6mivitM8TA+GYZe0rYciUQKYGHgNu86w7RrP5o9TxIXD26UOSa0H
Bokj5GzPwHCU1gyZ3LuO8TQE0oI7nMpcgUBMD9416G508NH39HUmYIiJxDarH6Ih
H6EpyyyOjyA2JKgm9q4LPG/BOs+Wbd3xrrZZqq6UqaQV8arsPLUuSOgh7wyX6gFA
1yz6R5FolVKq+90SD3TL6aiGorS/RZ4qhy11xTZIbNbbz2VcEKB4FYRkBolxg8w6
Dq78l55oNH1xf9nktFyFK1N8q44XjD9l9P3x7rTcUrSYDH/x2NQ0TP1nEUzrP9LP
5idy/yRr5h3V7KSmIC59bXEi6ItXk19fYEMmKCyhue3XqHp4Jdtvlvft/we7WmYk
0KAOI7VcFDSjEWs4ECrKId8XxW1uZV1TanVtaPDlS/mMHqswLyECBy1+q/G03ft+
szUpa4IAWgmmbZCtdcJIShZ3tDouL0IKrNw0kc5vD6W2fBDDiEmwRwpPJOTOatcc
XaKAsnxNjHPstkAJXMbqCCJ+UC1SRTB6kRzAumRKhH83giWCNzMz9cSIw2K9JAL0
t9wqcVlX15dMYRtBeqMxuRveRjSxB9GuEpJkubPxJ4fc8r3xdqMdV2RuDC7kb4Q3
2U0BJwAt30OIjyO7mYCVr+ToEW+cX6QX7s8ZhinCiGf34s3qauH5L31V8VhOogEy
33JcMJL6xIkXy25Z8umBOXe1EvbRtggcvmz3RBTzbb+Xni2Bs28GU54INF3ln8cY
6cx7Cdkn+kpNzQOtGDbKeiaal+U9cZKSNsJnkaMqBt88ae/R4XYoKm1wqgpUVZA1
X8z/wnYbZMrZKIZ9qEXEcd4cqSuSIb34KevRCyxeYzmlt2vG2nitwhPOouA9YnC0
PkQdr7WzD6wUH3y9AUrHixlvd7StcbcookvcdBy+0aLshLxhe3PutDDN5y3uqQd2
OxNUvif/YZ6rPEtMH7vh1dF5mlhCqda/2Q01HANbXC5vjB68Lwp34J0JgJ0TaY73
MSUpLAP6NWhyQQ35L3kpAEYe7g+mx5EIZ5XZJu+2Bf3V+L03cwj8sD5RSW3UFhSW
70tWvTUFpw0aTxRaQw4VNVxryDV4lGU/mX5XePC+HdPa9lPfB+sEtmWi61RM3EH2
tCCGQP8ThTEojoXU4AgR7MFq610xOaZ+s/UY0OjeU6SqCcijZDRS9fV/+3cIYDS1
yuQj3kNYVxFXMKHqS6fbP+LbKnjqR1MdZLkYqHUBvJPlXtjVO1DswUsq184t33TT
42S/YOK6rCALb9LLG2G9sOBcZs7ryOi5fZEiPsDmLuLt6PQK3RbTM5tLjjrNgXmg
Q0zDMFDaCjYn3yBRFP9tUlf8CptX+fLcQF22CHfhD8ZIh5H9q/wAyIpBimfcKLLR
+uFaFLc6ewI97KVInCvjw/GKePbJ86VhhBLgWTXjCxuob14C1cLKvP+P7CVGOdCI
y/pDu9LinRAfXi57PQuQg1/DbSh0YslbsmHwD7FW0RftCb5x9jEouXwu35S+Atv6
VGJiRSIDcZcNWPLmQiZ/vnSODHYmepDeNWlXxMwXBN6+xrGjTCda408hFtXU0nh8
iJ7hICSS8FI6B6+ygg2+HMoUPnWZID25EQEsMte6r5lMgcLTYmt7Tef/y/mEIKp2
CKR8QfRGGM6fHBd7OGbV9/+fSM67ICc7sA5/HEcQogIK1bMHE6WEWk4vUSneTED5
oqnhPnXkO4TGsR0w90yY9zP8Zu2GzGY8+eYeLqFNN9ZmdasusUGmfw6D9svsmadf
oUm8HhYQbquK7GsOBXDA4W+LL6MKTeqyvxot8T6+3E4B6cgrBfEQwVQpigtmCyRw
Dv3FQ/8QpnY/URdesqV6UGvdngjlGs1YC5SmTlPlhCI2UJATGvqD4upNxke9RxGR
B74oHhK9Cf4hZCNIashF2Pi3/yuVh0flyicZACIW4Ipw1MsWrQFy+f4bBn0TaA9Z
uLIyCYhOBzzt1WEwn+e+tO4K5sYnepNAZyL/ldYvA/yVOp3n4rR8n+6KwYqAmhuR
MoAOyhWPURTfTnAFnfzFu4TQ7Cicuyf2EfIWG6Ws6X8way7n7N5II1wqq8hc3QPN
+l2mGxqUMri2lliwR2DsjfhfGT4AQ0/+g67m9ROqj0Vq3D5wTbKs/nEerQP4Wlku
VIIeGO8xStH20X3YP+X/B2Uz19cQA7QNBxf+IvMsUzZQu7gQBrNGLmWPOe8JILOZ
q0o0RF9zCytsUrnDWMirczaMndM1eI5mjBEQkNEDAcHVYMcWMs9oS0bRFdBeXr9T
vVg7j6vNfUdKSqlGvBdpijITVug72hjtYuryhEbHdga3+6KLfDaVoMOGg9eepQ7u
P7Mnjb/E2D0cjOVsaGoXcA/bp1c96XzxqiktgnbdpHakVs15eyc+M2MU9HbMiSDM
Dk9SPaLZZ7Sx6tpdJmQq5RKnOqsTReBhGIdvfoN3TUiCAIAzLPFGQQeYyp0d5dHF
kk5Hdt7kFjYz+1FlZ/6SmA==
`protect END_PROTECTED
