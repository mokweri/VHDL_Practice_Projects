`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I2Hc/jciE2HT2qw4Dd/CTQ2h1B0NFLFA3tL0mjRqJ9qxO+1rEszmlOAYrVrLLL8s
4J2HPTWQD9Z194f3Jdmfzvb8rJ7QKY+wlUpQ+lTxX05+c7MN33/RjVsqSiySU4Wd
ljIJCisTi+i5z2Vbu3GXupVFpfbGG/TZCNvFCRapJcagfdzZlqfZRpp42pGmtKRI
gEWukspJRQOqlUXd3JPBg3Q7IwY2AAp6ZxLnRvIQTiCqJJbSsNo4U2x7O3hvLgxH
Dq5wFDTDpmTtTBOt/6cG+XywNPtWOBolaxifqGq/yzGUu7ytjQDCtREfJYqK86Tv
1E82IsNpxjhAM3tHMgouZ7LDwi1gxyY90Z0L/jtO+fuinEBlxLRtkSRrlg99G3SF
GjpJn78b46BiEeDRn3eMOqLqZldjD3cmgap5hvZinDeeX/UXm13KSKGW56dijB/u
GnGzSVRNSaTlyixKL5wfLXO0rpDE2tR4rTIujpvzkgriIwp7fQxSuDhilCW3CFjg
1ssuLygpypFNAvGsC3MjIr3Uo10ukJfcvLftCtHTuifLXtzmzFwTjGYZLODi+gm7
gTNyNZ3NCFEuAsPm1DZEYwpo+tzeF8CtLAfiw6mPTWUr+Rwu2QVW468ih6Z47SsC
xLZzw1Zy2eN9mgiQFRt3+BjbkP761BOn6MhlY7qp9I9b57njC2Uz3EMooWqYaq6O
N0rTG1U2yR9d9BRqRqc8dcOLXBuZ8CtUspm4Gh9kYbLD1zut2OMVifLrA2bdr9ZM
fqs+BE3869dAWSmuTM/HVYDACHqShPwB9ZEKz+pDtjbVu18E4kWvPmi049DOWdy9
mpRowXV6enihaawDbSM8T7MPW9eshHBUwNRBDirV6tvC9bxmyI6Pb7R39u64zXhE
w5+2NLBz9Gajp7tszbARuGJgKtyKc9+Dhd2tn42pxuwlK2UxC1ZpUFml03yLtrGf
av8H3zk+6cG7c2/MQysYiX6aGw/jpaJgKpCoFxyd6er7Fk3OG1afMUFKr2194Lgo
tXfbqJRBhpOg+tNvdAQ2KxotaFXtDvW1Dfuk6hLiOqYn3KO4mU8Be3Go5UZlnd6z
UDn+/E1kUP+CRNP7Kn9uSU1SbsAHcN1I7TDQAjUU+5Kuknn2wKGnbRHMzfPp7HJA
OKA13sWALLZ9s5SH9o7Dp04tEr/WJS8HAnH1NKmTRQ9NCVOtOVaxzJ93NUYanvY9
SLZ/ADnddh/HTaVdGXMVj9rplaVB6qPHveemBkN08tw2EUDL10Gi8WLiRoFuk0kI
q+TDi/h39ytNghacC2XIrqLPyovAdvBqBEWfkvjtjHrh2xXagb/13Nuy87IygOsV
NwdnF8lngo3gNe1u/OLBj4lriYLI9S1Rp61wU+e9BqOVE6jOYEsn00Fo9NsI4HAU
jW6hkNB9nWQ9LNI31xJLnOJu+GWA5TIONMmyAnmLoYEKRi5ptsE4PUenlTYpqCQx
eKcXlUkfkoJ+4TIbfhvSjeDTFWWLrW8tS1PtJtvhWNkSBtpyrLkzrnpU9H5wYkgO
qNk9ds+nMRlQoSttaWAdso2AxVuGiumqlwq06eHnssZ8Kr3atRjyHkSTkMLjdQn5
/OHsFraeWnZ61cgMQjnyzPVK0zby6lo5hhgUXqrWbaUHs1aFAzF1nDtpNLO95kfZ
oK62atzGdINginwuvlchcuOuTu6/PxYep5LWo/ghNXixxMJV3kCryTzUWELXknIx
mjT1t7v2gYblbkoxGtZn6Wc1m1iOwYLZ5JzLZpbBlu0aqW2YeAERbV+FouXnduZp
PUw7aikhlJNSBFty8b25zOhIeLpXnUnf6/E32hPuZdOy6ZiryIHk3TL5n5jDWyGf
af3X+8s3JEr7BteKU+WM2xGaf/RBzOFneOymCPoOJrPTGXIehUKA/Z3CgVAQDZmQ
4rTtrBZq6Nan8bbaVO8MGphfpFbF1DcJEfCSUAZMWMO4hLnU9ar6k3wVZXfWFhdn
4pPKacPrbys6C0RxLVmoA9K9umY65mjt578sLdw+mYLWYctODjWpK/yUcclZXCLV
1hZARPmjXSltly0HoojH1idtXF3kucAZlsyzbln18ou8fcwoi8RDrNNg1/JcjSQ9
vsvLfArwuEqhMuWyxGnG7xWIqJxMICFM7/Fh+KRyuJzobxuRSdGPR/CyFQe56JH9
WlRNnXU0knB6KQrNRDq8522CJ3PlqWxsVYmEIW9+RjHGUcPVhJhTNUgLT29Xrh57
e91PvUGYke9hNWF0iOAeBxWkb5NxiuOpBM0qSbCzNgNYoPAFM7Ti1+Mgyh7oaX0w
iHSH+wmctIqSH3nsYhRFWg2evNuXQBpPt+hJJzdxMkowa/BvKsHjzSh7IizCKJ3Z
UJb+5zfI+98eaqpTsrDBWmMPl9WzPc6uHa3LNrp212s8kxNfLDeJmAF9Mp5EmCFP
4zZIu0u0opaxeCnZpTDrLld4mNIFUyjhpuukhbPeqZHK5YNfkVCOle15R/e1Atf4
uTA262rgOWbc+XUz2qFjvdtQLC+QYGiCveXiQHD6aWUgyFEfr25pS8UYxEuGm9iw
908kq/vFRzp4yl2ZUaQ8IX4paL1C2t+zXKtpK6Arg5MaMRlIKmxnBDK3C+V5obSz
v9Bn4jxbLMnWjk94cJjrymTiWF/PYn0kAQjlVJbTJovoWKexIJwz9bcrTAzCa3ll
yzsjeaNwYOWugFJuamFasMReb68PaV/0fUwUIeJO5Vm4tMNvsygXwtMC+nJP1pVa
u/YpFsqQ/QfVmY6PgYen1KiZyt8yIsCS4WZE16K7sOHIu4gQhAZdNyQYPcrIaREA
h1qGMUEjqzJnHLfRybo2bKNS2Ma/M8xINfSgmc2e339fZyJxZ9iu/W1ZkRBm8+Pf
36jN3u5yMtZslnw32MUzqVRW22I3eOUagsiMTuz9azqLsoxaj0dBrvZt0gtuZjcJ
9pWel4jBRl9vzT6tdD8UZreqlShc8rQbg1Pk23Z2u5IUROkSEw3NAZlL7RoIdUvd
DrdM/5dCaJMaA+OmooTXje0IibIUW6q4F444rtpEvSVtj4udkp0pcq2NpB5v/XXk
TREsZ8vAgr8i3RR51FR/M+ybCaPwEViR/A9tRpKFz/sw0LcaqORRYgtz2B1JyH9d
3xAfj+iN1mCYulf3lr2TJfbVoms/b2SEeYE8oh1w1orlkw+bvzpJ8sFZweIorAdG
J9DxJJ2QPpJeodg5E3ZW69DIvcgX4fKLEyZbAw+taDwmBP1EIAA4G5tu2Vx6mVE8
HTk+3syLeBk05Jr6rNruxLD1QBL+nLJL7FdphLV3WRmSD8ZpQjy88irJ5ljZejzX
c3RDaOuqU9PosGDoX1DmLHbc8Nxww3aWvEEyUKCTTgjgziqbgOUtS9R5fgUAUdMK
ef5U6uHNCXuHTkg/t6Talbs4sgpPnQeLIrRqoCPnsqaS+c6vz6yjFDnMUUokBy8B
K73J4YrQmjnLTTE0AnRE2Jh0DGvZXvki5jD9TonZAYkZDlc0Wx2mTjmGXLL+IUPK
6x4Sjr1WWEIAkoO0yyfo7xfJIjoTrlrPqBc+l0oAcEa3LaYyIpDdEWn6AK+ABX4S
lB8Rt4fQrPjuAVEzcGIGf69slbdb2VWviPwLuXkEQfev2Yed4ziYUOQfvVyKM+Pu
y4YCda7Pmgugy/FQustxa6RgLpmfCbP6rSWxCRRv89NjpTrAptwTnVsJmizHztEI
DLGPBAp3bevqyzShCScbHbvTOWUg/qi3H8hbxwRjUKIgpN4lHmvYExdx+s0uCgjn
lMb8a7afXEIFzv9j4152pWhmKLwapj3W4VPhImmESvvdtA5OfybXh7/ucCYq54Vd
Dc85iYYfdOxhiAVdrO2SPAdDxSlnmXo9TH7BtbN5G7tHoXIU7mWh2hO1i3dRMneY
yW5sHzKcdbvy9GNFscWzd0kfKAGDjLYVRALDZssjBGXumGQ2zrju0O6Hwb2ery59
YhcCm9VzNvEM49lw9sqSj867tMWbA2MhztfwvbY3+FgVOxz/gGMPHZCa8t17T7U5
iFi+Vpp7JLABXMrW5S0aXWLBDrC/sNenXWCxBSV9q94D0igj2/Us0xxGdEfzF5cH
N4niSGkzqcH+Dzc05ZA5hvL6mQOFIEWf653y8AKMwpbAVqCAQwAXxlLS7inK8R5p
ScTOHvWXGQQszspMG7JEGmsR7MgUqPnROFZUBlhmU/rrKUwFMDWm1N4JMl86GWpB
16OEVNlaXxp1CPm8jhOgFBbYLOF2OAhITI4u257GRioOk4/HYDHhV3Gip2qrIFdO
HwhhO5oj+T+TpyM6a8CZF3Rf3pN/6WGEyYOJ6ttXsJ/FEvy+fwKT/2S09Z6DmoIx
y/EfkJBSTHmeHafL4CiEGN0mYA+UYCwPgmLMXj1OeGWO8qBEr3kkKoVualRN2RNP
f+UI2n1FBdiT0MDaEWl23dcooieKxz2u8b4CGV727NYGFohmwb+jIM4tyqh4pprV
joJddbzKESFoV9ZU2KZBHcCg4f3p6XZ9blhs3FGvc3To3KcH3FfE4j1WMvG1Puis
o6gO13dNsbnc/vhV3OJ4/lGYJQnp4cVDIJorWoYMBYfEcijBHjSiqWnP7vyPw0Gl
qGBPbb3SvhzF+zM2AUThZCdApYVkblffDOMyl8/lEhZkuvZ6j9bmpXJZ8ZTxg4a/
Y6CGJ4Gx0xejfFq0X1m/f1OsuQUMP6OWKaCfcq772e8qr1WL6l1IHM/yPh/wVpai
8mXv3u9uw0doJj9e4zYuzmCyxphk+1cXL882C15PqsAIZaIapfzlldekh+7N8eG+
lCqvHQf+g2s3Jcp1RNi88vOVQcOLcMJ2PkpOR6ZZi4EDfEkNqyUcz/C8n7jApkF4
mKmTDf6IAPMI9txR+V8Zz6IdSQYNj0u+vS0QrjT6z9Kl4PpZkNiBE4mljYdtU5Mf
hoDGAQALDD8+LAax+tkvxc3pIBJRAbgXfO4fRid7dz3YuZMhtDCyJyx6Vgb6g2fS
aVAZpn/xwWSNlZe5wI1JuyWQV5kAecNNakLkO3WDx8I1YOzuwHY0u/Y7cedYtTL8
2MrlKcMZsaUaU/iHHrNvntw09OFWn8d9QFV31txPjFx8mLKv5YjwH1KM/sqH+i9Y
BLts0xYE37QysnN0Z0bzDKqylwrxKN4MEZD1UXXoqUSjxvELOy+gTem2R8WP73fM
yaiOswHjDVS4hs8kj0CZo/HDveeY/w/JDGbGIUnQeDqb0WTwRDuRn3SXC8vwGhim
hyl+hbHtDFTPCl9B+pRpSTLf0xp5mq/CboLvO4ul0kRjebe25OVvw1qtgia1q2Mg
5yGsnmy6zcoL5PS5O2VBKRNJcBlV2qqrFIXFt9tsXgHfmRn+ijY022tgc2PrD+3T
OckT7p2G2mFVgDxva/bu15tSXs3ApxJQye9CianbaNL9liuccR20puWtuouxRdOE
+iuYKFiaslsLe733Ni0+vvZpTqDE8l0NXMib8lRcrAAyKXjJl8BEWP0vJjuI484/
trStUhf2twf4I82zAlLQu9pBoTpiVVrBseGrj+easijQnacydBg++DybZH4fNTye
il0h/ZXhgPnYt6VzlLkmIxY3s0ZhfcYqxi7YHyxW0KFwYwHKt+umKNmx1rFvcILn
QZ6bnedo01s4+SbG8+DiVJjq8xNspXawXR81w/o4oQTK3FLzlSEPY1x1bw/6aLXJ
Cd2PTMM0BRgTiCVRj3sudKMKzE1hpgiC1fCSQGj8fPpzh/cH0wU1+ZEuAwYmcxNa
wLGKoWaptPdjEp2ZO1Lfzzrp/pfhdwQQn1bh2QpnPvUo7E2Kl9iO9Qq7cgQstswQ
5+SZyotoRaN+B0bFRZoNv2otvKDe0ZAHiXtTK8IAcdUONIFTELFbuNL68D9zBQmE
2RwJAU2/xX73rPiaSlQfC68zDWQg0znpPAt+gh484SAmnj7+Ke99J1UxYQ+HRrW+
g3M9ihelto32bL4wQdykI3iZ2A9YK9/VcrUAFQfM8pjbWJp2Ztjw8E0eP6JqibMB
5/nSKhuiYlrDTBHkPQbaUmFrhS2fZbR3bUPldGvSz8L58FXE6TQG5QyN8R5go5Ep
kg6JBdLK7bUru/kKvlJt8Xnh6J0YWidqt0nqCiVb0hl7EOXbULXc3/TY++s34RVu
zYdCOlXmDbsSuihIGVriYWLsZ7esRPoe/B6MslE9u/sPGfOiZF0EgLRx8cZKQOq5
mKNqIKZ5PoXWrGUfPPFjmvYqT9bfSd02tBbthPUnzh3rwwnBwXaiBey8o85Ml0Ci
g7qwKV9lBMPw4WxFy/23ETZJjVV6Hd5NmA9MLGcf56+W8ObRTGn39j5/+H363t2o
oca7M/SZsia6+4QQB2eAHjpDRaoeNSNJ1SpmE5EkK0Wz0/41sUE0MN30gYiNW32m
BihgrhSyZ54hF2A176XurPh+i7ovj5aQ/ADVft7cYgSuUsXXjLmGzu9Zp7l8htLU
Z0c+ZKJwv8rvAAH1Dvm+f7/0W+Y5WTzHBw35tQZJhT4ZTEG0tbKelYvnXoW6BDxR
0m3xEst9t5axlMkwW2lICEq9ip+xmyremtzEL23ykwr3ngVqnioyYceJ32eFRzgx
2A0Gt/HXaF7NcKosTq5DwGK6nJ0YDT7Nnx7ajlKuy7dVTPhNqsQ2/aXrlwLUx+CT
9P9uaWhuKQpaIBaPcPsEn+2hiVZUlkURRRI1tqliX6xQ2Mwe1Xga54CeMMfoSLs0
bS1jM4Bm1aR5dAG19qoyYCcwyKWZJsBd95w/jn/ovgy/pB80aQRGBsT7JsisR8lx
H5n7gKBbMEDbC3sKapBbzFL1ubD4pigGz1Xg8vyKnOApSqlz9xlDzKOCrchCTwnC
pe/dfKANWk58iUC2NIPpPdQ1eCt+5/lnfO8/XYafYzkJnsJ9n2Cj6IuBo2pB73ud
GYRdRQLSGsZnDSY6aHQF+rDaASU9NG3rtM6Q+hGouv8ltLCEUqUCeQLRurrFy4mj
KeSHnpAoIES+Gk5Gwp/YcMltn+JI+PkW1FIzsUpFWf32NXfCrwlaJi076z//1zqB
nWOAM2MVHI3MABs5Uw/9mXzVWNbgLYedbBQh6nWM+GveDyDbYmqsUzd4ovRdyFaZ
ZYwPiAoJq63iTNokjiaVkqlI11gN8CzxSqQGAl6+EMkTOx1GgF84PBBz1DNeuVIL
xhyCNva5QSmpQr3ITxDdFoaAl4/PaRwF8dY0jeqdHSlnU7FkOFukePlHtnO35qRd
/biE/05eTXZZu4bgK9LGzvNzCQYi0b3bFgeWrIT73SSFWGZqe9f8vYa2dCC5IazZ
x79EXPo8qLNzH4e/YPuNOOjfQec7jqEjJQWOLyzAcsXMzoyG7i1K0L1iQI2DcjNt
Ru1PAvBXHM5hUeDn1zbf52oP3FQ2QYAT93zENDHFTh0FHw//Yhwt9ECmdk79C9Qo
oZru1G7SG++d+Q3msZwoxDSe0PbY1FjAWqT8qGQAdXDmalMYQUSoaoSu6wnnpzyT
JswkBk5yBjhtj/U3z3fYo4gu1Zn2dn9ziU00nqc9T8gLOAS3UjX43litDSyasSGD
+T3kq4KiTwETlnOLLl3IvwdhXg9lMNiVo68WU+MPvKZyy8INW4xCYXaj+CFuRMuz
aL0S53mTcXK/uujB/1fpQYW6jDTkFkMkLrFq1amNFI5hAR93m/bj3Q1ENMICKhs3
TKe4uCHsnjXAB5tQDq04PuJWOr7qtM6d2nEMDVCkB4dCnj4g+3oc/yJXhyEWvxEP
xYPpnY1529j79UHhgG+P34BCRIFF6CpH5IS8IaW8jCRDJMrOGNUEzFtfP5aAOvIb
4EnSPHvkTWSdP+fB9AnG3LBlHV8OlAJUUSVlQfKPymsFz4JM3gv5+3g1Xft4PyGL
bJeSuOeuTyvlIYyUzrewhJC5qoz0ioiZCdBarmkdXwajC9AugCurnRDLM3pHlgbw
eWLztmJ3wsWyr8nvoqFG4I7eAlyEyXFKrYbCL4DW4mTcJFXOCMbo5hXcT59bdQe4
kTf+oDoKyZYBAVn3VOBTZwlnkVXt3xsqn0JYltmulyquXiPm1uZ6ojZ5CFxHxksz
APSYEWmHGhFoATbuFbC1n+S2Go1AN/CYLfG3BOj2L/yRiI3Fv8pP37DEgBdk4NnI
m3knFXalzY+h9Yt9N9BZIVGL5t9RjqP0DQM5E+ILKjfKCg6Nz6U/8DIatpsnWRs+
YqTVuQUR6huVwlP4sLWJsTu4wkqj7xPrdErZquRCeaeoM8MTY5IEwLFu0vjGw3DP
+ojBFH3Q0dSbwaM6Ltj3pcOwbKwaLbFnUlKfTVg9xR4eshyvgHAgJ7HNbKvKbe3k
jXeWv4+Ebpj7Xv6Zu9Ysg9dZD3mNVnRcgZ//BJK8md1FI+/vfz0NmIeiNmF6LYL9
z0E5gH3/OUlCeRNi0xgf+mRpvcQ8CS25Oj92NgQULfAMeWKlDGpUplDaHCBh1SNC
6BB3KeW8umwawa+LZk0RHDDqUtWsXTxHV0UB5UYXylGAc3o7PnqlGFgUUj5vGIRJ
tS7VWaWpZ4nug8be4V8u7dktNmukj38itcu3zWNSkVRZM7WYgovv9We0/jCNaqQ9
wDpyZppex5ntGUto5+OybLRXofplLEub8Dbj7LwmAk+H09G8cmo6jSoiic50oJfK
yLZrpxUUof7h3f6Ms97uxuzEhBIE9z5kd5e5kxfMlfH5VmDh3nJ2GQCJjNCyB7un
kyLDh7AjWyeyCXN2plSJi9Dvtv1zM7SRRijckqG/4N9bkMICCbFQ8kg2XjfR35gp
hguR3nWYdX8xN4FKrs5Pj102aAZTdZkiRwPy2PtbjOwgQfN76e5gNwkc+X1VapX5
XEG9aurMeHdS4fIXJjflLwjBx3JmAZl4QQ0mQNjhydZAyfpvKTUm8bc3WK/zzBdF
/QUY1YQdTGbgevR5ba72vHnrO80wuEM7apUwfhyQN/FhoFYbp38xJ5EupaKEJ6r+
cDCNFZyj48ZdBvfnNAqpOHlEcXeRqg5zS6XhzGV3jAL2X2NxAbVZfZAp+ChwU1ay
ROgBiSoCIBSlxmFXIQpwylS50AzVKC66ssj5DcFhCTDAQ+4OVWOLJpZ19IYmzms/
sDQKSVyUhJwpk+cdkd+2GJPK/JU3t1UEPq2iDV7k///vCKNcfqueNz6rAtiA1gaO
ZfwrqD/US1pZiVz8gAOZoNAv3MVNEwwfiEUKu+hL2N8K4Z5JJayWIahzFeTvgGt8
O+xRZEmZnIk2MsU5Y2Pdz/J9Lg4QV586caYGDNi3V1OHIcTdMAjDVYpIjc4JbSh7
45VXj5CjdJP3n6Ja2iQXtmNj7suPYFQbGNWwu5F1zr6XFovL7IK7h99OQa/Aa3U7
MeHqsXUPaGcwOTCHU2PvddeKvLyC7BiynFCv6QNQWqD51MdtVvcF6Ib0E4QeFuLZ
Ajeu7jRyqqjPybUxufd0NuDp9FhafLNIQN3/4aG/0Ytt8aQRflJH7BCSNkxKMxOI
3hMlrWnW34bdVFPW3tcEhK9grryjdcdW19lcYTmSq3UjiMldGv8b2/V/4fBNSs3t
kSntEf3gsDM/5ZWLiHHLa5qHGVsC11UXcGPpBY/P4UgzdCHtCjIrb++XqUx8IGOv
eckQkm47fVhQ9bExLEsRFDYCfJRzHYCzenrPO1GokAX3aH3otXYJ06/ATLqtIAfs
5cnWEFaYoeykEWAZIqdoo1dcp29QrjFuQq2ocUYDFOtEsHUWE4dVlVbZxRB8uAC3
nquLYWERIop7mvH37um6yaSYuRdZEsyWOUDYR2nprmMY+Xp90E1XOSC42gyxxmY3
B0DGHOGSMg43dM5ICM1+00Wowm5bZnuyxh7rTahFNwhAf5aB12xOhSbn7r/ZmWQG
qPuxN4ar5j07GuDbLRf5uuDezQLANJTpGquDiAcs9rN8n4oX+zwGNmjEGReQjZ+A
PRc0uiveb3zkGx+9ZjdO6JsBejbhGT19Swp14EsUPEw8/1g+QA1HsDbFY9jmN3mP
1Ap4auL7Ek+fEPR9Dw3R+cTbsvDfqeB2sNJaRRLl/Cztj4sih5shUgDsGfjXhEAH
S8NWUCpQY5Bc/ozgkXecwhugjRQk72HLRqyXPcPpVchfpAiJOzZoXOIhoODSRi4x
tVq0zI0LIwGvUQePtJ1Yn96YqxqqPjxXXt9j6TcDGHxnVfjBXA102uAtrMkwiilj
l/+xLBK7ip1g1G2zlwzBVRrmQcoSuNbz0/1+Xot9MmaeGPxFYsCoTAoihTyWE5Li
Ha/5bsZ6/9c0lSbqQiwMo1WLfy3igrX8hUfjV8OA0bmgT7MwRAXva40qoc1lSU7g
A1mcJ3xT9hoxGqL9zcLIr/qdxk36jkRdX7qvFSZ1Fe71474qD6YwNPipJ0iDIcMD
g7gcKOIg2kfU+Le3wUeFUzWF/4/7c90DYrX4oDC3D0tuikYi1ea9oXkXLbLs10vZ
URJ8s6VSQQEvaNQCk8gHEf0OrHArmDe8w789u6AlqJ7B7fLcJP0UB1zVihVyqi0o
9DNp80R893dtOkk0bPxoMLU7jLAuMkVJ/kRv8M06nd09VthUnxZiIVAcoRAlJ19X
1lMGUsrYRWFVH37YW1S8gt2qCcYFZyj45ED+T98U9qCU8/AE/nbyh1VfNUwovBu/
Foux6NWuakQGdyYdMsol1I3VJO51pC82VB361JbUHF0CY/48vh3YSlRJjjGbKUuj
NKH8+wxu4xx5NF3g5/awgm6is6VdZXngHBuUfl7mLh/FiZSnbe1uljnjvb8L9wIb
lV4gQ1KfJ+UXRVHDKsjcrES0pCfkTt3cyh6nizIfL//6eEGYETI7wTcOu9QSXt7H
skP8bTM7sfyzRIdbeEl/wFhaIlnW/Jslz/hBKpTHBG9oQRH6uL8gwQCd9nWesgYH
ocSjOxl382vJxveYmY7eFH3oejN+nI436yCZnMeLZXqEbPjOKfwO3U0Zg2ePjubW
RYLOjwk33YabXOBqU4Bqx8jwnMeO8SSFsnCjr8gg1X9IRLTsbTGYV4NojLCsUdD4
Xj2UyWcC1Ba41VNgacNMsFW/unWCsuOcpBhhQCVmRudIB3KpLoA4eYpygzTA47FI
LhTv75t8DC9aLILX3cF+4gzWr3IXaCe/kIrlnPIGAqqJoN9GP8npRyCbZqjIZT2r
2X3kex4keYanuf3BUOSX+lV5GbtLG4uIQrSeiFkZEZ3QivccqpETTn/i9A8Nt5vn
LSSUaK6R/Cn8R0PvH+yEJqykpuckDoxYLQqdrfG2f6qKyMyPW8SO80nRd844QUyp
qxqYXrfruSPI36Rgz41KFILvtxKmAPitrkVKYf3E60oMuR57BjwgQYTvHGqtD4SU
fR7spIsCKlY98YR6NeT/M1u1TsBMsPo1MWx7/vf/jufJsQVfMeFLDwsekOtzpA8f
ZLKuCHo2P/6YrODVZSS+pG501zEJN0mtEsRNZNOMBKwsN6gL6blGIHvt694xmhJu
80EnxtQ+EHeKqmaJJdXHC2ahIpBkWA2wv9TjKgSlZFl+XSX4uBB7KDKMzvzCdq5l
BBEs6s1FzlMLbj8uc/ijrMtx7K3oDdNRvqi3Mzvphi+KAjWBQ/0U0rke/BgE/dwe
/IGOYZzmAwSSs5G2oNvclPG1ywxPgbUUbqIe2N82rPO3YfzVMpJyTuUHd7yhAfWp
yQIbx4UtoGI7mQOP8/eUxOSDJhi/zUrsy6orRWnDYVgR2ez3pl2bataHdl3bijf1
CLl5st84RHkNph2khbBvTL1KlbxmTKa6pT9Bav6two8br6DRkRllM2KRWX7P6osa
NOfdeFyetwBXzOYsK48lIhH0FQsxpuEeu0eo1DiNAjaseVD+KJ6FPrBkIiBwN0iH
dltiMt0dFzYTWH9G9DFvMFvmqO4DmIH+8HttenAC6+cbN8ntNyDTnPvSyi8PyjmY
DmpVjhQHGBbk8ublmEgUz9G5md8P/0zUbAfiqDszXyY7jKOlpzZdCSTGE9IFz1QV
nX+8RndaCLE28eRU/2rNLP9luB4bV1yuyIOQ5JHOaZW+oT2KObFmuI7aKZ5+8AIw
NKDf1953TObm5fjiolEXozJvQKSDIw2Ugai72mmbplQlH8b9FGHESfTEPry1QSzy
WfJxVuZJmjmtN8t5wRNulKcBK3Q5hlRrkjyNpS9S34KboHJH3HaYshhZYcsTNXSV
LMT2JxgcH6hH1yvAjYXn7vTUAk6PRdIG4LpCfc5+iqPB+xrvtCGHzOAKJAewV6q3
y8YoYZVfMWjb+3sb8+dN6q0pwjl3BfyD5/mNGRkxQp18vNDS8M1+WBAUgT3KYhwW
7XIBnB7xdfosPnfr/2aze1xaNXIP5BOMzyfXrwWvbPCG+R6s0zrLKMQoFtHGREQG
ZzrgBiBXTmICZZSaahr4+EGCUl8hjPI4IP/VbkgZQVDDzZBvJURdSy2zqf6nhZVZ
GFD+Cjlb2hMC3YuT4p1PF1hN+RAJ4STxBSQHCwFg8PwibqEH+h3/jFJv1aGlRqua
c3JyBRhKrRnLeKaqc2paflSDsqJm3GhEcbYuKY2D6RKojt8cNuSu01hM7dHnot6d
wUXPFigwiL7GQ5d8KagivKxx+ioJUrb0DogTmlm8Zt87PJZI9aExHITJLNam7O1p
QFvo1P4QynfVV/iPt1klUKx3+xmSFBhSmu9Bkwdsoku4MGUR36ahcuZTG3ElnbJz
r62F8eSr5e1h3G5fA9ggnNRCDZkWJoqZur7rkvZWEZ2SnALNvZu1SrYhv9+VZ88T
5VtrFY2zKIl2+4FEMxlVW+z7b+87ifNC41uo063rT0bqHF7QCHYBJb8uaVktK44z
Hq33J/NyybmQ+QY3bjqOLMHEOxih5bd1SlblKvh8WvmY6mO+KQwVYzWtX4ohDqwv
f97VbiHUFs0kO+KB4AJxhgxeLb78UV70GnOtD38+QBQ7tUS/CcT4QvnmdFx/nz7k
CNS09FdK/jRkq3CZYLNPxNzBGNDk+20mAiRMed8zgFIbWi9ovQX//9GMXdVyHbe6
v477RZ+ioZiTs44aNZCeHkeFv3lC7gUnZhmo/jlBUqKdu1BpQHx7QfK56CbQtFDk
6M4my5KfCoD1dHzvtTYSuOpGYUl/uEDP5qzxzQDIvKH0k0kScQggl7B/4L73UKSv
H8RsiI6tO80rtW0z8fcAGaZchYAheOxlfFLvCXwfZup2AGgcQkuSTXG4gd19P9NR
kcmCC1euNeuj324Zof7mRwAKrkvdY1nUQ3ktsSZ5z46sC4Q3ui9fdek8lNKQRaDa
6zqz1P266zS5NGzGpQEy0/SKNOX4U4I3/wICyCDxljGD79zRAymxW2SLtlbTBoKn
3+/IlgMy5XPqsV0/+96ospp1Ko3LtFNPuNo5JWUEQAlOpRxbI+4OV9cYaU9mAW7f
wQsGLwIykd+6LyHWuZ4cYOrokr+fDmJrBd9b87xOKOvGBkRj7ymYZPacZTI8NeGC
I3IX9d0euORHB4KPbmRu/EhIz4S73phufAHK8Ehyi4PrhhzhgJ6ugXiuHfDrX1Rz
ctfRUyHVCc2xadQA9NuSeGKPUTdp6at8z6ip1yEa7Rnn5Sx3BOrsN5NborxgDL7H
+eOyEY7Z4AgBPGBymmIYgdJZvQDfEWrLGgYHkdS7NvTT7nXxALF8D43IeeJ457Zv
n9n2lWo9PSfbfmtUm/57jHkueSeOni/NBQKtTlCiKvL/+R273VwfcfzrKXTFaUTi
dhlWrHyovJy/Z296aB7lyXA5aquGQJw8+8069SZgqP0a2eVRvdtg82aps4d5pbF7
XKfmnStuFqZ6zJ1qPulSKOo0uF9e2Dqumm3eRQ8VqVE5nD/5FWKmHZ8mmcVde0rp
9riW9fZy2o2R3ZfGdldUg0kfPw6LBd1aZ56t+OahAd9vBE09dteHvEyRgM/b8RM4
qyxX+P5C03Ewgvv5Cbq8fvNfS1wLvLUIO6ERjJ8QKqnCZvUaFfgOg6b8X8Zai22C
79DAhaatxIF1Yr8sRHHqORFUKvNDS1nRzdAQHZvyUYY9kDPi1iTaUTSNas1mhjn8
K/HIWeWO/0ELQRQ2+xtOIjXhQfatUluksgasuDxmFQzPSYK7qlCBq6uz2r2INi0P
pjjCKhR64h2NjXzajQGwsBvmpvb2htHZKpc/l0PU6frDrWv8kRPQEPcQ6jOth4JY
EO7MIdlCo4LblIWB+PuQMeywqkBpVnI1MdvhXSawnC1QZd6kC8PnMo3Yq97zti/0
m9TpEg7Dj6C0yeF7ZTHLgnBAi++kf6jEVCLhxACt1L6egh8C1ut2JYDXKMgnRTj5
GDGfPlh6dLA3ReSAitDxGo/vSXsZ+hJxeYSvns0ceWxkUahDbHbUDw94vX40spND
aYi+rMiMFoq3GJPNbbvVRqc6KJ7Bm7iul9qORytmf4bA3UEW+6rFdE8TKhY4Y4Gr
227vrMuHxdY+ta4JVw0MQaZa7XZ7hDySE1xc5EJoQ5BLNgi2WMiHWuQV76JBvNbN
N08EtAQOqXwbCyEA7q9NFkOopQy91sG2CyJoWXsj7Lr0oSI0pcZ1mvun121njW4m
NSiop+ozWlOpUAYI8V6nlex8p1BGHiXbN5urPfnNVyiey8JZ4NgrQRGA8xtu0JvV
NY+9RYi73spylSg3GUHGANLAQlEz2hUd52j8NNoYxqe4WJYrm4YG0XShrvbC7+gR
35kyEeSropC6HMpp3/MZg2fST18Op+UTgFPpOgCaJ2g+Q+8xyTs4/kzCzWeFxGHu
U+MJQgKaNyOMkDucqiDQzV/notX8f+eVIcoiYbpQbMRjsATBQSB7R8lvfLE8VbnD
6lh8TmQwCbIcOPDcRB4USoqPA4e+W/WbPvrElVl/3wmRUfXLrwvoB11xubnAIbmI
cwrMYFl2/omfNyPbS93ipHHBlEKs/AdGTu9jovR7+lBgiMBX9hMXyO+8/A0GNd7j
9q9p6CA3d7ixu0GxTH1qP9XZh5UAI4IHNSPrcVoetpPJqfpuMiXrzTLiz0JO9kBh
+7lawWZvFqMelnSFaOTCVawoLuttHwFP46kaVKd/RYnLkJHaqRBG8sx+GG1dXy4p
St2xSY5Xu5ruausaao5HgSusnzuBOpanfhTlEGzUUb+/HNviCtNDJYI1TNq+tNMa
HLjRYi1jRZxwhESkiVVlw6zsAETyeiQuc4FL5S++he0Q0fkgg7fBGl5I58eadYsI
E2QwpgXxN4MoSpjaylP2bDV8pWqraLdI3eZVERgK3DW6iT47qiguk4Q77ntGZdOm
EvqILmVUNa2iEpMiggGPndbssjsr+HoR36bC1OLofvDXtvluJOOU6wiY6O+A1+L4
F+FggXCZuf3cYhG0aURlSA48CBcodgM5eW+8tueh/Ma+1M3K/8+iORPSxtdveRmf
KpWtrUcugizvF0BSkNxX/Jp05bMsxC6n0doldNBPsQ0cd2NfEFhOJwJMRztPTAPu
5pvGkQ8iIjJtNrqhDZSj1VuWr0eUFMdLppPfkVLHTeASgeTqHRMm1oScX8DmwtZd
F6wHLpENy90nfJ8AsOSf5EYCxTm8Zj+wLyG7+Sj85Q9jm7uUrZYhK8Rfqntlg8Hm
Y7nQb2Gd43meSPCzLtzAhZ1V/OLjzLv/cSnjl3pSIiXd19awk9av/h51C7NMXQ0k
taJcnRYw0kaLsRPlS6Zh2tl97iNegp6Z0u+z15lFClOO31+WwtveQ/5rxEqnEXnc
kwgo/Suc5iQsvYtU3EuEdod1Zvw4y9GL8lAOhy6VToLj7fAT1qxMtkEDkd+EE+6A
J0GpBKnsXUw1AlpoapM097CXqjsAKODu54VyQacXIrJFCL/oaaHlRuXF4gR+Jr5O
tYK2KELWSr9NwezbIOx3cFNKhgNIpahxvkLRH/+AFN88sOa+nf9Z6LjdFLJU/O7T
l5lgbZp9PJGQFL+VLM/sWoH37zWHXqM2RpZJycr6HCnA4eElsUZAACoLy7Uqfdli
80h/VYYGTtGl9r62pKyElfMZLpnV2D9dVv+LZgknSqBMIjMXYEIpR/vlXlrD5A2D
Ksh7aEQmCTc3yIB/Os7RyssvEYMJ9SlC/ZJ2ComznkaOdp8xAXQd2JbSZwDBatJk
URth7QuAfXU5+JlD0Fy4UoCugfjEWiJwobnePzEWChEDLQAkAz98L+4HHKz2KnY2
TU8UBr8y29s8rC0SsG3XFYTCgefMu+Iapu6E+VjYF/wDkH8xEA15JpWYoZNiERNr
ioCDO7RhH1VF6aBH26IN60rCG6trVbceRBmGOTMEgMfSv7aJ+RQW4RwcWPL6Dvhk
wjvXkG66LLG53E7ySY+Ffd0dbMucHZjtfy1mvnyj8tX89yfk+xWPFsB/oakFkPVx
QZWafN7ePHoAiZe7rGttpKggGS1rJmoX3/jbwMs5QPqvVdDUUzClZgRtcs1cOhI3
HB21BEJPlU8ss/2zt1l2/SZn3pi3f1/6wTPWaJH3Mo0FHR9vx/Y7MQDXiD8JUTvG
gj2QYvhg9QkvTkfZlWY9nrVkCeArAfFzLxb3jcwYKhK831P8XBLcAN0KjcD4balr
ZQBzF2P2vyjVB2cO1kGtNMwKEgrAuTUPvsnrqXW5nIuTOBVYgO7+4JnAGgUmaPrG
mtrH1O8dr40b1/3uVcz9P8fdS+IC5nRuqzN14tlIAlb4/dWkivvT1GPMegGhS4f3
bpizhpRPh0duVt1xvtbCjMzEW91Cm2Y5l8Pnev7a4TUn3kY3IhRn9X1ee2ZI5+aI
4BzquF67X9XXvfFjwOQbk7X2F0rHy+0I0pVEGki5vSwuQ0OIkiXhsu2BJGAISPrB
AklkBOd6TDbQ883KcfgNNALNDrXLYBtYbE1VMWs0LM7819P8XbHdbEWCBInZnX1q
I2rZXRZAag9lmoS25+P5nza7SGEU5oUXcCUzlR9uc5KkpKdIJ5z955cCTVFX3L8v
9Ghts0gbcyQwr9eC5aMtHh6BWGpVuX4QC7q7syoD8/RXD+gs3O9HoHxf3BfX0biO
vdArPMaN88MQzGJ+ClbQCnyfmlWoZGLD6uVYvhff3BcMEazomvSpISVyGP0PrQjv
YW84Bs07gAL7OYbPuG2hpW4kNOdVdKxQxHBjKUvpA5o5AVGiP1qsIrNj0nzglSlq
I+haPxoZc87e15n1BXqwOY7wiYv4+Qr4GQM6qNEPk4l8YrhvyyE563mJty822Rzv
dV9WsBwwZQRGPSokqXqGxxYBWuOTirPs2C2dP6qJmCrtu+lDVzXMPVy8/gSOkSyJ
LGMyvXkGYgt8KNGS9S/ZVsvU19WWePxumxEaBgFaPWfqhgfGou/hLYN1KSPHKXNP
WiDCOtJcFNkM/JiRfXTboHhX3HUVNsOtr08i+o8iLbG5Epb/MK0X8fxvbHtDTIIL
TfuG1YzoEgpZnqLXSry5EKtMJqG5K33wSfs6Izeah7GpyF5aWfYPJfqOG8SrVYde
CEYJFC8SizVWVHT7jhmsO1GbSAX8dK2AFYZ/jb7N7Q3vtqDGCCrYJGokPdkd37mY
EL6Trmlmv2JcEuajauczl7CNJXZLLzMg3fr7ONQNmwysPt/LPrUobVgAItxeKdxH
K7Ucuj4Da06qXqYGjQUcMpIFyZJ7UnJPxkIBg68YZUXZ5UfwMB3pBpRKvgNvrJKb
u5Rgs9ybg4dYUpjlbeeXKI0z+fuM3cOv16FdLfgmvUaEw9eS33OcmZ7Aw8R5mDZ0
pfDuFUD1aSZcydiy1hpxSDLHjs0+XAyj2fjanYMPDbwXNW2aAEsMnD70q/AE8oIT
mjtkYVJp7HteJ00g+C+cs7U6FhKcbM1iGx7YPyweJl6RwwWLMoD9PR6DIpocA8Sh
xmSwxPgMBTZDF15/MPVQZpg4GjgAmGU+GRl32JXV0xUweYh/42ObBUMd+pqguIBY
DN6KdvgoPJ3YFNNtjH1tS11PTogLsTdtzadqo2sGy44zS5rq5W6RPtP6X/lSwl0W
q9FU9C2NrRg27xaS78sDlLkaBjmpCNcgmjWk0LcDALfdNUYAMbzRj+glh3Qjv/Y3
VYDyxzSLHbc0eesjUY0kjz9mSevp9RXuNhu8MEXOduHEl+vcsJMA9VutAyBWZcxo
YaCE2cEJS5Nz5VEi/MC+r5yQ3nvl20dPinafeC0q3vVnmj/m5xz4BJfyIqCswFZ2
8o7KI/+7iDy13IoZs23C320rh3x/UBQY2rrXVFGbOnn+rcu8YWcEDnpl9kOzMpDN
udc5cEOoApH7qFNZuskDnQ70rYopJZNGQ6pHzKcfuVYL8F9bvqArbKP19PU7pP9b
uNC17b4CxiVFqL5AG578AGHodNlmnHl9o7I9M5o9TkoxAfTsiOsUqxRo04C7HoYr
Hne6bqIJECyRcYfYTbeNtWOt97f/GmFFSHRqoONVjFTIIRYot+vqdOVBCSPhm2vf
DXsMRXhAWf8uu3aLlifWzRtNEILgXclIfDQipm5n0S6/PoMpR4UGIKI7tgwxVvyz
psERhORQokkSt+XeuJWcLTJl+dNlu+immJ4p6fztOL7Cgf1LkK4PW8czC21Ulwtk
u72pOD5HlTbBfunE3GtK+OoonuWxLKtEuM4g4RVEtHhThW9Ubf4tkOY2ev5ac31G
VFva0JtKYbAb2cuTOg7Nty/lXSEPf36xFryzsfEROKTaBb097YThbrm3ItY0l5ns
MX8p5vAuJtPTiUYFeLLTsS5gknbCWOzw7sRIcG3tJyzbthp4PHX9kx5kfnEsz2E9
Nmhc4hb3CZJAtJhPRlzPkjFmhZnEEvpUmZyzmMyKdnMhCNMhX7h8GZUR6/fxFA1m
rJHmOFQGtcldjkSpoo8ISl32/L1B5HFDXth0mkIPHObxGViIwOeHRrnTOMXmfzcK
lDbeU9jiX3zN2KJarJjf0PVNgHlAbR+/5GfHayjvfF1eHu+FWlKmwigE50BfcbGb
KlPaQEDJmBuyRvINXN0sRYxjKjGUrdpTgqCXD2nchvajKkSADPnnOY/7MY+PE2AA
2QDdv9OZPB7zV69HLADzAbBvPLtL4SHXSHQ2lE1cnb5HT6rFsQj/maGeHlb07ms4
MUC4t574c+RgmfWT0RIB3JYzuy2xl1uO8pHPLWcMYmdgvc2dj93uHOpd3aRUK54R
aSsQ60w5Fv4XlGPCv56CD/+PXwybcElmxOybqKP2ijeGQnfFKj0GUPS/+7U3D2wQ
V+tYg7Y1ACbCazDn12rcREdhCIEZzU7h0xaB1yPhGtHhY/bbCzwMONqgXI9ELUYQ
Mcx/nBMJh+FdR/tUFZFzQAfZacAwr/KStv6RPFr1Cy06tBqJ5UZf1Lg8WEHXWHTc
VgO/+N7iu8XfSmW2DhC+6TaYVTFLGvVI4nfaxOoIxS1CEpODudyKzUplgRa0Bqlv
Yt/EM5gt/hHCOGDOWQlg5aawYtfrxoyYLXLDPgEd/noVwnO6mZG90qBTfq2bZmPE
7+J+WFNhnCb1AMUpr0UP4+ZSacyaF9QYlzNqeP0umbc196Sp69AYyJmz0hanReqs
MWi8DThxHvOvXsjrjfqa7/K7lbwJQtUDdR3UY2uj5tYYPRHBJWjBsF3QYGbJvM3V
KySJwB7j7QrWOdJjFfdMa2gehDQdrJX4lfh2V4W1Hl8kw6NgshWkbn6gwupTc2Lk
dRLsGza1mDRz/psWgJrtBXibH5u7FUvLKOgddMwRNz2OtlyYolmE77ZOLK+Lqsk7
H6k9j0/PGk78XNlkdyodCzDEGmiiQOVVwAPMsHMNmC/8Sy04GIDpkCR0qVMUbZlA
nfiR4zQODTSAK26W+EdPFlGoZCcXUhpn1P/5hHZgU0lw+0mbAliUmDSPFvDVpPI8
1HUQjXgUSdrsXjwSiq5eL09p6J7KsjCyLuwkB3zaPseeRfgWcKTDDNp894hWZmI2
YCJbJN7T311FYMNjAbUA0IIf8mDtygYXpqYgn2r1TrYe38I+qGIZgP9FWqMu2JZ4
2gf1X1ycHoK2cZylBu+zrQHPn5FlpUnIz2Ewye4+Dm/grJ9w1dAA5MDNOiv0VFSo
cmhs3N6Nx97nrxdl72BsCdWcyaJ5m/EYaUGFPMF1pD/3M5U90MVxvsiGRogDOqMs
bjfL8oGdUfWIdG6IrGV65RnpH9x98p/Dscjpq26TqmBrXTIA01nSPj/0F6pFebw1
jBpV9Kx4GOW0e6MYChWZAZlJLex0baDrrBVIP80jketO3R1iD8xVeRBaox705UpE
rSuDULk/3yKnmmcVqCC9fDEgGIICjzYB7cmuw13HSAqselXzigIU3DeoSebI9PUS
mi2VlknRtdP9xXHUeIRHSW7FO/qzxObc9gzafmi5K4ThC2pt4OH1TNQ2XAmu9Snl
W0+0UMduTPvBJulBI6c+bkTNve+ObpVckqm+p7xg9WkjUIK7v37bn4+sbI/N3IZK
3FJcOcYPpfC2RKFgMZ+jxSTwUpSmo+lgVmD/n48SUPRbziHoTFyC63opU1v/gLiW
y73Oie4dTj0GgH9+10nftNRS2VKpY/7iqoUSi96IbA1l/HXx932oc3AbcFH7hsbR
b8PthYdAS2gO9x83oNiVWupTqXM1KmIbSs9/TYRWM40w4YrpFUSah6i++bcqpfoP
bSdaWUrlLbiVgEvDtf+Dx9yc9Y7c75f26MzfrrvULhdFvKFSx5o0OhNqfCX97ymd
G4gqJE8SO1qEV5WZNCDSraNu9H481s3jzTX7fcE3fgMBD047F4Qx3yR5izk3zXoD
WHyWiXJed4+j0dddM2xbEJzSRjtOmL4y7NgmL1BvpS6LYW6wh9dNKsVeFBZuOn6b
pJo6r7Q4H5Syx9o/DX5hh3V7aodKvdCZnp5/6zcKpaghw0TK35WgvHZbqn79+4zQ
r4YsynEO/BOEiqdw8nomzhLgA1/43ff4ntR/fIIeU4eRPuxu6S+u+hSz7SoV9HxL
h5WvqUXRITL43IrjR2kJbo/IlBGlmulK65D7TzjJLBLepIHkhTpGXuu57SCfmhlh
esePUgNaY/MflpBFTex+sIz2fpesxeOFMqjrf6s/CAkBLNTkiPniPmRnF1bBgbhZ
r32R6aFDQiFQo4MIL/Bd73RA1VJEayg5kWX3lZsHsJjvRPPxfeAgsRG+TCFMqiki
Sr5tX/43JiOfZfBf0TwGhflUZKBv4Y1oVXviQ2ktWjzkwHfgo5/M053AVtJMEOuF
Trbl/d+6343y1SfPH6Wh/nNNgOjZzvIeHEmtrk0pDDkUzIRpMNmdt8fsFu9xX5v3
CM2p7j9A9FZU34/i7X4EV/G46ccT+34m4Pfrt5HFwB+Fb1TgjNM4GQblS62VoCrZ
OUXGT2rkGycbzrcbFgrXESj8YmyjVAV2Im4k4xhINQn+fz+wxdMTDzzRGqCtc/yl
TdcLN/EEedT5zkAxAGMiCtJ8HmLBCxGmKXLZiYp++/cMrBQ2MGOPfc9ReQGfdxLz
ESm7jBDQarjyTbjzQ6Y2VoVn74ttdKKNsL1XjitP93GvoWC9PYgc/LTAyc6UfnqP
TBuZ9zoouswooqryb73NwBhiNziU4v2I29IvEDMjHQTn78ElHAA9cnWiU3gY1oeB
MKswL4atG1Ob53BvRiXyS56jK/OfdfbJoGRuMQWcpdnp6M/2nHRQqGLzyBwFD0xj
eYu+QZHdsRhGC5Kj5Bqf0PzqcZqhqmc50h2jNFGNN7NHMSBmt0l86/0puJLWREZ3
8pzgmVg5VqH+4iXWCLiNeZMd4KUFqP97J0haQsU3dTMpvrmBxTqNKRGjfx+ozIgy
RgWKcTvkaZHjbbsBlBIJeSkAhGnJbSWgUPE2MEu/ohHSwJnkTynSLu1/lGa5bJo5
9qQyyVEmYBbzbWsbszI2JuMrnTI+0xCgfwjEhat9D0IALR0ISwoQpfLBEe1VvYoh
UwlTkkIDJ/95b00+AfIglVSgNumDP4sZL8f7yCOrB2M3F8mtXdzGou4BPd1eb3go
1B+5mMFTFZ+PUSoI7C15vbnLJFj/TmGwk1GkrmIfu1B3rmMU6zKvodDWyuQnMZhX
5bxnYOCgqenE3nqN2zD9AEcoJQ0AYSqARvQPHpYsj3ZsmJ7AFmiQa/nnmk+GyT8N
Lk7F7NVeY0QwQKqiBs+yM9WevEdowhVMrSxeDG7BzJuOYTAphCY7mR9/U2ASKXhx
nCxuBJUx3txdviwunQ0QIz/w8yrVnQtK6IhmB6zpE+v1zKIstGtr2uw/CLRe9cjY
ECoTDqizYMSN8Aow3aLvgCxTm6n4etlyhAHG4K56XSG588Zh/f2bVLBtXkzF0XuK
J1fPLSWYbJ/dhiokrS+DVPJcvaAC3orhomYnsE/ZA1IJPtUsIfpB3kk6ysClJ4FI
w8u0f/Z/aKi6xd59c+otXGF2xU0A514mW3ytTcfR8AetpUUzxHQFR2qYHHKOgEGY
DJfaQQYvSCKduaa/ACQHmy59TOwfm+U2M5o0aCKyP1CxAB9BKeVn5comQGNaEICY
vLCZpvbQHiLtBtZyDwg2wzTzG3JE7HnABX5eSGElJk9CPOw47WRlCeRW49CI3QIG
7rLXUPsBSdSarK4yNbAEQa8i8oaPc/NiL9yHsaEUBNDNVCHyKbbJGa0fdiUj2cG4
pVcAW2YHSRTEGrlSBAr9JqSfIcCdbBlaW7raz4iCUiOPUSdE6fiyerktuZbfWXqj
O70wdzho/QyP1CgS1AGN+al4wX0wM5+E9j0fWdKsXhHze4gIcMyinXXYMbSKX9L5
cNA4QQaEnrOHpTomKihN0+JTvJTvdxITzhp9YSHSWSHXG5FSDlNqNmqqZEtkfbIh
5JW8UWEbaWniw4AKyVosGs+7xep42VN8WrFwHjIZG9iyNDQfgm4xEknN38vCrHGs
/Cr4HAChHJmkGpv7DV3+aorzOqnQ53BJAK9XJ+QUyK0lBoF8Gv0EmNZvk/887Hzt
4bZZpqmfu/+gij+b7QvMIRkoxxkB+LY/M+nvhr2wqR/iAHvWF1v19tpCv7yo/PTg
sYM2WAcn1IVcmx/zHjoPUJvHRZwtpD07hVEiW2WC6U05l099XW68/pY025RXh+GV
4V//k41Iom38K3+RtenMFeYu3QTY2YgrZ0nmrrb7zdoxHFYnb4/RMec0W7t3L9qt
P4UHsKCLjTOAdnaIRVa+LNh0VOEHLsryk3rzxETbSLs02oTewF4cX7yVG5j7fa/K
eInnhAl0Ve3rPMWHpj0XfgS18a+9MOp54gIvLH5VdMQhE/sVqDwHMgIk/aevpJ/T
bvFqEMFO23N4UBG4XK2sVeW1fZoNSeOrcF7HKm+ENlWyMRYxWMJrTMkz0dP11eKp
BFFDlZ2jTxh3Mz8CYKuvUTW3UB3+Y9nM1uzcOBdaAUlf+jEs+n71ynYf5QfSROGW
KUUUl2kWMO9LYzgTTIxkaRQpK5G2V/6syfcpsT3JXBOqxFZ5AjTAef7mPTVb1jLZ
VIyNcmLxfkhJ3jqzJq9Op+DRXF29M1UZ2QwO3qNek22XU3W91+dDdbtGk4WdNNgS
MViesNUsJNYokAjmJFK2sq86RdAJWQckX0SXEPqLuAUihWiZ7wjb46lxpJXc+C/6
7fqkJlFp0WRuCn6M3jWNEZ5HvSKVtmQNlfvfJFXuNvxd/CBV66YZdGCMUTk29tSn
QwZNJyqkQpZ6jdlV7L4oiT0ZGomW15Xl8hUr4dvt7+ET8W7E/UjeNmKbicgwumIa
ff/kDqrSS0ZI6s6hoccw686TKNSyFg634pseMwU+cBD59Gb9Ny6BrcOEh1kMoxTu
LB0gLF/gRoeQEC/vCwQT7TsiCEJmfgNC+slhdR2vwfiydUDLl8xK2Y9JvP14a0WD
80aRy7ftq8XXx4f7TKiofoNPYh/W2c1+5H0VySPwBY7kkoTtE6mb6cB3QbwRG01k
4m95bNjnQLfz4qxkQBeYNQtmjMYdqmqtK1hHxMNiOj6KggBsCqfIrWd0oc2TmkCW
JTVyU65meK7SOTMD3Bhq6ct+ObfuU7dUecS44o/huWC502LIa+6oaf+PsIMGfHrR
C3NIKkLJkt3O869DvW6h9WUv6KJUwlZu7cWcPgN1swrAScd2nqjZL8uTYXkWfTYY
23AtYYYc2XFdANTltl9r1Wc5ATjgYDkcpaQhQHt1wZXpcsYZIVcEqAwJgQbhmlSJ
XNgBbnECGqiDQdPZpAycp/6ejwcd881e8QVMgyqngbVd84s9EKfdi3gyjTVYDpS1
tCp0Ssle+sqO9esLuGoePdaPrILtUSsTMS+jRvVi1CyZkWpfxtrB0xalbkzXwjVO
C1eVzf1XoQhjiKPf53LXblz5TO3ZDFGpR9j3oLpbWz/BveuQKHj9Lw+H1i61Oi1Z
G1toceHgMRAjIy6fscQVzC3EEho9c0J1VvxcZNkGjA7oQyGIfnbtJ2lNg+dGX1FU
sXQ81YefZfZALZ5FqG0Ljz+pma9kNFOcpZZ/RAKcki+aCMvX6IZbE5SBnswQU//5
ox+qF9fTNPyAexK3MKVi3pfww2KAgbmqRYSDkgmkZSG6Vemmr4a+aHSG80lzkOAC
oxaCm4u1g/a1isUguVHKwHPdazzs1cMaXEEA0jNpoEPgZhMUm1yMLk01hjrtQt58
eKvjpEmDg3L+cT/8jdRYCCQIuaMRLIFm+Xisw99dFCRC7HvmOaY3N3lWm59cSzAy
xwi9Ylgk7hWcYjtwTGB+7FwFYYsRUvDiSgI/zDUtvRT60WUgTyhlJ/6RFuD2lY3K
xcWpskNZrMdqIalYEd8G5/qiyIJAUJU512Wf0mNJuuHsW+Bu4Be/PxRC6460d487
EDDDMdAsayy8qXgYHfRvWJ3JHUna0B4AOIfVHy9U5PI0ycayTuJcjPbkwN7H3Cqf
cRRwk1Fbl3dLDmSq/V5pOg+0NGXCf3RFA/pgryRb3Gmzy1TC7prRHCn8/28B7JBD
XrZg5hQz22XVNHM9hL311jGVT/xhdLJ1r5k0nlFwlfc8thhMEmvTUPYy2ETWV87Z
Bi1FTVMiEJWNSW/juJs3d0U/iq8H/x947yZCSPCLqTJEIcPWGylm/ekWsskdMeHe
6F2QbmcK26l3ig2gTpYISw58pZ8o0yF5KhBWILtXjPuFwjMg3+KZNXw4AziIhKjq
nm74XFRBi6MY7+38t6zym0EoEiBtzOsMTt7AMHgOKQXv3bc8d9JCx6WfxZPLq7n0
uEAeOJHnzbDNaEvHQGb3JZ8Yy6vqPKNOEhl7FM34QfrPkMxgMgo7kewEkckwdCn8
99KMtJyBBvwTVo0gomYlx7G2vClloJHCnDHW1IybOQbE8NBEhl091XcFaETS8Qma
pJr6O5sbD3xHR1Ek6ky/lxyB1dL0yM9pB+zUBM7jfWv8tBQa2xSFIw7VYq8yMsJa
1PK6JCj4e+PNKgIRMcmyM6mWkeo4w0kTIEc214suKNSNFPbaWbYaVPfaWysIhVl0
Iw2whJSGYSRxN+RfClXRgyLvwoTYfA0mdo9y3Brm+QIKVwM1OnCi1lUAV79YppCR
u5Gw5W5wYy41vJiie1X2A01Cf1BwDPFzfFP7itNudB5Gw3Oe+U9zl4yAniMy9nuw
Fac4qnZGLD50xrdw2M5wKox71Gv4LrmOFPDxbQ4Pbe29u8+sZ+aPRnlD7T1F78/j
rx5Hr/+KY0nKnhDtP+c1lunKdmAdUNecn3PYXUQX4dkaQDW+4e2T1m1XoZGMFGj5
fzSrR+LuFbgAnTow+iziQsIN3XjB5eZM/SSf39Wi8rZN4poUkRPJgzXC97ANga6F
Tx8hYl/3mYt4NSdi/jjeeJ5VexBTc1MxhGavLd76Lic0dz0dELH/a96AfDF3trsq
6Mv1rA/wq27irGqIwy2VHEFzRzv7wYWcVLhE34DL3jPK1/UAepHJ6f5mfDM849D/
/f5Q4JF2alMosZ6Se6+aMbp0pZroCFV+j/Evvm3rgZ3YQy3nElUgaqC283+Fzv9k
g/WJTbd8mPSyKX54UdBjbCaTtcCrX5QFwog4UeSmQKrNbErexl2mvxenNV1jvhCi
a8BD1gCzVdrS6d+zYVmb1Z2fv45V10X5f51HuhiRRRKgd5n0jos/wqWS5g5pd3lx
hugAs1CEvps8WURPcCMGGS0k6OwDT8SKflCpTOt5CeI6XjrB6v+Au5mm58FRMb/y
+CjYG8o8tsO7hE5CGonpproi+RspI+SlUld3ExH97F/fK2naH333GTrmlTEMelmf
NfZe6JYfpBloVf2FLbR0SaZMfC+Axlinw3rNHoGuMBilzAaxDd6uWjpxaxK6TQ4V
/gvlsM0KdjiQmk5BWd6qMdYC0K7kPMMDnWvjpymSiUxMBz+8akZW3vjQ6cFanzcm
I81NpoPTg5gTcNqb4atlsExv0IyxZeScfud2xCqDKAADbg3zhbzpoy7+ondtwyPt
h5dZM/QQAf+8h4Jc952ABQ7wNpqMc5FLYgMgDj2TH9UQ63B9n2EAoZ/C6YtTLNiY
GipC79EmhLvUzlG7HEfqe/0aF7tAp55VPCHSnWAQ2bE09h1jQNNTpKNsEJ9SCI5Q
SXmjCk5BuC8EGxpJKiBhNwM+cBByiGFhC6Wy4RZGa4zVaU5ydORCF+K9onpj51TE
npgnVqu959kWOT7N6cDvy5RbXdoT82wl/dguxsieBSt64iGn4qjpH3FNGhmdaCIU
GeRQ3GAGTuKzPh95HKLAT6NUs2y4N20DbiYl56tx1KombEJcKKOMYaMptHIzehQb
+OZNSRRrjefs9w+cxgjnKt7wvHLFpcvvqFsGjGR+3X4rVFo1w2fLOqB/gh+IWw6d
vh8/JmRkZQn5UMHjqt6QuP6NjT1rOgSMajjO+SfmHSiMxHOW0lsFGSJf0cZzNb3Z
TBetWcgh8QAvf1RtWafluB30tNvTBaCdga+jEQ9vSonSunolgdNSXrHOPD9TFNnM
yf1wKlX78p3ZOLC0bGJVZL3PMxWSKLZdmmmRjKfvG7L+yUBDb3xB4apyIzb+Xcog
MzSXoF9JJ6EY1BLHf2pBFQ+K48PQCwuGZBTUahlNu/XefUs31zVNfBV9eARb1iQs
S+APyun//nnKFR7SGDzRmzfkgKzd3BcyRuI0bnwhh1tapMV/L7TzkaZNOstisEFv
XvDdb9ZsSzTL4l//ClAtEgW11cnOZ8eHPNGF2/6sT9psRgplOMd32igTIJQUOOSv
ow/ZVtmqOUP8mvSf3OJjIrT6aWaABUAJwfvg0KgrLwXR17DM4Mw2ZRmIjrwQR1nt
38BHZNY6mcYa4A00mHOgtpfm2nyvSeTSsMV5Nga9pLKwRI4+JlvpZKRjb3CZxrVi
ifbuAsWYqCVRYk9O5Tgwvc0qW/AECzKdyzgzrlL8S4p2MfJNM/ltIbejC1ayp0aN
zAhTRaFTz5cNPafnzGTzIShFlY5/fJScZrsnkodRMomrFtq2Rg74M9AJXtlyyLMZ
WvoGwu5RfTfM1/PEWpnnj5cDqlgyvi9PAfm5G9aUpk//QYxpbOqUn7pmdU4qyTWL
1wiR5dRlJ4cit3pg83jc62rSWXv2MAGPe8B2aMN4JJTOEqBrXnyQz4aDWMtUZrU1
TAcmuWZQpg1taIcKY7QKxLJpD+uhHqNynlQBIdCThX2XalC5MBA2NdPkN1d28uBL
NsMj2yxn0tDYhNK+DRmM510iKqIfYkWo2WPkFS+/7Fq20MGAZHH3SDcTw5r3WmUK
WCzVWgVE81ejj0GY1JiCzL0ZhzsmGTO0NnDeshDtRs3v1+pY+xK5sJq6Yeoq7zBr
qSbPf8B03zOdrFQei/cLQJuVFdW11M9LMmECB90XnZS9XN7CB3pyfL5x030xeLO0
NmomUBevosaUUzaTz+qeRUbpKW+6JSDvOqqw6HVQZpmcVIAIpytvIiaX4easWT3d
eWKfjf4cFPARyodasu8fJXWFsAh/HtLFtauaSFUtEstGSco72ec0+15R0h50Qf3h
BNRwHt/c64svWH2IidjvKajQ7HuaUyriOEX7x5pwBLwToo8rDZso4vx2qf2025y5
Ni0H4Q17LBxhwrcFvV7AtfxZRm2M4HHqWQwPethnQL4qMsXrVq+jvvEgz4CpFd/E
m45IWBpuzyDQlrjBxaAnra+Rk9S3PQdeiugEAFSUKR6zR8luo5ofnMABMxzOU6do
XrJXrRuFCM5ZTsTVONsbfV7zXlgWZfmmlb2c9pfxHf+B+PMmqR4BNzJU4fM6CsSy
tUbs1nuZ2Q7aZFbQQn7I61YUYIB/h/gB95DFaTt7V1iBPUAO4RHzh3WuAoU+v5xV
JmZQqQIebgd9WgkKYrKi53tBgp9MZiLLW34JnB2A3QjuUVV4v0gq0bXCfozkuTKk
LKegn6Z+eqkdQWy9H8DzWipdJI6+veeVtlOrM3C/7Hr/qSv3niElcOPajj9Gx5IM
wm7qGGuLSt1owehQbHVTD9st8BkR6wVpvuTgASKdwv0I8suvg/9mha+SZKaM4yJz
LKIZjRZx1eRHrhX9zwUfcuQoj3B6suBwPHUVRKZYR9qA6SHwo2GR+oofq/WY83xS
lpc5UruWqUU1dYA2cEesdknewNkv/BlIQuAj5sLyWZWjG0HSC4pJuu6adWwVXKQI
uHwnUq2bNa+5rsrPWqlyNQETWXFIypsKl3Jh+GY4Rn55pGU9LfUvemxSqLD+xW32
aR6KgjuAL32dsltPlv8XmaLLnsPXvluGTXcxeDZt29eFpuB6ROHyHDbwmt5j4i/p
MVj7lzBBxwlwIB82rv2j6doCRICawlfhX8y9xrXEb9+4OBiSBKlgEPFYTxMJnNbo
F0sT69NS2R46ksgbnwMht2k7N9Ism0G+CA2cJxRC+jkVawagXqkpdENQwzn/EOTV
ZSg9YKBhcxLS/CvOInZDHnPNropahoQVFLZM78vpzlYYDxSTNs2jbVkKBJTxIi9M
MDno77We/+1WkoiFmAKjjLSDVBM1oIv8S4g6X51bf/mjEc3i80ySp4/AlFhVUr4p
SfeBGiy74bWDeg/I9R6SXw1G9nOaZlvssTp/XQ5x7RpUi3k5U/X3vwEm5B53Vja4
GHz24zCY1zqHPsvspQytG2uROlzDdK//FMecHSo4P/y4dRE96u+TdAqYGl8sX+IY
KYNUiJSx5VSS+Dny/Rj62vUduwZFHNQskLC37oAHYXnmCpVocFdTLHywYc+rpxTv
i1FUVT/tIJFZZWVOksLPvCC8BpNYtR9Gd1mI2PenJXEHC65ez2O3a38H7kAWClqV
5Bp//u6rtQijul9ok6PnBD53v0IxuEjRXa34jR7NGkU2AiqcNHjDtQUBzh8C59IQ
48VVXUbIhFx7expZhzPutr6mQ3kEBeDxnOR4EV9EwD7iCXTCMjN6W+qkCydPz67b
bJcV3C77w7Qxk3Ub/7NZBnymawpxIr1YPmT9eaSdSPzi0bt4Fw66w6xyLwJmSpB8
IE5JGRXqUPyJMtCxddvOLIuql6NBTnJR+WSjd4E/J7hXEI+5L1h/PcP1DErFwLgl
Q7ngGdQkevbgT8ishoLWQ2+9BbwvADWIbLadZhPAyd5fgOHcuy8qAI1r+xFmZ+ZM
AJv/0Py61g7uL6OY30/JFOBJuICuNWiIs7XRZwgl8u5hzryAJUIDetIhOY09Rr9k
cqPbHf4Hpx8kx8YjKxzz1VBmjIs550xLxv5vEIHDxRkrNBDBxbOnBWyB6tgZnRYp
bxNMWpF22wiuCijEst86afELohuL7zvUHA34uJxmn/qRN2fFmo4VekTGslP0cnCI
SczLGRzMjeollIjQNqczTOwex4oRkmcK7+jZdiqewEq2+/zYhGCb6ZXlcDutdAVl
VE50MFG4KCeVw9R2XasdCcb+/iGUu+mHOQDPWmQgd7j/iStT0ae27QTCs512hu0u
iVGJTMJV4JSCwQY+aB/8j/KA6bZBb0HAstyCWVkIGy+m61dueWdrxqF2p3gnsaHu
Vwxmtzn0QNzZT4hLFXqZhdRmqcKu8xSncHKnUHaB84LhQN1dUGbeW8o3chTPBreP
DRa1277/BbSepqO8D/LxJOyXT57Fbei5SmIoAdq5WcPv4hc+hOdeqgcKz4IW6kQH
ej1Z+yQ6q4Ar5E7z9JqVrk3OkeGwFgbM3iDuGYRracLkmTKOGKfOjfEplna2IWd5
ad+GAtLRLSiuEtrbQu0v6YNLVE2LS74qiWw6Ww2LScVD8xJGUvidHZfedny5nwi7
uUsZk26lRU9EWJ3gmQ5ESaKn8pRYKmzQkGEIldhoscQiz2wETspRAp3XX5QtS9ID
xls8TspjGfpFCx1RIriORFbhSajACKb4rm0HjAwTEhmbezVmV49vfT28T+dEUB5i
leE1yYjzM2RDeKx/oX3tGu3t4JfUWI56ZOahczToNzy4Y9wdc4alZDITpFOxu+5j
gUb1v46ozhgAmDOZIqrkqECgfCOhYwvsUIKIzidaSsE7akf9OY1FDuo6wvdoPO7g
2caWA4W3MGBe9MCJCGWSySzIvVpZK6uWSqgZTep+Mh/EMjwdQUfkw+3CS0JKiclX
ao3PyDotao+kNdbg+6GPUNubVhm1+MV84zlHbH5nklG+Hoo2C6g7JwNPmFXMA/YJ
iL/UTkafuMM6yDyNMHtjwtpHokIc/tlQHwA8/gWdsjFnZiESJPSjC99/cDnG6CiP
fohOuOq6w4BTyhf7SkrT+Q1jGCMzyB03tnAPtO/a6f4LB41+0FRcprWUTbql/5FK
XOR/9OQFaDuNu9UrPjC6xBZMz9nvzqBCEA7+5Ws380rjYOvhJolNCvMIZOKkJuCW
5/3jCzoISTnrW7GS1JGPl10AlceJcAejYNrePQUlk2ORTJ2/EHdreBHvfDM9EeVu
ZqYout1JYz/pB9UO/Aq7Lwvg4hZu+32sJA2XsM7Dmp1Y4YQkdKux8A/bS97iqjM3
KIFdqLgNJHrK04c6PWw6NUB2QhHflOvVs7J9P+V73UveF4+jmoZ59/4xoUo8VNBo
ytVSRGNQqp2tiHThIuKkI7voOV59G06KHcFB/gftCX5lrDn3u6zoOuPa00lu41Qg
IqjKXEMf9DOUgrfXlDhfNqJ7Fqzp9kaYQlZzcNGVOituEAItOu+Lo9mb7eCEkUPk
65bVJ9A+vYu/uF7N8uAjRRzf9u6Bs8znlxUUg3NbwQa+G+Ol/Xv9yn+PxhU9N+8n
dbuFl80oqIgnZWDE9l2RSZOTuFMYh42Avcy11CSxJ5if2BxdX2VPXpp/wJGdjgCY
nrbHOhITjtKayrwpt2WXSSXfyd/r0cA79IFel1kZKuGNFJ03C1kUEjDfi1QQ8wT+
3qwKApT9j0qQzN1dSdrPPDo/PBXKo8gOuH5invlDTAncuRLVIDnyjVkwUgabZeYW
5ufarIkZ64gEzSXr78J2YxupGJXxo+EVTf3FZh8Phu6UOIdnhnW+Wk/MKBW+TvUG
OmuAhcgsr//ITCZ+oX4m7uhq/uCMmkT4bBZVMjApUeAnISkOWPuxmPOaeCMkpEUV
uv6C4bLN8tEELgkqpld8XTqrpQUcBlqcdJQZ1MfVdJKn1nsV1Rexd94H+Q+Xz8DW
OML3twyr/242NTBWSn2Z2LhjxrOcBuAw8wZiTRpMmFntwvMCF4iQjP/MRpVogeeL
O+8hcgRLkC5+FP7Q6yidhTt+ViAN6+m2BBYfWskkHzlQMgQqYFnvFUY0DUSWo550
Le0JpNoIJQNLCaG3m22CjoO3NosL73ArOg2o3HVb9IFNekBnhhVtMSArvARWzzKC
VuND6VoOYh8HtQcltRWPhd4oUkGZkqmyfelwYT15OeErZ2F8BR9YuutOO/ziLaAc
TBY9SBj3RYh6+wgm5YLHQ1oysG2UjWHoOrWmJhA6cjFqdPuNcmXS3rF9Ad3qylk1
/ReJoiS5FQIIeDiKjL2uk7lmCo8F5R7LqSCrugfth4npng31Sp0QFjZ2lHKjOGDv
sxzPAPfJhNumtmfplOMDRz3guF43x2t8LpB0auKse+FSHsVMprnUiJk4S98XIRox
dN2KAay+kVKbvQhVHQmHhRnHQboRvqdWbho/ovboSV1N3Kdfddwjwur3kdDLIeuh
W6nz1K+90E6E/qwTZeA1DRYlOBQiq0VHRV4RtGXp6GY9/yZfzHfg1Y6b9TotA2z/
zEwV517Gg66i8a5YlLnQlhJC1o4Xn8kvbkLwHzEjyjWuXxxbEHhocRLKJ7P0Y7wg
UVZWhnr0VMxKAUq/Bez0hqayWxJdR+pvgrIXHuOyo8SNaOrxIYchtCes1Y/agAYD
/mn69e+C4QcWZ97ofZrerkqu6a+K+RL1bhpD0XyL2GpsQmks8/f2eTmvcqFR9qJ/
LLJJlcXnWqph32/YpGSUIRiySl4MjeznGU5aSUpt0GZM+2EkXVRwmteVuOOfTAcv
Q94yFNBnAvonGUkq8ZfTJzj/WpLSOZ+tC7xXdchxZXiXKWTTOkcaD4Rwlnzre2/h
taPvSADZu2dImavrhnMzBhbmG02tEvl4uwE3kgug5U9IboPjwlfeumzGFqXF7lEA
5QQPft2z6RfLz4tx0ZaVBCdu9nzv2B2iW/RJQJJrM9BItkQHzpmMe5GijCmhQSwF
L7snGP7XmvKJ7DkC8gEQPACQnKdlIS27r9Lyi3qAv2wqVTVw+pPMBkgI8l27Wu13
jULRVa25FYJ44gAhbRLvqEb/OXsMuU3BobZZqbcoBmGIKK3/AV61PqTlGbTlO3Co
zRAugPUoYCJ62A8tU/3r0N+Irgk/wk5SJQbu1ujCii9HYJMdI2BU8wcSBMtEDKIF
SqyYEUHJi3U+vrXzwI/bG9F5GPkb98Gyf45nBmMEY9pBnfgRu89Qp0olAoYxl6UA
FngdA0AExwO0W9of4bc7HY4pGOUzCuP1TZdhwcXeJq532YfeCgc8CRqajAuJT/m8
+wBOAJmWqVZd17S3j2VxtB0q+uSIZiq01iZQ2Gle5MR8TMZUSiM7WNtVq65rK52k
Ij4tPZwQ1Fa/NPXGICgYVdy1W5CMuK/JaWx84FqcFw1xviBP+7KLrw6DX5AsewfO
MVkmabIafXuUAXXkReYylfxrM0AmLpNo3OZfxT+1xTWAU/NEcLs43ZzQdw91UaHC
EnwI6lHxmnqoQRHAqZ8hTZxl2xthcCWGmOywU91XEhTOHIGKD4ian5qwf4ecgCqj
RpNQgePzPVhjVJ+17ZVv6RaheA3jbTV5PK9IJ5OBgUKNrkH5pFJh6VNttEefnLED
oZh6rEpGxA9TmbkOtUPuWaCqZABeepNOiQh2iE9pANOtFnOPVLEWddThHdUrwyx7
h6mgGrWBPh0CNVYj2xDB2MpLMM7h3OodesAJD+dfoWmhe5XPTb9/mxdgy2+Kt45J
OPz3n8ZUtf7LKxTUnEd3Yxj5wIktK7SsSEnvVw8kTDngiVf4l8Mh8vLkkfAqskHX
U9p/Pn0GUeBH6Kv85bBl1xrGxhVjuUYJtaFB85ZpuNV4dxUmn7jJo15lCpSU6X1Z
E7P6OglTRkrKKRa3y3tfnEzisIwkMGCx0CPSMAKOt6kBeQRLZZ/B3cQvUKFXMTDo
Ys26LxDiTwPNIWvhQKQ7lxHp5tucv1AtZznuWZ+rhGatvBQoZp6Yb0MB//nsCL0K
c6NsxS/s8bVbWDibrG7PGPF/apETCGbo+XngYt98qCbTJLWyWeJJEhxuPhEKOz0z
DIcuVN2iZgOWWE5tG+yWLnZvCcclkvL1wntqtDRklnXsghA3Z5ls/sgd0caQ44VM
rQZX9kGa4O1N9E4Kc5Q/YIwTpBupxj30B5R3hSSoRmcSF0oznr9+yf6gdCuACxX5
Xx8EIyCdf4B613kKWdrE8TbTv6e3Ongdd0a+KSAxXxDH4Fave4UziuEtaGMVKAiV
2j94npK4ZX9rkpR/G+d6p3va/kLRMT+/cZKmxVZkV8JPc8jYdYf/rfb9YwGCrSfs
hPxzk2XE72x40TgbXUkdKBMGX6Bb/IcCZFhrN4zj+uEutZFjTGAASmyKQQReZrqk
QUIh4/1F6hjeaTrTk6e6i0N6wJc6R7RpmbXBuHThy6JIjinzAq3ApZ0OWpFMjsyM
zRxS32xr2P82XcVYIWmXBaE5TjEs5HXRYrRzs1l0Cl88ffuoC1xPWHI6hQE+kLJD
3oNwarjMoMqwBaIZmlYwS4om2tynzkWknykQs+8z0W6taVNVy2n1QgiflWxa6Has
BvJf4dEUKTpktGtQiaDQIm2o4ookt5UhhPXNll/SQna1OjcMzng+w0P0+31BfjVW
/C0qlQjfO7eLbrrR6r73iTqPwcD0CfpcBdp3wYt2SqmtO2g5X8gh3EjRbr255pBS
k2uLtYqyeVpJA860loL/R8vbM1Szduq1cRQoEZ4HEFAE230V5QjCRwih3vS9bT1u
Bj5WY9x98S/XUw5iYFQnHlrcvPdzwMJLJlV4Y/AJ6kxaYxeCWEX1aamFDZrmvYJt
+m+4e6oMjzSbgpwRMXaRqLus6KINCuu0wqMmsP0dDAi8XTqbDfmPUUmKCnyHKDbk
IGZoGz4/TYFzfgRku6OmRXhGSq1uAtAnRttltgxQIS9Xwe3MS3K/cMe43NcviDtP
b3p2D7TSLnLNV9q78/sRglLkiiaZy6npZTU3Lplf81bB/FXDqJsKjj/ZRxNIS61s
HuGpRDIf6quSSMZwAQEbuDq4XCz//esEZFyWb/A/0XWemkeuGG3+jmKfqId3Kw/3
x/6bmz39rCrH4G4GTEJ2cRROrigWMsQ62uEoU+ZU8DlcJv26oBkFZ06MkH1F8Moa
KJnyx3ExLnCnMzHS87riLiOoYh7silItTfp6C+tiyHDTnT/E3WFr6LtT8+m+0kwG
j26oe0f9pXMuz2/QfZd+LgsfNtovDotet3jI83wYk+7T8o2cLaFd864BoeAV2egt
UDeRwf/3HvVYWGSviEulz0iBUOVT4y0GI9Qyei9iAjcggvwFnDEQupiytaqmY45+
C5eFMiJoS6QZHF3VJo39CGR2up87ob1GkkzTBoS3AGvsA57APTDnyi6mMPyhVfDE
oJV1b4shde36gOr64JN2mgWPH1a4AIKwbkYl9zeu+Zz9GC3aZYvJ5WVWIiX5Evs1
yhg+PCrWiSeggFulwzYjEjWNRugiublMDzbW6PBI7N6k5yNVkAAJaHCSMUgrHLYD
SukHVveANQNL5mYEVwkDUzCJkx8IP1yrSTKPYG8oBBnsReBJLATSpXuFoMtfkoyt
oTY5SJrIcflqEASxwykPiFFRFy1emgVGCJ0GutB7wstrqy59dz791i9tVWDE4kTC
tx1hTnuJ9VrSFgkReuvzkesMHNkSg8mIWNeYITYz54GykKn8yKm+xaDInuqSnQ2g
IGIgRsiimlxLaqQSwnIZCqcq+6IKETffnhpKjZvIaSBN2YQZ3xSphwtQSzsu2fts
O/33oOUZfP2JDVPhRcY4awQAClujchracb9cDpapfeLK8bo7uYWiw/AHxmfdX88j
1wLIX1k6b2JJpEG8rnaowTng2Pgyp01nr9AX7eACJYaTzGYfmpQcOUt+1aqQBg++
McrNAWhP4UV30oj+KdD0LkSfQbwny41xbl+4LVKRLEMHWxDBp7e7TFkXS3yGgmv0
tk9OGq4heoZeB3HE7/BSMd/BiWztHwLuAQdjLxUKtkTux648HyAx6jYqrnR+6uec
cBcbRgAm8Vo25sj4QE+0h4oRBVFV3jkQHD1IP7Nhfwba4nBC830vaTunkh+qX5Bb
QaewHqfSfowup9RUiBy3nYYQeqLU+cwph7Jcrji/NfA4VwfoYC5pW54Ir7uKDFTO
ACSbFKhORoEjlNnZWVV+IbyzGgGdEquAu/o0bdBjlFtA6crZysQ4ChHGM/9jot7b
XbyJySkD0nrtwH+zQO7YoiUAaLwYQtulTpwqFv3lH3ZNXcIrX9yT7JeboPyvJ2QE
Ww4g1HhH6dnXyaB74K8jaPIrOYancEw2xUSf2VHhTfEP436PHktHEAN52ToEJffb
mG805b4L+dminA/whoaSd4imPG9vDV9thFhboUR0Q/h8eEIlV1vnhceTWtPJBpoX
V7oaSevqwRFdmdCK6XcPDEmNwqauaQD1ZP4sb8OmpbGeGTQhu2jtGMk6J3DuvbCA
YOE2G1YE7kjAhrIujnh6dKb1pI7J3CW3mKYY4R5u8P5GSpblSVvaw258ckfdEhWX
yfcPcsfjVM9/pFzWDjjv1O50FCSSF2c+bhOsuwSkMH8KKlcHeGcmzuC4dfAheDJg
zUdNGtqWx0svt3KwhvDH7ubEbOBCdTreOOfvABp2IyPn7LCd74RKlKw7sSB+fOPq
W5+FlDkNcf2ww7NQh4ceUhSoVvGvvC+Pp/tEVczV8d69TyleBN/mjPmYhdHbqbz5
NV2MtWQ5rYD/nwlM3HE5imp2C2MhvRJYWelclB33LrTUbQnyOT7a2O8d0p217n6n
E+pugMnxyJtdbOJcTRp/I8X0VLuasbk3igRZ0QcXPHOzz5/SKaSGTDk+PuPrxvX+
L3+phzCboCNGCREQ5Xs8SyXviqFJRvXzeYxiQYPPg8+qxph1IzYazf1Te7pYH385
OptM8T5SXOFta8OsoJYWkL3J0JIz8MKWsgykpEKN4hRQn/vmFPN5U4Fe7vhupL85
0zm7xpJPC1gclciookXE0XvG/I4pB/EShIuBHsFGsm5vj/UdhLXcTx+mre1Qnuow
8THgVwKe1K7DmEZ1SbzCJojPhxEg5/x6FSFJCM2algI51TzW3Q6BnFTrqjzsg4GT
7xtO0MDC5HdrGjCcD8emQjBThKCpwl8T8Xq9TZzpNNaPy1DQINSeKbGHHTnEqH3O
XZaRIt7b0elOGuo7goVQCWo8sMJrZ8t5drpSq2iqaePx1t9yLOgC6Nn6djwjBaI0
GCO1gArAjOwW5V2LniT1tBqP3SMjsdjH+TF6AOawOM+JZrjgF5Y5IL6bdFxCBEpb
I7qpxeCntKEDAxqWDsuvM4sbsVNKtZs32oM/TgRgrZZ8nI2+GsZNK4IHnHlPzLqc
4+4ibmp+9uk9uRyve9zWQoeP22i3G/QvApOxNaM42Z3faP07cyNcM/JYJpKQKM3+
hSoK5PQ+z5MSzecvlI2Ennc/CMnikNWwufERHqxp4zWg+x/eegAeQYa1UbuvK4H9
Hx65iuDEGQFq2HcrLs2X/exHFr7K2Vo1h41L7brI0JcgzSp+61A96ZUcL7hiQnUB
M6/wtrkDDdO5+RhbGMQ0s/QJt6CQmI5LJJk0hJTiKiHNPXJboIcFo2JwPziyKxz6
aa48gSxaX0kcywg1wvEtIr34ez7tPS7MM9enxLXflOVWja+CL2oGGI01SZRkRiFU
Q/157d5JOu9HFk0B4ghaludv2LiBTJ5uj0KYQOpqsrfwrBFF4qox1YhZd33kU9Gz
laFRLoRKiYCvZagF9IrGEGi92bxBvZyw6ZmlAcrpXFnj+pexEHKfIbQRN/8mXxfB
ftdFKCAgF7IRdXVQaASQbu4pH9n+GFGl8HiUzC25ALNzjHP0TQUdf9RaBRF2xOC0
1/+5Y7LQ9648eUgN9kVNhwvTW2GIxa3pNf2uqsFTyECJG7arMcL2RmGZs7WSyaTN
/TQeLa2zoRCmhZ+cRRfgAs9JTj44XJrf7RLyJQcqUXfJZKJJqh5AwMZ6ywQnCiuf
cBO/my7kXp5T+i87FNL8sG/7xS44RYiqxqUQYqerPKYAw25pX4Ay8xKNVfwC334I
w2AczZcd0OSG0Aclom8WnkGzS4TxVmOeuyd0/JUo8DhPPPuyQKWrauR4Z0gx276D
rYOzm9AJyau0OEcaGcqwoU4oeT34jqocumB55GzLSqfcmMJ4VnhGr4/a1NQ9dm3K
`protect END_PROTECTED
