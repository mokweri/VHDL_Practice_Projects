`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gJI79phB5HDDxEZCkOslyMC9QItZjGOqB1p8reqK10JhHDgaQIMm9LbnHoj9zsJu
c68+1lyfcNBuTMXJ5UDmq6YtYpvkp5rTwjqYEJEbVQCASUgMcKDvHI7euIemtI5N
S25NI1v1FJNBh5g/zGvz6da6iEL3BBSFFFnIq2Rt03THXC11dD7mJ8Sh3ZW8632F
7xOPcTsy6Rwr0BL7DvjWNr/3I4bZNqrJ6uPo3pkNSneDm8klxv91T3M0vmRTI71s
6Kdj33KP6h1H2lpdpsOElRj/OIWGlplFdFvaZjJcLSqxjVjzJth+gt0ACjFLXHJg
gM8MdZcOIhypI1o8Q8jWP8fURVNqNIeOZFVDSF89WUmbAoBokM3N8ZUhBrKulWGZ
5olK1QLAl61JO/LrlstFtfZ1hs/Knhtr8RnSFyZR2wvsv9WOjbl1bCKD1mXzembQ
ghZRyeM0W0XjocmBP2Oe16U59EPHNYXJRbBb5iBfHJduaIADBAK8m0TgObnH+dio
sSgVy7qt56E7UWgBpIexfg==
`protect END_PROTECTED
