`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkstH2vLONl2kIEDy+kmzKQNd7aJ1tBie7R+/ToyGoxhV8er8vq4BRaZhhmS8S/Z
c/5A84OmWwWZXPy6e7Io5l2URrR0ha5W5xlq2y7jqvT5q/bguw3spWtqmMP/GyR/
DF7O1vL6/yAplk28RHBor5vg1wxC9gcK78KDrJUrgp80QJ5LWWAPTrq+8HjIs0D5
hjEdvm6+nr5vwf479yGp2ZtQQf4O3C6IFrrUtV6sPRI+Bz2f23kkJZYOrKafg79Q
3NP8UAvsiRo4eynlrVD6IW3wuVrKt2WsPGZQ0fk1AjV2a1XLLzidQBfDKy52hHxO
nASYLdm0oGFwORu4tNg0aiA8RzJG04v7LgfzdLUr62OYVbocrshTOyh2Z1b218mq
ZKmoIKssnEaW77NIYTV9pWo4mLfNv6KN3jOc2R4pLLMjnpsw3QHZtl1UjzOUQrtp
REQJ6cNB5+IrUxeL8mUwoc7S/QgMN6LtSlIb4N900lA5DjkHZU0S6dURghe3nNvH
P+nRCTVnjZFic2JuHZb8IpiM6Of+58ZjwpVe1kiPZUafRvQDL8uNT/Z720/9eZD4
jW17FCEaQcMe0Zb1ixzgRzrEFUsLaXmEqSaRLwNblQ4RCzBFIzq4T+b2mwlpe9us
GMGBCtvwp4pA5YyvUpGy02f3VngeqvuyYb9v4ye7zt9SRiaIRk+TA8+cD2367S0J
bjMcYfVOA56DKBSgqRVAgQCGwqpwOPYFlu/xIGnchs29n/s6LObU7NQqULD4ahmF
ipe2tnZagUFQxwap2tyiy/lYjqLP5Vy1RhU6QUBe0jE=
`protect END_PROTECTED
