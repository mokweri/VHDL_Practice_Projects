`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pvHcZO0UN1pV4g+lSdiiPRPjj6ha87rlLHuMZ6tMV3TO3w3VIzCurZzJlFjOitE0
u98g3omrzQO6RUEqq4P9G6eKLXmwj5oAAwuPIRfFLb68KO6Rnc/AMrHOWXwiuF2I
mNrDKSt0OSO2fuGAIet0XEhfNj08dAQ8eTdU3Aa6V2qxDyRBGVv0oR8BaaZ7yQAe
zsLocqXiIgLOLmzZSBfnN0zfPGPsfRe3r+po3XIBwPSC3LW2fH2FcMbD7bAPvYKc
cMz/WNyBSP/6i8UcUYAjQSbKD/Grg4+245KWrT8KQETgJCbyklH3txwLJMCnan9s
lTWuIA8pT6ODMpF5NY8GV05744U6pXyYm3jhbjyQ41tG6o2DsCFgDUz2vMeKUMfx
ohlJdzKEhj9TWMbRlBnRPXTZwzENccHvKUobxenWzKX3DKPjoeLi7rvXzqyN6/JB
ggT0qT1KYYNDoxD3OSKxwfw/zNHo7c84brTc/Lg0KDkB9seAnxFdzsF8pSBTylzN
1zgElTCHzFPKnJmeXp1mJqQUp3Qh4yd1sHxTcU1j11vbarlfV1xbRKJVBDEH2ZQn
m5v9xO4foOQHru/2f361zFkSKpVS19kljoAfXReTY15OPm5AFE4lv3EZ2nfnWA5c
6aAvvRjScwMthJkXG7Ba+65fQvzmD6eCFwXvr6m6mexkpB1BcKWaHQ3RVjRdUAmw
UvLuvPjUPzow7sepst13IS11nZW3vouMoP0z69Ttps4SLpMbLyh+35XmRoWmUwK0
L7ZTJI/QpoAIMrPOjnLLc1kdYnKukE1kf8SNw7UB6QvMwZUKEhDVgrYGSc000ztV
py2lv2ZfJmpPk3inr249oiOhpZAWmq5ZqJzSd1Iotkd0k2nXAATDfbjn6UmZNzSt
2MXKYM7dD4MebFYwY15YXWPZnfofc3cJwAFbkX6HVK8s6oK1iTzFRJf4NWCRG3sp
J4e8n4KbVIamrInePBHDOjvcHGv9bshmkDvN0mVJwSG8H/gluyKLzATgTmmPygY1
knBqW2XAn93lj8dHiWNBqhxTotRFovrFH83cklAn5rHwTfBT+bKHUnsdpMxCjcQj
LeiM9oShYllBW7KJUY7mRbaFYJbyMrp5HLx3K7thVFg=
`protect END_PROTECTED
