`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4XmiG1i2osau+8IaYK9O2oAYu87FRWcidAOxkofKOC51UiO+HMi9eRMpRIECyX5g
pN74tb3LPPdkDOSS3+opYZrMSWRCbPsvtMDfxwiRMRx8HOEhMdTvfW22ZDg+tN11
p385LosYgrZ9Lj7aBgXZJ7wHcNqCvFyMwcnapYXNXgKqOVy7VwkoG4YmScONZR8o
xT2ZIM6YH4bErqf3bMxQqo7Jg1E2YVbyY7w97d9FA6FURzzT0D/HQH6mZkcHqoHr
gXEYuaBq4aqAPFFLz6mqXjedrE/SkudWv16QY/Ya6yK/ahhhwVK9BJ5Iqyb3bAZC
L8qu6rAk0USV2bAoYMfPbbYBH+01O9wPpjqxhIlSqblxJpK/CHXB6zKx4YWqK10D
5X7LM72rXiF6eAWY42oWTKeiF4Vb+ocrkIFpG5GRd+RikRGWlgwtm1mqLxLaA5lG
dX7fyU5eKvkTz5Op6Eqx1nouRBrtVtKN2x5gB98vuH9iLUtB/rcJkJ/teKzmtPCl
c1WaGg8PihpnOOXEWE5trQd5JdwEibhp2iuiyIFpMMSEr6rGYAm0MGxAhrTg32OH
4TZMFZMJg9UjWRI+on8Yo8WKkPNgl+XlzVa1C34R2kk4B5GTzuarYd4wjVMxGX0s
6zJFl10jqWxVo8gsL+4+H+U7+Tp70iUsIxhfYxQv+FpwVaw2e0K5NjDYliAmsKnd
08EU0i8cdQNGM9E0PfvoXG1PsrgKymWmHFWVPxOOw9PZy8oyZeY0BFuxqAHMoYcX
nVByyw05KjUueI6nKvWmjGcnHDa7V1J3s3HrmhYPuUozR5TiNLfEMLqv319GEKYS
Py63SNh3HoY1Rd5lAEubRKG4QfhVvMw/wDljO+nscOoUhJusm1Ml99g8Tk/d0a2H
TENbMujuSbgQCnhoQDwY7Jicq+D9mtgTL/XHJUGmTbdFOWCot0Oc6Ua5QE9T6KVY
Fs4ohBWcl1KAVZNVNP9zpqGXWM4nLPZZ62GH+munDu7zhwRJ42Dm/zl3qy+m2hlm
EZLwshnfUquh+gJclk4/qM27jB1YIhKzbQ7Hr5GrLLWcQ/pBYvwYWkl3G37nhz9l
lrsJC+ccL9xjJ7sC47lVtSmqx5qYiHWD/MoZOhXaDQQk1eloKx+86zbqVATNvfxJ
QRfAbRDyhRIgKKl0sRjT0anEcqWv7shdGZQMBTIjYI48KtGRoQVtEwNDF7RRN0df
I7yufHbxJGuAVkLSxiywJ2AD2JD4k5BZupcew3EFrEunI0DRofGbQPRpe0SdzR6u
Uz6XAiTv6HE9YbWEDw8IF2/e48b8GtTIJJxJ1bFqVMHzqGb9U3GAHqlw9JY4QHAo
zgg6Z/i6vj+rsLcoRIJbQCsGcfd/gEaQzgUNJDrQwhvBGgYd09W10A/VIpDw+Pxz
ZtnvMMVI/nbL8Jf76abwd6+JwgLtI3zBEX7s4PesJF7Hg8fOH9d6Y0AdJFanURAK
ckM5Hlv8pKTTbaOy0ioBbcwhetNJFWJUWHTzc9Ai54HowENLo3+hyIaY5/BOdbA1
XaDVCwfeliqi9dxDrCKMlmp20tmngXqlWQMJdPp7ZAS9qiMkNi/1/HQ8SzSzyXXX
ZYLo4Zek9HEXvVVwjOmkSl8JeE5LOjQ8NFuZxFlhNRysBxEYI1N8pE/dRza9lAAd
m7MNeztPA8SW3O96eWO6sCP8DThKUX6OK6UptcRZ+8dIuxtCKD/31M6pMI2zMDjN
gGR/Iq6n9cAo41HE3ybv3WfKfVJOa69Qno3ZCCLNHXxyiTMUXnbX6fp5vUJlSRGq
EqBulMpsVE42O1GH2nMdv0ij9HQOVgburHzWUYwztKL8x0ifwBDOu7od1vQa1i8W
G9Kqcux3T9g59jezTMAImBO7SZ4X/AkKL23APof9m6GPjU7UHbojtddtBSyhhFqZ
9eueC2BLsehjV/L+WOF8b1Dc4g5fuhw/9eqw1bFjAKk6A2CFMMT1rIFbcW9hARNh
C0fy5hmAVnY45SGvbJ8MfNDtDi2AIeqh5SyyG0MRive3oK5Vatx0ZEyP/KBn3k+5
pBCwXRvhnbpwj0i2TZ4fFJRbhuX29ysKeFEyt+2pK8QQg+yg2c9wpT83HGD1hyYz
GJ4R8vx6SfeceeD/n2Pj0QTqCeocuVt9yw05SJxbwwcNWZj/3VYrt/0vWXSWUVt9
jQPQXN2pZSB3YPqEZ9k47s7+EKsDDXdi8wwGCQ3kKoHcmNTw06nQ0a0e9EpsuQhd
P2XBtbrd7T9eejefTHarJou3xJEjkC4pBT04VC+fRwKsen1tScleFlHugfcbewdV
QI036GIMkpRagB+9HYkkstJ/6T1+ZVY/TBEuguNaUduOCP1AzGep5gNSTX8TxgTG
XBTNqn66vwJNXxkjBE56BR78ril9FTQLxVr+4NISwdinWmkL8MJlIfZB+V+CbyGN
bgw2lG/9+GaSxSZCdh9JuiEyyS0HmDSnDrCdBTR5eM1baptTVmvLLI/WkVKfFIbS
XtkOvhXwPGkI3fJadilqlatqlcXDAyIWeD+lzYMuGMFL4vfACoq+HhVccUkeqVKy
aWqN1tyBXUO0QaAPkndxbNSLvP9417tE+8L9qfQSWraCXhVLbeL900MC+rpSqVz5
jyrVYbHOitRyzL9AYMy/DMXV+Kj6HB2MtWbHy8nKNELf3Y46r1ChQZG2ZN0oSk4F
6T4ECFbRTHqh9QyC3qBE28Vhs4AcQpOuoMtmgGSwLjXJWgaNkgM3CmGN8OmozRU0
q1ZN1vRjvHATWI/bgZQJrzSZFpDrU5nIdesBeQbzEAETDJrwKE728DN6fruxFJpn
PVH7nfTK9NMrIjd3QeabDJWEPrYEXQtC1eYP4kVRzlp0JIWs9WfYQmL9xZD6Ttxy
NgDmQhkT7lKZF8Vq94pr2SkhzbTil60GGsTL/08FcVGRCXHaIe2EW5/DKwcHTpK+
ZDfh/TxGmhfGEWWtPGuP58S40vjGvdVTG+E0JcENu3bxqQ9RNeHL6u8OLjnUgUMv
x9aPuCNjcqbK+f/Gtg1PqcEaX57LHN2wZ/mCUOYu7cav3PjmUkOcxjpP1rPhVvRZ
aps557lPWTMx+Jv2bgpcUMvWDAtAFjHyE277ywz5XVr/GbJ/WLQveXP5zS4RvCcc
L0s3BdVtQpIWi0Tb2Y0vBFj7NfHvv1DN6KAwHskyVCR7/UecLotEGD5twphpYo3A
MH6ybKom369mGRf4x5QAbG9AZBA40LhEowY0ZFxmri/b6xmio7do6EuJEP3s4ATk
KI/mc4v6LFFFdDEuW5MeOk3M7wr57zhcPLXZ9OGcSRUe8wtBe064XGtdtdv5NEZq
9vjNrO1OP1/Mi+WhL/EAU5fS+iPud1pOH6nBj5irCatdGDYDJOVk3IVsjxgBknFE
Pr23gPvPCatQeXgnVkUS+lRdsNQHUH87NAhYQKRHsSlWS+cOxeosYRFMbMTb5350
idVGw+bLWkGIc6Ri8X4T8MzW04N47Fv2maP/8vbEw45Gz56NeCkvSAmeFU1RZ5w9
aV7LbIhfl7pQTFqS8+fObFc7M81eYg+D1eKH7iW4QEW+SkBLEOicO1K4gDrISN/L
L5XoFqGukuNgP/Jr662Mk7CQ8I2/Jz9kLfnmDzRJkjI9bAPEobiUtCIFtgFVSkJZ
mvnZJMydnRVIJFe8HVbZ5Kd2QLDWuyc56FKkc33U5sLjXZh/n8ytEKFaLfulUDsU
0HH8QMlbpO/3jfbWyTLk3iPWpD2s7Y8yHp7PS9e4PqhpTRy76rvduUCrkoPVHoCI
w2EBL+xOvAVasJGtDYM6nsZ2c0WWzYCRw3cA+N14kosu3hG54IRXQPMVpf9lvFT7
NAtX4+MC2uP2LYERbuPJqq8AeptNyp0V987JaxkU4uANyWc8DhNdDgVH1RjPiS15
jeaCpCko8lYBRMASCvPTsDmoL3kCypnQlAGwkpKMigIq0C0Yie+eRkt2ifPqShcS
JSSVqk314T+UHnLXE3o7WkBRRlqDSwW7QbRJX1TDD+dIklI4Eu1rlnF0inY4e5nn
U3XMsWWsAsgin6eAklPG9aJq6Qd/Q9A+Cf0gFaAxzYIMsMTTgahTXkuvUe9reeBy
SYNZN1es8oVE5gP5hmZzHqjtB9iTxF+naawm0HL+NHiUQavkiT5Nc8GEye+jTtv0
N8u2NLa2IhrA5W/nz51n040ncoxDtKzWC6HDx03gjjz4/NlQXNY1oQew2bbFsR6x
I6gwMQ2PEUy2EbGAuaMt5P1PLlCRfs1v3JfF0A7klOu1MTt3C7xzwctmSCpgYAjj
lbzxagl7jJMLHOgem2JY2XVFyiIrm62EALVUZkq/DTrj23eyAJ+zjWAbnm0cXEbE
i9Jg2dfxJCtpkg2b1q5Tc80Bq8RAhEoKaCCptrdlZLWV21emlF6B+EZpPAA78ve7
Km6Po65mGiC+TWRq7WNjrPcutwibwPCtPVJBFYzAHxhFVLZCXto3Et/t05tcfsKK
1wWwwLImEQYM8Dwj41aroQwEvybNuuY41c9Gv31ZzBQP5tiPb5X+551C/eZ5TvV8
SC/yTPl/VezoeVzFpPqN/5pu5D5r4ebGZsURlsD0IkChC21OKf45YiER2toy4c/y
6wrsen7PubeweMIS7GRWYWzpnMGKh2wBhvgk6GCaWYz5f4gNMasyRkfKveHiIZYQ
S8Fjd0o4dkRRGnr/VJdrjLGGSRUehzUkXAj2ODYmVB4bKVstFtJ4Fxlxur7v7tzU
vUgzQDxpR75KP330OUgzlcE18Y6CNPzi06BB7+gKPuzWeoMDaZ1j6tpg6CTiIaoO
f5vkTKkwl3y/JxvzgJeh0QuJpPzhSJrEaGEkj/Dx1lz3JN+5NrJRQLH2E06B6cbg
85D0DF3yGmPUGx+Su1GWTq5IVNIVnwb95G9US7+jV/7uLCem8a4oXZzts0mJlYz4
VHTY3i2p6XH2MGgHyddQxU6PIKQTD8uoVCdbd2JfPZpaAO17p4GoOZZaOgj8v7J1
P0gVPZdsHFCVZONrj5rNZb+zqPg3SlRA795F2iNAtsa6s3b+72y+BQgyPQU6niP1
GG/Uk5Js6ln1sNjxi/f/TXPAoS3s9c1BfzN6hIJnDyd+1Auv7ChwYAMuXQTXmJkf
5kvJBsZ2wi0Y366LhDlNW5rQCowT76533chQ7r12CFPJG2kg9yoBycBFB0vwa9k8
tccvXDUjTq67f8lAZvPllym9qPzXMtWKo/AE3cQC6Qi6No/zWMTJQrmv8vWnkQxh
zVb8yQAiyLp3CqlKPgkDlmGYcCUX/MVxXNIDbA69pOX7DU+bOP0DgrSBIY95hr5k
3RK1+49WCg5iwGkM/G++Xzevuq+CBWdXAGW+7MmSU7aBp3oiGrgMuUfpD2ar4/Q8
rXlw58wwtSLEwQyES3rkxkk2WtbxNDQHMWvlKxH77m1Oi7zOpZ3Co7xVtgGntyll
BNKvWvnPls5uTJ8XwpnTN801EfjKB02BlWEVq6+JykxT6ectiKKnhlQAT0ylQxWU
vWPqGBB6SHhaKOo4ZRbiJSmqEFOv7LcesBX6QCllDbc=
`protect END_PROTECTED
