`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kVJZXVYSHu3ojsmA/7Cf4VrM7kDTwFYffKHm1S4z7xHBB+2LkKcUmP0ScQNjm6Dp
DGzAHedBzDicQ9KOR6NS+2PAaG/k53kTCP3pMW2XuJdUJZExqh4DQ+ny60Npzf0l
FAKUIzPo3kbacF0ktUOTE98LQ+jSGBHOVFIGc7981XioIabLtoaTW3Skmf14TfuN
u6wa3QR7nEUh2sJ2J/+FdL/f/DEbtFK0gTIaoS+9DI+jWD8NX8TlOXep1K3hK/5/
qPC6IVkpe6AjoYKzphjVFExWrrAQF/IToIUfXXADkMKd369NnIJWtSQUgB2zBbJS
Wcu6ztPzKsBkVYDj3dq5bJlqXsn8YgZhW8gOVK0Ccj/aZiJES4qb3b3jF4anzgt2
S8/kTou9qtV6nngv8CoQzNpsqsXY9z30Jux1YAsntGBL4BGpMGTjwf9KUvKnrgKt
Z0++JYPzJwaC8gY50qhme/cl24TSwqz3CsJ7x7oH099MuPnRnAeSbUNXHlDzSdPS
/hQGlXgFvHiVNVB/TA3e3R7W/RTCN4XofBEV6KQ5HmwbSWI3xCSCKuf8GU6AcO7v
h+TbELdLpCLEHaGumHuONllChGoi6uzrp5G+TQHYhmU1+dGJbYkXXid6+EzUOkPz
9xOw1awFh9t4c0Qf0RvKuvXVi1/7tfzPZrVC8njobO7BRt1VOb2Hpime388C0dFw
ptBQ/2qeIVNjZJ8Qe5Bnkj8B0iBm3kM8vESosPcwi0S9yMiNRzuavsnIPSMl+YQ+
sa2cJKakpavLwExoM524dwsimUcqL5BwkcSq+1AG++YTrT4F47BVcGvsBa3sWYfu
SGmY8b8Ys0ywlZvOkhVsXELxjoSl439AOtReDuMiWNKq34yqhLNoTbnqG28w8TyL
UtEqE+/bPzc3p+/2vahOTmC1eelSEXuPVxgnYtJRBLs5uqgQsM05TrIv5vEr1lsW
DzF/ao8kTL0wiXp3UIkGNFWgQrFHdlS0ii9LncCceXKvdgb6ZKAXb20tNfTvpNSg
e6eFD28p0Gk5kToxkgBbqTX+MYg+mI64LkrBwEY+dQCAVjHaC7dm/bHhf2H+jZhU
beX0F2aM/fj7VyXOymJV5yMzxWCDspcml0mVpMS0Qx0PyaCF5SGdLASMd9IrhYha
3nK21/W+HWnzfx/C95iyFrj7q1TRRRNk9b6Rfcz4wJcVMMSqwy5K4UUnQ2H36ZMg
Upzh3vCMwUDoDooX6PWFH82IX6y9gL5vOJu0qVJmnBzkab8Xi6m3Q5cKgUZW88g8
qlLBsO6HSorTBEJJshVKYZ5a22A1sNMR1dVaNa2nq+Ew3AFUr5qxAgExSrJ4iZA0
IaFNBAkh6REYdQA13zdgz3tmdqPYSrNn9mX6F9hX4Uvt8WxyxM1t76sPcSIDrwIS
JL2lxffV3ViQhH5LgkyVmMWuvpkDGL3YRTQ+/5noujVGhR07FylWUkK2Mjznncfm
JaItqmOyd+Yh0Fo29chjJ4SWtZaG0G0FzW/zNjy32FRXCVTN6AIKhGMLaZvT4jSm
j85vB1rFJZR0QJTzSc0a+G7d/ETmVWvVJ/+krZqall6B7UmovREbTmMNHu98RpEn
C1XPzz/X80yN6Cd3Vdh/O/1+BqX8h40K54G5U3r6I3LWuibdr+9olV641ww6rGvU
qm7kne1evfqt2iLkySMP38AR2BI4f37Ad5iTdugRKuMSbx5KajP7PpVK1xNOKRlQ
vl8c0T+fBSicn15b0zJ6hpRmmvjCoIkgzXoKKUCx7Qk0V5+rmoPKX12h8rIlCUcF
az1koUWKiBtfeyQJUvNSJOvdaAgaNaL9O+46fOzVeVpdlwGz3VqmxRBn7qYiF0sx
excv4U6/KpSsycI+4ILBc/Ey5mEGZ+JdH+KtCNsmzSHl14DVDZNGbaL9QEOlPkaw
j0U3eMxzHM5GnNf3pChhaYr4mqMY9jmj/ekJHzf+NmDat9jV7J9GumqjdciJMsG1
37DysUqQnSHYtuKrQlITazlHUgLNiQgqZlpDkO8CX76em7jKRLlgCUhmCWUdA8ID
PImPu/oc0FKAQAneTEzfYOSehGtcn5bJ8/gVAxggXruhku/5hQ4V2vaB1O++UhdC
ELsGB1diYF9IEKpivlpwv5JFn2o6zVmUfH6WXZpJm1YpE+hcYBEF1qxnN9FASMCT
LUcvgCX6MOp3U9RRFzz1gFpdhvAYW+PLrlBeOyIz/3r2A6P6SiEd7AZtVGOwwSys
8Y2+3y5Jkcz1tVQjIVhHQah1moLN28A7d4M1yWIQZWoDxE1EmjkyN7Eg0vodCtFe
gJzhycA2Dr65GJDiukV3wNh/TdsTeQZUZe5QFdF0D6ntKWrZWd5Hexq0nkNlgNhl
dmzZXG9YK4+G24mIQNmD17BczTntPLpHmM4Y2zF6rj7iXk3cAHN+CbvMudW29Nub
xAwwdQRE+95XTXS+n1FaxrpWXMG89FaGMv1bMWhai7MOnDGWYKWQwPtCqfyfTKoV
r6riGmNwX20agtkrgXBA5dHb3qSVBpAu1t9H400okUyofQ0Bl/Yx3hvuaOqIlput
ZiH6aJVnTDFV1Mo6D3qbc8GYkcFocpORwwpwXLSeGb0Omm4bqZ/lcX8suboXCq5Q
ivwj0r/IR4uC46rN/QixFx00F5rxub0e7tFM45eETy7auvwY3mBtSLkr7dS2sQdv
AGk+jVmXDkLnIc64ACywq5Op5CCWPlEtS7nhlYOs6UhO1pHtPlZzmtnDbauw19dx
9VpOFZQuCf8y809muvDFZrBg5/50gLqUryYjBYgY1+PE97vG3qS12zH19Nq5jdZC
l4Ehq4DhIex6VNM7bPxFwtXWkykvQ8ufOrakzctmcQniNmEDiZFP3BNGsTmZFVNe
jxhp/2qiRgZBfbKcM0SfFbIxSDVsrFNWAiC94dDatXADwaYfzE4f7FesTtiINSgE
8iHdUrhguBvIP/szraTF6ouPMzPEyCqHNw73VlkpQvw+kRknkINA2pVd48/QDgXQ
9O6QHCqJ9XDyGXX2GlQaOyU6QuNbshKzD2ILJW28yQLU7nC4LdHVbUl9zs/zKlCR
JUhbVVMFhRivRVJ+w0taEJC1zDvQHep2n1EUjf6Hsm1LaI8+FY9iBCcaca9RkceF
T5UrNuiJugJ282MrmvGrhlAk4iGNmDuVphDvP5vPReSY79gCU4+riMdhVRVi+W6B
fQ5BnawhQtlIM45yyv72g9gxdQp1m10VzrnuAJkObgFdStfGTwlHjuMhBV1k/dEl
sisLOqKaX9tJ0osoiPTun7CgnNjP9yfB+n3Lvc9BFLCxMsNUXgloZqjYBH/yxvJR
QT9vRlP5dla1CZhCkDObGwotkivdTEGdHw2lqmc1yP0t/RkLbWlOJXlw5IS7Max4
XsiNgCkKIYvSezwNA3ICVZ8qEq5uBAa/UIDAhXIhhp44hMB4UoYqwISByUyJvFul
mGxHhXWmsCwoEg/YOiu90Yj31Ov1jhIiGDVlCCKyZkdlBxa1tuwLTXbFKorSJBqx
ELMNMidlJxCQJtq8qsMLd7ocx6bQ9KBVbu2dDjT7ZnEf/PxWtdSXLoII1HAGCEN0
W6sGj0RMWsi821ZAI2a3X/nVxquBujcs7Q2OI4Gfj89XXlkmSPJ38v6sEpUdfXF+
XoqKYEMuS8zncVERrfatN8u8hZtrmrDK6khppHwwyqVQqyhtRD4QoKaJoRFZ0WE+
2mmnQvY5XRr2PFSSHNAxtjxAPjjAUs1alAEPMTM7tdyyCw1lSR2m2N6bvy5+Sqnt
yAwuML/yXX7oigxGn3OrSwXf1y0ucUwph79/Zok7ZB4BceHFywAL8jV5m4FcXgkY
1NgfSoKssN+GME0FmrYiUvPd2vE9q3I+iuGeciyfc2RGEhKaqqy/Jjwb5IwAKaeE
QlJnkqgu66WOQSxHNrGcL8DCFyMDAC6JCXwFQ+4RCo8D5pHpb2PD70nPG357f7JT
VdDSxF87xAf3blu3i/ROrjqIrp/nZ7kNRIojT1FWXtK0q3Nh4xoZ+7NPcQy4Iju7
+MShATojm60KUF07kgha2LtjixWkqUUf9uFCqlGwAqPMYhC6sx8F16IaIHS72wN9
pBLwcj77P6GdbHjr/INZkU7M1gRef0EZ4Kl68M1ZYcB40hbpq87YBruGBF+Z+xaq
2MQIwZCQ0Y9MLV1SQB1kteGxwqbEY9Ux6EjLPWzTTJdQA7GWoSciFHJjhO9skjMI
Wqpqbp1wbintLIefgfzPikzZRrirRQlzThwrt/SK7g6Ozv4mIGikCAFZ+ju8PdeW
nmosh0V0JJNqR4NJNyqdcqZ0JVPAfM6rfZT0tyKJ9qOkob7XqMTFsPRa8xxH2fi+
BswdDXofqIJaHxBP1XVWMPOOj/iCis/R/iddltn8uDWmd9lp/MjzsrnujA2lQ2Su
LsEBp0MXwSiBh3dYVJ3aoHJn9lEUYVhDJ3/+yEMNLb99VuM3Mas7f/oTXJvR5ugc
nrqyq+yDFB+K9gs7acklBPB2wreJwJiJuS3Nz8L4Nkid2U5LpCLMP7muYSu9sxUl
luthkkCPJj1d/QyeqAAdZomwaX58A+RZ9KjwyouQ3v93EGmlXLfJ8d3NlYnWS69F
LWfR9XO6Bu2GB7HFVqPPBzTGw6hiY1qWo+x4dz1pCelEPUF1n8rlMIj26yTq7UGT
fh+nflwMqDcbXyFDe+TVtJAeDBvyaFQ05U6VOJKrxPedONRjD7hxyBMfHo3NNJfw
5/pnVEKscF2JPGp/UPQ86xJcf02QwZKacgC6pzA6DZ7R3lcAR9WpvNyUWU/0M8jt
EJg1pKJ1Lb9QXdxWfqw/FjZSS4b6DnUfrGhDBS8OyeElgjpcwr/GlPWQ321cCukG
ihm6MU2yCi4U6yq2aav4iGDiRVBGL4cGDfv7mLU+niij4vkMKHMB2MtweMDsGLUu
0mR1FHtNeeF6PmiVuqIMPMeREu1fQF+XNZURHWyNqG976bUQ0PysjqMMfTU/fGUS
m0eLjWfRUUHWw8+2YNUVFt325cnzPTYqbwtRd3gi49qJxJ+YI42Ng/5udh67SdQm
2df3se7tnwkbayhd8hiO9SHiFVnPTuqA7Ipi9A+np+vOPvAPNadDaQqIcHekzMQ5
n6lc+NMeYCXBSVl0c6gB55GJfVSbRlnT8FFOFXLon2PtvBXm0dEM627dE0UGJlJn
BTfLnbQ1nIn/5PnUiWNxN628tRGizsJgNfajUnGsGum6jOR8G9Ryv0Hk6SHk3Hid
7zIxwDYIzQZ1uD4KeNbOQG6QCploolRiIcVYTIuxYWpPyU1mQAqMPkVV0TKd7rqm
iEPv7+w6/jq/p26qDTKyZ1AHZq7RaKC1WBcYF4qZARhgji3YmVRSDP0uYYShuqc9
8c2q3V5scSoehsjdF8D6sOc91pottPSJE96v/tZDSv1vij5bLzuP1+CJwmaRHzzg
fzt4MnhzGN+BDFeQBozFzG+VQyZsJD3xBhIvd8JwCx+wposMGt+xU0E7fiZpjfGP
YA6vo0MjbXE9bw4ifnWSb0NxL9OC2I1I+VpwbKkgVxLyipG6kZhcafblb7ksSi71
F8BWtFY5GrId33+i+XHXRSbkL+BFxz5avlk3vQ5QbrsECpbfrpgjlemjTGNAcJF4
mIqIJZJqo3F9QXQVKCbPCAIprkiwWDSwzpF2qU3YxaPKOxBlKwohVHRxd0uJsrJj
xog8f048mZbzAvUkiEUGKDx70ZYrTxHPePyYJNN6SG8Jw64Hzo/kJbMf85OSk0yV
A1S6/V+K8he+2zF+mbUS7iGyNE04TqEL7IU1yREBsV+hFnO6bGxpVExgvOlC7gGL
Rf0NYge0HZmYgtrXTS6xSt6StwknZU0xdN3mEVw/uBqiwe7gKKTbjd4mBBqeQ4In
YvZpw1/OLfNd1QlTNgdsJklvEBsoL7svsIaOvqDEpRCdHDqo6Ji2TxI2t7XIy7NX
fIYg8tTsH1aHXU/ZjaOCWLceGEKnJttXMqKOzBWIaGR00DFWbj/06qhW+vOhGnSe
fDfihk1AOMeBZ1B1PCkL81wy0oq+CKppHwSryrS3Bf5W7TXC2giK8YGpC4SFrt1b
6uQvdcHWrjY0dVajJ1yGTqC8Y9Q/O7FKbwhVD47j5NBvJKpDd18oK5BLV3ibtrAB
rpxOrsgkSBamFL0SPGFQkK64UiJseKWvE0bTBqnGB3KFh6izVb0XzEBV1p48qZ+l
k8dV8pFFcyJ4r2hMB1nl6dqjZPEA9A/WD0tlasc1LlyPD4HwBO14awadHHSp9EIo
X8WOKmk4TIeG+d7/aQu5DARDwsowLRGwJndDlkDta+Z7yk8g1AzYwe/SR+NK+c6i
xLYCCZbqjVcUl6xLGiP6Nw==
`protect END_PROTECTED
