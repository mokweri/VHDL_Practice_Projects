`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdD5/+GqK5USwrICshPKlvBltTEJX92bzrQYGhBxI/UlUzef3g5vSeDRbNAVECdq
NL/vO0TDLX+l02UrsvSjDEaio8R8yEb77qPMMjDfaLzIVGkzVI2ZpuXuozPYZTDG
UxbaaR5F40QI5xBSDSGBMoB/CXjhHsjtstV4d8KbDhtQd27v6b4zXbBrE73M8gZd
LyXhor38gTf4zyT7UDCp2vhA2GvHH28JqZVu8OGQyFBLtRcFLnNrIWY5c0j5Dxvb
jXcpTBz/s6YnXDgLtkaPczBfS8S1QblNEzciOFKJjJaxjM/Ajq+DvtU+09+/4jNT
xzxI+IWWT3mRbWKi1AYeDxio2dlZmTyY7iLwHAMUV2VvGFIV4CGcjPoUa2TvXz1b
A7Bq9mbs5dRUM7d1xzPbBVviEpbdIdA/JFHPeknT+aG9KltFl1A1+glk8umVhfcT
CuaAwSb6h/iklxPvywatR43YVVcC2wkICSmZ0pTkxi088p1nX56+jAElft4w627L
vf6+kqLnoewPwK0GlTgok6zANUzWQgK6ikWsdvmS6DhhxktskmRS6JJT1F40jgZn
e7HTz2pQmiLyMXLiW20Z0RvD0tj84UtJrgpNdTk8UbGQSZHv5SrUAg0ozavXLlaq
dnrpktGHtupRjMAt1BGXT0pqTS5WwS1wwLTEgx4H4MO3jLorXRVXhB7K80iJVpnb
t+xBphVjGlGqCi+4IU+H6+0cFlLlAI0qmPVZrpEd9ZV5xrMWq/iXRB/JqLjrVX46
ReQeRuOE0QRaIXwH0O7MV3kkFVPzJatCxL+SW82vHW+rNYi7PE0M1OGjarvC/6QU
48Ie9DXFg1quGCXzPc1PtWRln+scJpeKExa64hDHicJ9SNLhBtocqWS2opTbPbQ7
RjtSinei7dMwn2mTFVwWbnHkM2bmj7ua/rUfcgWp+hZ06HC4D1RvVqzL+98ZQpNG
wjWLjy8r+LKT65oSp3XmaU/Ua5vI7jhntFeR+C1BBgQ3kl4q3dAZRVNfJus669gR
oZ9lUZUQXdbHL529tlSqa5BOz687RdXv8PVUjTBIIfcsKikrt0Dh0JLN/v5OBGtB
4a+cPVe5ZYS+9HdogD6QnupVo24UBiJCFczJD0saCX+biqo05siDNHEYeniD5Ake
b91wGkJ45uPFETrAKt3yFWpYsxhkoWUx+hUdw8bLsh8jMjxi9t5dWeKjztoZY3nR
3RDOQbBOYIyI1DKTXRy+WOGhs8txMtQOdguwpyevqCZvU30/evbOv8jcC7hP8Fw4
LvbvQeqNbyjjakz2wyJoBz93Ni/XU05cohqMzDHXFGCFW5Le5+mlvcN//VVbX+3x
0V+uh8gkwbhiW7d4Ev3oouKQ+SBmBVtRPXRFhteGn+QsZF4xvczw7wx27Uc5BJI8
sgZ9AWR7xum34uD4hMupnasmZhbG6XYmXDu9yetiXEOUU4peZRjJpOj7KeLwavdi
QP4/s5Wd2+uJQEMH4rXrhz/Drz0/7CkrD1t05yOatiWngcwgQhmYKmSSblQI+sga
3sO+e3b3j9DybbcGVfGFrdgL4o5YTJgX+zXqtp8PIB3B3n/iM8iVSVs6mp91fRww
L4n//06bmaG7rh+//+Luk1LVMJhcyhngQSq5Jfe35ECDULoKnXNxRXiTAx08jJ11
ddRXWPI9WxI4thbvpRpdnFDgHbAFnCY5+ENRTK8q815VLLalK7Ccw2NtjdAhwXVa
ALr9dBwZlFTCebtlbmLOxpYyzx9kpATpoi26uNt4NGNHlL5Y/JX9HsUkSyLwkRmb
PNHZ7WnCwGQP8quZXISwlBqKy033uudkwZZoSCmzYtTDWPYWmh4vyfwu3I38qyT8
gKNqWWXnh3E4zfjoT6d0Z1NSzfmHobzJW59C0/nGhZWedsuHxKMIsMIFn6djpVqf
S0fe8Kv0Ag0JxPNA3CB9dLNzyHmBoSf4tv3pgFXt2sh7S8JGpeSuqDBFY1PVdT9t
wMggFaprGmIgPJH0v33tTV+c5V3d6onFMj49W4HJWnWyk3rjidZZiqsTNxIBQKqJ
inJYGM6qgOA7uNfLnnTWrFeJZWSGLl/l7cIRKbwANTDubMCAZM6KP523JBkQTg9Z
bw0XRu9W+5wnKxc7k8+9dfgGf4RlR1+zw49gNyGr9vOtnTI8y0ZKVg5SSh1hm7y0
3PSHxXvJLiwp/IGeA/NUUvDbwiuWrZDvsCiaBQ3Lvc7jmaPYR7t1zkoPWAtxOLu0
3iFrVW/ICIoCoTJxdATFerdZ5/mLtCRk3Hcw5Akmne+g/SnrGRAFmTkbYIOt8htE
jQ1iqLsKmaWPFWx/kjFYwG5iPIMSr8AMsnRsk5gbDefzDD3pn26vA0SnHeUlz5tG
cf87g/SBssDEwb77bm+BwkutTtC8cL7S1BeuO2stUvgtHMwvPM0QDBxH8PZg+L0s
D/2L9Ujy+6kaVKJoPtmWugyP+5cxs5mcsDF/uZI6ccuU20pyusRO9HvjHbVGGBG/
59r2h+ost98NtkUL7tihzg1roF+Yis0ybHlaYPgGCFCWg5ACnO9yd5kbUnQS30Qd
ceJa/FcTjxNvP51GI5JyqQhXtMOTacV0kXceC+zVbrBZ6Enmk5hUm9ntvRTTkcvx
rtzRcLFpusoSxUShsRdG1YpGqC+A1YcrIPFyYI4fzeM3YFt2CliaXrkK49KscNTH
HbRu88GPyR4snG+DtVqEL/ZAwA5QasQoLVZkKCN+hKjO8eFgLpUH4MJtxgUz9N96
+JMgwzmhT0mos0xU5UTH3DJjlzkcq7SVMThXTDedwqiuts+ZLTAv7xlhMbuXZktm
cjFoe9bGhpzABRABdjkdrRYIEtSD7DkcEDX8S0v+xBI5AU//Z2WOF4AwsDoHzqMd
rlx9fZQtpmBxS3YkF/58qt6NarZcDB/loKxJF2Rbi3qdsJ/+10sr1i5+XwfQ84ui
550xruYgLaGuXMrHSaUbhAteisbXn4qifQsCzj25je2uN1J/gNXBR+URphv2DlMK
JReoYoJ2sReGMPuUDRD1DvPGpy9qLjF33/qMTfTOU+Pmu8p6eCVY3jm2lXsdcxVi
bLAIV0/yQlDqrResaiWoGIwSgzB2kMIgQd3OxmWT4SZpxnjsNYuY4ucVIk/UMjTj
l0K15ZzyMsvKfdoe0bK0XCRvxP6+3DUG34msJLPAHhzAZPiq1lJ1imLNXD1/8qhi
7bbocecBinfJTu3yh8inuOYEn9k1hjQPalIkhybSWrngyZeyiWKt1MztWuDhJZy5
AJ+p8MaY5Hy3KIAdxhlK32bzuY7ucwWwEwHlA3hj5E3Bmkfaxp2U4eERUYm21UDn
MwKhjnFQBqaWSsnP//UXUK8kK8CyX7MJVFGVoIk95jmleEktdl6gHMhCifh+Agwd
5ffbxntcoY3dDj6JycSGQ/ZFdgEG4fCyvt4iptE/L1KldAY2JVtYItzpBpq9atLM
JSqql9qtQo1hla6giPFnm3VWiESQMybPQyrShrtTxnUZz5DBDqKPBj8MLQtkg6H8
CavkmJFJXCkXEs3+ADk0LXSjGQeoL+jraCtgOExsXVyHzbeysyzFff4OKhGL39wI
3Q0gzMDcK3jL/rxOP967V1BOkOEeLKn8zfcuaqcJ500IxVCvq+ichwiO2qxzMtLh
JpRj8Vv0A+xr/SdVlb6S/iiD1vsAvupHHt/GBJHoWa3gOh5ELswnxFFbohWb5PPw
C4LBYJ7/a2IOQB+5oYz/g27mkjSBDQialQU8RyaZCZs16ct/Vx2tHZbte9KDg7vv
e3jDm3eaGePHcdx1Ku4SZXDDDtrbLZO8tf6KLi4u36tECP9Dxqq42rQeRxy1tthQ
5roJKpzMVIAjLUPJa9cZcNfJp1xvLKJFHbDKxJxrD4JjlNm+er5IpPb1fbCHh7pO
oqLqXf5CUKBEkW1LFRf4iPM+qoBZCW1uutKixjanp/TJYjecitlAvWwPPRrnrBS+
aBH7Alhc1R+1sY0/Jrnub9dk33q1UcysiSTb9DLZjTlaTRJjWPsqf3EYUAdGmZs0
mXsAz5uXiMnq6YL0eUwFD/YBdYx8vtAQmtZP91LIIQcHYpRoe7jnTG+/YOXcq1HD
mkxjskDgR5VGfARn43dW6VuJui3/eiu9BOr+oGHl6LIcjEEJs7cBsbzi9JpleH2w
A2/S0aetJd5GM+M60ZKCOMTOmswM0QCFQYHtVm4NbOK7P4uHz7YTRE+7Syna1QxZ
VTC0HSS1p4ce504dsCv9CU3YPeJor2TAMVK6SPH59s+WSCAjfG2blTix0mWu05/1
Ff1BUdNbkOCokF7FnxzbfowXL4TVSsUjTRjG9fi673Prl91s3Xf1b0G7RxQlXSmC
mzxmbPNDuIGNFdz3ZcWCuGdw+jC0zY03nxdRLJoQ7v1sIEg6T+H4yp1OiDRlRrgk
CesdGLtCJfv8aGYz4Q9NBsupPjhW5lgh+bsG04yGt1KZqcX5FOAZ2cs/DIR24Mzi
93S8gtZOoRjOA7/00zXA6Gweh587Yycer86uQQ/hNxqgvYoPNCFm2ZgfBlaivNG+
KpH+aZcrj6REBDNVoRDv//9y31Og1rgHcEaYwDhTAFjCvxI1JHQGVyTU2CpCF6rn
SVARcBdsy/ZYn5UVC+MnLg==
`protect END_PROTECTED
