`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgOP1+hJqvnUZf+/YoHaV1TaQJXwwMP6zDwl7Q3+fL2mmgrHzAPdfLU+W89nelPt
U6XbB++Q846nEaHqsxVIuaZjHUq/vG/z6YQahphcdzHXAbutBooNsmCsU+c1q05a
cGh21P84zEJdvjBjfv76mCGSPXeGRROAB7oizIBrLR6TqReeumPJjbsnLdU1Ztzt
oxzEkDwhSesS2phP5U4InPsHI+wDkJmt3ujt4ZxB3Ai2CNY17QrQBnH9JfgCSn/d
TY5kaPtDQwUBNlNAzCB5LIMjAydLkOkF4nwvcDsPmyT/s32MpJO60p4igjRbtuR/
D8WGhsD9sHq4i4MQ0stT2/PkHcSZqg0HpvnhxEOuEQd274kR/ROFWVY631oQ26I9
G8CFc5g6vBj45sdlquOnkmNRK9cqniQXqJH0M0qf7s5LfhCIggLSY3NqqDiSiDZp
qGtsCKBxanzKdF43b0lDIIBPSpS7dc5qjn+kT4hxQYr3xeB/ZuKwMvynxi4Vwe7F
St70IMmRewc4FInoQrjT1nlV1uf3PkHWUvUrsSHLzBaNd5hDC72Jwraec+WWab41
RGM7NeKVhgTUlPxSsVZia8URQUKlyOgURWezgwmvBR3ePJ3tWBuop98kloKPp4sK
aM5TE9yfGeUj6vy/VSFtKlNW/itbQlcm+9m5WTsCe0dsai4Qet9BG2p4wASp//9B
CdryE4UU4NwpgJUkx08sdYZWyH7e15gUyqPrhbfmbpaGLG1mbtUeJ64/rINsYqZ4
d5tlxyBZo7fE4GKDgUND6ML3NFzZoZkyF38oo760zHt7Hnn6fCxfff6sVR6w85tp
1yAGhLjFW2JWax25U99MYZZtpijlf4iE7NKRUHkWrunJkK6Pg8L7eCOAI4CWlX96
MizlskzOHp4AXT6tw+Nbtd4+Sk/gBYFYxNKST5zH4h2CVYP0dDnxvOEpdwNRam4S
5ULLRkJ51NUF46REcYa6g//pkD0xrN0DpE4yZd5iyxwTG67XL23unBrrGZcq1oI5
aMkSWMLL+8h4OZsdh66jsSzDcKE5AacDg7dBRnNU8PMvhz8zuEySi9LN147Y4Nxq
beORF+9/1UY1b8yMQcCvaHmbBsCmYoHvbU+r3iXxinTI6TqTXi14oIjCbQLmUChV
4+22CZxrXUTxcwxZYjtis5Bqng3fpWHeZ/1j7zvcvAB3MN/yjD7Ik7AUUR8SkmXp
cQQNwD7fh73R8NqbzZz4QkN+vWq5+kEz5wlTW2eG5V3AdOCsn57Pj6qoKrAcrCQI
vjiUXHQjjo/gP/ioSdjaP9ER6swd3sB3nn7oFpEI9sczTYXrVxfSJbaz09HoN1Ls
LPWyv1a6vmESIJR6ECWxxLQLvqNJE3+UeEBI5O9t4g0LsHTjmlrRn2UaHKX/VEeW
vnCqpNAe5mVJmHWXKBCXK4NGfWiIhgw8pdGyDkYi262uApx0V13KvdncRWN9H/AD
r/51fZkLhoJhCDmm6LP7byu12ADHWkOAF5cAJfTpOOpBloPvtU16sS3VmXql3ICV
3C4oHxRKsRqxNTPp2Y+I4B1VrabwUiIpxBpQH9xH3iA32H4s1SJQPRqEroPu9MMR
7p3ERvxohkq3J2FOMSIImlEhCpOUX1FGnunrgHG+sbHPwYBiZ4bDFYODQz7Wh+uh
EyRuSf1mK7Sb7DY176UmDS6Z65nKuaTV43kntwu355fk4Of/oHaus6kANygFx+yY
izZj+4vJXZcT8vnIUAPv10Cu7X2Iak2i3VZfdnkXuZ1WGW3/RDl66MXsrlGwNokY
4CsW3kUH0HKYvhbGkruBSqXnt1bVbTE/oB9BS2du5/0rTffphMrv9mjESK5bb9Aq
kjKZhrt5895rpy1KpfxvQs+5w9LUW721SmXtu3KDQwYSCWrT6HEUxCr/2x4ma19F
fK7Hv2l4RphHsQ/4jZpFC2RFXRJTGo4sayYXWsS8kG7y3FkLvLM/F77DbSj/w8hd
FmpRQyftqpKL6a6udRprzYvKh+Ama55X8i0BG8inwJfY58BQURJkotRAkFaoRL8s
izWAt9EWY/JcuVk2FJ0tMNibNlO4q1bREOblqWQgaWawM9X0u+mOaOVRy7bjFBS6
w1QD/nXQcketCH0yKRg2glmLFERO8spnm61LaA8CjJnJxxr6Fvc1h39wk1XozR3t
lyhQFm0CfSTAH7ifS+qPRxn6BOYkNV+uZao7L/r/NJ4ocvN8512GBU8UH/12qC86
NCv13QXdS8jTTbSunXPD55oRbgijK66WXzNDDf1Lw83+9WujSiE6LaXWxPQPcpWZ
2C6wVEv5bPe/YC1XfKlTAyQnk9JxOJesUi2Czk+tK3CXpCdD6VfWqd2EeXB/SL7e
YPj8I9hjglTRgj8m4cg57ShNxFH5lsHxdzBgz743uw0HYHP+37Mfu7yxoMZVc99H
yN6zSJfStuPf79BbX2hI0VM2cXxjYN/LZBpTewru1tbe89C5B9S9Q8MC7QdJEqv1
nRMtTKwJMJvqHrSRAKqFgg5fMFEr3BiqWu96QG8dJQTYmZTo3t/ShsqGY/+OC9a+
M8nI4hTG9Cz6ZJ4Z59XJ87SkFCcOqP8z3Upj8C5mguJe3c7oaLHnzp8WPdTysJG7
T6QAMzhw2gjmjbykULaUvOyaj9K0bx/zbTsds+SwknQg6CyA2sdpaI6e0vKWAwlP
qZc7Be3Ge56usBzXKHuyWju1jULwwQ1lpUmqiCHWE6ZWcCfZidcNns70bdZYrbbr
sdMU5M6oq0nAh39FkCaB5BTyuITBYKtY+R26eC9cgCZkWT0Op/7yH+rLyhV1w1+P
tDfw3XQmmHmOsvZUQ7YpSQMxB9d2yd5vKxt61Mc3R6GeQtAqc8vFBqwAPAu8JDTX
pVJOvBo5h7+X5eRd6IARSVEQdBa7CZmEoD1DLjIwzj7Z6antKTFQKfk/5DfGqSaW
R8qgLTomzp2c85B5H5B2j80WKQBS3RozLKhOSWyaa+Der/bimYpEW8rwHAndL+tG
2nBCZvbcOzhZwY4DEZbX/8OfE3+IwRAQu68z2z0eLWHjCgNOzRXp2kXbMivpQZx9
YGLuEgzgMfTj+G6U2/0xBNugp4rHqvVti2Tobvljo3znpRKh03PuwrhOs9c39VjA
U/QMVgHmDgCZOGQcPFlfotVj3FFVEjzqVMEe2gm9hrio6gEeJ+QeNzJTfk0D939U
8VfbQY0LJdKJmnPZj0/unHXZ1zU8wxXBExY5EQh7Mh6/PcM1lNeETwXvMXlhLJKh
ptks1V65A81YgXRHRL2raehZty3XpdvNhQz7WX2IFMQHdNVfQEM4SQ5AW5cRz8le
OQGy8yrJq27UQviXDkjXwNbIgBjzQ9aAJscAWmGY1qthRTfEAEI7BEPyG7g80eQo
YjjjoSOv9DZDeLHHm6sYspC8z/pIGnjnMubMekHWi/VO+OuX7Fv0Grlhq+SJC2wZ
64S2dEPzQDlf4gWYO/67/OeTzR2dVRgIsdyb6WE3faYAKIo0biMMgSYw+lgtrLro
P47AMpo4Bj/4bptRMuDoWCGp8tWbS3WWyQ41cVqP8uEVbSFxJ6tl8zxI5fHon18j
XKR3jfMLFpo2guCN6610TG65kb46vOXu87TJOWZbH2zsM+3gqSilhahp8XX+yfEZ
7jHEhjbDeTG389W49fxsqqkEseHow+t8/3ggTIbibCZgY3qBUwLpdCztn3Jhqk/u
ZqZMqL2k7KM07k8HlHZ6QKKc3U7i8yaeb26TW4OVI11/zcTanZR1OIsHLiQBBNAx
gEaENWOv79Vc6WWgVEIVX9lkLhLbR/BkidI7sGSssVggc7x6cIPWb2G9dzqzQA7/
vhcqU7Di9ljs4eedjPB6mtKNwpq6tKOK3ArW9IFK2WzRT8tFZyjznXx5gr/aKOZr
7dxlmDhgGh1V2aoPKL81EiSXPRMJPoLVZe5IE6Fjq1CnyV9Q43W+4DFIGsSLHKMs
NXuDOanORmVb+0vC5LaxjNwaQPQM7uXzwewh9fQOz9pRRyqlnyiRQnKMQpg8MF10
R/DPt0nUuI/Y0kRTrgCCw4guHYjA4rHSKcjvAfc1Zb+zJlsMKe/IEn55d5jBUO2L
iTjwyO6TLCH/TDITAZ2cVqWCsFC8mLizuz8GwDFgzy1FgxsQ+xyWTh3Htrme1UCr
3+3KvmZ+/AxMa9ywP9F2tlpEM2dXwnu+i2LD8jbjJ2nZj96+TG1MQyiIzvwHTr2s
nzOfabLHlEadnA7/73BuzWV+VratkbB8n0CzJD7crCoGL0XmZBrQB3JNjC1HRaEC
EX5B+wab7i9zO/wKrit+99VqCe29gOVa3BJWfiXh28Sr9xar5RBrahPNeK6+wJra
9QowJVfMf0BGY+JP15apHo74gPNb+XqMpm7ClF8Xqj58TQnitl9yVpp/gMiDsu9F
1Lry3/EgY4q7/TRP63Joc9T3MI1pMvxxfIxUc/mzxAdz4hg3hQgDlBL+BgZR2rEc
6HvAyPvEBmIRoBD1VOySfKbkRmIotqvZVLhsfNmuOpv+RIEfeRz9aoAR5/RL5bZF
YnA4IadsL1Jpzvf77Lrb1PLPv2LNvrp0NhS0B/swSedcdHzQleuvOXAi7SnMrOBm
I/D5D7Jq3bnL04n40JXsVp2Lq5PiqWHz1CRIig3nTw909FKRs5bpOlNlPXD8fHt+
xSV6X0RAO3ml+eV3yvBBlbLmmVNbVQLvwzoeRUedOpMJG9ncJLKf8LrlgZQRaMpl
j8PeakzITYhxqEIGsOIOiNqozNENLAeFmyrKoqNQuUjbzGIJ15aVqaWubgrqOU6o
8rGTpnbnu9cgiykgKd+L1f5K6FpiWLkP7jKXioap63MQTWVGFt2Q1qzmIvZWMwx3
orRQrhv62i3AUcojYdlQbmBATJ/hhGXrxs4iZQhovJdVpHEd8iqiUxuHp82Aufqa
7yCM9vCp6Mc9VFRKJXiH0adcVIsw+xcRH/l1T8UQ18WjfsQyv1orT3Tq1DEgfYGx
3I1pF2QXC0sTOLuIHtnPq+a3DOcqcvi8t99zzgsSdNSmQII5oqq1FAD5vhgGwFaM
6h0xofkAWO6hICLsXXxky5Y8tuTAVLra/d/AR39fd91B2x6qfV7aAPLcjSMdaaBP
i4+AVPgrQ4Ze+viPyuXwonlQ9wbzC6d46CAEK1gFAROb4e9czgUemawCBMibmsOq
bnJ9RQ5aETlU/WfbUW4iMERSA++CIm0eq7moeVNIZxZtG68QYOdbFeWtP99RkdaG
07N/lMALSRx+LKpGhBVGeFRO5DEgpBsals61StNu6czvzxCWfO68qZr58Sd3UY4t
rF1kv+j1aDkQI0cTP7N58D+dnBtzZkk/GYFWFaAwIJ9F/z6e2YcQou+btrozCzOG
+hWT/LP/UkEX5Wv85BZlkL6WlMgDYb0rx0Z/vCEBAPFDR8y+BAyuWHsxffhlGi6I
BH3me6Xb2bdNo6OTdqigD5rUId0j6hzOlmlEptgW01B2ecZboZ/Uw/hgQfhHzx+Y
Hnwrxq3Y9vJL/NEGdFWBgU2dHDzqhzUrkdCk0I4Ei8I54YjdQVeOH1jpwNHar65t
TQDBd85MzIW+S5cBI/0vq2GvGs4rERO+6kYchGeEmarEbnMVmvhECHP1X8suFHsU
LkGvlkLt6fQBLUE2wiOKFiPlVvPJOirDqwJRAWg5NZoeX2NGbdxZpOBCZZO8OERu
RxGqGHp/+T7bskblkGGEeqfFgSpQP4mThxp0ML9wt7ZcnAodgt4y38D+8FQD4KdV
c2hidfuHOmazMpF3RqpEXbhOWrh2S7jfjjC8teDVteru81ByXwqN6l+go0Mx6tVY
U9TgtBHCrQEdrnJfVfMf9OvN8kIIr3v8Q+BCFgFYrPhWwUD6eZ3VmpkOmg5f5iUl
nIpwrf63IeqDevGbKkHEGFadLyf1eGiVrtumBKZZFvne1Z3d2ZL5gbyp8Lg0Iog2
pU7DihVuwf1gdgtUhLNvBHCSvf7JxhE1GLiNT00cRFRUDvV10MBww9qPYuXZnCUg
ELuMT4HRKFPixmv4yUYLBLvs/vo0HatZ5gsXXHLCaPkT1J/7b1cjG9GFD/d8SqJO
WTdZrnDe/jW3Uc8WO65ahJPpJr9qp8jzahexDGLmng5cMCXafw5JnxkEPMpVXjAu
cn5wR3R5lRs1dzfS8bc9URfHZcTJRx3Dm/xfyKmid6w6FdX6f9jb4qUcxKAgoZiy
hfz8ogWEhpLg6/FbKeeVPYEBLOAF1VK9ND3jaIoy0c6DCv45TNVpkhxXu1nmOgnl
xGBE9fbIAUT8ItYfFFh1de2P/Wpn/z0zUApAUV8HGo+hRpXnNR+FvS9B5xFqE4RO
hoSm8WV+UCgvhUYBfKc/uy5W7HeltGnL773whtwNRoNFctAz5MkD3CVzMX7fZ19T
rYjfnEznXF0f4yHrxrI4MMIid67jFC18XoyFpOGij7v/DqH/HiQi7o2pcZzhIfod
5Kiv2mZpaGLsdp7yVcahAjvHfK1dc2VH63vC/dmuVrTkxOm3EqMxTlAxPg6ezF9S
8TYLfsrF/CiTTdFgiETLJsv9bAks+duV+TaUwd1ox79CXlg6MNof4EjyE8S7iZnR
6s5/uZ3AHWOujBhvWq2F0yE18BFRuddUArF7+x2mc6VHKgfj3fC0rrR8Wr2244W2
bt+Rv1VHVjJLXjyJnIa3EPRhI0Nf6PbMH6hzPHR6SdAYSr91FPGQ1PStT09z9N5h
ONSd5ouC3UkUdoLCGc35wUwQ0mbjKJImVy8Tfj/lAYBa9nWYlm8MMkh58DcdqS0+
S7/O5GLZFUanfJ/NvFbthdDx/Zlaq7VvwbbRYmhRDBBC45ArdPZS8ehEy3NfIorQ
L43EjhN4Za0vogXHMIhr9IH/36mrGLv+/nzr/4RjM31nbQMwrDlM5ujbzkyxOKjF
/RL+JCfo491qHnXd8QFsWcczM7AghMac8y2x8LHhUtn/Skh7mp7Xx6qrFP5ou3z/
IGF9OADh6kQhskiuQ82e+fE/vdXDR1hRyoruMHAgKUTM67d6qCoGkcxnbc0LE1aj
svEVyYwYpsJ2M9HRdUp0MfUdqlwZSEKqKJCo0XHUrIvPVP7SXrO1pyiJ9bp6mb9+
bw/GEbHgPj9aG48cfpr1+rS/H2pWE4xSWFAVMVax6i4t9Uh9W00jjcVJrzcvXCxV
xAnaTlsJjhsXMb4xL3gHR4FqAKchZw/NIfCHZ4iR+s5asxcxcdDtw0RoDKPWfEHn
6jFji8jZvmp7xSvv51/+4YFz8Spo8U7Hb/syJw/5+4OrG1I6LK32cbXOsJid4NYB
u2XTe5X1HT7w2tgXIH6Kop9AzhDjqTXsTTjGYORNwTSkBQ9ncp0p4N8YPAEJxzOB
MWe7VUqiw31oS9LYYqpCZiaUVbvTLM9pz7offSfQgT6M0BzANuvb/A34tvujq/IQ
kbyE5zNhp4kPZbA4gnPk4aDH/9j29jP+AqnJeny9uGETNBlzU2aVsMPtYHgn3PJy
YwN70yCo4vHvdKgPatRB6W/iqX5lgLT7PP6LGBuYVe1oHFc0YxHlmACTmjcKCdIa
8WylYvjBqVpj/WkpoOkRuaDRR2XfNpCXY3uD7dyZ/ytKRCPT9ugVJbGNugh+KfmU
tv/s8hlgJlQViWQRLdyLgBjeK4eDeiwWC0pALNJA5XLdFQvhFWL33UC+PjPa2+Nv
zuMaGRDBhfL7P3LcwUzuPisQ8j0zLyBrdhqo3ztLJFJymtyHGTDtCXkxDmaHlmv5
GPBtRd/kjCzd9XbwfVb6Lg0xBaBm0hV0E+ZDBx1bE+9RRzxKahBqGvxcoOwyF0VW
pPEERWbamNhnZpH4KdyDU8iamoTzOMh/WkBJ8Ndxd4Cre3hSWT/wvCWkhlxRYNFZ
eB6ljA5BFvGeM9RjYozuEOliEGWHcgV06GbVf0i5/dTxmmYQZm7K39I+zVh9VKW3
/Y7UowNfWnHRIIBcmtJz1MyoP/wZacLrGlhWOduSV7VjSdro5tieNKy+ZV0BGWgB
MCfcO1gMLH0o6i9DDdUADkbLBeM2yBZ3jaRprTuTHGiTxgu8Btsmd0pBki3dxZci
KY2J4LzmOGL8k+utOmamWIigCHjUUe0IJIU0TfC2xATRwJbUs32a35SwozMAdE+2
hpLn8b+ufnTw19Ew733UtBbArK01mqBCf2609MadHRAXStNSc4Cp3P16xLVIsJQi
YFHdQgREQqg0A8y6QNE9yC3QsEhShixPnxtlS9+hxpzbq23anDacYcm6v71tlpz/
iCbQzzFCOB9ABC05QbAF6QIg9g+VOm0FV6Q4iXt4tVN/+Vvrf7PAI9ugcj95eMps
o/AYmbaRSuCfCOXamoiDW+9zSQ0V2htfBcpMzk/CngW65BwKSxNoC1jFHTV/9Ieg
6r1ZOTRF6XED4lloD7hS4WpqOXxuItPZtPQKQVNgu2+yNyU/+GdPtSyTTpMBbxb+
jHwYP6h4c0kuuGhcoX+rOrBL9Hf2cD4kh2IQ7nW48e7/rweVmBpRCbn9DsvZhhK1
eg8nb3ZU4QrhGEZzGobQyXWx+/w5qU3ridNxceVBN+OGeVNZ6eQ0qKP2lLUvHvGp
8UoBNKJQuTdGzee3yH8RSXVJRcZntyMsSVzEQJnwS1N0pMpy+sIvHOb15GY6ht+f
p4ejCOPU0L5vHXfqFbmelfoSEr22+sECIDyFDdbejy6m+TrLIxNipDY5eU7YtoeS
Ub9HwDSFwfxDE7gAYWmaKLdbuVRZVwG1oGKwSzkh5c6D+sk3N9g9djzdVHMO2n/0
VmxeZoRN2LW3O7kOK5/a7JyzIVvpmIYGscjSHRNZ2i5gnKqdzSvDRu//9yv1u8Ci
veujWP/FPb/ws1veVJ2AEmy1lvziSPvJvojDA/S5nh+ECD36tkI4AZxvZZI0kQK4
rtTUsqt84RY1PCooXP2GywM2itrjMlaTzv0cq9pLzEclS8/b6wCe0hTncCHtwLN7
M1VgareTEq/FdhYQi94A48MkpBklqwDAPkIwyKSxzT+29l6+xku8lV64hlW9QJQV
wvABIa7LNjaNFhxta4wceboSHwtqaLKeELAe/6yj8XFVNJxJnyvp2BQrBHHFlkWZ
xv47rGqD6VbhCn7aWtCnnRhrUoLUkHsVniHzvADrBXKo9mChHr3G/MorkiITRvJ0
XVQn7XS7+v0nObbDPJGSlTU2V6C1mngR37mgkdAuw8T228AJ0hrZyolM7jFSUtfx
adspP6cTiIjDn3xdnf+lzw4FKE/5iHbcZbYbu6mWTzZ0+VHC3I3i6QTHN2jG3oG3
yqXix9GWeCoZfAPZoVzWRBAlveDWTkk09jiyXaSKHQAYmKxsM3DBiX4b58Zsse54
+KQ6tPdZrUmQNB24PO1hZcFWsHgyF3ZOBDbVeWyPd7MCX0OnWMCIPEnWaekLnE4d
Jo5ZUFkymCa5+zN45FJdwrcF+XdUJ+rsQnbdJNvvAb9f+lmuu6mtLHAGtKa/nuUI
RM8N6UpEQl/EibHpev6fVKZEUxxRRAiz6T2EjAM+bqUvWl7dhl0+7M18A+7xOxHi
4W/HbcVDxeABn2Ceuf1JQ18ngZwCAdCBhN4n7lhXFKgbhguXXYqEHMI8kHRKSZ9V
TnpFfLlm43bEJrVCnKp9+F91MVCZEWzyzJY1ErgsRDJL+pHFyL5ua5p7eMmEcMWE
1l0QgJx6k0xFqC3Pzgy4baMmxbY4YoB0BOnPt+64n4UjZD8na9bklarQUcQ8oBCw
PTTTNvrWaM/t3xoefM16MgeyqyCFGXi0FeNwP8m2s0IUDq8tDz3K/JdYzaNkmSBb
ONtumN6Hl4D49b8M+CwZzE9mwyc5vc9yzFA4BJWOOpmL2APMNpE0D9qyWc6w9ob/
OjD2icHiKT3zJYu7+ruUTGEvbkqlUVDa2MurM4tdFfg/3le8VNS/bgQk0ds9od7b
tYltUTurRKAC59CXqRE86bcVWiMXmqJnjUf+SVEkrJ9nB5FTXqWjfeLi+d7vvo8F
2pulcAehEeumT8rmlTc9svYlIsrO932d8sia3wAB6v2NpEPWQdMM/CTKwRmGFwAa
RH/uI8sMON5fW05FJuRLxNSm/UGn2bCx8ij0A4vhZO8OIZ4IvHRrw6Hy4L+mxpE2
8XMqEDzrEIWx5rbWX9oXgwEotphMG3/53D/6+AsUPCH1ZbAri8XbRSqZV+vXFDtn
BFqc4FTduWpawALLBFzXcj0fyY2RUMewLkNbMz/uXc3hsTkefkySaJE7Y52JaZqj
I5vSLD4RLpMTjuCO8XfUlpTfPGc8ybJdl8NWBfuMFqrmMNARiMZbLw+Si6CP0nJR
shjYuXi+OLsNiWS/PFuyxGqWPr6ZgZYAOZtrDRlrVD49vIVquxxHf11N3SxdoC6Z
N/YInSeXGvogBt8LYumh3DM/d3MRBCIf9BNlawqhtJPWY2/9828nqTeSiEu9gall
e128yxt4CoABeATRYHWnRLXv38zfSJq2kAkKM4Qwf4/9pKH5GGnYz1TAWzOr/WBp
tbqJhzVk1A0XhYq+6Z143CpGDLOd1pLHr2YmvZDjqUNqawiknyTxYAdAUJw3+4oX
+oacqwlru47nBKWbVWUiMFUUvtOZhXiHS0xSYz5FRt/N4lMrDKAeO/I/a5Anfv3P
M8lgub6M09ozAP+mzxPBtLs1TSLXUrq0TwzOBJCmrj64BzV0wNN8GhhwhrqVIHKR
dbAxip4p9kIUKkBbmstnMlgzYJQzizKDBh/gCpaRVI/bxrqaGTahm9bCync3OBpj
WKzcwDKk9GIdr9/mqCEWFLf/s4lXc9muPj64ObxP4LMh47sEREwisbbk1Qgu2hF+
Unu+zwv6aKHB2TazT+SUbN0fUBDKx0gfr7gHuqiNIjz7NSAxZiJr8z7M9MGVasXL
I7B/IadDTRdJEEH6btDNf98qBeHJketxj89ouw5EchKOqgPSmAQD++D4YaT1HfX3
GPPLTrNX2pAvB+zu6iTuBbnc7NBaXgmrrDr5hJnCg5JP2gU9UDsfLIkdCMtxhCGC
NSiWaacsdWyGSOBS1+CE2uX1YPSvqQ7bodsrcvKpKIjhHX4KP1zK4eg5Z8Y/6465
tTHfGOEuk5XjBqkN8Z5uo35Tt5TlzqJuVDm10pzlkt5YEvQN3Z+RV4U4oD8VRyOy
itQN0S+qDtZc6bkzd30F8Rm+wFGUKbTNHz8cRMDF2HxRHj9MprZZ4dSJQdVgUHec
68vjl1HChDcSsi6tF5CuwYENkbZTzjB1dmAIuto3KjS+8kaUzP3wa4ezOTBfZLAO
LGWybmxzn9T1LDqAu1NvHZWCOeTqRbBHA3WHUPpEFmUjFEVKJY0v9htEK3R9K34S
Yc94fzzrqDqrpJtMfLjoPdtVD1IvmSX22Ew24QxU1KIUs9SpolgdhVtNtUFIGf+T
zye57LRfylTCH0Mz+3IHXK3Qs9cv9pTk/urgPa0jfloQUVBfSwtQF1z05oHaxi40
32wou12m0YJFbkwq1BCQVTELX3D0hIPLOB4CzWXnZnJPYaXpsW8AOmOx/MeT0INL
nwLYd+fZOvx4UeIzNVBWJVZSmvYAkwTD2Wxcc/RbW5YxY4d/0o62/JfbEYniWx/n
D2EQWn2g8kX5lIglAdhYHzz3V3SjcJoW00FX91IbS7MbnXhNWqfTjDAx0q7l+Jr3
ctC1IgbohgCzx18dM3K388OMu7lfghhmT4mHli1cau2zWF3qLp8LP9ER0DNNk7i7
+XjBhWuc9DWigkpdJP8ileWKuavOY/XBAsQxMxdzTifPDf9mOnKdCd4oAbEI5kEU
5M427Oswj71GLtOOIptYfL4WSVfk7BW1ExsS96KpSHdFR7Y8W0SMW7rgT5JYQTmg
+VOwx7sDIR0qb/P03W0VRbN2DFu4QT4+HA1Iplxd4GQVWv7EnZPChWzdYFOuTJpS
UdHOQOSdiV4cqSCeaxSxZ8CDPYLuI/4XHoxX7hf1WTLk4at5UnBPYMk6n13VNKzm
BwFBK2IiXvXcKWeIFNBgJO9uBHuvo7yhh5kSnaq1h+D2xaefDubS1t+RJa4EiaPT
FauqIV169prM6AUzoQc9LcH6qKf+g1Qp6MdozRhmi5otPV2/3aRcwA6CfrdooCvF
DHLzE3WJxtc+ylF7UhYDmGjT06PjFRIoKEYfa4cE9CkUR1e0f2x7JivpHF3jl7v7
tm0nfZA7/XbG9dA+2D5wMftFYPlDfuA0FwpAocRLQqMGRhoz6KTUpQTAUf9tmP3D
3LpjmVK59qOeSmcbhgCjI8129xw6066lURFYYt8OuNzx5k9hCCFVuJDPffxRvH6R
ak7zhc8cKtmaMwczLljDwmi6gk3ECIqPPdJ32y6zhAI85L9H1FjwwYZHHOlzmVoY
eS1Vs0E2IcKqlNhprq2iza/b/zwpWBLNscofomYXx+ik31sn4xbEleEadHw2F85D
dxaVvGo6GWKpi27OhByagaQv4QdXsfpFPhOFRblJ/3SlcaJMy7sNvEUOFolYjpXV
K6ltE9OTIKKgFZHGafei+Ln/Lxyr/MGoXfajh4CgXyd1AsON7OUKBpxFys8aM0Dy
L6wbKAn8/zxMn7SLETfa79apZnt/KlttMvMwDwoezU4f8jHBGAYY2S/unFZiG6+f
iSUEgT1O0Myfcc1HSJYu7bY7yJvneISKGOE/kfeDe+ILdIdL0n4MFVrJ6UO/b2ze
GehLI3bAhKbynbS8WxZijszb0BHCP+CAjiyesmy78R6Ww61Vzh/1OkPK4kh0DkDy
8yf5f+H6nB/8nDIMh6+zDDsbgJcn/F3h/xR6FPkxjrsPcoetHZgI5UbYMH1F9lUR
bOTv5qPOmHX/lFAhYCVD406P0XXNLsdXN4/cOeouiZkYV4orEkBzGb0oi8rhawMr
RwVJ/E4Oa5C/vkvkwOd8ovcJ4bKEBUQb+Bk/x0az0ZpZCO+8E/gebJsE/MmrKLm4
dSh6CyLap/WtDdW84h78DhORwxZdOGcFRpxyJLaWzjOqfdt/gQemflyolqPyFum5
p/401zo/RngxZRBH/IH80Bw41kL5EOlKUq4qLYAMtNIi98KINudHhM35dNF5U/dZ
0TOiXPAfBGtYqcYOmJTLzXf6DwmWu/q5Khoen3Pi4ojYdk0dcs+v7hhFvFGBEBv8
EvsPijxRglHeX/afxGk8FOKITKk9aQjRjmnGZgZMZVcPiYtPHOU8cV/eBrLL7Jq7
`protect END_PROTECTED
