`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4cKFEnKPvlUw2ie4exOp1H+To+vBB7fweSVJ8DCcdR7wjGrGup4N8xMlNlB9Y0p
eKm7KHS4Ko7DQEaBsh8Y6jnWIlNL7iOBM7+GX0+IpBWNHqbCHws2OAgJO12CTEgv
ELPgWn/iKuAQD8mR7/z/eACRYkZEoBVkABvWjmBekbxphBCUyNiIHxTnO+zJwYNs
dAhY3MCQB7FGBVwzW+spLXU/pU9ai1CC9J3aOMFxEqaqyZC5t5FQkPJTuX9sCZmE
D+EPvLylGdvLVCisrQbo87HExVOegHVRNkTGSFVIkZB2Q6MmjGv7phQ+kTZLjdeo
Kg1pf+gZ4gw1K2fXYxNaNnkKOiLv6i56eW0AbshmI+g3iaUisOUo/3F/rYZ8sGEk
vkEkAFO+ySItf09Wu8UtuzULr9PMmlj/lVShhWqTAuiI5YQCJ2YXviGkOGwysfdj
`protect END_PROTECTED
