`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/YjrowfC+wP25TD09siwpBzJfwfDI3nrGfCRJnytB9sWJOQyFWHW7J/SinRFOoE
/hNkLF8NXqOaVOFlm3XEY77v/DMPw8BMLca+BxHN5ubJBPCHN98c5j+M9uLuLy3Y
gTXkW+o6ac48Xu0if7ASbCZKItspkJRtPuCzkEjB8ycLolqqxEe+BDEB8YkXvXt4
flTMYUm68o1XOweCpJtSDRMcJUVUYg/eDE6722DpjsLaLmZ3SSizqmduwWYug4fp
X0qyBc3DAkYD53KztL8cq/QS7yTH6oCs6wtVyhOEQGn9hyH77eNFKGpVpa3fB6GO
wDV4JUhVaIEesW+GiQLYjZWHOW0eimr25DPfebw+6fXKokDNq++Mnm3hrKw98Ni1
66PoKX1EB6JZakdZymjPgxJ5VqoUnYHzZ+YMPdlI11GttxX8uVbsxY+WW2v+o/Rf
k5gM1+NcA/QAa19fhy/gdLUwM/0JVeJbYzUw24YGTPlyBN7h0DIToZza5E7t6cyu
5xww6YjAWhijh0hCmRPgiANQE4mNPmyR5+mrOSZcENOo/ON3sl+Jrg4lmHCXD6ET
oHy3IQm80shXZmFoSz4CMxZgP2P+LeRW7isbmPiZvya+1cn7vMCfePOE8MGJbraY
kZBwuF93OO2UZPKZ9Gt/mn38dAhijSRHmyEzLKSAoaXQfGKu2DqtUulr3XZk6+i2
4I8bKywI0RBBT1Ns70EQo081XY+kp3lEniUiSdxCDB2U3CxC7xh6MTgydxFt+Kc3
5TD0tGE8if6qRb1OLUe+FPyArJmaQQjEXv9nPU17yO6LwAg8B8rOdWl85UAMyryy
IM/yZtbcUfD76+GTtorS3e6rwzf+H3We8z5P2tqmds+Znm8Okd7l3Z1V45jloZ9B
jImb1gC4HlCBygmcJ753IoS5WG4LRkBsVMy+keHO9Ciwwl6ncYYStoFB1lXYmY9N
CboGQfvahYe4ZkY9oT/3QCvF1PUyXBDvZ8tfcCyZIJLlWXhBKAHclQaBaaJIFg4+
l6GPrvU/5FBjxOPW9B1F6wpwP7su4b5KrGdAspQgM1uGis3CwltQlhNw0uGCFzG4
9eTOTIVJ0siz7n0XNt0etYKxbbHqAOIkoEElWWsh1fKUKYfaxP38fOXj0zxNyxKp
gIx7R8L7XDpERJM9KL8tHfpvhbojQeEModq6ql8SScTEhprm+S1H3xzx6C86CE/p
6Ec6R9P9wbZvrx3HPqTl57xjfYSdE4fv+aekISw7jptJ6+JtLX4p0bbNT0Cr4kka
QdD2HCREDqSlR1zGBpDfTqE16Q/IoiPIsKwQn/f5KELpEe5oVbHTp1nCP4rmNThd
EIA0xjpIjOcr3g6CteEmfpGV2zLr/s64Q9jV7nRs8E9zxlFhBnpyojG56dVmz9q6
tWVA/fSgRNAPXIPbrDOlJlVQLFj15s3yQgikdYAnsbaYsKacU6CnEiNq6Xa8OS4q
snjnH4y6Q4Uwcb6qi8s2RwN/QuBY1xVLlc++Tbgzy5Yz2KaQVXVNcr0KfDcDnejq
LyDgrAXGFO/z4P2Gx2h2UU9HYQk+YE88Udg4LxjMl7iipyd/JE6nm+vYuoMmblNQ
KoeD/Ht8/jwASiIrggBfiK2gecE2bQD0Aa2GKUFSAA39kyEOCXI8mVoxcviqVJjn
4HtkDt6OooliXuXAEEdcJhiyFtVEbWiDobtSCnn7Fbr/Jal1x15EoGWiwCrq4L5B
0+0UrOYsogTQaQT57wxVdTnUw379wLA46s7609SZSj0CdAY8jvKTU8IDVXcLkei9
jy4/YK0izh9e62X5P3pE+yRsc8/n8Xb5kWhM08fvJjR3SXQEUu7NgpZ03G1QQNvm
wc4fO6K3t4E5dAyxFo4MD+O+JLXayv8T46Sz1NAIDShvAiau9KCLEyZkvTHyraI2
Gpncs30uZ0zFdVaxaf+JQxaZKIClsg+whg6QlRQRlD0aOm1fBIZIiKzt96iQ7flh
wGcGB/DG+4Efr42RJGXUV+OLi5cYkN7czzjSBvqogJg3XBbHssOR8VhpQFHmQ83P
2F4Adiixb00lxCK5ymizPm55ax36NoXk2HprcYXeiV5zSwOPbwDSG2/iVzgVCJ8Z
XaVllEoahpB82JujS+ZRBDrhCp44uJYKmpBTqHekmflHftJOCvGIFEtDhzSWb6a2
bkN/Ho40xXqqfGmxOQcxmEjkb06P/iAPlYOY1cOOPR4W/b4BLLxX5y65wgbTLWuy
SovNbjpNZ4DIO+cHyMztjs7tcGbwQAYdUYVZHb85hs9xvN+Iqloodn5PC3rx1pV3
Ew72MIdKjySokQu4VKg87/icKKWxFHPUR1YoNvbIQrB2EmcOnS6pJQVTjvV33Vza
+UBeTbhCzTjSoh8BQPJYesZONomnOWLMcve22c5NsP10yephgP1aDJEqmTtC9WUg
Cug7Qg94+e72I68gz0/1gv99SvjSHaR35ro+8LIHk/1w+EPq/zXdTufHQzxJlwED
/9rl4joqNWDYS7ks2uRsAV8TTFoH9sduIg1kcSHIG06760qgFSwSXp99q7cMKv3T
f3eVYFdMVItXvyQykVz9yGBFLglhnKKRKGCj6Xg/5814ZpDCc0gYnFDy4q6lXlJH
m/pBXRdBQKASdGAzoVMvaqr8P8gJi+iyPNHFIpSlzlTyUinWPFl5CjXP0H1EuR83
j93ZVqFElStvwNmsy5SNKFKMFy2vZyhfG3kaDBU1KHllCmq26O8Ws1UvkQt961lN
sHQE6nyX6JZ2lFRTEH8CIkzijpuPOA9ykpzVu4EBjHFhJL+4rj/ISpvAA9OBzqWl
UUd3NB1rorlUpxDNewXHFZPXXvNN5LvTvq1+osuNkXonZgLDd9aq21Li9Rz+M6mQ
gC+yQ24+Wbk4VfcKM+wBsBuLrjNYE1VcAhHa8pTDfX+SYC5FS1Cuiu3ydqrt42L+
eY5b8dw4BdJuGU68Xl5td71ajOTgbcye8KQCvFUlld9fB+geKYIOW7WfPRFt5AaV
Swn0Y3A569nN+j1Vd5TWKQjo9oPzcmZorbMQQ+eUaE8zFDkEwm5m6gA8CiJ/ZGCH
AvOx4stpPcppUS5/D1zUdNR235gLyvX7KpUPa3MCC+hh0lCwkbfR1445HSiVbIBM
ubnYkSVAGodaE44fFVcCPzS0gx+OTf+cZXTLq74NCaisGvZDkNkixXiHM6C1fqL+
Z4o94bT6pHZhcP/uBiCVZnEBCyqoNsfA4tdmryP/TUrDe3psD3TW8QZcceuYCosO
3KfgaqzwGiGClALUmelExRSmkpmjDjkKKdVStbQlzSBIuAyAVP8jkI/ruUF/njDi
8+0k/xCq9XYlMBJ/yKEaiMRGkh6wctWVHlheBi/QxNiwf+8oIXdow+0DfJNiAX/2
ZwRtbzo8nSg7IYeOD31JYDfrm9WqT/rfhwEksGGBEqlKnxlO/lpwAJhwbwzl5KmF
pglCFpZQpunfhvvrMB5e2mazOMBzX8KPIktTTNQXMFx+A6L05GyVrVe6RoNMXpWb
/xuJvnXRB3PpVHIWS5ygTnjduUzuccD12wQ6gXoHot5SiNZykXBMd3wWFoVj/eMR
7osYcRIZ+x3hYcJ60PSrUyWeyYz63zk6CmJQBOY2c/2bEfUE+rsWL6+XX2ww3p1m
jT7OUBITczsggIjVPWBloc7cpTcRmklL95YK2eblnWGYQGJekQqNpBxeIRJAf+xR
J8vWbTRKC7oMmtWE6mnQcdiNU2/51g12oaUG30gwBkbNGO6+XeVLKocPZ5cIVv99
qe/Qz1CRpoJmCrfcSQshOrZgvBux2SIsg/jBSGblrjob1/nghyUyl3IBdeD1kj8X
4vhTJGSMY0eTcDVtTHe/b/6ZRiQgF4vVk35fo45/SFCKrXDWZwE6/kts1t2/RB/s
lMm0gJMA15DY9XMk6V5AEozIJRgTZhpTApQUt5kL+1A1gTNv1gsBOyUOFc4ItMga
Q/LJZkZYe5yPrD2ym4b4B7kPNPgWOYS1qWu3+vD+P4OhoGSuBnVvXj3CffoNBSEZ
l2qtWQmPSNZhwIG5UQhNZeIFlZsfrQKA1iSfTPrGlztoteMIXOeg0ynGtxOrn6NV
BH06NZHxU/q4DnipiAdZuCRehxyY/o8meazn8V3lZNTt8oSXVIIpr76VNGd8XLCs
EcIIGXeFCZM1A3CQE5fWJxMDmkjZsBOkO3Vr68KfzNpOzztsZF1r198rUeBUwc4l
J52Z5JXXkEVnj3FSKvbk60XITdTv7+Yj6B2AxLNg/y+b8qrQQjaapvVXi+gC4GAm
EkxF+qOjkzg6H8K2HcfvRJpJVzbMWxT5fBorUrmcDoT/2FlqgLxUiYssRjW1xxZu
gegnrYXgawnUyVpY03fyHVZXgZZVCmJxdhTOkgHnfqvtIuBrzFvVFUV0Qnu1QFos
Sftx0dAWDVUjw0NNS363y5hoWEQS/BNp+gMJ8ugg48SQmMLds0l7F3lNA3OX6JbP
EdBUyYo63wSHquXyZgbK2JvV7Ol8C33sg8mYW1KMTGncLjEzwDEjmSW9kzPj5erI
cDQVskiOMjikbJIhlYtqcOw6T6jEkdGaOhvSeXacQaTef+mPJP9yFW+hotKuUX+D
1qaMOyX/0zC0AdsnTgt44CcE8vjhjNqktZm9v9xKTd6+KlE7b/Ty/K+1lvyQ3DN9
it472VjiiNvXKX+E8UNFUJ2AOq57hz17lk92ZzPhHYcwiAyZwJ0udI7M1FVnIn2Z
cAu3vgL5lAFNtgcnRbhm7ICDIcfsml4HFdLbPrwFsck6+9TSxLK2ua22erim1Hzj
5JbCv0NhSBcdEoK4xONt2/0rPhwswYqR01JQg17mfReV0ShBQEfPa9/YucA5R0gf
kOWqCEQWDPBfbBwxvrVNeIPTCK28UVKJ3CsvX8XWNQ6CUzZ+0A47f14016MBTmnm
REDOltHeeVD3M2fHngNUUbVftjGXa7zKiU5tyMbMzTpYmeUWttYVLK6ae5aZAoWu
uBEqH0hupLCDf2A3MKQAKMJDZDn08HNbyUOfOD4TJpynrLkp3+a9gvy7MC7ZDP6l
Ze2sN0t1Tph+YpbDl2ezjer363YjEeQqbGTEQ/2sj7neLjU1D+tE/AKsiIwbCmm1
P8MDuqWP7JTz0148+c2OBJx/TgBM4ls14Bt1IB+hSwkwZdK9FuyAGS5mmqbHU3u4
6B1SM3mVv/Pu40rO/282J79vzlWptm3R8ZFAzWb3+CoenDMDc//sYYXjBdKSWPfm
GzmaBuvzR2X8tTautXFeNtLwyMlE1QkegM+/6xhIBVWrOHyU46Ovwss/TRgQvOgm
NfmgUccC483xPQoqo5CNigNmo7QpEUhRpvskQA9l3pCxl5tNj1LwbXPrw3QgxvTw
T1PC6DTBJfnQNgg+ZJyZ6afQ5gbLaFUOK9AGAbzxoBO2kAFLwbQGk76PdjWwS8Zj
PN0Ib7cYmScPG1fKF6KrjjU3xQTRowI4fViCBVXsXWn4MYEiP7ePnp8LlDLeH28h
jQXFhzGtrWZtNdGKUaJ+8YX6ECo1cgTYdZBMtsrRKeNtr3cvKGv+9znbhHFvXDk3
rycwtlznKZUW4dKOY7xp1ln5K7/V4WfDEjvvb+F/+D2fXI1/VsGSWpi5FsisFfbM
5bYb+lPNGXY1eaDG7lInvtn/bsQf8KQAi+4fCdjxcG3Ye56QfbtgsmtQ0SVDIt5T
Uvi435HhnwybVxHMdmPFbAw2SY0qr1AVrQLWTm/bEKzzADm5KfCkfChRO7uOxt8/
Pme/Ylv2BdMS29pC8zmuEqz154Wof05QIvwYmP/uEkWAzV0lx9n6q25dVCzLXu6f
PSGqSA1JuR4jnklvGHAl1RVaaduBnGICBll2hl0SqI19xp1ssGlQwQo1zv17woWM
aFecKIOMiO6oUHAy+8eRtZorpCDJkfGrDkYUkgQ0ybnaFZ8v6itaBImWIS1cday5
NEZNyiJiOGqKjxbBmdizGS20sP+h58bdjpnQFKo3a/mq61XsPrAOxScmhRY7PPuo
0KO7CXQp6Fm24Rtrwuy7Y+B8smhIf+UI/arIM2PlPI7rtOT9fivQ06rdV3MSk9tT
1mCJ3aEW44PIiPtDiZVpB4V/WExfpNW2aW9w6wqZ5AYxUS/4llGKOg9wxXEL3ARH
bRXCrqkuBzMbob+rmldy16nHdzHbP51k0v23i5VuX1A0rOf2gXmDF04m+NRCFLYK
xVo9OXIKhQnWmlT1m+H6N0IK1FqIPtjdZWVU6HIBjs04tGsJEK/7uBN5tr8VMYq6
k73JW4Kc0k/XoZaZ2zPUsflQO1MFcgD/ncHQGvcjeNlJPUpip+ksekYFS5vud4zy
QKUpvkaImacPCRvA7eDwquxYGg1YhlR2ktAZql50jUrtC5YX89r70xXYLLz+5T3Y
odvaRBlGp6FbS0RhmqwTtTIivfxfDatYp3SFUSWfwixDTuFEHwdoQ1/vqxZKkip/
jlfYsi6jHKq5euqoNUaK6VYRii9hMEWMKjuCMnLIhpLFr9/IzZW9RagesEJwIHaU
bYTfiozkNT3471gLM7SYBrOSsM/15roKgvDEAZ08S3chD15KElq5HEt4F0d4ATT2
Xx9IlyODezdQsdNmcAg3o/rOJ8t5DuqN8ivzohkbQNex0sDyaDa2P4GAz0/J4EvK
32AbBHt2WuHyfvEbzPH+LdSjsT6YfyT8a3BgGefEMTDuw+/1JZXMScAZav7qJBkf
l/4j9af2uytFnVZcdHwarYeimpyQcXFBBLzr/mIBj/y+l0MRDcevpKWJsG17kuW/
2cKEzhDRA7/mX+Z1QahK1SXhxJwjR8mSjgPUQHQXOBHxijaNxlRIl+uIbFgrWdb3
0NHv5Oys/MYBQKErTcvuyafpXtRlNNDq6sAkRJvjkJS1R+cHpdGTrlU9s5Pl529z
Y8luap03gGZVc3vuJUhQ3U+Cr+c76HZw2Tg0mwFqjobYUmvxsoUF7/D/6Q0NxK3U
3ViBFrxU6UsM08B8KtRIrq1evwcdfsPyCK2h4Q5J1/Yhnpecs6f4BBVh3EMqmePB
emy0D9+5qX5n3trcttE2YsvGIk9qsUEcJ9bryOHOKdNhZKPPY5tER4ghlI2cnZ1S
Ht+zNBOGysfjCbx4QNjQkAHgb4337vp10tr0U4l2NYVRWCDJ7F+5NGrHHWrBqM4z
nRWGNNBBcy7RZ9vK+h3ShCo9bW1G47ENA2Bbo4V1t91mcOidXkj0nKjr30C7HfdW
D6o2DS2aqJ1t1SZ+ffucB/JXjRJ+0URnjLnPIZbS8cwOqO2PA//csFkikmQKDxMx
pvklXPlNOzQCZpXYqbBjZL5drdzH3ewaH6JRU35DvEJTGy86VidqmpiA3Q7F9s5X
ozuPeBG1omxRfZhRH2Q6euKShyVwcjAHz6LEZbmxa9Vj+z6DkvxiNym7HxSjUyLw
DtNGgFam+kh8kCUpDwRFCZGZnK3JE80xnQVXFy3Z+w8/seEg2zsXhQdAbjoGnWz1
8lINyMuefijcD7w9c/n3blHwnhPqRfPh33hEbUYPNra8t1tGDOtz4FwUzmbrG8oV
VZlZJjdJ+Q5Y2WLvsWD0wIvjpenkan2AWjcR/+o1ZWPl5VEqayRdzYJq4HVICHiY
uKaqyx0USpiHeZwp8ArWhj2vKCraPCJiwGfuhfcP0UfNtIMsD30WO8gxzxduD0GX
kC9A49Bno2h75AHdjib1MgFuIdetEtWIURxiCM151u6/G0BtzsrkxS+5IF+j/3xi
APn8Vkm2hgKHd6HC6AGwasAWJU6DxBnuwYaovPup/n0O4jMPR+dEeBQIJuWEfNZV
dwnT24e7W3U3WowersCrODZSHSBj0voFMAP7P0mI40fQk1O1VzRo1XCRCHjo+KUt
wl9BZCR1Gx0z1jHaNKAmegGuz+hQoR1rWMktqnn472XjJh7edVsIKmh9UQWaix6j
X+2pKFBaYu3I1fDzwLDzkMmC/i8xRoBXli5ytt6a6G4J1XenaESC41Kzv8I7/VAE
+Vus5AKXxt9v6dduNxTGZEQgyQ001/+olG2F+V7KbcFhhCLmN2ZX+/BUSyQneiRy
petiMxB2zN223JYT52pT1Gt2X/56xqkQWRfoV6hj4t5WcbFtuAu2rpCYUPxamAnA
IaKqN31ziBYPr9ZydzKw/LGmHT/fLyB6z2cd08XIvvqfxwn5f4d7i4LB/wLk5I2D
IPzXG/JG1R908ih8ywSU/m7V0Ix0yfHlQf1kFy6RFo4Htivv6YctU/S7wZ9AG8xS
vQEWN9SIyRv774zgyTPIoyNFXjjvDJZ3pOnhAkPbkhzYmJxW+vmTU33K5wHAiP3+
6IkKH92YS4WMxix5E2rBKkYw+tlyXJOnCllJ7rdRbRkOF1Eb9dfQJfmUnU5+5JZx
5Clq8Fp6nB+bZ0DKlPIJy4Sm04FDjQYMYRvfBvYsmREX/UuINbquriBCc1FA1jp6
8alXdL5pP6JPAVLEi5i91VsREX9gOKjliX83g+Ln1YVcFuI+1NTPQlFK0EQOauyT
HRGlJkltBJkRxHQhUKVFZVB4xPqkLRelwiL/TEh/r86j5e7W+pT8GTeTOunXzUaY
nsNbsJuEp6A22YjE3A+sO2tDFt053EKNyf0nJKNBC+9RLR+dYW+plZX69cJqMIWH
jxAfd/F7l1vTmpv4umPqZqR3TqkjK0Wh+VKwWIX/86f2mR+OTJRjKD04SsGeQOQN
XAnUkJQ6mUzPZNYx+NZoRsg2tvyDmKsoE7MrNRV8wHoYLMdJm12UP+yUB0TPIAt4
zCNBpuwHTuSiGLpKosPBgYgOIxtwfw5daxFf2aHMvGNant1zLeF8rNxwRld6rqI3
CWCszBncHu6UMbtn8USwlnhqyF3ygpgDIHpf0XzgIB2ymg2t2BtzwrT5bg8asbfI
AGOjQKqyxwi8VwZoaZN4ona2fCiFd29L3xfiTgaTt7v9nZFmPVFl8niH7AWa1MJn
hUXrTI7kmKIqIgT6woWTLOcTJshi/e3ykgoZa4ngxURqf8xNbrPrCUhgJBdOrDRx
l17zpkcyMMNSbGBulCpRjndInyJ05p7uMCU7GCFt1RyHEUa1nwlFUX7YIz6iIQuL
2NUwcb0BhPjsrSSSRBfJHTPgzN2sE/Y+ZHqirRqEHDaylxQVmelhMmAKGuunLEUt
N2ZJ8SUkU7V2YvNoSL/qpmX4gIwYtFojNCHoBLtSZtqCl9PnpnwRiDZ4+V8fWGT4
VUAKhL5DzurUqTDrvn6oxzworIl9QLVW/2A6EXrj872ChVXHAzcFCDDkWDy+tj9g
P975ELx90sk7HFUGEVyCPMsorBrHdiQDZxutk73nYLubIQOgbWPIG66EUFycm+f5
evdxFSa9pdhmDXlIXuKQyNeLgx9bWwpDzDJ6xMbcDN1M00u48t5ojLohWvniBuW8
iibRjHoP9bYxa9mmPiVU3SqWtesIIuYkz5woeyFrdNhmVbP4Vu9HvHojhhgwQakJ
nGPzt26k0VKra2jaNb5Y+XN1tKt43MCOuhVLr6P3UNDomyhqHE/2pXx3qYVJrWO3
yWaJVDoUhJGYywKmip0gHprwrEwKMg18LkaQBblHDbnmjpdHfcG+Vg4NK/vvTo2G
i65JoUHiaCXxIHH8HZ+FCHdzr1kABm8i2led4SfdCepcQJNHj1awA/IUzPh+gYtp
88xFo/bK4WQECbZ/vJ/HRWJti9pMMXVhFZb2q1ztMBydZnoXu2O5FrGpYcNnOpUk
DNezyOvRALDFKTWheixRdwM2leDrCYRT7RvGKPY18lEjDIdyY02IuSs4khXVfgp6
83Fi73klvAHFjFtv+T9o5NRYrwyIlQ5a92cmNV7vFRcZdahpiePzp4Ded9FvBNtI
oFxYdpHA/qcYDVSxdUFuda626RBO5FpKWlqr51hjOSOzi3pXraiuF5AtchvMTI7A
UZcM8nPS+OmZQUwtX5nZmH+WFQtybDYKPWu9FvgcwDl8XPY0YrXKLR/I5Rv4fHRv
AWVd1tZRlfg1wyfu5JtkmbZLKqCAnLE+r0cxKuUVHrzXR22cqfEY0Sok1P48CP96
rxvGGWUtbku9bTQ19usy1bnUP2Q0zfw8gUekFjNsHqB3opcKDqbzOfUqTbljsunU
j1cgKs3BWbXxLc7QjHCT4MTO2WqQcDIt1atJvc3M9ocwEK7KNnEY8UrBQAtmWOrD
/Wv+Ty4hJYk9fggYMzJZOnfooah4mw1Bz0S12J1dwO3XGKEgabR1eJiYCq9x6vB6
Ua18Gp5I1shlWzXfb2b5MPCJ6eJPCXy/acz57dLWhFor8bRBG/P/bQx7oHTQDVD8
IX06pNcB4VF7KyE1Wv1b1MmPCQNPQLxY+Xr8fI2sBXGRRVmEUE6A/3MMgKDQl3GI
3ZhtMWAFg1Fvy24jepJfVjanNWj4j3WMSUG1pg8iBNrBhOX0YaWLBRp0vGSgQ6rd
1VVKz8wlbZXZ/HpG8pJSWhY3PJvHIjjMR3jlf93HKlUZJrqHDzrhU4soxkZbVzYi
94nrRd8vf+FB4s7RGwKAC9tAbz4B3ofYIWK+NjzOFvZ4TCzkQ9taVCstXSSIvCQf
LicRZuMc2HH0f8bRd5SpNi+UNFbJbHEqHfNqfmEWFujON4fdM+HjQeZjP5RB1sew
t+BZTXV1Us1SE3CcIqtVGpJsojag7zMTYSWUM+9om2Z4YaDEassPB2bkKO5A83Tq
LsUPGPK4wOX4ShemQ1DIzmnwwe8GCSLd1RXrxacSjZfF+AnQz5eRN+FvNgLR6jix
gbYlbKPNH21pMbc1Jw5yDOoiP+Kc42G1g1K8sV3FZKOCj46nWrCxcrpaZF8soBJ0
8D2CtHeonc62IEO8VQkFMYIEksl6suTeaYAHp+lLbRE60OMo/AZVlcdEYnIfTFq5
nQR5YxsFqcZtQvpHueexdolnTfJzwdOteFgGFYKXl8LEVtrmIor3TuUmvSDjtHh+
qotIKjyiJG5VaIBMSDc7mvAjU6B3qSAZCIfNOjzmQ4qfrr1v7fUJEhSekeeb0tO2
KVV/gP8fXk8ZFoAlM7efpGqF8JY1CQH6GQI1jcIgUAxBIHA9MDO7pb1/lsZTdz9J
hLOHvazPIVoGAkSVtqaoAoIYhq1+lCCaYyoZhn6q0d1okFnQWa2e69Op3cPI0M2T
JVzm7mwN61HgQ+2ZW9nj1waig1e5rFw3ly3XDen0p5Kkcn3DsKs+iX93kOluEGCc
dPqfPp8ZLbtcniZArMJNvNdb8p2eDCgHdpofi4WM/MxHmADSTdDm5qm1C1Ppd5ae
P4UeednbByeJDTx6m1FzLXtwlX8qZupzFUO2I0d28B65bvxNIcB8SCGBC2BY1k6r
wEMbRfLdxQ6tmwP90abGG+VST1+pJudL82EcvfjWgOVGInwyhs3Kn+u4MrurPQ2r
ygLx9EdPe28Si9dUY0PbGDzbiBYxUCXtWYgrxyuO6l7cWuLzDchVZ3zAQHUyANbX
qXAWEj3Az37Zpe3XWVR/L5mJIX1Qhwxe4rwecVhe/ET/taoZdTCY0P5TMRPXsWzV
6X7wXRi4UffS6h+0OJfmETt22y3k2Q8cr0PL8Vyje6tx97v72TjS6TxghPaCm+Wg
FK2QQOLYk4kX6Rg2ELnu216pKmdix2ICxMdpNaTH6HIc/nwCslm8+JewDvkrE/gX
4CCtGU2lbbT0f3uQcSLPlZNYfDVkcfvEekH64NT2OLLPc3zEy/L5uH16Y2UwhhiD
oiwQsYxX5Y+0ZxNWieWHIrS2ynzic4K0kjr0HOjwRzErj3tassVpp7bCtfjgay4i
eqjQurbRxgol4NRHd7aeQaoCiJYU7dMyB0MgkksXPRNOwIlcHzeZ3SFGU0tqvGNs
ujDnPXpi1N+5O4fSgyDWyNvmnrXtUg6Mk08FD5IUp+WF+yvHNiOUMhOqT+i3vgSz
ezL9YX7l3TCxA4+F4HX24WPYDMkZ09l89FcYuM4xRaN19op7XGeTCvFFzeHQ+Qmv
CWR+5rpLB3UhoV3JtMVACggo38Mlya23O8lH0ioP6byxmBgMa56TAn875Nvb6Hbp
iYQaSHHMaAz252uRwihRZPdEFIwI7c+4awb6jZiTLIpETu2OmjjJoBmW1zgMUqOS
ay47ppwr4fonwU3qPQmF7yeHgkQdI6uOExYVdTvfuA0xIBSqBqvMvzRrJ6a5Ugdk
ieWx/lysmbrxVRIvpyniLCzJr6M8yWNqzaki0QXKLtyESZdWfSD7dHs3zhbKELhj
IcY+gATGBP9qCvBxB0ksMmxpIQTehcxpVP/xXEfxGN+Qexe0JP8DUtAqM9k2O9Yk
LmKGshpbzac7DRRd+1CZW69meyT2I8uRaKLdwrwyQOj5z1y0lAyqKqSMxrW2ZFNV
gmc+81cgQ7t+FWZ4cylkIQsaXys1SMyXYnEyWWD5b+pBK4HxNwSJS0gkDYCGpmBf
UB4OBBNognwfafFMYzrGLAciIi/tpcvR2d5nNmSrQHUSAnBwtAqGd4U9FS0e7LeX
YA2AB+7KlUbGSYYl0Hb8RbFqCeBQSJmo/reUEGDcXQL0ZqOL91MZhsR5SFShocDX
PDja/KDeXVXKQMw8jQxDpi+Sjj0gQOhw8lioN3nPXU+pVMWvhbbE4CQ6FMT1zQpL
2cJTQVT/8GkzmXRQPYP66bcGnlfVOx+aZZ7hxW6UTJfbY3sVv9lZ1ymznaG/D5Pn
7ig1AnQebrNIiX8Nr/1776wZ6egfYqFoHMN1CI/20XqOldJRmYxTtBUjna5tRMK/
3Y56aZNbzevGl4ua4fDlv48y495Ouw6C9YJ4r9FMJrjv8KGCTv2C+0AYCUBMJ/gu
UJpAugNBGOJQKcamSo+udyWdG67xJM5LpIXMfH6Hudlq81BRJ/u+ewzvDyd12zUG
LefJwbJZtu3gw6DV4auXCAUsUuV+tRJ5ZkMdY+J3ASBlGJz9vA1nr5PEpTJC0gKR
mLejUEYxuN0O2vFdwbFc5HNWPs6kQrjSvqpqi9fsDEtLy09VRTwlh1yJfQw4BdrC
i8oIWVElHK1d0kcYS+Jp8HX4Cm/Z4TFOExH+cokNmzkxQzmAXnPKd8kQ8bwOJ1sr
g70r/b9f9YFgOTQR5kzUP1lkIYBoCzb1jQjo6dhXrKVLgPhsWOxSFG0Srw8zew1V
HOv2joysQ1/vnn/guKBQDVaKDrT2gloYmu9du4kSc1JRiE2guppQgCvclmpdPTs4
StRDnNZnG//GI7JvZSaAN6AqgHrOQ1Myuw/7NumyAgqF1qKAxrI7lw57CuhqDGpv
hkLjPzitlwxlY1ZUN4AVMVjlugx3U2cKP/oK/72X5bym+QcGElVvpxVrDbus9MUB
Rcerh8cJ0HxlBzdbrHt+EwY8enNlz+3eMeF8G0Ld2gLgA4rZY+7UvvtBbvgQl5PG
29FXUZx7R5To1Tht9jbIPHXFvmi/hZ6oUJG2WAUOyY0SG6DJtzcNwBngmiPFyGY9
plUQn993n++3EDEupY+iib83WbZ6H/Zy52/y7tRFo1S0qJF9cekMAiQcK4Vhzhvg
ZGOLKquRrsw83Djaf+cZ85IeDLZ6KWUR0PjDQ2oItcrDp+sY1VweknKma1+KpUoI
vveS+psAGnmxu+qD5UURclswSon7b3hMsp9EgW8FKgBCXsv5SsyWO5yFSnWEYlXV
MIqTEkUmD7Qi4u7ars+JnY3taiIzbeMhfszy4AufrG2AR6EyiXm4tM5SoMU0n2rS
lT6PQNH3DCCMh1+jVNvuCrxkOaXf2cW2vjS/fV3gM7/+PcT4rgH+oZT05IonbXz8
n78yVjXGfxkqItHEimbCwhI43MFMPAqGoM+wmXvzusTivt0oOK6lGsoDUJSZWQLF
amtN2LoaNXIITNoxaj3+JUo1LhVAZLfQB4L2cDwWNe9avsG5lXzgWeRaryjr2BYK
15G33uFVqAnsI2hRr1Y7JOnT6W4ASPJ15jQOxlZCOL/AuMLdvATcCaJGxU3boKSs
k4oqLfdEwiA1DOWhFDKQH6V008KDppbPo33xEsxOquG0Fgp6Hm6AFWhUwlZFjXY/
Zlg6FjcPwS58KZTcFqfo9EMVXW57e6M+2bRChusoIA5OdwKuB2Q/+0jRheKQQpqk
2mOY4SJQO7ok8CVuUSvfyn/hlZvbfy/hicGtCb1Qpu4Al3EsvlsrKWTUZbmpDkH+
WIpbvv5+EHzCv5h4obKCYaMBGZOgI4gY4eIBcKWAPB/r6lQqx4TMimijedm+n407
DbKf0tD3RUSjivw10L1T+8Q7Yac+LPL+g7NVn8ItWnitcaAX/UJ7LeUQHbEiwT4x
Gh0T2Ot1tR+xaV1UWYQARATeBZrCbHqyfbRdyLRmzEzw06d79hI24ycYx08aW3Zb
QOkdkfzTn2jlxbeVyRBuJtgmB23T5V+YZ1EPZLMrbEArERAnDTOhi7x+zfzlfH5A
cD6+tw8ySAxMOr4vmtOY/E8mOiAy+O56sh6Rf/6YvSGtA2Em1ruIY3oTZqtiN4CL
1FXpqZ5tYmIEfzU9BT1foW6oLX1M75A0y9QRoZZzZDhbKxdppeIaNx6chVh/rZkm
BdwkwP8beFyVDDt0SCWsxF7GzF4Cv0HIrTgrp/GURGhpTFrW0kPsOLOQlReSmiWT
a+M6rq1UJek4/eckzDXgi//diCeek2/1ag2vo/EuuXXWy1zsvKrHzMJ6wBc8G+Ev
tyU0m1yz6VthwnFFxaTf1HjRGl8d8+pYJ61gCS0EQKdoIt/9wdHDS1Ifc+mi/T+x
DGfYduEKLNDgQj0N4eB3LafYvFKhmi67sM1uWhUxkxuVQGCdJhpYBbzr5kgdaHIN
JwJcOz50ekKToWsclWFeEtY87J0eM+tJ8NEhtf7B7P+eORjHoCU0glFkbd6Oy6JQ
J0CjIsq1Jd3P3STQkvqCK7PoHpknAvSf1Icp3tuUnA6CW/6OLuEJt0EzIWDpt75U
jOFwgq2t59KfMSohO1/ruq/1o8tMj6pXrG1pfaA5w/xEL/AgEfvNoeiD3qAnGFXc
NufnU6j6f3Ivqw4qA0Cu7lFHUnjgnbjWJLbsQqfUoCyX7w6J2CxSxapf9hrNP+5P
4eO/T8iGJ6Y9/v4+4ZolGpoUmeMLbQEuSXg5dxYwgp8omL0ilLQ4Za1OpREIwbYf
JI45TN7BIIThGDLdESIHvmvvxN9UieCsPsB0VQmf6ZpdWmq6y9gf4q22HZjEAhSE
R6CyuBC5o5IEDjBblyBJqY9np62oUJ8rghaOKFjpbXulyzeljZ+mOImc2yO4V34V
GI+7mm+pPk3rgHwTAO5YyXXn7+xhtDPbRtAQovG2Pl8uxKGorx/nnqTBW1Cz9/dQ
3eAJ8VBCTzmIX0x0Scx+NPhQgAVLIYor0YX8cHfNKeC6sCEx0fjdyKO0OddLTzLP
+byYgYip9ubagwsBCHjnEXESn5J1a3aPBpcItYz28r8LR8WK1uAcclJljWb+zAwM
OGVlNk6fHzi/drUNWVuhgQ/Y3TkGGu4zYa45nKMb1ES5hFoF9MCdAVVqJqaCQ+CD
AtDNgWOS4GI9FgKxv3l2jAVsDxvsYneetW/rrBIcCCqg7zCuWpfUyzzZ1LUZILgY
ko40Znllf2MsYc62r1RuMB8ot+iBEsQ2L2tuSehPWDHKAawpIFqwX1RYAEUQs6ZS
Wip6iVerCSDsf3VAqAm5fKsQDFJKllgMv0Hd7ypRW4gMMlZvZzbCFM45Cr+nsHKK
qs0tyaZIqh1oD65cm/ZD5c8Mq8YX/q5xiJj4ulp/weNbCZLsiuaYzYTkWXo+fhtF
e0y4KjFGY0J/sNIlUq/yqquDSP9k0N3cPzgRJARauGbc3/gxDlZVZTY0X96rz8jQ
KYsKPBTol7bkqHe84mvcrtBiq7UyF0o5xFehTCoBeVqEtu0arDgiNPyHW/rftObF
bal/vHQTvDsjM8drpFdsdz4HAhAoJZ2FRCAspTbe6sJtoBvw3h/YNdLxMlEsi89l
UiXpUYmjkPfsaJieQ5lOnziFbJiYWk7gIY+gB5AQxG3GubbrfyKghsJsaPQi1Rps
5KHXXJUueP6fBXRObmuVK196D0YzJYUWgNbdMKzce/MNSlZt5mg52gJxO5BLCHlZ
wverdF5VrK8pAYu+EGvIRZoXgu3KTCmi7aI4nHG6nh/qtd85/LVmflmOY/FCK5G4
mWscrjf9y4f91shkd7ILlH7/YV8FfRqGUJFkOZAXye66pKf5ETz8RTVMu+n4JetF
ymn2ueTBfRe4TA9l7T+dxEZG3efAeirmSWkPPlMkXHlQQMCH5+x1Qmk2oNB0ssdf
HeGplk8UUASmYLmOde4n3Y9Cpi+mEQ1l1iLTh0mGkn6m+R/sCGEM2oJAb91H3Baw
wVuvkkMewEoXA1tcDznHHVfbiOvMJy5I9//XFZEG9Er/8VmvaDFxSl43ytJwyQyd
iXsEoBZepSxDngTbQ2/JJhogDsmAwwflz2qjj7pVVRr/2K7Lm/78aLGQhisTPCOG
He+RIorxo0DYoghOv+JmA+aixGOcFbj3D1iXCYrlDTeV/raQgNp9xF/ukEZzbhg6
mjDGFzvr8yTyLS6gK6K7/wxtwTE/+/WXRRwQxjqQWSuuI6k5mv7kfkk8gSeeHBh+
76cW1H2CGqzejywX0FqSZdAgXybACCeMTgVq3HpbplkEM2XnRLr1mP/O1DvvSJY5
Tj8H1Pp1XgUQipkwVEyEozr8+AZ5QLKm+eFlQCC1tr8vn9aFuyIdiEG8tRLjUy3W
/HXxNEBtnP5XMnOaFhrn70dXUn+7gB2nbg2+lwEn/GxbTwZOE9l7iJrv39xDTeHc
gSVVbjiIVAaciNgE8zOBqL7oMa2LrvFIXB7XyTDVovHeVYCEXZSYMI7pXs2QKX8T
GMVymEH6yKw8+Nm0M7lOPQWVlybZVvvzDU5PZ8DesY0vuQbis2MJYA5YITuD35Fb
gXLtDytaHtjWK17XUscruXPIJFpxXRzEj4nWshxLXS4Do2MNLgRs7h92ZkTTkmpX
SC4OEq6gAu79L9QxBakNOr64Sc27M3kacQW4hRBEt7hYYHhBimOJQDwP/k4X1xSY
ClgIxVzhezLsJMOfowL8jRfM06JV1QEMiwggCK4sjY0n1u6BBUuEcoaeFIZhMCuZ
KmHBq2XxUFOBKnMIilsNneoIqLQDCQikn98r0DtwDLB59Jcl55wW2qi1Aax9NZWF
BHGMxPtkngPJDq6GcA6TRnsmnPU90W/eMOuN/ZBxf8Jxz1KHs1noCo0HqvIxcPkz
SJL7h9EcSssX7kVb+NYlElMznR3vlD1bFAJSf8TUlF//IzCWCeLENa0HmyGaZ/bW
eanl7udfUWFVcJf2JGadDULFMHP5xW57BEDeRmkd7Zh/PjpRV6I2OhQBilxf6qGC
4B5YFkTzOxTm1zUkMHtLikEU8x1M18/mYXVVvzq+Bq5fsEZcu/D1FXf905HTyR5I
6qrjpKMcbX2ShoRebP36h9mOysI9ZQOFkiJyc+RRDCcwkzcIkcVzlLs+KiJkUA1Z
Uhw5Xee5i14FHWWLScOFglt3Jz3FjJGGsfaP2Eltxh3uxDDOrKxHnOIL6zIesYn9
s8HnyWUSlqT1sdzqTqiyL/uMR/fXcuKCgn9k1FR3Bn+uohrqgk6Ad5hSUrdnMePa
suWjmjxEi7wNxw/JLaY2mXTxpX12ilAr1tfwGi7ukV9DhG3hzf0S5QOBhapM42qg
k4wmOXS+WOJ067CffTHaLyePnnY0BdZrq4WieMfoxdpH1Woqx7ANy7fFJeePaEt5
HFPif8/TFXI3gWqnHV/EvaXPn9QnbVEHEjLBEUtaKe+CoLE46/OZhZm2u2kxbEbv
/b/FTNqz1yeImDyd7vu7rWZjcLsThxdKLx72WzRkw/+BrgvxaNmRJRNcZZS5bRZF
kEEWHXP+ZuH93oQsmzXJxpDuuXmYlDp3DFPiw9CwdLD4aZNcPTSy08PWpgLK/XUz
iN7Y7w0hkNFB3ITmnTsbocd88jhpz2B+NY+d+KDfIEuNWHlP8MNFsJRtH0HwQm57
xY/suDcP+yDvKA0TbwxInOHidBb/MQcp0yFctrvNmZPU1k3JrrgBm49c2U2Zlg9u
Gj35IjACTNiGlvKNnq4moMiXLzOSkciQIKDZzEzSxwsK/Enur0wXXihok8mfuJVn
mmiCo/8AXJwQCtQONyKDHMzl/m/oguxcfEHSD+gHeeuIBhKdCGR4l8witARruYJp
Gp/twvnOP435tlIDf3/gVX9D4M8UTghFhMuDQ13QVpATLk81F5ANF5UTePtDdZuh
SHRHMRCXmIAuFfKLWIvXsYQD7wRYnDDrvA4F2WCQXAKWEyb0x4JsrQ30hTgn3vjz
lZGuuc5ZL4mrnYftxGyeaScKEvayTb5JlPS4dgzhLeT1tqK09EumlTRFbDCm2/7L
4XtkUpESGiSM6cRZ+cAMg2lNmThsrxXTmJnEa+i47Rx85HmaqB76tjDK4iF73cE/
h8/Axx26jP0SYCsP5zCjmIUFLoOuViurWZr9T82i797oFjOY4cPOfgL+eJ9wjuVL
GQdWhZ47qw4Ps4XzyRCCkPH1O/E4WTAWt7lnhXeaA/MlS9wFt/DL2lVMWQAaEZwY
SiBKInTjEgat7wL07y2kxKtDy3TUYoWugqgxnZCOF+jF+ZqcI1942J6yZQeGf/D2
+yMRAH6eswN2VN1PRC0hp4jMRvmgBKVCeUPEc3Ys4MEQqyLsxk6+q7Xn/TD4xX4O
o3MX0xcvhAR4JHrmN+iIEciI9XE6GozKcPiJ8beWo49sWsNXzZyyzsj3ND2kVZny
r4asvDUbVRgcQTcfdUhCpAxWZ/Y9qrjXM+Gl3GPyXdIEYCrsikf+ivTiZ6hyw5wN
l3WlXbYLvxT6q/p8o3iAeeRK5CmsLUU12HehkYC9xGaNR/jjZUpM83FvQRQ1KgBu
h7IRgGXWmHaCPXFkYWKErXuVGRS/t+kkV3Bvgjx9Vl0VeI9GUUGnBWWL8okoHYgA
z/JQZXf+soCkELVYKFNRxRgc6aWvuexjf6HgcsZgjZAePo2yEew4UpkDJREw/Q3v
+1S+tHZM6mRebCHg4DyAweTMlY1o8kygfdWE7y+m6m9eiaOIzOmdb0eaIn1d1/D9
+xM9tpi4So5emSqtpTIIkpRAUl5P6MorWp0g4HL5QT1++QbMsGYabxQ4npVaBZrh
tvtZ7AFJ4qjiAG12nDMo0h+nbda0dfMkljj8UaY0PChZMx/PrSe3guCIFQ3X6sDx
LEoaE0QMADgJLUjBCSTVlJxXoiOk+GlfUo9gWgZO2ef0eZbXxCp9sVSVbxNe5Gax
Mj457gR4H/km7auMdYihCgvypuqNkpBJwt0zRhi/jZtuMcnkieg2U7Znjde0hvvq
fBMumbNRwaoIdPVCheKuPwLxtcutQQorFpZTgVTBLbSM4mbpcfwJwhenjT8amtK1
/UXGMIxZT+4pWvfgQX8zO2XR1nmJT795K5mgKimNhbzw3JS4d8cpkF9NlSkE5WGP
GzLpv3wTxEHuNN03YaG6gEKkKJTNBUQ+RT5nm7SFWN1OfRmplF1GoSrossagkSYD
ob3Vy8+dCAraCRh0DqYEUzIt1MZHcdp0u8+JWOlJSZhzShVlh1FZQrtni0SMxghB
d35/lKE3dYOve9lAsH5FtY6/TLeFLPxwawQactbqwHuKOkPXG6e+pEMdwXghCHfa
7t8TgspgET+v7ruPDBh8uk+M1GdDZj2HvGYHsp77Z3BpnmRAp4K1vXWDoxgTqy2G
eUj/e9O7uqDJcWSAHgzyfFmw7LcMBRg50YcO77JWcN0O9lvSMXDa09F3qGqkz5iO
3jxRKrDIF815f+2X4dp+Hsi+kK6kWH0k3tmsCzmke49QJuqf+F/AlMad1eERsIKm
WEgjuxphmTagA0fWJ10Und6ZJjzsJ+9eVRlxifyaGuyO5tZMX2/3UEJqroeH2hh0
qXFZ5alMxOntH4lUX8pViEdt1cSFoxW2+YeHv4RLxo/PHxG5KR8cSTqymxAWUq9I
U6A/Ha9FK2721u0ciPa9+smdsF7AB+K+jm7TP1A1EqlBExxcOUERBbYQvlKlF332
cjuZNqyiMGV6xYkKld8MWTQZKBd0Wh34HXphtSC+slXd+bhALfYptOQjU3X8IeBG
4HkakT/LqSXDumhIhGdK9i8eGiXjTy4F9SOXmUwkelJtDACALSkEM88SFWtnoFjM
hbUjvO/gHEdaJv1wEDQmYy9WwlLYPRDPpWVrtXhp9b6/MT1LpjsuvsjRlWMKhpu1
vL22Dz6rDCV20LaCup1t/aQh/aS72yavZHdANgnBisWrM4u/MNNlZAQCp29ICseh
iVApWyk1yV/X+BUrYpXFPmdiYu3guSJ6Zpb1rY9YTrpXtqvV/ttYXu1WPYa82U14
LAzSoxh/et2SAD3F5vBVcc1FQ0UtI5F1o9wybCXXog3ovGDE1VHZiMqdo1caJnJe
j1NorVSihPucBNoFc/is1toIcCQfEXFWTuqSBxgKwgmrhXq00/L84+vO5ngf0kF/
w13/j/HHsLz3+ysPjb16qAoeAIWrYOaUpOr0yRNTelHeLykMku06UuqApWfcg+8F
XNrcAtV8pV5jfit4HgeSn1Q4XmDLWTJiTu9/UOPfFWrP/FC40dK5z0vwAXMa1Krl
yrXLb/qBiohrA7iNM6zBPJAXFDX75jZuP9Vha38Uvv8S/3IoIF8r7x2EaNPr6ZRz
Lq/Mt9vA2a+Z2IScpIWZWq3P9cipZH0vKu3MdgCi/B1MqPl+znAcN4cPMquSoETH
zx4l4zP/NLbUSdbhE5FF4d9pkEVeJmFdcpJYhTuGXIpnxuhOzQj/EtXGLXH/LsG4
7VEk8jMcnSU+vyRS4NMR84GLu1h0+NeJuA4kriMZNONbxXfUgcCBR4jHgkElieVl
9BVRxDBkKUG1SDSrPaewkXl/1LA3znYBQVBDNrX2Gsi1q1ylvQW/ox+8Q34/VKOL
x1dEaWnoQmGBxPGQnJ49QHsIjdkbQULdOXO5Lc3CHAXQ8Iz+gtfvlOxdOHJFF6oU
gZmYeEDWUILWeoCwjnsjPBQ4BiT4z2fehQZsxUJfRfQgUuhdWgFjx6yhBipDkhir
FZIbhJ3z/+wfsJA3KwPYpSaTXYTlhHkzxroDEwPn++QPc2YV6YMyVJxHkBqk5aDX
kp98a1P0ORTCsV8R+VhEw1JENsOsPqmwsIg66EYqo0VtFYrcOroz+2SkdsjOzg1K
fCwY0YEk1ykMPsOdgLwLK9U+O5YmQ3f6OdVHxWy+RmnP2fCMpIstFvdwTZrulgS6
A0vPhnl5oX36C+t4ZKIiJUp0hGzJmUI9iWEN/PZZUxoF+7BqqfWy8rxu8r5vvwZI
arjWYb2i8AD4QVdN1sKO92MXgRRHegEqTNHw8uInoDl+zi/pPggK+nQnWytVWs+l
gnukphY10det43u4oCLaEu/1l8trZ8mFTd9LVlckNbCxlyMhsY7RjiYJKGi6Rfcu
pS2PQmvvwgfrDyxyeOi/n1QVK+YZvJk/8aq7E/NAedLyAsmYULe/IXzwU2CFQpnE
lFEi3Hl64Dyvs81Mu2wK04X7rjQOqcd61YrxYQUBi8DOjm2Yxppfgi8FuVBgdjCX
YinKuBfJs+jt2c/2IPJ/NLmK/RxrW4eQnYsuv8WZMFjt8kC6RiX6cfiTMb4v/kns
RQ69fN5+XlrHnMhDAaOp3NnML52SDidoA0CmCj8R1tdujsqTyZBNnvLsSn4CGYWt
0jLQv5YfCJgSEdh/jjrPcSAJ14mo1xxrQHz5bGxVV4eBdTTFeDmQIhaRIWKO82fq
D2umQX3FydiTspJUYe8RPAp2q1VP63l+T6IF550rmqRFrq2ipx8MosltJmzgLN5P
gvbZBPLgwP5DvrkKcD8cUABmbp7N/DotH25trBSYnAFeDA4FIOx7xbqbflxRMesl
yxzZ5rSTLMidWpOEpa2xDPikLaZVAwaybbmVrtFs+WcVQHMhtYV2Aiodzg3W0JhJ
TonYlwacF1cJ52Ru5nKjL9rq70U1dGvm9SzoU1bLEe0mvLbLaGOOvSxTrjOttwb1
G+m8bhaWfpkk+YselXFM9qfOlqUMuE1vzX2GGU9pgrv/EbOZDJ+8L4+wx+YNUb6p
JilpPbfKe8JHNQLRLR/IF7isLJMClFGr5l4TorX7Ork38o9BerVFStNdgz1O7u67
VPHfuTrr1uk3SBUIsturWSkBhYaAwUKKOOtXztRjgnw6Mp5wnUcTut6upeLbbB+J
L+hkZ7GuLkNXtEMk44fm78BxEuA8WLzmnZSl8rPlegdUwnbbgZ6cI9/ZofDj+C1+
YvTGgrKJQKfDQYCrXRAvCRFz5UkbxGqtXBUtXSyBBr9JUyLsRWRyq7rlvB1cZ5jP
ELZFQ9IspMkRp50lwT3AONTR2pBT5/NW0OsrKUEJcuWxTy8Rli6oRXzFLY52L5vE
DSqiov1PIvSmH0MDFsqiYG4nSEQu6hiyG2Q6fImofml1Y4ykztj8x2UIEQFRgnX/
7gNC89oeVm/6AwBCi6h1y+YftHD5vqhL8RsBTDHtkp8rtpNtCSWdXBAsaToKP9nZ
py9nN2auqjLwDwmoTjdCShHvVIxWaTtZKvRGrIGtrPwWOxGRxQU9C5ZH8khHDZRo
YYMRO6IuB9JDEX+fy62rce3G9X8MmjVtayEWTR9yxcJVze1Opa8mgAE75K5J3Nz2
+KGfxqTzqbjCTyxiXToQrFCFIwiB/27eCvu5AK/lzkltRW/BAeNWrv4QwJ+PLyX1
m2mkubUGPevL1WWiAwuTm6Br5sHK600IVX5cwJK27v1QkKNI0zqZv9wlqAicT0by
ZTZTt/EkOwzC+R6OKyTfXLwhOAiiIrvMDAd8YJA6cUJVxJTBGzbPACgP13s+5nh6
HaTxpSZW1YPnqM49A10xd1bR2nNeUGY1Ia8KL1I1CQ8gnsklnC2kVtF2x6OELtBo
9SbTi8XRJWybTcYPLCqGbiIeNY3zPN9KJu3ZuvnSAzmATwblO5pORPMgloF+kKxe
BqPQHH0KcIneliMpNPDee29zGF5kk/z0jh1gVHCzEsNvZ51GX7vUQUC5mEI7Z2K6
KcFRck6hjxHSoQ86H9jvOHHFfxSASgGXimrS33rCIP9fkdkzEbdYqxQjeLuYwGn8
BjicRVxv7JuMxLnElwee2WGkmeTT/iuiPjkxHhb7lWbNqXkhEv4xWN87aYWpDXx6
mQUZfhTSvDvoiQxznE+WIlIiSuEDcA4wLdvVJtPD4/H3w92JMfFb7Zy7EXJoEQ/W
xIha7h3U4CtIiq0Sw99TQE0Ybfx2GGKxWatekz9KZGIWeKR4ej5HAdRtjO9ycGZV
ifMFYa+lzMG6pOqef0QzZB4kcfXNxhPcDshH4gIGkMy7v52IWTnSGYqvxFNfmgiu
88RSXOeKXKI44spxcDbZSNYy1mq+Bpu+7sPblhZYh8j1w1LkDQKZudipbnECmM3c
hXsIN0LWRzfw9ifyrlvdvAl0xTgG2EA8Z4VRYJ+y+f5F+Ux87dxfhJIEUn7k9oGW
EkPHmUbXjpifVBGxHwEvqpvQz9PE5qs589mDG4EUaL7qL9UVme4Zq4c7BVi7j++/
nIK7TH78IdR4dIl2uAkMxT0k+S2FSlglFV81Bq1uVoNdDzjZOt9vu62xv8XV5dEd
K6qyc3tsQCK6yBQX5m4/8Hsev9066tKLSfNb2EOULSgoUeEv0fHKksPoWRafbozU
hlJ/5x1GGkxA0+1cv8aScQ08mk3YfWxVg6LuVMXQouCSDuxlpIWJ3kpJYAR42EKy
NoCdemip5gMYjhpLAR9ORS4u/emHUnAK9Z6I/tPB2hXGFAmlj5jVirMYpNj/+Wi/
00K412NZhVzQ+WAkHEy6k/0QO/x2uOgTI5Ackf+Ij5wzEMpb2sy1cIbVcCbGqMr4
FKtS69q4/LOoH5oUVnhyBqVhdTW2aioRKyQJQnABKkAMOeQkcVlcX+hlI57WUaGi
MG6efbim2ZbcNSDJ9vdyqnImY4I0cDvP1Nqetp9CrwTbOBY2YR+SQRoygFT4LIGq
sqe2GzLiXL2l/buVCCEWZej4xOVyF72H6QGGDsuVcKor2r6eOTMW+rIsQsl5QQ/P
6SvIKxjPX8ZFQac/KyurOeHqW8flHV3ATZMx4SvsyfQ6BfEG90x74mG0RgaBy+7z
VI0VsFfRsB38DlFMJCeKuPgi5Pn38O9Vaz7hz2k5rNBd8bwOjFcRwkSS8rREKwPJ
uJOfhYGsjHBtxWh9r8DHfUwDnB53L9yjl0VQs7wIde8lhHcosTfCAiYDSGNzfUcl
adTlDMg5Wtdk0emhk/cTvq1XOcZNJgKX0tHJiktXtzihTtpXZnMapUBgdP9GzT9x
8T5aRh6w8iNtePXB4iyWV1LpMTebRlLApxeig+khtLPySbqzRNgImOooUIno1sYg
4pVpvlTCnqbpIbO3DZWMO71qJ0W2UeZBaj39b4vZcE5wfyksb9DEqnE466K7yySp
tH1I7xhIPcNiJcQnxGENxQ5HN8YugLX0vpWILvDS1qVRCmBJcrIry/OXOe3C3W+3
TytQKQtzNPIE4wlP9wPgVZnArn+QNboRoXEXuh4pefDkmd85HCUTsQE1eOFZSsXz
EVh/jrVPLdbulCFkqOoDpD+QYPUAsMrC69tvnHnkLnuGCCUU8CfTiuqmu1xW9L0L
Vu65kICR3l6Oop2ttBecLtiwlNZlxXn7bNhReWK0BfvIgDatK8XUBqWaGv1g4lvC
Qt7z1FZyhjLIPNHay9HJTK918FI1CDJ9wqLcsuLZIugiV6KfQhYmWpJal74/8uXR
9dKL4gCM3CI3S/A+2U6IUm82cwkaYo+TsfWoNshhRLbdXp5oD9Rh0O0wK+kLkPVm
vAdymES4CBJKlmoTqEQi7PcvKK1AgrPqmBFHLOPvhs+QBMTPFy+29SYM64nUjS46
M4Iu/X36k/CX70aIhF0Ze6/6N1UtyxNMfKXrbXH3s5Ca07p1I8RB+HTooP3as934
3p8Exm2d4WpgUnDrT/6M0l7ZYgHkwhbGpmxp1sbvlb+FgMiV5xhejVR9R4WS1NhB
BTNkDgbozeJgQjGHAd2zZa7oYmc/FGN6yIr08P1QhLHjrgFCO9mwUmVMOt1wuWwz
g/1L8wx6OBxGMnqk7cH+azTylE3pr69zY9BPq6NFfdDF5dPn4ZqOhUnnhUKx/esC
R6drlPoBB1dMa00Ah+amGovYVBmS6e8FqXbIzN12N3BGGIANXzvcLzIFKGHIJhBv
X1uzJjzCUcARHPYgICzYW0K9SS2s3nvFG4txzDHfuDEHUShqhdgM0ZDy7R2spen7
pRccMaO8PEcrzDSPavdNFVU3nuN8HLlpkT/d8qoMIVKbFubVkHrIbeHmeRrK7GPn
r6uBCm6LCbn1N2rmxd9gynSC9yjuMVXvowSV76Ul/w/lcn22wDXMxVtrsDUJx5Fi
V+/C2eLg2zQsOtX6JKTxQsGZj8Cffnb930T8eF+FGRUB2WMqkqrpfPyIcXbWB2ix
u3xXNSFQ3IGGKFuC10tv68LOYGlfwD+PcrNtRzUoL9jY1/1q7kPVb2blYX+AxYOo
VXDZiJH8vK2GJdL2AOgmJUHVecaQYuAlOOgFA+hCoS8/MdCtwAAEU/esPBr2mciT
AaOA38Orv7pfsoI3sQRk82U5wVxKNnOVmtK4iAXSC5rVH7gdtyycHmyOkNMfCjm/
wvdYF4UHaJR35yvBzJ1A/vIMcsB3HcE5dVKW/MrskIqX+qqFpUynxK4qDaorWm7M
f7gbxgI43FPLezYql6l4KfHZsyiutHryzg53NK3fn55E7u51pVPHD0UbKtXXY8aT
t5l1NbdNq9CMYate1bYrDSfzQexksEiE/CyNFlJDblAcOKwgowrtO/iDxcm/nNp3
0aPO1luMR+XPsOtFNNUwhBSs78RMxt0D3CMFJOkYlthiKBmH/lad3TJpLIqnjJsZ
MyTyAR9pwQL4OtlM4Onx3SCXklN5SXBDjE6pDcIBOO5gvV83E9dqaR1C0uZt48Ke
feeFMhvCLtETTAPgnbv8maBFOLvYqMIgzmxGIQHG47QtY3Ak9iE5oaveuOhZa0vq
PD4oAxtplpJTJrPRxDCvN0R1Cu6nvUdM/NkxNVd0hkssO3oPUvMN3ytXwhTa33wX
fEKK2caZVD7sASOeerv9rQRXHwl0w7MxgAuI5NoZ4L7tDV7OZdUHYT45nCiZVLwH
URxLJjyWZ/YQWfXFQBgXpvZPveXaV6nnQG1kJMKLsyZHHFJR6t4sVk7Uc+jPTkPc
nGCpUsO1z4L05US9oC/84An1wNl88daEo1qfV0JzKFW4u6dncKSX444/kb1ANko5
RvuZkgn+VWUVThd1ue27kqPPJz5yH87O3vgz9GYw8T85nAjx/spD3Ah6N3jrwILg
Jp9t1v9SMuk2qWCI3TLBOBP7TcMqpJf0Rw+PMB0hSor2Hmbu7EGcnjO8NuqLvASR
Oa30QDH8V0euvhctr3GwS59xpqW17B40TaZZxOsoo8bkB7HeqXYoIA7qA9dUl1NZ
DO474xWs/rSAu7QDzJm3TPF7KDgCzLO2gKPwbkDrB6xtrGm3Zqx0Idc+JYS8U+oJ
s8I0iEbULFnQj6zyHuCMWKMPJcymICsFe9uzFTkLkdWG6GljdrnHPW2fYZj2NO13
FtfwvaFHfhhD4XKp9N4IYfCTai2ZOqvarBP2T7PKeHGOQ+7Fpxk8W+gxr/80lPt3
Fn/wu9GI/2uiG2T7XctMjRFZyPdjXnaZ2gOv6/3LlK3eje1OoiviPVYNt8fYdHKn
ZpBgCfW33O9xlqmUzDRmHaOHqXFbZTDNc+meTU1eoQrbnpT2Hi1gm9DYbztbyrAB
evjocBTXFIqzlj3b3Pl7j+5Ce8iNdr3WYvFnoCGDroCFWGjRQxCHa1LlUY/dpb9M
Kn75v3GC9Xm50N9HeOV3vf62J/2pKcoC5L4UVt/4AmW1Iur/+g96ZDumxJOwCM8o
FwKvsHPh7tMVgWBdi/kKMKy4BfH5ERtuRpr3+L3HU5hpMcp3x+1DrA/x1WXWhFGc
tHcsmGb8ddh8vy9R4G3b77/wvYs5meQXsfCiRGeTvWAgEj29HNRvB8rQ4KXBOJ9Y
EWa/57BR0QHC/i4wFWq0kJaHWNiP7JETes69qtR/4JFqzHbNiy05n0+hzLK8x0AM
du3QNf4L4ztf8rqjIjj1v+XIw3Ve+ayPvIepT2T9EscDmBfTonu9KqpwaSQ4Wtvz
mLESWqK2/07eb97VfEbfR4twxLum2noQjX2etGNHSvSrUxRXLFzMGdesu80SLD1S
M+xIe8RgPjIXxY/sV1137AHCLxWSVJXXUTdd9FAyEMzXj9rqO5MJV+B/8NjSpP9w
Y4Qz6Sf18KDfG/HbSoFNEdca71g3gRn4GCQn9T2/NgiX1eZ0bLhEFcxguYfFBEYT
GTZg1yQ8ghSJl1BWmw6RIqq2eLEEdZaszdk6PJAZ4BkHt2SbYPZvTMSR/2WXlSEd
ui9Tm2nlJJPPoa0EVPHPJ3UpHW4mtdsuXeiIbLtPRmmDK8Un/nHo3EHjtDfgo7ge
jXUyeQgjBl8RsdwUwG3Pximj7QzpHJePhqNc1WHci+oIP0ukbDdYxqDc2T3F7Bby
HvAyFhPz032Cbcm7rkTj13D4D4EEFYmKdzSThCv9OFCFffIMJpsMlsr7epg4webq
3MhsH8PuiLXnjO54R32KYPbd4UovWXZ1SdIBDPEp9f+zJoBBXVFLxto4dhxuOwHj
e+Hs4UCuvm2HCNr8gjmPSzXmyD2nieNhaqzMWRxfdL2Tz9EF7LJUtG3flyPNW7UM
JJqmNsLDO8/bprCFlPRopTXPp6tAlsE509sUmw6dKTay6X3Xp5wpJ6FElnx6ebSV
5txy5UbOv+XL3xQzCxRMYTH8adSb4WOuK05j4FS1ca3efBVR5wrhzyFtoFeQYRxg
Qzajb/JcrcM9RUSDNQ7BNIsIYIN7V1vuOirUcWj8I3dES7jTOYq9+W+FcFFLQCmo
+jFSmY/qY4j3ydCN6FzXA8aalt1EiOLqMHbOln6wY1eFsLanazaX6//oj/USBiUw
TM+hsa6mapzl2oNovOBCz5OfOvqBL9UHDNGBSL3uWVO+HGE5JUC7aMn/PcUi2Lul
rxCCGp5mtJzi5FfIpYoY2LpBlHD05CXqZzLegkuiaUIXoQ9WOcLUTVPKKt8xNyrG
lCxdIEGy4MUQ9JB03jN9Pzevbf7F9TgmlnEx/2Xkc2olE7R9hjAACfwePB90neWg
alBBJPes1dVZ9U0MmM7/JvSuRTeXfnHv7v/Yzq/l1KfdSfXfSosygj94WLABHnQO
F89AMlVV3Ntb9c12H/hKshCJILq+qHwdRFwKqfvt2BQWjxuXs2fqAXlKgC9bRdZE
Sc7d3tW9thDWbDglGfwnAubdmbdaEWYhZ28JhCpu5DMyqV8LdhbdVbRRMCp2Aqr9
+1yZyGRZubN35LA4eNSA4xelMVKJ1wBVPy9MOjmgQ6qpFtvT32upxe3sTth0TNcZ
91CUTfeZjVmrpDbuBN5zyBqbmdF5/nZPw6/99R5A6qa6c4iYeohbQrRKWz2IxS+4
J/2030yum8d4qNZiAPKRntdZXDMBWMxOI9daWqYH1gUHdrh4r7GPuc4pH/HnU3rw
zh3XH5RDVZckQVzm+2ZNufUouMo0Zlb4uYJWizwv1MUiolvZ5wM8c7d8ietkpG9Z
abCJVfnHmMy9G3w4UIQoXEO3o2IurQg1rCAN+WlzQeeE6WN11vZLTYaFPkwIUBjv
VBheLCKB/LXookZgDC9Jsie5MXv64O5rXFK79U77L77qC0U6UWOTa2XHqNqRRITC
c9yN4+sRqmnxMKybXzv3pA1MjuZOtO5brk78azpTMwsHxAAEOF2Zo8X66W2yASnB
NnC5aluiM4w4pVw3ZeYA8uBbcurH4BejAc9PBsxWHliTIwPtnJ/vmJXfS0oe2+yi
G6yOGN+76lMEIFERZKB6CKwxwEy6sXqcaOyjkvdB0IaOngGSGbPE58PhF7EGHn8u
nSTwnJM2QF6v0ptN0RxcY2YRikyPUOjibAh8ivVbtQ2g6ILOFkVv6BldtmKcqJ69
k+tANPt+Nwb9Wu4pQ7lZGl9cMiIKHkjjVE7jyMnvZb721djCtIs3NQXFsOhmPLF4
tpNDHMrxC3AH/n+1vIp9HhUb/AQg9dlYTQOg4fuMLMWzChuCbqKAUk3hjUC09Igv
xGciK1GAQkSc9IKJLvazdn47y+jm7WevfKtL6lX/smSv6eJrzijGEzHGQU2eFoTy
rFF+uzTnSgilynQX4yIwZsGnKauVmJxSGuiR8Nn2xGM70H3ckPFCj9srqo9SqUDr
yOdPeZexuPIvlB8IlcnuVX4IpgcCuT0nNSna/kfUy9Xf9Do58T4aByRn7AThp4d7
SGAtD20Tx8o1abv+hge2elZyuuv3aYgPMmaRUA77InYIQzSvHxVU45tFO/rtbFmT
CRgH3kr5eSxPE50wCDErNBdnbMRxLKwz+OB0jHyZCWLYAYRv0gHDhZ9gLp/+lvoK
VBBMr/oQA2kTIP1jqlJiLT1czn3sYOKfermiCKJmhdSHIxBKu/wQzDYdKhWyTwmL
/O1q27TQ0sw2+W4NR55eLP339mrMFrPFwB7FQ9YCudPdiISIwFbxnmJusRVAaqX5
fGwWEgegKs1zzZ/SOyz04ja8uxEUiob9pqgjKRqpcKGYB97OQ3fWkbYRLw3INWoR
K6NfFBtTRfeJvRed2zevgaSbF5N1abTpFtmj7FC6rQG5ZPyKKmjugigAy/BY/KmE
GDM/wfUA8fyUpve96t9AVWpgaq0wzu8oSE9aspvBT8Jm9UqTUvBleLFqw/CO1g8K
L0xgXkpclbe4OS/Qms+fTW5U4A//UQY506EC+lqIPxlTZK9fMGlT9Tr28SeYcRvK
le4MJjzia4UHpz2x4GOicsY2rgigQrurRXXexymdOSsvqEYdiW52y4ElIjqA6qcb
altGQmQ8Hw8J/RnIB3GRI3VpqkO9t9uvGE9CWoW+3hcsk9HDqbdfHtKGgpxr4cPo
rd3tzaSiWHm1hV1Tv/yLixNFw5S64rkmSI5hz6kKVzfrdE/9bJKVF8gGMz5cpBRU
ZasLA3yv6KGsBhJEIh128qORneUKNDWI68mVXZHuedMvhkeNaGkTqQdCEqRO8eI8
AODYyWrMrcAtDxiy5uA/ghUlgikpLc5A07mDbBpbLgvltyxTrGS7vlPTxUNMLj2B
sZ1BssM9aMMCPy8SNEynZ6RaPej6zBtaW86VRdFaJNwdWAFfmjOlfwHt58d6pAXx
x68v7vxn8/6l4IbL4HMDWf5ehWBtmFXz37omgXSRGXagltiWugWtWmMvJes+ENSL
hyNcqBMvF1QXYYZeFNOUPMtnFY6Elnd9sfKLU8VVCrNg22sEeYx94wmFDySuD99R
uxi8imr897aOtWeJrsjrbjT4DoL6iC1pW64b0xdmG9lg4dlw/36EmbGxqMN3dNwx
BVCZ/jPSsWuy9quW54KucYskGFjxb9UEX8B+IgVVsi4ChXFo6fY9PvgMCj4uaSGL
oXf0mPml+sOOzpBNWqpKafsmJP5a9qjGcp29n8wxV+j2TEL4ivkIFjkBbbmRdcbP
VP7ZLsLBhjdwZY0v031tS7hS2JZyljhX/fbXsWo40jpoKg9K2LUPyq3jiimt8HrU
GWwnhMQvVWp4+xMhFoBKSmmzmr/WKeeVQmNR7OxEgkWkgvJqJuL/3pK/ndfOATBU
KotziVrfEf5cBRehNZYv26UBcsul80fJyShUs4bJRJcrE+fFD0YO7Z+TV76mLDDC
TcLAU7X6gAqZGG3gtnZOZEzOAo7gWElRQfg9l28Tmd2KmMNVnVoUhZk7SS7CiICh
mSOGHbqAsDvxhtbbpCJwpTkdz8L2AYY3OHvfIWQNQ61/MNbF7qpuaftc/TJ+kB4b
nweK6ppK42561ZelDlkEUrjNhiH+C54pekJ7HgJMpeCBSQVbJLOyi/g1fHcQY+er
YBI1o20RfMADsfTcWcyPD/v4E26hFxDfI1oPrUkt1DGYQa1JYo6BztielL7gU6hV
1YGmetSy37Hi4FVxu74CC8str93c9o22eMptOfnMUCAcgYyVbj87cx0ErBz4FFuV
W4QeMGAi3oPkFa7QUmKpmmDJtSvXWt9al+jsXMTtHV/Bh6HTIBaEP02NqXKaSsON
LO25oUCWuqyt0fJ+zYjK+n2ypO0NOhLlVvprOPDETebCjQPVR1mS2xx5x/Z1oEI5
SmdSMZ/RCRg2xqy9UmWhhWAUB7Od7jX5zzmitraaqBExW+GcbxvkCy9gh+3fK1rL
xLTythpcK2WEU2VLIcCl6pjT1KENsYKCxW+bLb36lgPnOIBqBoqJY8HGv5eSiUzp
ot+PGK0wtMOuXfUXGFMDU0WIfDahkOiava3tkHPpk2XV6HiG39n5manz6RW8601l
12XK3uejZLAX8CScUiNtiXlEbRNgrJLqrNzITv3YqS+vXUyK8SWhdgaa+iMSvrQC
guBVauJD4KWkXIxltXwwe6QIuDzA98PdCQMlhGSBHXsaRL/9OaO1cX6S88BN/Ps3
jcdfg3hMZc6MyDpSGTf8xc6+ghlJ6jfloEyedi2bT73LfAj6l4QJE+UsHG3JtMyb
UYaShl9mNL/HAjbfZqnIkdWgCEaRa/hIT48SuRGCIrKxrfpS5b4r458nAXmBt7i5
PDlHCgiIPrlX/XMNR6+l7TLNK8MLmr31VGwyawlZtyJHKKQaPxsUTNme6bESRiFv
GVUOCzzIljElxkqboa4ff/tIideK9LKthLaUm/OOJOFSD0Z3E+saBshdmqTHo6zL
58K5pz37UIfm53Kzm0QtvwnCrOmSeGPRXurrm+fMe5oJSqblC+L3CNDcUab65ahY
a7w09JDt2cMZmJAKGyeGwkUbHDYHhZB5gADTNjygpt/I6+hQKDLk7sMmy7DbiiCn
veV3g1wNbcG2NqEYYWZ8Ge5RU1PtCH43duyuYWKC0B6tutGbkY+GC7F48sz+rh9o
oOUhHaDOQlSn83WDBPysDFjFdOGfDil7KPAx2fa/up+0ryitXdbDDfMzc2+Clnl5
26tG6tJa5l2kR6ad+KTpdHGJ5i0HvM1jfQ45p6V3WoSevIIffrHgML6TP7lpEbnV
JS3ET71Xg5/xAgob3ZIoHUMekmMMiZDvGUxGaGDWhhUz2WZ/JQxEH2fyOWX9iRzi
mBK57+U9awlxebFa+cW/bKMzTN3bFKyXX/fst/rkdokq/C/WY69mMtyKeCbujpQk
Qk4yzZI81EymvPwnfDvW4LaYOnoADHoyu8EiM1vcq7zjvtE6rOmsWkOAbWkyF89H
4w8Uv5mk5FIu0uWAK5+FsC8tvT/31esWre4wl1d4Uf1Q4Cq4RzBypcpzvkDclKxe
sP+w60a7xY/U439NQggJtwVa4hm5pxCG2uR+GTuoABf0pr1usi+QxVUl3cEDDr27
LGGFR/bhi3BM8FfO7OrS4PeafAroq7kyblRfkYfsnIawkg41+CCQg1V2RSsnBk9W
raNcExOkUZI4WDik/RZzxkHDniUGuBKP4L2GWo+Fl72BLhGVekQJg98S3/u89RRr
dtj33WlVl1tbmbtpB0NvidunlRwOzwMtDQ9b1G/hLLM34koxcuD3aDywGCq1j2v4
IuWNpQUi6FmkMelzJ469YNSGvFgu5m4sSsaUKuWJ3aJD33lZD5t2YD+hkPlPMTwk
jHgBugil2FLe4JGmI/hVF0TkhzSIIoTzbPzwk68qakTuEKDBGUNDEfWl3PIK7p7+
mU4G6vgFqMD/Hm0uy//t64CLVXyXk7yIMPI9vPfs52InhKd815mTRBpdb8ErrKDy
rm3aZ6sO43Wdg1HWRTa5SsNXrf4jT0Ac81zuFW3MLVIqkNPD1Dyjly6/H+2PCAbG
4iWRYy/sk/0bqoIIAxWEhTZHQYajBT7VEHIANtGG+BscsBZspx7r7nv6RhAVleKG
jQNz5MsLK2NyaDgAneq9qOtAtk57n3EvxihZGEN6REa/Mtjoxo97IkBCF2RgbLxU
xbTqpxxsTsaqfOPMEvgAqY7r9rxq+82Eax58SHCgq/dzeufNPkl8RnnoEi5BYMzI
qHkIjQP4OO4NFaFm0feqqDfp7bCmPyucbC8L5nyLW9AknyNGoHe0eVpOwRDpxk2b
V2unhOfbSkX+ikAMHrVMqCZiU6G/Kw+UA/9Srqp54XsL623OQNXzcUjStcL/6CYG
farQe25Hyu/0R6zzcOQMVpQX5hWm3m1PT+IGAbwpPvAk6Xw5bdE4Jw4AmWYnu7X+
dXdsZfevyMKPIA1pQtpTQmQv7MfWfvLyStylO/b/5tq9e65eaoAFHQEEwmaldXfh
Bs9IHMIL1pZjTK/+E6raUSlF26KFqkcgcRi5C1ofY2UBNhMj3ICcK+iz/zNtkzQq
/F53jFBMMtH8UhgDCnssv40V4sPAdCJr45gyDpCTYJQMo9YJNsUV77z+5q6xGb2B
2Cy8SlPtMLxjjbAvB6OsKoe04GEJG7aV97vizSDCWH9VXAlSrqHd/9Qb4EbSPShy
zdYEvMYdh5q2dTYTQAUwEhJDXgUHSk5P1L08ZSJpjGfkPCdR4gJNSs49miCGZ5Ei
jlnMkUrr3P+KPV5P9MMbU4UdnyGaARzhDlb73icRUo91lRjkzmuEu2hmlbMMVbWD
fH5Dt191EmbQAr3/fD0tlsj8ShPV7cL7w3mWlTQ/C43dUw1LkX5qqOs9c5zeSO1V
ahlLWifX60Shis5h8N+ZoPJuAowCLfETUiEVHb4PWmFbw8g6V97Zi4akr6nf1rtK
KjpUVpjmeK/TLNkSt2S2RQjM2CwIqkOxq5YUYhwcmvRr7FC8HsFO8FhJmGMBokUU
wymbvI1dQU2vF7eEN+F8SqJsM8jjrnVPpx+3AAPRppPQggJgTVy52/bMyUraxjfg
FkkerQ4ymmdJrdPekw8lSAIG7EieEUYYqtBs2M7kJmwLWEtn9kN3NsT91vlDfbbO
eiznMPEx8HatsYNdXw5DyVXPfZ/bsMIVqMbV+UpFXaQlnLszJRZtoxjgEjPUNpMS
WjCtaDIq5vHF0OjbdbSPzgX+6fkqCLmre/bRBPBrDrFJkGeAF85dTe6bGZ6vTs7K
y6n5VnV03GsHyLgYxEgxHpYChCJpEjMLpVPoHRn355jG1OMf67Ks91U7D3G2G+ZO
EZuyktuHHqW5WqTf+8/B1Wg41mruiL9s0Bo7NCmywSquwXsTAQ+i2Ss/Nz/eiBeZ
eHrcW6kMLchCFrY1skEqvRFu7aSO5hVEhsQImQ2MhfidaEvw3ulRJZPBUrCKuIhY
vyAeOqWMYhtgkC0NR9E2dh5SfdZ5s8zJC4QebscMHhLO9M2THyK/Of4kF9Egxxdw
nMSwZXuftR0+QtfzY+QD67qjpCfxeWVoZp2Q46HJAMzh13q/d1p8J1Fh3ewEOUCS
G7bIUpxchYl8tGqEUADu3nK4t3iW/Zsnjjo5luSDpPunnvALves+zyD7x+P231eB
0fK+4A/pi1YzY0DnkDuU0UOyYBoj6JYUwu1/1c320BUDa2tEIjUYC9j+6avm76Mg
gMRmP1FrbMDyOIYPNeKS+QDPYvEgZv/cB4ctchklQxvG96sA+qas1MVaXa5rbx2A
j9s21sS/ARUQ/H0cpdYjZ9RSKGsxasQef3ViYkR6JUp6L8L1QdkbqSNaxnlbk6h1
9wNLvb2bd4VbfRuzBgk4TNTbcmUv3Bk+mJyB8n1VUnRo+fMTmQXaTb8lca6ytfwJ
GExg4gCXyfG+73NonyGenp72iup7ytV9v0XmgmEy8TFCUwnxHtLuaK3OP3L+JUhk
LXcm8jnJuVrhhSCgST3LTXfAN5W26GvMdP7SbDymFxrypZexo4wq/vIrCbxgREgP
Zauh4TyAqOVjtL3MaDU10zteOH02V5w9p78SUJ7s5gILkQoU6ntKZIuSJwU2qfBU
azdqTeh6N505VFv/fIkUd+n3fjfPUGaq+l/pyXEXwb6HjmW8rS1GF//eU/NOVNQH
zcBnVf5QJ7Fdt3+w9xonUNFjP6PcWAE+ggIN8fBDkqGn1XKCG70RpslcN9Iqayri
JoH+fHu9mads8v13o9NF3qnOuF3+sf2pZPTUHimWJUs/PhZOwVihJ0KnTMOtQCUQ
/t033t2WYF3j/QQc/KUTgzpDlCWE1yAhFDlSk9qjWEG/s0xQoxsV2XTVlBuF0KX5
M3lyy1bV0t0EHSAdwuOOlRmDLhRgE9fIf9vRuWrG1QZlLGOTy1tU/chOFco6A6i4
yB/0thwRQEjfFjWl8ckbsov+NvGHa1aem35jBic3jAPiqZxE8jaLSwAyDbl7pP82
2GWYKevke8L8L2wGSCqKSxlAO19RWtRTWQVnfgKxqoZ76uAa7DnOV2mhDKlS27F4
7rxncFVmnq2DBpNB4H61GySB3g/oAoGzFxgey1QZwSISXnEQizeS+w0ErmHxbWGn
L5DjzyeuzX+ub1JE6D9ziZZhoenG5ZRZ8kkc+rf7HW7ciRlZhKECF72k6/JTaz12
w2LiVQ/jfRCuje/1GhArf4FfGvxr8pc49mgOqdfKmjfm/c7SmfLYUalPMXzNFIAG
dSmSC0n6z7At7/kxHbxYfAaWbDF9L+rUQYahkUPk5cxw1fL1nq7J/jL6J9QjWoIQ
v1YthdCQJozI43Vk+CYy9LpsWGS4Aw2C/00S+ucn+xEwbItGWgEowhH4Uf5eZbME
zQ0VovdIAwBZp4z7HCgHta3z2hsziUXmANfrjvibFlbh0LTOHYwBpJ4j1hBPsGkP
/2ja67Mf32ySSDUYf1dKTcvAZI4IWPLUF57MBU0vrzXFBPGU1v8cIarwQASyC9z4
+LR1imy/F9DkHZ0GQNy6+0bkcGyIOC6FQLG10q+cpnP0ztH4/BgEa7Ubd8gL16a1
g/yk2LGJJHucHfSSLAKeBxPIUcQiJl5yJg0jgBPJoAHWjn2sobcChS+oGqBGased
54EhY68GodLPLBjH47LCPRuccTErJFdeIyO4vZ1RYD+0Sd50P+pxsLKjyLH5WsfI
s0vW4MZjrzCYgSlu5HwNbUbI9Mg4r5YbiAnLcWC2e2P4CSIfH/wqU+StG+9KGKgp
2rAZj5fYNyvzzezJ9eFJSnoc8dzn/x55M31JS6XXJOTmj/XUaDS7ydNAhd7D1/A0
7BaVVHUEvUidpxj6F8xHBNBs8ylaJ212ZLzzkXknznbxN+Tz0iq4b3s78mZ/h/vQ
mh7U9lOUfjXpQzNOkKx3e81VxE1lWzNmKdgRiEwe36VuSBY8lH+4SYHS7Q2294a1
Q2VxGszP9NaL+P921VdNBQYweHz4J/ZRfBoEdiO/KkHji5MtbkUr+WOJExM5hiKQ
SCyOY+2lxx6zzEntKNagANkHpzfqFlF8n73107qILlQog3uTwz3muwO0GbbzFz4k
JiCKN+LVxfyfezCCyK+QYEE+IbUsWjv/84yxOV4dQhXJKrbepIJ+pi/RQNYfx7bc
2yJObMo6Nu8yq7M/TKGC1VilzoGxZhyFJSKxtnNbbz0oOi+qjEblrnUMKek2pTbf
WqY7LNNeJazmsLnUmrRJVROzmdqjW7e4/PdOyrFeGvmTAbBwERTHBAFRdDkgJOBo
ilSuP413RvWPqrF5kOm9eaf08QkROCz51AIA/kXivBPOKF+H9JSTe5tLNHThkdlJ
B14lN8L5Tda0aVUjSgTqNzb6b26r/2MI18tWLHnRtZGA4mtllysDhZed3bgRuLNv
J50udDVtaHF/61lq0s2e2wtXXtbviJbewtGmOc8rCmLVO7rnx4qbFcdgN7QDSeR7
Oir/dcOk2sKzA6uubw7hTEYUvTZDPjiSW7FGrSLYQvxzRPRKsmcDTr5art+00nSC
BfXFslp4RyrEYlCXCQWAVpRl0EpBrZMACoBDvw/yrmB5cv66iFvvdktKFnpEgT8Z
BObWgzdRZs16JhcY8RvFZO1tvHrTpXstHQrPpgMCMSM3IuT93DMz8Lr8lsqh19EX
qKMHqRa/UtlDaCdKEBH2Ks5Xr14o7lYSYFMR/JxI6XwbQBwbsK1Bl2roJOG7GWKm
fGZliCzgVArENbSMwDMNFlXCTAAJZf6uy9z2WJTuKkJUvpO+TXjsfmPPTPkLdn6m
1OE55OuzBMHf0NHDDawZBcVPwVXR0RZc2xbJZDxuytjYkBCz6eLV0oa9xIGB8hcT
Yabe7vh4ZqlwAD0OE9shZ0shfo3iLNnbh/+pbn7cuadTRrTzzP+mgGCzZaRatIGC
swNlqUcNXYq9j9ACsMU1SyQbG81BbBoVVwVVhYOYnqaj1fwA+f36nKZVlrwqRkuv
3uRDlmJaA1GgZdGrxToPdv/0d3/XvJADHnvUoh6Pn5gKtP0ZXm7UvrW5FWEyCwZ3
CJaDHdiChbsVnD8h51OPgmOpHG1UZI7fHjLGj0sqwcl58890Mz3AnGCJTYtmbElX
ZPn9bzeBJ5n8Fkdy3qxmNoKyhOYL9F3szxQBajsPTNxHBLtxbcNxXKQ7OACbHGcW
8qCZeVLlebpsd3qFN9c/lbgnWavfVDp77nspchQPsBajyX/4qcdGxN3SYZs90E+c
U9JJ7U6/iC+kQlDiP2xZ1QVhwO72jH3VhiKVqOsf+vlD3rSDS8NvOYhX8Cjn4fwL
rdCcSIQeVRFCC7myzdQFyfW8PycJBOSrTl58PbeFcC0ezTyrc3jHWhYu3CiMNZRY
NVrUzhURDVUcXfbIitRQ8uesk4+rpoyV4RizaZ3DxLM+KjwRGcY6FE/wfCtVQ3Qy
XJE+JqVd54T7Ul6DdQqBCtWU+fhYEbAMYS6w/7FCnE6s6ZnuVGIww/yo/G3iLaxf
v89l+jWSMiaRQJiBVkpFKqoyzzvdeOFPcSVYiRPaPbRmsYuaZp3zKADCp7pxs5VQ
H/3adC+r1nd5dPs1jlozMAPDLmD90/WIGqHsSTC0oUjgCKOTO/+dNX7lSRLrdBuu
fMeC7uHrdjpmZs35K0mDDZ8OvRvKk2JwHZ1U+rZY/NGh6ZGLHyEm+W/9Qwg7Tz6y
BY0duq+MIa6WuKVOEwSwJaAlrgDUDTe01j+c/FVH6MFAidhUquE6HUAvZoIyhx5Y
VanSYwuow+ZrPPl8kZbGoalk0RG1xnRfxxiGT+K2ngvY44sOH5VZZUDhGswgcjcz
1AxMNdvIXYJtIWXm9MpGOWbwKZhUqiXOOHTpdnJkohjojHGuVx/cz59ZdUYyXe06
8pzlz7aQcz5J6IPgUCLYSy8bqOeRbH1sidSWiql0uSXzcBVcfIGokrXRkko15kgO
C3bu+pfXk8rPvSDdN/C52AIvC7OL5LKDwZYxVqOD+OcaggnEYv9LkZqwvT7TlgZV
jKdOzOfhKpx7tVs91y+5F6MmV3TFIIvRK+ztEoedwhkmzZyIKZYVXIuU7C98pQ34
Vak4kj/+D9NgWkEb0bpoAdYWF0lXSo+zSdrXZ4yq7EHHGhxJaiZZZX+zNCT85WhD
YQwH03ozbMRAdwp6gse6T6tvci5VqdeF6loXQvInoDSSlihact34vacDhfpqCRWL
Qk90aCbOpMz3dAOdK3KhBEXKGj+1KgATACEqTisFHzSBKkQF3k45in73Chza3PA5
mhQjr455avKyr3hHXY2zcPuOfLWM5v+KJECZvR6mPY5bFpiQxMHTVsEDN557Yrvi
nz8VQoQNEleveT5F5wuw9Qfurp2ydPObArIVF65SYPS/MxBB2iHon7VutBU7p50O
//FaQky4GFKf07pjW6eykpL9JSQRwstncLCcj1NpO0ZadKpVv+pdXuFmYLgTM/JB
7iVyjWPxB7EPwB+MoM9JdWCtCsaPgDm6QPhbz3vzsfJh8eAPyqM83F0dXGIs1HSM
ePe65b9vpZvFpizrxhujMjaFUProzFxYvt/wnj1WTxlATjjqiW3Z3MjLn6DSBKqd
/Yo8/d2cw4eoYS52TEj+fog/TRKYnW7CZ3F1aZr47nZCMTE78dD8cxG0wZsNj1Bv
0WKxImhSRRdB7Xh0h2/wGDZVwrVWH0YAikZxSGt/ZJlB0+J/e0b0Dg4F/CxlgVRT
YryqaOClL40oM7dk9Kp+YlolXFrnDYMKXkoqW+o52i4M9DryGUrqtFEONjtVJ01M
uU3NVzncoN0LC+tbSFbHAJMlAAiTb7Qh484ys93ZqiWOE0TFkWGLB4SXkneJzMsc
Cy6aQ4B0nztTVs5WX6YVaXYvpk2w56K2UYu0zxMFxMEjOjqvPWi/wRWBlO61xyNS
Zh4P7JvDnd1GPCeLuHxt//ZE79af20RElj3mI/NkCg1L5qePDbMjb0orpsC6ftnZ
gc6wIcz7KEJ2wYx1bQXOYpRIgBjc9jSPLcTA/kek2O6L9a717oeBy/FNanSmMiuS
alS8sAA/X3P1lW5MGJcGNnAvSCMFO+/tXQ5ReLvYREHeKJTefg1DD5ujaQWBwQmS
F0YgtO1l0bxNajmLVxUWnTIf0jhFxlnDZKsHxJ+IvKL3rYouZbsDYPmaBGHBv5ic
2EAMwk+03ittQ+Mh85IwSel4xFAQjS4Lxk8dV7Ao8SnwBhptl7JvNrOpI1Q2WYgy
BozvUCjZrVrgeNL2Xylufnb/g8Xr+ARw/toTJvm7BX7kMPwbz28QZ3g/6AmcJGPO
FA0JPWsPBpA5dcg3r6mqYtOSblcJrnz1JJ0JW2svpv6Ab0nthT50oy8RzM6Iw563
bBBXaFK+0saDHJ1HILlA/fd3apcdiuW3u3XxuFK8biRjUBc6XngOoGyTKVkjLfuA
qEkTQaG8Y281D5VX2wXah5Py/KAEL0ThCkPosCf8jS6ePorWFR+MjsBbFzt+FtGx
cfUIs3yDZQ1SuNyrBl7w/K/tdbd6xwFZGRYX3gqrcU11NCeGkEOTkENEDrWikgUF
upMYd1Cog5QTB5+RJmqD0FV3I4gl6xc6q9Mz2zaP0IwxiHjGlek0ium3M+Qfaha/
86iOehYsVlT9+sjEK46hE8xeFtVnuWc3OkBeVarJ7KnJ8o3VieQf1wnoSddEhlKc
KXADb4RuVeIi/u8LdTPXSPop6C4g8A6l0t4nT2cwcGHu8fwGEC0y5hfL1yv8iWtO
tz3CZsC0RyASuYD7nN6yrhKCvn8QBIbnNX58wDvl93N9jpQUHnIjrqAG2qFfRV8H
2hC8vC25QQ19CT3m4HSBPg0JGwZ3xgcRbRB1rsVomlSSr42P4U1bHezp+r128pn5
q0UgnJMbWMcCzcPZ3k68xcgmVAUVmM3afZVVPFGJypk1NuI2UXD+fpfaejKb2Ofu
Tk3oSD4RImw9pI1pN3C8LJJQ6KbzPI3LQVAno9slZCbYkrnfl/mTvLyofCWL+2iX
JpDGlkrBF6Vgv/CBbNHpSuAlo63bUHgWILzAk+gXHNepyFDuQBeOA/ECrSyjl7FS
oMlaMoNxPm659v9ixA5Ey6zOl55QUP/iShFgo61qSiIZwmAqErRG8SDqDTyHCWVb
rn8XCNsYreSGqbkZ7mGEeGS8kj6k0VpyO1597aGg46kEzi8k/SR8VvEJBZ99Ysdo
OJy1FhRUuOWnOCUE95pS/CGLc/XonsyFY0nUY2mFBNmNaawQfzB1vynZVsuy4RIF
5cL0H2wxnjpmZvUSB7VZGHoH6H+8dtXcTgy+aZXn6BLe5ooO7irnJYvp7/04Rayi
/EHYAq/LiGqPI2PVd7twR8JNeqVJchGjYg1gYoMckFzIU0PdqewItuedKZ6Q0/64
MMrC7k1QMPT9o0f76imm3mvXYGTVbMpuR7/HWr0e5DxvXwAJV0WEfHBJLQA1yGDy
b679uTGQrTQsyur1WSTDB7+ptDZZjBZa6UIK+t3Umbn7QD41UFNBvVHBpWUR+LdY
Qk8mTbiXCANrRPq34HXIdVt1uRC4ZdE/Zxw/AUBM6IasjJLpcPbAO8vXSTAkPPAk
xWcTw4UzDhTpWN9RFXIBD82Otw6nNs/3r5npAlxUAI4Zqs7hEztgb2Aj1bklef13
zR/6KYeNB7qY/r+Di7tmJjj2bSraAIY2S/U8MUsUQg4v92lCvKmqoLjWsp98Y/hG
TWv/FlukqidDa8n5rAL2nVV/hORh5s8V/j1wtKYlbHXmtb0M7RbSqoc0WW1uOylp
Ef4331JwifDiy8AoFG1DIPkbGXvNmumDOknZy55RWxn5yC2+Pxjxvkp3+R5NceD+
up1CQ6CSDprdOLQEICEPShXD+laRC5jAgJ8iIHGZVFXowgHG8clBlbyhnbioEtwU
4OtzXRxMfZJMaVh1Il2HA+Q8+tzbYtXnYIuoWD7dc637dEBTgnE1bhkOXxOKpnkx
1/Hi3unDn90O37YbhD0vuGCEWo0lKCelYOU06Vo7PWH0ovfTgU3AepYnejNqUzut
NmE2UhkhmxSMqphBkMlns7fAJZkTE5ncWfJu3X1B6y3s0ClDCWDph0lDd9eTP36p
bdUTm7ILqbeXnWwHye2UVmvXK/XUIITchQcZYdb6DiGor4Va5VZCROwPzqQDc4JV
+9DZ09+yuHdW/oD8Q4G5TIDM39pv3OR3T0GGkGXL4pFWAmOm4+tr6MIU5rEu9Mr9
9EceYeC7VEZhgTfst2+QEe5hP/lhRiX9rCsLY6YEPCOMJq5Anccm+200MD7V+YXl
9Lb5vqz8WKb27guQCq26Ls26aDmjNRobdxamZUre9DyJOCqLPiug+c67cZ4yktUR
huqEt1uKcGgJYetPamCaBUyuIiFDkC7U5GDf8oLkX73gJv7ovJCCTcmxJ2C44oF5
MQRWChOUZezoefBAuhRMQa3pw1wEL6/YHUXsDpNqv7MENX9fhSmvDtLjzrcNCxtK
ZC/pQEHemRu0OoVeDTU30aDx4Hdo1dl4Ry+ba7FABzqi2LwtkTt7F+tl0ZAzMGTB
5I713+S5BP5drSKhyxEIKm3dNDwJqzre8Yo6q4Z5Q8jxjXom8yhYau0HbQQnp23A
qz/+ASazjud2iy7yjybkUdAZNrVe7Kdu5kjg/FJhpRHdOxw3VA9JjXmtmibZn8WK
BW12OYR4hdBE7OCSMOAPDyDQTA0+6PI5L/MnrSkHQFhVMUUQZUU2t/D7S1/wmYuV
pq4fcBNJsx9HjbdUy4hNNlN3SHoszZCSbydTZ4bQtsD3wzYdbcy7lLWToVd/RQVb
d4wzyEZ/CVtDXbL7BOElJ6vthMtB4/kSP9x7RQ/xaJtHWa+sEAVUALncvg3fUBr/
U4XT2uQnbi579iTV5yidKMoN1zbQJVtFRWhZcnwVfezjQmZGQNj2bEn52+SX2RcF
6Ud4f0oGb3s9tdm2fVBtNCMXdXXmLFzAoD7124Tu7/OZgDgaDwDe9MEizwbCM1U0
3ZCRTQJ68JoUkfrRXGE91TJTX6Sl61zFkbgPYeL8aKINHqPCZzBxwuDSFEKxPzj7
6EwYYIVxfg0RlGhqIDKFX6Fl77X95U0/fbl7IMJMsz/MY8PlwSIy5sD8mHrOoMnl
1q7wq65FjaiyLkJDQN/T60HtcWwyN7w9t9Q8CqJGLNe1L+Y8GOpDJ/QbnfUkK/Cf
YRKDWDxiWRRgX8Kn8g6azJma/EY9u9rK3cSz7oPKlf0hiRJvCrRWPq5Vp0b+5QHa
H++n+QgOguci1B2XqBagWk/VqBtFS+eQWh9c0KEeDkYCTtcwWNOPFcwy/u8Qbjbi
N2f6MDKsgR1xx2KcXk1g4ALevv9mKmea7wLYD/h++Xcfo8A6ioU8tE6/OFq6p3st
1CTK2jThCoE1J/mh1l0I6bg+leisV+hLMjVjsSwQuU5DVwd3LXzfXwV+vxu/RbxY
KAYlsuaXux4J59i/jvTwoqvxCN72Xil0JNeRCxh+pX4eIKldZlLU31HwSptC0dkL
ZUB+apJJDFQOctTQfy0rnMg9pCtm1O+6G15SORlVO1Q7CeHyLsWC10qfvFYMjjJk
PB4wTk6jjWHs3bpIe1z3nOindq3WJBerNs1mOri79gag/urqxPUvFa7ZiAdnOFAk
7HVsI+AQuxI5DI+JiDlwZ2OQR8ILLkvC8K7mz/LdWX4ZbffyLzCWAFCmtz5s/cpt
dXbIStaaT9oQiOZdr2EP1a60vejHzYskQ8/wv2au1FbaPPLaLVdR1N47a1LjyxgH
pRY3texduywesaIuPiDMbB6XWCTDUvTFLt6JXCMQkAwdTQLHvK4L8bd2wtZW8mnD
SXGZEpLA91xyH/1nwyhXQcejDYkQ6fW81Wq3ShaUYXz7o5vnMpd3ns+wuQkjOekU
Y5+OIlNja2lN/gD63ydov37NMFH8dN+yVf8ECNKr7AdZY0LG+D+msOX5ocKfaUD8
/a+wRBqUTIkMW492kL1HFJQsqevMS3RywKgXBcYXrXt2jacb1sl38evM8PMwRCKv
6NDB7pa1fozDJUvGr+sHceiLZHLwFKqz7aCcNL7n541QjXhJNUV+rxkeOEjdecoG
tLPfLqyqk1WqdPjoOib/ALMz2qWF4rDgQVLm6j5A/X8BIPdCja0+Y9z42P2KFMBc
pSzl+0Xd3E9iONM4xsELEa+/Eb6rP++sf8Tanz7lTt7ZIqujPZXqq8meF7pM1k24
SD/8t3ilwXoJIIotxT396diq5u/bJmWRI2j+lFLSDtbc56vAmctKsXtJzkPxKEYM
x4kuJ4+0P5P1/orxhTJ7Vi2k3lUHH8qoDUUyhh1LOB6AfWZaxCzwn9Zfc5hbCvQZ
OnmGRjxV5tAUheOCDVQUF70UVT2FT77RtlgTWKBYQV1vdavPdqs9Sirga0UFP/B/
rlpyKmWJI/4UTDiCGygZHp7RuDKAGK+nEUFD9mqe3QGUmkZR3YS8CrtZPbuZerXJ
GOyQN3h7tY+JRFUZhIZ7Yp2dWRJ+COm1+mY0lS5k6O0gOP6xU90w/kCtexE9fLG7
h1OADW8FJL+YIB+P2883Op0GlZ0tlFVX7113T4BQRekMUhJOdMt/mhyl81ORm1UO
1thQnX+XNRheTBA/3I1H3Cle5wlYvdxv+JR5K6d0WTNeOQapWgu8tEpSmOyMMkFW
q8huT6cyz9iIju7kcBWi6s0QthP2k5jRAH+lksdetxSVGD7duVT0vq77oDRrrowd
4zhmF2s4Fn/cRHbw7NB5sKMjDyyBg+Q8Gu0ZWK7b3ObeXsx5kqJHdTSsamoYvpHr
L+WRpfeLB+Nhl+paDsHPFTCRkVO7ymq3vl19Nv1cvo2sRve9JL6CgSD2g/cSDMJX
c4vI5BEvSHhpP3n4XNv8RbnF0dG9FoogHBj6zzz+r9O3gKuICxnS+TuoceFduEip
+m4ht/6hpV/9xaQBtUFK4wI+oMArGPJ9W2zn3Nmgp/pHkf63FFCqcqQ1xfdlJ6TT
aWqO/HGzn0qbtHauqPbOtdX1XOPAida/n9b/Hm9vDtEnDMMxSnaRTpxu+xs+L37Q
qTNyD/O+AGotQBDYF6xYI5ApTP2YttFikfYpYQQCRLwKqwNds+cJ0x+dwjIaqmG/
Jtedmdz5xItL6PwyLjwMWZkOsYFv1ZMiLhEBdbUhU2TgqJCznAAys/tkVNXkqolJ
Eq489ED6SX4uNetlWRsQfJ8RU1/wZiKWhAEpZbKYc1GQmkTcRik6pJFE3NCObeV2
f2fMgZ6HfLRSskbewlj9VjQR03orNRmLRZUMZwqo3pxybxL7lKsyKeDjasG0QCQB
oNP3BSCg95WX/Vo2+7pouVuql/vQIGQC262W/0FZvhilpucQwl+Fh2qT9CAuWYnV
uxALor84wjCYUFVu+WX8yf3MyZItd36pYn4AP8PPlPXH3wvb8RhK5mYZfUiBWZG3
pIUQgjr+rsVdOmAlkxWYbDdkyrQb799KWV5GEhgFrr5WivOTUgM6WD6sQNBfmLkg
HSWrn5z+LqTVXjxXHVWOATxC5ffwmawJb7wl3xdwHjMuGHQ25rRl0/vOXoA1BjYc
hCH1ofNDoiO+vy47KnnO2I9kOIDExrStu5pMR1HHHvWrIow3ztxKK4r6a7e+QkRw
J2bL6WwqTB2+TnYDAQTeNMp5I4zpLn1VM7rXiUZvkJf5Ucfqe4uLKDonCXzIm0TG
ZAjUrSUaXhQNCeYZMxk85J2To6xJpUKx2X9pabNj9Or5FBTKIpKgoQA68w92pqqt
rtYS2nqDTEfngb0celPJK77AfK/7kdUSkPYDVgSpDN2epouXiolPp1GBNQwrDkpM
NXmjiH4jFMfMTo6FoFjjA5ScTEkukBQEPxcL8R4PtrK+HNoSL9zO1xL6zpZJfj8p
M871Vjk5mP03d98u+oWXQdndz/W1YRyXadtqiTQ6ooXYqrKbjliWULVHEk+UQTvW
5iYh0CYxYrJtO+53fgLg+VbdZn5ulSzgHEqSLeKL2gvE/dx8rECEIUdelfTqrFBu
o8Knb10SP1YHkH7yW5/c7OTVqArrRYQwRb7HC6geDF937DQiDqQ7OgwIPEhd1CVK
K6zIpA0euxekALNLOjiUQYUwFBzJQoipAckfmkElF1x8nTgeIVMACU9ZGlEdgc7d
EgcQsVoRKnEAcanAJLDro1nMS5AjWwDuEU/MiSZy1al2rwkpu/CijJQfA1kznklX
u3Px9mkeTmmdcV/IyX+gyfkPg9iWc2bWx/v/AVmb+9cScO1d/dA14A7UHAzh8o5J
U6qwJXAUlXHtuXC2yqjPlVmspHvw2XNz4DFm1OH2gp9YclJC2xirIHcObRudZtre
+2erMYCWvNWYuTYd07QKPYim3JII/ljlZY32jTFEl1YgwaGfZTqszh+jwtCkF5E6
8W5e/y6jkpSZboMw3BeyPdyg3DEo3BcwIozrjykwkopBcJiCbczt+P7IPd6DDsPm
j7QG+uvj68wskyiwYLn6Z390HgpCzchbPOXunbxDbKXfHzABsauFx1XtX7MI4GIz
z5/IOwLgPMUAz+afz5Ffq7PJwaJTynwcU4QgE68DU5ORZIUeKDFmy+H/saiQp4iz
THxf1giLU9C9rPfCjxy0x5nRfSeggAB9lgP1N6vOF7c1haicSaVErM5k/tLRbrCL
u1W5YG8kvOUwyvQh/xCHGk6mptUgGSf5/zA10gYdQWKy2DyVWXXg0FwMhE1PJeV2
Brf/rW8a+4DzSlqtGx9Wi2/Fe4WBihMQ5PhyIfAH0vmH1hdJANKqedp4mvIQBNB8
E9hKkogQ7g/jTMcexef44Q3XpzVbzu+4CW2NV1D375wyDMjVH3pwzOY9qKlg1vmq
o0Q7MzGOnL18H3+kuy2BamQRpMZEjLJjZOGDmKP38hrf7LUxB60lbTdALuBkogPE
eMsWQRx6ZQzNF2Ua0fdUayk8kevMjfm7gKZZdT8M0lNPHjfKoGtPiV0gTm52/ZS/
766CVHOGngbGU8zzJbMpo1A/CSjJ77yhH48wpkf96MWIyrS9m0M2/fZX3yBKK4WB
lZAp3AHRz2ki4ndzrRQzsmJKqqxGnkpOqSc/hSDUKXBWaO4njm5dDTWkS/QzZyPQ
1bEQ8MJJceV8yxzpNL6jOnxqTIERDFgk9Rk0HlvLc34g46DdV7j4PpXE9HoOK6SA
HMIU9u0IimqpLWGjZy8xnaRlztsdSaN8wZFEjx2VH2vSn/NsBV3QfbjSP4sQkQ23
UwSphK+JAY43+d9kCbQVxhbfR/912+qsIHy1EMd3rFYi5mxasSKAE1ltlgYIy5sE
v+ZD4Y5UspuCwMqOytCFt9hPAthExwGZP2EsHOKctrzgfB+2QUV6xlkJ7z0/k8Io
hrHMkmn63+CMvdfYk+d73G3HaqykIHh3d1y+QgnyAHuf2uPl60WOLfEoJFfMqfd/
JGv2ypQfaQPFoPl39mtiRHra65bRm/6BxBj9fKbQiQQN0qTeFWhS5MEbVPWhJlSZ
n/+a9wwiMwKhpdMHs+DxPKH9W9CSrbsoAtVu+f8aPPJZbm6NVC0te4bt9faURs2t
fiJubG6Hbpbcxfjsoj/M5WXn3I8auZUCvpqGnrDA0Qy2GuxuTlDWBAGtCA+5RweT
+BIHXF70oQD6hE+9pxTeacYZr1SAXap9K70sLxXp5RMEG7FNBXkAH5k28/PlBrI3
DaNUG8U/2mzx5f6iThoPoU3WBYGU9gAwr/MyqPEBlYrYJe7rXk3MRdvEodrSWiyT
WIzk36PDEw0waOIirs9bjvm1Nlb40A5WeN++/ERyKNKJBn+zVqnXDv8sUX0JfOby
Z4c0RaIi5Ora46SMBDuGCe/NRTbf4PvMr288t55+UhVOlaBMqaXiqyOCHlqJT+BH
bTSAAYYoJkT+e9/oig4Bf1PbDtbTSLvOKEeXrQigE5aVB9LxC1pHCLemHmA1cQeS
t6TWFIDma7SE5OSpPIOmtlXYD3omc/1OtVvnnliCATTCcYpP4i0aqlB48UhMeQ8g
0m3fAfGXfawFb2TjVQ1EM6DojZQjf4uk1KcoLa1B84WAwYIP/xsgfJ/RsBpYwOdt
ZgWPjlHoeYjtfr8xyZzmbRgYH7+voLyZewengmVcgfd9YNHM5gTjAZggX/0mPWPi
lzaxi0ycAJFN6uj6QBN7xE9zrPFsx8h4pIXXR/DdFpohBcJ+TbHkVNdXsAfOQ+c0
ncT2G3xtScI6XlFAU5sIVMdSznmVy4yewIlJwpFmu84HK9YBWwv2SA4ZQOLlraek
DUcyasVVWBPsHHLsZqCGOBYb4r6ht0zgwp721f5AADJkKp/VXt5+EXTUSACZcXvT
I1rkHLW4oKqxw/GHHtRvwxo0lTSYNxgimo6t/YBs3cYHlSDIzcdl0ZXLozKj+rfH
a1zxKniRRT73l0eCrVhWZX6jDin3wBFxwjbgDqeYphkzOunBYB/h/1O3cxgjL0rf
F0XwzTLzgZ8hUaazo6z4/RkXEo2krGpdHl1mIbx03BwvMoohKvbgl6ADvLhzxv49
xJUNt7T11TI+sYbc7aP8VS6fBaIjfvcqBXEM2/yIiwfhd95GHADiXPnRP1jN2x64
FXpaSD5kWkFICIbB2azxcH2BnJGvkukDaPaZbdxsI2P3SOTtDk7PN/GLY6p4usgU
Kk2lKmhLPIPvV4va0VOCFLBY078BMtoH1HqhtSuv4M0Qz7G4rzPzqGUxV6I6oaQp
B9+DMB6Zq5BpucBY3KXe/vTKfI0rTUZNZ98mWdVxNXiQ3+8mU+O8ekaZdT9Om+av
rDDR3rGfkxXknX1IbyNoCYAnhmtAOHdK1f1U5uhPYrTCva2JofLfVYyBUKGfS0mk
1vWVdiWSUYgiDWLGCbNOlLORC0Abwyv1gUbRpM1rFGESEPd0YvjQMzH88gLTBCLQ
ZOHtBcb+XPfHllwz9tfAq3VKqO3RdZ59qmGCMiJ3qWSsFEpeQHdj3IoNgkZD9cSG
mk9AtjHpWUQJbJHAmvEJeOzcXVlwaPmL2inwHJcw2jc8QQtSjJfT2uho4V6sPPmY
cYySZo8Ga34zmG5xoR2LxDsX3sUNMASHQhDSY3BaOjivWxjhpzRX1JjAUN766CsN
PRZiWPzBsiQJLUZ4nTTbgX7g6/zW+633LXrrw9IfkEV9nzTNoATv4WdXhs7vwl61
/Sk36nFqPhHpADAQTWIAPBSBnvdSEnrj97WBo9f57IOYASL7FjMpCSLweSddpDWu
I7/3v7z8vA7hKbvSEVwzEIaO+KpM7w+y+tMKHdz7+OYvr4mVlb9R8oYOSvBzViVj
OVLFtuhs+yIXclH4I7S7bb9TkGyHpZIHUOBZC52uNVx/JktPoSlN1Tn685OcVTAB
tEVq/lXKXWcDL1nJAw3M3weCO93X9cHH/8+//+xIMg4HE1P9vcQ7aRgpCas+Qkq0
uz6gyc7UcRr25K5wSFb8W50ltChyHH9aHEcvhyUQ1b8xDnVBLyi3OZ3JaF0Du+q8
tv4ahTYZBcF2Wgd5q1r+jcAcPm+zTzUg0dUeBMboAArbuJ+yl4ikMufOxlGewsyk
lBpFZXkMoA3pXQMwgoESGRTHHJwBxtBXtbbO/nrUHXV3IHwEHvqM5hVsnUNhrBIU
W/YjzzDByGhDa/VRawacBB+NC57ShykxYgZXu0I1ZViyVnq9C3RGbDYC9AIsXybC
Piq71q+bqYsv3RPZPdDS+rrecPewGpVD2d1GX1GILMTNf3Zpxh00GAfz3/s/pdxc
YpzWVmtN/eoYeqMUQyhyBZzN0uGLoGRqvo9Ngm4WvAeRbdi+Z1fhSd1Egv8fvgi3
5j6p1xEspNSHixygA+f//KI3towWavOzWe1e41RkR3Tv6AfbxCwG5sPgXPctek4M
Ywtg1EWrwpG0ZcNhQ9IofBSYTmPKofUBZaDqsQlE63PoipFpUPDWTEVi1oxXUhYD
/6Ebe4uvEtIWqKwnyt0z5OVrbDROwvddLtB6GXhXKIRPaQ3x3AYhuZ4K9Jq32JgY
xzVyK6BazdX7GedyXp1wa5vD/EOezZe7MRXxppiKWvcdRCosC9mQ9wGym6y8MTi3
c786+XhjgedTD9F3B+SxCbVj557O5nHQ9Ys4HFhF9symipSpe3ScB6O7XOoTalPH
0KliBiuBQf1KxiKaQQURVW/j1L/MaPy8GmtQFNRh79MGpzrjrljIbE7q5wR2ucBV
RfsTOHwGBQTyrURyEWHwCgSf+p19MgKr6hDfhFmo8CjU+T6e2s7dAo2GJUr0xMIE
yJSHoytNRkuPuarjU0O75Cin3t6xEzi6PVduwEULkZxEdKUhuFRv3n0mbzWcayf0
g0e6bnx9HEDnco7co5FSlq1GjT704XmOZuhW+zuebYGQ8z2q7jupREEAYWy5H42b
VRHl8F2OvoZjbTxhqpiNZTfCX8EMxrKf/5UA1+Jk5XPxPnYOXYTrqSujfEPO8+C+
siSRjiCwIJ2BuyaW0JPIuEHvORUg7gmZNjU+Nbp4df+yjDKkbH0D93wtMIdFHcYz
ioc4+MMlJH4WpKWOy1sTO3PciUKWlzK+hAmnAhtZryfxXm3JrQzzJ3eAetGNQJGx
7lGJnetVl7kAnOt2v0o/WOX9HjhIXEaI5JvsFy6hbcNd+9XwFQRRfaAuKyDMQg8O
RHmlHRpvwuU1SvveaciXaTwEw0zLtTyT55VCjvMiJzrnybBij6+rXKnNZ0iwnqcS
CmP1FupZ7KZA9f74lrLZMaWvvxoNriFTh1z9uOOhW13tOM//awNdxtPz2d9ZMpoW
F2MdJNC86PEIXsZ1JWXNOh/dOsh9wIZ9H5cdbAboTf9R1KBs5oKcMX8ncE+xmQm/
F/TDgLvUXzNE6jcBcZX1mvK/xODWzG/kYQtm+WXzS8S9e6V96tVQU9rlsyr13mXD
31nW69PVy4BHGKKKEsRno5JJracfL0aFvHW/ZYZhZ/zvbxOsGufwo6Ga6mhdn8x/
po8tf4dkjp9qKmFxmO/gtnKgC34cJnl0nIo/36Z4mCE7QLKARUnOEZMPk8weeYqD
9KG+nlMfgIFA8yqRZEsQO7txkzNP1ysSvDJvb/7EZzOSJ8K78lTrlEBFkfp1NfEu
GsovxfbvvE3WzJH3iSLHX92XPWjSCkrjLUMrbs3oYZxjPP/hU6foq4VFxv2eclHn
/P2HKYADV+Gz+KAwJRde4OajWUaFbpFVvIth+9UyHA1I7d4R92LRFFVEd0r0GlWt
T9qgQkSuwJM3ik21prZ705Mwfe3XdBhSu1bamLIDE4FFJoV55GKDDK8s+S8uvum7
hdWOjBArQiOD7aD5b/9Z5Ckt7ZQSzkxhtSP7ur6Q4Y4/+rJNCpSAlfngkwOy+vCD
0vSVxlxOYyaw/sEOi44uF3TMEPg5oSF9LrxV7efgDcs3Ou6BhXevR4a0RH6mn2u7
oTjK8JWPVa47A53R26C+HmYYiutyioxVvlw5TNYsiNAkp/5MxpExs+lR09agcoYA
pUJIhIxbUwxIymWcdlU5lTxpNmygTPZn7qTcWaddKiITzJpPPUdP982UhQhBIKdM
jXN97Kl3uZdprwleI9nkbmamAUp/gByhKnj4mbxeLmGCr0T3xxXTtx1sxcDqO+14
7UohP7HA4STn5D6QKlyOHAO9T+0hZk12o1lIkgZTJOQP8iWlCdSbv7tjawL6cHRU
8HFnU5dV8GrFW+FqUartrq24D55hlIfSUGLegT/t7L/1rzfdlfHHWqdti7EFDJBG
5FUZsGCWBDqpdIAWAS8Z96SN+6E7x7JvFpITLOAKiNZHPuNBmVkaNXs1z/GyqX1J
AbCXwWV3/ugrsL38Kb34r/QPEXWEaF/UEhxvmkf5dPXGTEfBeM4v2MifEz0sWV3H
bvTbe3c8nR4Kyn49REqkX54Xz8qfscyBh1pmNmuEjA+Ju43V+60UHP3GHo3Y0SPT
RIRJiIBBZpAue94NzADCDjxH0Nat+KZuT8uUwkUN0AcoiY+kcmOfp66yxb/NetBM
d3JiBZNFTXjEwQ/eIEabFgkzKmaNByoH++wcMCGkctxGfuLLESJv7Fmj/uOlz+If
H5r9BuKFAnlyOUkc6miAh1F0JEYOAyCrqbcWd9/YMTqUb9BkmO8sLtVZ9sYmT+eP
OSP0yCggg1K+X27aPv4yGXHGRNLV4/hJPM1i7dSQ58KMWvVhdFnmT+RsGaR9yj2L
UGRg288BaTos+R8NWxdSWpA3tF4mCNRFWb5HQx0nyrdeHLzyeotalsEA9Z5IPixF
RWO3hww66cYuv37ggUvjQ0adHgLUEO81HGGqUJ/Ct8Uqf6QuJCKpePLdg6QXLDFv
3vmR48L3z32Wr1sOVU977oaamUrYX/IOOMacDIAgzPkT9sKLeX5oDksfrNa433TB
oOwfNk1DDQ9KKT+GqI5jcCPr1KyZaBUvojHTR7CKfPoD8rWKrH12ATipdfocQ0Xf
2ukDvgXLADc6UiHBpDVYc3PJkstltAUcO0eWsNAICoEp555dnB1PTxSXpEEt1qMU
e0Ltx5pjdHuQVKv2PAiej8ET5jMkfZOQSsb5A7Sg2E6ZxZDFTdW+0YayYQs8aNpr
A4bU++2K9ZZDfQVkaZBbKjmLtCw3LQK/O3ihztO1W3oY37wP5/kCGTpbjJFT1skD
MvCzq6cTvT6otbC5fLaG4M7wi0T+jPRVCKG1aTiuFcShjT7/OFgQ0p++ekggjmuB
ThfcTuJfidPKTAJ6QbGckHLaH+GFJtEdir997VI0hp+H8v+rpQ/1gZ20orI+ks4Y
vrJkOnbj88Y2AEb80DJRWl1PQmY31f+oqfrrE7R/e6lgdn7dskXeNETQhezN7FfG
BuhmpG8vDKuS+cYNMlnwaweDkfBbljxRl7Ef0/7JZPUj3LNUZgdHqucuqKjsxnC6
jYPwsh6gAA/tp5yY9SkTJuiK3Sn+tzcUMwfgF++yvNuxZKy2VKyhGLaN3RztLjFG
EQLM4NVC5hXPnec9nW2ML7uWU6UNbbigtvZ1cM3uizTLQ3yi8SQ9cVS4BZ3EE00c
4OuumI2XTbs9NPgW6d4OX7HjHvKGX1vKtW3XYa5S5E4sB2ejQQWcpfhPqClMCDiQ
8AG6aZazyca1p2y6JyPyB6ARLvRR3TloQQYJYUsgdlJI8z2jJp9zsjPifVDac3Vi
JemNYuob9UKAsbuWTS3io46WChNaNYfkyVutlmjz2+K/l7Hn4pcXXJ6nJh7cJdnR
/8+6qK0/PXvpW9r8e52B9Wh1rAVtQwGczEX/d8F5HJYsUdPC1h+DytBt3sCbOkyv
wbYHcUvfcmbuqYoq/ACU5kNwaupWmh0PaCWgeEcb6SHW5VE0VegGwcGA+U3iCDtd
oAQJam+826WmXjGoYUOoz6Ruz2K+1QmXZFdUzFQOqhUKpN1wJDc71db4+KDzmtfT
dl7nq1ZkUL70o3GTd2V1swpElWoHrVUyAvgnwya0qlPXF1e5R7q6Im/Ul54zsBKu
KRL3c6AXzCxvyQ8tuEvnEaQiuM7szktGuo29FGwqma8DvgyaK9XtFv6OjCbMh519
HZTUiTrxuJZa20WrHFkoWFtxDnjV132ML/gBKYWLZ7SFer1193XeZGY1YpHmCyWU
jlDQdMqTk70G4ZURaSNhkSWN58voxbplt/Uu67IrcYkOgWBWNd+rCjeFx5fH6OXj
5sYUfme7NdUBdyLriivfRtulUQIIKMcuudu1yELpz+2W74ZnOv3XpE5DX9kaQpyo
Sh6AMrcApXODxbUZ+/ujupMwyFXX11ku6BQwW81il6DgQjaatRC/0v6UywbbuJnS
0dSMl/Jipdl5cVXlGf3GVa6ltHf4oFYIiJWlCgIef0BnYzCrkWKO0mIop8rPn33i
kJ5wjzlg3G6pKZCmFewtkK6+g4hJ7bSkXsYQAEqGpZ0rLKkDJjTmpJdgFdVgVjQl
L1J0EpVlx8ftloKGmBSBxgU6rzJkp6wbrBonHNpeK7VIcrjht+knvmwDpsOdAO9e
PLc+BXth4d+JHCPnYqrMCGpaV50mpwuZyNgH8qsumiLTq/5VDIG9xfFms89rlB18
JeotqGPseZkuc2icFxMjk17QYQj8h/HOTB0MQnzGTzR1xukVTKOTySY3ZaXnAcw5
cNoezQsRFOIeDQ0wUaGJ8iQkajd7usu8EV775FuBd1LulvgcE7DvTPlAqs4DwzzL
OouY+VD2HPGB1paAy9nzxUtmFgDRvvfSkAwpioPhSLRSMEL/hNheZ0yYBExeLyBV
O2W+LPr15AhdEXRMvxEF6lkcb2Qxnw8m5WSTA+NBJS8MwWr+IRkJInQoleCd42SU
QkFa4hxTNGAy2gwBf2hAc5UE8vLY+6yGVSeKH3myoejN3+dNCtAB6KNVQVXC3vNX
7PmLnLTBevgdDOF3Uo/nY+JoQmHKLM3trwvpV5zzieJZvXWEg0TrcYersOD2yrzf
G5V/K2q0l/USKAB61RcNvyq9gi2fppzXFogMhO5ZLdTDxxatHAO8e77EJJS/oiTe
zOOI/hq3HVmJbnz/Nv6u11hnqgafwhRRyrqICpCyZsVAxL1FzzO5G/P+5UAqia+4
Oe7Zh6DjLr79HMrGsom4FU1kVXT7P54vCIkIXgB6S1cCKYz59wl2w1ydxZ8TRrCj
4NM1ZE1u0IFDvt0JCTfuQJrATssouCqLpwrAbUTv88jL6ThqXsd0rDW63DiX2Ajj
TlabvvkhOLpVLFLP7yHnOq6ZDqbFoQXkYB/JLGMxlgqeBpatfV4J50w1d5P+kTBy
1dyLqRjHTtHt3B9Mi4alb138STzKpYQZOF9zfEczdV70uDe3jPqk3dMiwpOHDFz2
RUtG+BxFu3qZMfVdPEr2LI9DKDFHvpqIyyE41G1eMI5iQQZZIOC0pCYWpyz8IAlW
QHabj6+Q2ZMhv8/63V0KmgBRMluJlmEy8E2qksF2sK0J/w7QnEu01xIETJ9F1Fke
6bT8yV2ylA2zKYuPdE7kHpz+hGg7N2rGa9eAh/rDbkZWlrKibxt/wZo8ao4oRX//
G6LK9I5tvfLfi0CT5Lpma6BY+PRL0eqkw6DWD6ne/8VQX3AdvDhESfJn2SIUk49A
4oF4QqK06lGqYeDd5U4/zxD1b0I7cy5OXpcG+7glBdcdtZNiEggdGnT9/Gc3AeJW
1euRsI2h1YmIKwl/JsqcnEPSd5n2xMWvYfQGeP+Uv/+ag0mX/d2GLyI6ECD+ryOs
DZePEyG4CGwO38Ar59o1JVquZxXSf3OWkfhvLTSnNqnLFR2wXV30cMXpFpfHqftB
nxqTn3xxjXTAxPAdiaiOCtJk371HUr44m4LsRAEfyvakTGRspfI7IjILbcSGQG+E
i4UsFUl+y6L1dHkVd/yHG/jiK7TAPM4Zm9f3E/hmpHqnVi5u4ATL26qBwbvPAfop
hsvI6/OcE/+dL3zuzHKj1Iy9oaB7DELGm1Ze2Q9yuMvyJyigTUZnN+BdQI0IYYHZ
T7tCEWa+BgpAUWSbl+j5bZHLULE9aZOZC3uNTWa8zwKfi/Y2xTBcPyneSBZB1gyq
G7/33pj5di7JHL985eGZEy39virqjoDgywFZjIA0wkXsZVtbeB4xzA7ljeVhtyLr
tADbUFYtr3p6F/8rqm5D5JyAsxS2JLzD1CKnmBf33RSf8hUkED5KexF886+tkG1n
zQGTlxUL6NRDKu6byG0D5lhGahv3p7A1MIkEHXIjNM6dDxLjEi9nSa8ma5EOwNHr
DWMr9IlshtPq5+TFJ++7g/6wFyReqzIjGGiun2Ww4AxLBwzqa1cXHw2t77rVSrNr
GOGeFiSiA9bGJ5cxMTtdh+cXMzH5tjeQX3sqmsHpFeC1S9TqTvrrv01vIpJAzzmf
lG8xLsxb4PdNDtvo2w2sK50Z6kZnMJpk6DDchhu1pLGBjMDTQGobgyJ8Bhwlez0b
SOJugQPWcBnpPeECBtCGcWN8OMabd/P5s2YaWR09Yyw0j139ObF2B+yeFw2Qiwn4
KewMnBWMk/80WhNRSG15Cx0ScOZ7fYhu4bXVzXPZAeq61EnUmv9x3V5dDIFrmNxJ
w+7TkUw9viloSK15SncPAclGDof9VB6NZHeM7Zo9OFgLzKvITM0eW/OcO9i7xKaF
tMx80Wl9GLMS79OKIb/tEUpWDecs3v5tPVJNx/yH8nmn/j2tK64A/J5QInfIDSjE
4TbV67QVNH5wwHbTf9teyvMEyK+zqtSoQQV/g+hoaRH1u9PX98ofDl55g8BPhdYC
SI6cGBJCBEEL7l9Mbna4IxRmrj525N2VLVd3Hi7xcOWEnuw0zL9k6souV5+mFa2J
bWpXehP6v4MoCFJslnn9WrTs5AFpLBGlyl3tm7wtp+RlW/UQrHgcKmQ9Kqqlp1uo
L1A5aBczkMoA6nmRZO5kh288pPQ+KKE6pft/MVtVMVvHXOU7Z9/fARhmMABokXjg
1X4LGfhOOApEeL1BxE315Oy2DX029Su12cgXzoMeQMKSoUr8t625FxLUYBFM5aS3
vKlJaOrmlGuVAm4qeYBTNY/4EwE8EQlunw4gq2mdOGxV7Z1z//QVrSqA37eYjYOr
HcvOu47XILr0mD1A/W9oc6FUjBP7cEZiDsVDsFYlwKJBp1voz8fQSJ/ENdopuo3s
bY+KXweOqE6ODOv/btvz9WzV2VKUeIMuby1gnQDmyJgAxQF4Xb+bUil5yMSv9GLm
7hmqvFqVtEYp6DDhtg5bf1LrERxNRhesfJQ8QVo/YAICPMYGh+nzOhqPDsJEQSFH
YUlOukP4dliSr6JXxIbUthThcuNIgDSRBHphChlEeUtSM4aC1L1dqqkLxGUYvd1Y
zq+SlqMNrpPgXXsRnQ2BIlKarrVTV24c+z9q62EdnAzzyS/Kc4BVt55uDw63KMOI
PhXMmSeV/zdgq1HqrkaCnhK3jFPnBnyD3LwBQBVrSijsBhp5I9/JKsNfCMymLc9h
53528M3DU/8HiynsFIOrIbOVLlUmVbMosLb/32bVD/q4Gvn0WCSYbZDx3t/HdaU3
67Ox3oYWEI2onpp6WxlUNCgkGN2YzY3Vsbr8sjxo5lzfUkUtfaAfT9raesJjPKHJ
doR6RfB/5jHYEYgA9Tv485EU3owqiIrPFPFJ7HSCkwU+0BlhZmLtBN7ZHcmEjhJQ
j/sF+hpzl0+q0weBqddk+QGptk6p0ScJTo06SCdN8sB0APAhabmXh67TW+KVaYEW
wextlmZ8azSldp6r4MEFeF6NTbvoAWHnW7KDNJuBkB7t2hHjca+zDHaNcLVnP+qt
94auR7tALPqd1TzPb4EJHRzXdT6UH31hWcYy4Qwq5x32etMtDf1LOOzJAXIu/5ZK
pQuhVGNk/YQnYusSiVlBJvq6tttwY2LTZCO/GwvnhV88lXwcN6ElHhWmLiqf+bfG
+4pMoS9dISr/NZVKV3k1x2OHsAjYnTKdTMGx0E9uu60XdIv1oE5QcJMnCO9SWl63
B3oWJTcNAI1GmRtGU0AFhmJ397h87zU3CWO+HY/FVolLMgluZBP5i4yQPZDO6Ltd
8QrrI9CR5laxGINK+qH8TTy+IthgX66Hpzh3N/PMiIb1k4qogEZSTRKV167PXHP+
eTAQf1UUytj0zklUc0LnkbsIuTx5B55I/F4TpkVsrcktfm3u+fpIL2sz7OTun8jY
WJLfLX+UmUiU3aE077HgWYrdcrrkD8vm4U7mIgT/uJE+vyWHeqIYGSZmFq/xKLiU
JeSyDbN3zMppDdfoEyLR8WgSeoN9GeRFPiYGzth6mR66vg70OUJQnmFTNmA6a58S
6nzodph85Zj79gy7axrsv9Do0aOYOWEE1Dfjac8ahItpVqM/+Qnch76dV7n6XDKf
aef13od7wHrwOxp6vzfb20OX9atRHmmAYNcrwHfbaVZCuqNj7enzlwshGz5fPlRN
8zgcx9hNE+vQzeO2lpQ/PFAfBU8Rmj6KQ/XJdmNdk9WUQ9WE0S0gCo6GoxzeufWT
lUCXPBdKCDGYObfe7Am9OLQp3Ucgk8+qTet/bDzPwbAl1E0xTH0wKX2o+k1+ooqv
xa59zhrc9guwFwB4dPd/BixyjgPAnTCDMCIirl6Bow7rglgxubmPtlSEQ9PlQF2A
LbOhBA6zoU6Nmn4BDh0+FQUGAyFpbLgO8birzGgQj+s0XtcX6Gc4AObTyqGOY1pI
BuWG3UOaU58TbbttznBAym0W/y86qdtMPJrVWhQh2i0WG/VmOG87fRuSpLbIGFjF
ERFS8u0Ns8UI7h0znZVBkMV7gwxjaP06rSvOfqSyGVXdV2PovXqXLpfocdDKJeI5
zt1CKRo9Gtrw3vEZsvSYAIePzbZGnXlwXIPH8wYXzolpKPc19N5v7rs5z60CvNnl
jKRznMB4rWenoDBPXklh7USm2r3XPyQcgTPQxnSdSS+nEAHWLnB+Lk9PAgqCrddl
8lPFM7nU5VGT3NKbfF0dgHdkApj5LpMyP6uKlENiJDDjgLFln+iJrHqw9uHKI/0k
CQauqT7+9YNUsBQylysADIq21kMGeXFvYeXfsoYk3jZ0njHXZaDM6LShLs2Ydbl8
sOvnrQYYDLAuJPMJgjrEdeg+0NOfkYr9S4vJfYCE92s69a8JidX5Dca+vqv3eJQU
4g4c2GBRsFEjJlxINdSzyAtbdzhXARdvUtpmS7Pdw4YscWjrAITsuGtoGfbKxJrS
3/gN5gxnlCryyLsm/P/CTzwlMjKpttQcPs0bgmGstfzsIRNTpgnwKT7/hsGcxRxI
A6hFSM4uj81lgyH6U+GUSI6fx53KlHn4t3J+hituVixDF8uvI/Wr5FNmyQGqPDsn
Irw9/3v5shAF2LnrSW9KX/dOL9QNRj4+MxPwUkPr1wVe7BLPcFchE+edB6oiPyIP
L+g2E6fSU0/siR21BMDfwIgauopXzHlQS9UcXpr+o2LmrVGfxgniggirko6qpPn5
lxHT+Gixk/97ApjsZYiOCaATJTW0558yLNZO5W9sWv5gt4tdoHrv2Fda12g0Ywe9
8Yt/X76LE+ALLXjJvPpDi17gSO8IrJOdJU8CISbsiytrRgAySh5s4baPt3bB0twy
ny+uRMrgTZLG7CfNcWNyvw+7yEC2PwzzEtw8sZZYg74MqV1n+0Aa4zalc22XlTJ+
8iq8psKvI9F/iSIAGbb7xRkZW2gna2YWimS6dHPbkym+75aBQ9HYAJC40q7dW3nR
afxdaHe4vruA5EV94XyRQvWwdZz0upqj89mtyW6ZrE0AtHhUpQAKPhKmAvs4SXol
5ms4iJYAupWfuKwBOnm3kbERWO6KG2l8/vyXYX7BZmtmMDFcfuO/m9sRLtAthlja
BNdj1Ew6fAETXCtYLom34JDZwqrdJvUeAdzl3oqWK8TFvazO8SHdANt5D1SU0uVm
oaxxWox1iX0m1pqRpjF4GtS0qd2GTxfa+OuBaW0JDVEskJlrPhcvKvhl7TpCH/6U
mOuG36Nsbb0AgtE+q/3I6KEOx02wIE6gQAXM34nKYfuhuWgU8k8FfprhC40RhC6W
MrW1tpnZmR3tQgD2yK7U2cRAQOkAadS5rnjHZBzDl4irW3FLwJ2u2bw81D4gDUqF
9+UCxS1lQ7V3WrYOq/J/p4WXseJr9J2ytQkzC798+s78s96xBHlWPisGcbmA4fxj
pgA8f9Lb57BQu+mYy5triGbufeqAxq4VX3xbrRHvnODoEmZKYzgEr+T9F7vzOYv2
lMc971W8Kbf2RRiSDbCfceywl/WT8hmYlnDsJ7WPwrJiK/KcE1aJPMvx2tPwroPd
j5GoIyDewpoQwXm//+DWPXSwNhC/0I8f2RwKg28b0WOte6/chMpDKr8/332ouatu
45l7YFEAx37ywIwG49c/aRi1S8UoakWDiYP0nLutLiQRiSAmg6kX5TwYf6D+Gz1r
bIGcXrdBctXubt9oobQu3NTcldTOELe0VADSl1ILAiuCjDKAgj+2WIdzOEsiP+Fg
3rhodfG1fpVlO/spssAdD72XfDLXWVcPNIKa9SalanT9R0cpzVRDdFB1ASpPcQWo
tOo1I5joXc0MMy5b3y2bm2APEbFeFtwd0F/UXIWjY/D0PfVBjbeX7uTTTZv5Ecrr
BquuEdZ28ExflVIvk8asELXpsHIgvSkF0jC2SopBeZv1PupaZPzR2pDrHeteDOuS
WxgRp71GvvU8z2SrsnM3eWdPMFBbL2ttTtbzxgTs88B2gBuI+o7KXbnECmM4lhhK
I83ZXHRXft5rMKhU+4Rx824ASB4cVR7UM4ola5UXN1Sa+4oVWXEdERKu2hPMwuOS
trIRdv/clj/5SmjAGyRmcGkToGSnlAwTEvFJCI4LAL/0iPWrKDUyjEpuZlfqr8Im
HotIaRSBq9GVYXuIgoKRY80S9FcyUbNdsUhxnjg+KfETfkTSLd/KZ/gM2KFALESI
5wj0i29PamnBczN2iI/9BoZqvtJuY2xzOc6iAYjpzKhWIVkBlcCrff17VfmwFOih
0A/hR/Y7EPF6ZVIL9BRJJ1RYqZ23Jr6Lm5SQev2fTvFegZm0zsbaFitH+HapSnM9
rnZX7AkT8EPIRuB6ht+d5/TtdCEvL6KcouSkF/muNsb0QPB2RIYnXHnpce9jqnKC
45xeE8QoAHT4kkgofPjc2/tboydasp4ORo1HtlzCkBa7nvKT6gJyg3VRW/bmKsCY
7Mg3lXpIrj7/O0nbsDFWNiDofaVu9UwIpZ/nPcM5uau4dsq0iBAmQyliMnmlnLu9
DR04TVaFtDtKS6YdkylwIJf5xrmg0QyExUzByueyDM2Pu57Ff02T7KFesv+MClWC
WLCrGbNQs3ExxdzQeV+aPS/wlDeN6YWWCasi6ud7BF04JCyZ4NqamA5ccUdQ8dRA
ydJ7ujgj8h3naWsoLVbPGkGcGd0Thj/PniHdMAjatwjD6KFM3tyi5UNYrGHcWya4
0REzEDldaEBLSq/eCMLGF01GV1d52vEPaftfSUOgkttQCgj4bVhflNhxSovO9B0g
/Q/ZVZB5Gh/li07XPdqfQ3lfalE+qe5uFPHb75J945qNHQ6wcaXG2RD4ZhAZKtW1
+eg6MZ0lypgVup9PvZ3U3zaileQCoL1ZbDSF1NEKI8/5lGxHD+Bwb90vip2BzKCT
87HVcbI8mo4cR2hgIXoJtW496V/NteQIhhIznHZKhJ0q38QxUkH1bNmu6FZa940z
cytSVpTdOtQKZz0qukquSotknIfBmDUVJ0CqpejT+0NPRUzsRoVR1IRFBjUEcPi0
Ctr8PtB6y9rNPsq4crnoAbk4OADmTiEobjj6KRJvt9mFmHNNY1hVH90Mjxeo8ZdE
ZckKAOO6jfxoSDFeT/YrqO5P6ab506DMrbmsH7gqRcirekY4HRp7dKKD2+ogRemq
h0+Ri2Rz9iWt3udqfOwF2rA1ABRH+DAsdIROIWWEn2D4gtAHyuLSroodFTvtNTop
WrCCliP+X4spd3ABIvVLMXsEoGUF8UEhU9GHd8KfzSaZ/u5lrCIPLYHAjK2HGwBQ
fiXopm8bRRn+HFmSD20flCq5S9PEw8LwB8kRG8QfqFUq+iibaRvalJT6otJp/04z
D1vO3C9cZmJLsrnDTKsi9G5NAto96n4J5WNNIjjAJOzWUx4aFd1lWG3YXiwO4HYU
OMhbLED+hn/5BszqIyB8L4TZ9m27DwY1Jbn/l1YjLDiuie7fWNe5aFgPTkk6gOrH
mklE0wxFe/tfNGjpU0p0lTSW6CaaPGKzhcmeaUM9yX4dbN8mcRrKEakQsRgjl2U3
NVt1a6APxku4BYrDVw1yU3odCjvkmBgYmmHv2xlTskvMpiCiBoyTzauCu1CIrOQO
XwuGyTmBsXJjMws/KSGf3rzBnd8ezVPjbmQub4sihXgLOEXFptpJQj1mUiHao2tu
1+ZsGccjZYxlkhljKxd55j9pCeFIM9YrFnwspo5m0zPfK/ufH4ifOcDFh4SY+eAT
K+ct7pjgxLl42oPuR2+DK0Tnxi0I//KJK1YrMYFPfLdQ3HSh9DEiIR7KzTZrfxk0
ik8ORx/hXQoGAP0yIWtnPHkGoFlJY+pLExyO+yr4EY2QcL8QxVW8bV13NrVM1eCJ
PV5dDTWCaAvSxUUfJ27gzoBQuDeegA9av2jfXOAxNBqiV6CVSFGNV125GMOHucWm
c8odOQOpV/P+dbNGp7uMvV3uKk83DKiqvidVBuEO3LY1n5TFKBs9twaj8M00x8nN
ArAapuhzFCRPxAm6wSa9f2RiewJezO1oiJIvYBZTf2MCZQuPPbOddjx42/v6pz0P
csJqYc9U7XdJ5DQU9DGv47cl5Sw9Bg/f2uqB9N6Eb0hfOM1W4ML5EL+7qPcbdwxQ
npC/9Capww248r7PsFtK2vL5W8gVu+Mke1zXMYmN+MI/ldj7KJ4gP86oGgqIf4Oj
fwzJIDk8aIkbBkADMk6epl5IfwymfAC+b/B8kRGdxdDOnai8sF2NpDk6LFzl4sQA
5n/OS0DbfTI2t3A8Fl/57uHFQr4jXVLvKN0PsWzsRGuIZRVvNX329+Tihpnv3Yie
8h+fq4SOEAgyPhKYsTSQLaIIay2EfNBcnH/wNxCBEnfYqx7fTKeJSb+j0Jh88XKl
0nL6qJhTVy/pWN5CWrHnD7Li+9X8/51rO2N7aRWadnhsCX48+/Mie4Sksxc31Ovh
maf1c6NrfkLQ9zL0I2jqTsDEFoMvcUDwx9vFsXThIPPJB64+czZIBOZChK/Q4LnJ
gONPzzwtn6UxSj/Ic7SWI4KptkFUKhpbzj0YQ/xtQrB4r+mEDACyW7SPHDSRs5v+
cBMsZcW6x38JytKfrdvaQhu/eN6hkb+adSTG64yjBB1DuIHZoaA3rYdnKpoGlpOp
YdgaFjMzxF9waqe1MIlhei5zvQeXsBw9hh4e0K7SCXA1NS1KgEjDagjkOYbfQkJg
hql9sOKywzLXnVO8c9HE4DNdVRgN1YF0Srwqk3IeVVHyGOqkXThQxfay1FLftWDo
RO5rfDp++4yll9t0mmuzNFC5x/lOjcjbHwuXs2Byq/9Kvho+I143xYazuJgp8qUK
7BXwJx+IIwLJBFIpe19Lx+2MLFDvFLiYkM8npN4IJp+1qBm0rFjO4uIERRZNRtzp
b+j+/Hdpmahnf+br0uLyqWhULcrMH0oFwWlrO1Xxawjh1ybcHng8KhW/psfF8x3Z
xC4rlkRJOFXWK16zeF5DGEz3KTM0B/ZRgj1qTyfUdPjtr5w81mb6wvZueSTfdpmc
1HzaJHchyVFO4O4tVUbXNkkY9tDHnewBF3KavgQlZ6kyBOjypmDdNFXjEV0Y481U
VrY2BNNj5m8+ieA/sAd61gRIKf5nM/HxenEl9eXwYCYZ7SMrZNP37cj8G6VlxErA
fAMm32nnVNFCmQLjb4lpcb2W6FGLNBvrhejoqkF42qjc57OY+egYElCnvWXpRY78
/hht/ufnH3j54No77S5qySOhi5K5NtO+DSloc3n2fJKwjbP8+ovnfXrF2nw/koB3
s4IeNnWJ/ueQ+4P+EbJY5BgeFs+dj3NQpQqxCPHYK4mmH6KbQQKnI4yba7sSW0t6
XTR9fhZSWz5perS5Qo0sHBVKxtEwB8gpbStuISU9GFVfmXi0KqvNy9P6QmoCX7Pu
CTvEMNbQFACjrWzs6I4QupLD1JVS/FkVbxwOhatsq7ScCS6OFbb8+cxXApLDEt67
3WtY0t47FlQd0wtbS9h7JkGwZFTxgTFsEMjkFga5wRm3FLQFTAM8SD4Ja2MAwQHv
VXfR1SU3xnryTxe5Q43a7rooYL8gLOqld3m4rnI22KB1FkaE1ijpym97fePGVoWz
rNYMakS51xdytvizSUl6u+6il+JMydltz2YxuWuwdYyQc8B5A2gs5ClMI2+7B/y2
c2RNSXR+ll6C68fB+heysfwbbcgUc4unXmAWYcYru5Gy1FFUS4iUDCWTcqDFcoSx
RLE+9Vdj1x6zXeQ8txQip1psrfZ1NZCm52f2KkXkt4EmCMUFiEEWm8BLEsVCJuRw
0U2rQJU22YQyNv0BSmV+2HMvHrWRaiW9eLbm5T93yURtA5J6sc+82U+MT2/3uCYM
afqZcw/giin84AZ9qe/RSFuR3znup2I+47kpNY51jFKhERGTGDQA+Vy7qI/4RFCA
ehSLJucDEG6ep7+YZEH9o3uHrsETHaVEeZ57+kj5RC4FHUDBveUXdgmSzpn9CvtX
IIJTeNVnHzKdgTwhOLLyuF5mooDo8zt7/sqSDKxdPXGK8SXarhPh58yPiX+Pttod
g/YAx8h3SNLxlaJMrsus/ozczr5SdUHJbjP24KT3FjVfid0Y5R/gCG5TR/LmtwKO
eq2iftK5q6w/H4+pMihjSD0ryXgbBO+kW3RPuFjXojwPMM4JysR5oxauWOR5OpjG
4LXw1/NET0LUqWXDh+oPdAqA7nk4J7ogZrvOGLJ3dbR1D7DiOSe11JhURsoPdd31
Z5cbbTVxGHHoiq/C3Ki2QkXeAOTo8/651AU0rzF/gCg0C54mpbE5e72Ilz8ZbYZw
jalwvpffstp5+scUTHK1Wc4m9zKm1mDhhOXJ18MKgURRh+RdIj2Naml2KSS3mW8W
SEcpxL4kR9LszqfRqx32nPTAp/bQoZhllO5N6hK8Rz7pU5tbPVtUbxIKSGWgbZkL
hx+Cat31bRGsrzzSBOrYljatTId843DNBCBWYK8bDvKqCmu0xsg/BFWp6WqyU1df
JZUzaqFCExS9CwM3cZr8wTdV5EwriFaI5qHT0fNcxNy6J+X9SHIXWzhyXakkE2D6
GVdR0MyaI7zi9JEoOlHWBceoVXbM3LXdvHJvI71XjJJbB7au1401emb4TyWFsHcV
16eB37rscreWEhs7KVs7cs1SFxnC5tpn2VD9zmId8e9dlpPay/0tlnZXAN45diPH
rN2RnezpWbVJR6xvNDsiREvIaygjOF1/u+rCeJnnDudOME0hcX1X21pbI5dhMBwL
djUH0eJMVuKB3K5PA9+IpKlKCDN04u/ThkZlcL9fuov0j94ACotM/fy79gPVrEoz
WbB/7VL+wtbPn+hSr7J7GvQrLjVCntSPkW/2/4x6TBo0Hw+78/OlbWvN1kyDCfim
fMCpwKaG82io2fx4XiHuvrfg+vvX//Yhk0qPpQ4Olp03BPKS4BBXrqa11WzuAwA1
zuURYVZEtJtSM4T8IFxdnq/fC09E10Gx0bx4MotK3XSkPDqB3DBBMZ1r4SBn2G+k
oUxxSmXB0hFDxfUsN3gYsHsDICpCqcRXnNh8VE1LLe773uFc0YrPeRK0pCEA+aCv
Kon5zGl6QCp5vWz2BDzZKrCM+ZqxuvzfIyqOM12VrCyOftt9qU7t/Ph55Q70q1Xt
79JLsYEuX+FENrNMd+m8jjSFwMwpDkA72YvkNISxvDwmd5Idsv+J2kP06cfAhxjQ
c1SX22h6FCNzm3W3WZ9sC2gcbGZkxlFZh/saoaX/QVHFEOWcJEyDGesb4yqSDN/z
wI8K3xaXnPcp31w8YY4crZZy9gC0ETwXVts/Jh7zRBR5HzJk2nJPKl1xwXA7rgox
R+VMMgaYUYinWW1P/M7ZpGUmrrOiWb28n7c0p3WiXf7Pz7xK3tsxy0/GFh4X0eLK
JXihfEO2fj38cZ2qtq75gZgcsMC2ikz3L7p9balbNeIzvVXyu81UDNTuvABhHOdn
7mieuRdOgIqbHLzmpQRdb0ez5Gln4y9ztbUJtGUkJC9foXjxJrn5/ex5zZAUQbuZ
KlQT01/1STKeIxloKRCm4kECauWBOji6HzzqA8zmII1b/ccOCh8hfBDS0MZAYG+k
iM7BxK+JiFj0du6Gf8Ohu+Z7fSrVQw2OfYnmm6BbaXZ9cTwZY4i0N3qwLuOIBPkl
JFfEwF03lmHgXsr8Jte2c9fiN7U0AMtARYb+2M5pfQ2XvTRknOkFN2H6eXYrKHHE
ovZUx2pOnLbVvx218Hj1IKaiWxtmE/QdO2SDNj5LbPeYcK0msJDW7Y+Z3BMGNiqp
b0EjmwQhSryJmzituO5/inNNYxbJf+zd1p6JmCfxuTy30UI/PNg29+C3k8M3AGhH
MnA0z6Sg5mnJ56gkmk7t7SjGxZM0kGd91RShyIWKE0sGp1TRCNM+hZB4ceT3vuMB
ohkmz8D3no4D1EdIyo6xD1B0RW6ATS5hcRWFqg4DPLvMx/p+i8xuyjcO5ZFt697E
SSj6uLdst6QIqjYeMrhfqa16Qz0CSaHNfbwJy9nJUtEyyN0Ds5kkYqEUkf00G3dM
wtNGK4M9ofObZI3soOGCVeSKgPTf8PkzYBjPxNH+8CPVE0dIQumth89yuyx0QGLI
uqp94rjqcuQr7s2tkYPJSVYp49IriCQnJjGJh+K/rrSBLSpkUmnB8FNZIvTjJDGz
GZQ11Ns7TqCUov4V2dbCeY5ncVVkskeD5D+ogSUadTTY4TJnJsTbCuJr6/mJwlni
0lzJp3fnU27euyqZcZ2vS7yz7BiJ5oEQrdFIpDzz9QLk9xDBndxhSj7249Oj7+/t
hKyUBocfpnWIgNdhJYsiAeSUVDk3wlfiaSBzihFVV7oL6Xc5370kcnXhUDW/mUAH
ykPvPsEvpTRULyoEpqMKM4ckgb51a40TD0rdBTXmzyoY0HAy9UYxhl2j19nKfVgB
IxwRcn7xy2RnIS7yxkk87tK7SuHTZhdPBnFO/rtZlGpNV0UduDRxwVQIS7BNr1jZ
oAotseo+lCqO8Ienk0UUm2mmXpxZ7rwOXu3otd/P+qNk+pZalGX0wDrElkgWBSQ9
ksrVBEnsGKxyejn8U9frvT4fQuLl+vVNkIk5VDzRfNC4D2etWipmckQ2yxq3tF9y
SyKg6m0i6YLiekSvMrl+oBOrPfD/pd90LyWY5fr8NSHZjp07vOh1TTVffoljmGU1
OcHkrZ5LEzMLgCuT4i1TObTOQfWRV0pHVtC6oJo+DXHMBwDbWumdl4LsOcHfBTsW
z/N5wJwDVVRC6Y9LOlaI97xy212QzotC8lYbrxCHdRyV9cCE1QtNIjieFK4f1gWg
YU9pFznSrKrVCcTzG8USZV75REv0T8hL53sRG/R99USHgTMokeUE0aS6Y73KMa09
Vp+Crzi0IRheeGVRoLQfpDdLUWKEtmZPETs4zsb0QHKTDWipiuqghC6WwyCTlcs1
Vgc6ZbXDJXt2VlxqmPvdlF14HQ7yhTLolaO//MdQvbJz+k+aFb5GhcbjeZqNOGa5
kGKgVwE+I4nmjSHGBct1cr32Qyqu1bVdzI4NRI4VN5HgwZrz4/flcbCb0HyZfQCH
661s3o6vN9QqvfGl/9ChCdvlOTvHZfoT3rNBXhEBEcOwVWvXoJTtnUASyeYuzz80
heenkmogDDjJhMKkCeFj2zlXWDmYB62Gbu1+1OGbiVMhfn/I7CXhqmNda8Q6GO8F
YjecHVvW4vp8zp2CCkSJTkmoD756+1Wx9dL6RS7e6z0zQVAVhMLh8rUvnkpsnwYh
6TAS3Ky6VR7D6pSxkENXUe/xsgHti6E46Rc74MK4LBA/rkqsKhOUNMxUXytuPkkT
vFO83uUOkWNAjTcPW3jcfqsqdPNqpV5cHYgm9kfWMgJR9XM35s7UeJbrXwfmdBOc
5KafScPT9RtJT9oi6RoeYjiFTnKPOSqM67c/11PwWK+er6RTgaOUxQbatdV9Xn69
riX+yqg1s2se4G2w5El2lN7udr/2Fcx44M//0oM6qCTeJaJCdn2L2o9VlyGYxp7J
fUqVgbWQgRy4Yx+KpRsXe1dg6hOAgA2QEM/T6HnCIHKdoJNKRMI+zM4tFgjRqHxf
jh/MpNQWFc+GrgZma2hcAmyJSTf6USwHyuvH0b/5caLPi6Ma05FQEAoWA92FCPL3
9KpQYk3aHq2+S1dfwdSZoPi/ZzxwAmePBkSCcSdtdd7Q1ULEzNkoRM+wXQeLUkGz
s1JjbByZyfCw85BRQ51crFE0NK1nRyFxOVPwCp75UvjM57ZBhx0w3v5Nbd0KI6H3
NQ2SgAdhpJvtcTwzEZd1xa3F/xbRorXYsY5K8Kuw0AXbbSeGb4oZoco2H8XpgxrE
GwF+zYuwhBddLdAJ3hWxdyirkBiQPmLgmPUz1EBbaHzr7k9vVTw5FAKUaENb7DPc
5f5TMbTFCp1S9FELAO2h5PndkpTmQjrxWnPj7cIUZ/tATiH8H1HmK8nwhHEyysJL
UZcGPPYkGpGy2XxFTr+5ysXnXdwb5igxMm615OzlkjO+NfxLN7nS7N8YzTc88npI
3CD7A0iT77vKTvLrscG1rtl+wPD6VBOQBuBP4RL7hLejEC1hnIDU+xbnuXWr7j5g
CdG6zq/YxpvS6S9f1bKg2AtmQd1diXDiYBLela5GYnDu35X4woMSnteARU60y/bU
G+/Ezl3o/3gu7ZzMceQ3CWC0r8jLPL9kicb/1OX4460keeFACp9L9j95hPHfCH1/
pL5MaMZt2yb9OgXfL6INuNEcY8puwx0LycHrPwcQYl4SIzDFe6xD8vu6+li8JNAF
t0QRqGCj1ejsS9QyRkWzXh9jdVw3F1A+pWlZt4wdlB1sNpfCterCkdMC1tUxs/vo
ANQC7Cz3Nl2JFIZ8tFgmMxWqdHH8Y2Tnu8PJNNaIkL6CjyOCk6PHvkAweFIDAXGG
LmGlbd96E4bIKsnxav+cCWSZWRD0NBgE8YsSgmyRnjRjaUory6bj8JcZcaQjVMgO
AN6phy3Nm4BLm/eOfp1Q+e5B0gPsUlJxdoMz3jZi2aaSu6b51Nddlwimuc8yTGdT
t9Z3//4nd/HngDLePJDdA3JI4WMJ4A5Wzn+2CxYfL6LcA1CCklEDRy4tHxsY5yOo
riIOqqPXa4W7PnJkLSMvIjIPlksKsD+bH3neVKHJahhwbo7gbsfIO/Hz8Vx+Ku2Y
7xQqqKHHfn75iicCvuH82IokhZzgbNiRESPup9ZGSBWS4UyP0HIM5RObJ3pb6/cA
spRUkp9in+ON6DIdbMydPrC81h7UiqS/YWLPbnyIocmJmUaky1teiP0aaDrpRyXN
rebhua4VMii/Po9atR4i14Mn44u+nF5wBKtYSWH3oMry9uIYfYW5lQOp4Cm64IVK
eruMR4wkWZQaNWRg8CJe7er6zjDvelOHi6nZ/dvwlMZXSEKJzboAG8Doq3FMZOev
wcfSEBV1n7mlWxts4au5VQuVCt3MsxvnwmQFiKA/PuVrG61VoA3aENmnVzG+x7ie
KJM57VjUjyKk03RLTfrnFAIPDDrLhIFofIoyL5gcK0gqxhSDsl5PtpKs0WkVid6R
M6+UM1E+IT2gbzwRTflqn3pyL2QkyMRzeg0XieHL/1j9fjk9a38VAO63cAKJFUf/
pd3Yam+ZITSmt3kMAHXLTFufuffUYkb05VrVoCerpYn0gzHkip4ZDxKScTyqlFcm
a5G9r12yvoRN2XdWPf61CCGUEi3sEcaeM5+rgqU0IeKVfXCQa2wR+A1FOZeW7o+b
38mGhzbere2T3GlvHXRCt8u9UI+6jf+F3GZ50Iq3gu4yEC17ehHPW5tK5jEYtqJR
psQiIfjTJWIsRhHxWh5CXjBeXAmlO0bAlr06is5yIgmMdwr8VHYjJ30ZfAhswtwz
DCHm/qOPVEyT6vv4U7Q5RF4+2FEKBr5ervM4oLCWLNEMnw8J6woDYM0IL/sM4YIv
nBelpxWIbJW78K94V9p1m/uszy6CykL0buIn7Hg1gF7qkMcDYzccdNerzm2q2FYD
RGoBAw7K2oGWD/fqgTjJoxvylL7ZLg4dFEyrw0jpo99xHUaXuawXhQIo5v/Tpe3r
SFuDyw3A5gIXo2TNxl9YYRkU7vWgv58DG67F79+FG1jF6uFdBsB8npnZcO0sYTLZ
X9q8y7Iskz9fcZg9q/YBYFD6Xmb7GeBqLG6YL1heqwemZdy7ewUBqFjWL4cqLq2A
TmhQ9fB1OW38sjVidIxSg2LfHZLAxZIDuWvWv3yHv9A3nMB924R6uINL7cr574e9
e+JjAy8eRUnhLW8gTQjgadJhb0cr+CjR1oyXoAsRaOh93XU5up3Co/ZO5WhQnvGo
rnw4AzX/FrD0BAeANReD1lGoTP5YCgqUbz57jkAhUKhE3DXQ97ZPN+oS/tRfgmUu
6EcHaWcIjEb3ptjqNCft6mIObSiEu0ndnxwvgFGN0rxlKt5hLW9q4pCfYEdqcdjb
pwe1k7A1V9FJMsd/j1YkiGw84hkru40b3ioLoJf+3L998UiyfZpM46VzalbNSgHJ
XUD4jW1XoDHMFaEtYCAI+ZRGnXwb1pgOdDW23TPzDd5XlvvUUknEaO7Eul6FLyqY
KH6oKBYlnyJwEHwit9WP+o631e6M7sFkDxn8qi4MGD3oXbv58czIaP4GThb71O/H
5BRx4z2IbHX0RqJTaUQIQbjkaxGg4IMzyRviy/JhNDb/5xd/o5YFCHh1yCR0QpUP
d7ZnfqbKMXrkHIKaDqciJ5As/xxooen4qLNXVCxx8yetQ+LCi/LWvhqm2eVZi5fT
0/Y9Bh1CBYG9HgtXesTxqhI9PjPs8N3upxswJw77NChBHCWqIsfRn+dCT7YhzVNM
k6mH/jfmWAUghzIA/rjrthtu0uKaCiFDYnEfYqoOdZFowjOylflCsU1QqSjX0ekP
Ne8Q3h+G80bos49WzxCu6q1TrMpgF5+MdCrbb03o2Pql5w4J5Vh0PXZ+Gx4+3v9C
rqm6YwKy4Arh2H8taGIZ7zWeVuYKO1dVbs3MELEsn2UfeZkxstKzWQkKy/tlIz8t
b7WVYkXP4qSTOkheQnWqFc99rsNdjL7s8KRcCBdG0c6jqk9DOtyLW1jAbYF1nT/U
5Gz9n3GxNcP+xfyVa2oWNbJ1CTqTY0PZom27WUaNL5PbuoNNTW7HDGb4wvD8A8/B
QqgRxXVh7JKRtB9hBQRKcJ1oCwlZUIPkB4wgcZItAR4yEgkYOdl7trFrs5PfImH/
Kz9Ux55y1fe/YAFgUiWcDKJxitoUVORH+dhrcMgZkD7V76DbE/rCGQZerKK0sHNG
p98TQZzUSrGi2cRfqnT/xDHeAPiodBLl4QIGBKrJlR1YpheeIOlv4569Fo8S+W3G
aMxKR1CeA4L/4IFKsSt/yHN+a/mRlPreemF6a5A1NNw1uAJVWgnpWoKw+TVLHc3V
SoErn+6PKXAV1/DBGWksjr5eIZOy6eq0LqrslWV3J1A8BwXjtHJUkc4vM4WNOpPc
b41NB2qqoQZhBRCTGzWoIpZBuICZRdO8Lk0d9MX1oT7uz6+w2TjJky7HgoUI7Tbn
vqoKGt1KNXupQ6jmCzeUddfIJzN5DapzzXYwHIzyh5mxS7GbP8XhlcqkpzwA8Snr
ZWnOICHgCGBCa7AesAYlB70FbORxHGhyi3gq4frs3JlcKqHrqlgX4BXXHuxp5iys
5DAVHQoXRR1EL7ai2agyC1hAQuy8nVZeaClZe26S9EsnwoAcQMCiruc4GZJZ1X1q
0Eqq5AoPronaqMIyrJok7XQ9bV+uZqw73tYYF6rCVuc0sAMmYtqboG5k+Hnbt2NA
u5drQJcwiY2RsbiVoPfMnqaBzmlqSS6djL2fc7jn5zTrpzXqQ72HmxnmIkzlnQ8D
auDbn2w7/9y5ARbSjqVYIAP1oLMRfQ5h1mJYjVBfPJxFqZC3sNaDWU0NYSX2yYug
EVk/GV2jh/BCtS4bZXrd9BVrAiVk4qeQR4a5Rxu2034zQr6tmEYEJQtyDeq7fY8/
ZT4ZoSHaAQr76V4WH3Zox6dVpRpvRr4ErewcsU/9aY+PChfVYqZpr3+LCpe1hZKC
tOBXGatYpqPdsDDKJMzAEyBC4rY73VMw+xceAVmN+JbKuKzjdCdb/ImEYGZUPVWc
LSXAfNplUcRpJUnMdivdc9l5oZ6QgnqDRcwPlnHM8yqV/nl41k0n2/sIE3LiQ2qR
pbwJBG5fudWpl2f2hHutNLrAuwdcWVivDbnSNAayDYQ9SNrr6x99kSxLeLYQCa1K
y4kHzK1QfGNUuxDt2jG9MvC1jFPNRqkioMRsbtpZqhQqoy6jwYKCT+hYELmWlpbm
/cHZikS4HONalnW2oxHwfnxQdewyUdU9xis+yDGBaKCxvfkfo71LzCfxqBAdBNOT
+mH05mUWGY/Q8KoSaDjl7U3G9N8NvOMHX58Xb29w+nnt9D6AcUjok2f5k9S57Oys
BuesIrcM2shmwbiFXWt/ixG1H1D3cmnqZYCE+rof2c8rT/dMzUeNdJaCjz5SqW50
NERKWTaMTdR3AAJxO716qtk+IwR1M8qU0AJteNF+sJNnl6FXEN8TLqKCSiMBfsmr
O8n5RnKTQMjkahHmDOBMySJl2AEROWdUavLGgqxsLJISKqb+8bt7b4FhKe8HDdoO
VPU1z9AxmQR0E+VUwiMxAWSe0jvNgQcakne5lRKLU1t13tC8aCJdXYo6B2oAiUQu
nboP2spX/Yl8VUvxQHfcOde09SuwKmW+SIak2Qtbz3AVwJUUJVT3r42ndsmwDxEh
kfcKwxAc37YTu+sKyzIQkKbKuCvEVWhPbBeX0WKkkOLm9vhIcb+ZJSp37oakj3/z
ks7D+TkqYxMicchb+hkZvXoL/O9FehCvcu0RnwBSCme7iKhaulPlWDe+fHQia5QW
SHjNrPeEUKOvHFdZqUU/fCUCiIekBjuuT84eAkSHQb+GlhFdIRpiyqbSsedYWhDl
+ednrUH9Xt0y8QX8+GZKkmnIZE3GN4VTNqsei4NU+nAI+mHNGg1PK4Wd3cw/Lt/W
C2j6NHyJIXnI8TCAwy+kH+OYdn0MdJppTiTCcaEMSVAevA67QDKQX1SG4EsxIORt
AFw/LcV0m39ZHJ+wCFeGi+ZC1BkpitA3xdROEi3lkdMThAp2ttIS97daFxLDCgCZ
I7rbAjkdH+l6uuqpcHnamDxR+UEfeUO7r92ViWs70zd6dysEyxZVL0GJnGoT4rEl
ZpjVMw8dA4NpYsSFuBvQaR84+aPv3J7pX6+NktbkDwF43QaqUz++8mY+G5iu0tY4
cNWLG6zKnWn4Vqh7QLwfYPUJ+za76ajdJky1X4vB4QcYbQI+jE78X2rAQ7cStUns
BW5/HBPDBWTBJso5JruY8BXr/lfaAk3qLlkY8XgJyEsAFq2GMAJCTPmitzhdMige
QzrdVFHN6KUfITK7EtJ0r10XzJafqEG/EoAZI0mKmDYqexC+QyDhTlG6IcdQl5fr
/dIaiJ8Q9uWzotLYA6hNiGNjsGC2jt67qC9CJHhFVodN4aCSzdOXdQdLmcfYawsx
KNQrmMwaWxwTPaLB2dkOJiVXyN4Jg7X6hGGLUjIERIym7BryKwo+39WVnsDqVmnI
rvDhC4zIfDMfFnOoKlbxSN7rDeC2/AvXyi9OpxXPJ//03g7GKmmYKhbRvcj1d1rd
WCVpnT/oPgqYBCh2zygLGMxE+aR5ETaMbpAzsGaTkC8QTLHh2VyFgB1ztSl0B0Ty
TOv58DUuUdxCZS/ZLSX2Z/IEFo8HjmgxIzb7fTPT63f46B83NfnMUuZYEZPNqVlR
Jf+vUT8Md3SqQyeLiwAbO2gT+CTY3DKn5VWSDrqI55NgdAqhslDepFJs6Ju8I7IK
DZ37yj6slW68e5pK9N++aHwegYLaLbzA7ZhfT+/nDImd3VfEl0mcFTjJlAlOktfx
Ewp1Zoer/tydK8OyNRR30byUbO+Ee2ugObIus76z/bOLJ47rzjBIbvuhrWOeY1o+
Ff3oCWHgEHJ+WpC1pWcH/2lh/CrIZdaWDsuDTOj3pI9ovgsqn98cobE3n/pyacr9
rJWZV+p0hLhFf/Ke5U0vaArMROtR39mp5SzO7S8IXlyFL9nBLPvJFWzK5KRMCEA7
el3doO4jbep516FiYE9DopeUKumQ12ynJDz7wrmZtiwhNpi0RkGeIaVjJmYN0WMp
F4m5kb8U12DzMuPGfshAYrKzmuAxXA75trKLX2EAsSGrUwNxJmDD3GPKJNdST8ik
WwHhnLzyKgy30neQPPxmvh3EW2bYYJIyRQdqqddz5wYCbwn++B2uk/ysDV59kHyK
x8hDuG+WQAkcLosnL9/ITwv4hkRzfT7ucT2oMe7ZKYWZEo+rQFAT/LlOjqn+ULN4
6AfQoGsku2xa4OwcV2Czn7Gdn95sE6c6h4hSopSwK1wPkFBRsOnrtZyqrKaZTxNS
C6OBwnHCk9G27hIAvraNGi32HNFvxd/t1bwv3TEcNlsucsai8zeJNpirgG3HnbLm
7OMvCDqQvxe+S/MijIM/iyuCYTOTYs4fxOrzaZzNhOzEJTj6Jf4ZQaaQkCGQ06rv
er2FXNE4y3Fxk5Fylu9mm/isd6Ew9bBoXNDog+lL+do=
`protect END_PROTECTED
