`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOH1zw20Tt9RCI4dtjWlvzaOYWkpaswPkrurHfZJZY/WvV5gKIV7mFTRzdW//VS0
HeGifJL8xWXhhx6Hv4NdzVEkzZao4n91nczfHYQBvJTPd6+JbhnF9m4OQ0KvEhh9
P1Jo3QCBT2snHD025kFYgU8ygOnliuzWiVmMV6wt/YByyYWoGpfR1/gRwz+il/tF
vU5Ci4DAtsaCr7aWJr7iwXrYf9bBO7Yh/H4/PiCXKubXRHSWZwYUZTPSX4g5lno6
rIUi6CzoZqNoOamK9VgZwtaaxgMsuGmJpMeT9S6nb0b2bjL3eg72j3d+n+HlHJGR
kRrrTYDSQKq+MDwXoTXiRl5vyOhsHvkppDW8ojzaTPsu1duyuYzXaOHNExMiqYPt
StIBOEVKY0Wk3u2LvhL8pg==
`protect END_PROTECTED
