`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asUytlzPyOQcWkezka75XkpepG0LZkP+douHr1C8PsmqQbukmjJTaqHuZniqyJs8
EnPETR09XqYR4I9uP3BBDIxP5CAq+bNbffM+CSRVDWn0/K4tYSGH26LQg6jAITiC
f68Pp0tWgbbH/P8Q0mF9WEt+9vyyFMiCyGHNsPqdehEa9Y0YNpqKg3XZgDs9s6BF
zLsAk4ppWcmJMqgQP4rLmTH0ZpHFdd8rPi+2N4BZ2kFclWOF7VxmfTil0QBPI1IL
7ShVbKkFeQ+DyUe5WA9/+rtCNlpDdS5MAGYP+bi8pDxYpbFgFeaYAoMTnfEGU9OH
L0xak2KapIRU3WQyLLf1gH/UcGvtFyIwLbtPOvjaa4tJ0+U9EfrLhuTsyVlo8vwX
tqWDcoyibw+LxNG6N8Tyxr2nxYVm0RaQW/5idhXl1EHYQqu/sQvSQo8Qosm+vdWu
3bx7Zap75DbbuyD52PSPlEXLlrUTVB/il00dnPmeYiOoFOzDw4xdBKxGEnsrfCaf
PfmqfyKjhfyGKermcQNUDV/vEZA0JJ8pCYw29xXH+LfBmqumPILUKgDUdHsLKP/p
k94iELraHmvaLrb1AMLVrMppLu0mJJ+4V/lhpHshbBmDmlDLMmtQ0j88GxEtAFT/
Nax3AFZ4fM/v9vuLfB8ANBxnkxPQb5LxBhw44i7OM3qBuuW7dM6462V0v48vPPiK
yi5TNqkxbGr0V3tbOSz4XIaA7Le2xBNuV2xrRsXATPqQz3zLW5NUSpsYfV8aeifR
EyAeh5h8ncHM2qjeumrfRbfwM/PKfAnPDb88pDAR6F6P1kH9xMdhEvnkWUB5p4iU
aHRm2uTRW9JA1ObIAQB7ToYw9/aoKUcY77rxE2eBq1BWV+/PtsYmaIicGzNQvt+h
0WDJ3y+gX8z4dc6mBYTbpXb/b4ZkoKZFS1QDAWLGu/I=
`protect END_PROTECTED
