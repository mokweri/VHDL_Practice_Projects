`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfK1BhUNlgX3vio6VylI04jTAkfMn+msiNibJFcACRMSZ0xD4VoYGv5u1KmCMefO
AWIr737z/FnpstiBiCTCmVetBy5y2+KVqoAAgOMJRzklpwQKzGQoEAEoeV/EaBAO
u0YrdNUMK7osFsCHsUA/k+d9G2UCy2a0/7ZNUpCaBSBp8+e6yn7WE5ckBAsaQjjH
Q4x9RQO3twMO09nkcxuXvJ+0Lkm4Oc/P3eAwxBx7cGkg5nWt1OMWq2+lHu63L9MC
rgii9DmvtpJMqSh71n5SSB+IYDYC45SDZLoyss7bTPBitJNmnBZSrABaM7vui4y7
6jQgYtaUrMBGfrtrtXS3XLmd4FfdvEstEwV8OfwHGXuMTX9+JSo7OYz9coErP+vh
uZxHzgY5BgyZWJV4TW1rKG7By2zoFcJqbdg0nWe0unJPVYgg+aU1L0JMCMlDsttQ
FKXhLDG2anxUAxU54VAzzqPYho8Y3ehNZT4RqacgvFWKaE3mK8s1IldW5Vqzr3j9
wxZq0mrFBdBR5zD38n5VfR+y6yEl03/+Uj31X6ozUpPz9+MvyeP4nO/O/9KgULQY
avIa6zqDGylYjfks3JqbH84OxLsyNzaXcj6UQV2ma998dj5aCt09twNTzN4o0ywj
nHwCoPTm5e4SKxzF+XJB01F9/PgRxtMup5IZ3BkVoWrsgXrGexESHsHF11wML8VG
jBwpiAyX+NvzeBsOPP8Y7qq51LtJIqO0spBShwubiFTB5TZ6xkqzAe5dQybAu0S1
rmb8nerGGlji+Bz41zCzdDkUCopbQiWiqJP+XJr3gSCSJlAvfvBJ5pQzjZ/uTZID
0Ak+8ySpPwEFttTo4t3UML3Tbd5zFduOal3lHTt1HhrpHnZHA8jlpeTFp2LZBgOw
niBKI7oMegdoYMIZWn5I5eEOPBEhQrcixA+yt1R2B1frzdt5RlxPgmfExoLtVl5+
GGYH+SZ5MI3gGc0F8iM2M29g424Bjq2g3e+fZzzCVwxrpUivgJd5JllofsGiO6L4
BoSgHnZiwQJtj1R92notU6Th0Q3FRxGJLpm3GBsdfL7qKIUNAQ9KElkuhF9WHXAT
i2vCxrrK+VbDYvIp+eW8GY11/jxasAzfN1lq/MrzPJ8Pg6RPXPbOf+Xy98+T5vLM
Fcx6zqMFYophTyUQGRUPjJg1TAW9ZuhcvkzrNS4SzNFznHSMZfwFFAE3S1E4sx3A
0EHlKPDWkF3pgL0dfJzxgUOLMdtUlwhLtQf8BoqiAzWIuz/V/33BrUO4nrqtkE4q
5xhF5K4Resmt9XuMd6lNj63AUHnZmlY4gmzqEU2+S404Sj3yu7tKyvKUtE2lds/r
nY3Duarj6DfBUSJilxa018RolAlxMfO+x090qUX2MOp3PmJ4m0UmdXeLivpv6Ak7
qOxJWmZPab2WNhiYFoKHGrBt6YKPPxV4qiuzDAd7vJ6Deb78Lu6aGOsc4FQxKuP4
9zEMs/7IrLY+lFKC/yRTXCnz9MKUk9SU72BDudcRPNwqDFK4sfMmAGWMnoilGXw9
ySn2cZgDgPXmTE6kF0wbLtZ/EMLO9y4kK25zDCg0Qxr4v3lx5/gdoLLEL5YMDvEf
UnQUhUPekjnkFkUMArfipNP9/rvLhrjrzGYFm5b3BLGX1NSUKmn0S4/9w8BTZmI0
`protect END_PROTECTED
