`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWPHNClM7NDtiu8aYmrMFB8nUWWZRiLVwes2+FVHDv6Czg0wwXnoR7UC27VLgZXq
kL4kp6Y81kLA/MnFYrpcYX09UXuoSlUg+rwbsi0NSy3oPp/E9KeIwPRu2XBsIXsT
xdpr8StZIHCytxXGDn0NajOJckc/TCfTD2+oV6j4twUtkcvHMa4RxKA3BzVg48vw
iU3qUWwnaEnYCwqO8Bt4D7PUtchpgzUdMgn9UxjACQ/4fNgUBp96zO5SXtxhL8Fs
53DKlZd2+5RbXicNh2EjdSMmb1Azg3ZzuI7JPrQjrHLERKfh+zT7B+RtXo2XqwWn
WBGUGg+bBSw1YcHGNGp70p8xW1ARuMXTBRqhomIKF6rjrlREcN+1y/BgiQykDZcu
OYhazNnH3EY0EHV87FTrDRvGjs31yMyzFCTCJWSGzT/sDFFIRhu4oFhYNbFYDEq2
HZ7UX/PA+qaM1Abfj7MO22/meK0QAGM0jYW5HI8l5TxlOQvit1iz5lItw9m8nPnD
`protect END_PROTECTED
