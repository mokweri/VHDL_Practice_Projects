`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WK7zhFZllVjJ8pIKS2BzpNOOC52I7Tgq1kxG1HHSFL0U9bjD4HEyMZ81iSD+5mP1
Lgt4iTkXkgnIfFkgrtpcs+6qf8FuAZN7gV8UZhQK/43sXWvECLKo7I6SviV2c+H3
3zXfkexSBpxpy+5C4CC36kpXvdwM+AwIE17+PmDDHIgBIvZNJJxvt6W1DzimWMDh
Vuq8zHHkEQZoAw7vj/f6Z4JKq56DXPZfCZGM4QwnW4J2dwRjSMoEgWw3fOL+H4Dj
XjVIReL8RIzgjQev3FbnB+2DqgbRC9yUqy2usXii0I6EDapsLt0rQBynksbCXd9d
nzvjSsdzMEzKVRfxZEdjqRcI053g034efeCwi3PmhZaXxcmfviKsA7fI768bb8hd
6vmc908czb70V6xv2ButE3l4+dDH10wkJdeJgqxXU6BkQBW/6J4pG2pR7TG+td0B
DsEcv/YKFAzR1m/R/amd9JJWBwag0MedU6UMT8kZLWp1BkR6K2d7EYkPC8GfhkBo
zz550lZoqxnv5jnKbFZ9tjYgKJHEtYZThCUQvACn3zNZG31MufiQUl60B9yUhCd2
ZNuFYSNxt1/zJOXaP97GXngHuYRy9gPVfVy3ZfjWPawC2doyhlb0EU/fDyoK4ueK
iyEKY/aGInuKwI71QH3CqwSU2LrYCI9lnhEpbJQO1wNPfYV0kVPp46O5rkUs3f2T
bYhGzYx8Q+csiyFEInzYfhFpJgGjhqr6gqDuY8U8J5KCr9De2fJX7a211gwLitdC
CbXBp59BqIFy86Dy1NGRZyDCfbdkD0oB3FilYEntUd7EriuwLmod0SP8QoRXZKiB
uyV1aK7EgpB5Ed9o54rZVPYkHhTb5GgACOs2MQ6qrGVddbcnEmqaO7lIgcIG3mEB
kmh5D0oEulJ/P0LXYBEx+knuGHysQW6XP7qxNeFrOOnjI6Xg6ZLq+T/m1jEYlHrj
`protect END_PROTECTED
