`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F78h5VUc04+HEkiKzlONwKxz9Y5fy7v9JyOIS8cOyHEDSxgZKbuKQ+quwdPZEXPe
HvGhnfrBjsDF7BygZXA0qwf55wzJeEpTGzLA/ao/XJJwXymZd+0cakqhYTQMnxRl
/CWGTyZxfHr9lp5CUxHLOWHdPClCrmHl3rr6+cW8As9xZ1Xsvhez1QI6p5l7gLcn
9pGOHO/ZIYxkTQkfBN7ZhO3q/7M/C6cd/emrmzSlhE1so3GNkGV7h6eP5OSiKQYY
mXnWgIu0/3sLA9mAnirmVs0kYFnfJO/psEszV1cGo/h5Oh5AYPkyLpaH+ioAbrZd
HoJU5EAIp5ByqVfxd5laD022DY5NHMU221piqPlefDgNkdc58AYG0qw+lSNE1irU
+lNpAKRJCpVVXUVf/CS9Ciri81Se5CS2YBN5tm+7FjkwAYEvP4JWDcXajL6DO4GA
8rkNJ5yrAvNcX1as1nJo6mZdPFSe9iiAItPyy+EgCawcCk7ugmTjy8wwI7QOMuf6
v+KF/GIGETp1cUM6+36dTBu5drq0dDdBdH6y3sFC8plcf3EkNkxRru0ujayV7Wwi
PYKhaZMkh1wVB+txVwdZPaRExVL+29LxqeTnaJjnq47Hox1AKemgLbxm8f3nnujh
KzQfOgyNkNGObDF3xNRa5ivjvEn/GAYHZtyAq2sYGkQnVpyA4m971pCaKc2uTRvc
f9fg0E3LNhyVGUFJIp9zwjYufLD3nfR6kiwThGYJ3rr5vbDRJwoEUy746Jv1Q0wc
4Nh21fxqhOsTt38OOT3wO0Xy9Yb1CXaRAGNtpt9LO4mEw5mqvQEWHqiBA2Kt6ERR
suU/LQlf4QTM+QrLNdnQEUr6K8rrMF9eihiNSu/m7MrcT8JR71SzyVRGg8QcbFaH
/3+VPEPQZRgCgBA5P+vdNOwqccBbNfB1MrQhvQOztNQt9kxgARMBn60m9ee9yqEw
KTTtLPfCA6hYpbqNsCKHzkGqRDdTJ97XmKMPjq1IQrFp7eBFqIh3FniYfRZ2ZTCE
/JOc9Gv+s+AWT2p4YXl/VP8HHvAZbldqkn7DtSlqwtYKCXI7GP0jJhBTxTSS4TZC
zsafs7Fa0JcEI+mKpnndawlpfs+nOKOPD9vceJqgVGepkIqUC7tkx+bTkk8djQK5
zr23UhPwLAVXrU1bXus+AE7JjXo2fX7PJpluISagDY2YX+AlPQbCG0ea6YzIR5Eq
Tb5iK0Q4PjEhyerZn1NZkgUnRrOb0+cZ/NgL2EVcglrFGUd7Wtq48P0zVF6Mnfqn
eMk5B/FptlaKR7Vt5tAAwsirz0T8PuajOT6kTu4w7Uyba0veS95JS84GfA5o36a/
JXh+1lBY3Y7b67YFOje76B2+hZwLTCeyVwtHOZFf8J2LMZZmjwWeIYJP28Quu3Ir
LqJZfHYmfASP/u+yHQvquiRdvBEVIVAdd93ZCmLImZP0088uZYjp2l+JKRQraImz
Z7maIqYG0Foh+kkkrFdiSBsxc+DJ3x0dHx19J9b3w0YTRgGWwV1lBDCrwaEM4Cxe
xrOWy1Dl5FwU0/JMaCv1ich/qVomTOY8DOjI3xKThiLH55xTna5A8smneHC9wdmk
+ZzVKyCBxR8r7f/4gaOtvxaKFfH3bB+CosiisnjKlxVy8qOvSQI3FfOxvtn+yKZR
DbQbSmGY604ruGvtCzPcbsxwtvkDGBdODoVXybxTDTYk2Cnsxc7/YkbWXhSKHLvN
F76ny+p9n3Bjyqp+5Ut9hGRWcm8DA7a0wlYc12a65/sXslmKe5k+RKfSrN2p+fc/
AKGGMlf99QKYhMTs+17OwwIJM+9U9X6eWhfGhzy2GFcgQtC0TxG7q6M1/0Gea1M5
H8UfiXPlzN4prVQZBsCiYvkOPcS+MWbN/zhcTMjEE0okpcJo3RigDICYHwprjCUY
kxa8Y1oFm58C62EO/+A8wb/pPkNMA7+LXuiUzLNR1aVmGjYIybU1nNBKjcKHf5LT
gHJCIFgib/GqnBAWusrn/VoJ/dgdr2LElpxkkmG3SZwoBTjy+eLcJh/fbRKUw+tC
/ArdnTAyYzB9J7iXUVLQT36PHiZEE+VrXYL5XUzoqiUR4Euqj2XU7LP+7M2bg+Pe
xNMxekhbvNk8tYJed2U/aihE+5fSvj7fuJbTG7TOHEQBYmgZ29QEhJmMDNCCHsKl
2aT1004XLOA5HNpOZZrcFNsadyQF3j7R3bTsk21wSTdIRTZawXuAvMpGdZe6S/I2
g9fltf5lvZEVjYPrq22ytldmnOZOjVfUfMtW9DMhXiLevHLUFPtmV3mhThs33Ih3
OMxDxrSjLMSVzflYxfU5YA8U1Yr2HtK3ZTEQrn7IMVDTtDTLWHCpv/tm0EXwbSjt
ts3LVNnNp+de0Gy8k+mNt+ODCFM+HVLzIHEIiEQYnG9JvY/5TfFjAgdXo5+ZO5WS
GRXYyqWKR0FAlcqpiVKcst3k3BLHXgDyrns3E9tRsexuBx8qz9qRYkj1OXAti3Z+
Psd71TwDHKFbpwIPzbk83IoR1PBPglYYe4JmTXWJfsSpVJs49MWIwBjpuTJzC0ZN
SlTw3VogFQqnRh69ydGhtFqFk/sz3KRdbzfItvMa9iSBL+ugGSHPV/gWN86zlUsZ
BbNN+UQFLXIs2Z0J4qVlJLjTGsfiBURWUoF210wgrxhW8KkIDvl6d5fstJUYHXJa
O9xInbfJRg2sqGHvaWIplp7RB8yv7rlHaq2bOSRF83EHlm2NB3iiPcjGgAjKF92Z
6qk2g9G9oJCBP0N8qgm+1jjOtECWgwvwZ3fpGvnRb1Kf17Ke9tfQufIPypeWDlaY
0FIZPJAxvZq0HSUZ/b+lbL2k075AhWSaok6mxgV5Fq5vL0mmzoNqhHmNmsw2349c
uOYSdUStdObYWh7nzxtLeNacDy9YSCo377mPcCrmoEe/UxyA4TYfDy+TeoKuDY+1
C+iMqJC0+SVDWHx+Bc7kQrbiCGCHbzo/O0bwXfICSRm/CmqXiI1+2kzn/wMlANSU
fnDfxiamAbATrLDWVSUiIdxaS22W4l+vfX9TfaX72lo0d7eiqiCJRpYHKgOh5IRJ
BT+VNAa/Dj7Yc53RyQ6T9hWNR6FRWhx7fUU58npR0exXJoZT+CVd5jQChicS4XI0
SK1XRiH/ZpHv4rERYDh5OMHG3rj4ynyfX/ISsPSYs76miawtCYI/uD/26KCpHlfn
E+OHj5uXDdv4emWkEs6Ch6RmXTjIyTOsiIddsDDpipGKhZu6HKsygquTuODH5bBO
Rww2OYClrIa2osGJZKPkRj5h/cnQ/3yfg39KYnmRaFnjUVqRYtDpdkJXz1WCsSAz
wua7idIj94Ukgwtn1Sdkrl3aDeJXR4+1mfEV2KKOntu4ogiBQgftdiA0Y35yyB3T
Ie7Ocg80YJo4DyyXhIrD3k+yLgaP+o42T6DOq/qK66kzBCZ8ikgevkuQYVcHqQV5
nLNky7P3erWfE3/FzLwEiggb6R7BM0/Cg4XaQH6pK/DWY5GbehVmrX009LL3HrQ0
c0O1H+wD1/Q0+XgeM2C3ZKYeINkY5Bx12HfAQyzaEuXGivSSER/lsuP73AT4p4Ff
m3AofYdlwNqbwGaQzv19/10azvAgwRzcUtc2O3htlwL2nRgPAvhF5GdeCKQU6Tv3
fsezjexyyemGmqjwrxUAXlRFVuSBDWe8utqfdtHbYvI2kRDJCk9ZJS4x09sh84Ei
m9YQ+pTYAt2G2mZWKADR0bG8hXBMaLvajJtnXxBj93x6BiGny+D6BLZZNi0+Bqzc
pwcFDCGxmlLDcfV6u/5LtPifLbeFKQ6jM/8E9oS9b1fLsVXyP0r6e2VOGQCIRo30
W2zYrnS5Wxd1gqf+fMVL0hKTJESqBn2IO+oJf0p4yGvesNcyQ5CzJjEM/91n8oMG
QD7lJqIIVsUoyeOnuisKBbFMNsk6vaU8LqOzCMlcK41bOTMDZkcMtZpg1znJb9Ht
58SIIS56GnN508kRe0LHAQ+RjQO445ml0lKhKKhIgF2ug0T8x/0yETrCidi6jFLr
N/Ah/dJKMX3ioWmpzfaypyKzBEDEFYcLi/umg6tezoh9JAvVPb7m64jLd3eKuwuk
/p/9wpqZ5+yDL5REtvFqLwPEqrU+o+YzqQXCFou6RZKJIiqvLBhpY+RNiLVq2R8F
0mHHCWdMRr52fg/KVBAVPIlx2xXAyraxYVGs+TBTy9TisA7MUlYwQANN3xv/nL+V
hZ+wnTdvP0sw1CPHYF8YNM4ooCYxGJPGQtp1rAGN0XSxZjif63/JyshhrxgUh4YM
otvmibRvpaZUqIXqLVSM/TjGwNqlR44iydQZiS38SaVanpJ5uFmGkzK8sHdxXmdS
cNMTZfjkxyTEODmMAzwJsEMUYHCrusWfvU9mJlO2ZBSNHlU9WNJ0L0+Bp1jZJnoV
whMj8+HvHOKnxCbNhf39lazYWoJedtrQaeryQo7YEGHifBUcScufELVXlqMhVirp
7hOZHNcdUJ4SX06lX/h7GfxrgAw84I4NLr0LrS12oP25pCJppemqVzMpna3OkDSR
YiJwLYM0LY9AmGiO+kF13ZQqPuDSBhcBMqmJTMK1OVE+FsbcwZwFpE+mrMNuWi0n
FLwB0/BuhGPGZOWZmaE1NXfTMvOTtnDbvyrzg+U9fUeLrCfrAu4DMvLiC4mz/hNJ
gvo9SdcyEGT/chrS4fMtYC1y+wQJKK0Cuf3RcHWe5M7SPhMFNQJ15Mzh6aHvNiMD
NBYo4+s4GK4eRIYvCSwsD1J8orKdGB4apkxyd+J8/TMaAQ1Xio2MShuZspwb9GP2
4fOWlP31fpfamKCth7ce1tLQg4ByEOuRM9I/0jNFNZzgmlFwHHmT3f5Dxut6qAJj
H2xSobfKXUeE8YO+vMUdGF3UDDrcCf5baYi4zHmFp8DK5i+lT6RZpMO7JzcIdU1U
X55bV1CMT/CdkD2DRCiYeVxnnlZ6wGYc73b/8O4Ese8cfNHD1Ow/6nD/FOJGd7vI
EJJWeESWbD2JWLHxHLp7DgWU1JGbxszNgSIW4proDcG+WxfWMSefuzghTueiNc2j
Pl6RS60jKTm979ziyJGuj50aVyHHAxHGtvJpKxcYGTbbHeSqEjv/tGb5Bxzi0mJH
1KrisYhRUZI1pQsbn3dHTwT1gH6Nf/RA3fNT5IRcng/21xS8yFx6YS3MtHZ3jhN7
ZFbC4rxk/wUN9nG/kSK+X5zbEncKxs2wCM5tw4DdsXUAbccPDRPpZeC/duKG52NF
kSEXGjEhscHEbwMjtZrgrNwghAWX5/C0+v1e+Rgls7vnmHfRL6+xZbZjOlncA7yH
cD1YXP4MXZa9ZRV9DmEYkSNKdpITXPND1QcE1XXEcyVcihZlQaw/QHXEooK9t/vA
S/nEjeY7g4sZbF3/OSeLEQH5j4cUGv9kq1VxXX/F4oS/NTGofJdPACimbZPgSsdg
OwzHR+VJ0RvpKLUk7W4sUfRio3Xj1UNfV9C4UZ06M8qCUGhFYcBMuRPzTSY6liyV
0mUdxJlATYLvMZDAgexcb+LGY3C1k6h9RcnVDTRXgUhvI7ql9K0AkO3Y6tVaqwOU
1tFtIdNTyMOUF+AYhQN1aWaQ/Rd0H9f3gZJ1HncNjo65n7OmVhvEf4i/Zrgbdcl/
bUF9Jj/Brj6JaO52UWmoe9qeih3qjS01XTc740uIn68YB7NQ8JOQjeCurACv6HR/
fO9fKuIaR0edkzJnqA2iYBsQkL9B7ARyHsIaGsSBa6rswXR4D8JlO/eG58Oz7K9X
sS4xAlndFqegn+SfAvANVRydO3QWNaG6x1WKHvPj71dmFgaylsIyXt2E6PO75aZD
Ok5AMGdESXH985UsdkU6smREVNceewvlvp+33FTQGQ/SxPPLKh4+PIQTULub/ugg
f3+cCGry0Or/Z5NhGbb/LRKyIxZu9tTFakOeNxhIa5V0/60RKxsvE+2HzuU4ip9B
IfZt3yOKL9QV4asuoWtHD8XIqeDLRSAwk8aRBKLsCVRLcxnXm8sm0inbpGO/ByXL
67xFwt4Ed/w5LgQk1yezLQMsf2dD9mHKyRTHYkQnF2s=
`protect END_PROTECTED
