`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qB5J0KYn9voeKL+VFkCcZ9+OzYPiWiuW5Ux9ZWjJgNX3dRwW/jlohZFq/eVpArV
DwneuEl733MrbSOxnHO5bWSDJoYzLTJOmRgmU5mcKB5ULvukM4JLfOAzRgAvyonW
gh40N6v9wRYgkfyM16HmVk16PykP2lAKdlT/zLccaDOK+ggiReNNgdWEqMI2f/rk
JJGXjDc6kuS8Mqexsek9kI98Xlf/KjRfIkC9IftzHD+s7hPmoR+zZT129t+dknVB
N/CxiD25ILpfpOnGXXETRMHnpEsbUg0Uxhaj7EIT9QOarKfxt76KYzFavPLhxN18
YJVsMkhN3alPwrtSPe3TjteSM+gPYWKvTYRKW72OlU4v2n5RgSVCBSa/tF/GOD8t
9NuWte099gt3k/aV5yO4qy6JvHC09dT5krsKfB87YUdwal8Qx96vaFeJxESjIbDf
`protect END_PROTECTED
