`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naDH4xDcR5FSryoS82bkDQgdWndK0gd2nqVxdymZvDSR5it8hKxbpzkw8yxwUtUs
qzqw2vtU72iqfIm23vzC75bOcoZMFX0bOeIEzQhgwa7SiSxKcNXraCWmoUA81Bfv
N6ZUt1KSjh8ijg1NXSdKpbgueVnt5qANOaMo7sLYTYpw3FX7CpBHPieBZdiVZ8vb
JBsABNQsTE22A6lDGde34YpFlvtufDI+vKWrHDJ5k3gCu4rlK9Wlds9U3mZO2lTu
Ltd57n/oIlPAT/GCWYDGVzhcdw10cjmkh1LjIRL6OOPMRKVkYDUIYIebefl6YDuX
ArV3G34N2hEcq7fYeKQk8nV5VfGBqsaTBdeBUopD3oIGGFeHNVzbtJa95YncsiiI
+h+F0v8u2fZvliz9tkAcJAREJKjjCjuoxFkDoUknGzcYOEFAEkQuJuEXGWfOCz+n
2IduWNtsQNfpi6lhZIstUXcBsdxorjkOBFW/srFuOQThbdmbAx7v3j+ovaFs7ZqT
ak2tMJ6H8808bCg01yI/NrOd/PT8bE5Mmhwhf9ReaXFFucHq6kAtpkr955RHeyLI
ll90q8nTA2cW/wRDmtp4CydqvOmcMZA/lGb1PS/r23mYCkA44wL6OcYxmY7Xha9U
zuW1CEBCs0N1eK44pcRwdKjhb/fGHCYWgPpmf7JGjEJobkyhe7G60C10AiDI1DYi
bn653wkrXtmRb/VYRjzNcKONTktSwZFtxz77hNy3EW8oIT/ks4yi5cA720MHsWXv
B+eWqSbe5U5UR/JkzaXWM3PA1ciuIv54mWn0kpCjm9Z76N7yEFwt6JT77cbYKwvb
LUdOV88JgQd5dkgKazfZ+g==
`protect END_PROTECTED
