`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HZDT+4xdkYyLrqgOMDsUaQaJFXYa7zj2X5lgS82SqU284HzLKXU1ZKtkVddVz/V
ehopLCMfQYJDLT4s4K6CIDW95IGiDULBrg3oRJpe865a8HXRbH292AEgUe6HEPOk
o4IIMYaskwC1min//f2fbBlfoJeZGenO2tR5lspFyCffO3T/tcQF41AL7CbMvpTq
g9jMRFK5wLx2sD4jDf4APPFvN26q8O6y8bF9bX1Dx81oNZcWad1+CM78/qKLc5wb
x+rV7pRMroe62vvB2qklq3KxNkripeOYUbk/LQ6p4wX9EnOXhrMyeuViZs8jDjru
MPmhYjuv7kITjSHyVrZCAxRNNSFiVeFa/YIItcV++Jpm4H+G9wZR6SIiti7UvNku
9mk75mE5HWCiqekpI6kQaer2hWv6czJB5nTk3UEkZemjDrsLFxAG01ogMHVR9+ei
DH04TNv4QU8OyzuqAXYrbZXra5d7n5DJeuyoo7ik6TeTESuxBQQRj+Dka07+UEqd
bCOXfqnavQJY+sZcNdI5Kw==
`protect END_PROTECTED
