`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Obl8PjVNqWqvGVBf00QIKCSsAFTCjm5oawC9KZ92gCuHiNSwIdqkQkiT6x1lQLv
GlHQczJpnScOdP6ZZKI2w2byxvxJCVTOBY45ZAgJA5BB3tCLF+LHEFbuk1aAmrML
u7r2hp7kbKOoCAPdwDS+ZZ8buyC1oMpiJHmJJwzznSQuXpHpyNGsHq0NTPEs9wA5
sXWwnMLVodpSH9o2HJtL3ZS2ByK3gJLm+vEFvOyq2O9+TFaFT4USvDrtXX2X/uKB
cdZHxyLz1fiq22R5Egk6PBahE09HAFV3UK3dMDqRX9TLPw7POXmG5h0d2ZhER002
UNPlXupbqg32M+pslc0mBuDEFyTyMTjR5lxvAvgoU3fznCWfty8wsfmnNnp/mWZB
bgQ9kYkSncLnTyECv2ZXiEV8hfqXaz+6aXQLxiFxe9cK7uBeKTbMe6SAzP6VkDoh
JaZMQMiXmfWj+5g1Yu7P/b1/4b9S9MxhAOsmYVSulEdzUrivpmrmnUFF29FGRlGP
27N24ugq9ZItLzclqf+z5tjrjlORMpyH22bS0xnATfPM7yq9ZEQCVyxF2mxbuceD
Zp+5HM96FI4bDQp3XnWBis6ZIKAPasFuttIIQVJjFR8NJLhdQqGiPpiFuNY7jDNj
aE0Iav8y6xDU8umO2MM4iCc+Laa7FmFPECJnJFtfGig+RGToc7ei81v+ZQUsAZHd
jmDLX40HMqSIsdqDbDU69WX4Le5b9OMHovthxyapqwjvFu/t0NmEt6SPevmXegwF
LlaH0GM+98M9r7/K6sOPaVMDf29znaJgm/p9vib/NcFRB/GlRzu8uU8x/K5ZBBY5
3M7gYIH5u9964tCcmUDc1nbmo3Rm38HxN5r1Q7eWc1PzBMsCI0tM7xB7O5GgZyLA
GAyEQKfidaqUjpaE9lS9ATXVU0691ho0E/McTR+BiE+T+zDAx6NAKx0kOo6Edxby
g7Aiu20a+IrGxznyMCKuYbOlsrqIQ/6ILseNKkYqqxZZWMEwVdoADO24R2AFGywQ
6olLQbbW9Ni+Ha5+3gBRj7x6cX8juZuhONiqCfCE7RN9TEQQE4VZjrh15XQDd6zS
A0dhxI1lf+qqZmEYm889j85pS1gVhrGD6XURSQrPi4le4c//ItBHlofnMltJu3Mw
luasELJfwF3bfxe1PET2o3dV7t192KIhfQTUTCfCFrYBwd1qYAK8xeuv/VpLMSCC
tBHzoTk1g6f/DDf35oDtaMin/QIEka1Hm4fiH1fQaMZXb8Nt8XDXU4NlCA4HpoyD
nzJJhDHg5/C49MmNrFmb/pLQHxq5L2xRccBE2o9yAs9o3uDOKNmlyjscnAbS9SOy
UVMpZjYukqLnsGCS6tdMXVAQogwMCp6+7TAOByvglgwk0lVxPoByGYqazouvN2FY
1Gw41ehwTjC3S0noZiw+18uyY2T8dbiVXclVINi07Sv725YOlyz+LaEKuJo1adjk
srhDk3dw0ZHcTRHuvTZ0boum+VG5bx7FlyZtulPtuB/dQAj8jicxf4H0Vv6IbDdW
m2n0Hq6cw7cGV4gAn1aidwGl14sM5bKPdgd8a3KajPm03Cmu8pxesMvL0hOXb0ni
E7gQMESHwlBC1CIdJZOzYtRv05cEeWaHk6zuh6GUlAjrN8jocJ4micsNgA5K0m4u
1tFd+122E7EvmFPbU8YYRHluKvOa4RrZ56VHTFC2MGm/izc6TzsEkqecZhiax9Gi
mhwANq1Uzz2zl7MLE3fvrjoIj6gfHm2cOvC0wp5tlVUJYP2c+yr6x+P4ZV/iftTZ
BYbWn8cKSt+gogjIYktXoRvNSNgrll9AVxf2l65lELEeYMl8h/fHLImIQNsIG+Ks
eiCCx/1dTGkqackamWuTFPeSHvamOTAp+Pm8iNRcgUay6M+MoEFqaazV+E/UcQbM
KKLHk1zSVSTFT1MEDAptcHn14aNwHI/5EQy7+klinqDVudbdgRttrlJHS/MAoAvp
nqkMSJgiDv7QUWGltQdlSV4ybr1AwcwxWVJpwvpdCZ3RYe68cj6ZK+U0BYZ6Oy8l
LDORHFPoScv3Gtqym9WcjQst12B+8el1keRZAvB4u6b4ONIBayRnR2VMnZDd/ILE
914rWQd7KUY+KWFfui1YmTKTqAyJd5zKpqTcVunLnXdqH2Ov9oU3Rx8H5sX1TaNg
32gIX1Wca0+CWfzrnqp2O+mSkEoJazR4sWcTBk32fRrk4z3zyW/DXMpLBNXrmJzB
Eop9XPBXZYQpHT1pPk7ygyDbvqdpdMRrtWUZwmIwP4Doyvor98KzGh/SkX72mcvb
1Cuk4mSkSMSX5kKYzm+vwFlxcjfchwOBteS+b+XPpoztxIme/iJgTNEFMIV8EMe1
KyQwIgYpq1hGslS+MEpUN+CZWENeKTNplXsIrWCozOniof2UDqiXJ6HvFLuTqgme
0XHCJ/gH12zjvsiGmLO1CG08S+IZXX0Y1mrY7XkXhQXfBmuHj5rTMF0ZJqdfrg61
Kdiu82/RvQsX4fuPeGt3/Ng9zwEFJibo9eO1BE6PUJIqQQaEmH/DzCNtm3UZJ/9t
yrt4bgHfh0baVH68kVJlv5mN2I3Mg46+Uuz86MQWXeKJFR9GIQGM8QKv3ranOipD
rzJfzVIMFCBW7Qdo8eQdd7IhP1JXXP2VO9/S10zO9zLQT/zMkbAH2/G5VPJEuiLx
YbxC+uvttr580b1kxuk3YWINU06tvGdHCWhXCArR86GqsDIQ+zp8gJ7XQIz65QSL
qQHBVTRcn3FzSZlrgdy+YTr7uZJ0y2pjDTGdA9u9ZF8yg5TCGzNRhxAsWRV2PyrO
x960Bgyklp5j7OneYCikqlUbPAHKpt0UmiWmmEjKetxf7/6Xptqk48zl+ZGhdnbI
RH6Y48OBSvBdo7Q15vcaU8zM5CO/f84S3nBM8Y7DpO3TDQNlXR8Nl8L+rFroYnfp
E/8s8NFKhq/biHzq9jxDc1Xh9DC6kO+xeiAM9MV1y3EhpesHBeIa4D0B5i6I1qxr
crS2J/Yd9tlBhNM0IzInvJtM4qhUIiDTrSH2H6b9Kcm/N+13iZOXuDk14mtvU0YD
jdJRunk8ahpjVHpNTmYMC04iTHtPiJH96GLo2RJOO21ciMA2eaK1nKLmtbFQUWhP
tF1wHknQGpws4yzn3Xqs4aC3ebGhR6ygNbqLqWmU2+C0hClrnjcG6UNuFJxDUsyZ
JIbWnDMQXuIrtGGbtUjfOGtjqYU3HmBT43c+z7XN4sJeeBMRtwqKHBZX3Pa7KQ5W
9QMg2FVQ8nd2NpC09jNE6p7KGTMTxysaKS6/fgIu6nUHvXUxXRvfv7VkHuPj+B6y
AYxSUrFGE4ANW0myACyYQPP/BBOKmZvKBTa5pxYXZ+mkMLhM90HJPhPYwE+9NUvG
+R9bu0u6vH39GSCyX/XomTKq8SlYSxzEnt9BU9Fl0M8ftii49hKdogn9GJ7vspL5
mHlNFhEOhD1GLTDAY1xpkLlm2Rg+Ma81k0jEqQCTzW72bZtpBbUB/QWeyOv9/2rm
sY+rQzqV6MJKmErSk/YfhGPIa9ntlT3cBpgm/BayYkT/Hv6mbqCNq+HHRUDYl7X7
/QA50eeRlLMOF4NiqrUYfLeORie6JYi0nEdO53EwvDyoE74iIGyQxDMldUKwUYnQ
uEf3pZQHLCV9pMOjj2G6bvyR82Ph5kz00sFvqNnGoLIb61T/TW5HuVOYR9PZE1GV
CA5nF+RLcep6CsXq388al9F5rVB8hxMojzlIdUt5ElSzYisVqdenlQ77PCJQYksu
7rT2iaV3OMRASq08A7j5FHFbo7hIJD8DU1bshy3qE3KoKfIU8cl4Wz3H67IUrDYL
Tn1h4KyRh6J4q99nR1E7C72U7aBmKxNcX7otqflUSWPsTjdIQYXZv/04+1KIJw80
lLAq4/QRtzDQcBqhhpkDjBuO2Z9RIL+xEdFtZv0cjA6hO3EuHFn4IhchVFstMRdl
zRdbvdZmCHGQVra7jMREw3sHJIgN7JernIKgiGRsHbEDUquWCD2xjzm4O3oZLkxP
4AgQ4/QBpbvceS+WUD7cHvsjaIYD4AKoahu0ZbGGaOxsIAEy78lIhXVsOdjx11xL
rEHisfCU53Yxa13E6D1zP/fMosIKbM/Jaj1lQ+syRSnmml7E3iq185Fh9hwXwng8
WjWqWA223HfYWTW30wx0I/WDwbxVr8nqmrpYtTymEDhHmMdCW7+TiM8TXj4x98If
lrWUGmOJJ1+L2k++KTEXGCftb2bLHCMdlDIkgjLCOvla0/hxct7Y9i8IuqkbpKYl
7/E9ODf8jG3EifHMH+V8Vfn/PMQSeWM+DzxzLUz2XsH10WULIAyejvuiO1xvN5Vu
rRQtbwutVR5kL0Rg7VeOuByZwESEZhUzaq4yYcWeCtVvEPOYt6bU6VKWKgn1Sr1Z
T9X1rH9eOIkdkI7LNYPwkfP4ucX5PaZqyE6lrIJ4iPELSYKfNPkBIOJ5C1D4TuYN
37x1WsxgTQdJkZD9cWZPnSTYBkb/QPT+kPj8tQHqRF6NnC2iNLWsw6A89YR7prTS
tyTzH/CiJUlp1F7muV4sQacswuaHIYRnnKgqUXh0kg0ZAPoSYOVcoUx16y5hkaSM
unpgmBJqccyiyplwKYNh7D1JdGq/ZW9NarNgFYdWGiTR1ygPQ1nVDt/d2e4TTEJo
Bk33S6UygNKAUjcv3FbZY4SzE2r2NdIdpXzZl8o29AgJu1g4OBLZhdrsAEC0WraK
PuW7rqGzXxSSp1WJgWK096RJl10EVajP/2MNtWFErwb3W7PVzLrs36ulhEqzUgVg
FRbQaH5My+umCndJVHJ1/XSbX7jMzuyQHwDauwJxyqYp2CeXFx/YO9w/iyP5lRZ1
YdGbIwSmM8GOJnMv4to3vmY3N/VFwxW8f8x6otg+6YnzjhcFEdMQlRhEIx+qUw2q
D6gI7EFBH7UScBfOxx8xv+Cv/9C7QGJ1n1mDfvPRx7E=
`protect END_PROTECTED
