`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjJfX5i3HNa2Z+nXVak2iCKB5RSkRMvCnJpjoUvDIZhza3qXGpmZxj0PMJORGxwk
8fh99KYdYs61I9HjtWeSDC7RjSXIqfzRtc6XNBcVb8ym+0otCSwuk16K3kI9Xnaz
Tzf+wT9hQlioICpW8QX9leyhrczMFkmPnyo+BGMWK+kmsgxQPq/ZVTNIxAFsANe1
KT7uIdHiRAm7vT/43Gf3L8uRTWzQVmIrGY/U0/bBTXDisbnUsdcBCJgoqSvN79l+
EHccE6uuzw/VqdWdnraclY5dO27PNf6YD3VMVl67X2V2goaSZtM7A4+J+yd0DF2d
0/38fMa1mWuVkCOp6tDkDNnoBI8m96KyNLYBow7TH+f5fme1iTJz4WFdRzupAfwJ
fJKZHHFv2P9G4w9SC3AvzIHkkjnct6WilLauP5S6GpbhG8DsbhOi6r4eAHKShVuU
yOUBedoviM9dQgn+ZTBUfN/ScnJ41GG8q29LS5AeYTwgflwuMCHXUauCn7ZrrCcq
bTQqHWl7IepXa7IMzFPyhMICb401D8/rL+pQ0CAbyv4lC+BCixMiUpPHGaOmxg5W
8sSqyD5UxUhIdVIK+5efNvy1mIPS+4/ZF6mDd+DxxvvhwQy14z2L6R5aY0tMfBGT
sUgrlZnLbmeoLXKakPp/M4fhMQyQf3ZGk8iTdXxLAPd71ocpXEGudzXd0G6qCPvU
w37wzBA8vqimYdwMqbLZfIp05wvWpZuHHIsR58LjQkcJCwtsn3ADHTqe/2OLPq8Y
kouP3ymqNHJfDH8cqeb0ZLhyP3pOpIWFgBhpceKeL4yZxbnfGgBW5eqgzavP2d+3
OdzjQAnrPhjvzjCC8R9eUmwlK6ALwGcoLwq3ozvNFiF+o06wIlDB1ah5hoDwzr2L
QhN/ao5bMY7SPmAztMLhBHYIc5kvODkoUboULMxR0AB9MCYOjqkIZDJK7Q4xwWJi
aQQfHEmXP3lc+frj/cMr1HgpNTU3RFLALfmbk5+8IQUuvMogeu59Zn7jUuPi/qQo
6iOpxiNI1cbQRmAG34/nGtyFXv/yu60zlK88ezLv1m3FEqf3oIzurwTNKgWiEx3R
pG53vS9ouDzqgOgSZOZMR6hXCXho5gLuHCwHU5UcH6k=
`protect END_PROTECTED
