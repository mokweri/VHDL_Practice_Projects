`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcDjRp3EcBChAOD4QvsngSquo4T6VUxnI7hGrjZE5Eg3ifGEFBDTbpvOoD7Ya77Z
IQ5oUvWBYfA6O6XGT/5eOwSTf1KWHvqhoOm4rtB0HjqH6YiTdHmI860MZZgochYb
3x9oxCN63G0EkudOgbYausQnz1xoJglUZpQS5FLkhNjWn5GSdqDAWsmsSRKVYZ6b
QRAtrQYAA4RYO/m6lsH2QVUI3t2xD7avoG0bM2nKqbiOAg9DqQi2N9oD5GBkIk+q
BsUdEI2ppsYdH1QRegDDvENxtW348W0djN58wdRQ2k6nMUSriND3NEwEGDoLzsZB
p4ruV4xi8lzacBY3ni7V3i4K6PdmxTua9Ppp/4UVU0HevoNgOHeIDILkmFZlR9Bi
u0caGBQuiaXmqzPSBiNEXvVAsAzF+A9SOdyFm4l+zV03hI6NDf09BttZWJAoTBeh
9QvqAir43vXuN/HCA0O7XxTqXJH7rMFfabPtZh1oCqfJGvQXMAPyI79sQb038MmV
7vzwLMdmaLrDDzpJYE1vz5S7ynYkJV605ohJvEwmhLesAGNIsH+Rb4oabWtRetSJ
BlO03hNfpro6zR5fB2K80I7NYMAh2ltoXoqKvGYJzYO3jcqgIIxhPt/renUugRgJ
Y4PhpGCUATwkR+dbq+yi/t0rEaqCoindaE6s6y84cKgGXqo5kPmbfB/xSZiLObfj
U82eE0hqHeLwJjp0XT4MV4uAAwYXynq7Ck84wQd1LX2yS6TPt4vf1f/TX/8n/YSf
CFUSf0QKW+t1aenHY2rOB+aJJiTBtm9soUxzrG//vkFl7kGkbUo7UHUVnZj3JEyZ
LL3p9h3d8vc4zUGfuaMy8X3wFmD7zaWCN5XX7THDfAXEr9rJgL/CclqNFLUBOKHG
vsbYYcP3cYAmGEh9Web5TB0/AboW1/D7H7RMeWWvmprHpPagxq25M22LUh6TMm7s
NhnAyukaQYnH/M5vLA/V+DVDkz/tPuhvZrcqd7DIMkKxHcV1l/53tO6NZ41rixU0
Iyr8ovcWpCgQf9i0mJD0RNs8fbS5fBiTbFQ8/80aUUIUJeI98msvgI2W4ZFQ0khX
dU9TUdAzxyOWHZcSAlXVXqoFJc9G6xf0GY5cZDRZsVZgLRCJEnoI2bG6IokBQwT+
OBvhn3cX+64GjQxyrh7x3pDMM4/cMp6+ZYXS7MYoR1niH2YesiUUmmuqqX+wOkV8
dULTmt1JXU7phiNxGyHrbsid9CfZph+eCb+2inSRqYiB+kFBHE/AODXCdYmijoO+
DqxAkA6lCFX7v7Frd4HAb3YVHHqR+auENuCI0igQZt5yANjjjA8hYyNmcgFVYapr
E1cddNkC9k0yXUiApUoitlF6mIginme2z789BVz+RYFauK+eW8duCUzJgaJlh65g
82L+rJLY8mJuMnRjxuqgqxVDhRzTMix3lC/hNTpoEYHYPWMUxwhBNB7av3w6oOZc
fcegpIcTspt+5gLl5Gn3VZfpJijMxiyzh7GUiiKc19c1sqr1al8AVEgYjz5OKMVV
Es+9aJQDfhf4dhFJkCeU/NEcg4ShRDQrqSugDUGcuwe1saYtIq8RpNid+wozEM1b
k8Ipp7P8PEyf/H3rW2F51yojXKhiZR66A8z5/cyTV4CVCDKReSODSC/6RyJSluv4
Pft+h+1ybfY9yXV19ezE1APbGXM9T9I7W2T/KIbXA05m/z7smiNmGggrZ8H1Xrv1
9WyMkv188mIKfpixNqtOJ4gqAcxX2HIWTaicYCjB7i0Jj67rQBeaU22+YK9nRlG/
kgHZCH5zSLdZw8ILaOPjafFrj95ilo+Cb+MwvVNgtHrA0yQtoUS7B9ctN3PLBeTM
UzjrdYaiQ5narVRbWqX4/LgT60D9VxtbJEfJku4Ga6BO8G2A9mIiAB8hr0BsGse4
uhEzeHjHEalqgxBQa2Fv1YObd+oJxYXA1xqYWCqu6343aWPs5PBfchREuatzNIg2
pKndCVbgqbtjGZm0BIrsjOKlNiIBSAJ96JkQOAq69lH+WwZW82SuwOB26EVfsv0I
rfVKKAKRONYENhivhg7vvecsoWU+SMEKjMiOd9OJnb7ot/82NdyO/QiGGWJnsKQA
XOToFxumPbmnqeXOcFj+QrHNV1JkWJRZaQTaA5ONDoKYRHuy8eGb21RXfw37m7wY
uYW27VIlXZa0OBg0VqQabswIkP2ttKGuASFijoQhe/lZbP4iBwdK0HvJV25QxWG1
LndNganiOHe6p/Ssa61qndMaOrdU3hWWEB7CShihGzjrx8WtYszBD/8tKKH76iwn
zAPZQ4RzTS0wf3OmcOsp/eD3gbBq2oR0bb38ip+c1zEuE0wPwqNUIqDzK4E/Wszk
bluPsH22JAD1xtK1t9A3bPVaIR/6EWvtDU9hOVH0ztdmWYC7Fi84OytHiGd7tdgM
Qe6D8c5DlkDjkADgKrydGYSnUzIdJRyOtPiUDx1do1unlp4ObPUv7lTl9setG8GK
l5v5jM5GeSvaRO4ZMwtyU5GvyPs5ETwFW5ZB76wiPgPF9kd8k/o1dOYVuPKWtB+r
rBc1NM+8JeOTIle3iar8omMQrtSITWGMKkw57J2uUWBOAnGukbIJhsbHaTxwWlOh
pcAr0nhz/hnFWfgDHgsV2ZpAJH41RiAXCvfZHi8Nna26TFVLfBOSYphe4T9E0Dcb
K41dgagcwb0cUQ8fmh8dp6Ee1HDwy8S7f3BsstoLJE41IW1CEVNFsprSKt/XD6Oq
2Am7SRWMO5PujYbAibrkVD03klSOgiWKnYd5w/gjLvTxy7FzCWNSgNhVchwjOcTQ
oc1rQ2KrCwiDkmsq1DmTiVIAzllzoQNncJfH9q0wtr/pOvl4CnMsqOf7XTNJRqzL
Bz+Se/zU4WtTIZmlPV+MBKfivaYgOXMTR0Dhi557Bik7Vy3Y/CEWVLNucSnzdRj2
JxnAMMYCrgIbiWPsxMlxz6IEdoeWcbIdGsHVw3PjXMkqMheppxuPuuYyhEHYlBdK
MiJa3nCqC/eYPgFO+4+JePFxbNiJo4BbDQtuBIBNRo0OZMuCjRxgoqBEOcJ3QaOh
yGUIPjGEtQaohGTiBiB1bUy4dttpMPtvebHyT40uAMuYG/g41yAfOPDRhcTb2FAB
ObUeXCYglfKRWj4lm9CnO79eniuKbUKibxgzTiWQGKsgr85exJjvOa/YNdBFsc/m
Ddol8EgJSlfFzuTYUoTB4+cbpFP6QuNLN9XKH/pyI6nXCiOjeOxkLEfgd6Yd477Z
2lMBLrcho7OQjGxz8BrFCY4PwhyCjJMg7Y8nqOC79nqtSBb5PtCge/kB5o8J2LZq
65T9oHpQmOCRNVs1niMVJ5c/CgBImNuF3Q6i1nQNjI3zwiulRZkvCoH8UFw1/KbK
VTzOqb/jQhTNPndn8XUKJMTBW/bN/kxddBo8uJHz1Vz+tkEkYZMhIrcM1XolR/Ds
`protect END_PROTECTED
