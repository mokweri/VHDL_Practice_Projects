`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azaFzAB0EuncJmS/XGIilSMemKl+8WHNOFdWvV4TGHWmrH03xQ9/yQuzwHnaVG94
ZR1Je3tHJq4QcuP5lCd7Z71UUK0Ag8+r62IBDyX6jnZyBPq/rMOF2X9iNSOGfnK5
q6DVr2JDdLys+QtLulKcgBA8kPO2ejfbUa/8LrBWrf0iDke5NW8/WMJ9iL5OAN9O
pG6j9AuXeB01uicg79O1t0VGz5jyy0HQ7xdfZFvgctc8IfVAuWw3pL/v5awiNjpJ
b1mwLOB6wQu/ex1tL4zKb47F11Y+xxOzMN21sKgewNHviVWW8KnsOdET3W07nmvI
Ty4Y4XwS5DxLzwBIcn/Hu+bQp78l3U3J4ODQo3iu9/Y0NLeVpYmhxGFn8rrWQ//j
PzyFmRZ/KOrxixKkP9perOktWjkHalqvTawro19HzvKZnPBIt30drxjHwoVqjVia
zqS3azH/yddRBVr7RqG93GsiYTRXfBua5sSUyPTbgxs=
`protect END_PROTECTED
