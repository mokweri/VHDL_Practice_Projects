`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
thTmiua3QXUAPUKK4x6RDMqndI8NBrQKC5NbkwmSTsbFB6ZA742H0SHZCu86SCxg
tCnjV2MXgSnPEVEc+/UhAu9+DAuswE7rizV0Nv8p8GPVXVJQZfZzTUF5+InJHbLi
LWrO/YP5d9iqWspuiLYvn8Nj5L0kQ7jrtlvf1y2QfWx4kAREnObshjWACk1IYKnx
DxD7OgeS9Fw56tH3Mut3eD3MCoMqLce06dAWwceMfe9GwwOyIabR5sb6W5QhmzqB
yoKCJUywEDbY7WzOUMuuhuHuKIDSZM1R/XkLSRjxQs9q7HcCYrPRFVmbZpoXkGuR
FOV+2NAH4VpLgVZmKd4XlLx1nnBl8Go3+TFACnpm296r7NsfbY6DJCyMX3m60Uqg
F27P+YDH0Hwp/abq0eSkX8gNmUXz1fIWl+yGBboGQovIWvctGZnpY0k1p9S637ur
+fr1V5H402lwOYvPHV70nI9OPPKnZKqfmNDDPm9IUG1pMF1dRh1iJKBukyZYbiuo
FeFVxS0LR48MxsDS1leyGxLai3aNDlWDrJ4ICNvhUi+uoYR+ssLfuJZp5KjsIub5
K4CBL+4FRIYuB+yMbJI+OCNRVrgxlP5/ztUyUQhzZdfplMVAWaE6ba2NHpgblFdI
ZBQgOOdhSRfBANhUscJBraX/Tv2IUCEQDuBg4HFrnMDdLyQeQfwLY0T5PhhIdqma
OctxNrV6ptG6yZQQVVVcLiGAF7I2ZDNAm3cJ0dUNN47b04f41YiM/o6PU0Lw02om
7LQdnezkwuWpmdcQqiffARa6q0MlDaC4SzexMQJKEMuLdWAU1GTMJ5d2QpeigMt6
c6DsV905wbKu0hgd7z2vlNs6ZwPDhxVDfN/OttKOMxt4YVjAMbknukKpJqhZIV72
DnrhTgA/BO7wUoCw94BtTkt8RlF4/51pW+akNZIdYvxVNimV2U9zXFQbWHN1oq3e
VFHEydkUs2KW5s10OmEmf49PMdyJCbGJjWTi0Igy3RTHQtkmK39/sKQ0U3V9UsWz
RGO7/EpSmOigy401hBBTWLwnFRvTrxLKkA6DWOK0w/QSA0dpVYDOH4llk9oL+PBR
tNyF6/6xDJ6omdqTmnBLw3HolPebAnyfginoZX4fp8Sz8OSAUfao9d2H4KijbGZm
wt/jvLzzjO0ihkZFcXzNIdNhmFB913HB4XOMd36CmOh/RpaHQOb4t8JeBqfsHhGJ
fIe2EV47w2+D1mem7xdlOxgELCrWvnZW63orlboU048Qsq4aCQbPkKNFqZpBM96q
A4MkUKD/MELmyJxWr67Y5ysFhotp7jAf8jP3ejYqPI9pCnKmQFU6ZF3uZYnvkYoz
N2Rh9No+nPhMH53THreYtiBwOSpHTqPcnknODfjms5VPhlI1QfgF7Llv4FV3Onob
+9Ubw1DwUCnTGgbCZf+0KYUm0bQtT/1RN92L+1K7zR2bVWxXnDNEaTVSm+yqtzeK
j5xh/dW+P90ZLIAfbaoE0Nxstujyp1RwNvF0KXEtMt3LZw9ncAT05spkAQjkIeVP
06rUv//coXuWJoO78b8H6AS/LJ15wo2KgEU1C5syors9wffbB7M9vXfo3R5s2ww0
xEPPv6CIL0T+Qye6h9WSqM0VIZnhK6wCJXozRxCKCSlgRisJQnjMPKw4+iWYMCdf
rusit//9/j4geKQDwBZX1jUnt6eyggc366NpmJ6wCKbLNC5a7QRLe8qgPzHJ9LhK
W6LfFWk2HBKhcoYhZz8qNG7pw2IUyP/f3JgGaBo73FcHCkibi2tbSekkBxlLWPOU
jxlZHXMAPXw9D4XppIS4Wd1Dp11PF0plbZVAIfESJ3SZDLRvOBUVilfj01z878vq
F/wpwrkRukiB5VeMjf0Xb8L8sFPLfeaNM/Bo1Rf3DMHKkQBOYvV0RR2bBSrKeT/r
Lk8tkydZQezxnEDWxh84oCZaZ4fUqjEwUkLjC1YMkuGO7jka1IYTBEXlY7zvkBf2
vdsv7QTCrlC9AmogD3j+a7zaYPcJDjXsiGGNuc0jDIgysZPmM49sba764eTTfEt8
QQh7f4tvNcAratC1uGn+yD4/SVpaWk5WLNER1rRIVTGvIKfC/AUSmi1IOFtceKLN
bdLSr8Mewi8NYi9dgf7WzuJWMUQeWIScAdchVx5sIVTEe/rGrriSFz3RKv2VNOCm
Xvxvly/8fD40xiXJx6c800ZC6W8pOlwakRZz5BcJREQy9kYv1SsCqyU/sex5EDTe
th2VYpjCxq6RhVCeoSqO+98Ybhs23ZJVVKNQOfsqHRuhVrWZslbSD9xva2sUTyWZ
z6KfBUMpK3Xr3f42eiBeXy+PDqURkU9rQiTjU3XlYtQwN5uatnKsvaweHI0ilLpQ
MMYIJAHBc9ZlaUCKpg33pY255cchRAgz1ej+I7a6I0CpnPl8CMQm0jtsiSspMa4+
ouUfbvZXalI8RMGqglZ91EPbcs/wBIevrnHtNpiuKVQWoqFlRWvltX1EinRgtzO9
Fu25h+dbW7fJ9Og5wN9ud8bFY4juCBIXi8kOebQ1MAMNbucMG3l5KA8B70qeQbbe
o6Wq2Rpa7te2JpzT+S/654hFi+6rRT+x6/8c2oX9umh2n07wVvlTAPF/of2yaRuj
1NDmpEU/OXw58XnD+HPuBvxc08Mt88bWkfY9TGphlSLwPEu4Kc80TGYiNMdkwz39
Cd5n6unD689nj/LybJDD5ak4fMks4fFOPrL2mdHKzIICRSF0cwyB0A3X+1eNnA4E
0WxlA8nleDI4o/gF33CWFG6lut16GtIEF3AmmZ8Mn2VbwawT+8ZPqYX7Dw9gqdOV
naLKlGtmCEPq19/aK7Xf7OdnZjEYZR8gKvdrwVVEp3mHX4sDiimrg99amrxq4rEr
nh3zrUg6kjXP8v5DFEHjg9LGJtpPCx9Rw515q3Leep1+yxjBmst4Re/lu0yAF0Hy
vQLLoxP373KMW3N7sfs55CW0YZtU1ZO+5uywltj231SDktN9T5CS6sdHyMAzuLZh
caG8H01SXfp4p/TWP2HUHBvDRLzgy6znfQO6ZtAQDe8DCgB/vQj5b2LV6i7E1TLX
5AW0ckebHcxJGYFWIUpKMlKd89FuaED+cmX6rCJl/9QVsjdNkgJ3NHU6O4acshTy
IkLYFZov6fPUC8oEqZXMv5+oX6skQLzyRJeSSMg6tHkc1pd5S0FBP/8w9ZnM8VV4
+2xyb2owuHTjn+2KNVNfrTZYhgOuHaUMHyD/gtLAf6Q8Yot9Quc1RWc6XFlAOvLC
daJ6SFziRGqXcEnaNucItml4X6HwySucwF+55FOl/TG7uk81plgsbiad5XbJDRo+
Z5p8vqicsVzjHnCHHHfWrUFt5HBl0hkXYGEudDk7h7eYDE6bIlC5xxLVTiIWpL6o
yJKsonkMB2N0G+GWPwytVhiY+zZgdhZM0m5PLC8h6RH6BHizkYDars+5OUlaK6Rw
vFXT+mpwQVrhdNWzzuLXwc21MUxm+4x41IFthX9ZHDtYk0KezM5L0QMxBPOOkAuH
JXVD9cTOJoc01pNif0/sf+kaUrpu7A+T2yoxCPGIC2qWQjIAS0sF5kO0JklJM+b6
ePJ7yLDVTSWly230h06I/qARhgjOpYVCj6/Lfr1zDZrpRd97epeL27ALQ2OTJ1O0
E+F6Cm4iyKIEFRTumQytewwkJMTW/P+l/8yNA+enogDWkLqKF+PE9V1mlaUlVf+i
z92k53/pPcp+f22L1YzH00TJ3zDqDudSMrWcbC7l2h+tpNoi84bC7cyUtjlTSQ/Q
bFvrzCdGnlyoAg/ej11cfTSSJHM1ifjdDtEtZOIVOzkvhjgSbaRloQoWcMXBzLRj
Q8NbEnxH5cRitbbORhMP0Z+j7M+8baE9xnrTpK4k8op3Za2HU7iCZ2QAGsluj+84
PyWd4Auog50DCQk6LcTZntysw5hi3o8wSa2HtfHKxOsDnVEvytMN+kBCt1WsbwFW
ugnNpCHdvFRHN/1xq7z+8d+i+Y8YNyUUUZoXSSSVhfWjb0gcywRjpWaxsyVKwVdO
pQoIEowxxx7gFaMYSCgV1B9vouaY7dGcPpO1i+07OobnGPDhbdqKIPAkH1i4+hCv
Vfci0qosDIFDX/V0I0ulVCBF1QnOmNZvspmOuebyeonpg6HjztJNFxqtL7wdG0d3
MjtO+xhTa4Dub1cYBL8aYsfTYltbRDhtBCCWx9l5qVmPUaAYXTiuvVERqf2eT5md
kX7Px5uuzRNJM5YENRxp/U/PZUAxzX42kURo3w+VTK0wjrtksLERnhP1kjlrNKge
Ez7AI4YqtADcQ3V5qnmHDrIhAF6AAWqH+TeTIw+v7bhmOw4bDNG+L6OHydvRnYDt
LNbOho/enVPzYqkMS+259l9uxJtzEL07uTLlIrsg9r/OxmIaJrGbB4hVAGbaZREi
9TqKUNPfTdCie2YyTEhMMJgmCiyUfwuKkAO7baiS+joBbuyLflt+KUskzB0GH5Li
RgF48enxID7SzYB83EKZTAy/W5YTZUUT7eIekBklqIAtpjppbdxn2hlqyM6O7ORt
sLi9OyNhCfSaDQZrhUNdLjYAWK8S+aAeL33qwkGTdA1AQF4uQsGJeuqOH4/hF0fu
jA4wC8VJqU9APJMrDPVtmVNODx4tlHl1gZ0+z0cYpjlmdNtrZrCgTffwV4OuXxYU
ZEkODoyM7B8lya8c0Dm+KCzOy5pnacFEZEEed9c70E1IXJXWcGaoOvlMZFxkQKrs
dp3uJWxUQGu7868xAFWAvPE3gtyouMLZikJKtriPCdS0054lt9EmJOHKbvVbJuV2
0DV1kCNPwOOmeCZ/ZigcMlA8uZbmvXIHqpMZ5hZZYGclKaiyTHz4a5WEDR/4KspT
KzfvpTtX4RapqYuY4VHrIIT925JIa8GP2WNnN08mPUtebcfkvv4TTWJKOx8HlXhj
mFiWVDw0Ls6CTrvJK/xvfMzLgBITdYcfL3XUB1gQLMaO7U4qQ0X7myIUxrSJhv67
JRJvGlIwyPx7QqNYTAbrjnkDPEy5z6RrPZ3e9gm7QxChwAUzHiSDbQ3Z41WHkTDq
ES+KzIktAsw/hoIIfke7Jur8ctD6An4EHc1RKgJxKMefV+WQcPJGx3DNAK9WtrXY
DGpS95Idm4v9hV2olHUIrTCbjqn+JkIsnZNOiTNojxZMCWTUwp3Frw7M908JhZhm
Q/Z548vvVsfyRKG3QncubgEDZIzT28fUO137OYz+iUVzIp7ZkRuDH2DhI0s8ZuMe
NOLKXWh2bXCEjpIbSOrLTxU/wO6TF7+oD/85vBijcYcNoVhfd+f9iTw/gLWCvRSd
AfaoP6HnQWzM5t/o8OLu5LboBpbjRDLhbln85fxQlN/VxjAXvT2IRpP5eD+u0gaE
D97pRzf1S5nNtyCtTyT0uqsWbmTfW9QZ4Z40d72Zob/teR/9JDG+qkACpHLhNTzo
9iwmPTq2EgsxA2LAAwV6RXslhTmuUEvRIbDYHRmJeFRSswG8PC9FgG7PvEp0fjQj
1hrHgZCNBPMOGo4ZYs8trL+jtNtCzENbAD2Uyed8ejblKdwoX/xGZz/xAxmbMcZR
7vcgLfu03s8JNQ+xeAY2BBtjtQj6/A4MOsetcUai/GMTmAketDXPMqpVnYuroIRU
jlaXGOabX5+TCrMYbkO7DJsXEFMOSeAIAzGUSjoaZyJF2Tpg/BEV5rHh7UUFNWfV
AInY6p4OQ6ol5f6g8WCg/LjmRA5UH/72YKACkRit07/7Qr+rKhqjAN6vw2zhAvHY
6AP8F2+98SstvSdzkFS00MmrrKIk2t+q92O1eCTa73VzD48AZX2KLIwwvUgou3TR
cR+FWZMAifWizMZoI8rPjMzJ8r+T5ovR7soR0xsImtFWUyKFwjhkMNm0DGZRJC49
a574kG8bP3EcIzuKhk9Xn2+fO3byQ7sDmNEqwEiPvYm9u7PkdfYxcDMlwyQjGHhU
4qLC787bsuQF9lVlIaDfdgWSpKGweVfE7F7KgoM4G+CpR6DTK93HTqInVYwb3up0
Dx44btYO9YXoHwO2LvqsQdwHCHKLFXFJ8VskYoVgIdftxGFuXQWZrI/l2aKJryIO
yE1Xd/5CI0HRBgPTL61BYuEtojwoKrEun12VTQ+78XZTdzbvwIJgTMCo2IZtToE7
NtHYb40E8521YRH+7T5H3KSYx2vW88aGtBRqKwNUJa55TPlAJXR4TqNzfGBR9HFZ
30UyIIdW5XCFbInIv9TilqX3XiOjgvBQldLpPaTa9e5NE88eWsTE6kIVL0JjVZfK
aRfqkaOW75odtjOrJaA5ITYfcUzVw2uTZyyJ4UFMgLXZ2finmvTP4s/dkRHk07dZ
f2A8vhY6MrKUix4n+tK16kNDpyM9t+0s5yHEs6nL8pa55InlRYuwSGyrzapZtJ0q
gUHEMmBfCqlupKTtvUlOPn3Ul/lRF2penA579BO1y3hXhYBrOUY2vJo5ztFKL85p
fFoESeukkwGDMUD1fMrXhLGD/YENeQRiD3VMGUyWP4PT00iXbANHcT9geJTkHboh
Gi/1GHrlQsTKwU8T0NrQWgYmmquyBdrfKObhr0fl9QOO+t9N/XMu+TIiMfbjgDRZ
788kFyA6wnTVr4CVNA4Z4h6PvIav8oWuArgHJ+wuu6Gv6fOEI+7LUFjE8HMEGKH1
4ZodO6ccCxiwKIgOP+ztIDrmAGszwi9HyOXPP6H+QyE0CKlGX+evknP+EMC7FFeE
ljED3h8Jxmdbc19mrfUHVhK6mRMbd4MRVApyb3apMK1jI0d0OcOYdwq/tYzh91W6
Pt5pgw86oLQenwlAaRiahK5vy7xP6refSjWJ281GQohav5pBXWRvZDs/+DQrJg3w
ltxqqNJWOS26A74ad3H4SiZhL6xfC3oJtvqbJ6CYtcLrCqU+yDAtGjdauJX1xqYT
a2Mivj5Cwu/9O3pkP3JBO8k7qv4KsBNSAaKlT/YjMhSSQFmaUePF3FLvbEd9cJfg
i3mHYuCzhwGyZuRsh3fT6P9noOnCfHn2KjlwbCPSiA7xQ+lDQU0Wpur9Mkd7ypVr
uBRjmSpv8WM5VewVlCAPD7QVx95M9DjNOGJc11xO4wNscrSaBhatr8ZnpOKhKII7
rfBO2na2g9py6EF/koQF5JZeq2bRW6G647M9IMgPQGJDoKDA/x/DVVuFu1JYylkJ
dkFqFBBrjvEHIgmj3NahDfiS07nLY7FtoGxskXkSRTlPPP5c9spGXTHgQ/gWDiSV
geUzuZHtcdVxF/SC4faN8c+8u9gKiCapg4mKmzkcdNcy2AnDFDNXQrmzEgezWL46
RQcazgwHL1R7YI2aq3afPdIKjhYCqQBqT+gRa0JE0Ibe6tUrs2gx/t+0NnZOQEa2
FCAgbYMaIdLR3ZAm6rrKzAGGhT56XGo67lqV0FXJw1fbSBg9pQRoKNqcBglsAQiS
7SAsDAFKYCg/BCtAA0r+2JeFSVddToWU0qM+x4Ow64vaqnMfvR3KN5oKTebuSFuC
SrtVVGi1fu00gg3U0XM4SwnG3TGA+cegcv7cFsEIvN/NarHSal6ZD2lolfPrnHRs
FWA1oYlomNCTpyH1yf33AbUNvldfmjP18N/pSvanGXgojwxOOtWBCDCvnva0keUC
ZCildGA4zkMOhF84HQEcrMfy5ZiaAGwbTL0O1g527ZGjVHOiZtsd33nA/KsIkDIS
HWu/pso61zj4KmxCQkK2Ikr3PN2C0/6HynFauz3kfydPsV+srs8Sa6MC4BcLjXKS
cUP1XCnfp2sDUepLcMxkaObsMX9GaijhgUkWB+QWoF52dP2PSeXpYZ0itF9M6XWL
Y1s+cOY7ExQg/6ZyDkHvVhGHaMWtVTKqM3AgyEBN9HD8gN/lGKUqH6ipNrTFXF00
ewrnN9K4hXT73oIBg9qMvRc9FsR7Y1yMgRZXF3CcFq0JpkTlpNUy+eLhecwp3gdx
OI/PO48T9mJVs7dSOjfZ8KV6g8iIHfaYCRyvYTFs5E6JoqgfyeyC7Rs0fSe9CuZO
4D3w17wGg6baVM7cXEh+BS9Vfc2X5k0v9RR0zlp0ZkhgumeRHnm0qF4AFYBz3zCJ
CRY0vN33R9+LKZ13bCkWLwkOC1cyA0UzE7H05ts3UMKUZhuh7AjjXf4g/Ok3DEOS
IIlfkgDoj3akaY2dt9Ue3iUDZ0QW4fGCO1QiovoRPHd/zS0XmNB2/t89Buvw1Ygp
Qs/0lX9OyPVnhlETOYGUvOGIXMe6IAiKPMhoQNsGpmvM4suVLQEcDdyWTy7kjFtB
jvwkgpMZSNNVaTf6E5ArKmzeDNwv0x6qSXnvsTctPK5L3z5ER1MwvsSe1kacyCWX
cbVF+5Et/OaNvkZiT/d3jor6LvksCUSW/hGZs9e0aSDaj9swan9IfEPFFGbYy5NA
MB7nnuuiAUoXTdWctiZZ3ClwwSpxO5kCUE3kxK4Ay0cpO+u7z+GnPOpaen0cI6TP
flLa/4so3nhzC94WDJQbUkJyqsTh/nL7/gkkDPACRRn3DoulrpPQ4KvHY7Lb+iri
TCCMt7GGTw9QNuxMqT5Uy9CtrSmlzg+3xXWHdT59wxQZIFnTJTwb/5yr5G0VVLyf
nS7er3nwoGwoyhz76yHufw==
`protect END_PROTECTED
