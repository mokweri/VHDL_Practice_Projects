`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+p90tXXEoDesq1L57X3gFoefHNDc4qA198uEUJ9u531JOabjnMz/xyqXU13eeojB
PbFhDWX1X6IuTOj322t5eogzJw58JBuG0fbv2tuHqCPrVTenIkvZUbLlS3X1r0Oh
gOWrR8FrTp5GKqSSB3K0J7E++AXq/vt+Mvplr/IMhzvbezKFJcOlJj9VUOWr2dTJ
I0U563HGRC46qtxNnulf+S9i6zq/Ibh7eK90LtucXzVtpK0BjELfKa8vZ0Y3lDM+
x6avYBHZSJ+GN8ifSRaTovb8VHCh3/gC+0h4Q/mO0qcIrpx5baPbZ+VeDrqMZJLK
tBrFRauF5/buKmx5btgnCz+0sHP34jPmFwQLxwem60ui+fVYruHBuP9PKv/xIIik
AJw5pudvMHgDT79qbGdn1QKlQGkaorNUCpA21BMCjchor2JUNYS+BtNK+CAFwlD1
0m6qdVucmj6vloWjfoYYynVfz/HpSb6md98jvmhDt2w24KeG0TecR/6/Gvft7XnS
AqxHHxxDVahCcMsRDq3taAnrt1IqSeXarp2/zMofgC92dPu5yRJS4h44XjTGGPVj
F2exbWZnr/0RDc+9TwMeHQ==
`protect END_PROTECTED
