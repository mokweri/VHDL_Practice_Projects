`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+LiKn8GOYF63yh+qLg7vcVI7ColWm3Uhpqo75FudIyZrXdG1C+iffPDsKN/gjoHC
eF6+PkyY702nwIJlrv9NwyQq+wkEauqMGOep55sR5raLgWsHM84SBSIrVt1qb/BL
bu65sJ7LMGdi9/oQPWZUm91PLU3GrFKXLSEYIZwXxQAeZeBfVFzEOzrDYQ+86Cnx
s0H+kb/RQtQ2O54F5L8sGM/8YbRRS4g/Hp/Vpjua/bFlQgwQCBMz5MH4qZwTyCLr
gEDbvcjzptoUPs2IN2imbW7MAkCUI8Pp5PLoDgIClO2xDRfmn8fDwEh05YaRkFXF
SNoxmSQloDARVtuilwolMHyD90D02qXCAi9XaXGXeFzk9EvFofbVnqw+h1eDVJl0
WS4sLeWIWTZ4i2RXTtqIa23W3NTaFvLlqRGPtZ4kSXKy7+LuVQWwywoiDcNGhR3S
tQg0KmLqx1NfpcFTXkby5TJ1B42ob3oqZ4jGasvAAPsVZtgyuO7pGsE6hVUSAY8Q
zus81cmXXB7+kQ/SgCAaEUYnfpQuQDSuKmzfytXHTwtG3MIZRs+U8N15J9AQ7L0H
uXJON2RcS6iSaiuqHOHzN61y+lXSeoWax1ma4j8ByRwr3dLP+Ab11WcTBtexCxmE
I4KL3mAYuGDET3w3TZO9+nt/OYkLzrfZu5J4X0NSnlhG/YfUhHjloEtxjQ3jHnc5
vpKoY5IqOHQzgxJqmXkLhoWprNZjPZ5FlCUCckB8yTsVcabp7gzwbjnAxZA+KwRX
a1laIEL5TszQyJgJX0+OHF5Uu6I46tTKDT+zdUzGgtiDXwJSfseVOIAaGNNGlRor
uC/zbOhoAn5obHOMqqCIdSZvNCNhfjLaBuEzMCpXL1pfIRdpITeRfLovq38gxHR9
DdBD4dfpyS8DY8d4V5XfOqe0kqvYb3gk65zKOSsQEpcCRqsGCCc5vXXX1SJuGjWW
gFB0BDqkE4/HT5c7oLr2t6ydqgncKQY4+l3wuuJU78za8UUYzvvmeGnGdYGXKYRx
m0k+SmQETQpH7pjnCXHedRsEqcn3zDXsYyZ708qlorvxp306WaTWhmZpSbYGq5BP
V7zg4+7HcF/Xu0LynFR7tJ65lToM+2iyv7rhxhtkjdNVv1n2saWMJhMmH4AXOfM6
/9A9i7PviZdMuy6t+LW1nFG0zphHFlrY6cHkGJukdPbbsmCzD7waLYW7szg3ejpn
i8EzbfdSczhtjhIIrk8swb5NmXMk6Xvy1J68u2gfxwXW3juwixunCmpg9WNlRUqu
DskyP9IYiJuLt8hpAcIYnju+Wtro1Fq7h0Qe0tjV7LjP5QWzjhamtlDhLTgOGj2s
XyzERIO9woXfLtGf5hf5OIns/68ret766M6IrUFqlqHQSPYYBL7GOA1Znf9MiQzQ
uz3jmDBCdAuusxmvZsy3e3049OVAHD2RR5+lCTLbEvoeW+CkvwtjD65zutclKHO5
DnEJGa44nzCmaMSTa+1ZYfLXsLuo/EOklGsZ89BZtQggf4TEQBlaGjveZSYeaOY7
PwLgy0Cy/TVY0p1l5eAtNDxM91hMUlk7GfuD3l1ffFIxhWwYoG0fnLemxoW27Hao
QWCjSZAFNNj09wsTK6kIB7J7f1SkARBOlER+BwHFMvrhuwo9kbfM+nUVmgkP628a
yDaDbisI8TbxZI7wAb/TdB6CsqbSF9OTrCDayDqwcleYd07aZjqkuie8JvT4Lb0e
fuyNqN9QpCPdBQjHD6KML0wyt0oS/I0P2C2r1MgxKouWO5mEPmpq9rmnwm8coozv
Mpy8orzJpXpT0kYx0DVIrP5aTFR8oK5LsjB5Ehp/M05cysaMCSoX7JREwUsH8wKt
dckeXPujpc2pz3fZrDQgrw4wXFwzQ1Mtcf5EPQ6WvXyWC7MjFt3Wz/ezpiE49oPh
fchWPWZP0dQI4lzKTxCX4EimbN+7ae8nkiL8vme9SxRDJJxEiNy206i3F5jXl4w3
mDb/d9j28o5Nq2WYQtidXSVBvdGf9faFxNJEzKBbWKK4x4jHUTShwHcHw7LvBmWZ
fYY7A2+RsdkfyX/3zFMi5XCRVTOmmPHabNNmF892hjEJj30pDQVJUFnVfcM6XAk7
8od7po9zODSZp4pAfWXJsY9v9k95Q6b3A6/1CgZytSR0SgSWXYKJwOE73cUXT0gb
UlMZpN07eWQXiLe6ALDP9HrCEg5mL+mug9rTi4ptXE4WcneSe37VVA7K6gXs7Bz2
Af4DZIZbDq1Ufp9I/QLfN4coKj+SoD7RVlT6uCD2ZVEvlUM21KCaoUdXoJByh4Wv
7oLdS4OBS2GjQ+vXPJYeVjs+b1QWuq1i6WJBtv26bOsq44wXH91BMGw0Qgy00+G7
0aallUxB944oibVg+47Y/64sf1zf6p+IH6ZVYF4wc+NPf4JNCRqnzINkcHdnXOnF
k2TW+PcjtRDFtfAJ2B6LcCh+mpjK42JY+eHLS4LaNR32Xji++K5dK8JP3bpwOQXY
5fRNXwOvA2u2HX3ObgErh4nwjvusW2sOuxsZVrK3WjdHKPYoNAuT24jEAYy3bhST
E+1v8QZtUlBk9XIhHRqONPEmkcCLchDwLaRoooHZhfJuM5kIN/aw19BzqgQ/qhMF
8EWsQHeB3LNXUQXYPQGP6MtkgUBJO3CWgjcDldpVxyba0pWz4+Rz5TntJVTdZAhV
Hka/8swH395dll9HluEqx5AJXSI14EZjrhEzzQiEFQdpJ5uKlL9QiEZVctfOR0Vv
X0oIKz3FUs7ZygSCoI5dQUxLdOwKHyB6J9LNEsdtGJlSBI04IJehJX/OPOc7urhT
oEpA5nxi8FXR4V8226zcB0c6Za3VatlmVuQ8pGCrqOhlqKHx/IGQkHdmusrs7CGG
wEpfzI3sXrVg7pgjzxokZ+6/Ofml1EZTusyB8XysEG9WYUobUMxn6wgrNbDxy9FS
y0zsMNqBy+A2BsL7djX9I4nt+ORpaaXj4sn8fcDnpSpdPdHkYTsplroTnIny67mI
uwm6uoj9yd2x9r2CX4h249eObm+PR3DIgPMsKX1Bdpe7heJgoeCZzP8XKL9W9wY9
RYC1Cvnn7m7Ko1760G4hWVGiKrniPfv7qygqgIkU59duq5ay78+8XMBALIJOBCTp
Zd+aTjNveiV/K5wzNbs2/jBnamqFPVEVEubAPfT/tmLUE+Q9ZB7MJug6+7knydsv
xp6wo8RsOzl1tK2urLIXf24XkHbo0BZjF9FRGQjGhCYAxUVtvKwFwdFpnJeHbynV
2kF/IC6wE2J3X6wBq7Mhhr2vbPtQTX7WTflIjsekreU8vzJEFY1Sy17uPQUhpjkm
WhXCJSIy0yyK/dp1fVEU1h2MlIpM/4l8aw0SgOjcYXKRBHBLlKMSzBNlxLZ95kKe
4O2vKGF/rQGLVox0X6ptaN+/1P/AwF4SGoVD5f6UFcDtRbwA27Eq0Ig+06ygKZtP
cB2s2F0eVkd70jy7aNb3HqfzKkNZMfelDVpiIjCQA1UQS6jrFjNDKNcTeEqgPW6M
C3LPWmpZK7UgMXomedV1jiaCA3ufVrmV+AKYza/8hSb5J483CWr1VbQW207af92J
31QRPciFodtTGR0/cyBky97KE6vQJaNiVQ4Dk57BxeDP6BzEuZalJkF0PLx3qk+f
L6gibrPZDquaW+BSSELvihnS1JQ71cRoHCwcJlMTQ32SdLQdDllvlJZaxeOnkNdl
JJg8HK323QGquU7DAFudKJs/elTQpRRzBuBZtt0iVts6fkhMDld69e4FKq9h3d7J
tsgL2LZ+k3doeWvjC+ab70wH+i3aZRhB2pBp3f9f8iET/n9tnlPg0n7kflgW3XKd
GoCwB20Hanm3449bFPShEyHWMSDroiNJwznXIafMbhWnw4eu1yPx8/Ek7lDApxpQ
PgWdxTAaPIiZZYsFRCMXh40hbWYCJ+Qif3SjZnb85SloVhlQQ8jUZ2a3AwkSdo+r
moPecYxbNRWdrIDRU+WiG+zxAAyvY8CvqUmCu480MX9frYCGcn+wJ+F+19Eu7b2Z
BpiqWNKrVckmSsiWYhaMGJS+2OYUjXdH2QA6PgkI6UhmXntjwJmoeEm3uUHimFbQ
b6deHF1yjpk6x7NbLb7bZl20g4Tq0f0IkNEI0kdyGR6pnMzvcFHv42Uy/O2Z1wY/
d6ubFmqyt5xj1MzwRd1CROwCu8hxEFvgQyixy2ee5MV5NarXEatrrvUZEc8MnpqX
2vq1heN4rssWOXv0Qv0stbAYoVcb7uYdLiA9n1hklnoNeLbw9E0Kt5AbvbkH5ZV3
YIUqGw5lGpzq708uq/6ZaOTij7wnEcX7NDjB/7ePxsOwJ0RVpbn4mZWW8BcxRxjo
7jd2LudQg4FfxkaZxapT/TwXwqq/Ki0qmgJWv5VwE9ogBs2CxLeM9kDw7HoFjAMu
OBBlR5s0ziUGdNnPDx+upT9P3mC/x3JoBWEIgEVSMwFs40Pc3ZGnVCyzF5QZGGR1
XDXdu/QIFsjveoTOq6KCXdTIVpdA7+W1FUkM4OQ9KRyi0Nr7W0F9fZZrSdsnks/u
t2MbWyVWYyfuO+toPykdKZE1VVLr09eUIXKdwom+OKUEOBeydggePCOe3Gbs418Y
KR1L7UwrNycFNlahy2xqz5REBZjMsG1GDgrjM3bYyTChm+uslM2frUBByFA/AYn8
7igWgaFTmgXa8J+OgMTiFinDYjDVmUYkpj5GlcvKXrB/TqWYm7zJu4F0b1I6Tt1K
iWkocxBSqRgG+IOVU84qloa7Q4UPhgEGFaw00BT1Jw+p0fzeYj44e65NblXGJYp4
cRF5z5qkU7tSFrlFADviwiI9MWNv/zaPtKaYSjxY6t+tpWqhnBlOEvjEF1WcHvAa
6NUXEZ4vLOZMrhX7cks07z09Ywhqdg9SrK5NOX3xYnoK3V+xg3J9TCV8vosdBIsd
VX0pKGg7bo/CzzHomWdGJw5k4YhYVF2Lp6eXlIpjxA+u69mSd+agyRKaQEzfjihp
8S7GeYURHp0YGBAZIVEHJvivCnarfRF02uuIv89/qngfDxJe2rdjwxtN+VWBBc6q
r0Z6uIKX4sxkap1JTG1wi5SAp1PC5xOlP3MDlue2d4tCFvViL6jYsgAO1EVkIXP6
KgThIFepJVkAwliB9Gha+4HdldyDwgsiDlK9ypG5nOfaI5+6L81z6zyGhRN3Yc7/
QOqXr7EXlGpXyOhRtKHqhpEiXS5wC3YgvwVxgNR4wKFimHBMcOIHZxdC4xT6EwtJ
6by/0q1ZTlpC+p7DWM5+HcCbPvuEq75UAncSE5+2dywtD65FhV5t/vLi8bh3BDG7
LGFnZI7tuOaJ7Ui6eUs5dsE5vKnNomuS93OC380hzuZXgjyZvrR/fIyLvHcriuUY
5AG3u4qHi9BB/gw+sXb5G3L3aM2d+wOybEHJnCoJ0jN2FdnjCx66qkV8PVVUJ3lM
dCo4SZxbONDD5LXPubTu/6CD9/AEflYonVNl5Bu9izLnhCV6vVevZJsvVaMTglmG
nSzPKXiuiIYOv/WYcCD488w75UxcnLSjpVMZPMeVLTiOrRJb9UspmbZbcythT2jx
uEEedItToKKDAhxwbpVL2Q4o/BHM4GIUjDRILSjDp8K+xX+fisis5Ns9ifmJceKJ
lJXe5RcSGsESkIsDiAdVf4weA+uWF94bttRAiD11Z4L0A+g/6E0f6g+O+Pk1trVY
5poNSK8s1NmPfkWoasbYdrRnWYO72qX89sA9qvOuZgCS0aMYWwyYn524OdBKG+mW
GDNgcVQmk250VWwfxMpcXBI3dNT85lbOhgq0fc4xmEVj1idht5lUFqO4zBtovNdk
vznSw54xNxMfCYGyOrB0i6z/TmOvInVeADKa3ZplE6U3FVsyW4yt18ChR1jO3iGk
TzEvxyoaG3kaZW6xuXX5XTAA9ThvXdNoXal/3CR51YsELzw9Jm1Pi1moZ24+Af2p
tc7ObX1Ya+YaHYybc2oBLZW8anVe8E7ozWcW8QgoGcK5pJUg4Pq/kgEa6j4hqNj2
69oNbo16VFc6Umsq9am9tHGdT8MsIo7boUgHBO1eYeC6Dw8+4dorIqwXGguhMkK/
HX/0PAXWq1oTx2g9uBFoOCTzAMRkunp/AfkNl5H+JWD02lkpWE+7MD+5HH63uraF
r0meqj2jJ7Iy08CqPkcLsvp0cbHYBl11yipgpYODATDa1Ozp3geuJCGDTHdISWBC
KL4K9Mx60d0I5duOtyhspmUjs1aF68I/84XT+FPPcqahRQ/iBP99+dyIDbtp+0VT
+nW2+Id6ycZViUGwE0kqrXAR6uJQM2b75uxymS4F7NbcLiOYmUBu0FghP50gYeiE
FnFUSqm5TxVkx60gDvuHbbgGljr/86syUEjoKe9NlVM0QUspAgehqCBScZYqNlq7
EzOd1oqmsg/4PriM5N2gFtDl5WWAs54JRDOH1T3r99f5o31YjlnUrGpxIdombFEp
kwoNUGsEt2Itvk3BT8bRmNw161h0Ley9rMlRa/skaVFfEq6PgL6ByIsOq0KmdMjT
imPxAfA7c/dtvzlCt4wE1T4fpR35as5KpW/NlDWYkI4512JBGRySPCAEQkxadZyv
OIGpXvV2JaWpzSEedjnJEpBxlYdKSHOPVhxbg+MMeLVkg3qQv85n0b/A7NXJH4LP
bIkchWNULvRXCRXPlv6lWGWLVLQiE/i12H03dhKPfsqTrqliq2/DjjYg55CMw7JV
ADrY/dg1FeOQd9ydfmKS5Z1qOIkfv3R9oV/ozJpEBB9rKmgDND4RBpFKDMH1s4OS
TwP/IFbuANLhk0FFnG87z+1UNvW4rBsO0RZB79GMVjzmcF4gYuIKdg7MhsB25KEi
Ucp3xudymYZPrIYHPnAsNwKnxL4CrwZGvAd1dq3Msc7rrUAuc7KRK1ntgciZd7Py
ZT5u0y3ZwTwMO6aCKs9iztVmsdhlQpGIGz4pac8DbBauNMGMc75FZvN58uYw2/sr
MuB0iQfvWwfh1Q4KmB6vmE7Rl8f0nfT/o3XcQR7vpcQzO8g9Ag7JkZWuh8H3FRBO
sktzuFIXMwbROLljfGiTsb3MK3Cd4KVJDe2m+pzot0YjNbEnQKYeVjRLaeTwEYRP
OCPeSmWI26IyPG65EFHqbf1WZWDmnsjZCiC0nDY7wbHigHboomzyTy/BER53qTf4
vq34l6VMQY8KEpAg5iMWzfT+HEooiubInUTKVv3ciZKtKW5Rx5ufecCBBcKNLInT
VUFnVlAGXb8OYisPbCOiYeZgOhM6Ryep9uy/93zHSdNYf53/oY8wawfZL038VLly
lsxaboMsg1QFZXwEcpMQo0UU+QKnjvAKNwboMIwVt5eLgjZSS+dSD6SPlYG1Jvrf
VlXev+mtT6Id8tYJYFJ37ZY0AynnAa1mrgz4goZrEMELRwgXWrERBDw65bFC6SW6
JNqwswlg1HZ3KTG9nErrJSvdYnxsqXZHerLVKVjXlvdQ9u2R6RpnJoPCgNFMSrNz
RylAcywzJgctiBvEr7yYx6/9S9fO8QP1zc8wEKeWsV1Uat4wDdRjeBOSpeFmrUem
r9hxjJFS7iO3UGSQgQX8hAuzfIWTVSQCFdCFWmiqIZFPkrderhXxJNMNkEC7W6BF
BRchrEcSa1kBUhH6tU67k/pRG6nH8pEqEc2de4a+8vWJJC7rCO//GaexCmlYfRmx
4KI2ewDYM465VrhDwWyb9rpJBDgdGOYNyeACzcpVYW+IWPw+I8dEC0BFMPrls2yC
MMTdQcgqzDm3lGhrxq4/Ri1no6kEy+9Ox5KqIBFO+76wAEtjo3iD8vYUsHoqBkwS
BWKU5sko78ACLa7LM2wL1//QisSie6Ic/LDiRltqFJNJwH8iFmZFdsJtMXwynInK
fL2xiGqKrp/6HnRXfL7WFG9/QnNbOhTF4mwFrnuAT+oNVU8gHPvAswEbB7V2hWSX
OJbbHpdLhwBaqRrXMe6jUJtWTyPa9+GWp6Fh69+FRpnLqco3WxtkAtnXiVydedA+
uRpe3IFuZcW9tQ5l8/opr05xZMoA3udXEYE2hsRPmeeDk9Psmj7YSQ15UNhVL8o7
DiTuPiRfLkuuwBUyoTS0Et167HYthGz8QiMkAGH4/Ync8WpeOvQb4ycBB/Wodq0u
ipvpDG62e//MUxNvm0SzTmoH6Mz30W/QIIV/56FkwnAx/5tqNVbX0Y2wheWFzV+M
dG6iMnoxuHsScZ9U4zMB2Bmeh7YvGLojOxIBWV1wRRw9OfEnsqvStpZFdZENFlQ4
X549xJaxjr83KpWQyWmXZHFFr7AZ0/VxOG1IKXSbWM7P842DE2iCwZPYI7Vu7cAO
pDCp5SXBFSLv4amsbbzzcPa14Vz2toYpYvT1tAWnRppQkuMZnCMlrJCf7pGQP9pY
bnpT8SUZhQxOtHcMp0Um8w3YCscls8512/YFU1vd/R1lgS19yOKxJsJlrAKKPOmx
KiHMWQgVyOhYlFFS6teujFHKeGTJVRc+6M3mwtrsEE7cfCdmHOyk9WLu3ztolo9R
lvk17fYi5Ng2HNsebnevMxYtQxSIUbTsJuGRdBHP0hJZCkA26N1gr0x3sqCVo7Py
/gFYzDwPXhbulsy50J3d/g==
`protect END_PROTECTED
