`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5bkn4lLqEigx0kLG/nwOU50y29hlnhBjRIfruOgQv4Z5Emk4xg0Lb/5h9vPNtj0
gWZDsjitVWE7nf/z6lyOwjfyOA4cf8beHKR3iVd1+x6qvZB8KHRRdhGCV/6qywaA
zFB3D+VH5pSBy/cA22ONofxD0gcbqWpX7lt1+jJ0/FyaNDSVG+X0ekQZVViRJclf
0FXQSvROOPqitcmkCMv2meGD5AMLD5qNGpP3yU+SsXf/Bib8lZuAYSA5SsgCSfqW
UqL5SO32pNqUZDju5poey1uh5qhjqUxc7Ocos0ttoxcwXRJAMLKmpeVqkgqHq46y
D9etBl9YyDqsnXYKyJfDBuduJYduzESNouNQRHNc1PshpKE1D53HbaNVrHY99Mcb
k+CKNSxtBbB5ujTY+d5iBWcE9FntTqNhux+82Ew8RD109iPCKTcQuZRjiqNd1K/G
RrtvDTcqrNu6lO5NdJFrmVal23CJ/UpXZ/4NZjJDjWGAyzUw8RI/u7QsYNUG9sE5
B7KqSthyeDZPD7rxaGOVYAnKS7E8UMggRl0Aff9y5mz0iHg0xniHcbGfniSw2cGz
YXQEbfYfjRGb6cPxLgV6jpg2X/I3Jbv+xQxrC2kBzCBHz0cDLE8r9gyr613MrZ4B
BvHoHlj41ECl4//NWnNukP2WX9EGT16m8N6u8WsGDzaV6GeRt2rqqgxL/Z64MzEz
jhnbdwudp6GR/TsQpxlP9eRKYnssGOzrLAdKrtGKyKngo78/fM0L5eFy5Js3o2XF
TEac0MdI3Ur9oWjltbZQA/lpth/e+zLopTreOA4PMl5m3Iq1HD45A32lLcpYWV4n
fHjPfG2HQU6xMdZxdqTTG4rTmTirQLsvImgrYIiAM+OE377q+k8H73ZfKBfVmAdx
uEpOs0edpYq1+AYD1R3uHiQ1rxzxNB7avauSyE7lS0GUs5V5syU0HmkO3J0D7zWT
eaVjs8paKvzWuDTdmYpW80InSiUrE/5bs4y/nq+HK7decU9zCh+iNEkS6ftD2tXx
iEgoPOeaGWyuQhQuJSu7uJMjM6ekSUeIARJwbAwpRk3FHW4loXBDYusOLW3lbVia
ilQtJBdPirmF3kVclO4B0F2BtdpR8FW8hg4B40N6sifu1B0MaLvlXujVInPds1s2
VdKzuvahkchUDFm/O4NnEXV6kqindymI2d8/oTbtHYYFLDATDEJE1HL+pQgj+Csq
W6EZ3GfV0Sawz+JNqmcuZE/er15ZaMueYGU7G0n1WpbPwwwlGn5KYjO5i5GiU+n/
bHj5n/yctMByTCHxDK9vNRrPKm9ccGSrttXh0qeSJZ2hofM8dyT6Yd/3eO1tQSyK
qeY0KcHais4uPxQUsBPxj5PjRwmAYsOyMm7Q75WUJ/hn1GlFDoW94/4dLO84uV04
JViHNS+HTA5tl2pNmu1DWEjh+Dsr0xa0PqKHlLY5A4DpkrLpxDIKFaznCX5dMSOX
wmQ++nUOATps4NSgKpuY2/VJ1r01N7WZ4eA3pTzE607mQu6vSVCScRqP5PLRJV/n
g4hxVoEWEyKwPPqLBmfeWP9Y5f3i6SP/N5Am3ZbUhZTnZWKgRhfoElCqDm5vdTb8
p3yRv6Jg1fyvxbLG5WjTwGHAGi+30bLO+wgbiZZk3cSjCjJ6g1HK8UM0TdqoENyw
gttSkfsxdLLgLhtrtOeFRHhbDKX3p6S4gzPEcI48rSDqmJTeflb5MyQ9ztoscX4z
/EMd9q7+1CBhYU8rLQUUyhkhvD4dbkXQw6VG8EzDdV+pSBe7/jNA8FRYDlYrn6PU
v+r3YuJGt06dQGzrHKtlNfLor2pAtwDBToDdoOM+kuFrSSsxb0MUw2NJ8cni9uyN
NA4ujQIIoxyWPY/W756rbzrQMpDsNnDaxu2aFaZnFfyQ0ByU3ogtA3mQxqoi3Ocn
HBiklPEb55AiZYAVO2ubRjujLqfedmpunfX4VIbxQFk/yf9iKnfrHutscdWY1TgN
g5qGc/U3VNHD4R1GUy/4Tfmtbc7Or0KMgatqgkmQ89V9yuW6kilFWxfd5DRkJh6v
6uZA3Wwbcl2LzI/t3RDab76FzhI8wjpXQ5rQZ5brOGsXc/ALuwKLqRpAX98Zl+mk
11cl0gANjAn2vC47WtLeATwTZwKaTucCSn3BtwDJuyFvyZhYBsJPwondtzYbDefG
1qKAJWkgfXE2a6sgmmzSrbEWu0bTFFIms2Lrxn79gQUa901EiM0UuUWJLyoul7y9
zX0yRh4kCQkCdOTOG2lmvDxVBD36nERxNFNKZNC6AoZ4n8+fcwA1QVyj70kADsRF
ZHLmAX06OIX4DPwrBkLRuNOBkj43a/PvjAAULejfIJcb+hKABpjXj0RLHa5xjnYL
T6wREPfQML1WPfe9Q6q6mi+G1A/i8d5N6n+UCv7Bn0xLuTUOZ8IDEXhl9YSVVksI
eyXn415VdUkRThVoVdnZV/3TaUsMBCWePx6YX+6vJ/lHGcenW4WMLSMnzYR3yOme
L4pUC63WcsP7P+tl6RHy7XJEfVRvWkYi6NzvZ7KRGnuzKb9USKjo1iW2KL/+Fn12
ykVIcKA4XlT8dUtq2q2S3iTHBrhT0LoC67p41ajDy5jOplotabVV30hCClOPEVG2
+tbqlMPnjA6ZjpmR7w+HYZJuICWutAvdGeTgUfWZ+e2yMJ9GND+M0A8od8m4sgdS
roNxdMEH0eJXlg9L0l2d1dvIRR6tyZM85i49HTKNKPQUtiWiJnGWtcYy011j2Kgj
2HOch9GyLzkHYlRynGp1l0PntPzgArs541bk2yFGwhOjvvmRpVR9ZCXgJzn9u7mj
vZo5/OoRzY/l9euBCsWbBwmIHkII8b36csvSMZMJALnFehEmKUZld/TAjN2sywI4
CEmYLKcCu+94e9Kfa++tR886AMp2qu1MRwYTjjCSNlHumR9q5bHEIGgMWHZg4mLM
7CZDDf9mqfKhOt/ug3V1F5z2W8QtmifTqHKN14Y2joYZyRjPE6FKXHvYaC8Z4qXD
tfc1vIVcX+sLxPeSYM8+dN7Dmx5BMfdn8GOoOU4k3OyLok8K5ztJYagzMgvrLMIP
hX8SFwhaV0g1pNsd8y0KOxA3l8ihswxnJLNiYOcJows20TtXpOm7GJMhgXsVtF2k
XadyNXBjtqhCRYoIiq870rtvxv4i8Oz6FxESvo4AoW4k3m9kghIESGcvh31Wqzk8
DrOygYHpjuCvwU/oITUFfRydYnfKPF4ed5BiwjJXcXMyjfbi5iJAM0cj2xrFPxjW
TdUyhz+A0GmYORpfLlAIFNSGbiWKpB4vTonwqMQ+jBBGb6K/pnixpHNripI5HVvl
c4BT3ShmQk0E0U43J9D8RXXYdaPs+5O1438q1duP02cqoGBAX8isqCgBhAJauH2h
FHomQRN8nGJ9/TgFftWH3lP+H6JfbxdR4PDYO5dA84F8NKEjpOU24Oar5YTVDG6U
NYuJ6K2inzxMUbS+ehqjWMLhsNiSI0L2V2ifOqtQ4JopbnvuDDfweT63+bhtZTVd
S61H9UJD5bOadH1IBhj/8becTeWz1MYQeH8SloYQqgNs1BmrdfG4WaP9rnSFLR1/
gidx6qD35Xy8zpaCPYF4lYTW5+qMb90DuK0ibRz9t2OcC16GE132M4UZgcTsF4mu
rvP3nXbmzLpKrZ1q+p+i32y0i1tCUrkdg2/iUE1DR/OiCVDj4QOKe6jNNNnUIHpl
r6kO2l3g378MDh+/s+6U4/SxhWLMHe7cmts9swaJxeXjhAlcFW8iSiUHejeLcof0
zmLlt1rJd9q8K8ClkJDVbnM5FuMx5+ilrf4xfmEYoPL94YhAd3Yja1ls5/CUZMTS
JrctAk1EhpR1lJiG72dh590ihZsUdUc6YsrEXQly+xoh0VAArRvldxM29AP7efXh
zBCvn8Is9izFs8CSDuUoHCqTam18SrgqGb9eYTgzokQ/qEaHj3CtReoXm4dyQBqd
w8xxyE0MQmFXhQ4UUa4qyQU+It4+E7fZAtotEEsVUcTgI7LrRJFxO/IRupT6cvfj
8q2+Ni6Maw5B+JI3UstJPIw2vsDbabxvdnhe5qxOvxhkqTiLCNbzjG8s3rxgNlDv
laYruncrzYGt279zmALkrMDV72PmmTVpZS2oib0q7BgXrKm/Glo/hef8yRm5b2xf
kLYCQ7nTvezh0D9yN8l3UfDNGYr8o419ckutBuMGl+OXXGRBds8BR1kPPH1fP5IC
QCPBpj6PH8T7m5rXTGhhQLI+2iQZy/pySofUFloJTkerdN0GUTVBYj8jLZ+mZgQI
v7z1d4WRjfr8xCe+/+w6EhscKqkL8k78V/CHyyk+a9QMymsroNKluhZyybILWeZQ
+3bXI8wNsumG5qFRWuLN9Em3yhPGPX4q9pPAOLmdSL3Lp+R6C7npWGUF8mPtrMm/
49wyD7rzzn6T9bB/lPkkStAXSSpoUEOKhPnndq/CDtnnA3dTwzq8h5G8UT6h7xiO
ZWzyYEwiRytm9XkBJBNzmFijSEzuXXGaik2xKjo0v4o332R/liBrCsuYAGNB4HND
lTXzG/QuwrBJ7mbeHv26HsefvGt6bLbylZmiUkqXat4SpUnKF6iV2gP6jdILRBQ0
NywUNaFwugdCEjfkPbbpSw==
`protect END_PROTECTED
