`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/nkpNWjQCgoE6Te3wRMvZNfDDuedhHLsL8dmRSkO1TCbtaMZTyw+f7aD292AaFV
zQYwwQ3BtA0speYRrubzI79wbZ150H38UdA3fMr69l+3OsqxHtVKCb01wms39H3W
ieenBQGBeGmr2RilngWOLlN+G5PCJQtkEdnn1g6BPuU+0UIYBWM8A/JowcN2rjvC
f8I7IASF2AJmHLqZvEJoz79mx3+8z9R8qV+LxAMti6O9+WHEIDO0MPucLhSf7KFO
4o9jLT44uHqUnGS6xp9lHHN0jV+jjAGNN4cHvXYymPbdqmVdd29gbWo4WHx52ly9
I6hg82X9HVfTsdtp1pWNfT21ASq4wVQlFTF2GutvxFcHm/zHjKlzMA/xJGYlsDWA
KB2HDH7idwuFiFACXZCRnNnwpCq6QJg779vdRiC94R3vNTKrHf1Sa8ywerSJ7LRE
O+6R+ndumJmPF8BFDPHxH0XponC5NdgaELV3ptbLRSYaSmeOiaBNNBnZr5zuDA/M
DEyWvDhZH7VYNDHLhIg1q0L+UaBlOfqrqLvGolS+YlqA+l/YsJ6dlfs7Y+lGVfhK
UGSRI6SeHMHwM5+cBDSN51OiTYWp4hAeDV1Dein4xKZk2+mwP/elIKUshLJEvtSC
FG3CWXz18QStmgdQaa34ciHthWa7SFtnMfUyMeBMLSQyYsgK+ceXKJxurVHWkuKi
8MqnwKwAlar35oLNFENVnOIfTZTnLNX95PkeWzW1KoG/GCl7q+RJgU0fOXJggryR
qOuQhpJOxaYA+TbGtMwfamW8U330R23slkGwkounEMP2clieKHtYs9utNeLEyzGo
eRaTnx1sRyJVbFZygVHgbfrsBss19u8lD/IEGx257+YqoRPl6yPQ0aP9n4QMrat2
kPeSh9wwkpVoroBOEqIQ4gBbg+Bw9wei2ndtnzIMohbGHWy+3PfaeVdD4ZKpYSBw
Q5w3A3HSkgGFlYxHCX/d/uSnNrkwbPJOT4UZn9Dr2v00h6MTK5MqFaCeEFcCcOSF
Apvrp7ck5kRaWV55OZT/pc6jJ9SCFSzXu02b5Ztin+2ReAiQAGhQfVvmXvFJqBKb
cXSjuNemTgrJ4Uwh/6N+0FxHuoy0xdZB3cX6ifNMHRNZ3OaTLnI1HNs4Ad/axyka
IjSuXBTkfbClXaKKR0T9f/8KLd++UsVSQc3r3MeVMIwMvdHkOrhoyNAkRvdWfLMI
gnOgSlsZoHmnXcAaFH/offleaKbE6u4i5754erA7HhAtz5zZMTaaRJibzywa+j8C
ELQkBNmnrUIg05tij2kWDv2lS9wcSGi+1yQeaQDjHw7r6/ajE7RJBza+7fNx52ut
FlliBUw/32/xLssJGJwChlb0eFQxO+0B+z0gZeOgqZHHlH1CQrKTMu9jwwv2jXcM
S7gegzMHfssRBUSe/Uy0IvpfS2d/ZeTyQpzk/xUy4zs2P8pVz+QcxZQPBI0culMT
DRWOl+WL/ZV4+rsrfcUsy6NDtLnl0Gb4YZOcpZVkWPUivWNv5I3KXTlkr9ksZ2X/
dhc+UZD5R/bjBCYK9Psctg==
`protect END_PROTECTED
