`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZKP3WL7fCUtIc/gF4V82j6zaNtIn/TEbluHHGDjYEcZXSx/PClGxvnEds1fH5ySv
5m5whGY0lltaio2cTB2mxFnbmVd/DRNjjTsYDjOosBgcZAykGp6dnnp9Et3y+alu
D6oclwRB7KZ1ORAwqVKiM99tkZCORbHdx/gbzjlDy1YEpKiDMo2HGZ7QKyWnNhOj
pI8ru8cYwJvuiJRTdojZOVbzNeSFSBcZ70TzWMeckZPmW4CU0QEYm7y/s89ElBba
q2Q8OOqrYYk8lK1t2Zt45nKwGkGy5O/GLX4Ifhg+oHZX5aH8NJl8MJwsAXDVd5sW
y5Uo/dvmM2gwV/M/oChdyYRhfalW8E1C15eE5jEeaNaD55nBppFsQF9SGUziV3lR
9/jIvEwDAUDbFYGkyNzpGWOcr1HxxLVZE2etdYDa4pnHYFQbgOBnCXQkBTbkp3NB
TQNwuB86ATFgAi8eHZtIzZMcOvKU8z7HuJjnbESTwxPf/T01nKLJ2Dr1cAx1fFaJ
tbJYmZJhjB47+SGzJ7AZtgOqPHNosuFvvZVvtKOznrgmd1NeGWBm8yM2JLSCIG/s
pw0IYr9ZHkOx/fBeVBQWkZ48PYgjjgWYH5/1xDZTCioMFQNIhfDUHLKNTBj8Udd7
WPx1SIsxi80kwm/0CvUGaHZu5AfZpxrnDCkxL/T+HE1yXhyaedrHSGqrJJsrm6fu
Zu9tn/HN1ZhwXNprr9VqOt+tdEBrELYaJ+cJteiQ3pxYe3h2t1xhZHpTFwv1HLnO
8fC2jhWLqM7NJz7ZSR14O7rmDe3/jd2VeCflytutwb0qLEpAre0hD54/yv8Lc5Bq
8/6jJX2XyZxQdYpEWxM5Qk4bXwwECMemSyhYMbtMXK02pFA3XA8tXUaH30vKZThD
DL4JuaPeKRKQsUrszjJV2HTIq6EQnIYun54TwY/R+aL2pYI7j63MS53UQyICXkv7
F3X/F1zOaw4wgVpl9/kRz+liPosHXGe62wcswb3M6j608xLKf+aPWwmZb25XlsPq
0M7CIBHlKWqLfdWYELQ6KGEV1L0e1sTF8wy/KDxv6af9uBv8+CtDTi1xudB2+GQH
iiIocW31mw6OjOK3fdcZU4Afubj7PF1UnC6wj67VHS30EwusYhaXL6I4G5T6cnMG
OBUHkz0Jzw9LOuIfsWyQ9n3svJGcgNR60tcim7P1SUVbzG6+fYTXeajTqhFVf6HX
qQeoj6orfilkLTlX/us405TLhxyvIN/5YnCPqbaED6Vv4y6eJIXnIMIiblBr3a+2
aRK2Ok5EM4z9UG4UNQvSVZFeWOs9Dpu0gc7KYh2XCG8Ymbf6YQufTJuq8Bt+LqvS
7Zy6HdVponrfkAQh4ucOx+HDITox+MrHh39qFVAjVmKW9szTD64eRrf+RO007QPx
QSIN1WJ+ie5HRvtrGqbA7N7XtVuEVbr5X0wzGQR3X/jRFQXqChkos4uI2RC/Orha
dHU9B5R5W9fqDZ006BUdDe7s7KXZ1GHfsbQpY1m0BUCttzGDzolkhBuG7U9VEk72
lFcv+tE/jQTs42UYvag2FNW5qxZlq2VlwJxocnZauLy/st9iu925cuE+i8uXmd4z
j25A7dfQYKmnhByqjd5j/+vSefBGdUQ7TQY5tAs3zlCjrQ96ooH4zTLGqcSbjkUu
3+Y/YnEzBTRJYXplkTJMCJZu1nV0fMbYmyNYD7umXjtVokOFrV7O1J9RUTGgeYpU
FeTaXurpVWtnBV6cKmhVn2s4FPzbzrjuzj6QZoZnVrK10ki5XRaftgR6UtYhDOft
1y+u6UkA/OPDcCX7mefWTBUJCj44LkYOFM8HlH9x/LVx5rYbV2viCkTMJbReAuIs
GSHib1//1jOES4svxOiExE3d+3BWTuWB+Ot892owvAQRIJbeDUEXBSXV+JQ6XElE
gTn7SvNB2tNPhCJ8Zcuj85JktiCHWC9gdSLKYWXC57zI+zkgJ4L+jJT6Ep/IccVa
YnVUwN89jJtbSBOVM8z5nXXD6zsENbCGqUx4x/mLhYgo9DXYHvz4p9XbNpt9nGYN
jRTpyDCjuGnUos+zdvNcIqlsUJdx+DQrWoiI9VOutbVO4+C8TI3MJbiDyBP3GElt
EhXdh/jjfYxEt+7jRXjRYBSfcTjsTx3GuFotwIrcZyZBXJ94b+phHseSFoC93lRF
linkwPNB5GAcUEhMk5cQybbiin5GHgshelF9rBGMPUYWpMpiCAwaa2/B6ZXu3ICB
4ax174FX/9rObTHlIk4F/vwlN6vc0IoRK+eRFKE4oIqtOjiv3IcK0fOa2/o6SjKu
bNWMElaGTuQafRLcufQAxjxOhaWZTlNcE/R7JO/pvl2CIm9Ui/KG/WqJ8Du8UmwR
XJ8qgm/YRTeI1Aed86ZTtSz48oWZ+6wM85D1Zc9u8WNENjx/a5UdZMlfIfGEc9ci
G2/aeTzcS8qt2MEI9JLl328qFWyXSpF40eBAJucnyXHnWmELWgClMv//p9hPZR5S
7UcscRMTmcvv84QP/nCSVQ==
`protect END_PROTECTED
