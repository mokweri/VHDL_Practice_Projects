`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLkWUnKtVox38klIXOuXfbmSC8j1vRqdFQ0cgPX7/EHEyOmZbBs3TBSxtPJy+iEz
WJkk4CLQSrIxYndwnMNTa1O26wu1Io32XN0MwLSs4p/JbAZP7PM8QnSwkvHVHhcq
AAH/8XiHICHQZVFdG4jJ54vGBss8rN7RPFzVd0tCZyMZ2ibjs/8IG3b2f8lH7I8e
TPxDX8Vac+JTKmzeWCgre9XpP94V50xhHSFdbUXVKdh6cRB90/TseZ8DrXWQhK5X
dVQS8Uoi22g8AmUtxULo6GXv+QUjiThv/kTgcOnarjgr1A9wXuj0xSBo8AcSr3Qw
h6/L3WNG2hTqWSKus6VA24OEHPe0laI5IchtKH5RwL03SfHzPQGQ2ajo7Fu851nR
OwGLr9G59r7ZWfVLV/3wuZ/HDTMqpy2q7bawq3Te1/DXTlG5tTYy/gNz1rsaeQdi
InaGoYRuUWrPtt4+TmPCipOj3DGhzKLu5Veca7XpzqVFrleYM+wq9/8AIrwQ3dOd
ww2avcIwhtUHAtBWa0pOw7UbYOmRWcrxuZ59f2tOBHzndFp4FVomiQkjkaVtw344
rXCIFJaqRZBfyK72iQFML5vTBGbQbDRRz5C6tgmtoAGoVZunM9sNYwobP477z1NN
grIv/jpYC3iyfMApOYPhi5JJpV/gT0LttLtK9YmzH4k=
`protect END_PROTECTED
