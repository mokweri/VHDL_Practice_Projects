`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uxh4UKFPUlQPN5u6/N3tk+0U8USYRtcR9aRFw9xRXic7V2LST64eOgVo8Y1Ve8YJ
3gqvZytA+QTzlhlvX6se0IaCI7uYfn4hy0nEDYvmW+2NuyP1aPqrjqCCmQ8K6ijn
6M1/kIgRatRT9Dn+3pVJfai7MdBiluROnVEDnHTDTHBeXU1sYspIF1MKTLA6Ais3
nUq5zhN2JSqAnSQM+1/hmWw5VyKgw2ty4M58Gr6HOXOUAePi0kF1WpnIrC+h8kn/
uLeMFDTHQG7bFjYc5t28SUSntyAt6Xux0o9+5EkNexdd4KU6LGOccf/zNBDNR1ah
FYGHZ/hwOxHq3IOeMM/jXWUDUGlpErhTbXEA+IZEop5TNGFpfoB5Cr0A7qnRJHI7
GQgPn/gW9FbF6xpkReYtiGqxMGX594pgQWuAeg+WA82u2Ja4G/03x405XXJieKGV
DEy0m1CjR12YIr1EvYQ5oScGv/DyHj+IkOtrWYtHwr8o4t0ffV3PTzMLfwxXxvsZ
7gYIzMaiUMAmTOzHd45G/7rJCcoWmewyFFlaXe3Dc36f7dQk1ZX1YswvU7R+r5UO
8YQZ5bYAhwJrb2Cqv+K4HpdV4mKd6eRd9WolJE58mK7KfjuAZEPPrJBCR6eChvd2
czWd3Zq0YYXO1ARGLVp8ezp1v3Ytn6291KWcdr1flD+Bjgex6J/9EtUa+fFxi0Is
bfNQAy1N5M4tz82C/QeEmJjYqvokD/o3TkpgYEkMS+MawxsgLIMlSHwUHQ9KDIxE
sBhkJBwtD5f1gbEDWWRzAEjwnmL2j8q8MHacomaVxTGaQ3zk8x5RvNOW1grTx26N
fRhOTC4PNL6+hnPeXZggq/ZYHeCQiwjzlziJpe954jD54EtBqGM9BNshnSJYNunZ
VNPg5G3nUfxBZmYEFkmpmt5xK2DmpGvSNbavXo0f7FjbAlBTbSEOFtb6/d3HLndp
Dmvw1kk1qPO0z2ecL4XBfncS7PZybfZkcSj9CWBtwe4XBJW1/zlkKBGcM9hJ8uwU
Dy5IOYwXj0M00e1P/W+Ynf4maz8KZAugtTvWFqNevhG34bhoxLKuhedzuUn4ybv9
KvAYeBUf7aLLloWlJj8rW2VfK6pO29rdneYyg6LvMPtika3qJz7K+jaBjqocitGp
z7qBpXnAxwsmSEEoMWqqGEiDRpP9WcHJVasI1Q/lnQl3P6N8asNBjMwiMbHN9mwL
zKR+AWXaYFG6DraTxjv2U0LVv+9XbVQYXWS7XN/iMSVdzkwZ8gxSY5gfZqUcYNm4
RKeMVEOe+4DSwu3rx2QUOTJc8Jy5a/Pi/aoPmaO3IqsSRRNYhdJZG5vvb7spbltT
nUi8cngqRpAg066nRAVPqkeFLsteMg9F+/J/i3C4BEaQ+KI/PUm0YxwReUeEAgSz
cp+XMFLERz+dcFZLxWcjIQrWmY1B6/DX9bSMRUaSQx3kiQP49P0stwAw6W23bPW3
plTtuW7GVU6R9n6BB+JhWX8BIJfUDVrrfcmMYlOGPf5hlvU/1d5IK8b/DPaMv6d9
aAQ30zzkbRj1GsceGYoow1ekJyRbYc2n+bAQXxRptkveS/m8KK8QRziCQzusCtC6
wJrPwJyNKra+PoTvF/YWZdp4sk99e4cTb97OQ7NlXe7xV+nodkPqBfsJoTcXu5Gk
pgrK5wg1goSB2Nq1jaVZOe3+Chbmqb7kOgE/hhIOI0WwdEQsRMsC2z/ix1cM3KFw
QJjFmkiiyYQhfKrMQaatQmMgKIzCYgrvlTLpbTW58ForWHQ5rRKk6m+nlSOe66NM
x1JfZRNq1vU8HNGODnd+frvKRReyOu9yUoGtFDi4CMBdG50bXxdVoa36IEBvzwsp
gQ4e7ED2KelsA11eaZbjQuD4rO8FjS9jNYaEFEiGvrQuiAv3j0BuPufxqbEION+9
MiWouJs0kHWsw1qnfY1jumtaLgjjXGoCjYU7ZLDGGFiB1Xrj141KgKPH0iHKVTBX
FmzH/f4p6fbrqXUkFDn/cnZh4C0/eyKH7v/ovFSiAiPZZzyxoNnjbdEPq2oi4Irv
LNmWLUoQn5W1pQr/ZckwVyN/CPSNMM9GrjDerEYtbD7+igtgJ1FahIy0dn7uoyM6
LZREl2NRtYuNhvvo6p11agcIFtRDwyD/AGNA60bpoSf8/rVT7PjBWGfFFdfZA0RH
Vze738l4XbFHL/rS+xGElYqWKWPun5+AjGjBQF4GUsnygzCXp1zLg6jz7MX5elji
jhefilCHnuDG3BBuvXM3xIG2J8iz7RSpZUogV+xjtfHL/Kl0dsyv5fmnjvzUlpbo
QETuKU8Bd0tRkFMdRKyVnYlKeuJBcYLqZ67C//jowRI4AQRIIH7SL+DOMJ9Hqjg8
jqnLJEkaAreVUFtbDxIIthmHd+qge4yfKbvRU2wDrfeymSd+R9G/T57UttuqcWLy
WuRmXy04+HwaSXOEdBDZdk1J8UZ5JCZKKnfz68ODfyKb1eSI+LNr8NT/h7enbYRX
jTn/NL6Qmx+zymJD/gaUi6vfAXs1lmpw8eghbF/dKseCWJRcEYDYVG95Q+Y4lzDL
RHtqxf9xqCk8JQgbxm27uAvcettfuo83QXHUbi8kRWwb2Bz4euD6nrGz+fnXDukc
NNhVX0Kn/uHHnndk4exgmCgwcQp4YrlugYH9M7GGB3VfcDs5P5hdbu2Wv20lnNe7
2Rqyg5Oj2JUlBCRrnSeHggtMDs85YOlz/aWrOZNoevoUcln+JTf3r9bToiGiQlTi
plBQmBmwSHnvXUjGVlJNfxe+5xJhDVsUu9oFNN3G2psISUVKADggtoQbGxrFf/G0
+jHrTDdXZc2hTy8d1vm87rfk+2w7Tc07EbjCv6Jy99PqXiE8h7eMnuslNrWwG5ch
bQGbDrAXigjI25llrW7ZCJ1hgWwPJ2jS8ANqFsB/NDe2udgp7Cit9BfQZ867qwKR
CTQqlyisyxXLScCbEPKcRzmFuQh/OIMVAOlV8EBaRJhXtxAgrYM93Vu0Z9pEyPsn
XQO05zCu+cAWSlsYxLwrVI6vdFhPnvwDvqp0p92CIK9EPFx4+DZqrpYYyZVRmAvr
olAUs+6OwtZWffQ/4bM079fVFa0nELNbyZPglV9ylfJObXy6OroSC4hpyUtyorjw
LpiLqBpPSiHQUqq0tkCtDy3WIBC1QpSEaGyMEVnjPvwLrK8yxMBI6yFKzSHXg5wA
1Qbjcs7Yj7Xzs6z1sL61JdOSQFqrhR1BM6OS0FrcoEOjtGVWWtIwEqLG9c3bk+bq
vw+5wicDi30QIhbB8gk6xcHlqHBp4aqab9YMtjefn9l2NkqYUvZPQzf22VDI2wQ0
5c2umPb1YyE42rL6VasK+Tdn6Sls05cAkIoJyZK5XPtvmMQAuVQkQrmS8N9MzvXf
90ssTTdgOSycsOg6MgxXb8GfyhbqvhhkxjXeaoPgs1GwEliEYQK6wx1T5sovfygG
1u93rPjxIxL6DsX2Fu7IPZ38j4XmClA+llk7bf5Io24cvCDM9X5varOPbvuShrVE
jtz0aOH+yg4DxkrZhu9d5gS47QDSb2h7af24Azz76LDR0HYUR1UXTiVy44s3QLed
x+xnjTcAIkUabnfbI/i1/Gb3FEI0cuqazgmc8g1B7B3klUunYEqj39kKreslsQzi
0bkYXUjnRAOSnKc8Mgd6vCmgATv9qwymT/Rutmijf4TxwIGHpEGFdVKyYADdY1AE
LoSE1eID7/ML0ujQwkgkvgJTCbTnTSnQujvWoqu2z88Y0Fhn9KrvaSTctgMXi1Ei
wrd9j4i5ajmHdgGhR1sZtkgfBH2ztjttBmP0RC+I3zaqxtAGTKXIlCfS5Ob1YtRC
rYsQH0/8pkVxz3yU5V85CTjdHyUYWi8r0hRxliAuT3VwMZuaoYp9dtoUTgw/NAmh
krUiv2BKQ8bw6vglOIh2zgAFFphAx+wP4msSrlKMvM8pfXDuKtlwndcQ3PjNbmky
V6MiIQMSOwcGQzVXUZzwK0r+QPW/CXRidQPdInQ6qkB0gN8HEF6Z3u79K4IpGHFO
stlUOkZRC5jaO52biJSa06vPXO1FtbCrakav46IQ+qBwigNzxI6Xt6XwB6FboDD6
dA2EB/dHZvvnsfNGitDglWVfejKB1S3J1MgzYKELAYxpyalD37wXdksWa5TaBDys
7iw369HyIxiMFWYwdXCgrsBMEvhxRezv8keGpy0ihycp3g9t8e2xSgWvashVgvPE
2mZGgOXWftc4YX07bOybqAY4hlefURfxGcpf9+kMLmS+ukvFc98rDjILRr7JaL2F
b2D1vaQyEvOmjirRO+60k65/6VSZmDDCqQdweoUpG4uzN/vvgAtsE3unjI6nmqxt
3vVTTWI7Lc7CemZTZIXLv5DhOyfA94PV+tCCXdtzDBWBrdZAgK3Oxrw7MawhkEIt
o9MtoNz1cVeRIrzJOL3PCZT+m9XbC6MYsbjiqVpN89SGDi96W/V/DywvJXLuYe0f
GWgBGfYgJMucM6Xyl/RxTIvViNfieFFHt70pZCCqQrOvTGihPfR66zZfJfnKc4pP
YOq5jJa2akjPHuCqtIlTp5GFAH6uP1P8DSqUrntfPejlGikFcJh27viVE2d2XiTZ
gscc/TK3khgHQNYacHTCZJdKQMelvbTZVgowHZJI0Hp7GrefnLHMAuWa8Svi4dYS
fwUgHnsaoWfPHZKGrLQCrAkmabt+mJQrKH6zb666nMsLdyfGzc0NogOjHOHfHHoj
xat5v7lnz3qQbVWXpgP3mNSSmbHtHNSWxco5Pfm5z1ui0v5z5Vy77lCsUDzXOXne
cb+5eM61CI4U672d5qZ8ruVXhgG1hJw44Z+/4LCYFLpZiMgLW7T5Jj0ZNG88nIXn
afQUKkHKbfN/tE9lZYU5D91MMm2sbXa9ZmCOYyx4EgQ3MYa3uOpiT7/hhpFg7KF1
U10xXSsKK7rI+sRQeRv39T1JU89IZu5GvnDITFjqFIGyZ/qpWpMU51m42GRYZFOm
uay51FQQCBajaNx9EDcEWBdqpLHcNBhHXNPnHKeztk27ULoEvt1fLEuadLhHSksA
IW5ypmK3iYfz54QhnZEuoX3afpXetIQmTWpPdX++jT32tG5RvNIyfjO19KiS7oaz
OG5aVq1OkLs1FbVbIbpraUgdzRxT4ubLm7zH2XmRQwCUIvJanV00Mj0bDJF2s9gI
NB+jorYhcyJ+0KGWxlt/YVuRh77Wi36dzNm2I70yEZEW+s/or1a7elzBeDGOMlJy
SE3mmZvGXBVMcB8DVuW4On/5ven9d/RdstOaxmI34dDQCppCxEGyC0T5h0T6BlcK
6ECKi+deoUkoiD+CO/05/vXPSf4h83Eugvl+NABUWdJQ+i9Yv9BsReJn87OdLQQ2
YF6qojyHSslvNoMQD7RLZUPui8nypyO0xeEXfl3i5tdY7SibV41lCgV1ImETvyVL
FyVY3nj5Oel6cj35gyuyqPrMOBABq1SY0/8QoCHema6UFUKhwtRWvoUNABpM087C
/btxFbLK4g6zrGYfycuNcXzY9i11siksgNy0zRTHCZWWGGWbhvs56gwpfp0Uyvv3
Wc1C55SHZEOdVdrY8qe2EWAqcTLnqT9cMyQz3zooAEGH4PB5lYDtJmzqE0zW4b2A
Ai00n/fu6FzkWF2cEqiaJF8zQwL0Cb86DG7M9Ay0oh7Tyzu8tRmzNwlevpFzZMDo
2S6JxxXiUzerNJeViae1LzCr//RdrKuPHkyBELpt9UxDE8yiTkZ7yOKRGrFuC79w
VKOxDu11bqE/niGMVHw5D2MoB7wVrOHWubUxvXDL2CiuZETGNjCcGXre2o4gyGoD
jK9ISj08jPzsVuRXo80FIBb2D3d88iRNWbG0WDOxzn0qbf6iUqOjBVE9Zgetkore
YzaBZn9Mq/1QLk8+hDi2/C4jznBVv9DxKou9FngsdZ8hNtVHggcfQI77EMvzGC3l
DqJyR/rJw/3NTVNTy1OO/jYzO9u1xiwMnlsk8ILPIzq0I7MWre5Ui8GWmltn/MtH
pPDJj+hd9ZdK+6usxLEU2bsPYEMBQ84rw84mrBrGpqmR9pQ23EX01MwOOhCfUHkN
2UsZKbLov1W3DHOfB2mMXcvHc53ZN1CXZDgTfOViTA0/cOl2n9P8Tp3qBcC+tl6s
bX7FXJXznmyQCPhIndmg3uu4XE990CTwoXdGj01J9gwPzq7fIKJOgD5E14Y48J7h
TIjvMEIfkqxbxf10aLVW/PqvN812ZpEa1AYV2CBX3n/K8yXtGzn3O1i9Z3SiJQSq
t7ASoeumBXaZ8RJ0h19c2kzIdcrminEnYs3Iu1Izx+EQDQX4sZhV6VDYks4YmIMq
N/b+EC2bgV5leVD6CffmGWz7bFg0wduXAq6tmzYBFtBN37hPeCXcMGoPkDFTqHDD
DMim/+3p8DXC/STuos4GmHnGjTIrTV97EMtZF3EqF4e0wUdYNn664KTel6Dfb35A
KVswKLP/xCJ8M0vb9Un3o+/66XKrjLPUrOo7px9chTHxoY+WKkCumwig7US2CZAp
8/7FkMvFeadTJHcOSi+YJAKBELMh4ua3fXHmOWD+HMFMEKF/j8hEPDPWy7E6K8z0
Hfio9OOVhoG5dpxAJx2rvFQv9lKXveMfEP+/a24JFfUqvq3Zgkjke3dqnRQkaf+7
JZJ9ujw4sQLsiY3y4trwKtb9DMLNNrPl+lNiH4cd3c8ehjfTvtebEpccIhCAcYvM
cQix1ChFQ8DdUxK5rh8wpWWBXxdTU091LHm8MABU4EMfuSvsAjahCnbFizLw30gi
If0u2zIMea139QpnSPtroAka3htlGF41HIipLQRT9BdMYFNNszI4ewH9/IAcHzIw
88oRg6q6ys/sSmt0keYZZxZZ86V/WJK2yIR9JPwjug9068trpPWkXxJyeXte4nzB
7pLjS9/+q3NEDBJoppHlNn5iBuGHJ7zTpcGmFDlmGoWYaZ2sSrd0eFhWXDNyq8aE
nhrRd2gpHdVK5w9tiPcRDWQuuBdI71S3oSp7tmKmEXylQF04e4/y6sqbA25uKPzG
8ppq3GZNm3ZtoLg0AtMsRTIZar+Ck9RqocQQYoQJRHHxI3MzhXeNwl1xfvKOECAy
jZ01GGd/IE/vMTCd6LJjTVx3orbk2awKIch0Z6cm03F0XIKIKrq/hn6uWt+pE4Ed
H58Ycp9GIa6BbCI5BKs9okghTCUYCx+2X42qzWfsfTOLMS9+z6rvfjdSqog0Cvvr
QnA7q5/SJvBBPdN5kgybxv45tHC78G/vV0tQy9NkUwyiw/KzB//yWZHIre8yYAIB
MXLwUSkcsiLNyKSYGwOAF8dvEMG766swgC7k5mKxOUa4/6A2rPcQLMC+Otsv5EI9
XQuTBLgIkXOYV3NQr1/AA+1jMyhjBSKJxlNT/hljYnCMEfmIztloYHxlcRHUgfbN
rpizAuAIVJQmNgAyTyOlseMauq3PpoVbIZR7HHLDTIhCKbx1ew8UxqaP3Z4xDSE7
NewKKolTPGEmcdLkHL8CJ2U/mfp/Bu4iAGxipoNw/TYSl/F8CcManqqIDipNNXPZ
gYl/Os5sReOcNPOAJQ7/6MQAfBJUgVVUHPPvUCnAnRZY2Forgn2fD8Y9HH1/XGU+
n5Kax9XlzftyruIW6cfEMTru6MBuFQM8038ywyialFE3OEEEia6EbA7YHL0BrtF8
IOhSJFon6tdWUA34vHw0AaoAfd+fvuWjpPxkL8kdDBN2C8bFgW9IQ9rVzj0wTegp
v/I3+hdxMHefSmAAuI9rCVRNcR8XUMYweeWgtzESRj2F2tVE7nHWouhw1kAYVV/H
xC7ccuhfnlHXb4l8r2r4LqEpMwbZrI73vezrqkJmP3ItDdxN0vY1A+0TU7E+zm3x
Nc9fZOx3yB/53ww9DxNkglzA6kYwyj1adP/TNXn2IgYPnsxZvUIsZtbpflze+wP/
nf0ue+gNzjPkc3Al8qD8k+TfdAeT6b8G50RdRHTH/cdbzpWQBfaqIX8GG0tLVPQE
84Ku6Ideqg77g/QVX69Y1p4nU6D+VC5zVHMjOQik3piUbhdA5OVkJD5g4crRtyRE
5Ari5RtdTbYxqzZlVEi2yUA8irv+denHXTEBLDOUFH6KOFIC2Esmhs0R8o6iS0rp
30RJVuqHl3JPjEUmTFx7EpWR4d94IyJhOKmu27CZFWvG2tRZ395Q7/qHovuGc2U+
ou4dilVzCIGOUUjjxtbS5ohxSDRwEEZX81djCJdW4YtUeuBFBAuF4cz+mpyz0Wto
JNm3UJVoE2N0uhC06AmFsCjSotKwy7LKfVUhXBZcJGA1EuZkxP9CHnuTqM/xLTJ+
+SgEkxe5/WJbDbw3yl+veU2hglw7GAGEiHUeitLgB0W9XqvNsh/Fp22pzBxvPFZN
D/VORkRL+h3o8hYokDrt7Q5ueBq8POMZCu1AupO1a8n3/Vc66D+Kseo/dNatpOT/
eyS7zX13UkZkdPGAGfoZuU3WnxS/wUa5+wC8+XxUFO/6d5jEamGgvqF2tUxqJGj4
sU10JFfRkF10+RTNpli1ESH78FqrRZ1O/QMYP3KEKbo9e0fSGWiiA8GAJKdU1e1F
DjNNz2DCmrCYll8+PvHP5j3l5/8m2/rJ4XJjxn/RYbLWnguD+dEy/wXNWIPlbfup
ejnYMQbSHRYMzVchJBs9v3x2MjYgPpwNp1ATJiSCHbFpaafxpO79TX3YJii1tDeY
mKy1j0ylEvlsZYFj0LKSn5BDcCV9dFuQInvv1G+flkUH3eoezWLyUy0kUvUv+lhX
wFckYkgiDxImXyDnTaaMktQVEeCKvvIkPs6DT7/C9hYVu04gi9OFq2YKLNXQ7VJg
tr1bdeZiRJS7OMXwXQ/JL+OVHWRuItY9QyQvyzqR6jcTxMlP8vcrIBKWPS7cUxTf
Kq9LZN4QnuIZUukFsCzBXfmcWAupS98QjmvewpFofLYRAo41RvCg8y3M0xFi/Njf
wwVltWQ7Gej98iyA+NR3XmP0db2TyVuSZ7gnWR4OBRu96sP57lMm2Qtl7l1V0PfI
W8OwWhDrfCNZrEzSZHc4F/inSKh4Fsbrw7p81MZTlRDytSYrC5ADG6J5POrIbu6g
9aaneRntPrTlNID3aciWQgxrbbnkm1uBF8HYLBZvB5FYT1Xr0juPdkBl7etvJnLG
O05jEnAe6wUivCkACqvs+F9D5Co+gTXhElWeGMSg6rqtpaixyeS0SIn9vqM8151v
OOi/bEfLjYXtrXf+wneYp3xfESXFK2xqfsLvttGIpTmRC6dNuHJFdLo8vzz+YyWF
iQqo5Ys8WGRYC7CzfC4D9eW0tWupk1hB47CdWoHeJDE8KfO1A8tdA3fNh/QkwhEO
82mD/O3n+OkiIRgTGkXrdURKbgE4/oSyF9pvK0jhst30x9BzR9WhRH8gxy7qEGis
NFPvjjxt4YJa3zpb8Xsab8sLTwZ6Y6JMcI2sqFy8FhQD2C/8bjhM+4UItOpnEFMM
TaH/SlgVxvPynP1r93yTHythZCSUYt/rnx+ihRyW4msON7NevWqkNL3MgkIg7Bqc
P9KYTtnFz7DLNBApe2rCyobJD9YXHhcRWG4s9pdWPfHfDzVQ/qNWrC1AMBjAqKe4
fp4SC7B+S4f4y/TigsoWH6SWRAF98S9c8HE2ejUYf0KJZlP5M7k8WnUgMjyV1akb
ur/KeUrsBfR7B7pwKko+4KIcr+QmkSVnEtbXHQWgogjMmrAgOJFhewI6TyePA7A8
gHVNLvyZ/+vyYslmwr4WipRzEx/Ci/LpaviofZ/+FPq6XzOd+OzCk9BkPFL1I++E
N9wuqd8Nl7hwXbudXg8veGhcde9mAk5DJHNjvg7CGaK1ZcOvKXk42Les9S+BWJU0
SY6h+XJVSbVJkWGF4Kld6m0pwqyuxZWm5in/+ooQm6dx+Hujj+2JJFbuHY0aCtMj
/ptrP0RVWNpfKzfwawzvy4o+hjPDMjXKDCBsC3HqQywZ+b9MSatvaWWm9hMEID8q
AwMKDAaG6rre1rq6lHM3WTfaDG+RPO6jR+iB5ooRvIMZlE+Rtg5aQNpGUnmk38s8
QR504eBFiAPZz4ojUNr25Ac3Z/wMs11i78BuH8b82RrwDkD806O8pi+tJVXmbigJ
+8lNgFBbpLSnXS0KOCmdKSy4W/+L1TIBSFlB9VkqZ6qmXW4JHxsuEFpxQJDvOWW3
ssrjf7wMVtHraNTjayJFoyForao7dr573br8r9HloUuSUIr9dgPg8H5X+Gs7Fg8P
C13L4Ty3mGUWOpl+C4zMQ3UE3gx0LZPW/AILUiO6eLJUxHFNcj4DLqk4aGtAsgdT
e2jorkccTkYChZsRSgCncS07TDYttTPlGY75TMt7/zRP4dci7vLGInZKNuQfnjS1
ZkUFPbspXNRGrmA4N4SIb+y4vlyB9KiGQe9u6wKzwX3M44QZIoGFRsYrBnu1J8Kz
L25L9Xvdq7GemO6a8eFeCH1jY3kZRLtiVbgEecpkMCzKPEyUoIIdFcGjnQZYf7Gj
QA6Sxe5JDJlPBPv0083mPerGXYUn/01Zo+kolswuFAk5NzAe1BxQ6cJCzVbTrdCp
AW5XUuLC/tHGSyYU/GKm3Oy3S28OOnRNRdpwPhxJUwhgou09hPbcgZY3sOgaxtTn
njtr3oI/nuWayTsMjbVlBtUFmzm8UBkoLEAZQwSM7KPTsJyfqGUVijwVvS65gMmE
mA1HNHE57kYEEhf/iRQm0eCsR2U69046e1gvJZKwbcI7HljnlCcI+YGUIISPNyyo
a5sPJjRm9OnHJPnJgZvH/KPwEgo7aaluLIo2CjFXbKu9QeGFhPcqSjHOt4EZ5SKk
l87ULIY2Nky3V7sH6kYUm1EipVMAYi/PffrU3r15m1vKD65blaB/zx7a+B4CGfV5
P2+sPI1BAaQk5Ky62g8UcKMKrPL+44vKtBsZiUWFKDs7GLtVjw5IZQfnMUbKlJNJ
2FfpNtTDjoEiZZPeH/Rqx7KAtLoqxvoV62+PZV9gXK4Yuv6GK3xUnyYXku7gme/L
7P74W7kKx760XMyy8SZZV2kf2VgakC9JxccsavrvTZBiitraFZReRqrRBkO7eZ00
tXLW+YljrkL4L2MsYALlh9qayvCu3Jask3NrmnEgXU0akx1GLJyNe1xnfNt3z02I
/MV87zUjtXAyUFyo/ZdiSZySuLKKOuWm93jHwfsb1zzKhIiD2oiq7it/m5sq8Aab
BkSJ3P6m9Dlb3AvDbp+ofrNwCajNcp7oyNGWlH5d8gXxikJ9YtRIo0i3kBkzlwJf
cUknwhmN43C5jcSTrNF4bd6UyO4j/+Qx01ahOttDy3o4f1/ygMIBrwmg7AySKAwt
PAy6pYaPPGzfejHVg5NCZnc1QBDsfztncurSs2EHNFF01PZVR9dQdTm2tyZZgABA
49YVbU9Rut3E3W1BJlwxlCUHOu0Ou43yk8KJQr9ucFlLiV2Yt8DFQOjSLL2fyqc2
XR+3x2W5fwF8eTuZHYCwoQdqa3u6FDWlp9EzhDDz4dTjvz7S/cLMjCUVmtJ8otwG
Kps0X5KbPXJPBPs486n0Ipiv2TYafZ8MAd+zpmx84Apb1Ifaa8C9UL1bBFt0sgk5
1Jp9tcGJbuUXg5qpP8Y10ASqaMCV6P9hAgXVuNl/fv0oWAka5F2UHjvPQB3vz6Wh
pzzMi3Q0Ag7wqCI+7IBWNFogGT1LRBpsDY61/0mAk64NR0G4XxzWfG6JY+P4uAkE
NRYbjXEn9YNfn54j4ZVsxgn4kzittBMHbUnZU/MLtcAXSBKDVuivZs6f9S+k6p6e
4jaROEJfX4P3yxikhRfwPbYypgiAN0O3FuWxhV8el0E852JNb78qlyX8wzM6u0hc
NVnY1B3T+l0DJf/5ritbUjiiV8jve3rX8/qEZANNLLMfLhF7TirKRfX7l7+i0y5a
bHqdgLnx+nczjQLl8KI9tgs5Q0N/aODoFMPMylHXrcHs9BPj7OYABSw3a/kO4n5E
L5nRLqLFHe6ns2vJW7FNqASZt92BWwrTfkkMNQdk5tFtImyJW2H0NA2bbXefyEgl
RpeXXUixjy2W69RZJ/N76fdxe597L+l7AV0DfLCOQ1vNSMOdjQq2xhMUqwcpJcz3
lJitT5yTP32hSNbsYZ7mXMXNp4skAfAMIJz1togRQWZusUMGkeO5Vrtupc37+T1/
XhuMUC6HFfxE9wCxZr4eud8UTRnowc+ERtEvELOed2xBiRAKfR8OdJkN/pkOFQ10
Ru2jh3bsDUTiQ2rgnpiyg27lfv1Td/BwsIk4TtcOzhr6w7lxMu+9+whtsUSQvNNC
X6DBqZbU2x4yBhK2DgIrscBHfO/A/warkelkrYfxks/us7B2+qGKevi3CY9Drcky
jVyI+6eOd46vhtdl757Qzh0bmE+YH5lRiueJ408y7aoLoAJyQePO2NwWYMcK4qXs
Nu4GJo1bnrLwpEo6kp8ZLxp6oNLC1dBun2m/DZzbeARDs2as4G+n9b0Ola5FpV6+
AbjxEyjG/XaostogwcqzuBLWhpZij5aSKz+e0lk+40QWQgeGDLNsJ3V9DCbASR6Q
OCE0Xyt39hrpGOCmauztuVSQGm3qQqH+7+iglBkMxVCwAGeeOjojQqDEKJMpjr8M
wsUnXi9f9x8xAhsoNyaQyvSIGgS7Xr6EG3DV5e3j5xqzRbnqvLkkGOa/K7r5/dSs
x7MWPiSmb0RuogUxuHHLHyNfHlprEs+iU8ZN+LC2CtF2exUPVk4XtoJCXs3NMqXR
3XgVOU2hYPlRjJzUa9PBPageITCiw3ZYDPW3sdNrHN8o/0KLtLmZoRcBfCPfTvc7
3waupSRZ2ojhYXf2us8fqGzMEGiVa2O9admYKtBihK5Y5z03ViYUsLR7+9RSzx7K
Rcd5D7GMOEeLJxXDjEbZ/vly4BJvQ4pvKmYNtbVuChm7ZjH6hwBpsWnUDoab6AlL
Vp8nZjVslr1S9SQxj9Puu0CkEdcVS1GHs1VHbVVZHSOGlpVaO4F0TtU/zjSm+awU
qPIMVG1AYPHHK/K/DLfzGiiHTbXttpZ3d+/Lg/MYAPi7Ba7vDbM6gmOxXpve9+Jk
oVNKcQzxZx+z6fPlp2bH/BxCvGAaa7v2rnj5ANgK/mwK0R6pqcVsAzC9NVD1wCTS
CxvV1kPIYNsdHlT11C2hvG7XdUAdA5mBRuXAYJ33L9MnLr25T9fvaw2rKvKv0LRX
U4MWLAJ+ovGdDzTuPgHgxgmJ7HlLh1DD9RQNC3SxY44zqt5SKI5tihK2/X9xOykD
Qc0Kck4AJzsfmRMQiRn4UhM3lcF/w8AQseMgAA1hMIGA/gQmpCgi3VDFV92MLo4b
BbMen8ZsE2Lt6QVPUytruaWFc5EgZzsNCJDa5+yKaWDXLQh6ztqB9HAwRB+CR2lW
ynXsytvqbbsfNJFc9xaqjpr1LmvpB0V+lbMNxPwDjk1dbGhseH1a0C57hA+oXTl2
B5P6HP3S4GjgxKjGJZYdgYvYQ4lKu8FhsUkjLAUac0cN4ANKXF0xvOMvS30uJIxt
kqP9eM8hLrWus+fTAN7PUkWYvZNpMMLpfLrQI66tZQOHQYOQef2ZO40JRJ6nhXwQ
WBnCP16bE1DO+DHPoOp9KaXtg4MNQNMROlE3Uc7na72emcG/mRAO93slIXFILla0
EnWs1d+2+zciHszi85rKxh4lASWkzW9qp3aARtSxU5MeEKRE9qFHOs6+vFjqPl6e
K/AYYkpQPB3qX+xVfE9njEkpia5PziWK761pC9s2Y1a6iKWpyuR5MYX6neoBUez6
UMLx4mkotana4ykaTqRar/Lb/iUeMEXuU+j+bnQDo/BLEvUUAfdu4WI7mByIzuof
ZZ8qmMZMKdy2tWvJWYosXi0M/WDweRAzhnRKut7ZbP9JSbQKzNfEt8X5K+a/Grsq
NlGEpF1TlS2ggVA0ypXXCMUo2xhlsdRj6uKgGH07FyGQOU79lwGdphWUOW1GGIKQ
UPRosTP3YyRyGNeBAGYlvMTKg90rwbWmoY1WEr3x0mA//ohK05pAUXL4KwNwUFj9
8AtDmvka1qNySJ+3qRxh0XReACxcfhvF50nI79Bsd5NWydZ9Bx7FQvinIlvolcJf
fKK6iOr0h74cDaJVLdJWSpyujdwGVZYGfTta8GbEtPAIPNjtpytYW50Sf28XFjmi
TTfzisqs4FOaSQ8YfX7oicCmnG9z8h2xuiRAGD9EFMOTmsMkaEisnUHHpeWY+5a3
8+6mJoNVpWDHXjoOAnFdFTb8M+d/j97qXllGqlS1XAlvWrFIE4csXpzBnZrMTEyN
qVR/39FD/6iY9AKPvTsI+4hvepkSPplstKiO+dQYommrtQYdjNzrKSsqD1y1aqLP
OPhoC3Lbbua35aVsertR4x/2MGvEGrB5jOYIpwcAmhVgF1NWvSChT5ultWwEvaAc
SBaspdkX8BGKFEjd6VTbwH/pEjmlI4+h5TqJu+sb1POPIqGq7R9nq3DBt6tAgZOo
/KpntPpbNGSY1b0yrDRc+QzNiRupeU/LXNu0xfBSLTfsObQ5NDg9HXOV7pcOzxvH
65JkSXaXSZrPq7dLRITMYt1sxrxPtjmxDxMXeRwBaq31hbTnILUZY4dWxsxvqQqK
36OeRQ5YfvDDuCtDfFrvq9Kg0Gh+KLFSRSu5jvbIV8OqyDUF/a5Y99Rdt7PzEF7c
39y8fMM5ynq4+QSOU0Yfr1qVEKflkFiSiVkPh/3xV8fvxDYLSww9oWT3MaNPYuWj
PDFALT7idoTLXWQ8CllwnS9IEGfjNY2iLWWzbP8M+P1/5XNDg9wUp+o7uuXbCtRc
jPmKGICFnHK89BDOgzvmfbmd4v55FcOy0EoZ3Fi/94l0G9033MX1i3eQNYUqjgwh
z7O30qQUN+76soE1T4V8Cma8FGg2nHw5KTAxkJpNkq5p8cht6RZXO977CHcj0gxJ
G+UcHTIQMYtRc9US7Nld/+9iNjEJ0VChtfSj+IXpuGskZn0FPH9QFp/WHqBqVtle
k7CJ2djrgCPEsUTEf8mSmIffVn3sP5eiOwYsoeVAqb/Cu0jzAHx6wJu6xK6UbOCu
HYRf4eLF9rNGOaAmiVuD5YZJn25tDdMthiyUg7SdR3Z06+nnkxB3Uv/oL2A5fOXW
GvDX2uy5XuG/c42mmyc5u+9tB5P3fINdi4uK9bHKFvowPL7XvcWVyLFZbTBYj61P
lzVSdYh8h7HK5nOlVDq6973kI9DMNchsvJdKTcL217eOUhHCuk8lh0xg3RfIv6wo
gA5SCifXUbXTmMYjqp5cqE6Mg052S3bgP3d3xIiUiWmebGUUBji6/HljMtV144Iz
ySZJiShavKI7QdAJWsDmRe2sIZ7qm0vM09q0WbNrKsbgJxAkFpXQs3BZP+KXEIdo
x7o1IVpM3NtkaahtXGsELURvcSXs4kwt7kdlbu1e8OC1Ck1ibrljTPg+ry/MDYpe
faijFyKqZoQI41+IjWgpOWz9cho2y8vxU3itDGgna+DLuNRjtMgjiKFv/vHS38lw
g4X4rRgzHPZ/qIKngDIRgvYERgr65X3YScHt1gYJk4BQfp5vO5J3GaD6j2yCObWc
nm3U6KLfSf57r59poOGwlBaulVNirBljxBqmsHBRijYwe/BQWtqPKTimk/jdnSP7
gOVvkVIuDJ+BJBL5jAbt1JOSBRxc0zr88Ern+A/nmeLejZAk6QkQU4BGE3q0ZhhV
WWyDmAZzY1aAe8uKAhNsGdIcYjWY5dgT0pw+MdXs0Yt69fGzAMPdO2ZC+VesID+z
pIfbPSiHCqbWo7l1d1acFSQtzS7dAz/DqeeO2uID0boQwmxXpRzeFlisQOxn5ETC
513fxHKUgNIIKxoeRagFXmaFPgSjQ2KqWJFUCuJgdbSjNwBwF2m45SZQh9HLqaV8
a3VNo7CuaCIcfXmEiv9JaRzEGJPa8AoAsCCgw+UrpZTDldy0raXzNSXFCQQ2Uzsv
J1Cx9ML8uDMGewJWG7Ktv0M1aBtGoams6RJLU2YxcAaEm+5bKOKzE08n6MXF/AUq
GWQj3MIJFi7GawshnYawOa7mp59iT4wdVBiYUKMZuLSoUnu69BTjJ0pkn2tD23HI
KcLE+pCp9RIxb36eNLA2Id+7rZW9x6mxsx+yM6CStmUzJfBVpO4FA6JAafA1hh2h
Wv02BUr6YO5i5nPsCZBs1tZG0yAtvWjyBjGIWIk0MMxnp/UHd+egL+WmvJWoAcBu
+ve5Cx4G8kER5cdXFGWjFIE6U8ior0peVTzXsmewNY4jgipVmbrIOh6EBhA4LPko
qUhz2SuhhjaqoQTjGWmsgXpaf2Mn2JBLH/JnHdGVgjfun7XW4ju4HuV86t46xGKd
4wxrlRHAU+MWJI9izpMskYZ0Fv932FVuW0Z6zI/MTHyjQTL0I9QVvldHMh2DPH5Y
v4EyHu5zpkU3d5bV0jK4AQ1rr1X9NlwodN2sX3dnI+ifK5pQL6xn1/4PXMw+77tM
rYFxPGiezWk3nmoUPdMKODXcX+38yCAMxNMA7wD9P52lJr2egkqUob+5/HXoX1jT
HWB46/kkIEMDN4S9usTim6m7pqv+GJ7KfWWBkpeEhZutaU5jeqUOdmIBvwoPk0FZ
Sik94FBNwgryfappaS3sLved8ygH8GlzB422AnKPK/Pek0uUpRedTB/51tF8gG0k
CPvGlEIGVjTxPMzmuHOhsfUXpx1ry53UmWFTGG46LhWboek7SUo2f7sHTlBzP1V7
5jac7WnLcsUacQQVIQ6ayCoeC1ApMq+/l3dh33V3Z5798rwWEuG1g7Rc/D09IW81
Hvj2HU9Iy6U9D/Cb+9/ZyCwNSSdJ7hawTxG9TpaxCktFnBSJvG4p+Yf7ALFAOBvg
XChdKvr2zUmzda2NuFT8IfT/y3LZF32OJzN5f3S+E6JRtrukQCWiNj4gY4mJNp5Y
j3Elhmk/DvyB8JS2Lvq0sx7UokEplsvnkLPd9DDG1pStkPa71qkM0APh4m7IuS1O
4cFibsg1BurFmmIp57JAayLRNCsZWTL81O6rOemQ5OJFd4qGDpNGMNROnvoWe/tD
OCXxr0KHQE8NVV2nPa2X2/HAxHjvtNX1m8WAkSm7szv2OLA7UUwCctSXcaPeMcek
75vVnAJHnY5VI1UeCxX182yV+d94CO8R5prVPJL9FOZEFe3qVCkHjeWgtTlyzTGK
LT7TMAgsQvPuJq9exNpuWD6gmek1NACqQRKY0ttCP7+zkSP4Nuvzio77YHgQYN9/
pztHJ/wrMbpxil44hq15ZdS0pV7xOX8t/MnE87k/LvrhuJVKB19DlFUGcljPgYFK
GsZYVXWCyqjArl5h5sf4/WoPhc0uy6typDPO1zfk0PAKNzSE234YOZyd7dOY076W
mU3tVJ36OBpUCx4YnYG8sG9M/9lK9aoD4kkiiNSyyZlleDR6wMhId+wKUqm5zOyc
6mHqKlBCeALliLh/+rZKzRJiUE5XeOoe0uu3+txsGBwRJfMAEireRwsoFBJDNqDv
aZ0yyhDp71EEC1e1XLh8/rkEukYDGbBG1oQsc1NVH2ucENHn4QNiSga6Ho4EA5Sb
f1noXHwPCmr/lZ6iZHQqxVvko+j/AvCNELfEeTvHuAPzcsVxOXe8eqw6ZBT43SMb
ZNXzatP/NWR4jbIUirp+ccWKnloHENBoVX6DWfYK5aAOo2g93A5JWMnGFNBk7a5w
z5OJn0yausvCpWkJFmWxj7haorT5GaNGWhyynsGrNHtlX3g2G0P8GqgjF8Alnbdn
JJrNChSm0zmGN3UEDJUm4KK+ifEMICq1cL4fQEyjRh72nqqLPfVHE0Cbdjdv/sSf
Zoh2xaUG1BF2g7HMglVr78XmRWvwomrWFhCvfBAkN0tZC072o70Ep+eRXdY07/A4
+CxV4nfFvlk5Fif33uo3Qb0sotH1gGdkec3eLhng6Y95d3j3d5lV8mYs/gyGX1wj
reCXNnbEaTzTcni7Np3HtDu9+fhw7qwT81UkG8YdJBtq36IdZ4e6en+vXzsy0GBH
9OvNoAph/R5T80ZYSgBVLqqAQG35rKVA23sRAkrs18Y8qCDr7wNRpTCNyBoTzS4T
Un3Vl4rWFmo//hPaeAlz0PPOXZ22M6n8wA5leKuSGMY5dCcbWTHEB7XB487FGG+N
93iqP1Ueyew0TZPvuVrGmnGZq5F/vAr5FFKVZhcQmdYFgRAPiL5nYKHIYX8FzbIP
DXWeaJz5eesJF6VIq9dVyJAlrjmF/3p0ciArpzr9ofWgSYh+11Jv9ODvZ1rDlXVm
FA+ruLgrz//nZOOPLXvkFlZ5XY+l7CII3ihoVF8kp6lThVzbR2ekKlxg6FAQpOdn
ySP2GqFpQKFYkIvOvEu9Kwdas76hVqY2DHdHgAtt+QuCbsxUl/8ijlgBMPhhuEES
Wcg4+7EA5EMg468Ve5raZhYif38KaVbVveJqImC8f+uOZNo5ITv2hhjEa5IrjQPB
ikPT/R8QtRGoG9Rcjyus8QwSoZp7Wp2YGlKfg6B/9jWtNFSdfTxllojO7Ip6dnIr
OysNs8QQJ9HZA351smFV9jZTCbNMVaVr+MyrMhAsWjic7HkQhpp4GxeiJ9WdlqCX
xpdb+K1eS4twkur6NkzNEC+Ib6bk0hY5YQxLDMZ0bG5+BzRUecfQQPmhqX0KOpzn
y+hTsJucwg+POZHYUXUeETptaw7BmNEKzsud4Yw8L+jk+ZXAGdzbyp8IyEI4vIFM
7jX5AypsSXDXLBdn009/5BiSl/EP399ZKjqiQ8r6DpVJZIQOTbeejo9T/58xwZSP
kB5ifVN04iKASwAvjW1QX1QWyntb/+L4cYr+7WXwOml5IKuTzoUJcahDl5RuL63Q
ue0uYlOVxQ/JsH1JY6p7MYP9UFkiaKaDk9N8oFsyKDVJJ1qYnxXH9VSfdbq+xgWf
67tfNbhf67ujMxJVV1ymlPHBe8lpM0bDnYX4Ul5DIwJadV/iYZKhI+lYY1FZwFku
LjZY8bVO8JfAjN/XVKayh5WEInW0g5J7w8fl1Gj9zFVzcJzOOLITblLIKYkQI/dH
OrO6iUsguYx0dgF2MHrPjoXQBXFByb2ABfAfHIZXwBZ6tTmerHCh4M9Or/sje/hY
Hwqqq5CHYGxXzyxhhbC44FZtVovLX8jLv5k2QuSf8x1iEZWqqOKp+3SPKztSHNM/
HhuTg4HWAO1M4IiIQZp4D5zBE/D2FVICHuOgi927GNcp/eJw1wwkO/6EBoPb6Jh/
v4UOpL9PVvwXPbvVWzMXfuJUKG0LP91HYBFDhskS99GdTUiFiKmDO2kjHhkKU3Dj
jjxrHOj3KB7cF6PpYs/TVaxPlsI0hEHQyhHI+k7hpRAVsByUClPUSBJCTXayLcrv
CtUS0r8vm6IOs/xZcafpWMmfC9dePklgnFEpcul31Obq/+uvvxV4/fTgekZpS6/7
LIkEmBStk3wHqzJEtw01u8Kdrv/JBQPQPb+qZEVc53/buPhfTOsqkOdajL2i9A6D
1sz0gcVzunRqdDjAGGFEU02TJsp/S/FU8Pl4U/Nb9o/XfjKuE6VRuwPiKy2Z6ewU
rf8JBsA5VAj9+IvA98zrWfECHipL+ZjS5aE/GXHoCEnE8MLQVrYqG78Qad4W9WIR
eXb+opAUOAAqyPkL9D+PheuPnF3XiZ+dVDWquUQ9ZT7IL1I6Eu2jgI0jQjrKvQyI
s6NxNZbsrolk8HiK9pN4B+88ZTIQ8Aa/AH7Ti2kqLabUrFVMfa7+pnIBmm08b/fM
6dyGk8XQrslFRdi1MI1M3vINjeEUmPlqDAXg/0QQgXEuoA+iSNP0F/3Ky/Po3zhZ
Wz+AIZu2m+ZMotVrSoD4X+MJKz5YNrl1ic5TvNldqgo9FyIVnhsPHOQeFJA5TdaM
4+2Mytp35grXf2yiKR0/2J6ccfQPvjeoyzPjS16h5BP53CUyNV8NaUK+gJ2czWrE
2VhdhA8cgP6dwvlJLyPrWxQijXrtRoqKhMfjtsLtrKZV+/XOLqLQJv8Zu7WmNhnj
DgZB31eovBynIxZCAWW/IYMngDPfL3MG+w2r3f5KcgJrfmOOMuUt0XxuYTqmJN+p
wqP56zKNc6x/Mp6mphRnZBtvSPLTLBjO4jz8C/EkeEWcpYooBX3rgDB05tXFXbxP
BcF4M2DYNaDmwUbuUyV/TRt1yGG+84yPOyhdJ2kHUKlY7+SJsEfgMCwrM1b2v0yJ
0oSTGJJDbJ2Qn0j8tPJN2GcBQ3ObckgzfVgVPmFj5TYKXhF0T3Y9KVnn7wS7oF9u
tzW/ytHvXjVge6AMQcrPZ8Zqz9fwNQKQ3WMpEKyTeLniSMky8fVCPxEePhavyA9q
DnNA3So9LmzDPMvbnoLCuvo+1GUPeTrtnjcQwR7R4N3qVQ5zhaaCqlKgFDTm9g5p
SNE29LU7cpIPpsxHG/A32b74NUiNJT1gGRqZI5BqZfOvFJhI1V3l1LFMU30To6AC
b4Iu4bAjTHg4PVdiiBOWr7czVAK6yvtYdkResVM1iyVvyuOBfkKAvqrXn1Y92hWZ
gwhtnStSUnV+36plK9veMIxnB9tRIuP0PSmcgivetX3pYEZV2wdSJPGt3FPLWb+3
GNLcKPAdKShVI1gKJoqEr/G90QbFOr6QiKoxGMB4Q7sHjVeSQamlMOWngKTAE7G6
qxX9ZxIGbk5xJ5bxYXz9WDxI6u1S2jcEqdFMq0Kgxm5+nT+XBp07XLEggf3m1utY
9GryU1zIVFhFKcRVfWPqkVBjjQXq/4uHIs86oBepdgqF1/3aXgDGgWnfri1uj7EV
PEH1cq7va2Qthcwz2RrkykwFS9DkIx+JDRMNNN1Ir0ohh7rzASEm4lp/1NM0qiyP
hL/i+HFdhEhv0xHLUOd1AsLTwnuPbpFKaDspUHuZJB/5x78iIG7bmHavF2iqIFCn
rZjJ41u3sr5f2nr15Ah7aZrqL1jhHHCPnOgphHpoic0J3JVodAm3WkhAcVyPJaPz
P06Q/HomZJiKNbbU2pxWfRDNBoKpY7LpDsfIGddZiATivZInFls37V25NcLVad3y
GOabMv5waoNlDSrJ3n4weB4ceQqysnWvkavhEha+54YU3iODsuAjGQiLMzDpYH+h
DL4Dn5v0vwdOVRfUULaJVmYc4aabbRGsjo3BwmSZPorHpG+Y9k9xruBeXY0R+rEx
syj/q8cN6ZwK/bqfdIIukdcklN2pRInlkrq3vGu5cSpdoB5ZrPTyXn91A3pLjP9h
BMm4NPagbe1+isXgUfYmyZJXE5gABjpNyucsFZW4T4hZt1G1TP0WsH8dvz/XhdP/
JlJpH/N2VPg0qJQbBj6peHrrRQ1Do6ktwdSt7uWOYbCmto17cW0zl73fh1wHuDJM
MJeO2E7TMOm37T4vtTmBGOVyaP/6xPUmI2rrSGiK5xUzzBMtriHTS0K5lagLnCzX
VhBDdblC3/iZ+U26n6fJYFcNyvHSbjXhjHT4rOMJHn9JPsN126Y0slBH17KsYwLF
LuyEExqwsEky5YIIEVmJoBAUQFGqTfcxoP0aHoL6TMCHaKTmeLf0bja6npFehjT4
etJ4Tm6wmsRw0YK4Q2XdR9Vp+AugculzWF8kZ/eQIYu3qPSEMdbODJM1GCSdXdlO
PMIIPBTzhrY2HawntqFoGGdd6M4oFTrUSxK9oBGCzlmjA8fCNR+/W6XyoMiv1xrY
IzxPZ8IMzcijqSUVtL4jiEi36MPTXT6GdjynoDBF72CxkBiDngO9ATIqJSDFCd9S
wxtAipBj4rF4K/rTJBsmJSMWLh27ImdkmRtafCemCmFBiLebxrKCsDLpZD/QcND2
i2LbCP3SxnpqQ38uZ/dJ+TpZ8Dj+kDS773jhxu7QXVnUJqh6nNvVLLwD1LLKMNaw
gixTVFYkIewRma15ybXOBsIe7cqEh2sCjEKlc9A8cIyQtFf4+7lqtgVrDHIHEaLF
+uI0nmraSo8JE/eBf3MWLIyaHBaTiCx1gLKF1UjNaDEultWTj3n9r7aOGkSYudE7
QjpBAd8F1YB9+xVD5mc1UjH9s4mZbpj2XVTWz+GQ+8GyzBepMNodIS9+rCD83FDT
HlBzQLEz5HArVLuAwr3Jc1gfRx+emPxRzYnrhe+okvC5HfPA3mpFBidWxWmOZGvv
3aZtRY5OAmJPqUsz5hG1YJkKF5k2ZRLkTw0X9ehUZQFaCxVap+79DPqVoLBLYQZH
VIa8ikdBCrX4uGimQJK52VQSKorLkDiDgv1oM0TM4ZVkOcvxnnrrdcRssnw4RBYM
uZK9rmB0LmDaQL55iS+gEl3SGq7g9phe1teYX3caIMKLtCUDog2bsbUzMuR20Eu5
YpCT5M6kYj1v75nG53wb+Q==
`protect END_PROTECTED
