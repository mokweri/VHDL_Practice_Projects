`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frDLHvG3DUeQEJy9EhbLiqIDxcQcRvIaBhtV9/IahJwzTjlRLoNUDmWemmpSsjv1
+8z6tQBWnixP28w+QK1k8D0cvqL2Acy9X4vPJTWDNY6ME5NTLsxHd66XgG9sWlDK
1e68SVareRl8BhbWYRpmKP0ASet+T+7i/9cLQeGc5aHdngRflmfM84Kd/+4O78Jx
qf/UGevYV78mkZmsM/0dD4AVvqAQUaeKKb2pctOukFvuw4LBb//yjO0449NFMwk0
EhtXNXMQo8QuH7VEfxeDg3Az7XGB5r+jiothSIdPDFCMqThPOEQMco/+tFYRsslB
0iBanLyR+hLH2wRNelcW0I55Onb+W9gkIE9X54Jbs88+OFxM0FGLRnNQFepGWBA9
94aEQkctY77zHNeX2sDffU9/vJalO0KnO+tQQz54ye7fsGpjmeGZA0agB9miCJ+V
YinL3zHLNF0OwMG7Jnsnb1xhVeWSi7eE1F6XpLliKEmZBbVa69yPtF2jHaFgFO40
LP85WGiy4LJFDxa6qG8MSq/OuiIoDB5+oZvKJTUzTfI2B2TjR/ua1DjC1vZ+imd/
+DNUjPbUkRSyvSqjxuQDRmKJkzZs1nfJLWM51vKtWKG8KyMmIfbOr9Ijn+LfVsdi
ZtjHHM7M5Qa51JdhH3az0Po8inLwxjjYKaiWzgeJ34/bVsFeiLzftAIEj/+Acma1
47zy7KF2NtfJoGocTtIT/xqFNdqG7zT4UAxBUqGqoMknLgA8DIIVSKE4inbWMbsG
Se7b6uNcirKFXUcDEwZnJ84YQRF31flqDPZxvXnEDi/FlyCHVEUSNx50h/+jo5+A
2trN1qJewtAhZ0EBwB93NZvyWnuJZQSBYFRL9rc7z7KVjdPOtDjQezH7Yw59aGF5
e7ayQIeMr+mQRBOqxICczgboWsGvig1W5LZ1FPTuJ9v1NeWRjfHONsNvBywL9bun
tdMaJpylmNJGQ3NMYsDjD5g73BoXbXT5l5kJ6T5O9UAtvOQU4ssHC2RZ4eAZUILB
yMFU8B7ZUNiU23RQ1IHVajKlprqZONVJ2MP0NUoBVpD3FswqClS9VVzD1k29kRvm
kMbQHgX/ytW9DSowWPYNncTOPVbJdkai1y/GEtFcSA5WC9JCLgLqrxZMoaRV9ouV
GGXulDwf+7Mge6K1iJ5VKWdAfCoiEaLp6r5mEo0z1TFudT9I5lDxxOgSaJA9/ivy
KVuz5CgGzm+E144QVN0yMGPjV6ZSaUW8ghrSQj6ZDEnWl75gT3W5CwYyJUUTHzlR
iOCxodXjjy41f3b+qRREJoVVhApeWQaq+eG6n8XxlxdJXP7BF7Wqh7R/rfbpbT6b
gilWlJ12O8EL9PrtpgKkt61V6IJRVFa7o7Wct6/NXi+HLjumXapOj6lmcBQM1JMK
fNH5438TMyq8Aae351bvwISwWzl/TbUTt9vcqgamEIDvv1gmnDthoBUlKo2GV7iW
pu+XWm9w8FP0ZiMZJhIvliAhg8vEmP2VwBsW6C4iJJ05WFtnAPoq4276Tq6XZYxe
sRUpfx/Hvn5kkgnBfbi8VrhP9VE6NeY73IhkmvaMUygkOLjsScdV4pZdbsk9SQaW
oF/2NjDMCdjIdbDQp/rNlxvYaNHfSvlnrZAKIVJnpOwaPxgSxxEgweoe1Jt6HUut
ahcoxuktXm/YMYwEVYu6hDcmxUHvyKbX8QvADoFpaKjzkRIh/3Q8BjNh5hsq45FI
7QPr0Uz5eiFQ2dPfrhdzrQHuAzRUhSEgN53hEriBx3W+A0CpnbS+RCYq6n+dY8Gw
gxSDgFTIOGj5O0FMMLFLX3ylmOq5kdzqPfpZuGd5pA+0NrCEvwljGQkJlFea2YB/
CAo4IMdntRpye1VMNCGTUxwJeCz6fTSOUge0MDjHC44SkrBqBRYBFtPN4HQQYkNf
A+kUC7zIsMO4t3+XsEm05B0RnV3rFtgA0+R1NJve4rBU/4M9h1R2lIDi7BOssqK9
HcUeC//+DRnRx0vCNA6Mo+6tRPT3BMWbNMnA0Cxq4/Q3y+f5ERgvGU2T1kW1c6Sj
Y7M7U3Bd+15WklXGok1G3ETPPxcVuytkCuhh2qOGC7UlaM1cSVXl3kGjd+vvq7l/
0ANgGFh4rX6/mk/T4Fn2SUFPrFFUuXgMc38jENVfv5HtBIoQRUa9ahACAVKPoxz4
z4p6oMYnksCm7sYffcWBtGDqkudU06ua7DIAYC4aGwzHILzmKPu+IGkeMt2ATavu
inQC6ORGfm3f0xtH/mvYagikBxTcwlJS6QuWiy3JxCfw4u4KOVHX2mPzHbUzdT06
PO8xItPsB28diQAq99WN6uDCdSzJcwB8IKoCZ6AFWJuUqM5+BuZXaSQk4ZjSsZpj
IFHQOeVP4fgv5fviNnZqYSXOH2c1rD1KInMtG0FxipWanzx0KdXzRFwtja87SI8X
pmrLV5uop7uePobgkAXW2ps6h3ZftGmFigkgJdDUQbddXb9W8gvHyk4QaS7ZohdY
79ZtptddVce6PgVsy2ULSD76Jw71eR5cqV29pFdyBXASxjW8s/jPaOp2pIjHpT9h
s4srYQSrzAOQ5p0WkJdqew4fzilDzJQ6B2FEllibpLvNuvRgiSZE28btDojTQHGA
Zo3PiZIHpoDxc9ExiynUEDnooC399lIJW2gFfu6f3VVim5Tj1nggomUVgre24vhl
eA2ZKVyKLsnVJUW6ZfZEP+3vM+zdmkA2UcSV3pBf6xvz/yySD2UyUzt4tSfmyhnN
jClCFwO8a8IdCEw/l+wmtsMDjssEBOb+CrnK3v7yC7rQvYIFyzCNKTwyLp+ZfbRo
JBvEuIrMLS4Q96blXj2IRUCUNVwl4gdEAOve1LatJoVAny0vUpjhKU1FYWU/We3+
rEvWZiiKbpGl0ZHdBxMsgHtckFuBdEMOiDeDs4beYs6DtkTG1ExtVj/lOmA2haDI
WGbO3akQ89EjZPirL9JWOvml13dfZXCVxST5alsdScOXtTLfwCgG721WDbbMsBo8
wfMPPoOAeOGc1l6V53A1m5kZUxGPTa9fU/mK6LbeCp53uS8UflUnUub6PZHTSFPL
hjBabqcslyotAuUra2MjEvuWtLSW6qooax+Xd8Clk8MeTtYffYIZ2LDtbdHGRl0B
fJDzA7MERjm+SKo14jd4vHuTefnIO5Jrn0Hmpj3DH0LtmXv2pS87RO60AB+MruOO
QUYAhcNB3v5yS//+ut48pk5SvTv0KhEYTLV7U79n8acXdVoepLp9ezVkP3aGXEMX
HWP3TNJW6IxxkEZ5qU8qrRyoBB5XHMaIrIzb3x9fmEG5yTqSoy1LjvHSvIODqJli
uaPxWvH6ftpQyuH7SvpcQLp+l4jyxUUxzZOoJOWxt1jJw30uizU/3B/UJC5Mrqt2
mUxIPEdtjkUDXD1o6FWeVUftTKvIjeWXcrUhm5Xp9dMhVdI0E97Vlruo8SiydT91
s5SYzSbiCTzQ7TSDjyliIs7W67eOXswIPH52VE7Cx64B2XdHbfOb5+seddyYw84a
JGOkqH8xOSdqpzFF5JTb3tphX0fZicQHdU6MiOOrKeXk9qSi1/IyEBIl83L3mUmH
aNVEjZpUzjZtjat0+3CtYp6iCtayghyVj1GXTtl5Q00HsrnUbXhwiHikXAkkUOq3
PgvQJthwUSrIh8Piab1WkRAfQRdrjD7V/KHeIPxTQIfedOQwKw1QFN6Mm4c/ldBU
O/fR5xCe9NeqAqSmbgkxE9bPb3+MCLQTURB5IgKqHgxijOMjeZh4Jm2dCNOPlQvr
vc734uqeeiP/tm+eXdeZ8cT+nxmmzD9J5HpLF81xhAIgjH+lmMjesmSaROaBXev4
IF3I1C6WcJuKXngHZplJteU4KIlJ4THfcIpzDZQMdKfsnVIOdGfolLy/Wgmazc4U
Niu4BlOP4mrrpPc2WHqvOE2VoACJmaECxvUYW6giZh6Jil1eLFpr2j8HB6s46VMB
UkGbdtnaWFvwe9zvjFjbjKOefSEivCItO85NrGJOAzqEJHCoE20Y1kwQ3RtZojEz
hUu1RMkpFleVjz3Q+c349UgUDP7Tlju5KzFCzXwox996084lM1iaHgB5hwFVfzCQ
Yg2LhQXUhsn0FFw0Ln6BxSGE+hLTDfqr+yB51EejJBLZrSk/NPpZ+EZALRcHEC1T
9e3A405+rNfnWs98rSkCbXg2x/w4BKD21pEQBfrRm/AV2c7CZgCj7qUR8c8bEKaG
KGKv4isHAUJ4MCti6mpt8Ac3zkym3LrDsBdvSYTGziJhOoP2EiyYSeTsfhylRYFu
0xuqb1+UTGUwYno8ENeEQAmnLyMfNKyil1DsdVjVJll8Olaqi470+jnV8DTw7Aci
XbelLUkLSYm6aGjNrPl+vw9WdnHh2WqMmmKwq2Vh9Co=
`protect END_PROTECTED
