`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y/FJ9HhzrPH+wCgqPgNPgWT42OqzrBRqxoQZsFsy+Er04tCvuZAGOO9yPP+doSwF
eveH2G9qquvnRPNaMHpPDUWNXEBlhKMQY4qCyDeOmMWiphDPgNa4RRwqTM/4DwUL
rabrPEJZtgxr8cg9lVZSX3hV0B/ybGtkn1drW03BdGKuvaqG2+R8f4HtIWFxFmdy
cjRYMJmuojviqqWhaUCGaNF3UN+djtPGGItCu2L4doEyxWHhYn+35LG+iW+XF5nK
2FDqUN5/zoTMr9ZXJird9SB8iolcR3wkx+xtOxvJhhQioEaEvUxOoFlfWta08t8M
gH//u63vLSKO8oOEm+dXGYrI4pu4gB/suymuTt5S/kUILcZHcBT2wxTD/t/FagjV
34f0f947uWelbPVazwrdyPi1WDM26EKRi247rmavxQRMGZZiKmzjw4OKphL81sn+
+W3ReECbICHnrk5/Cr3WnTpEUGO59/BfZo1oBZLOCAjQChb2ROU2q8a6jMQI3kqu
GJ/t5gHe7WIsLTs96T31jk3XB41gSjndRqNRbT8Jcpn/ejL+bclsQVAbtkEXL2HU
jv2vuuENdckNsBifqUXnmWSuMd53L3xPGCMjWeLTnhARIdjgg9kQSTaBHB1cV+24
vZBCQ+T7eCT7MdOxxOs51YRB+HJCAFGuVjXHsHLgOQLjvpYYBI5SIDuibd5/HGqv
FN58MIcawofIisi2T0thS61Eowfqmu/1O716g/tpr8+NFz6V0WpczzE9fFpSyewo
3kvsgG8BVhGxGLPU7DWTxZS/Aw6DQOAJq/QJ1lQ0YMX94Ns9C6p3dlstw/tjB1GP
r6dSQDb88L8Bj/sPofQkmSIMJv0Oq7KLv+JyLxpYBpRmZ8ZoqpSR8VO59YVT+kHJ
JWa9D/M9tdpMu2eODRNM1jNo0CZgSM7DwCWgHYapS6YV+RPZuP6NOCVvENrPkU2d
/XCN/pWgRzcK0XlkKfx0acLzW3GUNDq/Hb1fGw/23jpN9Tl5ILkLHQIrLuP8maY/
Ee09jD0mjorlvJjEOzRgSjqjxpYZKZ4cYAfZ7+qu11XrGeDE594de6P1plWkx8cg
hF0BI1WVj1dNC5L0wRrxASb0IYiH+uQbqfrsbt7lTAolkNQckq1bKtKacJof85X4
qYBRV1ODTtjI1XgvxXz/QThJEW9ppNsldU2OEtIsvpUNyK1X3VgKXbGD2H4UynqY
fGYxTZHlviviyo3CnVGXYd2NqRlRQOJwfI9UH8eFJSfQ+mio7EzLUGfAH7smRN3x
+OleI36fgwbsNUVhtlygbnLyNv5hk5KVCp5/uum7wFBcwabM0uU16eSzjT09fLO9
Z1v8I7i8C4/h3OV1UrMIxbIjOb2K+Q//rd0/v3JVElLozyNtl/rYiqLjnfplkQ4Y
SG/Boan2QhdsKW7qgHBspvQdXdfqL4DZlzpMrmk85LCTQxHCtJvibOyby2MolgIe
SWRlzY+7cKYTRttzbR1J+aT++MYRmUDfVkCl3PXebwJQVjVKApgVCUHIVLLc3WkG
xlhwOpWahZD+duKr6SaAZVaz89dA0QxZUrJlrMhSm5N/fYiOrehnXQQFc2vtgONm
`protect END_PROTECTED
