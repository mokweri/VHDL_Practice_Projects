`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+a7cXQ9rKysF3bwlTbeNgTPw6yTGnPP0O2g+QrlrIPT4TwKXHnBIw1lFWgrb/Vp
fukmSQaSupnKMRGjZXkzHn/dDccJKDMcv0vs0R1Yzl57yx2lWEkwwoJRwDEU5dCF
CxEgJ0ZyYnHq1peEHTxfwhU2kA7WwavWQ9MCWEyeX5WR0yiwDiGvvO6YhoSGLmgy
Kk4iCbj7FkBL0kHDDqzetFoKfDAlrn7V1X1spJnNSIL1G3G/PhBqXv8PfJdbfhSs
yiOcOzq6OdPv68Dlbu8pXVco6xF9TDcY7QPkJR3S9r0/UE3KAVhqsMNfqYKCG7/C
y7gVS1Fz/I6Y+hibSjQqJ0uX36H9tTV8lcXpPrvpIByEv7uzxdfeh4W4bKNY/ZRF
AEJvrcHOeCnpyLJ2236v1HM3BFtpfzakDYRrVAXqasBgBQCjfJlFALyM1UvZdwSP
PPtly117nV1rJi3rIJ2ztPV7ddHS2I30F0Cd5RWPLM6UZanD8e5INXxk6bd+Ys8h
zpdjYWXWHDLItQMlo8bSwdeE5F/X6IThvQ7XA1bt9nfy5/wLy/+/vUVJ5QffqSuP
Spd40mV+TbSh6ztH4rbRzQ9sCh3J9ZeEBTDlwzE+ZVPb6z408A4ph/WaVeZ9E552
kazVXKg0S96pC27IpBi/8Ryd7mAc7yHSmRBaolgpyUihLvSH5c/oNZu4yAxP4bQv
TxTPetWnwA6Gkyk4To1XbcO2gvKAMIC5tRWLmx1D62WWcrQ889qnVxxzcmOEjZqD
vAa1HcYp8ASplyVHfWK8zygw5UqKEXQeZz/1OzLb4/xmospgHlHYfSPlwY+4pntO
RtAWLBBJvrNGH3Hmo3rkPeMHvSa7trXKHkNZv3IQRzPB3E1fphdS0ul8XnjyX/gy
gdtiOsd/FKqE2he7y0Rr7v7lCyi3wROa+Y3QhyPEDtGayPpaIopmIPQOY/YzbrVf
ffaJHhas8gXzBblttuj3EdjBhXzX15RoPRcQQrbqRNMy6dDyI8UVBKe30PBiUGBe
kLMdaYp4KSSJgPbnp0VdsqNb2JBufRszqDCOQPJAMb2ossIhE+jX78T5GZ3QdwmD
lLVkxJCejhB0EzlXNXlImUv2R5uS3ihzJ6+5nqgDPJ/u5KjEkLh9+yG3ZoFu+61v
hPsh7paDvw2FF3PFmvdIoiOdkSuNkij0NkTDrlVdPZRQoY6yj0LXDM/c/T8RfNX2
W0r6Ey+T2V55JplGaZ3ACeq830qmIy9V+a1RyUU2X9upn1TbqAIt17ZwU/aklZTy
sGC9mewZu5zxwnhfXcFirv+uaCgcKTtDjWAyBvyct2q90m/4tYeY/o0QPge2QKSs
b5925QVb6cbt6Y8xyMkiljuzfcqIVrLruMW347M5RzAlYQAxO46/owuacA5It5eR
s1w6s93QFimnfGynbVg6/LjjS9KdeZRc6gtYt3QBlja/0THaehACVduoWtdDyROB
bNuzPxpDKpD49xvn4cqyDucZGkSJNrP949J5K4b+6kfIFw07kLxIY/4h1pkLZG2K
xvvA7dnJd4afyp0Nf2Dej7BC72vwDlT1busiBpTpejlFr4bEwjC7EvYqRUwbzlt7
Cl2YuFHUccVR/8qBd4r1w8E6tVxnIIZ4DAHnCLX8BFWfTyN6GpsDlpPMFFsHAABJ
9l8H++wt0UymbtKusTZ1kql8B4cA6NXHHZERdlBjcFVTxosjiS07Vze+Y7JUXmNY
ODsroOgK+0/LXcfCTOgFuvkw1tXcoGf5ALPRfJZPXv96XiODDu2UcJbraJ6ECBr+
1OEBXxaXeoCCZNaWB6oGccKbO70NZ63qbub3s7RDFcgxKwVNGX4W9PODR1oll0yd
09MLbNk0XsV2h8oQ+ivbtVetyocosGtgNqj/i5dQM9wfNFsd8uDxspYkW/eYx9dF
EsiVXBbMIERdmbN5IQU4nq6VZM2w+mkV1WJnZDpft2csDuDRrW9AoTpCPPTaewzQ
ibC2EzZFtA4zhjlZ4tlOZ63poeiBlGzWq3jc9Ds4A893tzItlWyYuyv+LtGq7LQn
wyhpCLGAbYJUga8R3+jRlZWtmRHVWPeXcjgVZ6buh1fhC4TkrKXokBx2rQhjNfnc
SvnSDGhSPTQfC7i0LLJVtnQ4NQFP0OMv9D2zgl6XqwU6wz6IHxHWuqNwvZmSLIIF
+tXUypZyE+ZjVReCQSFJZPe9RKTOkIIB3z3tXdxl+VORkPzxku9uj/mBiNz+bpDV
9WXJ5ZGdD3dIjQCw1p2TMFZZxx6cLEMsbqqLrbpcerEQQeLF8XQ1LFD/aWi3CeXb
W/g/bb23USAsOqBzaPNvzO6Mo76FGYCGv6KpFJtSh4E3D0Ttr2Xla1nWwSy63KMr
k2THNxpEDkOZO1FPzvrDDIYSZofwPZ6wYhXzgHAlnSjfTRtC2zv1FDX24MiQrKAL
9w7qBUJHIHiPlLlQLD82llPoseJuvoEnTAp7XrDz6lmmO2SL1wmR1mFzXlQ5t369
H2H1gp7VjQRuEYwMLu43QCmt1uSZ/8tr92seE21L2ZvlcUznSlVLJEt75xe7fwkt
NQOoBAPTbdz+X/mE0oOI0Gp8fUxxUqszOAF7iHV7EQIrzbno2fazqmFeXDBSebWL
imZ7h0YrtaCC/E/+G9HmeCaC1pf0sjv89Ys73DCRCS9zZFbgSoG/MEdFFIA+6MqQ
NMANRNz1dS4FTJvuqp+dNYG27Z1XWSKe+rLJwCjB/zzzl9h6Urvk1vU0eK8F5Gkv
2lHvhw61RFdvt+2vPCupGi2dCQN9A2e2MO1P4yv5hPRvrrSuOoxW8Aa+5kpM4FYm
7N8+lSeSeBC3eB4MgxcCPMTAP4A2yAZjV9NMSxi1g32o7aJQDV9aMRo13W7ZAnj2
TzSZnUiNKVgleva5NoN3loA4iJZ2fwhdWMUDWB4xzxqWmvm2iV8dk2RKfvQKXh2R
GeGdwOWYbCQrD/SX2HFBdvBP+W/BTWJwjnRbr8ZQlBQQPtr/ybT4y+zFLxaKtvxY
IubrVt0bBuTSWcOhNX7mtYZRH8HIH35gUhq8AZefDdab1hLRrfR/fkHsatSi2Jov
EWeHkGYIEscTGlpSzfQyZUyNrXSmP5SC3YmXXCXUjDPSPkTEyelmu+XvSQMrQaac
X6G3hCrRSBwBbTcXE2pCY/5s2SeH0D6q1/elQaKUQ7gxxZsXpxRSUthhmyxcohVo
9y03vR2Mu8PPe8yIELTPPvDDbVByFAKNZiEyPLCO0+KGA/UmKMhHrDVJW9T9DWQk
Nz5YvzXO/alFBCwy4qVVz/XSy2KHewmvyVrCSqiJfnTL8dwvR+Zna+7XncwmUwo1
/AlXSyxdoo/PvcafUU+aVb1/jnjFW62iBt/paQqgddDkRsDDLsEt1D3NbuPH6cOk
n1Lu3gZs19k2Rb9rRIG43D8DJRr1MdCJq59zEPHUq59/Wl1x+2Qez45qXbCJd6lS
E/OnZscnuSH9zP4+YfXpiqy21NJLBbac6PA1ThEDFXBcPivQAtedqyRy+hTt1VPf
GCuNFGa+9AkX4VEiu3qfe+qWcOmeluSlSQNK+sf+bYT0xNp9YIIY4cyo9hvkY/Wh
HZjtSX73DCDeQ10oUzcgaZHRxq/T31KI2MsYTouECtRlmK2jGXU2cF78GqMvb/b+
9Q3/oF62WhT/eiDuDvDQ9v/a6MWMeCcB5u92fa6TCXI=
`protect END_PROTECTED
