`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XnEIi+7VR64ce32DtHQnO8t4FbSBUxkuNz+2wiQHES9mtTG18w2/laruYtYfHDWw
TQ4Mtd1PwadOLtPdS8DeY1Jg5TZ7SZasJsIhOXIAn/bIaFZ12JP37C2J4X6jqmCX
FnxcblM11Dq/wuwG/egRWm1W2EzLSdVAWlvZ0+tL4mC9Kpd87xvOmAqh8ijgNbhK
fPdEgnuPO8D3DSFKiPPCAs1B0xaQdOwZPnqvCRL/Wl2KpTDxGqhZ07/+0BhZ8P/H
zqzW/cawePTcvMq7HqXNVCq4ofVNDd3liuP9iZ5HiVNaNVENyumvcTxm51/p9DTi
SsOS8mcgiOuIUs37wruP0toDBcn41WDYMUgpyGiJfuLSVzE3x6+Fw3wr+jmZsylH
o4HgDFNSFPVXDhjrlIr47uk9PgcC2HmJtOAfqNJvwwbTadntsfQkGW0W1SDeo+fe
8L470O//qNvvKR3jPAEUGp7ma+jd7EJmEabfZfmjIdpVNATaIvI6+3a0iM68mYmC
mKZEArttVYN/fZI9irgxvjolACvElyPLPzT/RlMZg4/45EiUNwa5y3UqF/DUAh+5
9uCDlZoIEXqt/cc0TP/B1rSPnpn6KQDXoe98Wx+PLOz4+iJgks5j1W8+x+nlK5TE
eA+fy11xlZhfv1rJnBOXhXQGw/SO+OLAHYOKSMHjZLYFI6JppZpYPKyA1SFIbMBg
Yb5IMlaGMHABMWp+G9aVWJEDCBWFnEVYgxSkHdcpnJXloe5z6va2A1sMpT7aAEg6
aW5O1PBr8/BXCDtIkmYwQsS12tv3pz2SRq8cCH0kb67ANLkn5r2EveSxnu5s9Hia
jxcp9YTDySFq6TAgpnLX7w==
`protect END_PROTECTED
