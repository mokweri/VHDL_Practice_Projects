`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jVuZx23HRUBVDn3I5udX1h4Cw57yUd2xWH21N+uNRLHCcwHy4lcGbYNnjoOdMLor
9jQLUCobf9NO2+PkvLgdlDpADcxxPRDkZLr+qAelhMdbEtC3AevW/A5AmqX2lvQt
+uPoHgi/QBmQtTDwutpx9kUyqj/TDZxp3frsqOMZe7D1RWeNbhYBEKJvNWNJ7IXi
06J/+F3S04f5o/3fxUmn7GK/I+RQliBl2GjzEG0CAJADw1RhMwn4ce55EcNCC/SJ
4KL+vWeX8aYdJZYnptOOQ2q8TE4jnU5+aMohQjg4AA7T5RI3OBsH15PRLTj9N/k2
W7nwWZNiBELWhBduANWT3Zoq/g+xUq7JoIjfynwHOzPif/47AVPA3kzrg3qBAjKj
V5i3PL0xVU/wbdS1xZhwku7OP9f5BSgwfwfH3CcfVegEA3WA4aX+BtYsHyV15ZrN
4leOeoZ17SnSks7KwCwI9x0UnC/c5iKrRxJcdSoeUGozRkSMNtbWm/6sdv0gURuf
lC7GCoPH0KJ6xlNrfn34MXoS825d4epYJeLZyeY6P/wgx6Uk29/NIH7yei267FRG
d88kzkM9YWKuTa/cGC6LbooTLg2AtgwU0jqPe/L71d28C/YdiUa9naJkZWcB8KZK
WI0yqCUatmxIfWrP6SmpvAQXRbS3oTpxC21weu2uknufyKuULTCsh8PRZBf9jXRJ
yoU9XHm434ihXJgIgbMcwTmBrrHyt7iVb4w8MN9CoSFho6G6FdwTBAvDjxevM9n7
Ft8PefFsk5QtgrelRWEKr1iwOS+tJjP5S4FuHupRPQhRnsuvMPFHHSsPMeEEfDJZ
S8bfLDSzrmVWToENiLZ1iDx86PKrFdDP2alsVxcC+CwOpXVBlqtyhFxEXzQK7sVQ
GMnIG+TNEsB1taJRgtS8gUJ79CjwQosWpMBCzszDTB39ZdLuEPukNhS9CfqlndLV
P9vmtslmDs7cMSO+lPH5H0SiY34QH+rc4G1YCRq8sonGVO2tnEM1Fknv8nW4p6Fq
A4kOH9GV8bfD6zUB5rV5nXH2DyUkQfjg62PHNjgjlvhFxTEGrN2ePhkRysy269y9
`protect END_PROTECTED
