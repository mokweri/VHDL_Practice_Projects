`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C2B/3zKfPGLOpbqmXa/IOhZ/n+rnp/IQxmza8cpZItdEgVPIo4vQpAd7DrswP41k
94EXMLKU0X3T2UlQe/nO+0X05WR3x85DrD0x2ZYEKyo334l8vL5+Jp9G9+1tv89n
P4EPDrnwtSmIcY8An1JI2Qj53tjmJ2vjhaGfEOtvqSnIjueDqXVzE4y5ZKb2I5WL
jT4GTa9faz9GYQ/H/oAMEg2aPoTj7onW2Uv25VwgeGmUMtm6Dc5b1NLaHAyB84E6
jxUmKJ+FqEAW6JNzlmShDA==
`protect END_PROTECTED
