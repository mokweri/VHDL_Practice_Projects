`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkH7U/0p+8vtVPt3NO7HudMmmVNoSsxgL8y4CnVfUKaI0pG2tcXmSTPZN5ofiH3F
irssPVDLWZ/VMPhr6naXqyNblx1QsSJ32fWLu3QEL4NxceXbu0hcQyLgPFW5h1Nx
bsmiFN42+sBR+7kEh1qUib5j3c8gr9nIyIcLai5IBtApTRyoiVCuDisCZWzKdgLb
IuAzz+PIFCuWpUMiHcqdbu3huXbf4VXdjv9mc04wWA0hiwmtRHpPqn/cIemCTTXi
4LzQUH7TF8E4MR5NbrKzFOM0nW1aJ7mYdf3Z/StMF2+GOAZxXgwXNgWoVp5uWi3/
qGEtkU3IbgnnyuZib5j2X5IwyCXaMWe1EQDdz1nQnK9WPCAx23G1SfQsbdUNrV20
Y+jcDthqMLxuva6Cn03aj9vxJjLfPJE7J3gwO4Zzj/2Ot8G3RUidreAHl+su9HUU
co2XPMVrg5B+pkjLCu5UsM9N0r4qiU9I5dh+W23AcSCZMbVDZTMDxiQ7Wjny0X19
DxG4azQcjLm+nRrL2gwlEhhEPa5fjZaYvELm1kXfJ5o=
`protect END_PROTECTED
