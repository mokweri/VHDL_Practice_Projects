`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3b95yLnisQAXVcZdq+YozB6usOVDhi1pK5hOU7d/9QtZun2l8o5MHRSm8+jlTlda
eCjVmYIknbr/k+dIbttdi9Iyx+QzVzEXvTeOWklk8WZIQylhnDvk5FCrXMrthyfk
CrK3B7wdh7SQaKqOHSSGaPEewZtqJy7jFqg1C8DsvwhR0gQXfvj40mh2hNZ5RgqP
Vbd/H+A7BmVo8OTmw/ocu3vnQvANL4lc3LaMCsjn7yevlrP1AQf/1uHJ2I5sRVJp
0EZQkihIRUuzDkGIbJQSaUo8SWr15Qk7lhpSHw9AGRAeog1jcWhZ5IN7VeEAAyTr
onviej7lV9mNy7AH7Jg7IFtED7xE8l3JcOSFiT0cKWAv7DLTbijotNd3taTZj+c2
1DgUM2z+9588wKIVdfn7UQQzpGkzwc4Bqk1MSL7RSY1PqIMMUbfy2pvrDwyZKeDx
aFlyNKN1CHM9Cpj9FGt9Y+UVhm+t5FdpSAXoRPiv/ZrAyHs4NukEIeMZNwwm9eHG
rEYtgY7UgmWi5Zasls0mArE52ED70wWvFzHBAjMzzWlKNmrrfb+cWFnmtS3FU1CK
jbMxmy1ze0c3u1pxHnKFIr1doxSmlMI9dyl1CjysEpD87vA1pWaoDVxN80HHiPS6
klC/2Ge7RYqco3UTxhUYSPLpgB0P6hiIL67xVWLYTxl0dvFZYtTnU7EsWfszN1jE
A+KE0Gn9sAzjiIPNuEWikN1UMDfaIHQnCkXLjBek86jFDphEnFGc1M2HACRz9b5z
LkFwFRQWseVuaqwSbfiigfPHEKsR8XTkv4VPVPj4BgXDJiTE1BC68vioZPjEsGIL
fub4Ve3eEAWzMNArq8CjYppGwNQ+qt5sBzhiRkB0OoC2lyYuH4Oo27iGtYViI/fT
ZPPA1NjOWzSP4SzBKp/G+jFuJJPUePRWkwZpTSLg/hFRNcD4ciCjX51I43KohINf
NC+K9ttP3JrIBzh2nsUCVGzHzUoei42ukaYy3RLgn5Aqwa9uem3ZWTqexf00un87
rgBJVcxujjmH2DOv1sOG87V8Gs1/BTqqvuM7iRQ1tbNPuqHVtXGTfeWBeFfr825e
1lac81ucqMsSvhfo4+KWMxF8PkRnSGMg778i2M4YLiAroXVM3wOlL0ZKVIRhfuSr
pYfiHxGYQ3kNc82WEVrOUBgHHYiIvfTfbNWSJCUQwXkSwv5g4lFDr1ZH45AvZDM0
ba4ncRsEomkpx8eXhFHUwKfb7jC5PualIGzrsuFIexEDiimnBp0P2541fYODzWcx
1KNPK4OP26HG36BfLBlEgHI00MqE458dKPHH1/kcmdciFqjSpr+3dA1rO6Mmn80Y
BAl3Wo/sWZpy8sL8+tW/kmGgCBlwPUVPc2UOr91vx+oN/RJYc256zi39PyYKWfwf
IqMuZh6BDSJq3MNG2F7BoXA/CW8/ir0uFWTSMMo1kdATREVcdI7auYrHzpCmqdJ+
hDBljIB8MmLOxlX2+zWx1KFoYmj2wUGWD9VR4S99cYAIgUDY/OUXbdtVwNmG8M1d
ttnVukniqy+OyMs6F9c0T8WXLv4gclOSzb6/WZ0GvHw4BJM7X4905vFMDsS1nD33
NmWWP1DFQETmPXUtKhENBNB8EKb5LDc4du9T1atLnl4i0A7qbhYucS/0cXBi5uzx
b7IARR4IIKPzBEj11FfBI5X68cn12D73aayLkb2c96mlWbQdEEx4upQd+IETB1xm
Y4w6ci9f0qGhO7Vacq5tWHANeYIYnQjqtVCNRKEaJ1sxhOi00eYNGC5kdk4qLzNu
`protect END_PROTECTED
