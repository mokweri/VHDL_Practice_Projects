`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymfN8dS/1bIVWFliZGE+C53skfHK2vkFTsItjsNGKMWTSMejGBk7HrndqRonOa09
OBi4lGZapSrdCcTne/jf11QPAsFaI1ArPvzIaFUEWfJHEboHye01/nm+mn0sTc7T
tF7fF4efJVdto/1pCF8+w2jvJ/tGoDJvcoNzVKqiBBapEqiZKnTCnBiJwtwn/LI9
dBT9lrv/h1WIm/FB7e9tHazOO0bou+rzEwmZ5+eUeLyujjiMKoIr8XjugrTJJ+P7
duQReU0zAUS/p+2uSwPjLun3nmPzJzXaGofz2ycnNXnWLe1ptCJ1RuySeqAZx7rI
uU/1QTxVE3ai/dL5Dr4BQ3LWZ5+Iqdng1Db6yUAZMwreo5YGlAfuC59vtnCz3ViY
iFKIr1+ChHM4xvj1U5aFecqd3IC6QT1YCbaoKdpyuJ2rlgMQKp88xN51jK57v1y9
PulAxCB6iw+p6MKBqJ8UQVc+83lSB3I/YBMdCkcsGwLddNHvwilUmpOJ8L5IaNo3
sJURLS13aGjoNBoDdEljObE3A0v0yvac1ieLHXJKbgYCcD2gdbxBRZ8E2lx5lH4u
FQRE7Y5OoEl+7BalbSOP94ZgjLh/u8jTjYcPzbWgg9Rn6WIZwrlwLoi+W9APCM9G
vhz540tsY3U+4OLEduIXL5bu4TkZrD9TD0grjq11/O9fHG//1N0zxDkvdG/HBFn/
+F9bKyqmuRgqifsqVoYBWZIvVXVXE2Uyh16AKZGLd9F5GVNz+pWrGXGhERw7tVF/
IT7uJyH6NhcTOvhA0mCbyT+2swwvt/0H6ET9pnhPZ2kJuiIskLR3TBoc6CsZ5Dc6
d5w9FCnzJyukr9XWYTxQXYb30MENQhWTwBr0exVCOZeeoJSui4h4K6QMuF8F8vfl
RDZV3HkalzZu+QI9bM9wq1+O0K+DhSAG3Q3z0ZZOxnIhIU6S3iC9SQwOmczM5y5n
eACYq0LucDlHQYvP58RVzCLbibULefXTwFZu3lG6Cur7Lmj1UL79NNmBrmOLMl0T
F1DI7fgiB868UjTQhrGnwkRZCBEtEGKojGGtDfrnMn1lPJAhJyvaNyR+Hai6IcvL
a8zTl+IYDuaYr0I0H4MtJgxc0QaXi32uejdfesZc9Mu9gjq0DFEPxp5+oGs81HYS
x1LG4D395epL/sfLr6UzTdlkYD/tfJlHwai3LjjP7Ftv/5YqlS0kWUOZq3OYVI3T
gVDd+IbIkdjWwvzIYtRMymqFQmNX5FzRMEdUiQ88aciY+f977Hdy74RA+Yp2Fmma
f25NypoxoQclHBfVFqaFCVLDJjmUEp3c04/zumKxNDZbkHWokh95BLf2MqTvG7/D
DTcXjaqk+ge68s56cRuudCwcvXqLxpJ1oB3Frmm6b0raC15tkby1/pK49/HYZKU7
Tz6G0+KIjOPz+8Lj+GNqIxuC/WdUeqZ9qjVSL+YfdHzvWfpQv6wv5/3pPWNXLNm7
XVEy6fu/zhK/2NGq3bWQyMSn/ReHc/DkbjqpE1OwDqRNderd2ndzMG7AUDK437jV
oTTfAqtvyJab765vIUCTi3MAc6l5u+fuAooiAt3vBT215C9nzmEbPF5WOzRia0TB
slFu8DO0LPU8IXtWnTylSQ8pH5YzMKq8fu1EHyklRfL11CHZrufT+jPjsIXWxoZ2
nPbSwE1P8jX9eiy2qdYhtfPpBuD7y2AEAmrg7wxXB23SD/ggff9vTj5K7w4gsoDG
BZL1ciEI05ODajUOll51gFTk1QTO6ze9vnQmFjBYFQkFvvglkVprbTWI1U2GBqcU
qK1C1oGHfTdbOvU8hxwa8fhvalNEXwtzQAPvHNv1Zp6rlBwNU+z+x6R607AXw+l8
fYFjb+QFOBJxzsjCJsWDLe0pqRlnIrL+nTKcOEEw/8ifb4w+d78+xp5T76HimTjN
HWizleqzEuh3SBCzrmvZYp+UhBY6IctbkCSoEmIx25DWybjewgMqNxlf7FxTog6k
Q70Ru7eUh3bYrGSjW0bnzjUYFdxQPV4tZzTYQOVdf8bSnQLJYyI8NTS1zuVaZA3J
mX2kmGDvuCgGksNiApbqVG60lNpvNbmaBRgIL+562GEvNdRBWs1wg5A86ct3H7Sv
3MD+56Cv+kYj18evvZzcXS2jM//+sBV9F9rSXtbk1LjDbi0aXCDSOClFrS5DcE8I
yX993xhBo/MVW/btgq6Gb98p8MSCrVuRxLkbsQ3xnJ+j2DwecH+0/ZR6MkD8Q+v4
YrvaXDjG7X0fiXky8kktPvhItO1cdPKumbmp3qopTaPwA+deJkfbYVjtcPzzm9uv
E8J5DKNssjg3RlPJg7ywoOj+QqJe7s7j01SruM+WucqxOWISMR7ckmJl2vXOwLLe
eC2SSlJui4spxO4Lm8BljPx7rj+VMjqiXcxOCGqliTP0tcrtaRjWEtXGO3iHDHmq
SNieaWiWVj3tM9l+0cgu2MKmkZkbUwv8r+2V5lz8k78snjaUr0+o+Y7rLWIC/6eD
uL8TI0OzgIl89hhWfPcNe02Iy0q7tQrtCnYpxoXZyBhuFhr3Bm1YBU+PZR1zLf2f
VD6LEkxNCbMb7NNVz7J5ncjdjxSOMpBXNF2jEnLq1yiXgz6ejsJ4ZaBFlHoCkEdm
1Snr5Rk9RjIoS0ySAK9wEw2kShcXiyKZsYQCKWBPJ64=
`protect END_PROTECTED
