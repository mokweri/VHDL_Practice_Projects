`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vw4MCyOes3ihfwuNUNwvFhKFkuyam+0xsYcc+lMfWdjMYIaRTd82ihkooVcuNSAb
nBwCiZ3QRO9CAofkGT3Z9T/36tfQZbm0L6gM2LkV8wiaP4BysLrLboD1d3JOI4wO
Qw1oDJqCrZMeANl/PUx1gCChPMM5BGoxqGVIlLEV8eBUd/plg2CEv+L8y3ngtQHA
fUa/Z/BTNBGqYxbwQd9GOXfYW6diYYaotkA8LrBjqtlSDf0KlpunR6EQiFhN30Fc
HttAbyNQhmI+9X5PuKrXinSvpPvmydOn0vKniK1y+TNQEaSOoJ18EDfSJVrWODRL
Zp88iZSzPGusTf4PBgXiZuvXDNwoS0jc6xlbveosb+PgOJrz5ix14RiQQw/WcVD6
Kz7yUiroxbsBtCEcVVudGV8Dcj+D9w3od/hau4h975t7wSnEu4B+aA3xV5co8HDJ
0lOsF7amfKeBlUlAmO7vkJR+efn7UVrkfX1LWmB5r75ITmvAbVZJ9XHh/Sbx6KtM
wTz9Gj+3FjAo7Sjx0+S3MtY6bWJ1zzQCibDp8kzf4PsbxdNBiEj/kdqXUJ/5uUWi
EsaMQTkqUn4989ZxBeSZJv1CN4NoHXqhKmeF8kxj6FEAB90fTj5S9VKoh+VXNFKQ
F1ID3SHVaomLTFcxUh+VVy2EtN851JA1umaz55V60AsWjT519GMSfD/j0SSBxWnM
2+fWZA/SmXA2G8oUYTepD1jdDbbfSiloNTTw8vquYunsgDgWOL6Phxcw116cl63I
AoCkFm03QkpyvYiKi+fmwjiKp0cXjXzfReEoQxDj75tgxf9ZgYc/dlXZ6ilOitkS
mgmDMGmA89xW9VgdT33pqAmCkc1iDjbH0RNZXAbNO0zOjdZApBY+YY58kPdbT0If
Yi5A7rY4/U/ZSCL/YZSadFfwF0gkdA4boWA640W2+bB19dybonJsfsAYY7jTimV8
s5baPgcI07A/OJq17JK50XnKUuK/tZ58maq3ZQrtaVaIPQnzn7bwuz5dyp/4ygRo
fam01Z0ghfdMQhTFXLMQzkghZcLLWwkHbDoDU+uof6BzDrdoog64VhvPMofXM5dP
LbzYMHgztsCzL4B2QoBHmnWa5x1V1PYfM67XsrZDMc2x5y7EVw6undHInsm2yC7n
MTK2hYWvuUk5kTWLC83Pg1udYzr5TAUIDTeTAuYlA5JJIwlrwvsnDCn32fKJz/Sh
Szf/y2jyLy2+4npaUurqUt/T8lOD7k59Xcg3xiDaystF79aa2Wjp3Pp/9mAISsWx
MHFPOQN0TiSNFcwVTIpX20suodkKqAZuGtN6c8jXXtqNsq2RCPYC2vaHOMPsqVpk
xmLjr0eiuBBg+LLCU3t20sM65s1h3hXlXvW7W1VzgjJ3olB8Fg8q6S4fnHQrC2/m
ap70y9lPumDXc4Dsv1syNZ+6dHVJfQ3OJuta+jULChLEdcIrDP7ku+aG5bnjVQhX
1g0dN2HdQw6Dmhz+JH/PG41K9N396WtBymDq5DNNKQJ20Rc1fSe2z0kIrJyQujy/
/0YZMH/xUO7gd6h0svvy4z7P1028qZIOOS/clIbaEaaDgqJ9l8ieifejpH/evoKs
4rjgFQYmCixdJJ2WgJHeTgtHWAJSwhIHgY9YIsxuUstrdM9ndvZjPplkcd1mvn0t
jG6qvMdLOlS+GefSzeOn5WS9ui8EKVF5nf/R7OFfnKksvAyD0vzHfus//2FvjYRN
1oBg3+xyxkxCN+sChjM7DIIB+tb17TZIIfXocb5RNFX9bF2eCbbFL2W5IBJMe2r6
VliVByQVP0tJ4K8gcF5zk5p4+UwZ4O4aygyHfPc6y+f3AdB2f6nrNT2y2tzfWBUq
CArVFKCYmxvDTKuWEWGgIUJsgKtXlhVYw7QAQlEiDNx7YitC/nlzFRlWdxSH5z4R
`protect END_PROTECTED
