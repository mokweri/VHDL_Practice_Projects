`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jxNrGw609mnQRu8uS2A5r1SoJjFgNWUi6RtwA6MCtI2Q9ry2uLZDKCObEDiHAtMU
fvd9i7/dpCLI8wCN/vf8uxktLLNthxMp82BzJzQsCuEvdJmXIbGppq5sxjJzQ2dw
GpIMYMGgWtZ1yTtzp4BhXSj6nmRK6UsF7finT87o8cAAY9O29XIDCCqxjk5KFzax
HFMcWfz8TgkjSVPOrmaHJvVlEn78qYbTo9hu1GeuZkLpjvRDg7eGikhjolmOvL+f
oR/Y+UFbb6M0nXv31M07MNf8Wq0+rfGdWdnFBz6jwZyLjwMMwguEVyQJvI8dg+jS
g6oBQwNOOR8MiGN3NNQjCOCR5VwsueJiGpYYg/s65ndE2IsNJzy5ythyg1hGy6qq
y7qu4O/eeDLkMqt3UOqcX/FqxYKEEK2jH7d006HvcNWZucb0wU6OzHX2kvtK5ptY
KRUG6CX1XCti0mEMx/eyip3JmRzUQqFg2AYxPppkkwb9IOjtKkTKe/82eBBKWCua
Gokv7tbPkwWL98EO3q2PFQQ+z6G0g8gf49Cfws4vkU3xXKEvin3Xf3RERIDr+VI/
ll6gN5Yhj5cPQnwoB4NgPeuQtDA8DWFWB47X8p6Q9gGDclz5E7SOayq0jRCoBCW6
WNQLrDjlW4bQ+wjSJO289n8eKckkuQHkmUVI3ezmvlPWgmRgfOCIHVC6Tfj8wwIK
S0U0OZmhgjZSAgR4dQjUzHQx7f0oCW98fDi/aaprzvM/pFxefs6LsWpOKktjzn3K
8CumLEzVOqrUWl3uez/lItVdx0Juct8P5+0nlZiVsruZFTsoKAlT0MQ0+ucHukwi
`protect END_PROTECTED
