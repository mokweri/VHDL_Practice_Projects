`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h0wywfgevYhbUwEn7/+/vMWCZg1BFN/SO4hgG0EFkbQelAgyOWnQMPtVPbOdV1kw
9TzHNQmwZe3eCjLj5JOF3Gk/lmzd+Xc3a0iDl4QJVMIJjLWWWvJSnxRvu/s0stNk
gtFwLtNIgoUyHSXb8NsHDPq8tNXWCALGfCyOx4MH+xkjNRi+Z2ZiTL2Z9cIG5Mk6
FMX5v2ziyUmdwhtzGF9fe717D7j9M/XN4R8torQXbi3IjRd/Om8VusTkit/PAt1y
z5nMaKHP8PqUTpk7fyJgP/fz0zQdZMUy4YBigSPgmdBdbOmOaEBgbVPMc4STfaxC
6/tRxRSMwYznmTB2b+H9aED5fzyvd4+1SK4yO+sB9xYWRKzC8OqWeE6efz/6ror4
nNZomMVGpNLXRQVbNo1XXvAoOI437tBy8RFgvPV0HxFm8UIz0vApLlLqLuxPIxLS
xD82zILZ1IT0h08blo71TBlPjVPSrFYQx6E1GPUkBpQpl9+ARQuut1QMKRAhrJuw
/tXPW503sgth7EUo7uiNqF/oX7NzSUcp1vEOkXcx3b6Ti7X9KdN8w7dQwjXkEq4C
akE92Vx530F9uz2/s+7W+DCFOS5+8Iy4qFHijll8YoCfpb6OHfLbmLU3eYZEFyBh
Tc3XcUkPpAMiiq8w48fjQE7zLkWa9VtmiI2PUnfYsdS2vAPX8cuXeontJ0VekSeC
zUf2nA8W6mfnhKniKb5GhRT8bfWU2/m58EWqQCWFMvVNM1UXImWmZTgp2XWECR6/
x/1zoTyhoBC6J8XRE9oyWRafKvbmMHyJ1vsHWVXxjycLWK0si/Rm2uRf8+6crXk5
RO21yeexAFF+ChZMD4UNCily3uEnsEUJSvYfntw4Qy0MTo78cAPdvXddFe5OIRqX
`protect END_PROTECTED
