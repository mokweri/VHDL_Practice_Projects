`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JXDvcG23T+IWXXrtpo6oCp01xueWxjzQZ2we5KjXSEOHLyx+c+KHRh9C3tdiEo3q
P4ygQUf8FrZ4eRL73xoDy5dyD9gPNdReNW17QtpLefA9dJCsDPCx4ZiEkMtgSQ9C
EH8x2C5vssOtXg8bhm/wpDczPQfyOBLufPi3TRsaX0ptus+MXzboDVc/5WpH7Olf
rGJYyU4nPBMrX51HqNecQKbYCbZoe6k29i/IeAaKP6ZpnfIuODn8rtHUbBVQQ/5C
VD35n2KJv4Re0WqjQNK/1cZDlsT0+E6u0/tzTXRoWdNAMCd8Y8GFVFizjeybyLm/
9szWxU/Od/1N6kQ8P0/ii2l7DISmWCjryTU3DDjB/5vwl8t+zpTJJBwCgbCqYd29
p8nKeuMqSwlodq/NSSXK38FFyPd5KJW76IAHPWWAdv1dHWJF/iDlveXeW36zT9GK
2slwtS52bhOuUP41v7wur4wX3QDnI2aMpTLrMuLYdBo3pHYZHQfE03xPbQJmbT4F
cD3rkN2nSstAChfuba5FsJ8Wj/K6efA6BHcSz5eKa7Umsnw+wLGkRH1673RU1940
6hFicn4voScHmtYc26s4eYgrlweNUHPPbmAwzx9s5d+sTUp8oZC8h1NDx5SbrelH
j60CsSdLdz7yAsXxcSGL3BLD1VMK8P38IfKXqfDHa7am69gNkqQPabXF6U1zZ597
t3zNzfjUtAAsMoGqi9DkIeyhGLHxOcIKGUMVRIEOf2rtRqa7dBtZfqm6h5YpIdUZ
9AZ9u7z83ySdQc/dNs/tyg/URDlA2cpjkf29ZXdnHLvQeWrRfHidkgFfnB5cNnJE
`protect END_PROTECTED
