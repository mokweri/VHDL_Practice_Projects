`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yA2GsYBFjCL1kel6gzjETScfc0mbZumdH5bml/AkoMaPX38iIDbE7HLSfYctoIyv
ePbtdKwUEF24A6ENrZhWCpIkLQ5Iq0xSh9KC4EiRZ33fJkF5WHGP6rK/XO7Y7jjr
ZT4GIqCz4Bk4rFHQ92fzLpASfdzyi19vAmxeY4T+fl5opOouhUgYHLLbqiarGocY
Ho0R4+61FlL3YayeWo5eCK8YMmTxqYbYmlPVwCthHMikX1KtBx9bL0XqlPdVTt6d
Q/MXemULFu0u8Zrw4wCpPU6gJoE1iYKcLRgbSJmyOM8DhXi/MxG5MtfdYuS86Gh6
L1K5vcUAfruw59NtLigHuSjl6q6AkSOFtTAp9VlTd4ZqwJsoQgUoAVuDxujXZhZ3
kQR1ep1pClvmVexO5Bn5R+exOmTQYFTuyaip81vRbb51I0FRcSSd+MYYrzq0TM+3
T8gjl8plVixZ62+EUwtjidAkNdFPWbOCa3vOC1jPB1gD+sm1UnoYpzDFbELmmBOp
OQLVO5iIqGMNLUUJTyHDsg05A6tKJEqkdGYSjDKN7VLYWbQIAHa7eEerp8IhBtVu
pyIqregceMp7V8xv0jg75+NExuOINvcMaknEbpjh5Bm/dfVlw4sATc+52eCGTRyZ
rPFC0wp7Nh23Bh+MYuhO9KMMJh73xiXXVcgQPLZXVTSBM75RsK2He56YrLwGwr0P
fpCcJ80BGS4egQYR3jYl9ZsDJBXcKICaRAru9uEyWjHvjplVukytOAQu+3wtSB90
5nQT+L3c8lzmTiaLHP+5SopgT68mJdMWEKuVs6QKggxMuy44LO+nZ/8D3y39aqPJ
XTVj/aU6k11pXpIY38isD5aoesvNNW5xwt8MgMp5ucZH8g2c+igzNj8GoAU85n05
gKduJ7cX60KalIdmRqJvbZoGQFT58nOGHGUDveLDiGKUAXgGxqvd2Izr7fS5z0w1
wxQTpZR6w+u0WCA8k7GkiDPyIoKlRKgtZlAnLOKQxI7vmXvLNxe4HeNpddpfFfXV
jo76ESK2koOo6PZPMbEAO1sZ2zbryDmHJ5F1QwRwUR4oW0x5YvBu5gZ2pEPMw542
P+2Srk4vrPcP36me5wbmIz7xliKnfL69hLguscehkDOxSvhwZ5poLzz1oB5ZnboV
ZknrDmiLk7ASU/XiagQIKwou/8kTTbOLOo6zTz5PIAIt7vPEn/AjbhZDS8s09T2G
p6hw8nu3XX1jXnnOK0WSfRjRhDOGD13CyOVSNeiBQl2zVHawlEA9mZCYTMr3hOa6
HczotU55uTEcNt9bL6USluUAEaNqGTQkrgWVNalZUVIupJVCJekQdn2QDrOS6bsu
QcaBXJuvnrsqeJquPIQqJGe2rf9BiQoGIRst1QO8zuoiDChNTfSxTmHK1aawW4IM
ntekin5HfExYLdoGOGMEn1Dcuhf1y9NnzaZj1d8XtCC+5Dj5kkg+VEluNyHuOebL
y8gSKWv1M3vfuFnS5X/uaJ868Js1OT4+G36PwFMpfhAPsLx7L8wNOVXzIuZxLD7I
eik8Vu45o86L1ZYCvMnCecE5eBftVT/AM5pZPzf6weRRblqMhUUkNItv4l4MSiKT
tuJW0V9EtBbCbKgnzDjKiiCcr6QVYd3g7dAJ3Gmeka4YwdkfY009/ne4kQQM0nx9
yp5H3IMjkm60iq5hq4KJSAvKTPX6t4E73ySNEj+QJlOR2YmIN5WAObg9QiJRwRF+
dqNOPxXkrxEvwBAQ3YySwDDxC/KMWKUQVgnGLyvbk+fa1QceM3UscNJRJkO6PLHU
jJzM4T6+/ZmYnILRJ+B5Pp4vL4t5X3GMyii+u59/L/sTCC7Rab0B0t52qw7UJfNa
mCxqB5XG2We1ae8JYFaIt/6QHfYLlC9fgA3kq4Raf/B3bpRTWxUY2beeImOvix6V
W/pY+QSpD8Uo2MMd/TgT2/rouVh1W4XuJI99d2y5adJFK047YPuqiLwx/teKWI3J
2orkRDU2pMVS0dIY2BKT9YQBGoXU/+7L2bh7T0u15XjZtUtgP5HSowJRUyXZDm2u
xd6IfLqMWdYDC3tGyGWb4dFLwgstdCanhwRN9ZejUx4dL8QrwsRbNyg5uXXjLLEF
Sl/1cuZs3Iwa/GKbEB6LKUy7tS/rupqhs9hxROmWi0Zu6WDzC4xS+/wuBme419gB
E6Aff8z03H4KDnUoXNe9InM77c94OcxaD04hDh0B/fPvIckSlgvrkzOmmhCkOYOx
nC3c36noV1b8Y/Mi+SC1Z4W23wpzM5TDYynRuXlit+80awDWIaOuLEeVIro53h02
zwHw9ZbVb2dJowoqrpVH6zuA8Syf+UpWYiPIGXbuzjkZDeM6QoFWpLNonSyyqrF+
Og0tZ/KHoO5lBc/KHYah5GExcPNflxrqgs4fOioDR8llv5YMUXT85I7HGvoUHth6
PnRn0z2kdQtMRGnoVkOFx6NPL+6kKDucdNV/07/ukSaf4NYE+GvY2jdQr06BZsKY
6YGMM4kUMR8R0wSUZuCW0EqlaQUWacsA/40+bbDZF4jp52Czd1SLRmIKEMgGTVic
idiVPwtmVoymZyiWnb73t76YwylHWgXAQgWtfq4YRFiRHvZBhxhvg6thfhhFnZId
+NHN/EXIZaq6vJvuqtE8FULUsugB89kwPe/lPKA3AIhJ63utDWk+dhWRsmXcEqRX
XBFoQ4KNg/vrJS+hdDW28luanMVro3Q/LVaK/znyRUicDWHJGBo1HjZT1BFDKZhr
PcYL02JXx1kd5xfpyX3MJFB32PXcSBmESY8yhCE1V8pnhnmSuBSQy0jV8I1rVeb1
yiaVSCeHJGwsQvjZOXI6BrFu1FywJ3nxRwCl4M6SncevOmEZHf5VxLtBpUf5u/wk
wbYXysrCvjc5NO+czRx1oHogPQxYgjdKGNxvZzRXIBYeCVbkYn64W2jYK6Zg90+F
iajggoAwBdXDroCkq+GiybW1oqf+NJ+dxxtkNiedTC+RL8n/U0dCZzCfryxMgDS4
ejJsvnfGW1TPvKPl9RYCgwgxZFRnGJ6OXXacftHOW1k2tACiE+igN+IAIO87dP0i
aN3l7tYlP1327zac18zhgzVgbLlvXqjcvTjAwhy2gvAoIu5PwAwoHf870MzNuht8
TyC2N++Jw5KCmkgaKzcFrMfQ24eXtjb37znxt7COnLk+xbLG0Idg1V5KNGlMoKdk
eYg6b8Cx1G6WZkUnNXayhFkrChsp88GbxhgKI3XOvo52WCYXXeTqOssrhXiqqofI
a96zEZuU5DjtlZWxmRL7nqpr09qh2J8ZfAAMI2RT7NXE2vs9747DRw9/WIQAFH1G
r01/PA3tBaHH6t1koqGX1YhNADyJxWzqpP195Mqnb3G0zsBmw9CniQzGNIJYs/XC
VKm9aIY47CmkcCImSPs6mHCUV0LP+vXrDlQWtW58GUPOwmDOjYXGudrG1vU9NAZa
Jon3xII7IHOVyom2wk2mAXQKe5NvFPuUKgI6X9g9OpPd7WnX8C3pYjDf8xNm1EVG
WOjVD1E1DejHXsqEi0r9LmEp1QuZCFkMGZSUXEjXqmT+2ebeccxwN/zfyA5SZqjb
xTmEEd3BpnxB0q2AqIUtInMisQ6+DcoZaVYdy6AJfQF11vyN7SxhlPB1A9Js69MT
TkgmZuENzJzNpQzHHbeLtQtKeA5ckT3eW0KDYyJ8r+Uqu9KJfFh3wtL+FYeAKIdw
yaP1WfAfH0u6THb2zHY+dVQDINCpoAC5GOYjKPXfSPdnKZrWNkiCJ1l/uXS4uocR
6zOXR13CyzrV93O1FwtlHvzYbhAX6rIULEJOLXQyR/cp8Vgrk9ei1e5Kz5HdQoNC
y+iJmEs6BZyFTu/RdYaK4JZFGh92EVixIDNQxN+cVGqVt3XaimJVGXh5JHO+d+yP
qMHqGL77eL7r35uJ/0QXynKGYdlw2XebPaxDhbCmpl6HoOZcmiAgWoYvm/xRzP0n
3w0/SKrdQYUKXKwIYy6WZs6LwUNd39UTPszdQeL51qWpNo/5kE4HYUcF8f5EpxB/
OsEd+pme3JM61Li6ubsAg2CWV/n7n3kBdPe/IfltPFezKbyaibPuc6rdbvDcEJFe
BPci9HIkL0KGJNQsPWDgSnxSY3pBbmELNIDL3+GLPtQeC7peEhnIZfEaQiQWAZsX
vbQ5GEjgY7wcmxV4Mq+C2CAluvfi8h57OIaDiHAFbGyRcAH1eL7NO9+5LX/1PZgE
NI3OD2/aN3pba+ueWwDdrppJftvbUQYCGvHyQ2iI/35OjxHAnG+6Xesr7PSBcPEG
RqLuqGCFVfRkNZ9xRUBYYkBP/tP749AEkvoymGIzuB1gOWJ4laVM5m7BeaZZbyLw
sxwDA7uP20kPht/n+ycalgvbzHux3E9S5rbKKonFmehN0vd+KQ9rGRi9rK/dhogr
+HMn5J3s8iLBitzvxNV8sNVy/h107BPAEYn5QR6GlrftI1JvGLp9OpAxUfC7cXUy
O81oNHxKdtkJ5anXNZK7j6uW2i9buTVyPSofcs13g8J5LE0EqwKFY1uQYPg5NiQj
RjCHa6K2VyFoSsn2g+USPmJxl/IoXk4PWT6AtoYkmJJa93z0yntMSBtNWGitimO2
p+S80/9bdX0PlDWZoib3kRas/RqiQnDySGwTJOt1kkBdfFqRozE69HHWao2Bvi/L
7niXi3dG+oilQAopcqyzT7O1Y06eQyDiMvyYzfli5cW/GJk6VlaZ9l0WtuUOeRya
5cZs+voDDzrz2KmgHfmEqYXtRyFwyaCa7qoZmqTpcOoGoMWyE74d+XylMlvVzPuZ
giORhJJEBsQMcR6cP0zBTX9xQtXsuUNO5MfZv6yBcouFf70VWm5R/mLE+iNQoiiD
AxnF57kkMMtyQuAJwl0e7jurk30ufElKXE+tamxjguMKEBuI29jr70HeXdIq+zA5
jywqMjGBHm1TMZhfUamGZrMdxCQcQ9GzsyiKsTJ42iX6m9vnQYPR6BeXZjNKh5O1
0n9g4aN//Ow6U/sUd8+tX74DY/xQIJhpXCrzjdJf+SkVmlwhlchTAZln7pLy7QfM
ssnNTvb5a8DIclfUZSMFfIivxE43rE1W2toOz/ZXmLf3N2GIWp3vXkmbH50TrHAJ
JDCv/6yuLIoN0WpDZRy/h387NaPs4fqYpa3m29HoJPXZoZGT6tZDCJDz+q9tZpke
1aqn01zqhLJcVlPTt2NKIBPJbm7j6bhgb/jHyoyHBJCWY8HHZEZL0L/Dm3Fohi/z
Zc3zO2vdcSBadICa+NzWjYmsE9kYtFyVdKJGKAOL/mIzppc8ve+gaJL4qj9YZS0r
ao1Xy8rd/FAq2yEl+subTyS3el8ZE0ZLZF8iNuMnvrm9jfIRvND5BFCAW1j/CWRY
0ixSEKbmRKXP79qD865NoZXowYUM5oC1rIzull1iBO0SGCkfzffFI041cWyneLyL
X2IToXmDoy18QEzN+NqgMpeeI8vRd0wpjtAJertCH1pXXeYolaNK4YJmsJO0DDDC
iFhUQfeZFxKiAgENJwkNdMXBtrCxUTdpOUNt+EPHHaGdo6inW+5eOExGCgUtRUC9
9UC2krnMoVrmnQb/d3eAzMBknseVBa/tVehrzuPeDq0TTrx8+h2xzorRflDFalLr
YzsG7gImCVs+KrfGMmNYuj/uSbG1Z8CZucgL3vDKQu4rmBRPK4KZpa0W96ebAyfI
y1or/8NcZdt1Gwwrt0lKGUO/eUP+ghyZT9LWTCMUgqLBUAb+PURQiFGBCVQdSl6M
ODb3sYADcMT5s1Y1EEWrnm80aQBJShWPp2gUUxz1vbdaz2nD2NA1Wk5+gUVaXjP8
pWgfRT+YEQLZx3z5JYlTETNV+8cdeNNObilKMlgXYJ+Y+Tz6o12H8a2UEHOwvo/v
1rpX5B/je9Jm/JkHUtR5dWdtsUuJhalH251kxl2thG01RZPx0A5fvtkXafnze0nB
ozUuQ+pO2pLRs72xb9VSJEPTfRb40FsV9+l3LpJWmu0bvaerzPF0J9wJDUcFu4zK
kTKdLdOzbb235Q0IFvjnCi75Tb+OUgN9Lg0T+aG/l+XAl9JYBRWuksnGoxlyxb2c
KwSOnD158UHojQhnYaSG0bhdRQ2j6H8MoNZ8dPPuuBhEJquZkj9KoxjNIQWnsnK5
/fGaW2JUrBE9cvVLv12hklWlkCHxNizrl6w1s/krOPUDQCi243ieH5ieVmn/qviQ
CpgYxgEnegXsHTvx0kG9nSALFnJJFNefB9Jhrwqnnyl4oRveMVIwRKLa7zF/sNmc
NG2hFUmMnDUsOlQz/Z9K+pEM0JIOjRZaHTe84PjYx8GDyYWk8+BnHaM29ShyE6rS
4C2XPMv9z/RQJYbBeXmXfVMT/l6PKkiB0NilyIMpYOtsMIyOj7GVt9ALvKx1klka
X1YYx9AP4Tk3+HfzfjBOIEDk0XKjOIH2yDiGUpuGI2XARm7bDsSKEN0C/D5qHjti
PqP2wpMWE8rmIHChalox0OjPPy5nHbnEZe5ZQiYns64iBByjlwJTjggcIiKyyGmW
foZAbX5T6cBlhfUABCXJtPyZCSqy3nXPqvSEZWFX4Rhm/SiutWHmCL8Xre+hlI+S
A9ae2taXNgOy5WyaWYrwHqpDH0a6CrM/E5+jvWPbSI3wlqpDfZM2c5OtuddK7gRn
vrvcbInnHjb0ZGm5EddVGL9eX2kKL1nQUZlooNRhHKJOX9XrLTp0AWCXE5iCNFFG
ck+1VgrVcWOvRl5qktnPX3D1Xgy3vjrgz/Y/OsN7kObMSetmu+H6/q2DJU7wAKYe
4lRIQRspsTqIRaXfWIsb5WOx1gLMX4zN/zW+72r+czdScYWPJM0aNM4pV9a16Fti
N8365oA9b2vCIJDy0/RYn4oppPuJkjoaUY+6eV8grcK/9SK1zdxl5Y5cHTGRC1t8
g3tzGxG+VH8B6/FkWnCpPm5MIzwWZ/Y21oZTiaSZNzpJIxBZjQlllpIG8lMzuoO1
gAJdSslAC1lqh7SEqTA1TopGoJfuhDGiSSBCNOdsGf+Me7tNEjG00n4S1JruNQmo
D5Qjn5vYIo9jHXyLoxw3GN4gDb/jworgp+7FrlOEa55HQyDChl8QRgWFOltOqVOR
25y+6CAGnoZH0Y+lwlkbspPGP93T6LEVPuwpJAsHodmVtZTHZ7kSB12dq/k5+0OQ
EXEMjmbsRT3ZNvxWD9IXQIzYJV4w1UE6BSDoPrfGV+pGm7sF6X/QyFz0oCRzS8Ty
k7pdO7ZCNPIKVilAOQZVY4mr9T6tpf2JOqZU1J7vii+iI6dGfGsxywej8qs1DfnD
qSvpOtR9NdHhVh1sQmAq/VneCBu4ldeQxalSaiDozZ0PhdTwBsxUNLJLBMko4ehV
Ko4d64bFHqjrUc8H8BSHcxcflFfWDhTNgdZt3vRgN8fMeQF8URkuz3zI+5yRoKVf
wRJOF5z+4MV9VLLDj9scwWOWO3JUA3Rsosxju4E0cYehGs97W5CZO2b2co2vkK79
wau3U2fHR+MpD9rwVFDN5UK8DCzMtQBAj/mljni5YWX2WKuPGhj4CMg4Mw58utx7
BU1nd+JrQj6d9tW2i7zLc4mo+n6McD8ODoNGy4pZ8VA6zUooo9irLht9JCzMIP6F
pGTcslbgtID/OMUM1twLRAlG3ZLrJWkcBHUrmUWrlTrI6LevKorbEwAdqwfZtfAw
GTofOwKojxWAnsFqoUt0+pobwF0ER6AVEXfzGeFF9W09WXHEl3fvkyIB5x0Y/1zv
qZiSx0uhUEJlanSCf9226TcjLwdnivUfIar8qC/+e4+44K3/Y6Z4NR2/O1ln9NlQ
o3ocOev37nSkmpE+HORWW4LMmlJDNeRz2iR6i/7zCR6lqH0jme/nsw/12RzKnpdJ
E1t20w2pXTd7yFx3l2ps+TRsjJD85FEhZVYWAc7FJ4zBnVlUYGNP4F0ELvFyeSfY
zEaW96OJ+p1AGNG7eaNj7tTiqA7jiys4HJhXXhp3ZCDet2gqMsmA/zbu1IHZ6RKm
DKoi1qa5l3iYlqGTY/Hg/wX1X19+SApff00zOdL07JT1Wg84h36zKf4ldiHIaDA6
QQuGtqFEX+G8xJw+KRFOm9sA3OU8EiPBvfH0EbURqL5iRSCc8rlbwClPqRoEUkAP
twQv1RqTQxkHoGccRkmCFQGOslK5BLKgGfpDYtgB/oyRsBVM7AT2ph9Nc4JUo1S/
aThfWvG/T7+IHQmMhj6VqJzjRqsOpta9ajIp4HjRGj7wpdAf7KLJxE/RIecOvdAk
GiwSt3HHcdEYz9fVr1alb5MoEa4fwU4RFUBJ6SQYOlw5H4m04IuJPxKwEea9owKh
/eY+ppWY+VIvwULaiwNhrel+G8LktCdplgum8GrJ7MGROCO1aOTJY8pgaWcymF2O
s0JwZu/Ig2DB6YCm/R9UyuPOpfPVcHblwe2lX7b8NZCVhhRhipsKZtV1ZwQpn/JM
oWgSUsnJAM4ZJzKC3ErjsJFyL5Qw3n+nS1/pVKWN7lU4Sr3kLXIy6qn26uBladQv
Em9+jH0ycsA9rfWdeVNeV9xuMxc8earOVaz9UCQOqM004BAqTUxA08U9/LXrjmZS
M+kKRoeZPyowv8+wd5/KSj3r1YtQw7UDsNOI1zGRXMCNQu6OYGg4GaWeN17kOBxy
hnaAjQ5i0pUFklK6C4GQah9jR7E1020TPj8EYp2be7iJvzQLKeSW0qFMolJPeAA/
2i3JIYlCAuGwgW4l+t8U0rGiTArxW4UhoMV6hSELjKvFUInJI5jLNke4OPySO0Re
jdGRvwRZ6Bms5c1aVy4Prheka5u40xufa1z2MeKD6Mexema56C7CzgAMJzNu0Awb
Ft2xCSstqWHgBDYZeO2/xpFgdAmlQw15gnRDaMsNESWox/p+qh5K47takNpNtvQr
2WRyG1KXp7vTYU9JcVCuJ7S+USdOzbrL9G7O1CXp8MkCvuGneQk9Nvq9h8yLO1yo
bRgSrOyCI6comjMJCRMBx9UWzNDMbuSg//EXSNN6F5EAqXaDhaYcYMzRoMCi46jD
9c6xm41BAy80STFLoUs9A3B4M4kXI1+Oo/HJZ594sJ/QOXQrPeU3gRME5JjVI/kR
xdupQNYfv1T5cAJK0okZ3KRfgqgLCtBeH8wAPlg8NGu+SC/XyDNT0Q/r9BzL1BEN
ngmDZ5cYilZX8l/y0aI6Bkg3dNqeLCkH7kvsEnOVtiE/MJYubgiHviWHfMm5nv2d
HxT17+aPXvIqqIvU840bg7Cq506eV+xxQaUTnAhTXoKH707+M5BlMB++aXynZ85b
L2pjNeEB2AnIqVeA2kRTv/iIP7KWHAFWfC7AE62jFI4SnMdkAWlT9JqZb2cnf4UM
gSp7buvatoaN82iCK4/m/gJV1Cu1tHNSD2eJb3XJTGwhXuZv1LmTYvz/edEVgydq
uIJQn7WXTpTFRYfqVGXwsDHlPd3B0UHdyUKs9Nw+7Ao8lFkJsI2ym599/7v+wSRE
T8lWM3u17n/PdH2CqoFAlLK+SXIOf8FognbgYomBUdK+VHtS6wSvpnZsqxR9OSpb
63NaWCD3iuvIDE5r0APZb9o6eobr1lI7/vtuPgUAHZvGnlzK/haRdlPAi/MGWbST
iEDLfFoY2rh88i78sXVgM6jUYAmdM97iseSfSGkFCZhhIa2f8ZdklUbZU9QOvkoF
ixUT9bdcljQv0W8ke+/6ui2V9fQsRKOcYh7P2nuNlvMzcMT/Hl4m0b3bWEpqJZPU
smVdbPBJMJFm6cPPnWhCqpihLzHbs+w87KjHIqS6Kx6hSV4IdAv4Jx6Oaiu5t4Vc
dD1HZbNPtyJJF4vny4TZ9ft6v+hSJI8E61fIrNUGhF6DSNvxpRP6EZiQ9JAYpV4E
xgEIlUl9n9lEcQ7wyLMG+LIjSniL2omNymi7xEEkKtiluPnw+gUUw4P02ciIAieh
wqu7HrLq9nkDfxmSdUHf9rh3Rsr1SGnOPJEjc9CrY3o7utWAGEJ1Fb0k0zOYwZdm
peALauzBu9c+GVqWKOdy43C7pz5lpPCE9QqcrpUFpynskMFHqYhRwlG0PZA6fY+n
YjF5uFPGzE/ZM7GMREt48K6CNuvT5gK3Mf+4fE1bGa0ytZOt9O4t8fJjQCAAKBye
3aeo9eMhTEGSThFL/8gDRdgnB7u43yBWi+BflevlWT69Tiv/BAOwSR0u3nEKWNpo
he4sNKKpQBe8zYy4GEGABH1pP9ozQMhJ3mvaH8cWb0thY5TS1v7P7EdgwYdpnQyS
YDK++WVk9i1WtuKhXeJgUtcmO+s4912df1iPHHYPVnz6lwkbgD9CzMN0r935opgr
A1lMx6avrFZYF6fQrH++zgAJoAuCvHDNRNXfSrr089g5mOmnbBh61GmoRoAN37wS
EIs0/14ioqb32TQlYhfm4tVCgzjJJqxvdzeNIvYq3VptBPj0CO4OYA2I2UOetehR
jmHl/OGT5NlpbMDJsoJMcOqN48ZmWOXzu6Q6UUXFEIIKKMDzzBnOA/UwIf7JIGgr
n8fHn8cUeWOvfLoIvsiu9r11xC6FYeaoOU5/Jd8yUbigd/b90rKotnaHZRt1ydE+
FscEZADgmrTClk830xOTDjbbokczPUtKRrCLh9/HsuckSpjxnRTf6AJ+OAoeo7H/
gvzdR9H0h+yR2GiqpV4DmM/1DPMCyIU5B5nLo97KW8iGtzZ3aUyMKQnTEUKaM+G2
SONo8Ry0JCGsFtj6JUPCALbuqvi4wgR7X6iqP68l6uM3+Pznq+83+kDbHe/MjqkT
XtFIdjhH7pLX6ixIbxpXavuumfoef3PK35RxvZaKN3jODdZLKZKJVGq75AA7Uf+3
bp35hTLgRWuCEGzwZlPvSFtDFeWbaRt+SnRfq7KvlpIQenH88MP2FM4hZYq8Nssm
HkMLav0eN4d5/zsCOzcDp9x+NFl7hiuv0XMtREr67TKiFnQ0Dt7JsNEV1vKTlk6u
duqRNFLYXj7VLvZwCltnSI5bSdmmHokgTspWoQfH9e8/Vtilj4NcnnpIZqS3JUW6
NO5dPm4tLe69Q5phju3AErAfXZnhAKgoVSMY6BeIsakXEsuXFhgg1xt9uio2XVUT
htBtvG/Y5LWvcsQuztAL8LzR7pk5CEdTRKeU0eWTZjnTkZeCm/KBavK+OrxBfz+0
bSHDtxysz+2EZYcnubQG5iqPzrdeyp2v7u5esoirIBeiO3jx6T/R/L/24K9EkLO6
2l+3vmF2naU0CNLIKQ6PCXyniN16UmKiibSQI2KiTl9cv9QjKosA4jwolYhwnx2u
JUNV7zHE16Q4op6NDDTmbE1rhgGpEUMHb2eB7lB1eQGiDSAX1iC5IXqEipqh2tee
Cg/NFYsYxM5m22hdletSsGaPMQyvayl4rR55GYKOU6G6Fd0XH0H5b4x1ARnGPH2E
JwucDZ22CMgZgHpBMCEOMLHlj2HO728ZsV/9qEY9wuXA4oLu+Y3R4ENLlAxrBHtl
4lNU4fwvNQJ0ahDuD2QWbV0vkBwb0FPxlRjdhMfuCVa9ZwiRsIvjsqm/BofZr5YI
YRPHH6cztuZREYb4MCJpMhScWfZ5pe5GRpI2DDDbNZuwG5Pb6u6eMHsOGvSICL8t
x8BXNuTnNhYYpuzcb1o/6f0lZ2QOly7sDyHAM9MG9qg31BiypeFOb1csoJn1Nn+/
bRStb1IShy/iHuud9uyAyK0tV8VcW3XPWn7Qcuns9evNyoBbBeOfcM8G9mjYC5uV
U/wA1ch8F9HSmpOtC4mfH9GOlTJSj+VHcR0Rck4ktJioIHerj+hl6CF0WxChDj/8
UYtMG4MNPa2WGway4Fc6vCb13sqKEiINrnf2+nCqifGMVmPvIVco/MIRNdWZelqr
6igjfWFgpC1xa2rfrnitTc7Wn0JrMgq6xoUkJoRW45Aytug0RjMjqyF5wf/jHjqH
VpB0/y/4v2VbHNGtHnUqMMgK6eq7Wk+NYM+/mMnVrY0L/JwueSRwdECDHnFilgYP
+cNsNQqalwXphZW/phE7/kegbja8HKZ3+2NK/5dDUwdThsBUgSLNCj5tIDP2pMA4
uuUEUovEQ6w+YSY2thjiN7GNaZlVm85vb9chyakzmVcUtyiSHDcHgvxZtnpWD/hu
7cu7gleIMp7l3AMOkaXb5OsF1VaJbht5cv35eq7SGErpTTCKDou1moP/mt4kyoDk
7LgdMFzAZDp90eEZOr6iNFPa5eO0lHDJfUrYPf+qLlOOUbQo4OwWir29AXdlVyP+
voUQhrHhzyOHXOTNP+9N4SzcwPgI2rHl3E49rXkpjFKj8FSWoxsvi0SAzj0OBOc6
lYMdsL7avLAmvVk74qTJuHI8GSefwlaz+YX2EMvYZdc/zpowtzlfwWmxT3n6YVrB
SlqtGstk39IEYyq/W1g+Wmc0iwlnV9TYWzC0Ku/k40fkcTVxR0VO0CsBMIibaDDR
5hR+XDjkxJR5exORFjFQ3LD28vOmfTK921l/bYBI7jLJj/NsZ4LuKFsYcfVit2V6
7M8vB0pI5WgBYQdL94PIOhpvN4YvJGEtPGDBOwXNmnE8jwlwMUvJtq4sIFy0fqJX
U18k+wJTRDwfg/3hmPtM5H0sQIVo0WSOll9apjAlq/O5AbvZTSjCIY2JKOF+hMY+
7Rj8Xzn5vAuZ3D0qqz/TroqceB6AaX9QRTSbzof82IaZ9aoIuK4JYkhyxoaVb3aM
iuj5bhMquxQdAl6OPSRcbf47tFqnUcL5RHRZIUWVxI5hKRujt63OzsihhDXMMFAm
Jq7l6yCgUujCSI9TePbJ8HhFjxmc9xd9AeTrrxCa7FWIIR4NnZyfVgLJE+xf0Gha
ls8pS67n70+K6FHRclIeN5MAwitOfgimwV6QMptfB/rH0tIb9IbNX8n2GMZ35ysN
YHBQDMi0Vw3rQwqxZMhaJMw2MVlxzPe3D0dQYTo2UVUWJQJILmkwKyN2YR7nMXf6
M4v8JAsgc0kK60tFqEmak9vWl9vHEGVaEMb1z1VsoEmHNnK1aJM4yJcGV4bTzZAF
ZPex1Qo/w5ohUZ9igsVmLQtMcrjFApnuELSFrOdFdJxKonjHcisFCE80b+Ri/Ac0
OostWofhsl0kp/NYKtkH+ZQ62ChUP0Ia2oRV3M2NgIg1Z6k5hzlqqgI9fCmSvbb6
h38nnWqDHxLMK3ojp88Baq3/3Pg6dd+14g5ueO2jAO/uA+feiy17AL+LWBa/xbaG
dbH7IzsGoF6aO61VtlactdN5KXMdjSwDn9yosDGiQ8GosDfZBCZnU24Bvln0kd5N
PMtjMwr6VwGpPin4iRN+Z0LPP4eGCZlN5LmDBlKiM/g=
`protect END_PROTECTED
