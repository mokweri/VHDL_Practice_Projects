`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcK2sTHrySmRerNzsn33Xx9yzYPG4BONh3+CjxInreX4M+KzM2lMnYW74nqtXoMw
b0YWrylNbMv5KbVnBySfprvT3seB+wf3LFYYPqisd7t/Q7/Isn0O88TlxZU3s9gB
dTnuBTl5kwV9axb68OuRRWokqhY97Cfe010PINR3fQjzKsh3iFKQRWOLOH7cMark
uIcK1bis2Wyzut86aqbdyBN3EFyV7/joluTWQJlaIE5ZxtS7GiTkyI30fuEj12hB
za++eUq0mNwzcGr4larWx2filL0j0Ktx/7z0/pVHA5OOJvDWOc5584i+luTAYy+i
OtegXuG6uDG47O0trljr9qmiN3wFCVMNDvSAkXjlji5+BHYypXVfyM/d2/U5gr7g
MLeEO9y0GZ7cIk485ngB5YyXSBMPkMBQ4u19veZoAgPZVMcS3Aw2tvWrtnnQ3bMF
PUMVFRKYDZA9eELkp8nEgm7dYlgMEcQydrMG3aMBn+FJiOcbQ/l1keJMa654F308
7gNOJDIVMEy/zWf+5TH7nvBYb6YdAToIlSFqMMXT7pXQ4EEzTrAMGVuEV5oOlJ+y
msiY1XDE4Jyjow6fk1ZrXg==
`protect END_PROTECTED
