`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9YQojH4KuKJHBPTxR/6S9WPpBZkhdqpYbsgG1ukyD+8FLGvmAlBRDBcI0hximUa
G3YJDlSlf11K6hGnuBVWQR5ydpkmq2IeE6bX43JT1bUaPVNw7qM7mxVsnP5Vko7z
sDzvKUIRleu5EEBgB1lO73mQubHSUPgd/FSHZX181Hy0IVkuv5XfXApKsurJFhOe
L0att5u+FO4O/CBEgRB+W0JabqO+FNmfSRupgbUa++RJVJ1YXGfSAZh714AyGynD
f86WCB+7ViQiWjiVY84JsXsMHvM0UWRnBjO5Du/tWP1MOb7IriKs53d4iz/qWXpl
YxHXCXZTSS01qHaKzlGm1QA7H9FYBvaTCgWf9eQcOnP337adzM5CZqroJp387T7y
NohAKbGrD83ZFCbtrk6mojpqRMEv5XNTFX7fOcoluCfOxoOVPbNX1FizurYOFfyg
Std0ICdedHODh06L3WDfBea6xNXk6XADP9fFVvJH70gewlL3gGF7CP+oy+AP2fYD
laxom8O2LAlTN91JQws7yTrvW73DvHn3f2nqWgBHia9x8OAN7AakXrD5qrvY5pjS
6pW4IfZUai4iFwfM//1QtC48GlfNnYThalEPJrfnjM2fmvMiJi3R+GgRQBPvR2/o
5A9WZO4ZGuGzcvOfWtFniSJEz+BBAm5iYMPaAcodLdytLjfNxx7UwjQlxlEVletP
EWcJpk6OF4zn4mwcR2EoSM4k3r/na/Tzbvyy5AeN5PeB63bO3TYhsYcZi+he2Dmq
+yiCQztXLiNCjymPt6N8CS1u9+d1oPod+1JQ2ps96uhDkjhENxPY9FNgJy+Fngv8
jXTHvbcx90AwCgRbOhBtl/eRwJvyuxWvhIq3adQmW0FYf5IaEnLNMVF7QYYY2Zjz
Wzpy6KycLOD5XnptlUcyvzihffbmOdtnjRM8U/JMD01ya27swLTFGD/prQH2pPCV
v1D/dn0IyRnRzUpXT/y8qyVSXdittlaWsYJI03cwv/yLsfJ/ySGvyeIsOk/AnMq3
PPnp18mkePfbeLrvQuZoQsyjSwgG7dxsqnLMMUqLxwxf3Ib3jF8EINl6uWadwbcw
tw/eaF53WQw+pViNosIi7pnYYYXsiasLIbbf8fQMEHdCxmZ/XRWvkJoW6BXYEL1M
xGsmPTSkijlooMVz1UIsuCn/nxBO8fwPvvRKTeFZNg80aQKRyUJkVRMRclzO+NzR
JFVM9y5qsQJhOrmQ3u3qpBkScr5j+FNcQ8jfkvJluBOmhJnN99BpNv5O00QcEX5r
ir2LMyOJZlbtFCniVEuS+xBOy7Q5UlXqASACENGyb7VlpY+OTwHK1GLhqfRBBWYk
jhPSN9SU6ZTfQUO3AGt4PCOeJaQveGhVsD3588+ArJvj8f/ha9zywZL1QF1bq6Tx
zuk4iYP4m9nY4PS0mUap7GLyPMbpFbFdKLaswApLdkQjlxp4sI1CmfgzvTueNI4L
FRw4ZO2qE7sJabcS1/c2eqdYEQEL52qXA4c71cFF/ZkGyW7NiI24kyRwAG+fgE16
R81OgMRSao7CoB20tpWD/VU/RXHT+5st1rN1krnlHO2R+Pb8XmICNdCZv5Z2/L9Z
+rEVurgejkXP3LIAK7vSSQdjQw3lcS4IYnR1yI4h/vH7khLCenCIP5eOGZjx9ve9
QS/E0BS9ioyQxQuNa160TYDTu0/ppaYI4RVYnYmy59G5Lrd5RebOkPVyjZI60Qk5
bSJc0khFA3+P3UDexMOCzO98Thgd9F/yuBSV9OQcvzWAZoIkiL0GrCoZsNsONIB9
NLdXeri2/mU5kJ6hDqEpPb2e5wSksGJHin81OUp/pElEhc37FvcgZIgLtOAEzwFd
smiflA9NJhI0+ZV2i8Jj3L9gUCBtFLC1A4W3WJSMhj7x64VMivoqUxbC131QA/SE
mvxpcSQAhsNGY0kRS+Ree/qRuRlaPSqwJzO8F9/RdAqJ9FBtDnv/pwCp4ikXKENF
FUxHl4ULepWzM0GcS/0gS6u50QZHQnUilsXWd/ZbxUbGg6FPCBEJGklzH/qotGVn
EyE9u9XuvdCCKHI+h0vqvFLe1MLpyV9gVDYnTzOFRN0yJ+x39dAEiETcWKfZNhGY
Wxkp26gN6VtTufrAQio1CyiuvvTgHAFSo7oYiN9CytBIVUanMlQfqOS90tgUQEBU
q7Pz3lm+keJLMDOfwTypiGQyrI1iqDUvkJsCPik6DNcZnnkFW4dU3YPmVDlJKGw7
+nBPmeJCPioVMwnTb2frETYzeJzInd9b2D+NPsO+topxSHJlWdEtmiBHLngBMHOL
3bmenb1Wqx4bpRYVp4F9aRgtjTOHB45eNsh4/NumaRTcViZyOiNEudeXOotdZlI7
n8YY+ePlMF9k20nC7dFu10PDSw85kjw1GkmqLDsTTStWd9AJXKXFJVhai7EZazQd
KSgGy1us50NSpX0QxbMBDHclHV0wSZmvPecTdMkCBZs3cU641vTbV1sos0S+LLHh
ASGOvUUToCYjsKDTq568bxp+dlRO3sHyKNVSbJRPTs4bU5d8+mEhpsvTP/7465Df
+r0EiFO8mdTd98GPjp37iKrhGSOsfJU1HFoDDzFD6T40klK/IUfA7SZwplWiMjvV
3miVI8IcJy4wSJr9uOYiqZ+2GFmrxgC0Apm2fapDOAvV2ek01HHmF9qKZA6N5O8H
i3/60zToWlB93yrQh1qtRo7e/usLhiR6KANX75hB1Z12Mzt77eu+hkumRAwK9/6R
r9kBSkaUVuXBiJPRykSRlrmouNFQfe16qzC578kHypdr2Ly+egU+wNtZURwG8MGQ
M2D7TfGYytWaeQ88f7shlaSizOS/3In75VrefubKCpz4IhSCqLUSk51LmNLbrVJL
AfYa4lQ83SbQT8mnH4qg7uq3wTkvrUXneDpZL4PA62obULCqnUueF1jtvRElgxWC
E3aa9mVH6MWtkJMzijW9v4aKhvxKFl8y57pWg6u2iBRawRVZZZAhJ0GRjHQTMYlz
whsX2QflBLKOh/mqmtLSA2CQUGxaf+T7YJEK67F5n4Iw4/5Y1boetUUxqTl+nUVw
NKvRdKmFSy4mIZsyKLImnvGda5HipPczz3XXnP79peVAsyhR5XiIaR+bKJ15xBVA
XwzQRb59Vi9N7RwWdrF/SfUQlgoS8aJCUCULvlQR+puHvtn0W3WM4h2H0ccZ8cOA
pDj2lK91ITRdReO+dOUZISajZdjgB1+NYkJh2bYnNAs+U9Avp1ghWLLtZk1R2mGd
JY739UGhRyCEyyLYiXrL5oJAOd8md674Ub1PaT3elRHy4UribcBKSyK1eogpblzg
yGhu8FWwAGA5Yq7RimGYVPMqgApDCxkKN4bX7LbciW2M7RyGBKJC4DX4LOQggkNG
0N6CJkxDRTkasdSENy1eAkQUQhraHy6Olhk16LMJNXBRmOlJyTpT/5DsAGtDfhez
PAOmdi1g6GBBdcJ7vtMaWT1Q43jdyJq6XEDiGp8R+ZbxPH6Ol57yXAfCBej8Sd3D
UCUrE3kpk6BeMMmzu0tsYtpbwPjWaufu7h51vZyi7jNRyFC2x613Uo0xE2atjffN
XMtohow/LP+tDCjHHh8lGfFrBRp5PSJo7YbqFE4qCI8aeR59/PQIEHWbIN5QwndV
gtYG5xisWxxG9zJGvdBXwfxn9hnXw3xY10aCY3+dqo3mTM/skmrGo9AOi58Ljxsm
vOKL+jSCyioAK9MqpLM1Xw==
`protect END_PROTECTED
