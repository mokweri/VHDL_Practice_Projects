`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pSlWpn38RHWpzi/iZs/bJZC5lS4L7sgfDZOZtjNAnjJD3yrlaw8auE3frAWoFJNd
5DSieF6zSSmkxSmo5nihbB7o/P3iz5OyhopJisJl8jp/DFlk0g1BzzPOW5r3QCyt
WaqBh/O6NskGATnDhtOg1AsvTyjUVZZgpim2sE1lnGnrSAMGthlaOd+x1Oio6+Mp
rh/nogPTCFfh5UEIE/T9iVolQg/vxpA++/YruFwmHImW+O6RLyyNa+yx7Me6tgXP
r5J4Pd/zpKc65rKRzyO/psjWwi6FM8LVf1xio0Jyaa8BCKZYvUb9M5H7O7fEfun6
PF1kL5wum4Kc+6uCBHbRSrdIf4r/fbIVTXr95mpAj3EC9kFGnCpNeYkQJrWW+27T
kCcKP40BhcJXrBV5SfbNvNdAtoaUCfzQPmZ6INt1u3CgSm59gD7a4HUINW25nwXX
Mrij9b67oXnRe4BC7fcuEpl4WMJon/itYh1rf6bKIP/KEr8BwNSBtERpbnEeGrKu
RX+QSNSVat66mZcM82lvxk4a9M8F52nE+i59iaBVmquMxU4J93LDS4m1jyNnkWwM
2Dt3I3nfB+RsQtxDtbl+g+7s7aVAoaEmsAw9lj3ZljXbEyAPzpBPeFeH3XyoHS7Q
3GdWFhPhvMz3PG5+gJXxM/V5nlYklBmhqZB89i70WkZ6gtr+4iJAMoW5ymjiqSqw
P5OKL5qT9UT9+jWnDzAGz/Q8uxQvZBmwTL9qQaGy+CZHp+hSFxSNfYBo+XHn6edg
sGz2hHSf3s1S4ksMj1cjexPX6I13Xzwfo8/JH2NNXGh3iwC85udWbGlrewtUJhiO
CGOKw/qQkxbtTdbhelOYJ2R8Sy/tkocgvajTFZd3UMdozXrKzUkLtaNrYfSk8daG
GfHno/Th5W6mN+yh33IzjtMEtLAMTWUhsRXRKOupS7ASDT98QziZOhlrsoJobsPW
WbbhCNO2QFzyioRsAroat/3h92r4zurilzCZWY+jusplMCp/GB2cVjGTXeO9SDGB
4sovB8XK7u0O9TFb/n+MIPij4nHInRKLV/F5u0/sPtSa57rEUECigedjlnhgRxS9
KESgsa0Ng8LM2Gd130WVJOYxzuDcXoq0+L6Wmu5o1A2zf7OcFe2AZmfUrfsaC3ew
iC3TV6YbePmoT700VlQm3AsEC02X3gT8x41gmQBbQsQFAsAVPuS8zPGaXevX6KyS
joWZuKnOD/VNCv3maOTCQhA7Wmt+EWO6uGJIDvbijqHFs+3298sbL/2M9h/jDbrW
UjJKrIDsAXwPojwjLYudhTUparxzv1R3GPtnjAdoyZmgxEVthQxxBbzegDIYsH8D
tla2siNcNXAS+TXlju7XoFUhZN7lDas//gzeZcm91nNnLQhMVdut0cCU5BZ0A0jE
t6ZJt5C8YWXbdyxV1PHHZt7O9oKqAE7Or2VT9k8K/PFy8HmdwZ/pOOqksGdir/w7
vk87hdqimsQTQNVpE0aTsxNoGg+nDhHs3ilRFY/Iuh0zUjcu6V5evKGB6UV26sMG
ELtFIsr75YrqR5rEHV/yd35PgQhZ44iSRhM3lsYXtAL3WevwjhK/hYz/GAROVeJJ
Ruo1Z61Vk/7YAWA1z/PbZISeYdX1y7OusNUqi4kCc+xUd25td9CWSJ4fNT2S9W3y
KCNPBGRd1zrnSLqNn9P1AqjKt1D6KQguWOYhiNZvodqLFqWllkJjvdlJ6hPzKbdQ
rE6Q91UZwymUVLhPh9J6yw98lv8TOBeMyWmE6wR4FbSZieYy2FoNiPBUyJLgHrNn
iNKckGP5Hj0DMalrVMJXubYALgJyuBGl71w22SK7GRmVhK5NgpjKoY8uXJMYrGR5
egX+g5f+xRWz4Zluq1ad11YNOUFC6jG0WMN8IpHCucwnFo+dDvmiLqXtYzi1jCo4
tTy0PZ9uzfAr3R0EDx6ku6hnvGEnyS4MowgFZvJS8vJFfN+IDSqxOOXKimWZ+CW+
fjMXc/a+xR8K9N9+CYnzpUeYZ5xOT1sraeXhbuKqbq/Rp9XhM58IfsZj85l7teXx
1BUz1FiUrhC8RqYk0LD8U1qR0sdaAY/g1GsPXyorO+Vyh+91YMwNqBGFkIUfw1FF
/tH0MaDlDhKugQrINXTo3VZZXrYKrwUgoZA39Z7wkfV6oiNFFqSKlt3BXNCQfmBX
5gEDJSEaqfiwgPhVcY920XPy+1xpUu0E3yUPZAxOgp5bdoGmoTqREkJHY9vpC47c
ZeBRtu5m6Dmt47BBE1krGbunFHfx32ImuF7x8pmRTHekPFE3Y8lthQGIDeCcF1uG
bpXcGD9QzYb3yitjXLWs+G+g7/wYbJ/C5zxzi+1MtnsJA8kk6PCIyNqPTtp1y7kD
W/J6LZzZDsFmU1cWRd34l+ijoFH4hncVB1WUF4IDSEd6Q7CpP1TQdij+PoiVIK4G
k9ZS0T07YzZTpJTgCtoJ/Y2DpWRrzaRd0ishBVDBDwI7o5xzCvBo46pTr1vdxpSO
nLLp+T3Hkf8svOv/hzud+Xzq+h9A7OMw5EEPOmG40Anv7JkR/yiNlirTZ8Yls3pw
JpsJeUNzvL+8m6qjkfjfl6RuRmZzg1Qe+j8NdPaocs3JM7uiI/bWkgWghSNwVDQJ
N0cQrbIEc8MTevfWJhygA5VBej2iA3kXU7+mdLr1n5QTSqghwpHpUz1IAIfUwoOz
CydymNxuGECEPCZMeXJo+xapl22jVUw6/CdP2cUnObWfqgkNJob6gD9hg/1bJ2ww
ETxygrEheQHfy9tOzDrx+O8WGxpXbxTf3Xe8OzeSxphKuLj2TQPbXkHZOXOsUJln
y/txzMDPcZ7yBK6r3fAFRjYbF9IFG/LZoXZF14I8asaM3RGCFHbJ35zM6RmUix21
8LsSpQRxTVGmpe9mwFuHaRaagVglF8TP0PLQqjqnhTIr98A3YL0dCzohqOczF1dp
ficsIbWyficZTAhFcirTyU9CTeFOuzfCVnVBWafuT49yevts6Enea/s9HGvoeGnD
bdvz+m1q4t1dmRHvLSi2yNOmRLRIGYAoVH27LwTVbf0zeC0jtnqpZJ7EFpJ89jT+
ofoytf1Vn+q6v/+viZk+oHkf6cyH5mBx9mB2yfhVq5rEls467GXeKVzi91mS88Iw
InBT6zBL6/491fpy23EdZ6OuXjjKkS5wn/72tywx/UA8+n6WG+5jK+IsRF2idKil
33MdeUlV4KVQOBepr+AD1fjqJJEjJ2HY3yoKjU1TBp1mp7XFQTUZrn2wpJF2Fbu8
Z4PnxpUXt1iPI0eEIUu9dZPM1ILIL58rQJJsNVHL75Fibz9f3nzPxkFyk6iS/nMS
/pYkEBTj4PbIMJG7jqma1nddVtOAn2SDgzaGrkpLgZlOS+S54SPWdFndJ5luturz
M+ax8VIakIJTUJFrpPZ4xY78ddYikhV2vtQw0CjMgKl/gl1DYJHu59+4IK6fR+U3
wLXmFhGIvL3sFTHKrEKblw6G9WQgdu7S87NvBO9/CEoMDxyOiGG+6eyq8r6lSm0u
H22rZ/cxQoGABr4y3OkYYcHjxBOIrI8JBGDaCNlYA9RTQhKDWEAkje7p82vdUbj2
YyKv3TdPDAy0J7gyRgRqwW/AvOkOtQ2KcWuVSHm7KF7Mf31N/kXoUazWTR5H+9Wm
aUeNqwiEZmL56NBW2HUPEIHqQSYhwIYi+ZLzHkAku0Ek8HuSNzXeEe5z8I0gNR+u
5Swsn9BtkTxYs5u+829shkwdvhr23SMOTFZ7ZdwOBcq7rW7u7nzDKFO6Y8gbS3Dr
C0kap6z6AIDztdeQi4r/rUd/ZWjzrqv1XJZ2evx0YSj+j3oFRhf/Cjxx5cxjrUZb
npWEYnKiRgu0DusV5RuRwUPk7/MB4lPt8MmXchJTwC2zCDnS7qyr/lnB7dvgaWOx
rF33wJIKxXUqTqjOems8jl1bqVSQJ40cA+sx39BFCYU183hrPvt5KihH4L1z5aeG
GLW85daKipOG38uWdY3EFqCfjRyLzbqkRO5aAzQbSlHqB7qkfwDhL6lTUk+p2A7U
18CTSP3TXb44IYS99zf85pmjdzoVunR2LjDkpnWRIF+tgsHlqhRvGkdhwBtrltvW
HJ2Gt7Ep26pVNIacfbx2+/x2EPiEJBpqXNjQ5xwjP4kSWNQ6flipcnSYiOHT8CAb
a8tWzaKLkfxU/R0jnO+u2H7WyIbjnpkAIJ+OGv+4toMKUb5pFU12JGCns8hP4yu4
dF3Z3frgRxVrTvGzMEqwBpgjfQ0D7ouMKtmgLX+9Opex6KLgwSilOGqwLSrk1vq+
CzLKc2XRgJjDYi58guW2oxjwLgayGpKCUp/rbm5GH8tUaIRHBk39dDAgrAOhWba8
4uHXCVTM6FqMWhW4sh0sYeupxulV/BrbByYbse8idj56bJKl5neSAcLaataBQzud
l0zpZp+siu8A7rB36el6/P3sbBzrQjsB0mVgJEowFrq6ND7HMsMAcbCE4OBdeSBV
v5lCNMda1yYBRYMiQElta0zKVJZayRZ8UXrZJXd4KR1LwZ54nIHXiuaoyDfhAYWV
xDG8slv39S2JBQQI3jnlAewfWk8ALze1mDvz86KXSzg99KH+gLp1+I7UHvhEXEiS
x4dh3fa1ZxJOQH5iWJo3HsrSOsb5EGoQR5TH+dReo93OyiFZHFmpEiGzqxPulS0d
p7Q6Jl6jycnX19ac8WweqFsWDUM9icvTR/TA5hJkQF+VCVlHKc6p1wLcf7CbltYA
zXGOlMXfawLY6EnAt2RomMtVxe1v5y7Gp3Niu/ubnbmoMlprnG2yg90B0WnMaOqF
vsnJpKynEWiTKuu3bjJCLOBYXYvtxGoJ0ZRY7kdBXgYn6dh1O+E21m3zhaBkjf4Y
zscK1emtgfTLEPC1My9iuNeaXIjLBkXWFxl4UZnG3VTCDcCHbqscCd8OOcwUrbsH
eDfkMExUenhWzp61QGb7kqsKfwv7ZZF5+7gHj0VB2zxxb0iNNZJ4IuCqDT8ZaFwD
3djCSJQlB3DIU31Y9G6hHIh4IHKpsFs3n1o4JHl275d+1TcxxksVU4UARtKXlHA8
Gl4cBtajp+AkF1gQc+DmkRLTKqv58/aWD8R6UcBfkrpbYB/F72BnjOpjpXpRcIQ6
ACn9CGnUSyWHPrVBjQaxqaHrWLKIHcUFNz21Ql7C07phVvOA4wKoXEtwjzAnX1a1
d1yYTMS3DTOORjP6BOBmnGD6oKurG/vBrLdkzdnar8oTmQTfkGHCe0uoGOEJkDGE
5BEsek+iZ3sHvStEKjKdz1Nm2ZqvgniX1IVT1fW1323Hk6gFOGLKnUv9lleC99ch
W2wDK31mZ6mkQZhNSYpl6NjtvyjR3fgAc3Mesv8/MTM71t36UNS6Ie7HmU/pEWZ/
rt02pMkKNjCgLAfNXlwVhxqhIUgpN8SqEAISOnsbNsE5moevu0WFzin0Odq7r1B/
AzNUstOCLI/rzmOFbo16CiXwOLjVieJ9rqC7ROIvmd/NuGJgaJUyxGnjOBGzdX48
hmYH5ewerxD9FMotLFRrhTPV+FULEr1ypv4CbxhRmP6LOBc1dozLiDUv50cQp/r3
Go4kPDleNxRUf3Ba7Aqmm91UsjpbGSvMf8/gcNwu5QFDrpbDwVgsTkjxatN4pYKF
NBbWtu9XPpqABSSgQTy8LMK5XmCcZ50WDF3ytVqWeWxTERLESyl300FsKBzZvUAr
eOCKgJgg0WxyFvLAuiEQeq/YOEDCjipl01RCngCMNW+wkO80J09yLYtst5+U62OL
a1kA2ac5rvWVGqJqVqYLtqN93YaJVmd9OfXoE0MRBYbsnsSEXgYhsubf1p2WlmJH
iwax1OxQ8XiUp5MEnYKIlquhJLowK3i3ZkG3kElC3QRxZoF/TBF6GIDwyfbhHwyY
Fbh495l6ruJ/wnH/lTuderOyzCZiePt63z1kpyOhIRK5924IW5B09EGddOAQQ74s
tODsajxvJIwowqowoFfiTT7Z85l6hhckDsNdVNqBHHpV+iCfPx6ks/50miP8jah+
st2VfZ7msVad3HvIeRGr7EU6Ufww7WAI7naQ2JomDnbCcDAIhY0AB57SCQWjBoX9
t8fUaOJZ48OkzXaRrBfW3OeO9NYu8PVUpO3k+lmy9235ocJkjRv5ffbMGwuKsdp4
PcX+hkDCGrKi1MyGB3sCFfPHxXVMs9wnNJTlSOoGtJJwI8Mbhr78ylRmODxrXLje
ZRGj1cBWRUiA6quVNRK1NWj4MW+LCQOUKN/YgQ8MMXhwlOfBxEau6b8/fx7uFsNp
nrHjvJGDpgga/P4w7mcB/KdqiQxabdWZAdbcJ8q9KvVCgGlfRLq+ECmz6YWaEJrP
EBFSG9euitzP5/YkHvFVviBrPPZ1dXxpx3pUbmXbDUfF4EQWA5FUIrHuR1F1t6Yd
G56jU6IR8dEhnGyOBJTFBWiv7IhjN52Hg2l+hE4VqL/Ofy4gLS7VLs3LPnvZ7qNE
7EgUlDeJ48DxeghUj9aWxTNFC/6Ml4q4ihV+YVxYuv5DWHZRf6aeC4g0AtaTKdDO
Kq7jxnH/HDBlaQe2obaEXmf7YZygTyEWUEcHdaThclSxDR+fz6vkS99VdavqLR2m
W8y9iGd+Pf8FkwMb0x+W7QxT7qe5Cug5qvULnFdjSMGIApcqcX3sE9NVws30IRgw
zmGdnCvLNY1N25Adc65FqCMD3kqksWycofDvu0vLS3AtmdGmh/sPe6qKEL4R1Q4o
/artMhpcxsog1IxCRpaZrjqs8NSzV0GmF/+v9FLxCc+BNBRiXTHaaIiTnnvHLCzu
3OziC/tYvg0R5QGCdY7ZYBQxr12roL2yppQtrR/680cxER3hfDVsNdBIxYjSIpC/
AWvUJCqOIOU49ZyEcQQbfZrqAe8qfuw9Amo4D/UIW8H8KZBZIvMe9+IqqNytUhJJ
+QBRLn1Ms3GJDVFUH85e1HGM5MecRBXG44YqVdaZpurPyc60fNoMWeuXETCDixSa
r2lKW4uxCiqyikpDj1S79mVQxys1wtOAsZkuxrqbBHnt4NJn7/bItb/2WgEQ8jhn
3BMzMFKdC8iPl06WTwY9Q/IMzcMbbAkYGtSpap67yZZu1Yg6l2LX7Ie9C4zLwLBl
oxgdxzobhmDTRHWz9oHDCNN2G/d6TaxEfQJtRSguEzPjGTc5RPbTe3ZX1axxVf5c
2Rd0qciXjreQeFraZ3V2a7hMkIX+Goxn/6BB7AUIRKNmtn6XJtvrpoQtqXJa4pyH
AD4yg0Hksf8jioCBqo/rNtqqU6/1nLHc573RyumXhl4Y1vgVEUr5qRqBOjz0Pjr5
FoITSRXu5q9ztc660gaPa6L/nig8g1Ahj2lJrTTwGo1eJCAgVKMbW+jLjHCXqSsJ
cgZQTdJYzDmUaZqmKcUvbtOZq6vXcsF6Ci7axCJ0wQVsw8GQcwvpJbFm6XlJXaks
QBzdkjWFwMqeCqPqXtLH7yWu9lqLY3hgUd2P4OtIDLXQrBQMVOIr+c2C2Id+23xk
ltBH71niBbe6SxLSV28l2IPEfG7ukP1k3slXPm1nzPqJBxlkiN0jHAbmqzdYQQA3
5Jm5jz/hgiNJsKBnNhNqgmLah8+suiixjJI2g4rsH74QSpYvDb5DKxObvURJuk4m
GI626XtrJKThFoHh3lI3fSrTKuU7bS5qvxXb0eG5ZL0K9PLunUKwjN1cv/foloxt
y09i6PXQHVfp/P/0PIiSMOtejtz3F9an5ch9dFvmT3hU3l1CoG+BKxz1mupq5KWl
jg7APDH1QLH15ZnQpsd59P06QhQdj4luCqPglaZi/0kv3JErSgnY+XquUy6q2DST
OtGpYjMrFhr2ECErY5B9C80HztN+J+hCN+QBuN2IwvgP9yxfsskmlF/JQNKaVs+e
tc67q3yHjYlFWFzFaZHAanX8SBJXW9ul+znXaH03orl/p45EjyOjSBXW+g86x3/E
A7dMkXFJ+WZz4LbIukqwQjL629X/YfpNE8Xq6U9F8T2hZt04nrWJ/yBC54uIvX0s
BjbIqPePRlZNpjwROT8qjWSPBSoZ3NQN48pQN+FxoHct4mVKuw1D4sbIf71gOmLY
xCIxrvB05LVqTrNy8RUB470DFO840tX/jYqC6qo+lPZVYuiOxlopM0Zr1f/4IQxP
8XAwHZi/JXi/bl6K8LEUbcK6XQn8ZUKuLesRJvzfSwC9LuhJFdGVXmPLDzdUid1+
v40G+wkbnzTjb4rhjDJ48SMaz0HDt11O9kSS4XOhMPsIPa7dC5nQQM4RD6UMy/3I
2rCkKfHXQCJRacZrh6BGOefeUt2/aOujkilj7rQyOMkasXz4Z55vk9a2nuXdWXF2
K5mvtroOawY7jdXEVwJ3sBQEbC6evbDnRn7sTGftj3VwfiVfi0edzLpvocoJECqU
bwPk0jHdvVtuScL3aFrqOgmVBkolSu/Rnajg27PgCfAdB+JaM7lGnUhukA7Omkp/
CcobwO6l3+HQDyAlHGwN9LWjWz62THtjAlhWI+g8H+phJS1gbxw/XT4kAP9Tep2H
t+S3NxNtvvNacGhX2EIAOxkMpUZZ3izg7Si84Rqp90faG5Iq6F+PVtJMtJT7UIJT
ZYr5FrHTvDneTpT4HsL9eYFh0s6l3l5YSpoCTbcJCQgej2tcQG12tEl4F3skcZUU
UnaOxFlx6/p42Ep5eMJDk1fXkFq0/O5q4YjOxPOSHDZUx2PeqztpcmP92QTCJ+ZE
LTvAlwuFoikZeqKg64tEooDwTeHXpgNKqBKY/zvPznSIwU9WpnvqHj8nQq8EZAmn
EoN2GmDS8rwbYYES6edFe4dPHWrjPleTrIVeQZ4yy6w3AnsxyRN4SEuhZDwajUPg
jgzaX6g4KVvjUUbQXvnKNdadE9Ci5TbqNu1bQYKJJIJojwQNW+BMaceGad9Kb0L2
tvuZrQAWNdPwF6295LFEMCV0NHdY1rVnA6GtA1NRSSyW/Fewolxfjj9cNGpZuNdq
4hpKtr+OnCxP8LIZ1u8TZQpeCmTuA77GlzbrThHkuPJEm/39cYPuv9bmVo7RDNmf
ezm4aIzE0TdCXTFBLY45dCQxPpVk5CjrxCoaNjdKN675E3MTHFf0ETBGR6YSVjST
VKgsd9gJLza/zlc7CRbyhFXFEQ49o6XTvMCvKDK3fCsL1bXhKAi2KjTOJZJxae7M
Q940MG1708hKbgHHgm7SrK1F4IrMK9GVEL88S3XXIf0roS8khOILo4tGmULjMpch
c2BH+nDO2dWzgLRmX5ZzgI5kmdQc+OBtKezzphAvI6lxZdm4qo+GvzJ7CxFMfptf
cXDkBsR6BuXCvH31HO/dybUAHCo2wflxsrVJRSpEFwyf+kWf0PX3oAetM1Oc8ysn
UtkXXRFsDZrk31LwDxWXSrHD40NW9O6MIBkRRXQFWeDjxUZL0Ff2I4Uh6xURJE17
W5rZc+7t5rVvtFnkCC7U7mbDTectbnuP9zlyuQo4+aAdYA2Tbiv9Gjw0Ci1LxsHO
Gr1qFwXdZODtz7HF3VRQHXXIw3mICiiUREvsUl0kTtOSGXYCEqu1xkOnwMY2SMhu
Nnh8vYZ9HfuVTa4qY6ikxhdo1RHKYJ84bksrzUhx6/NXkqUcQTPq9PXgmg4ZAb/G
BGmNO8sJtPHcaUj1Owqtx5YPI9An9FNYNcq2g8j9n5AuzpUScfWCvO1gGCafMwMg
HhKTEUG+8W0fJlKVu2pQ7EkswP6dgxoFkxdtBly0YEnArg1t0RLISKmVKH1oHkvS
I60krMrfWhMmYZsVW44coIz035T9HfXWU1ECV1gdBquyBKWm+uYzj0XzZQHztlY4
De0CvKOu1TY0wldf9pu7V5oNOTXGkhqbIexcw0WAuaXH8OvppX0wKZomvNpT3jbM
kt0yvxNYxB/RZpZhAmVGyJv59VDK5E7FXMJ4OTq91vwMReeBFhOBonMasj7va9dn
7pDhl0KGC+lD6aUk/qpFYcbq6KXjpUQfHgVNVWT7ssQT9LtVEDC1i1MqG2e4OBnT
KcalcueUetA0a8FqXCN6FQ6NS0DP5fHotGeETuuvudEi7woHdUzXi+tFSrmVHc5C
fEpXkELB6en8r9aEIi64pAdk4ddBZs+tkuMxEXKKVxUqVcId2VnSDar80NoiyeiJ
wivrZBtHjTyHlHXprLjDzKwo/h5SXXVLsZoYBxm2uLwMb4I4w/myxZSTJrTiqmQn
j6qN+7C10N4h8ylNh3EOMsEt4DZECqktQHprQOHxyjacVMm7gMs7anX7bWXoVuv3
bA/lO7jRVgebP6wB3QioRr0lIIXiqKUSjkAYq6uZ2z95nDgPkIv0k1B4bdmvgVGS
TYFVWAYlJc1elkYs07KhRCiuKZ81T8BnyVO2Go2cfA69obv23pHVLQiflot/dSkn
iMVmOM+s3cdoue5gVqF40FmFMHQfB53vjZS+ttPwhSHd4TqihdPqqajKZLKjbU/3
0LtU7NDAreU6fUh1lSDkAurRR73SYQInxIm7pn+ABAmlw2I7lUwnJX22oX4OUNy5
iBRncDOCPmoQx6q36r1syMXr8qvHdm5FhsHkGZP6iAJvaFbQDMTpxHTiZVu0J2Nb
Ig/bCo3H4VNq2QHwkkKf/aKEUPRiSTwsCdZSX6kAMZaMcRcVURc4pu7H3VZgovjk
d+QaaZklhogz5kryUStFgdaDp+pww/bc3BAEz2nHVnwQSQPpQJy+f9oolZeyXGr8
CZwjW0gPwqXZPIF63v6tEfnmS/9YKBiaxZ4ihLZVa1qVAvA+QS8rfH0abmaTq340
9csG7a5bCcXeJSYycvKkqPR5tvJcHJ1P5naSsu1Jjia0nJWYMNJ/8nyasPMQJOj4
LJm18oza7EqJExDSgYrAuquEPI/nepMp4Pk9g7ArfH14IrjBkVx8anD/tqodUFle
s/zzlGluYx0fJXf1y0c2TOk9gUye6o3ePypBEvtiJxlpzMp3wlYSmNLihDTW3BqB
y08TdZTJMxO7VWV+Io3YqUyldM7GgIaJ+U+fZc1p2ksMZNfG1UxggEGGavzVUGtW
qFN+RUJghwV2uPD2rP/6x4IzL4Zxn5kiTwKPCB6hvYw1Rl1bhdS+gvZS3ZL0MaZy
EhTVT7iPYUJat7ctzT4GAeJfUMAB67ocO1sIaBwV1BFFmLC7xNACgSbj68GX+vmY
g+o7SyLKaHYs/6wEb8uut0gKsE+EkFZGn7HNo+hWOBW86Jt+JUivtHfBSvMsjQQZ
lJpYu3Pw0CYLrgubJm8q3pjn6kXS7mJYRpURq07QHn0D1iap5o+hHfQDdXdzciRe
SRJkP+6DOOcWg+EgjUzI3QovJNuFdW1wl7tQtya2RcSaSJo39wk0Ejd/G/8q/wvn
pbce7R0xSbOtkczXFoZKnmcErGqSQgppLeQJUY0+oo7I86fquoUP8jQ63yITK8Ht
QxTw2vlH8zrbvgxGBE/+ZZeiCGpTFKg6ruqI2hb0HyehAQsR8RHJtFN3bYBt8wQG
XqNgGs5RFJenIHG8mNqHFu+8rK16cM30uRDCe3EO4Lb/wTUxG/B4E7AqOTraotgy
JZUTayHQ+CK1yYz8yPIuHiU/gn7d90nshza/FNeNaoIeYpSOnHCvwhIgylao6Ohr
j2RSOxGwWoprLPxvrL3WwvtWDg/DMc3l1z4zJopbO/bLJLz9Zh6H2UtFykRNbWBD
gMvz8tZeBt/JkyqGq3Ummwyy+f2qufiGLJeA5YX9pRV0EG3cTbTILTrMFl4j9T/y
QSLZGLJAveTc/VFNToEwrN9zDYL2e0CjjQRghACV/HOKRpKeqlfq10D+Z40Ykx/o
XdAMDdgNV3F9CrSo+wOq9yGi1+5rc5WcMxdIasY2uNkJEyv1S7+BfrG4ijsHSw7H
tvD6bftpyOSOeKqXh6VHvKsmxbgpbEZiqLHYytQQiop+jbj60SX+m4KD0kliQusP
AZCRbXODEP960IFdoLoiUMcvOprp3EhEj7MPFQI5WvUwv4ftUPg0UXlxHiQCyKJW
g7qjB46q2nkb2RcNar9mI345l0bsPvx26yQUF12pD/Mlwwz7uN5cMEx7tk+myFkU
wXnmfxG8TcG9NXZxb9RDaaIQPyaT6GHBZ5alf1tBbZabrJhiuYVJ2eRwYTrzu2Ih
ZP+QU1jDJzLCfXVNEQY5za7DDRxf0wnnZmkG+ZTusSiaiUjp5aakk3ffuv6E06OX
8B0Eu1/ROJ/dR3GNO8oFelVAUaFJZCylqUGkNWbamOUdxL12XQYk8+3hheq3zH5c
jeGff/w/feAxmFyASogkNiX1qQHHCunqIX00gg1c++wOPbyxQXs9RZGD0V7ddj3L
gUnWJiVeONQZv8fCE+0WHMf6T6EGzIjBBNny297Dn+Z5CVHef+yI0rsVibyg8vPE
U0by0rpT+Gzezv9VVghrGwJj1PlmBxQ9G/Zmskvi528sbI6KvWxDk1iqZmudiLNf
j/XU1Aes/eGOmim3qRaWyX6wUWx0vb5WXrNzxHuIcX0kdKfevZOEAQziTWyDzE1N
VBLI0g0G9VSZ8Y8/yOWMa/eRCr01fCOPghB42gz2gzDWbh6Tm60ZsVK2sYw+by/Y
/NvvGZDob66JylSLh4qgV/x7jOJ3Oyl2xZte8y6aX1O74Jfh0o6HsPXeR9T9OsVE
UMxF/ptyxaFVLCDsA5mmmLzn37aKR7/Kn+hgrECTtvX35kTBsX30dR47pXazmRca
Vs7176bAStNtcvUvDjD5Da48H9oXoIkgZch95YaRgSbzyvL35mEcr0banOA8Ck8h
ZIyQxI31ylBP3UhICUlBd0pMdOqMSKaJ+x3qlvSrc/z4WqWm9INZJ3BgcfK6bCO2
vESVHODNee866s8uJBMNlAhNUGwyq/aTCTuBKC72ekCho1XQTQmvCRFwSwlDLBbC
GLZFi5cwFDmKIwCOo5s+cNiRcgf+Utmc6HMS6Sx9ab3rf5oicrnKkz9myW+4pkGH
JGFAXqmcTscnG3eWARnTHUVJ6mwr0D73/hnUuBUhjx5KwINiOXgcPeDg9dYWRNIg
XAl7FHEBsX9f870LmvCC628zmpJ1cfAVZFVn+oUnLDwcnKE9BAew4B4VR+3PPYJt
kMGyqb0idTsOvgcR4390Dty88DowVqIt4OPLCL1SjefeMz+QkYwR7M0KP4ZeHw8b
eDCgUql0HnSrPhzYl1n8xl9D3zOsGm94pI0Qy/Vkk9VYvBrTlOPBrGv8Q7L3SdjA
dVxtYb2CAm1G5vBUWiWJN5YrC1ElFXL1drqIsKxCWMeN3i+SEVouocBixnQxSfvf
z5JQS+cSm9auogf++9qmrisNZs/j4JaEg43Tb7m5zRc+v5Khs2Z92O4A/bGt1MM0
DTg3g0felT1wInBHG36lI4BRFcNy8ZF65tiG1h0gzMGBu6Xwz8+kUrxY8AbCsBH3
B4McBAHzdV14hPqtiJo2igQohhCVYch6LDLv3Kgw5pgtg/URG5GaatQsjtVRWFXa
GOJbnKxbtTvy6EBGuICHICWoEPKpeCcI3WRneXRrCLhSjoHcvsPhcCnsGqgGVpuE
vNHayRDKiPHC/tISdicTkICqJYR6ZIHgET5BKy0RKFkJUHW/uLa9m9PI4+7oHoxu
3JhumklOyqj93BSPb0dBuEc94O2SK+a3v45iyWxKSx0YYp76cXNDoR9gIJMs8HSk
H6cEAwVssO/zA9KSGrvp5mn4qc5Ry7QcPrC6pl0GCj778P9loZ6y8FVrl+t5jk+7
XdrhV/QzFTK/Ljow4ImGlFxPv1xK7qDIYJv3ig7FKxgzOjvfGBHYY2j7bnwgg2p2
wUSH1EsuilKZ+kN3Xzt9995jbKJoxSP4Tl5ty7zs+w6RkkxIqheICdEh8mJbyil/
N6XECo9wYeqBcYpz7SkOWpGbnIqEsOkvF3sGSmcKlH8VuM0yIVy1xJQr0U9DNog3
bmsFn5MQxncyJsvfONGchKplkYj+tZbSgSzt35Xs91QkZS+yiXmI7rntl5TOkxgX
EstOHG7X4pe1hxSzjUdJpPCSdr6+ICsMzSnLjM/r/LrcutbxyNL1/ULDS1QdoKMu
E73oP/ZfmXFzB7qX0HmO7gtBjmHCPShI/x/V/wH9wMVdDV71HKBuH+XqhOT5o7Jv
fvrIP86ODi3OZP5U53BV0Ru2GqDQ+GCmIqgoXZ5zWHEYrm+44XlHvwF1zG1hRv58
/xJx7GGrL3YF2iVKu1yJnbwy65OKlfvMcyiy4NNlTJwqBZJfgDWyaQfF8SoD0/7/
1MpjMPCW/XTOkwlFhmTKXIsVAO1APQYRwmLmsntwUQMv06C9ibF+ua1zrJ904n8f
0mFct+nxqGJrdCpdDW6UDlPgcQzrS3kYiInSKG7RTput37wWdMlywz2GW480krzF
FH/T7OMyQLWt+D0mAmE8I01Qrkz0khJl28vEvVxxtHIc0v90Kv6NmZYIBG1bO+iQ
i4mc7dBJp/ITL0IYUQLiwVHv9+4sPAtZChAhLaQv0UmoZ4tYPvRpcb913yLluLHw
Ut9O7C6/uI31TCu02AwWjiCElnG/kfK9cEgce7qviYnBW5axlPlPFK1cigexKTyt
E35mIxs7mTkkoWdnoF92XcUyteaeAEaFPCkoF0RMxtBiY/pwX2NhIwq3TAg/u7po
gT4fqjRl2OpVYCyQdm+HoNWeSxGT/c9WVGTyaArqw64xW6SGPfYqWvN5/cJpkWyw
KXRsifnukp7E3wAmPjPMmVT1Lq0b4Dg/slcLEcZDgIWffUHa2d6lKfAEZkecYvA0
mS9fEk1Las/9MbKIMEurZRol89cFJOqpBI1pT3fMl8ksq9sLhjvryEPyi4WxFKmz
KF3K+O8o6LSeadnrszgtVkqTIAcASNRJqvWmqNTQAg2j41zSrn7yHBZL7D+FebOK
DCTmvaIdkBQkrHzNU9JjPB0mtTCaqmFmJj4NXiU0HHqRcfvrZ8u5/0siGYmFSBo4
c6p0rbUPHIp+/x8fz1lpm9iuUioh5CNeJJU6Z/0AyqXvTl5f+z/6fEnkh0SADaf9
eiZSPzbgCE0+kvZxjJwm2deaitotC/CUYx2MGq0lK5BqLolGKwutfDoqbUmkMa1r
6gEUUw6ry0Y6v1UzMBEvkSGFvElmb5ki9d0lvIvpFi2FZI47jBuxX4kg1NgFJRhN
YfNzBvnj9RTNFN8xUwQIAq3QabmIvURmgszARifoC4wpTLjmXRcT10/Ifj7Sem1G
lVILe8ICqhtMBOajTG/EEIOPR4gwqMqkMAYw3nxZm7PZMwHAmWldS1Sz+9hLtek0
WEOVfDIEhDNoHm2nXoT/QfsHS11rhnhHvGbq+rudIAkWD/mWt/fWpvTV3ubG5Swe
bKh7/YHuCE62rvzW7+F2OwpJXee4u+zW/oK3o/9cA4G629/gD5meUbeEXKOY0GJB
Uoj1OrmUusxFuKIl61gSPKtKWXj4uhFKigCRjdsLYvMxdwGb1HXSoPOeedH0k+tT
mkZ2sIKSIebH190Uu2ujZ2n5JUn/ArIjehSNE4+DSpkshie/IfRsq1aZRhKY+z/n
Bws9i6NmqcYHJDaIXB6rUk7eqzIkYtCf0Fs6jS0DAdazPJ4TQlbg9ukhuNe8vljz
ogMujgPsk54dZriClDfy7Fni7a7GOvU9cWUxL4ulfdmcVMyzupYrckhwUEQv+Aur
OUL+lwtpDTu6gP42e91uXDEMQ8ulFeBEwWRDtjgD8ZckbNg6tB1d4Fp2FrtXpuWQ
e2tigWu0RXoDaBF2znSi9whzOL0dwN/1GHKZxor7aOwMu1EJLtQKaNUxqplI6kB8
pF4PElBfPb2+dqU229TksmODjHvb1q358CzugkxtJ5lGspIcPooMFUPpTFZn8Nn2
1mXaUf2LkluVnRUnlk2l23yCKPRUaGU74K5PmmV4x1qyDwun4kh1Ib1htlAo4ovO
3Kjh7JtH608PPX2OBCTWHnCx9VUcHq5tSzD/m/FkgIZY+Gpjp3eE3TwI0HkHalOw
bZrZ1AsujSbUyqjp354bEXyetD2l+1LeKVY5VdMCWySEV2jsBXGQwM1RNA1vu5q2
tie2jT4iDH2383/NYgvLvCUo0OPHv1z1FOPRO4bRrKvzZ3IwHV5lAKYq1t/XocXz
UlCua+jjtXoFfPFukCw+4xzmsdbTwh93iPpmD7F5bPHJQPH2gtdShn1hL2bKmR56
wnnOElIfE3nOyEnpIS3WtevCGBHgZ2KtifgA2Mf6w8bZ/+VVRu2+B01jqFa6dhsa
wlOaoLCG0KBE3E8laJzAqmdZ7GH5oy2Mgt25KOFfw6Q8ayuRnGe10gCrK3ueDX1L
UMWwHiK6QUmnIqaCxJ5qlSrNgtbcGG99KFd+tau0159Ol1AIfQ5I3JK3fMgl4OKk
Qs5EjwqovSfoyT8tALv/G0qNHLjI2K7PimOMED8/RVlomlmQQKVGwpcl0dGbNob3
km0CbHsijQZI7qAhPO1A5+WwRi6XT2ODTQL3uwx0k6gYlFHHnyez/DplmjHUzyRy
hUx+MiuU6LNIrFb2p/LwfXLgqNgjfQkjJPXCSl77Gm1vk6BZWbdfQZdt+N8uOv5b
RJsaWfjRqL2qptUrg92FPcQxvGIpPSIGI5OndD4j8owsXxTLEBVuqI0yUotsOwX+
jT3/QI73J2nF7ykNcMe2XS/qSpyYbqx3K4UJvcXhf06NOwObjxMo0bp0j92Qp0mL
9aPyUgB/ayyxVYcG7yk3RtiGwnTOx3yzkPop5c0tfu0zZlyWrgTlwbxIJI6iRdMZ
hx1tZhYpuT5YolI2hGc1dIsqCIWK7hDjL/wUPF0BIdcrCkFwAIoxdnfF7Izzl08s
ai/8PNiN8TPr2KfHO2L7T2GuQO0aTuWJ2bWSnBPis1PgUZgyDR4UgQ/PiHnju3D8
eMHD2lEIlt/3JzflUsATAeCzWPJ3cRH0oPZz7e4I7uFLP1tCBIXcD0nk6g7DP4yP
Tiv0ui2uYXkKcV92aWvjCIrCjXN6t4CAZ/OAPgba3gPJkhfuaPkgjMe5CHQQFugZ
L6/gaqEvdwwhb6SGmwiKYpouQJy5ob1KnBdUm+8Ne3gY04zvX5KwH9bK/uBOV4Q9
vBi/lADWyJPgn4Wg/Qu2eBLJJR8l/KXSTEy80oW4iCJXVADNE89GQSX4m73y/0+6
ZpKF1sLZSKOtvatKPNVe3sr14g0d5bkHs0cPaIH8xZW5IR2lbA5jsIya0X8/OIpG
N6xYn9h5sjOY1dh6u9ykgbhvIUmHYQuSJ9bidEVWqxv7L08jCecSAf/5TEJYgcPs
Qo4qGW/maWYiMyYTrsi22BI5vCHS3BuwKQqrz1pmHAZxAAeXXHZhvzEGdS0Xl4AM
Mvnk1t13D7KBmbjaOepHF4wftxEYuKJHxTRnrSZ09IzbX2EPfwXWqp4Ptx2tbZYI
mp7HF79bqSAtNrpXQs4WUC74F1RB/seTD0U47lUKcDgbQSGmDllLcAUuvtuS8nT+
ZTaf8kURtZkzKZM9IdC8/qZdjZB4x6PjVY4wsbt/cz3MPMEOnlA5W8yvdZuf4M31
Fzbsk6XYKHXftoIJ02IMwh650T/dyLiA51XTy/0Rg+s+gmtZuneiuDQ/5oHGiCvg
+iPuW+CGcaw5K3TNO6EhTlI608EyN78VibUJBJ7ctoNz1fCQrijNT/tlzeiLTOGW
TNNggUB7Z7BTPlq63kEUuo/H8xJ/xy4InuVefN3E3V5g64aEj7IwAfi+EcNnByN+
U3enqlgLJyquVyqzf5g3MJ2z+uRvMB0oqD9uyT1sJGwPNDcMg5hBg3hvrivBcTfS
lKxm84FDbw0yBNSkCRT/S8ltzaYUvqolie2FfVTJJroFZIZKbmwFDBMMMjgGDSAR
eqGR6c5kmKeEslFg/knsNQ8VRG1K7bsHko82mx4jakirNbG3jWdyBl8NMcXLYqr7
KGPA5caac4Gm+jXKmpCXrUVYM8ZoGdvVgNDY5gHBhG9cDbr2NFsyxD4bhAKnizAK
9PwZUcZxFncJlv039c7PvqC1MQNyzD23fU9Ra2og8s8/JRifKEDy6bCnTPYIdnlY
O8OWqbA2ZyZUiO7/Y05J/8AJx31pImvqIjoH76KWgz5PdWvvyzXTkwTM+x7VPX8R
Xb4VQO9jVjwR2WLyIOc+i8q8TAoMV7J+kek3LgPevSsMsy5L9mPkNnAhAa4tN0EC
nWt5OXbMOxAyCc9N+F1kdmNOY2KE1ozqaB5j8ftYfIwKxsJ9XRhY0aJNVmbunN2Z
f1zma/lM0eF0SvvbPpkF5qQs8E0ntkSywl6K295/cQP5m4dZTUtuPm0fwE2fkxof
tVXxpmmr0kXIGAElkk0Q/84sU4ExAoEJNwI31QBSV3UWZNlOYN9iWfixxGQJvQha
TOSGXU4taDJqkXY7Iqz83UPQN8XPyn5S0xB7IFZzBaetnw0YnfnGx1ElFEM4Itp9
m8M7yqZh1FkKe8wHsx2Db/HeQq2/lxcNFQGgT+G5Gh+gAdJRrepuiMX20IUvN6LL
ZXPkj5LNzbC2b7yZIYLPd+65adnO1rit6IF09LUWjTZ4kNFsqgkISrNw5/+oWg9D
9GkpNbzwORht7vHiGjTt4MRWnOqnpouN3t9/CRlEaxep/EzNRFYWvRhKMwu5GH7p
L2nejZc45kv1D1WLjcBkeNlSo3WzfCZqJLB4PnqvR5feTmcbnOThqwKMsLuWb+oi
ZyLfDX8pbtjHsQZMPJxY3YMRDOnntJUWRxpGKDsOsGGg7ajWMmYqLMipQzfpKP1b
GuXAKz4icGHd+LtuvuNOZX4KGgpLmw7at+I4CdL58wyollNcA+iAR77BWL+rSsfz
+ENBOsas7POa4R5RNY1qWYwx57nMpMmnAMJcAUDxVORJZ7HMWHZWW9wfVZD8jIua
pAwM8luEnPG5rrtFUIgmacD+Hy7QueK0lyUEXWK6SXB1E6FEubTCbDSHOPaH3XaL
knYb5B+jhqgthbe1sM9+3AbWflzMPLbVNOJx8FizXuDDuyhejzuo+wOBQt0yz9tO
lDQrXUAJhy+LXG4DuKK/E5Dl+NXqh01wWFPFa+eFAOo8HUhGpuD5Ma+8YtGwFdie
8DH6dtk0f2O3c3OEar+fDWbTc0iFzoSqZ+yLHxPAiWihHBLw4/3BqwQC3fknOfpG
z0jz1YX6AX2ooqJwfkvvE11rzS8nQN1CFxtqkfZalDu65s/Y8E1VgEJ8tHLmwbBA
yJo7NpS6L8HG+3C1Mg6LKaZ9L2Pmmvf+GbCN3tXT4Tl1b+e1kdbGkFbKVW1FI1ZY
/tmQBdyAPyS2c+/ufN/DmLShoEKNF6T6K5avLjrM9p+ZOeB6R+GKClaxN+DflsFX
VgQr0XlcbUkimHP7JgBpOqFHVN1bbY64LmTfdjdtR+O051gRRGEyHbrqvZAJF3Hp
Fo8cb0plS2k1MCt9tG0Uc1Zht5BPm31WXJ69H1l3ogomdxsgKVyMhCRufjbEMFHu
bQr8u2YAUUtCIuqeD0gyM689cQ511M0AY3munfiWYDRmD0g504FZEkMLpCTQ/PxP
v/tDOYztjHYUJxpHT61VAGyOXMpWC22zhx2d0jlYJKB1oE5Npp/41lRLxEJKo0Wt
xa5fK4UrcIYjISFuJKCQSOvVlciLb6ArIo3ibmRUJtye25J8hoyQnduDa8XF4yrV
btCxdmiVteK+0pAJP4tJoiFRd+XTuWPmWtqSYq/4qoK+aGXRp3eN9bDURL+6GXel
gY8tmoxCNFLDNlW9EMHChk3VE9kAbgyY9QVhuiqvk97qD9puOoQ/lf9NcsPN8/4t
dCfYlJlH6veI0x1yCwKEYfhKGra9HIsf8P06O9ppf80P3pCQLsVKDijHGE1Vf4I6
oYg64i/+Fb/ltLkVBWqw5INQTq4eQIJk9XZBwtZr2R7u3C0bqW0bN1mbsaR8cb4a
/EpoekuWGPaiELawBz+GPdn6DYd8Ika9QGVFIrRr/dUSWuLJuyS/UfsUSKJ+ghYH
ehH8xDbzNWL65BhPX8x1LqKPS5Jh4lyAGK1PM76OAXp1hJ7+jvbPCZgxysxXiPdS
4LDtI6SEKXAQaADEUWmjEoWVEVcpj/OqbXzGDmwXzsBtcjroAs7OI7A5UeDSRrdw
FZmUJ4HU1D/1jnikY7NWmI5nkdWdgKdlFtvsivhKmyblwJjD+3MmXB67HWh34rYk
2ZEBYxrhcxtQXshIHIXh9z/9Si/UqJBzzZHm8lWy8XHDNB1VlpGmSqxpUWAGSaTG
FK/+rbEnxChmBOGYlHP511nA2LttjQWi+KZpONpIQPs2veDAgfnJzgeQvBzTyj+r
Bupi6dUZPQ3kXIZ0eYIxSgl94iviZ97+kFS3GBC+qjJaz5kNlTrUInOtieShZdBk
PW/MECrwZOtJ0UIbVLhRP8vlKHIhUZ5pk5rsiYmn+oFy5jcAZqRznoFLGTRL1STM
pTUwYMqdvqjRB6yQm2tWm5RgjZA8+Gjs1aXdDFGNKCGXa8HoDmeyiV+pDeGLvmFH
ee+bpioQmGbO9kOyQJcol7nAQQxPbGWGtAiBDcEBnXBXLnIZKGWprgtqeJ/4qqMA
uV9ooHtSFgN2Y+fy7ZalcvunCfhkOMsQqhd76RjiAC3HZCXhfY6NEYeOpHlPO56f
6ZEG9UTwzNWdCcKXd7V4iVhumE2s8bdcJvLJBGlQPymtA8i18DD/u+nxyqqfbuvZ
YcbsJTM3wabtQEJa9QyDydNe3vOFlL5BnQJ5G+iUtb5xY+ezirxAFn7AOmTRXUHS
wnzgFIfJgK2NXASiILX27WmukiG4jlV6ro6AmoMh+horJADa3Dg/w10VHhEEBmOK
8L1+mUKYq8vbUgfPEOY2C1f5MrHfBK3LYxq7ILAvAcITygKzj5oCxEtPQjBkENrn
CN8g05Uq7Po9a8uA2gO8NHRAraM/Dcja9l24ovy1ffBGqyP9pMXEzQphjJbBY5WZ
Or3R+JWHtcsuQjXkA1sodoofw70SCp5yzMn4menN6HPjeNDNj7bMsFXthkeVS9Uv
Ip/W7X8JefclZbEGAdDE66uWfW7uK3ge5EizPhZ2EHyES4INChG4N/ymLlX1RKEv
i1i9ogFlkRO6RdX7IJtAybJwV9BkU3Bxzw+c/xOKDW5aPZNo7tlwKNQ7GSC/8TXg
3EJEvstyJUrJLxuSvc4+XCJ4+OY+A8F79o0CuD0LXxdE9/PMk17tVGn19U2U5KbW
CR6SL3U8LahjYEvJHbk/L3QzG6jiTWzrYOrC0JOjGqq7lamEPMr2AhtfGP3dIwSm
2NNQ2Zlo2HZOYkESvYcRTtWWbyPKqnpI6TPkxWN9sQGrNEcc97hd7iHQyTtbcPlE
GCqUisCWAyGOfnCcmRn//gPkMI13W6UO5PcPPLaSgH0G2j9n1isQhQXCyFf+COjX
NfXB/0sEFMdXT7Y5EWPPfBWK8BHipBjOw86P6+JkSL9cR0GJFm2FMOQi8z7I21d+
wwnLzubCXsEd4TYN9RG18GIrPu31NTMLwEoVJE9/TOUZ7vnbo4iykm1xiYgDQO1y
x799m/csYuYSEwZpmnuz7KJbBIWsYrsnyeJBJHn6+BNFykeRoM/kQBxVdtM1/kaB
Oc1+xeWQNk+CbylsXWEfbJctCUzQpOc/ZdFJ2/k6WcxdJSDPWU335OUdx5e6N6nH
F8uvj9P4gg5VXGcNtDKscPxuNLeF4PtJrxu2tGaFjAxryjyOHsmIVuZROx7SgQtK
MVOVAjJRJKvFIIbB9GllnU577HymTjirhlstOSbYIHdhHPZe/suglMTphkJ0rQTH
tBUMmDJiYSfI02bCobCNJCI5KEQ6Aau+/2fR7EM2CKroC0h5oxevYhXhYj+TUm6c
V+GCOfESIeGU2FSDbhH36RzicCS47RfnTCWRtmcEE7EJ6Hgj0peTv5lt96Uz0Bn+
xl4MNB20XOtJWQIGcpfuujcrSDR4wF5bDSBUYxiqkMJgoxmBwkIA6E4lW2KWFtps
Q/Wi5+LahfcySor8vrwcis0Egq8jWBXanXdLGmX6JJMXUflKtZLgoAFnip2SrenA
ZnlNXCB6f7mqpjj2MtaWSor8tsZDk5YUtG7r5h2WDuqVSZXPGaY0sLRh7MWQdiGA
JtGLfGVyWDANw4H3pA1Ylf6XK4nkpEGIsPheogtghiyrxApzggYDVWPwc7YeEghX
Y1n4sGal3b3bYxD6A3b06oevrBmwHrUzAx6+EcqdTofR6BP9yia4am9wIrpyv3Zg
6p0r4AqUEJPDonOr5UZ7LHAvf2O8PBl323F6FSnvkI9d+i6bf2Z0IZkDEtnpLyJq
5HzFQWwvj7UZT/RM0dHe/rqMW0+fOvfBSpgZ4b/2g7wYgSwe93JZjPJyULOJ+jfn
nJ5Oxv9Q3XSgTKLatMjV+DEpaQ42DmKA7WR8qYda+rf4W+8n8eRjXRIQRAccYCOl
PukYZ7+FMvSklQIP8dbXnmOIOrdBtgjtQ4sOH2YbvvFqfnas2q3/8O7PTE2yM1Jb
XMn5nnVYbo7i33TY9uCRG6Y4REwY90rZQZuA1KzKPP1UICq78q1aq+XS02vqCX3a
AxdB4XVnELMn9cmsn0KIXCbJ0O7GQ4s22Uqxmy8Tng/7OO4q/mNl4ZM/aoa3Mrk+
UbVINopXA9gQzQkUdQB3zqDBpn3b04/NCh7ytwE1qJvFYnJ57NClo7TXN9Ax2OYX
tDZ4/8jfnwXQrrfrLRb6GPKr7Q7/xt9paZj2HkHIPcGJ0nUx+Fd5WEcubTid29tN
f+ant/rVFpK1jw815mFogVgbemRF4pXHbWEotee1oVdc+b1HGakYfdRP/Iik68wp
kakMEmDYPxZh0/5F6RhYBcJEQYxhSOFDhaPsaCjx6UKg4xY/7V6nfL6F89LeD182
FUWBlsJ8+EHUl04hJJLXY8I64aFN1p9I6AgQbEH5A+OYvdODYNneLhBR/YiZQ8LF
wDieyI5nhK2wg8BizM/cNYlsjlCKp7ywb7dTkxdHzE83A6xEFJsNmuJ7JMdCnals
ThFXVmaZf41hL87kNYOc5EmiQ/s49myh8ie4wfbZin+/UCHOWadEMWnlBgoVACo6
Yf7actUx+yWyfAs8GYF6qDsbyn2VSbn2afuEjB9R9iuwQL/Slmc+OfWNl08iWRE6
gun7UB6KJiL0E5GtbJDLF8L0U3mqkjt/oRwN5VRdpDRkpAiCnsC64x7TuagW8R+Y
yTkv2/9PXPD0rzDYW4rDbiPMNX7rMlzwGFYudg32K1v4ub2SvIkBCNHYrNS4SnDF
eTnZ9oM6mEhkFlu/jB/EBO0SHTSav1iOyTUVr90gq1L26xH7WEb/Hebae4fHLIR/
F4imZa00Hz2O17GMgpaohbY7/XHD2eyRaSwpAMznVvdcUOp7tC8WBnWjXDX6lpSB
LqoZmkoESLIrnNlGURJDczZS5NmHUqBcXxxTI8HD/0RG2i+egvOADosP8i+4Plxz
HwajoRfZjp2Uw2QG8ab7aYPBKIMYP4DUggPKZyxmBcCKypE4C0Z2NNeuAxqsaLbd
YS8O9S1ZA9ycaH+TcezZKH2XuzEiylNAlVl37l1R1WxV4B3mOUQfa+LgEOgtcbvQ
KczjoHuVL/MArbOAaQQKeybt4Bb95SdbaC24JvszTk8WvXalu1c2I1h05D10Qj2r
/7jYIKcXKvvtsAnJoc0pJRrYAOKDL9t1N69Qtb87Is31rCUHrFROvYT2kP7LtrK+
39o79NtTFjiTwsven0g950GVs+Ie8WF5Zz/KJ608sdXToUkMcPC2ss/prSjgd54q
YpKvzQ7paCxVvl32chcD0QOWgMCB4xMWdxM5Pcqehu8rqCbTr7NJdaBhEgE8fyR7
vQ61oijr4lE9otFyNB+BHx8YGX1ljGlgjnTfkg58an+AiLkM4ad5cOqHf9nPWT69
yJzBO7tNuHAnWb/KdHLARMqSiCKaQU5/oDsWnpO4xOv/hiLuFLV0QC+JXKSHyxzG
YcjxpelPI/z2xsZqNtHShaO6KmcsAldMxcVYXxrJJ5KlXmVt64xPVt98PCy5V0x2
rnMzfNx5T3fPYqlSTuCFk2oQtZx3q14tt4ltixo3lC2Ko4MKInVuhO5oLZWiSGrb
H7DI377fjDoCtVWn1QzHlSyGfi66EQjOQHBZPk0miVGoX1xpyMDLqJD6tkQjpwJe
ATlXA06AhY5TY7gQzOauRwBjt6jJJud3PseZDeeBxzCf1fTc6rP4QBoPRwA/5fKX
R5+Ug1VqMCS+W/2oK86jr++i+WHuriby6JQ+VH6oo2lnklsEw+Z5ZpyNYIg6d6Md
gN/u3Lqcm9zLYCIIq11isauuWB9HyMyzS1XqKT3bm31AS7B6x7FIyvVpFDZCHoiX
n/cO927WXcejcjWvXiSHQmYHadLp50ZXyORD6Ol44WWpZRFqJzJiG8QHlxR1nIji
9ly/pMjD3vv43H2ksiDiMCZLNdYIJRaVbNGXcqhGZ5SfwE8Y4IGk1GAUNToFWcvI
PauAsLqMerfjiaqjr3qvzEfbDiy6yQ/uAZEstSz9UuVUq4+NOKK6xros7AXtXk/3
SKEt2QMBpzPKR07jYzKQ3WfESL2TmWa1PiM4ApxM0HaYfom23YswVeB58bJOkWi0
UatBy4rrYPyFj/80/6GOeeqMKWc35GrzN8i9E1de2rk3zbBzr+hfRWP/rW5Vlqxv
+kaXNW9Gyxjg4QRa5QOQuncuwollM0bxkYHmGD2oG0zZ1YDgiy/PKeY43hEeIn0j
kyfhUunmpYHG5N21Z1xpCjNNDqrixjJXBBitj8zHrDWki5+PsE0QYJhCB8DDY+/f
5l+PFIU8GZvnnVSixriYKndGLdVnv/XZB0VDhrQpSDhtf9IHU2F1kpOPf3yAu1Vj
jC9YUrG38Is/LAHnGARfXFL3mC3MzeSGZ3/cD61WKYt9glufP9HmcI5B0S3ukQj6
i9rE9gXOpe0aqpyi1H6Szq3jk8M4xEe0QwQ2//8oKTGtTdozZtfiCpmyzJ3A4hGA
QvLiIazNwGKZ+MPmt+F0yJYUM1IJcOG5wSvoYX09bITPBmMsWd68WtpLVtxnUyl0
jWbk5wfDYi1sA06mO0UsX91PLcwM+95VPdIcZVzByPa3XbZB7wJt+yuGMvxynRXB
8GbTpru3dUFDCzUDAzIKTRV3HPOLtblAGGIb+6j+PXZjTnGcsqUgEosmHaDU4k9I
Ta70BrnIN1vn5ox7cseiurTHXW7Zrhb3wDwGldT803G/JhmVV6F/Cjyr22u0b2+T
NaUHCTpuL+YGDBivffmzJ21lGykb/FXIFoa2eFbXRb829QvA3reQ6LFyjHHlgFUs
hwXfCLIKQBQnDj2Bgzqp4XZGER0/oooytPkv0Rwa5Dl7viG1L5EEbRHy9HlqaCP+
E18hKxtwpgspIO9IZgBxNhFWvfhFViaalvJpSCvIWdXj2HWzSp2PDiFIa9mEfzqa
QLV6oYiPcmJswMtv8OsggW8Wmj/32MYrFM5MA0PC8L9aZSPSiad38+ilEoj8AAiz
kuew2iYccqUM1v3R4qDCmge+yL3yueV/hHFPFarzo1k8Zv4cxyJry3CTO7Sa5ohn
Y9fdEs7u/WUN2IdDkpTc9iGCcR804p4cLW7XVJLUxFE8zLim4RuTRlXNWcG8T/hz
Ie6oPgECn7MQgmvd/x/rLvV6chpravvDY46hq+3IzU6s/nDemJn2CMuinEbqHGSy
XvUegf1ktb3kapyLm8szFRFcq+TY/42bjP86w9AzhCfLyJ/uL8eLeaNyphB/jnia
gEi3lDOTvizdvV6xHvx3t5rES25KaVgExn+9YRWEC6u0731noI1A2T25/jJT8mWj
UmBFrQiPGCon8DQ4Fq4kJuu/cUw9XfZz4PNIcj47jyG+HNgH0RyON2rxbXEH+p+K
awhMwA7XuNNzlBD7hcmgPzNgaYVnA6m06e9PlCkz2hX6HdfRQ4ZcGZacqAUcxmmF
+R/BCH/7o5QCkM0aWl/lTxGelCFCOGlziHuIpdwhFD/p1koQYqZWrY/dnkxU5NBt
VoxdWmsn/F86pezzt7KyakckEOv5lZVux98sTQ/77uvWUuJTkSrsaBvh3bODqZrt
GTDAkNpgepSRMbF95ERHsdl0A5/unhixRHaogAZKNBnghuzSRpMPFqE8l0SocSOO
CS/Zw1aU0NKoozT4Di8KQVFrvkoFgJkMd/gHjWPbyxA65WyEUH+PNZR6ssO68+Cp
5NZwnYA2Qa0mynwxPSppKyy4KRNn5rLy0wvVPrDv61Rv14KkHO1ViLBL0G+Z/qrG
rwF7VIwdEWvRgoYHCN+uatmdtGmPm+Zf+sLEgmuYyYaxQ/M/BjEpm1BTk4n41PcY
7KRPGN5Zyk24WG75QTiBKjlVYin8BEB/mM7lfiqpt2CXU7l0d7eto/9V51tOsVOn
8W1rRTr0FuxEYQCbi/VxGn3iv5e0/6peX7dR8y7dNEFeRNsbf9GDZKo3YAiCCtSs
1z3pNl8GcthK8oLmCnavi5AteyFSgISi1R2j8UFVo/PNVIMQN2oGGIur3kCOztdU
2M6Ulnc1zKUckHIHCRD8qijAAxq0mUhcMi78uflALho5j2hj9ic6Ewbfzd+ZDduq
RLpEns3IwLkbolo6pVmWY0gWNGt/aync0VSmNlnR6RCKpIU7iEtG+uIWBAIALyY9
CA08PQs/RqGQqRozg+LDnHIIw+2OOjY8MTxl+meV4z/C825k5Kx0aQ9wv9F+7mcw
ppss1yNk2IzfhoF5igjEgA7GVTURV6ZuNYPEaVWMdYAofEvsSbOSip39KhMow9q0
8rplrP3z58lWt1J6VfjbBwkxfLM7UVJ7DlOI5eTNdJpbgIlHQFhO21tipMW6LDMC
DV6u0TkPt35wUDqsCmaAgBP8410agmj9MuSFOHtoYJfiaVHP3rjLjcdROHtCs7te
98byoQ2E5xSDHfd302HU5GhAlt+Z7FlfiY7tI1y7LzPx28uEU4c1/jd+VQIjXlxD
DlJoXzk0CSvzvBlqZhtEJmMESxcvYy7w302REolMA0B0kmy3fyAywgZI+8ozSmcG
BdoCMYjxqWriW1UHGsLAVpvsnunbeSFLVq1EKyENFHtcgShZkj/fYho/PxQmIF2t
f1SKQlWffWdRlVSw5x862LMGGY9UPqVti50A6ms6mJk49o+KZWTbZ3+dQSMtnnAR
9PW9QY3dSz9Ri7yuFA+jMx8GMrm8Doyv1BXpB2vcnfgps3aeApbmVqYpMmhAevhu
EA/Tx5mqggNwmkvzn8T0CwBtj/E/efaZDpOo/dV2WxxRGPJ54YHQ++vE52CrumEK
sBPLLauoHQXYMU/2rUvqcOlVxsO21Blvmuh+cZSTHOJbQvcwLqj7RB3lOpACDMZM
AtvxSR/5/UaeQTatb9lpod391JquS4H+mmFSZ6A63gKotn6fRRRdgOao+viOlYFH
E0YAak2kSdfbkm1+ddswf8wkRD8QAhgU90+98racft5SoAcypLU+qbuozjdWbloJ
Vao+LvVRkV3QV0qrELJhG2UBjR5hazeoGi98M25QmUy6qBYl0xl7u5MT8N40ToeI
KYgEN324TZV/BNZRcU1HNhcqnQDOGW73+BclZakZZ1+PE5yjuRfw0ehZTU+xWf7g
Bg9sUtQh5l+G8e0Rkjt92vRxrnRjBmyev9oJIGPi68v4xAQrLgiOBYOaT3dNM1aS
QxUzIO0rHn5hhQZ/BoINQerSI4aomXR3mdgfNGUwBZpCr0thL55c2anPc7RSwE4/
j9wb/3YI5WL+m9mFh1HBYr0gFnhRoks7cYiuT2l8674TMDl/rHFu3vg4/wvapIsQ
IZiAqgUM0ckyl9LuX2T+NNNerlocSqFjW3hVKhVse4fDifRSPi68A/ZeTehcDTBZ
0WJB5w1AzGUMiJb+/mI6Hd+CWlSsV6HUVZT2svJMID13Tqz/pxyrdLCSTXg00YRt
HLATbgkdWOaMD74zi862cn5R3+Iu+g1So6HFX2iQEUpOzmaTZKkS6fiOO6PTeDlR
vODfaFwYPMp5i8/GM1efKzUitAlvcB9nLxxDk8J7LBQ+wzztuYHwpkeNnUgYxlsd
JIsUs/SOBFXsRv5DdbF7ZWoq8XD+FatybIMhvbwP8SpyXhdEZ87ELE7uqg6+dgxu
PjD87XlG3+Sz+/uAdOuED74BQEj5SBZL95QTSxvCFcldnlY+K+xNKgZdXpjsC9rk
qXhVgwG5rTQm34bBQuyWqLy70HnsYY9A6S3vHCvYF5X6XU/FIsy7Rxr2LIoJElmu
Lp89m6IR4U2WSWoKvEDwa8oX870J1BmQbtZ7GmyY2gfiOIcRtODheM6Gy6kqiHh2
Ud23qdaCvjdYEVy0HgpZFAuQlG8dEMKb/xlGKKqZMw479jEX3tknRty4clCBKC2h
cOKeSeZSj4xvhez+VWsweUc+k//BlJ4kGH5flG4e5yVt7OiLeW/NFMUt2iuGjHzD
RDid/JrTbPsTyXObWmyi2tIJiR9HFU1jyhQaK5pBLKKwoVXGv0U0cWCQ+STIiqi7
A8I4iETJ63lzMwtTkncDf06U9eRBimdBnRFuaVrNNk+BTHCORlUZfh+6TqXVo01n
CCLcBXNBnSK5y+5vjY8tOQrB7rHu8QEFrcxDx5hJr+7fiqh8ZSA7H/iYIvEDhe7O
ZrZs9K5y14EViW/xNtVnajjJ8gkPgXHSdvhsOkk4l/fV+gJtoF7h1hIn3IX3xtNL
gobRzkUoIOw2Vyvlgbn6n/oKrP5eSbfaw23LRbo2RawLTGCWKcEXIbeSKjMbG+7p
ZdfmMGK18Rm77TegPrg5DSMIY9c1SP/Fq3yQkIYFF3Atgrt2JdIoDggu4CQiIY2S
qV0oc4ksdG82c6nw76hRagU+GFFcbCoB2LpW3/xqggVojvoBRvi9qlS5mBlDb6Xm
2HQTZm2w8NoRh2kdkaJaFP2txtrpUsWrNwYuu8MK9lC0DA1lHdy+Jw4ikB53JcLl
vxkxAloVVOo+l7QeMESh2uhAjd3W9aChIckj+iuzD/B/eVshB2wkxj91uMDay0jF
n4xqMX8thY+UbXM+Q5/Lucc4yu9WT46X1hdvg7I9i3Tghyzdxw8GsJiZdnMUMl0o
tGvP0XVa3FAJllsnLnppcXAcXTHpEaf+hNdQYhvZSVM89UaRe0QUFHkZ67Uwb5sI
tu5bTlEe44yyjR2E3xpTcYwt+yUTwZMIQEdliXMV7yPNnvwLKWIY4v3KfEsmBzYD
nFOT6MPthP7TjgV1vIW1Pi/AlpQJJhUaJyNbLL6zMoQWk/5PJUusgBFCUHRa2VjS
xWvS8p84IjZOQEbTneXYfJeU8XTCxfEeLedjIS2vEUEmP7Mn48db4DEDSkFEd7iy
d0Ny8G4NDItD8WKx7U6UNI3Pp2TqTY9bma4uDpSD+BdhiFkRPwzL/Xe1AfrjjDd5
QSPPoqqIiSY8Cj13BItAZ0LJOs4dX/P/2JDx0zSE0QVFHNKB0Ub55i9NCu6+YQtz
LJBo+Ra3WhcREeamsYPnY4S5/65K4u1MU4QhrZwpM7j1lsQ/i3JVg1KFt1BCiZeV
IVOtUsf72YWDkXkA/Php3hnPGPKdWL05SatczK7lUO3TSWCOzMlewuU+OH+5HYDi
m+KnfSoLCGvqEIhIGhZ/efNStJsFsoP6HUoPYTfDtoQJwA9bI4usP6VB0rd6OzG2
o9ac+s8wZt0pfsWUaSZpBbXK2Qkm+4UErDstmlVTSNkwuDEeJfouvGemaZZJ4+mo
opUnDrqFa2fIM0igUemOpAYdPT66JZR8zPMx0kDd2EhIFoKGfe6k0/f6kWtPtdWv
j6xbsiZ65JgUNbfL2j3iPAhr4Xe1IaS5Pwl/IQZgTjia5x/LXatrbkpxYCrV34CC
fsjMTd6kEv2/ZnlL8e5Y8QkDA7w3BjHz49z8A7mRjGTRNImmRiO6nctmy7JX4+cJ
hJGic/d8TUcq3oL8RylwX7Ex3/WeA4lHsQi49YpGD3NQVCUfB21IH2s6DxE2utGL
iBwgM3NHd6EQBGxcSVFSb+R102sbTTIvmF+L7od5sQKiJugF6YdiypUMV/HQkeUA
SmGH7cedNTKY4RDJZm+xoADvjr02wv5TwE5Q6k6YcQ9TLw5gVGXIYSQuER5T1QI1
InbuNi1FUS/xwNzC18UlX/WWJKVCXfKyC+ytE0CsMVOzFeel/ZoIL89sZdxWomKA
ZAUQrBc+60fqn7L6o70duKUkAhwTX+Q6TllNwp5qCI0c7Khp/WsIlGC/pQM9E9o8
0irfG85Qm4l40oJw61HLppvPtRCHC2PnytgWj9XeaUd90VGjxJFiG3560+eyi+rG
6Zx56u8/E0/XNiayjk1oh6oIFoDcLKqSxk7U0It4J3HmInWkj4S9D18yE5IbcDEC
BYJak8eX5GhvTibtda0xuBT07Rs+BsncPqkFuf8JhN+tZRuA5bx1VMG6SN/WZnEV
y9J8ARoVKKStEnabyISORITKPn2CdnNISUlnDOHzcaoym6kHwt/FDP5bhCEh5+Ui
7h5C5hmx22Zr+oOIcv32d7FsvBVzvv/SgehRYOTpLXOV10r2hdj/3odIHtz4YDVu
vEL+sL5EnxXSYVpmaBKdgX2EFI5D2jUzX+C9A2n6c0QO7bzzAMW9AJsOa8Sbf0J/
R7luf+nKkN/zoiNIoWSA1jdPzkfGVJaTe+Pmsy8EQvmB3J2wwriQ7dlPC6rwtj3O
vXgqaAk/VmW59DXe5SBQ0WIUniC7Z2SeVlQYLusjCQRt0FRgn4CDw5iRNAaNcgqv
EEPaOIKX+oDQbMTb9ZT5bYClmMzjMuuPXYYLIJOlG4wkhCm+Dy3Rmp8CcYQ517XQ
FAETQYcY9VIxhMJDdOyNRNHGZuyFDxDqGP/VcrCSzgGWjiuB03OM8CgQbLCP/hRa
poXJW1mxGb8TA2rftF5BGkwaIqUwGWW+k0TBrNxBojgHT683xDQz7iLaud9o9Ea6
b5aDOgobfzwZlTCA0O6I6Apht/+Eo603dwIKvX98RKTs6NUJ0+A2Glf2XK4Yz0wf
zM+wb1jTWxcGO8YIMgH9zBe7PAzf4cGRzqZLyQfeDbXkdP+u5nUlvSfc2KfovAUg
eRBAwFCy+QXz9EMmooUoixWnG5WFzTu4fRQZAhZdJZTN/JmGfI2z0sHbZEc9IkyB
aBDfDFEZ3+hyeXuSIvnf/IqoFKkBzZxWd7m/rkVfo4LKcXy785tD3fVWhKIXPnR6
vfE8TOd5z44xBbs8w4btBx1sDN5dJ+BMk64/1bqimLZj2kCQEynqRBSAE2lxSMok
rbfmZdb1pjLY/Lsw2KtutB3Uc/NqV60445YByLLZPXDH/+eDq90Kx0JgBHyGiivu
WMnw2isMKwFka5gYggCZSHiIJNNk3NKa3TgHM5sev9PqDxa70gz4TgGRPVsOeueW
yH5wmPlzZfCK83O19O2LrfERpLOY554SRt4SctBvvB0RlfTRLP5XG1mhrLjcbQdh
vxWtwDtMwJUIPknT4mCOViWX/xUThquJ+bM2RftX5k9bkwv1H9MjRwDhS2ixe35M
2F0FKlk6ID8pt6LslsDxW2H7cB5/AqFQ0QLGRXOQFC0IJxNCrCZfuloI1t7TaZwg
pUTTvbcFvEDL0uomMIKGhf8jUbOJdntL/imAoblICpvMgpaBSsRpMO2o5vEMGBBS
NdMdbo+59DugCK4JXDm8t0d3Ril89/MDjuImFsx0qaEfnYmPCekL5B2yKBd0596Y
pnU5rkv+xK/sqRIShYjrBLl+zTM3E+1V9xD3SeuFfj1//DoosAUe2GoKtYA+xGmK
AVjPkBtV/90h4pJfN5lDFdjEsqqFNPZHfpp7J+NwmghQkBHWfLTHQqpylZpbPijM
fxjnZ8iWnnrs82IhZV4hrSmmI5PvzrXeG0aez8MX6ofxEoyvHfgYbztUoPHGzXz+
rF+T70PwhdMFuwF3UiwvNvd2i6onaqiyY/xLvPHBGZ7xDOjZGknXg3R4OmHHzve0
Gj37g/LvrPpYdyojwJWLG6rmKYZ4Z4FV5ch+ZkFcf3i5C9tZuOwEjALEJv4PXXj+
8zhxpE6RRmHku/K9NMCOXg4j7AoLDW+xTEetJdDb1cg3ZJKR6iAZ1RYHNmhblgF5
vqtas1k096Im4e2Zzro+AZt3236p3G5UUPrvVgoWtsUY/SDSPOYNrczvTexuBih/
r7lQuFMU1ZZT5AP/eVlbywWN84kBZOv/29YJs1igmgsKVQqaUozn2602DrzUYLky
nCQjOq/6sJuz9hE+0c6DtDemdHLHE5LPRPr79qCIMvvdAC4e18ymuo7LGzxyOUph
Q9iMNjgsz1YdStZCd8jOPI5uiLWKgVqPEcvdeUiW3G97vS+arbuGJPDMLFgdpjnP
Z/KQiktl3M2J1rVN6z98AqLFVZrjgliwdNNmm2CDCFqdjrM2nRIkDKao9MIQ07fr
FLb/+hsVAn4tRMvE+OZM8bz4HqFNXlA6+TGUJJ3TYMXp/dAYKDluCK/FUK0eW5GR
YIFCc7qk7uoKwoTOIJEb7oAG2uSh01esipc8ABbUCyWlia/XaTf1eWpp+LAVPtPU
EZ2YdTXAxhI8qAU4mdtPS6Vas296+ScpqoznJCBnZPVmvHoijVi7OHizrIUQ/Uwi
FWyhSrype2nfNs8dkd0e5yV3oiYCfY1Q10pUchWYV6K4aZspoD7fI9eVGwTxOKvt
9kKKRmsNlmQoSwoGqX/hYrEeOdXjCf/PFU8wgN26qCPbbpUcilHYy8VXlwBKrfo1
yrXWY6DAMQorzyyB5tVBmJ3o+0TpRp6gMp0kid8LN4bmvm6QtUzEe9sDJpyKawd1
Rcvl0lJyhCd4lLIzMpwHR9a1hP6ccmj1eQR+CtjTKxAv1APuE5/txgnD1+QuCfP5
x/i+uW3Reu7GLYQgye1IJVnsZnx3V/bfYYD1RYbD7+Ky/VEkS9Yu85GKIwhc56b+
EfvyopHwj0q4lOGQhl6opiEqOvspie6QEH3Zhnh/cAJhwdqZHH7rScxfU8BRttug
nCU6ioRe+P3DjD+ied76PqFKHLSMne0xQ2sQg267h9hc5SLHR1VgS/0QVIu28HHr
ds2Bq8aguoM9IlVdRWPzMXHQsXgtg37Lir2mNuZ5ejHpHHX1J3E0vHZqPyYk55qZ
gHFYpZRBlW/fMRzOBteb9ph/0T8NUrv8VmAhbzULtkN9fbSwxTkMd7xChp5suz/L
wkslNj3npiGg4v5T7atCCEdMXHqwpNiQgcHyG9uqKhsjYRwgsaOK3S7eI5KSbbJI
krCmKLtAuDo2pXA2vvfGsHjhIEjqwi5DDLrsLsiSzz9WKno2+pylSpdt/rCsSIxD
8l3IBa9JDEpfr1yFmbvgF/w5FRGz2dIzotEfp3Ymm+zCmyUI/H4Gt8cQAYj4+NRC
poW7paofXj8b1tHpCHMjkbnd20PHFgMYm63pZhc/dMGiRAeOY8SLSMUph4TF2JJo
FT55DMv9h+i9EjA8bmMQAgmhO2PPt//ZnMCQC9lrJIWS+kV343yLX86zE5up93ZC
d6+ZRWbxXZqw0KoVN1XVy23HftnBvPjjGaRociyrCPd/a34BgsrC0RhpSJi/eEHO
Ju/sPsvlra43x2H97UD/0IzJibczKAo6qITgSGHeb6oFu61xuVixFEzWZMMP4NTA
yb9CvTAuy68SxHHMsofchn5FMQnWRx4wLGF/cpIGp9OptfSyCDgpO5Ucr3APShUr
oT2rEtRxgEqN28J43R3BcG14Qhp/ZpDAUY2wpzrvByYVyAuF4lhPLXVho45sSdx4
tvhz1kgIyOEUkC/VQwl9kX2bbMFdXvLRazuZf2dvzNBRUDh0jHwR+ajnosyR6Imv
KpjtAfzDxI8kK3ywK+hTKfnkbYEgIkRHtD2WZ3J6SgJY5b2Vx5n5LwqJP29SMflw
TwB7NDKJjznfnRnYWoYcL/d4pEktmQ5RDkXayOGamvA7NXeYlQCHk+nOb577vxRg
2wTttTTQDI1y3R69HqkaobTpsVsu5bApMHGM5Cy76KXmUdMW19i+7+Uk0eW2GwLF
ufVeqm2XjHDFToxK/24dQQ1C4nzzNyXTlZbP68xUgzuCFOobW5A8ZbXFTUZ30GVE
JYHCUZ9oiciE0UeEqrb6zeSiqTWWaFkOh38t2xUkUXnQ4MrEoRXKBsa3XTNrjDoY
/JsKz/B9xhDdQK+bHOmjyEoPycWFL8lBMPTHtrb4Oh2OT5CiUprBDYr2lxvNniYk
oJH945AwBjGFx6iGn8aMue+Pqyq2hIvqb4mUsCbZ8XzvOOQFzo7TZnt/6nAIaqSS
ZbV9qgScv+ErB79iCo+wfse4V3unDLMMN4caLI72Gxu3j/WF+Iyczawty9AJKnCz
KToHWvgcPx0lF8LJGAUmB8f31efapU6ORogI45CegftDv+XO1MniA2pDAywlYTfq
JjcGCEvLW94JUPQ340tZGVMGgkc2eWeM/RfAZt+o4lWmsndfwXdlJQEQS4Bqm7So
JAZuMBlvZi10dMre0jXA+LeB6cIY1SVS1bl5rf55EdeWolInXOiyYgs8DEGJ88sC
+O2PPuT2eR5SlXyTmJK+pNGfyJPrnRpJKxIua6GPGwzA/3gBPS3i7nbNc+k0ml9N
q+A+BPl2atoWz2PFs39kZCCkKf0uxsC12VbLlxwulFRMMNP2G0Xeu+Vsu4iMk06K
GS9fSKDlGR93ayrFAA4dca+7uTs/CVQV+gsufijNZcvrqRtsLxNr19XICtJvohxW
Fa4+LnItMCZcsY1cuMz1Yc1jp+n6AwyzhGsyQN3c10dGBsoofrJQRBlLl6fYCd4q
ArxkhdWFLqUotj+nfurFUKNicMuEuhZV8/GwTNlePBJeuYufLpPWT1Ukxe/YABEi
qfFRS2t/P+Br8hmN+Fpb4Y6KPb02Byw9BLotgNpxrVq7CGx67geU5zc1Z6XzjPn9
9QDGAFDpmNPA+QMqDxZjYUUmOIxHYS+fRCTU/cEZEI5yl2fhloTiXM8P35Kp8XAq
jI/a7Q/NriiZd3DfVKLkQaJuPA2yR6w3jpd6NMpJmrelpfQNtJ6OM2y1drdtQlvY
9Hb0h9T3FvBCn1C4MeBitlF5HuJA1sbF+HDWzSDEJshorl7lovRDrVCA2iYIkEtG
HHJCveI/O6CXeOH2EsV1A7GsVWrDjrhSwhrs7H5gu9iCstOyHX1GZyiaJ/GetvuV
r1cwxd4xuAxCWLty79N4EDd4WKqHiZezerezrJKvPZTAlmIvJMgSEo5yzh2slexI
pFHf2k9Jj7YVsXYXVLDbnmc8Dx/tQX2IdRCVS2kVov1QXABCEkuM1q8UtU1UwCBJ
xIEaqCDogzmcw9gv5PIU4OMsMwldCq3OSpKY3z7wB3Du/MQCoS6KpHOxgw1r0gvL
Ti2a5RTb39MdLjHNZpSfXn9gOyhCvFkHBoUhzv7aHorT74AJ3CMveVJ12RqOXZx1
FK4l/FYUb9rHDsb+DyI3wH+0IVXiGD4RimkxjpccaOI8dKfGlw0Zdtr/ReTZaxxr
aN0sMyoQEl6cSDsyZYnOotrHHPgBmrN3HncFLzDRZ2VhbQNm2HlS7cxhMlD3ePJ6
xbUfgOkBmydvJkpIQarI6PsFrwG2cdjvJcsXfZBqTzG6u1kaLf3DLJDrzW9FJw0q
oNJER3vzMFOlF/XX06eWTUNAU+DF6doPH7EbqqDqcCV8dObilvVzkkMDgFguLmLH
InjcZvdM4sPvn/JlRAVDLiSzUsQqkrWlSRuiCjv1F57oEKO87/KfgX4+g2jsCgBI
Yrusy4LYJADt8YlGVyUTiuKXczywITw+T8X7ZJc6WyJOzBl+2wYyAm9GjhjgK/dC
rYAavtXwEPU9gp3SBPU7SQuYUKck1ccHSwWp+uqFP0WCxsSfqPMfYJL7lU8Gskqa
YL2DcfizkUGua5HoVWSM8Bw4WMaokuKPm3YzSdMGcO5VPi4Se421VVwqYQQ5IzH+
2SvkpRDIQ6apY7UtXCDp1ZVYzpJg9Oqo1BuToT+Q/1ehWPHMYTbk5GyWJAdaPhcC
tCzFyIHFyLP74Gq/BwTemx2Ziu04gBQ9A3kaEqnDSDl+sKzEhb+4s8vMZu8sHJII
r3RnEJdc8M6KU6z/br9b2bB00icsq4zsvN7fHUN3Z3cEftasNQBpt+HRTU4AZ/OX
yzie+Zdy9AKRvkr8i7SY3WDxc0pdTfJRiQd5COhW9aHaYKjonbJp6NsSSR/+8e4I
WiYPNOeAxEiZmWxgSqFu094Aa4iqKka5uzg4hKF+hOGHle8ppSuzMnHPGNoUcMIZ
XxwDa8D8s6q6miFo/5WeNdh9bq33GND+dmpuR2nd+IRoijINCxktl26kAr3vu5WO
WtuQEF+U6xj5svgRdOc+hkYUeOtWEzqdWyd6opXidxLB+Q24Qif1Fg7aQFlotduG
1lyCDKqZQwlxMyN3GpHyN3WQVlOFpdxY9bHee1uVUD96giTwbXL7jRpdnSiLAr+9
yv6JgDfbdmUHy0bwtVQ3kG2+tfdAPGIxmUKiLcOf8b1Pt/Rjg8KMhtkCBAZwqd19
A+qeEFYoAZG2sbn49kcyVgGLrq60I87loSIDWWcfmbgXGSOJTzvDQPCxn7Eth6mq
z8zWFZ8MGvj5mySlEReZYJEg0KDLEh0Ts1DT4AMaFFO5EK0ry7gMlyb5A43TpeaZ
Qcdr64EOkBoO18czBeZgU2eoONZi3wLfWbQNaxZBmtTvHO2ehoB1tpFPOJP0+jrX
bNeFRltzpUfHh5SHWdPYRWp6E3tfRi9iqjgzE9ztgzIKfyI6UamtO6yD1W0KVBp5
kyk0mNbEaqk3q2otV4C9Nd6ISqupNhaXdBfwWBia2lKKPMfuVrKWtvQFBb4Cu2NV
PmdTsY3+MY4+C4R1ktFhy9cnYquO3y1wp9U+mcBYCBofNXZXX2jeTD4pA8xxpVPl
3EOcA152Rg1kydlqI4RzWLhFs0t/SqvvEDSiwUD7yg0F6xQIj2qmD+lAl2V2OQvE
wJrkB+b/SrHvEGR6ZxD8xaz0BhfMGlCqhloEvamfsE5TqfeB6+hQta/MIXMtJf8/
VGJ7HMDS+FSayE+Xhq0P16tVPStQvvphOp73+kDkoa/lG5B9B9zkEs3V5nL5y7Em
J9yjX+h1qwbv0f5/6d0ZYj6d4RIBrw7BSpcWX9nOqTCtjLWiobVEZFQzEdWOj796
c13UX+0QC6O3N5nsjnA2SvQR+sQ0ZWNc9Cdyi4xGCgd96AUrhM5sqC17gmDEuI7D
+uqgujXUU92bvco/nFrdB++qnP+WTsU7IhvwWpwuiV2DCriegZ9kyO9C12VDbjb+
UGcelbeqyuDaEQVUgUQgFjQV24ai5Nl2s5XaMEeyXVPGNeM4/cMze3TBRRb7UHIl
PWrOYNEAMLXPcW9RWhDq3tIkIWQTgnykPBxGkyaf3LtFSu2VywkwCRbgxfv9M/MO
bTRVwwYhjJ09AIWNRyha3SvlaEsWV/VK5Yk+DR53lOr3JnQECZh4ufP6nkrbeNWr
T1LvfgeS5ROl4dA+LeXMYJQafYwYB41psNFfhbpbR7AeDn1p4ovHuVKNcp1QxkJO
qsnxbRKfPF9QmwOYXc1q1ajxnxquAtaXc4YXt+keaKbkK/ift/uvzefmuVwcTomx
6YE5RQh05Gwd9r8rsT6dfMENWgchDSYO/mTUUI6iA4lTlyj1LD84rY20mLmOK3j/
6NC593dQS6SaQhvagkRiBIIL2tVtzmEuwM7MWs2CQLSseCYfiWJWWBveBkXACqb4
4FTQiHRj/VEyRVe5lNOnhhWPCcm/TpsSHNd91GcOwq2tLuOD/Y12zZUQwmpzcpe9
SI9Ta97F0JZ7nx+0XHuX2STQtkQfuClFrgOQJMcygb56XgW3e9Sq1A+qkFF+1HuR
z4bfg+74AyXC82uCgEvoj6h3eFXMIa804oeK8zDUxi3JHO5R0opr5/oEMce94VDr
0Fjf8lkuGwG0CTyuTgShw86V5ilMW8tFwGL5Fe6//0xWu55ag80gAjwHyKCGQyKk
iGWzTaK31cDpdugox6GNDae4CNqrJOvXCTv/vCOW018a8J3Mi8J0T1Qc253I+3pk
gRrF+CrsEToyq/AxbW00yLnGJ01CcDsI1vFSBB/92amDfGP+xxghxfCEh/bWJ7WU
6sKL9ztFt/BmDQ3uavNfwvyUZoMDyoel69i3PA/1HpNeaarGP1IYHlWmaWnyQM6C
7nSIq0HoD1CTiSg65C4xN+pbhbNvoSZW3R8sJXqrAnT9B9crL9EW375hUWq1kYFC
ROWoQxzVw151ZB8DHlLhtUDQ8urACSs2AS5d+fHX+1El2OprroIHA+EMWW2Gyr1I
hbHRS7pTALmlDaIcRKZ92cKQ3AtcKeaBOUtH0zf+zY4xHZnBV1WK3q8EvpIjFsWl
JcrEVjGCHfo+rcNhneeEbmcv41POS1eLp79tu1WtuEyu0bAIJt7eIdpnOEn7Llqf
u9rWRqSHNmE2HxjQJ0p6B/w9U/IxGn4F1bZMCtx+9TImDuY2rJlUOErJryBLkbp5
LeUV+hVtE3FuAGZrtB2aBIVo+wIO2S3vtcpXmaoNP0+YD2+i21oJBX+49ma+O7kP
WHlVoKqV2q81DKfT9KWIrVQZ6hAl7MwMdxSLePfdMfhPSx65fkGGrybcRx9zkVLN
Nc9720JfOuRZr7+/zUMJlySZPl0YvqL/EwNrv6LMewYEMc+6MWweyYEJJ1X+nbuS
vCxZ0oP9JoPYOXrT425aWywSjAUmA6skaqBXOsH/zJi4bMIOuXR+XO+tfoys6Tdw
hZLPfY+wUaiNhxJaTytARX8C6IuSuamVdFyCI+CY0AHkjxQP2a9YzrHJfTwfvQV8
OKLWAkmnB6F+YrZpoVAAUJr4ErGml42AX8nrehXhBtoKY+865IMM6zUI14pjt3kV
G4o+Qs1rEzoiGgIG9VcQpJJpwBpi+XYQJZHUCY9lN1Lv7rtnkGl0oJ3uVR8DP3z8
Ub5tFiLqOmDrtKLAB3GlJSML7fho9zARNHqzDo6C7qqu7K29KTElmNd4qBExy8oT
e3ikteuIVBCiFExg8dyEf+YVo2E6LttbSFLXnHnxvsvsn3Q9oC0xgcCBhhGgeqJ8
awHZwG4N5PKsgWB5ohRVsSB3Z/AOMKBNrCZ9A1Jn7hjpBqWBbbllBtEBtoUSe1hI
6FN2XrAvjiNGIj5FZdtJ1b9cnVnRkY8j0Hq0xzOX+Mx1Ls0oDQsVCqreYxZU1A8w
Bd/UIiDdXGthW65ord3Wfj5UVIT33L++ZI8oOMj1zF/tLoNSHUgjs/z3Jz0F5EkR
skZ0HlyRcz20TqvF72gOkOwfzzCpa5ZKzEAxBCTdfsRnF78nO4DAJGY2t/Nc+S65
akNsWbw2SIEoLTvXYxsvmSG1lT1eIq8/DeGXvali4N86DqckE3bBym4C8cyy7/gh
eJoOvN40AG+kFwaoJt31JfHEHQDS+HR4yAgTg6QfNk3Ws3mik5GYXsF98CAk3Vy2
NrtfcfbYRb8i0CaRVGB0o4iUyU17q7aTYWBBvAE5UgiTFn3zkhpRB5U/+Qjk7ePy
VjyZiz0g/llpYkR0dg9htHYYk+7sQ7W0nyIalzNs2qxgNUzVtSFu3q8KCHAGc+o4
1AFlhqIBfyty8C2H023G9bScMSr5AnfzZIqvE1MzVfXXnceNbG4ZN7qvFLBe245w
nxniQqhTVTrM9vsS4tBHSVrh/pqpijazNo0xA3fVA9ypvBf7mrHN+wUd+XzTAjxr
cLKIekFEYh2Tft3mFVHNT1BORuxLw7rzpVgXw5xkQobP2XQd/ceEJzSSwPBlGXvb
uauvFZrAwaIH+4ugNbcaf8ulsxMWGgkubTbEjnXVLH78DeP7rHVBDi0mEQQdMPQi
9MRPEKNZTBAB7RTbxdFnFDBo7M/ek9Y5mjoaR6BjT7warQIMqj6Vg3KlS5IumqLX
JCNrZR8Ss+Q07ptFBQBevjSIXLIZ6IWsdr0kxT8znsTI7/rRXXATvVO9e1Skq0V/
aWtKJR3cd/PsmfUWCr8Lbxoh143SmjnWGz6CBi6kcZRWCTmH2ryoGnJpmnhLXl1V
hz99ayR0c3ADWDkMrocnA4XFxBDnNT3ijpA19MONMCzoE7BX6VPeHS98/MS6Zo5q
ZxQ9u5jB6VmkTMA/DTXP6zPrKk5iz7e/hbg7GJsqW2FVMulI5VKkdxXI1FAIK08o
uKMkXypEU1IByMStD22vvIGdnV+gYEvwxsWhAH8XF/qaUVyvkQRyDFcQwNVhEuhc
q0h9lNMB6RutJj62KRrgpDK1xgXSguhylCRRgjEyjZTQmCJmXG7y1GgxMv44VCF0
aUWRbSJQast2LrnrtygopaQqVqwd+8jiS1LX7A3W720ke0JFbO/eiAoyju/maaOu
eAOjKwJc3VIkjPT+5D73TyFHemZOqQsRlRdQvKu5WqRBRORa5UFdxwuAyimY+2f6
vJNH7/9QCL06KRKNvr1LTuIyHr86jXIBHoiXaFdAqYnlPqwevbg+X9O8i1tp/VcS
oQob3c+aWxj7ks+AYnXAgoQYR6M/PonO3aiAdcPCWsJPg8h5wAzyRErH3zv70wSj
zYi40+olVHOfYPZhFKpMte0om4/8aXGpr/FeSTN7NOOQvGZxlNpHAPycoMaSVsQP
M1rXCEdPMiESJugfrbDoEGCnC33uQVheqv5GEZeSnvCAVep4a9lpjJM2CBK/pfGI
ex6Wi22+ebguayilx28gWnFvDvPBvW0TVg4R5XuZtIN+ZDJQ+o5GbDNqQiO2kuTe
3mcHAGlJaM5msV8RDXPbguEF4nQBjVmyWw+yXXFAktxorELxtC6oYubNOjnU7ibL
dK7j0isDMQHLrkLFzRaUtQscOeAgjSgxJ34W+CWJBYS0kvp+SHpC8mrMc2meOeVe
t/J3mCSg9Cph04SSjla9TlGrCO1RIOgFEycrQP9nDvUpe/txtazX21ZBReD6nOHo
rjxNfwqS2OpdXMuRLmCyR+JBC4ShlXJyh/U2rCOdJmNpQw3q6PMh4SDzAp3UW2MD
yHnKxX3sr6tfgR97oNiMm1Ur2Pr/GFElgeYENUB6BWb+SDI2/oh6JzXA/zzFTAog
GASEv9eIylUuhNUYBSFzWZJWfNX0MBmhYX2oVvuQRNFEHB5IGaX1KitNz30jkqVz
qwreDic2MkEVUbIGMIiu0FaYAuW5nJDZ0fJutt6mMl7atamfWwASkft5VE1snTPb
EwZhaaWfWFEeptYr/181YeKxPv7eRv7YFz9VPVvpfcMUfmKD8YkmpAigupx98CUg
m/SVHLAX6S5Fkb8p+7mK8sZ7ZBnxGs7qy/8nzLz3pOUoyVHjI1GFMg/QP7vyYnYG
KjHmA/vOQqkAKvFvTy4s+BCD2BhmNOT6CTa1HkI81ugj3vAwpOTuaUU9VDMlxlv1
CLfjWOpPcYrx4k48x2bAKB5kFMBRylJ7AVG0y9In0SQwlD/QnM8qzEUHY7nsVQN2
e4hhFBWSWfypDhMiwwHFEhk3OaU3q9UfHSqlAtZszl745vCvi+FpC/kYedokKtYX
VW1uMnDobjva4l+ywbjVaB5yio7EoQxahgCSu3k0keVb337IK9aIx85EK3npUtqI
oL/jvqEKR6tOEfaBOPIfN96JwxfsZg1LszMiGzsdcx3PQdiSTqxNxaiNScCWBdjh
VBn8XR1fmWG2HxwHPRQM6IQ2htVQNTJooaVhqBuvpQ0AabbXk6GitJy0Pd7IP+ac
p6kaXM6H02T6kt+SXzhBGiHGxZb3BQe3q0CuKxVtI68+/Z3jfOsSW6xRUmfTX04M
p1XEbkRSsRSUXuEC19F0vUlu2LU0Z/cWsG5dt+jqrbnJorn5s/4OI7K4IrU2SFy8
JaEHah6jqMJENtQ4nbBPFysNzoWmz9hGWVopwXsM7tCk2Wp9wL+9H83AHzfOo/xH
q3llzM6+PX2Di1ZNV1YR7RdUEI8x6odtaW2l0n4RX9wR3Oye3JuoSl90GHp7WbBn
+q2C/rop8B8V3GbLjBekbwkfa/EydnZzH4rclXLpCWDl3wuuo1HU9K0QDBwpaz7g
CUL5fE+YeqtmQRRdgyjboEOUjAupW7FD1BohRCo8llzacGMDssB6uO5VqOWkhydD
lBtV1SclDX9AmKxgHXIFFEspWndoo+5HLzbN/cu/23tLrOXiPkSAnxZnCYVD7xQD
iwhF1R8OnVohlwAhwc8+hn9+YzKZoqpPrl5N8hX8Dm0FoAA0FtAaEsftpO7GGY5E
zTyx7PlMbXrZpgNyhioRKM+w65NgV+/aNJ2PnexiMf9DYQvSd9P8cKxmtj6Nu6Up
Z3XpEIuysH2Pk0bsonyZN0s7al0c68vC3cnqs8Glwf6F4F2oYOe01uwU5PdXExzZ
bPJjiXC5RTNYV/+KrbixT0YiXgft4jazYtKqzRC1a7aDd0X5eLvjLKVHi31qN2S+
uXng0CHKpum9F5PG6bo447z6c53kUAhbqlbEJSwPr2cs7rNPq+5Ii2zJ9mnO4DBr
FogWy7jYfeLd8NtzdPwpfA5DBBYJT/7y5BFKk7blUBG8UzFAAxSnwjj2O++x3qAO
22C7ks2w/Ozhbgu0ZCh6U2a2KX364hDWMdt0MPekDC1XJYCXDd5m9QnaO4T707GQ
pt43f7eeM8YeOoBLSZmosHamP1fECwdqvfp3A/jmsQTmtzzKBomHg4z3B1A+c9k/
2hW86MHaDUWFHxWwGmx6wb7iHuUXvnYriBcmPl7tL4gW3+meZscFvU+E0ssVpfPj
QN+MabS9JSp83c/YGZZdwxvIqc/9uh0ZvMXBBxtPYuPqXAr2p3Qy4CgFXNWBjluV
v80MnDAkWWmBX7PYtuEworQkiQP/b4a6RnWxu6kaIPkDzSwEP+G/FL3L7z7pXXBg
B5T8keeidK/v9jeqxAaBwi0GSgUwiuXNnV3d6ukncfp9/xgpQEKLItvkLfZtTcHg
mzLoR82X412MB/CxFeVmIZ1gkEA5bBC2A9YriF0ahUsHNjy9X7ZwunZVKsmxWVYK
C3/xYqwMeI8S5qQSG1P0RlxO+c1+x/AC2jStOVTR3+BlSp+xNJI6/mByq38L7D8u
8VzdNhXjOjb7TW71nV/3eFRLenbCHIDuYFS1n0UUyyCisrndcry9FecxKNLX3nut
unrJ8EEBkxCk7g9LLHWEuIyxNDXT4pfSWAFSKAhMXebRvcyijq1l9UB7f6GOZSgY
U7/8TYF0ZL7M+Gi9WK/wW/90mJ4zbQOaZMucfzuLZwe+a85/aNzNZsTYXhZPbmod
m/l4PY+xusAHJTiuk+1EX9AorLFYI+cJmbyt5QIyjihfSD/FPi6vsfExnMvJkh/g
iASE9DWOVLsUtn6VoTZZQrpBDiQHPQIkVb+lLjpHBhznOWjc+/5ZbO/jWuwuTkFQ
y+wm2wWyFpPlj2cT2WTQ7/m54E17aKFgbQ4M13EVLVmnpPbAbS1r/kDGmqvsUPsq
HJ/kg+uoQmNclK9CZDJC/U8Ln0uH+5+Q9/K5PeZ2L/EptSdpXdcbSu4fa1yalBn/
hAY3G94SwwL7aUeLpZqqLbJ5rMXqMTzFIL/n1fOgw6F2ZK4qCBODlENOjUU5N4LW
/+R5qOuR8+krtRJFhwVOk0inh+XyZmZCMzh3TuxhIbOPhw2qWew968/gY2MuoGr/
oqVjmJnV+1c1BZcu7vN1o8tnW+87lloY+Zfi49Q6+FZXPiOALLpSOdokvaWbZMcj
LBnUdvRH+t/HeGjlWS7Xa5VbnMufqc6Hs5Os10grdVcXbv7eXbs9M35rZrIgbOEA
MgGC6/RtMpkaKUJrz+hrg2rqz1IIWvASlDiHgDwAKTBNOBzL5bwg6c6vc/eRsqk0
6Z8dSkNY9Vdv1ymn8i+tuP4N6YK5ZKu11VBovuy4raykBTogt5PxXzzdzkuXQzfe
dE47kc6iaKKUzsPrxWiFfauUMuXAFZR3XUqmUzBVvsVYbvAXlH2HzB8brj/fVt4r
QjxEqIPRxO1eNy34RttaQ24Q/pYu+SxCUt1OuzdNRCxpz1iLGzJH5SC8PrdO7BTQ
dveKlqjPXq6pE7dm1s30+LKJfFy1Kncjwby/LQZFL8D5rl3wbGpEogNDgWfPAk2k
5SM+ByhGj5G8nvsh/x8alJefEn7lTobTrxI0S0JUzUlsdDb5P5gg23jIOChz1ybk
92Mrb3oZFnE049XncIl8FvxkNXhIIxjQvjtRGtSCuqcof9rtXLCh9QyZjR+3P3NT
x2LcklXW4+bApqAIhdCwZWVnBSaZb7/3yzxumHbqBPkA03+sT1F3SW53ThmJkYmb
IoXRdAnC8FfF/Q4lJhp6W8+4vj25HBFlglLTHD1cE2xCTm0PZqL6bYrj4AyWY9Sn
yHGRkCaWN9hwArmBy/QdKWtIo1SKv0ToQ+hk4ntUIoFO/UHNDb9x1YdcU9vs+AJd
9xV2v7zcMF2TySV9r1IyPWOer1OCR1ictlai7eOR0jq72pVQfoHUdDwIXjSryBrw
Amtr2UD4OVpV07ObwL4sGKz6tJiPVS2+lJ15GUNhSwX09otZTK92OPnNTGRgW+Dh
PpGaz62DuSrgUNzlN2lE3N3/idxGULNEnRAhnqooLGWsmSqCd2HSufNLzIDB42cv
y+tk0JlZ9HGDwcCU9mhNiQvaef7un4HF+niK/lJL/SlGA5DHvtHvT+gHpGq/C6XG
ZdJebVZMjpjTBpGqRhsdmzdN1C/7jRiropFNJSG222nZTiQe5lcUWCDBm9XdTWTp
L091kQ36cCCsc7q0xPP4DvX+EXRexNeSyIcnMkS/Myg9jTBQ0RuNg73oe1Z8AzSW
F1XksQccczMPfT4aLMMWUcFPWrvXQA4jxWrHyQzgujeldK295Oqbhi0CFQUf2UCF
pkwpRNuFfMj7h1Pxgcqnkf45O7tfjYDyczz7IEi4qswNcljRh3OrD3s37GXoo3sk
O5Dh0/ydSi6h94qzNpWOiukU9eJbUWf/l6xAIDuHy9tV0HLprfjX1zbmsYew9Gni
r9cOhWV7ruxMOuvh0O72LpcHIHAbfmY1hX1tXAuQ0zfcePvuYGeR9u+IYkl2rrC2
jmg51O/NS0Kr11luOp1UI8etMebS+jEsnElaxMsNhaqA9Ere9C0KN/fw6mWTq0fz
IsZ3lmeMcOeZ3ceZOg6xHhYtTig8qZo4LkB+5FnWk4WFCFiXonhaAn4w5VDC7rdV
GCza0pbFsCAgPRSe89qmF/cLHzzAUSDYTDyu+B8XCWfOG+xAXmQMJZnRsmLYW7N+
Y9fW/vZ/nXkLNQ8c9hODV6XICq+kJLfjKzkqCM3+KJixf/UuthZG/W3QXf2LNHh7
2Sl/NpgtwWWYgdgV+C6a1S+RuDuJlVwdfIraRS2YA22T9+h9ziBcRwH2bJHpm0QK
GQtwgFMhK01Btg97e/8Nmrvj435L+osxEqeAoQL959lFBIimhPCGoNL+x4SsV/C8
2vHylvI3wTYEn54JwrbMVpxeTo/h3qv73S3SV3yMbXLoTIbrjoaYWCeOHbvYpt3f
hJYFLsYEcq/OwWz6cwMG+8QLGxweNSD/9Yw7oPLH+tyfTw/Mfp8dH+gP99KkGPA1
Lq4IxwFxuOkt8PLxAEGOvsIcJa12hyUreNYR9pB5b8zLG+rnOtXvTf3/OH4aHyjs
z4cEJh+n5wJ55Y2hEx8o/IFaSsDxHQfLF6xQab65D5RsLuUoWulXn1Qr8WA7XWH4
p4cZg/C0UdkDOScQbXV+yccilUiDVvV5MzNA66dQ6tPuKvizY3G+tpzw2lzozMdr
Mi7eqmRR2GdY55N/3+Wu7irUGgnegbDeYDbqfOYn568ePoMzz0TwaQnFS0VQb1t+
C4yMH2mICZBgyK4C5sL8HXwOCQhkVL+zVME63ZUSmnRyqd6aaI0Y91gPaQo6KR0b
6cdkbNU+ul97e7mJWU74KLTbwIwDh5q44xfC6YOUUvoDpF7AUTb+1wEaWBFuVQcn
5e99CjfaTsV/3cA2aOiPdsLL++xC9jVRSrdtD54LvEbsseqkxcilfhur4YWjXjq6
S1D/NcOLlb+aNM6+S2wxNEjqwgpHOchiJEeqkyYZ8yGDtkb92FrAQmcSo/QZLaTF
j9gwzIK45Mz4wYQH5FTHqTHqNxLUGXA9trZj4CUAW9rzrGs1m555Xkmh0IYmrBpi
bY51l1MWVPS7638+on9VmFgixYPhWHY4dKCttAmFuHzsXES/t+nHr3qMCGiXCwSa
PeVZ0QDopQUscbBG6kIrMgpMMyMacXxnoapSmlD8gYnD5Yz8MqN8Co+8JpWUSOhk
3RE0eJRy0+qHWjEMm4SfJq93ZtAkLceVKc4wjS0LvJqtuUp//GpO//ni5h6tlrS/
jO9viHtOYreh0aLiHFw48G1HOk2qC2aRotESaa/5FNIB9Gu05+PmJZs630EWARtT
GQeaxMvOT4aWsNOX1gKWKNRM9ph7Tr7LjUGBHTIeQk8aRKpcLlF91HAiNE5qejsu
Pz9zedq+/TIiRQqQzUn+SOv1gahIBnMCPifNYF22D3qCVq5PF4qJEhIEzWPRlLDo
PI6SxaHOJu/+ph7KXuXG9XSVXDnw80gS9wSLFujiEl2OOPucdMU8A1uRI/TTIvh/
avNXcbLPcGwRBnIs1euoNqGCfvadahJOhdtLvDJ/ygI7/eQyYwk5Iu2VKAsYzIxv
3VXu5O59Kdku/mabDKERZSKaNeGW6GB+6RhLoDkZ3sgn0w9PonncZQTSz64ig4zS
qpqFZNLckRv+076tZvu1O78Y88vCgmrLLN+2sw6B2WbMUcQiLIZDL1otDSgY0GvB
E7agP1/VVSvFWBGYGIoh61C9oUWzFHCU+SGlFkWgwaqk99XSQy9vf7wLaDuscA5r
IRlDYwgV8SUwAg2C901yL5PTO6Dd2/k/oYYy0ENozlio8hOuDx4S/rWOH7DGt+Nl
DARwfCdRiBFQFOa0wIq/SfbQgmYH9pz2Xe+Sn5oYJBf2ittdyI3Vai2c9fAnjGeU
cOub5ObOY0ov2HwvLZkqw174q06FCOYgA2lhwZAgOKFSr2cxCAfA/WujzDGxBFx7
dRURW1FvEH8eYiMwoBbQNpSHmI5XMTEe3ntj0izUxrb4IW53Sv5NyH95RTfED4HT
QXGdO252CJgbLNmj54rqAQPHjdoYLLRKkuFxTewvJiIPbaQ7ZOTsjD4X7SE3Dk4j
XrXA4p5ImxCSe01L0YzPGsHyhxd6mmQshevh9F8EEW+wAvnCkO3v3k649d3lVqIk
UlZfTsEny1FnwaPciDdSxCTpbUBlOBVq4Nz14wnmk8nPBwo3o/OGJSJCyPXT9YTH
plY4ZBKVWE+Q3pwCsUaP0ooQ1v9QWSiX8Fc5C6ESy6Czk0c2Wbcg2X1xe4hsDoeJ
BwREORShZwTZByqBd3w/7VW2ZcXYZc6NRfyVlu8T9dHOVus5T0BKE4I78gg74j4V
o8n/Z6AXR82XcOWiVJnd3AZfKmVP2tqjwaC0OxAL98s7T0ArMkPMoPsVcGWV5ZbV
q+i11XDGARbIgnSezGFg40iIKbWeDx2YXOVqVHi2YB9mWU6gh+eBfAnZ0tqj1LU3
YWFdYHHJVF+tp0EW69oLI832qexljvd2YCAXGaiEnmstPhhwSa1KBXZF26/mzP/5
/jBUnsEB4i0FlWI9cCeZt0X8+rFwH+n5bNCv1lDsoz5CRT6Nd1Rtw5LM4A+mNVt7
HTeHR213HTz06YDTIksNR4WL2nzy3Z6QJlCL0ZiP15x94aSecTlbNxDbj+Ejiy4E
cKpSfMzOgqbUlpwTo+LkBbkozkZ+z3rcJySU5E9DR/a85LVf+QBiXJYOAB2fxG+4
ShfBCWkWeFuNxWQuss/TGEuMKS3KRqmg5AblDNPiBGKa11a38Kf6n9C3yksaAi1N
LRnKRKP5pUO4az5ALgeJ9JcPlLkV+ho9C06sGB+qMatzNCdBJ2zPUokWVcFACHKT
cAymBI7LV/ldXUJ9P5iuNaPJ28LfwNOLGpIwMRiLKbcU04JHZigsdzrEVEEJBGDr
2hDwYaPQT7ims0Czr0xwKMhWWgmuGuZ1QnDAT+C9SImtfaNebfuM/Iz1F2KNNO13
X38M4cMp7UEUJBb8MAUCYfNhU6gSSND7sm2qPsdXrn4R2CylMa3/FYepbCGowqH6
SQ3+pWYJv6MOQpKvf0O487YJkvuSQTsevACXl4yNZ7G59TsSRpM93GJ6oN8YLnTI
MrSO1YwDR3ety6gXpZouZebCHND/Bfk4CMrWfOG30m3bqqIqSt0IuHnPzC3IvBUz
Ho6/oeQfs3rmttmiMHHMU9/sjquzDGyikXPL3njTmRFfKSEb3575SPlq12KUee0+
y4sDLbIsDGUV8IqokCfIbyZj5d4MgqmVOjoOJHDmOdgjfufkS2zq500HwAhbJe7v
sE3WhDtWoeAFChHqL4vEJTfaMga5H7Tly0MbDCbnqoTVqKOoffhkiPDwpQ3tg3Cg
9I8+cKWdMpurAGX6WicsGKzcfIGfDnOAbySkxXBbqKgdyyWB/faf+wahDQwLNQ7h
00Hchqc6XPZEOHZTt8Ydblsn6FKwm2GX04zRsApg8IBK/0nP5FBRsvhZwJiLDCQJ
BfXKihL/5aGGUp6VgxLAtyJDYe1fI1XBi0inPsDiQxs4Nz0UUSRriaHY9l0i8y4E
kT/f+cDp9QMcAHSXQiC+icCX457Lx7QkydESAEe2uKrm4fdS8xBanJ66LbuZ0ZYZ
azgP8uFTXdthl4xQ/5Xd8Wz02Z0HVU+vNrEThw13pljhrbNKwbfEys83VBPWzqpT
7V7HfQl+tNA4zpB7tpc02QSh5CP7dsdDNtxYNn/jRIdFBfaYvNzqOpDd58JFaH3Q
IJnTpKcV33j/qPnYo5g6Y/RZw1rSD7lKO+A08zfLC0eIaP4z59FwMtjBfJM1KH73
VA95+76GX9KpivtyJTBJNoUr78h/Wy/9MCfMPljn0BDCpHV4avLjIMJ3asJxEt6P
YozPiXpTZ6cFhs9v8ERt0JKZhb+k8AYPgVcdcftWVUYd63NvZdWISvMS9r8hzmfN
2TmXrPnzziVfr89njARkDuW1G7wZrWuaKlyGk3Nxk9c20/R6nuEW1l1TsRl9LF0R
bKwKFIqLW7SnzYfWDwIPGItO2qDAhjJ6Oa7JnOm4KOYXbn2+H6XIKk4PRIFayO08
Pxdd7+E13Oo7lDdCn30BAEono3lEM6l1Vw54QvZTTFZ950ZcuARgMQv8KTVreWO1
gMDLIxIoknbzRwQkpNYRs/6OGhSqE6YBIQxOOr8wVMEDsshCd54ko+udfF/b/MWw
OPU/6onnF3ZHWKG9+r4n5ZsgzGItphBLusqJpxs2kMpG2eXROwDX0HEIVioZn3Bq
EHLMaA6CKgtnEDx+B3mZma/AoGROhkOPIqzEw3qwL46ojF+Fm1boMF6dAzAEEL23
mkbFfKs89q1Au2Vn7o0aBAWPJFqKUrwmMGfIt3KMXiZXLDf+XDEwVHi2pZ4/9VqC
5ZlQt+zaz9pVHgEwBpNl4E0npT388St8olP7KNIxKp/o/pRdHDsTAuf9UEyd1Obf
A1EYgEx1IKbXHxJEgSXhMtZg2oPIb5d2DxDHxUHv2/o4Hm9utyTlrXp5/MzNgjZl
0puMuo/BSJy+nZ6JnuR9uavdGCSJBnpEE1kk4JzvnU4gkdCIsOFRJotJ/9M/jmbc
Ia+C+EChhorM1oi5kpCTf6264XrW8/5hDh/aFMOGJDmkJpQ5wRyCTdf8w7lEXzXl
nVZr9wdfZ99JI+XUBm1xhZVqSfvNYOZhsmRgVlkWnHhMSababSyuBYc/Y8Qhhdz/
lg+Xj+m32em8eGexaJrxCNOX5qZxCHzMogcNdx3TcknZtvg8regWprOnrc0wvsWk
iMLeXMp9g4f8kE+J5FcC5hH1QEyuupdWjQgPOVoj1LWqv0y1AE1V8rkYY/3GKTmA
aqdI2t6PyMOG5ZSKMEWvg6PjJVg86F0eVD75Lvrwy5azvdbwO5CNn8K67bYKS82I
LLGZWynTTUg14O5lyt1eawE/hTFj0XTSteg18BF/n2vBJ+7vGA1UEI7Y0sljquHS
IDQDC8mdvQWC6+vJ4JAljgFswlSAPTp5+3ch1RLNnHRulqULS+ve5msR4C2bfzGM
uwnSVoRzMnIXSDxfgfdjKRKMYu9vTevyw+wPUZwmosYd0QU1EafDuUgvC5Lhz2Ce
cutvxWDydYZh7Bv+19CxmI2rXj89U4WIq9SjFtrE/6ivknGvTHmtQLGMtBYkxzBB
W1bmmjLPgbETfXFnQalBGqOUk7X0IEXZUCgHHdNLswECrTFG6SD984x20oXZoZFI
u0AcadNddquC7OV09/baxWZ1+Dr3DlCXZOc2gqXDjHEq+CyzAJuwlMtArM3s+Dfc
cdNzoXlQJ2vDDuXBUOWURTQkMn6OC6wl+3gOAANzZdNpAR5Hn03Od2U2N+/QXX9F
2TQtym7G+J71loqZfrKVNVoLXq8KOtDREqBP5OlBZBAxH1d3m7Wk4HRnC+TYEhUC
8wML3DMiw7/TaHlEHOssFUeiGzzm5PXNI7jTLFoH2CAFbrZ7C/j7IveSvPRSE1Mv
pmOm+ZkTLgNjPrDHtzzsrhw/wB2MAHA7WPt5h5MjLX8KdFXaiPiNqDcQrgt0rFKp
VPpUxyAcC1u0vSBU7ol2FSwIqmB5dWpmMZC8k0bkwZ4bLSmRMNmsvxn56pexL2q6
WQ7/o/4WMdzU2WqqApUaEBzounkVXacgrpldYK83RHTYoI/xNWM5d2v8ov5iYOwJ
ZHKFug1Zd2SctXTsiKwiFRh1WhpMWSodX+t/b25SLA8hpTxs5xQHXv3ozns1RmER
JvxCvfawPnLroKcSNDpu1aB5iLoVuhImP/28VrCntywSZjwVlvMPzjx/JunHq9UI
OVTXuw0khbdYh6CPJefCW1/R7W9kNEPnM8AZdujvB9gEOMI4UL05rmLsj6B2evtJ
p2a4AgZNr2bgK9F4H/4eUsWd51+IBN9KcqzNwdJUytSD0UMMvThCRW5+pqikHPBN
r561gVUCQ90d5z/qc71RignPm9+HOksNGLt1uWjbD+TyM23w81Qj+8YJc/P9ZGRx
h33yeeVpuVZCRMESarY9YQjddPd6NHQUKPSydwoG8uVut1lkjP6bfOvLk+9iawTG
pMgTpILpPNY841mlAzZU/aHmTc81IcVrgKew6QL+83N31B456S4IVGu66rAx2nNI
zz1l1RVOom4+wMmfdrLSy8o2Zkw81l+Q6WhIqRrmf8UHSijLw4xyxMtLI7hIA8pi
5UAiM4nRRLrgFBGftDYplPlzBXqsFCcxWmCsg7zWzWHzJfBLfv0v6G8W7oeVZ7bG
nBiegXUVkFuacoE2R6KBLI472iZ2dNwwevEHFa3rc87WLAT13aUcdr31C6RvbJMl
Dlnpd7xrZWBC3B1ox6Zhv5hkGmQ+8qiiEgT1oXas1u+TTU9/u6Da7mKq1i7xMCUX
qjQ7Gussw0VGjcQJ1McpVB8YQPnnvBi1QhOm8nGe2+TsRenhW8aFqD45AqUM97fN
aL8fuF4YWwVrWw5becDOXXbCqSzysc00qm5VPRvh3UHjcwvWawDMcgNH6C0MRLIH
pzN29943W23Sjb7h+AjjiVN2WjQGIW2uHr/ucU15VafnjZCMhP1kYw7HZp5gCqcH
Lwd3XWyTLE6IxyUxAf472fZV3hctu0lRnQrf0dHtF0LtVMRTZnnso1Lbg+8HfRaM
MNyeMSlGBSgs0PFGWY+Cmz1/xb8/Vrrce+QzOURMsUB84uPKPzq9RIyyIYRq2u6X
QrlEk5ZqiK8UKNp6+2WyS29Z2nCC5coQZCKX6s+IqB0yBp5NrJX0rc/fqO9vRW7e
QD8ja+mhqzJt4mgeBIMarOtS25zOkuhNy6lKOe4jf5eM18dl60a81kaeIHxxcYC8
nw5369ffatCqjalTZOwMggUsx32buXGH1Wm0pZUA0XgHVQNPykPffJjDrqlbVe3G
FCBqn8+NTvtYQpgL3w2kA+QFHZEnfWhwKvkj4lNvNCXBNyl3GP3Ee/bQsSNFottt
cQ9EcordlVDewHlZlx4bG3G8KZiOYOz8L9OnlgJds40ELB+OqOqNrHQqYxh+i7U/
6rKhBCxVFh1hxec5wz5RL/tsx9VO1Mivwb859YV+nMjt5AS8Py3v3M8KrjbvliOF
3V+9Mbo7vkDa1B0kJtefqPST3ZoAwGWy8hVmtgfIqv7u+oSBK+RDRUOITHIrrvgu
u7Plb7GSp9tEl8aNchaUogN2Bd+N3VvgTHCTGR8MNMCEvIK4gYrXjhRjduNHnxG6
sfEbO2BSCGybfsjBJO4LGinzD3h2hjiAekvZrnnN+TxNkMFCO1jrcIG0FXYhavdM
St7WBt6XMWGLJkVMIvKI2OIpWb+HID8xzK5BZEthXYXsH34ru6oPgliUplESjifh
yv7FPXH/gdKNCKpVPyhTheHVQCu2/2o6XuzTDKL9VB8XfscYvolFJlLL4OFUV9v4
qm9nZDyUkAm/GIbSu5fliXhrjZ4lGrD63VnUTodhPi10MYCv+3Wcau0d56O/+PFa
D6bU5nG3qJIRNAVPn7lixGPdD5laM5jLckHKrju38nG2mVUemn3cC4GAXWjQheQ+
B0tkAonQhbu5G5pAIJSGQ+JprPTGCfygaw+pmsdrABkO02Rc/P9ip0bMbBxcfPfw
iH7O1A71YkbjFi4AVtdkgAPP1AmYZfQ+Y2kVwmnMBt+B2lc88LEN9eUT2haAg5ZS
jB1IfcM/OXJM3s5+kSLDFVBxQULwd8KoQxMvu52c/ft1X/mXoIARKcOe7gEb2xAD
thvxPdE5h8/uU9+pa35Kl2XvKRrlS4fuDxAyM1OLWLFxTSVd7iYrZk7vqLF4Wl+I
b0qwp58WDRSW5K3qow6QXr3bBm89z42KJzlZs/1bhCbz9Axdk4kKAHdLXYxtkTDN
++mF1hjnsmlI/eQQFQT+LmaxiMrQDswXducbs1jwEQpVGlzWnagHH4Vx+MBkPrB+
RLx+ukF42JdBKGv1IjIH39n9snSRwJ62O3Vhba8LR7Khjvatrk9jd9F1hsp9lktS
Ugz8l/bwcH+wZotqH2NC/TUfRWgKff4w15cO3eVCraLsCjINGGTZGH2Lz4xhjYHi
OnNz0Iy1YWzeTWFKqUsXOz1Cz0PKrIlyxGitcIbWPOgEMBB3JSeccun1nSNjUZsr
3ZEej75RmWfOtCGlthW1F6q9GDo30hj/Sb4HMi66+012aO1WnvD6HrFXw9Ibe/nh
q6AS+XFyU+ErSKapZokoT5+jsmMAFY0Ne5shTILG/82h8mK23GLwdhxKYbgKgWZz
43Dj57XDDhfpX+6qrTzwPz1eKxj0sHyWprCxh6UtwDESl50CNmQOPVClFCkXBTvY
dEtW1EEHS/Dz58zkd3HZYTdGeYLAcHYif4Srd3igNmu45XJjSrcUijeH0jXoqati
i2IDXUig/loYVCL/+BcVwF6B21WuvqlkVCi/3nxXVFZE2f5Vl9wroYCaAr2iJtgS
UuXsIUCIUrdtlHqcMSObes6Hcf2dO0gbCqMcGJRZxmH/a0gfG74WtGCc3bDLxYIL
60jJrcD7B0R4Alqvp+/1GOUfUMXP7OOLDMdKaMmzXUzw/r+93aMKeGuVUqLHRijN
Y8paaU52SqkrClCZQHJB3GY+4fRBnW8t3cxfp8tHRlWWie0VmWqdsp/5RC7UZd8c
8F7n7Y2hf1mMygHXaZnnJQ65IHJaQ92yWmLkpzbAF18JtkHpRKTtaE81NOIFH9zI
lRFNzktjFzD6JKdukXLhsLryjaEqyO6B4VyRSeQ/1V22g1Uaqe8PGRFwBc2qpjKc
Q5+b0MVYbl9RKdnxaVIpErdpKywyExjbwSfSy0Q62WqCduwQ9RhR85BsPBCcJc+O
SCcmuLUZROf82J1YczMyZrvW7wa9cvPw7nPS/Y5tFsRMUyvAPBEhYDYzGJZOEkN4
XvRZdm+aSTeAOMtFd1nZHQvrFqj2tEhj520SYsLQYoH5r69kx4dzZgD4BhsSDGdR
vtADFyC/Omw514nj6fsCOX/EInGKJSr+aK/bvlHJzubYDdZhcmTU3VOOaXWAji+K
dLbYnkF89bOfXkb2VOlgZ9DfApi4pTq/ibChqhBrQqFRj5dBHGVCN+7h4FLU+MYX
INEVy3zfqz6CksKKuHiHpFESCKDFqoRl/+RUvuquEKdsswDqtJLGdP++YdD/N02A
n0WP3UPMFBcTWEue4O5rjeoW/zcP5gzC2oLifN8izxO6Cvz4PcHC7Khkrd8q10DX
fwH7s0Ags+YkcKRcDuE2w4h7fO2+t0PCFN/qJVU30UHRsVSl/WK8y8BZT474JNig
dG1Qf1IBNbMvmFOqEzxfGz/JUUf3DO1kkT9MV0A7ePI6qtt4f4yr1Wm/F4jcPJPO
s0GMA2Dx0lJUM+Uq1FTo/a/tx5YMETjqQ/BXCXf+vTgMLYnp7vsVSFOmQ1qnuz0o
GcKkkeZKMP1TIUCzjgW8ZTzsE01nWy15SfF0LrxRv0XM+PDRX51dF7Lfjqb/f4bR
58WLlq0354J6QGkYrLfIH4CLbkFofQj0fqPVKaRolBC8wcpEI2l/D3YPwVNS3G/K
Pp7m6eWwETeBCzrlFjhu/7db/ckJnyBS+GT2/LzH9d7IXA71XZ2T2gjIk3RkkU0j
PZitfp3SWkdr/gC1WdZ3IXVOo3LcdsLz5jxk1EnXqxgLByI+OKyBaKLOOKn/rC/I
dzDMqQVX68Y69LAAcFakvmeZHWVNH9jg3e+l2gQIpL7ulHZSWdKLDtIEveVGqLWW
y+LQdWjxXjtqsSDwZfczPQ98VRZlpZi9hy+5WQwHpOA5YqUfT2FyjoeFP7I4LYmv
RufmGCuIM5pVdecvVWLgG+hID3dUwkDYcw6+rKgieMH7A4LB5KDoHHwscIW0NO8O
nKxl9djMvctEpNjJ4UevmzqKdkqzZQLGb9LAp6j8I/LJNuXwvlKHiuEcrKNxiQcv
T0LRX3A8LGxTxqyPsHUi+u+xmU5ZWraKn6lY14gbt1pHJepB7KZCio2WF7SuCzvk
I+q6oUcfQnkP1wp9CC748WC5s4Hf2kxQNYpmbBX7HZPxqgBrl6EeYEMnoyHR5OGF
abZzt2ysaTRCGIPc3KvTCq9H4By+qR/Hefv96S9eg5jyDjB78oYJCLg0goPGfGig
UeQLXLtWjFZzN5cTgjQa59WmKE+mDlYmoEbAb+yVigoVaCNUMdumwDOoY1NQzz1R
YrJgMkuF4A1fNJrKhfohs4E6mMst6Kjj0DQgzTb6JhT4Btn/3y/jAQhUvxU/8FOb
LtRMdk/oZ4N9Y5qFsJ4+qPB0KfkRH05hKP7u39eUevhmGhgr6+AsGO2rvaer4wFc
XuGdRAAphEfb2ZAXhj5tDdd77I40Vb67T2BVJFQX9H6KDHnbBEVT6T7mZwWbF47H
QBlnSes9GpxioEEydlS8kfYyP1H5LS3tgsF6aB7kAkUxRCDZ8yPlNQoifZNJw4ca
0ezvUBvC7JaemNUnoG5J+HNal9niwbU4OoDd41hdY1geJelZkSvh1Vovb2OCgFP8
lAhRIi2Lqi9jEsHyLeQOROT4xZn2LhBTKCnRUKONtSEw+/zicyCcRJXJVL1L12hc
n6AFMU7FM2ls9H9xcNBLn7E4CekN37Vhq6TM4Hd2T+U0s4udYqQl05Ymcv1e+o9n
Z7EOL52EJsxOWT1MTODQGIIHlNFFNwPS+6r45Qg88xYcac2dioDrGPB7K3a2snDB
W7QWsrv13VUCeGxA6MXmpwgcJy++Gmp+5lQnhA7azo8hdw6t8uhxq/aRnjEFjAZk
4JQ5E8+Tg2uZq2SJmJpXeqsbbKbwZFPaK7fnWjJ6BUdpacRj1Z3a0Y2qmVeun+EH
6wxLrIuG4Ccn79UxPBQdYn0lZA+Hmfdink2z8EjUyixXX3cLNGhJ1tv+CgZ4nYeF
qW3FO7iXbsfFMgZEyRjwEzu7ZLhc048jDCPDoNHbsUk5c10Bey+fIMBQME5EDD0A
+rxr9c23/ZNvBClOlNPqBTQXtnSmufXAC9gw1gQst812+/22e0OFF+Xx2muWypOi
i4NOClAfhlEILaQl0iP1ZF9s78PG3KIkOzY8Vx8OOJUGk0tPWZTPMXa3h0KqpJUj
sdPOuzy/T7987vsOWF27XQob2m0WIaQE9xSsexNMdyx+XsJsyDwlz/PMXNtpmu8i
tO4gpHYKz7o7LRZAbs2ZAT2Zki876KbSG23OK877HW0aqrRjpTSJFHlUmFZPwsdG
YOtQsNifxEgFbYXrHMJn1RrxGYAj7/elCfVoAmArQhVVvXhoUnet/g3H2UnqtTeI
FOs0GjJpNJGj0rEBbInvrBdwzGegffmhZwQrrAgMHUqML146U7iZxkd6d6VgNsrx
u8LDBbDrT2OFpHawP1M1tSc8vX3onTKn+SQHXsSQXI36foWhUzHz583LLa6o6Aqw
mjMmbyiZ1xry9yzmYh8B49p81AHXH8GlpGuLTMGXFdfSjLEALjCVbRYJNYMiGAye
HR3ocjKkCg6FrsJmI4SZUm0Zm/Njk8QYlEGNNaE8v6aC9MKzAbfdxQKJAwbdbXd3
jJHfeMe1csOCev1UbwtZsasbHsh59PLgqlIuEewymabHB3suy7SKlmViRZI+17X1
k2EO64A1xFFLwLtQrc0gUHN6L2ZIrjaUjtcJu0d+v/HxGuHASG3ZK1CvjjhmgghV
B9hvwUPPjsBBCBjBiSlrsi5Cf2tY699Pi75VHVQQDN1Mwhim9ONIlfKW79uWvTGK
bss3IT00P69EXvEeppAJQ2YxzEaE1nwq67shkfhSg1Ln77jZjdoGw9E7hGqnOlrH
yhwRq9GfbUkKsMceTp2UFp1DPGnu4ASwdNbIkfLba2Z8WppunGCHpLhAMcUiGd74
aQrE8cplx3RNUb7AxiZ7Ev8LAi0Cuh5oWfoS9yj6H1AX03TOoJ5tnQTinTIZ9FKJ
mscn2qCPQpGA6UuvDJ4l5FYvOXOBOQ97btT3Rmt1zzJEOu44TPSGbpKstvG0sTVo
L5niQ+1+JFSFlg/Ihq4wlVcFfmb7TxTeC5WnnTzin5XJIyHBAOcbm5BCN/RWLvRG
qL32BjZz3LCOh5ecL2dSmXzTU+kVHbvu+rhbmdN3lFL1+QbOMBBW/We1ZLKhHCTg
NtoiaWNj0sWaz2HgQcE2N7EFiCT+c3CeeAOBVE+T1lTzxAmPB7qoUy0JYEEPU8LP
O4V3d0kLwpcBJYVI0YksGmNy0FmyBSjVJ9ESXiLWwa7DKEWmdyUfYFnlUickSACg
WGizY6zLxfqdqJc0vF4rI/gGLsTweMOlZoyNEtzZ5sY6AofsduZM0N/HFw/CTBGi
5yeQy/EgwiuhiRuKYyF1hQ3/zjC3Ksolwc/BvrTqlk0CbeH18dsElPeZU8Qc2Ros
/ICiJREMTyg9+x93NJhUB5Bmfy4TaZkLoE173ZwIiSjw6HAV/NpBNM1tPhK2lY31
HuacjOVJ7c9sJJWiCIfEv9ChKpbNeAw9fpIt/eNXSF+tWVQ2YCpV4b3IQukqcDlw
BJALEuYOdDAUoKT2H7dfLfICmg5169r1Ktm88Bg6NDN4rjL73/MVW2brW+XCmHJ5
tysHSoQMtOPJfHG5WNpeEsN0ZDJVoCx1QET77ZXvVbZyaThkFMoDYF4eSIl80njL
CgB2znfDA2tpZ2YrcO4UmsZW7jdKQs87riSiIO5DnOw3Q68CqhOHkLPSUtjpo5aS
my8CcsJyk2kNBo62US1ZbvHf8f4btZI2iVCwjoTfprvKC1+o1XbFSehWQROWR951
LahIIvL+NFlmacxDoS+Y6XJ+rKdw5ps5tv6wLUCIunrP5kZCmk8wmWXtVajKYWkw
/l4gzr1YaSwfPx2DDlR7oQmf8qyluYfAXJR7medssHrdH54yhDfzFWj3tY4/7D5g
n5ckaM97hfwcq6YNwq34CJg6uvFAp38U7u8PrJ8U1uFl1o3NdW86DMyIDhixbvyd
A3SLOQqzIMy1E+Twf15BMi/Rj5qcbOhyqYJTleMibKc8z0Z8ytImB0ieYOTFly8E
NmGZy/I6Qhmaa1kbRw6pOlmzDK0lzmP8gry+wLnL3v6gFCw3AybL7CsUeC0CrgsY
5xhjb+FenIljrZ7y6nXXIbsCESOSNZRDNTjniT2gC5GaTZRPc/y1ErshmBfnfyZ/
Cdf0JbQ3pgnhnUVmg4vtDes6HepM+Q5JYTNSeacI+GhL8GkQ83dAH4mECv6VxBw4
uj8dq9xEPiu9tN75v0MnCYudjaJL8NF40g0Cs+WRsNx4SxxYJaQnnZTxWU0CpqGh
sDA+8SEVGmS7qoVV1pdqNtLWmz8qFQ4+4OVX2MxKDdx1LPP5AVj/EQLw9VWeSe7y
EQa9Fw4y6u79OgF32GAIkH+2krTxrtFp1nbqZtlAW66mp3MioXG3cFL47X8VITZw
3V5jze5b1Vt96pmehjMD5KNX1NzDbO/xwqp3+ErKiFXc7vX6zt1Cu/J9I76voyPb
5YvewerrOsf0GydiDb/UNzRxXXoTL6bECV1MG0myOC06CSf3Bo2l6vlL4HMGliib
1RycnzfZ7+ciiEUWLYB2rD1TWKyMKPnaKGTSNUQC/WO4xwxwr7yHg4qQKyFJuqc4
W1SWjWUPmW/yIZ9NCQvc132fYwO0ZehTGM1GWHBhT4XsWDEdXPMYdxszvaPRSGaY
j/OM6GIrZtvJbgY8hnIe5u30dyMee/hsAv2Ev1CqUMoyE14U0VVtaOaYAA7a/Tj9
+e3uMszKwUJgAaHQHQ3aw01P1DlPDKJb33ETudajR+ogLge9KhjqUpxg3grnvwBs
z9N8teGFeh5Ri0RSZyovTNyun3TJIcCH2uorhyiW97tC92+G9/rvmRau73nW9H8q
jDRVkWqZ1QH5cVmEXZR0YsW8nuYOUNqAjPRCNxh4Q68hXos6c0hwWo16WQ/eCxBP
fC3VPBAMQR/9Gc/8Ois75OPeI+Uk4kvikno2NkEQQSY7A49ZkRto6qSF/Bi0DP7Z
GiqExX7IOe+qMMXKViZW9a6+mmapTgQH2wEHKx4bObxU5VQgNED8WJO83c+ygQZQ
RLmJIoThpezl42GXuuT1+5H1oMlMXnDkDu2o5KKtw4x/eCI/bTxBstJBRBdYofPG
cCTCdbweF+wiX3Vwwca9KGGVhkwrzsiR80PE+Dqk0yuygtjOwl1aD3upsyOAfYJ+
/vWsMvoIzpOnvMARdWV118YFLhUf9HnBNgnz8880MKt0hll/PZBjQ320KH++l9+R
ypfBOkybJSjm/r9sATowSigYzASvY4UT3oMUfRhz0Ttdi2D48uF1s7BhOPTZ3z3j
wNu83aCPQ/Bp2Mn93kvUD41FkimCXR2wDzUh7wnfBPSziL3rzG0e3ueQlJfmChIu
YkO0NaFpLqfijFfYvchPBBFwX386P6LxLAKcxo/wJlt5RzyK1fe+/ZvTpvuKmlAo
/yiMCwmnXx2iuBXIuSOWv68YbrsFid+91H0tyOumaFW6FbmBqAFgIaeQsZ3r671h
fmiPMMHXZPlHNnPD6D+D6Z4NNfwC7f+8A2PAwAsIYrxaqZB9rTroCeXTzuJ7Tg7H
WY+FDdNkNmf+iDiucD1bsAsGzEJLB4RiPf2lDM2jKGKXGT1vTpX/wY5jHKmWeH/V
DiHKYah52OfZDvV3njePBVabNNW7odre2jT8ron5X1dWg5VxyvjYVL2f53FzOG5f
l8ptxzPsbUd1nJuVRue16uNx4jJ1EFPDmQ61t508GkPjvj3SIyNx1j/R4+Radn8/
uYNavvxRVOJBjkOAJAJl/s6dsF/mf4gLD/Lx3tyPqaMQZdPDwVNhTDn9IeMy8Z5d
60NzQEEP5ZBjnmMFZf+QQ6f14XMGl0E6myIOkihBPfwcR3t86t57N5HIkmwZKcol
3iDEJ3/LypLzsthBVR834R+BPjcmJz4eLaQdJs92cHuJuFunQPGZnR8a+xRfxWX0
4HCpnq1O/gbQA2re2xV26QkjhCzRhg/mixbSpmqHatFMt0Ou1J7LLwtlKU/X7IvN
y/t+mebL6VNnZhn0F3qiJLXYjDWHpAe6iTYAimkw9bAkOoRQg0jJcFNSr56vpgQg
/hoq6Jkvfx1UZr9SSmeLQglnE4BVXkkXI5v0q5OUFe1UzgqcrT+bTTeco2sFxJEg
jHmtgKHgxGEP7XxiHg3hIM2oK9UBbmtn4kGtPSVr/Drv1KcHAOw2y6VmtvA274YN
TJ/V+ynfe/1aapyTig/Nz0QC5gIZhuNbK0sYwP0R9bG48rSsmJfPm6c7hl/Zgsaj
I43tJ5ONqS5/c/lJPZBfo75g5Z9/3Q8TZFMoqtjJAarRRTPaOGQ6w9in3z5U7XnO
q2wqKH1ARrnOjL4fGgcY+CHU3vMWTwtnFDJYaRCC9ifb9Ha1XJ6bn89hhVP0t8kQ
peVBSOwABM2OlV4mgC535n9cJR8B0U80yiNf8tMbJUe1k8z1v92yzYnrrKO8Optu
CdU7IzuG2zINPO+Nmd0lzig7tEoAupRD/oOUkV8KGAT7nOBeKkfNjttfeMBQNSEK
lOWeIQI8tIhfvsalf7M15elK1JoIHX4i8MT647fVTsVQGW+os8yMBHBnVKDrz9j5
45aHeZjo8tekfwknKUkyPF8jL/TPX9Cuo6yBIFdAI01Sv+60fBTQ1dGkF58t9zDx
DzZYk9ntMH0MEVGjJ78h5x8e3vwkq8mP/tUbIVlOafwO3JaavHhzQz3gUOAYFson
ITaKfaySRe5I6fXCBfhIQF7xyhh4ML5P2ooUjYQ4swNoI+17bXW01gVwz2gXuFUS
Vva+PgIU8P6ehvrvSzGyekzI7KVzS7m2NAnuto+MhLgViXBuuJiNZsx8KhPdmguy
Gd1A3BsialaA0Cv4ev4S3wFGD4QJXfpDAgqoPwyFbavwnaWm2o8b2VGwZsTzNHQ1
zpxN5Jg9fGBQTB1lrZ640n334mXppSHgyEdT0fvbTQr6Wpg5aHwWbWvCh4mNtExA
BfDQ3ymcQeiaAsVL75Py6FiM4pklXM1n00eZvV26kQczp/XZYDVBHnA0I1MXAw6m
ncFggJmrvTe2KReMTm8Zp9ErqHvlaTyHsmFWfCzToGIqh9yjt72epxLIpsegbjdP
EQwLP4OkjFYgpgYF1L1dO3Q8IXaan3kebmZ7L/cOMqi6okKzZHS+ksYe2CUQYY4X
qakzKYVGkrn5LbGl7X02wKZGdz61AMaeNzLmW7YESYLkBeml1hI6HZtFFzT4cgzO
xufzJFUevs9l4TlyHr77btvZpaA6Bjl/biJvmfNyFZ2VOJYO51LW9RvN/Nr9Ymo9
PmJ1O0Y4xF1fXiF+F8doQPW2/rLGBnWx65KH89y868lMunH0iipaN+6kt/4dS8HB
iQeJxP7ii67VyuOdryR9qPpmgBmF2+lKGZqm8qXy3a1PSqKUWZDGUGJdvxhxvBEB
9yOhYVw9k/RYbJGS7/Lt4EQVyqBihs4pzTpzNAtwDMS+wDuvAE5JAeuGvL1p/lyW
CGxPB6/ngo+AhwLKxjYfQA26BwI5pS9iQG3A9IX1aaQvZq7OVr1+vT2zr1PFoK+S
Qw5g+u1ualn3O/flk6xk8Ua0+kK0/5UPU31wUhAZrdBnEOhsT1PrVJSb6tjgzsNP
c+dKguWuvfusyxIfiCKTDLinZp4OFeuviqRx0ka6//loTdVs4A2OFWF72PxEwnpE
Jl6sZFv4dUfe23LLidqjbk4hPd3vw8QM+Vq1mxmkOdNuM+QOI2trLLZXgQ7fNQHj
BiF7p2YC5cPsKRtjMEUrvdfPMiSz6QgSc2gPfrGnfNwKNBFbwbmawTmWNh8hPw9D
jrX/V4E+mpaRtm7614CyvOI43UEci30jVQ0b8P8Wac2xmVxfwSZf0lsKpR5NHLfQ
/muTmPIu/iMmb3NaPLJkoAPQCbD6uG85ZTAE1tOpnnu2vAJ+Hg0JZMItySiKEllJ
vP5vt9syYayix6lGWZd8o3BqSKAlvgy2PB9tkdNF1pNkBQtwcswHlVkvTUuPtGh/
SGuPFujor0PmY690ODc8avXMBIOyMLLpkRKhPH6/Q2w+zm9q5g7FY3dDL3Mw17Y1
WBhZF4kqWBHhN1PY/Wigu9GQgO2t54rpxRSEjxesjIWUUwjAkiX2FUDFiDn+aEZr
NI3YjwqC2KOg9D82aFD9AyJvBqtXfHlFsiUsEJFPBwyvGyuZQHfNEpiEFtAWXdd2
1olF1N58XQo4VwsNc3lwB/86GB6zTg3uCCCveSGVrKrht9n0nikuJM0ezBBRh0Yk
wUsHdyHv/idyH1C+fheEEL8aavOekhOmN4HXKTWP8n9f5Ltty/xynAef8NF5dFDm
K5mz9+f2i3l7epGamZqesMVAzHtCeIxhb8o9nthZkDtD8pkUp+4HDEVTEqv+d9lc
4MCx94KHbCGy9pYfprPGwe8uA2Typ0hxDzi6V4l7uRcoviOBVqPEfKFm0vIrHI1v
MNjYKbq8Nl9Fa9HwQEt9FcRWxIw/fQteJGiKRda1IxlH+Olx1vxuWpRAfo4D2wy8
97E+PHrOebZm1YLz8x0YQSmLspSzAOxNaKzPEBOPJ6N/4bOBfiDfK/gCQ0qhMno/
n78BCfk+QULOyFxfIgZ7ZLygmC4dLHrAYTpK3h1xqTSyZwd/jdaHs9J9XnnikaFz
2B1lPzrBNgWVCay+y6JqAx+SMeMpsK04Ic6XkatYomsNo1BObefP2aK1Qoeqxfik
ws9n/q3dZcerFLTrxBX0nn/MPh+I5RyUIxP4z03Cm+R7awKUIG2Lu7ZLS4dX9bnL
bQ4coOKGdSD062hmkoVtHQKn/N3/LsTWPvo4Y771bHEPaP4barvuNNOEvdxl9DEo
4yFTar833oxptFgA4ggDBMP9WbJVY/OK7rLIP/cR+UtubSDTOSC6Pib+FG/wbKnO
97ngdOHo12E9Pq5+/m4oEpDTTxof8prQBjEZa9U+LiNvSTbQUxF578qvlx47+GYG
Yo9LvOLCB5I24Dr0zLeq64QCGmeQ5bu4aVY6GcvsXQwCzmthVeRFOSHstLUNy89z
gDB6gxobz6a4wr1aifiWJe9N7oNefmxLgiLKe4oBahjKQ7yCYmIw98J6RMHgYUXU
Qnzf62HyQYFxM7wkLN8lsgj/DHwltvWZzinkIFGdjV+1IcrTRYb7NDjXIjySY/VD
n3vhzFG43DZdMUHMzSrnR8NxuYwvEcBmT8BKVQ+Rt7vl6mZwWA6+ZxOOeW+lylpU
vQhRWM0OZ1sHlI7VVyuwUTwssh06OP90OiyM7+KWQtqMIsZj0W1WrpURhuszSs0A
SCEkPd3TXrwfBRj9tXNBaNBTG3x2gGSX6bU3iiNr4FFLm2B6npQmo9+moplqL5jE
KDpP9JtSpkph9khwAwpGvqenZh4oye0xAzIDkqMnKjWQeiEmL+6RchTbzKhPrmhq
lWDOpSFYY5PbPKHlEOPrW4MNE6jmmt5+540+GDPbDBXxL1VKWNapTYfClxm8UiPH
xolPrUb5bXSlh/klbGkjBdu2CdrX6MWA6Bqc8zA9Og9iFe/X5g9CeT2QcT/emZSM
OEWYIX5cNeKm0eg7fRKRNe/NIc/GLi/c+BxiXoWQ92DbHkxkncb4/YvmHQC0ymvg
eNERlR6HRB8Azlcr+la9WtRm5x7biNfba/LuJeG9pylfdmkhsZobwfw3S65w4nI4
41ladAFKK3IrmotaKPUWc3FikM4zrintCIKmTRsbp3cu4C1FL9llXON/O3TtwkV0
KL3OS4gXEesd1pgW3p35xTv2g79NlsupU+CLT8uvu1AvS9f+emtDZPG3lEbZb0hn
bb64DyIsTN878drNTFfauiizDJsK4Xa0Ik+zRwhoqmjH/83fkwkBVd5eI9uN1hjS
67y2dyHuHETtsI4xgQGw4+41Cy+CiU2RUl530qbS7XGnmfQ3wfmH8TRW2o7pTxJa
ektrqNtY9UrJhsAA3GUXY8mAEYhm8VDfMD4c4Y7dBeWa8O2WPgdRYP6mF/vtziSF
c2dQdH2GS5ym9Az3kGhqgTtMUlUSSD7duFLDpXza2+LF76LZje0saEhj5KgNixDJ
KsEEuzxU5PTl2GX1orUqR1P9hn+6N7Pde2AqkK1pno7xvs0gG/2WRBdHK70m76Gr
T77u8qB8Sl+E+zSAOEwX16DbYFmPP9W8wZcexg9fIrpMrk5Ox/iS+rR7igXJd8tj
QOu/6xwwAy45UAghOwxrAFBJYWTcAQFlqhaSr7vID8qkQ5oW3KC6oRjNPe3IUppZ
cQSfw43bp4VtV1G2NTZMWlK39g/Wwf44Ypjq9rosGR3y420q45Z6b+GxWmER6vMF
rjDPZWyRH2aCOuuvHUmnsT9qhqmj5OHSDJ8yG2aDuseh0jR4JEjZvnS/YaKqdBcy
/UR7xIml4nO+7l/3gFqG6HsZQAUo70604l+s0u4+jW9jPYpaCkXveVRd3ntnnEfZ
+Sv2LE8HVfO5r9GaQ00ZF20VB3/rWByFRb9PhKJxYIpTHoHZ1ILlyKISPJZqXVEi
BA2GezczypWfBamX7aTW1fIMY4VYy89Mgjvvhjiy52Lhr3LICICW77ENdoj27v66
wXvy8qZr4Of+s+Ict0C8yenWzGvVtR+HHcBlQeqUK9QIiTVQfvsxWnO01pgWI44e
WzoQ0E1CMEDrK5q4yqEGYleCZU5clBUKASFw7HUyOKVB62aZLbbV2QrrRh8ai1Iz
6uI6jrGrvbHMuhy3wh4c6JLhQT2leRRjLee34tzHQ8Zmypbn7Hv8Uz4MyhEIVkm5
5cSnC5Ev8PbqCJiFyR8leWqNi8iUHBIZf/kwFgjqtlWfAf30SkEHHV1BpqDPvj5I
/37u2m+svM7pTKRVhHtRRmaXDXc0Oh4GzNvP6Qezn0xIrUASMP+tZNONZqluUQ0d
cq5Hz/mXcmpBz8YuQrXii0RXAxtpNYN9LgfaiCqfUvwp6XxKiQKpw4PDbNL0q8dr
FBQkow6t1S6B4DwssVtwxMwjV5z6hI4HtPUolNDWBAcUgOaACInQzZbeWGDf0lp4
ELZaw3kyHCz+qPoJyZMEnw8iCcT65oyKsBip9UFjiycXArZV9cbZtRf0aGWrcJgb
Ccn/7M7gBZDyO1WQoyZ56O4R65pMG4EeGWUkO8xEyRUyaztYDEM4F8Bap0YvVElr
LQnbHn3xaFGrIV5tzx3z/yAIH1qp4Pg4cQ+lItovzzaVVAdtR/K1CbDsvudLcFY5
CD7c4fazxh7WkQm5bJ1N3xLaDE3PPFLM3SatT68VbC/yVd2L8BeI4ZdwPde0aLVB
liGf36p4B0ZwSkxxy8qDPSHwXpuctTLQ/gvH83fmPDjRN3EIp3D6ua29iIQy1DPO
7BaYmGDkcKlxeUvzNPLxeI3Y1wUOl8vCD5v+UHdpRpmUX4C3JM0WM8YTUXJG49zb
g8nxnlYA0Hy1csrmaEUniDK+XMFZ6gtaAhTXiQ66DHrOxhNCe6MX71RiqEVmzneu
cwSE6lWVtjIK9S9FHR4AhrNDiYP06atHEKAZ4q4eqSbjA5nOS82EWOL/0UAUSbm/
E5e6U1+SdlJxy1MfE7z3QKGSY9P/UCD1PTfxf9ANtv8MtUXDA7kOm1y6CUarCGpg
ZCIPQ9YecgVn8XNx253N3koTHBvrMVgfmedvzNIGgN2hR2MmSJ4QDxK/d4lKLxSk
kFMi3YDd+rv0V68UoMP692BIbD+V5Rjk1+RU2+Y4N4HzED2FhhxLKw4yJkbLyOVX
2rXSfeOr84aK92A6eLeZTmbH5rKZxTA8eg+RHyRbylxvHI8zSEgXjI81MPvrKPki
AgT0Ym3YDc7D0XSNqSYXB02cQjFPhMLyCfmO7XiX2P13DaIDuJRn6DgZZc7psyUk
P7LWeYozqyeypTmKu/+wWse3av8FLV7x6sKVwMOARP7twpgCPNPnxvYGnpwFrIB7
srdZgy2q3Fvl0s40G2wKgB1+mUKgou2Qwig3l2UHChn1echdNkbS/qqSIU/tXRT5
yUnkNNTQuHlDLusOlqK8P/CEvRJ5/odfBHQhmD40fJbhGwSgqxXvUWc5BiYb2+jG
SF4/02S7iZy3H9mLVOxRy4rLqgYw8Q49S3Z+Fwzz4J5z/mGrOI63+/nLRoP35Ral
ZzPjVI86kivZaq5X1DVpMjpxmtfm4Hzt/9KIiWIG6lqyiNAznXigQEk4sTIWaj6L
U+U7HXNgGo4xvAcGA6ABvcxJeElgkcZzVOPKOWG4Gf/tC8qyYdoFy8+az/7l4DLc
TgKmFu+zyg9PPd0XPfN+d7y+/fVmIPlLJVprz/bsnGW3YQdGSy2rnj/AQhoW6xzR
O6oVMbVjcKwPa6qVGjkiKVxXpfGxZWCQ6wbOEY1s+VJzpuQX6o6zxM5aCvdHU6WQ
gZ5sPEJQOtL6tULAWhdnTVeVrUqhZap3Dg1x3dfWeNzdSkBGeBgWectgH2Rt34i5
pmEIZgXOFx6opDShJsWsWa58WQ7vxyp8Ii5AxgHm2WEuBLZWvPuEbGDy2v8U4gFu
T+/hiLIvo5j4qyhqu5IlFlrNA7laVVBu1tvEq9gg77TYXtc6OOFZCSE9mQs+C3FL
gni6tjqIG/Dmon3RpKAxPpmKdKkigvYlkBzPJWVeHNgJ2/+Zo42KpvW/Dl5i5OZ8
e67YJc08DG0n2lZpMNSccK8J0QHC7LYH79aYraq+CE9TCRThaSjF45c3pK7ukXvs
af03tJSNaqjdjnPTj0y0+6itXTFfyoLQ3hl5lI3bZf+d57GB37zbI5zjz/wRFryb
my1dmi/gtis+oqwFWKDGL5s3TzyuCJJsAuL914eKW3ShYANwyvCht3AZujEvfWk2
/AbSM9rvkO8trRfn83n6jMzYrckdQVBTVD4X8s5DXKeOPy76OC/+13QNmTtpMH0z
lzm6O4knV8CJzhF/lw3VgnxzCJf88O4Yc9QjwjjFZv74IC7Y+JHbfbxTqMIlwfvU
sy9H5giduLWmoB7WieehMmIa0J4i1PigKkfzVGyY6IAd4KYiXzFCZQ5pJB8Rfz1k
99y+RrIzW+xjxLClV7jmLq80mpzSMqhsiHPfVtkY4Qd+v9u+H0J0NFM9/GkwTcZx
wl3qdcy85LK1lSiBQjPbCjJJz4nI7EhBISqqJanjgcdpDfR36z1cLL/IaiilIYD8
q012rB+FyZWir+n6zq22tkeomxlNDIP2+jO22hf6894ixRLw7MpG9Y3IxGMw4g/k
vVncOnq3xMxofdfwLigdMVWgcWcKOQBdWRzOfbn6RXILPSV/6pXmElyh72MRrrWN
CYVGeU4iOleU1HeAxoEMZmUWxTkEGyzditXDsiyzBkf7gl+6HSy3NRz7J8JkcJe8
VuP2FNsqFw3yI14AK0M4xHrPgGuh5Xn/gPcdoL+cGWGxraBxDDTAjCi5huU5XOut
sxvLIPVBLXjsjeAVj/vZDZsU8qRmoYSLAlzn5ii4CKDYldxq0qcP8hALD11sUj7x
1fgfu5fvdLLCrkpLLs45uOcx684S099uE0m1bwpbD57FEg3PtVMQ+gGFbvFPFx1g
u2bRXUMwz67CJFPN0A93ViZ8jBKpSklKJ1cUUKe0slc0XyvK32lkEvbFgfZ0IEGE
BX48KNxDE6BQbv02SmwAxV6zafEmZuU4qIZa6tQ0iuhwmL73U/N5Z0zLQPnOcx8X
YiCggG9LUz5GEsWaon6Lz0HNITD9C+82IGehBJMH9xJXfx7XZaJHN4NY31hg/Ni9
VWYM8Y209zHmlEeu0CLWoZjbwnuvbK4JJZsLMwR3YbNsXQEljHiYm0jefXjf94TY
58gvAEwmBiHoNqo5eHI8baBMDzyqlhVLfcJJT7xMcjmlUGBDVyBgWG3SXTqzGJUv
B9fJpImwGiNQvLGJxfIVu+KBrhbXXuJNB1Kp1ET6/o8l8UWbb8b7mXaieQtqSKMS
8z6NX4RP+2e1GLb7206a4a7/OIDNRBZRSUrsZHhOmhZ9xxHBDMAbly3sLQO9xrI3
y35I7sdr5ytSVwUZ72veHbWHNwY29GNQWGcwNJnMkeoRzuoOwEejNqy5tZOjNuVU
wGsBp4iU32Aumv1NbBFlCoWXpT5IVCSrTXL6YQRUTxhC9jq8n3pCmFKCKhBT30tN
mo0+RFDnGyZO/E1ULD3L4VDv5aVUG68toZRStMreYnY/HsJ7trPseaWBplv3jIJH
QyCeTWIDX6J1Rdm7EaFB9Qctvyw+z1Yw4EnxQ/5II7dcjFWXq+srLzwTLJfAy/2T
crfG7UhMMCXGq79qiojOqPkaByrOqTFIFWYwZblgmwPk4MvjMdOLvNkc8i1mPw02
OprNCeSiCCkqhQSabVUZunkBu9QQJMh2y+PWvwPbAIpKUYEtJ4bbOj5KHR4CXZfq
WhhYYhSH9fL8/1tjmxloXOY08erv3ys1mw+plThZFjU5I9b+lGEGsR92gvNpF9Td
T/N9/Tf7MRVBzxnXOlZEJsHWX+f3EVkSkuUSqwwNWOThTAxDtkZDd6sHuOi8I8Yu
p8N7M4WyKAshbpJhOeFQ+KANzKa41ntzC0GvlhVaU+RRW2hvv5NjUUlfDI66dN6v
fywg3EOFaJCtlrPxb/48Z1xS5Kv3Je9qHkA8yABOOir0SUVKZ87GYgfbJwmFLIIZ
n4zwGshEvSP/BjoD2XeU8hLUHtUfSLb+9zcwMof8aAO8Hfz1pvpGT3rCN1Hl+/Nt
LpzYRZaCu1OHvGxwGcTHApNlGyxNx1MMY8Maw7pyvVmCwQBddiyvh4T1iCvmdn5m
C//itB26JnrXqeI3pwp+D2ld+QTFih0yKGTHmfKJ9Z3q5yMTMHnujx2Arhtyhx55
0XRwybuCgVhT0AbsS1f0w9JPz/OJTaQ5YzuKmwEMV+S/8xHw4qQle6mp9SijpV1+
E6oLYqs4Qrr70Iej+r6ys1B8DoE7Sv9b1IlhtF7DkzzHkKA1BIB/c6qRb3WRg/eL
LldUkK8w6P4rS/QMlSdAv3myxEYOfMqFtj4NDiceYdZT2O/KeFm6yXeF53ygcWCV
mJl2FJg7U0UjWdLh+4eqy2nr0/xtBmX3zBY1IH5ZqETYQN0rHgK4jZbCqsgAf/ZD
2isANzEr+AqzWtX28/57AmNbXtqkC79DNBvxnHLFyqECkr7CWBFWyeTrDwbpEIZr
my/vmiSU6m5m+kSThoipj8wD3p9xHxhIY4r8Xdy/aR4Th7cDSgE/MpKY4kXGMuA9
kuxzRNSbNQlxjwSS2i6UAkTj/sx2VB5slh3fw2b+OmEF1RSokwosOnFSA13cYBM4
TnbVNkyHl9YYeBSjekuQyPBj0N9xURrS+mvnwMlkH/gTc3eH5Ecz2s6IDYEf68Sx
Sh9AtVFXAQojKOmxXWUyE/3o3d1G4l2pJkPbyEMU6c/to+MjaO6DQvU6OkktCo0J
a00Hv6dUyTtVGqwSnu2TTQbNpIiJSzO3Zub9snBnuqL3Nxnny2459fn6zCLBVwFC
IpiN0FglV4pADX84nqUAx+MvedZPfJCwYHcR3Ve7QQ7UpIJ/Zun4tJKWb8MSA8Y/
VIPAydyian/BFArqamOa+jR1VaHTcF2+6JBpdUulrh4KfUKWwkryLXNrKcWrRtIs
T06jhHj86En5klWj4Z2NkUF1o4B3LYLJKykdexTvsqgm/xRU2dcxiggvm5IH+6GE
UuXzjyoKfqAUcQcv0nXjISyqxpN+qLZDppPEikJEXjVgl80CXV9d6dbB5gPhsfp3
3aoPgT8jYT8WIbYYTVsBKIICSculoCwmYxcukr7AeVDEhJmBOrPr4oDHWc0SPEZc
Bazq4R7deEJpt2uX46WiXanV6z9ZRSGVdDo1n7ckuqqe8l2Ux7lh2AdrMOq4BqaH
UH/xRp5SvKnXysW/3+KoOcClrCakN5UJf9DIuvX0oirEcoDNoV2D166Nrbj67Tij
SUZl1SZOzeAukFlHjHHfRKAif6SZlXHfh19wnVfSs5HcXzKoXHDtwiM21bjEVRAp
U53EwbS+3g1cTZy/Y3JsBn+jDsU/0r2Ky8EX/D4RhBqwfFJ9DRhAqqqgUWv8LzkF
XUi8/OqDAo+liY86PcHzhuFP9sRLG4KZIIFWd5fYxd94CkwCwO+94YV70MaduPXC
gebgWI1vsbyYDvzl34AXiEkbrFLCMWqapKHwFs8y2HbF2k0LilBCtKbDN3kxgTy0
+4Cpv8BrNsnoh6Cqxf5E5+3ixO/chSPDUACbWZevChW0wv2qYXkcEMRwlji2bRlx
C7e9Fkdshv/3lZp4K7coiQVNTomeT8rJHO8QOILXmLuiayaV/cvfFkQtJPLauwRy
jjBTtJWbjU98ivLAbSKhRrg/b7P9Ix4rOuPG9oVGzRT5qnjPKBSe5HAUJ/TQ8pvj
eQyzg3iLVysp01+PdOmsw1sOziG6x2dhwPMPgKKOCf9weOTbcDMuE2DQgRgfrlMV
a82fvhUfH61FBTKpw3CwfoLbNfstskUHP1KjQN9WmSv/vkf55JtTJTjrdLavynXz
4EXm6bl/NOJ/Jah0Vi5kBay2k7IfgasIECf2OEtoTsKu35h6stnRaAa1tKNG8/Mu
/QM30s/hEXv7dXmddb25EreQaY9Mxuy/JqB7ClmmdHKYlqR+RxVV192jPDKXhoZH
D/y+tkpSFL7N9b/6MLfxirX4oT6JPSrmFslsYx3cQyjFIXGrmbL/mh8HLGgfzJIP
5fzDmi044PEeUFESgVFQU53tzNlHHTCc4ywuid2f0ETPdUPTeeo134s9GlPMRqtn
LIiPk3QQ1eIk0GlNF2JXfXSIb0QJQD1JMT/IGnSbO7b6qbJMvFF2lbIjx2vGIacY
7snlpkWlmyvL/Zpu/kaq9YdnvMsyxHyQOnaQ305HFTrSu6uLc02CdzLveCQXMxBD
zSTU0DJaz5LQwv9WRrarP+rpiurfcVMTJvGgLMlpIyHQA2Ne+A4nJD+aCTP6Y9Xx
qBjzmdZO69u4SKT6dQ6vY8h7fYbc07Yj9nrGVODzoW4eGJXZEabnTTqECDjuzjyM
K9VBRXZB0W9hGkd5xHckRXFOWBqnaexLoyoNtObklzX07jiwydPIPKoPODSyVlbF
hX+G+tQtDzb+lVlaQOTQNnjs0wR15MKOzv/VRX6jEZAMjXmsX6Gz4Wbq5ktsZKa7
hvczZQoqedcQjAZWXj+pPK/qbhCCDuNxD9cFudWAkYdV8MUBzLj3HI+rTO2DGva7
IZl9WN6SIy2JFQ+pMXxbo+MtYaozkGUYhVQ5k1J3e8F4VQKelEr1upASN9My8hAd
dasDpp+FWrD4h1FnoQ+5rAU4uDGxCmqNjyT5/ZTnEgwtQ2WXTmHKoE65CM25kqmd
xIbbfHZzMDgXf4SCLUPdJMjoQF/bR0eaQf6+0lVHzqagA2bi19Ps7W7IuXaqOaSA
L/6gaAun5gQ2CenV/Gg9CxO/051Or5aRRINdt0JbB0wyC3NbK/ThqemSgUOgNOzZ
j0/4TvLxXp84ihDSvOrzc8PmsEp6RK1aLIL23fmE8ejAB9ANUZNJ+S2yCJT6NVHc
+6Bk+2QnSOIsHzJo5xFi6Qqo0k8+2i84AUT8mlAT2UIwMb3trGepg9q99RMqRRN4
7v2BRdafZc1X7wLzah3IzOWtRajRmdKe2hNQVshX/wzYq11niJDitmEIHbgoW7y8
oZmXzmKlCOob3J+4IEhUzn4Wpn5gkYoLIybHbHw1nL3GDwFBj3EdJHiC21Z/tVsK
JDEA19COerzTFU92DV5nwMIQtpLmY00l4f3s99BBcnCqZuHLGW6DJtnDXalTlE00
DbLiPI8fYkvg6lQjanec9w7hr90XEokVovwsupPsxAP+LIQKjeM9f/rjlEHtcvyY
rGwR/2H3Zkrk1UPTrfagc9WPxxqlbGDPrxIVuq7QzHLEFmT5wR5s8ah2ZmkXK5vT
aLhDBpw0Rl25VUw0azx6bjVhrgR6ZZoc6b6p3S07mVpSYR0RxSLv5TMIOBi/sUf1
MoXyrxImiq/PgVeyok0Zsqez9DnWIh7pHhOJaBU3EkqcecY7ULqa/muG+1Gs8smH
T+3b18Mbz/gIgvgGxpcM4vL5IWhsYhZV53b39VZjGFIoDdjIAjvurDTdDip6v6pA
7+e3lt3RtJ9LbUyT27LX6vK8+WSTktdYUeqS69P3yCergo7McaT3uOGUFi9G2c2E
8sc/STGu5C8asOIOBARB3CdLk83o1M0ssHsu7kcsWfgJC4QHwxADWpZloW76RAVN
iz9dM+iVggDbmJfq3dcI7HysmnrA/XnR0DCpPBlTBVjIBF5VeF1quXTa9yAPQ+Vh
moMl+zMJW48FqJwoDYKsdbUGO8KroIBxOX64cLsUG6lOH3ASphM7R7XyVcv+QiYR
ljxW/tWNnc4+D/CfDtH0X5/idgWF3JR8cwnMwF35vHvnhmOi03qFnFbpp/CWb3pL
OBfzGi06rda9lPzQ5pDgryhM9XGywQD/bFNsqxD8dDyOgWhDKZ2EppLV2KRK7wJ8
SvjkwyeDHC9u3qYnL7F8rvroZ9IV0vmboE3cXKM5q2sMUK2i19LTYiiuli1pg8E+
AYkEXf4yMJ75axHiDhP4kHNdSXM2SxKtVVyJxNknmoY9mrClOElkxVwZ8sqYdRuY
jTtUPfbaw64japovW56QWU4rHZ8vxtVD2vvZUiC/mFk329orLTjIWyap3+smngft
wiXGFjNR7oyJE6+IJungarheCz+p8i77isPFKLx8NV0NB+J98Jiz/szp1TYEFka2
uw+UKtbEUku9JKshE5z6oP86NEYaOOgKVpr6x/HaxjCF7/x2CmeiPGBCSycyHR1j
rRR2RgzTzeY/9IAAGugbiUpA8M84iGg3DbUBoTgz+xWsMipvqnVvmQn/kCycn0qM
TMKTT0lipcnzLdLoy2cGeTWFC4PgS9yK7mzi5JWN3i6lFlJTHX8icAowoPUhLvL1
p76jFEJjIWe+zi0HZWt13YOd+ET6/hhKEJTYQbF0X0mQ69dI8pzt1l/glKYZvCg0
v9ljStmXkwwd0MV1IMDtthuPa1UnXCkftD/yIrrE2oZ5XgRTlFKDggQHfPkpzHeq
oDbH3O1hKRSr3NGaDO1A3XQDQciSLY7dU/RE4OJEI3GivaTpUsNjrM/hdNfrkC8e
YfQj1ucF9AY1GcwRdlyNoqg0vcdQjSaTOZzuAQAs/MaBfG4VIEeP8dI+wq2U0pcg
20HwFgF645jb9Hk2V7Knr3dwMSKOG+bCHU1LrBBNTttsHAXqcA7Lz/M0pZHh33w/
WlkiTWM9FwVZzHnzcRywm/erfrL4LgRnzUX0vb2swu2DJqL0YfrRb12r8wfcJNp8
11AW3ThGrgqTYwk5ejQaaAwabZaMTx02TW2FFRlSmfVtMgNFuVzpIMwCHOJYlwOJ
koOF1VlzHSzhz4ZdOuKIb4csOkMSwhnxTj3U3b783RroWfkt5dXdSJjK3N5rqGmA
dBEbBuQ+5ypt2dxn/QwshSrCBJX2dwr4yQ62mQzOOUP9Ow+AipjRy/VLSlzMNHKg
/cSMS9SfG+GQcz8NwS4qwRqUBepBJFmjxVdFxHMd3IEZI9Gx3+aTdowWLN9f6V9s
TB8lqDUX2tpQEjefcakBPrnIy2YjKVUW0s5YhZOqg2Il7lp2YDms/SCJgaY1SChI
zsaoT7hrgfAFEEYNMDZVnYKhytEhr/jddguhhsE1rbC5U2eFY0NWorY+fD4cGh2d
H2bopCf/2CELuWESkLZVTf3KdQn0c7GNTZi5vq/Ql2AN1OSBlWOwAfR+GafgaM4g
OSguB/gVdCpjcbgL0Er6JNtdYr4Tjm+Be3pcepWzB8olNF2fMveO04DxkyNMe6aU
+0pVrhWoae2Tb+kf+9/HdrMvI0zSj64w9BTB5sFNGXKi9Dde5oG1L7l4fRIobHKp
kkLP0b9+AAS1lUvWPRyLj7+b8ERmBomeJOJFyYu1pQxzOT2IZJH4MQ+QqnyLTwe8
pcWd0cu2APeaKAsOP6flshDy7ghTEOw1Mgmp/UefkrCEgLqzHQSEF3gsDx18wrML
4+6L91ombzSXXVLf9GivpZwNbGNZhtpuGtWyiX5R/juLJFS4wD+1o2cn2bW9hTLE
XGnboCg1eFt9JjImWcuhEaIU/fKwplwwYEG6qtlqdCGGHZVsvmYS8Br0da6SbJET
u6Fmig9xTX4JFHPGOYw4zDYa0GaBmwo86T3DY2AnHVw01F7ZD23o42KFeviB87p6
FyYdmWU+6vlnEJTsiKCg8Lx3nZe0vxyTd4dCp2UsJlXLU4ybz5GXqAGRzRQQiSJw
c+tX6OvidRZeo6TugNkqwXz8BTa0ZetV3Fcb/kh0qVKO7SkZ+mkuaxhsYLxAkoD4
XNkh2A5IyaQUMxfmUiY+BLCzOKsd2k+wLMFirlsktYkGQfVtfTHYgyzPkrs+CHYi
oY8Wun8uEtB9z3xHHT3rJntpG1xtr1pEfrWIV7j2WYN/LjCHPcCb+FjK7+/d5b/c
bq9pd6MimHTvvh2iRxNTm/uAFnTSpW6eH1i3VTEiiAMEpuyrUKMTmAYCB8RkpYFC
q/2sZl1cKOLBn0x375yJx7/W4VJRQcC6ijBaAeP9+C8bK+cc/9gHiDpvjGiBFjiB
txPTQ1xCIPRCs+Ub2lAIV4b3CL00iuo8LQ7KEYbMWUivkWt1yEio5impV2n5aMdY
YDzm9zHOAkK5fA/VQ9JFigtYZCas0VBLhYjK2FvZneWLdATvURIAIdU/KtM3kz6p
D+uKL9OTHOUkcTpGi9AZizgwzvsBqImBLuhFgJ5A8/350km8lPZR7US1XWbu6FKz
T3+zme+u6uXYWR8ura9KihEOHsqvq2QRZyVZLSx1HxsflrFMgZi7CoRFluVdk9vQ
sRG6WwQaVqCEm5J9wuXoYK6XoEMc1KSBZJw4NKqgwJyr1YUZtr0KTIqmBaaA1nGX
Ma6gjtwnUSpA1gjJP54HrjNZpl9kDWqQTXs/zL89tNQHFhqezz1wdqgIKrz8ROCM
39w/+F0Xmiyskssup1KeOorXtKhHJOlmFqpYnD8k6nuU8TAfr3VXnnzki+1tg/l8
hzD99XUl49pcsVa2kV7wvDWb1eEEOTQZxgwQPYtuXfLu42R4AeAq2I1xR0BFm6CW
Y99ZDrx/96XPwZ1ZvEE3bwW1v2naXz/ga1v+Ewc9UCmsrI9HdB/gJ+BoZ505flKf
zaIeyhdIX1HHxCn01wGBRQvHIc9e24FLzG4D5p6YsyELQz+HcxfDH9f/whxR690F
pd6gu56p4PbAJDhs4/+MgfICbYMpjt3LnJ7SMPxpDBk0eekrE/f7hD1dmM+o9D1E
5Aio489/uoOoAazyo6hEfxQAAP3a/ZSib/YuMKyHJ8f4lPfqKXbjJgR4EpdOPEog
t3g2vca6WuAuMjtPYPCCieyPWV6gPKtZIDQT6dCx+t+bqJMu06g5j9x5TQJEPrbd
o5nfNKUjvUzrC/2GswEYJxXsaob93naQgAZIGwVHaoWSxXyEXwwtXv+2CZGvXUls
tp89OJNZHN9KdRBGmi6oFAapJFPcI4OAL5Q2Yd+Z3WToNyC2PdOc7gwwZ2mGCecB
LT5hydwbN6nxwzG9PoM3NK1VbXv760NlMfZ0g1pJg4fSnHJGyVyP8OP/rqo7FiX4
qevLpJE8wCl7107+0JBGuWJuLOqau/TY474ABUxhRXvGMBhF88Dc0Nq1QejfCytF
fdub8UEMaGxg5woKA6Ur/fsyC32XTbwIYoCciGOg1nfFNUkCnqRB3PITBVYCkqnF
0dUhl2TQADy9BUD3kq7Pv2ALRw9ib39H/+z2v3z/AViA7HIuiezZYFTL5rLcbxV7
26EpQjhPsb4aIhzOFQJMEEVKDQiD0ldO5rs9lStyBidfrQ89l1gktIMBIFoJE3ht
1c6MaCksQROBq6BCTxGdVUQbH8Ks8X9Z8CZ9UAxWQwZyaHaqOptVlLsktiAHuJXx
D2oEVpw7D4KlPxB9egQ6vBf/eOZngCZuYy+wcjJReMfkuTDujRMmSHYa0sa9EnQR
6n1dRYXP4Z+vlQypb83l42vhi7Rmygf53GPFDH/IfMbS1eN9La7dOm3fJT8IKgqV
vbgJV4XMZ6QQUvLWb+W+Vip4KMcoJFAcGgQNeKNKbV9nWlZ2MbtFt8i3gymHxHt+
ONO9qYDLG9QtLd7NMmDHelRDEpHOq3Wbcthv/hhjJ3M3PaNaM8aEsQb35wVzGTVo
6Lj4VbpBqVJBZ49yTYUY6lOsXwenLKTTOX6/8OI6JIB0VYjs4uVFasiHa6DXRyV3
LMHL2eUXKtzsSNVnPk5OaPrZoh1xn5EyLtBmYlQHfNEvTP7cwdlk3r5+34ifp5EK
cas4yAqTUB+Aecy73el7soRWVVt7KCMIWWstzZkdBtAzFyZzS2DMvzfgBf987ef/
xMxRlTz3ojBoKSTw8s1IWeO+JVdBMpNoZg0+vA0cgq4mJvaPKhDUHcPdJ/KPgZ1J
RQOr9ydqS1FZ4WTPOmRa0XisgXvdIs26IF7U1i+syE7ApnCKIJhLmsWTwa7mD7qU
6NzEQfRbRxC63NCF9hCE8sqS0c+H2cjrbd2ct5bF11wGH/AoG1hrK7ogMhE9G1gx
WT6N7cInNcpC3+TDDz5CG6Csr+1/sblHFrFj/6lxdopFeWy4x1McfqdtczlkYavJ
1Qfm4zHbI27c+715wVNXtVUnF467l2+TJzgk0im7QU3Xut70VakSXwS3RK/N3nWr
xsXrVTdWqouw3UKh5eCBt5q35XAP+THzp2v4NmkmlJUx0JUsZs1EzWBG1wvMRURM
fl6HlxyDb2NJVkL9sfox2+axCwfwXJaTOCLv+voNLZseXvHeeunAaMYaSw4jpgjg
wBOhM9LPAa24VQ69l5RWvNScMk2EEkTBpAMdLjf6xn9KBtNvGe0v2HVMPwOux7yZ
PUwNOHqsXtgirO29FC66YrMVslrq/yeasOUj/Pze3yzH+umfxjjNn76gB3OEsdMi
EJVK+vxCKLaNZizwPSnzcVBqvLojnj7Z4O/lyXGWtTNAGKugx/vlWB/42l4T7W1+
tmuM2CNEDqP4hI8gKmbXDYUQmOVrPSbmobJPPbH5HoBet/Jua2knpN0xggeKxtRn
ukzCFhUsUKBPGkpAzMD/WRMS5j+/I7sSWCPZwrTwOEOzeGJknNR5W/PPLbIz7jFT
qUDDpcLjjWpltcL1/3in4VCzVNye7xJsokGeozq0mrY4yitIhLSPJHz1CAWWEJQr
gdw+lxj70EPMW3Q/moIZ3Ts5Y6gwuX2HQ6MjHnaS2vsRQ+nu/rB4yiNbzvXfl/yl
eRAQ+uKKFk1qEoAyTJvc9iZMrXpk+5kv2hmwhQN7e5Q4iGW4CtklyxMFjYV1CGD/
EQbQ/MNYUlFbIeG189pxa6k+LFAmgYgZixR4tagQrsDUF2xnvJKftjxjtM4/h7vc
qPh8YdRpQbWVjd2FeZp+SfMvzz62W/pP7X1mZxdqZV3X/2GQ4pc8fJ6DpfOLysL9
35zAZIwzTB4PhhMmEIk0n4VxmQk+N7A1W2znteMi8ybWY8SUQcEtDRg+E1Rd+bvG
wthyNkfB5sPKnZU1kOw/VTv+L8SSRary5/rsVKKYCmuYy/CCGoG1+AR1aC/MixvS
IgfFFGV5QOyC3jw2iobdy7bDSf1z5Ww32+ZX6iEVpXMIZdlA8yHWEN/hp59iwStX
jbm13KC0SEWPLre5uZREuhC7AQVShZUDexlvokAIsJe7KwwRBCRJlgEoSSB5gJzu
foX9xLFeqRTYNRsFRSGAhmIwFkuNGEl3pXb9CMe59Efg2L6C/LFjPzqu/iOaBwzY
Gc/nK9DqLuPhc6ZHipxofaxurZeu7i8dpsBQI/EBiQuyYidpjVp46j1loD90bNVa
Tj06rTYy9gCxRDSKVFU0Y7k1/ZRw3Sv+zr+cetGWJCjkdH+RftZacjsQqdYDG7I8
1pz8Xomeb/CiSNvzqNmRwWMXw7MbkOZ3RA/inTMUw0wzYm5ssRge+oXejterpO38
u0vIp5L8d5xIYJgepq8/Fe5pNIlNOXqvTrP+AQAhrzfqjD/Gu+eukNrXyvhzxWi/
3KGph7M3/2/nDq/Fc/hIKK3hfzZaLZB4t9Y7BhYQY20vS45X1W5/6xtfF9HhU/L6
bFo7Zz8jwLMqHgTu0UgDAOswIyuuky40G5iRp0Jrfofc08l8KqwGgyWi+ycSG3lg
7yAaSKQo7DzJAwf5fq/PaVr0ndixYhQ0h0VywN+T1udnxqHYme2sA+6rXw8wHg3g
Sfrs948egFzcqrQLrW0FNAOp5QF1jzWYmDTsMZb9H/hUrNnK87LEy+VCTQb4mw0x
RRqhFwfRsOWzQ2YNvdhwj7OAeCCBmrM0N5mMVQqD9lWa3x2VsYOGMxEZ5SExSiTy
Myoko2lMGIA/BKVIqj9aqS8EET0JyHBIzuuID72P6/ikRC9aFx3kmuv2kP9quFfb
u8tgbc9nqGrxcY5r/wHHvuJ3N0gCQUckFCatF/70oVuVpERvJojKlyYajnW32LoH
uOdBtHAhZn4xTtHEjVNcCntRL17Nc/jrfsGJ6m1XMch3rjQgVvSlENlMXhUqhvgE
7my4oYGCUvs7JBQ1SLQs1ATq0xZNZKu6tdO9mDuG1Ytqcq2rvuPJZyHR804mkmhv
lsY/Dg99OfO+D2CL5pLg1hc+rYw3zO4Mu1ZhKpYOXEB6qx8j8u+FiLOlJ8ihkOfc
NWnPTTUveSfeQ1WNwJ0gJTVMqIX0S933oleaLCHFcEhM5XGQGKH26DVPWW5tpdsL
Jo/JoHx7e5DHqbIWiCDXTOetSbJTiRCMcwD8SiGFQRLQAZvK6hOSFPJVRFKYqe0i
a+cMzkcmWTUpwI/yQB8Qu9A39b2OOM2HxhNqIw04baPLwLUVrSHV5IpwFC0K8S0D
ssJTsESVluLl0WLqKLLVfPIaKZ7WEdHXBLXR5yHTLcHoTtQW3QKr6iEvjkn8dovF
x9eEcyMGADAkHuTxVC60WTR/iUbxVY87sBKtP52UlpBug2VLAAiKPYfdYHA/feYk
W8jHUKJzHOW+5XCLyhfki49U1hXkiL79vwkVj0YMOvXa2ayEjWmgz/bW4vJVnCQW
eoLu69SezZ/qBdq6amkYvnuG8zPqOtb9rdTQZCfoQF8hktvnursUIsuZEzNMo1L0
wSqfDRqRC+7mDuTKM1/MlsFlu6zG+h1WkXjPdViPQHTL4uuQj1wh7UsEx5xWwVgJ
ZXsj/GPyKlP+/NfpvwMzOgVHPNICKYDnvOnhmojQlTLtMX+pt8uKbUdB3o/yySvr
3rrXpJ8JIAbVHjJqO6TlNlzaTEsHCXJpWQp4NWRApkhrphcR9C+/Zm5clopZV2aG
Vbd7ZMqERcWZ/ovfOQLbkqWlpC3MUYtO4duTtAsG1dy1amlGPedVE/4v3nForopY
hEfgNFgy1GdQ1M5SS1J0KbJdXDORyp3yywX3c6oWAaT+Bn61KEdWbGrB6puGjDDj
a5k1wp5ut15W8FdWl8KyJ0Zl/HvphdcEHHZsCKWwU4nU2AAInaXcBObZvwed5T6x
pYxElIFSFEzLqHRQApzHWtG0gxnhp14IkncN1bMbqjO3EVTfGrPnejL4ZdGdxmUx
bdoZLYnassM1oARNkhIZnyR5mH9v7sQOzYRS9KkaBvi1Mcnmm0z5Q/8FLJug8wbU
c9k7Kn8BvZk8UrdgNNCDqwmEYuR7MO0A8oNMpWfG5d/2IVNAXTyTxVBJrH5ho3w3
O+UpLdw3rHQtmNtDV9teV1xS3EQKTQFUnFvtTI1fG6vHCRpo5inQsGrGQsXCPfvN
UXsKIWm0RgHnKsBYZzZu+Gs36qAItyxbC4aVgzMXZwQ+cZ6UC/qk13SnONGx5qBc
3ZUJAwGAefgozVibSD0HaxRYSfSG9kq4lh8FqwemxQnZwvxH7Hf/Xt4ZQbpkm/q4
ybPWiVqkj8Q+SxsLn4tXTGXuurGmovBIacmccwfxr3/Kt4t2rHfOjZ0ojm5LOLSG
cl95GGG4XzdXaDfPLENnKAwsUzVrj6XhjgBDG9b02he+6JWejhx7VfFKMdDKp/q3
nVvxKG863cC2Pa6P5OMLqARpGFITlFqE7hBGnEDICDTGYTbMDzcKcz6/RJk3fpIf
jHCYayLIZgiyzB8BMx0u+gd5p2b0rpcxHHk1HOgaVPs8IfnJzEet9Oz0fqPKijwA
Mc5oc7Qw+Td787+yKW4leLiQxfK+gUall2TU1BaERtOb0mO/vNYVFOQpwTlFZT3h
Dqa9nmUzSgKvLa1J4qxjD5pGdnfkgJFzoH4Tlx7YBcSFHFfZcXny5w6+Ote12PqD
ANotzpeDBEIGOCJWBbaw6g7Vik0A44z+Z1hLG54MPFks9zmiB297nPyj7RJTHkHS
Kijamp67RFJA2nHjRnHpOqqyEaNIoXfZP9Y1aWbxnLPt0E5VW3crsLw229Qiwo6F
YRTMvk7MSIWc4bm55BXPFdsY/vBDjSqZrIfYduXfYa9S4XXuKb7bUahUB1eJmB+v
S6ELBZrSxPVVCT8XlyKYVbn4O9tj0oXxvaAYLPKKief7ER1jhn4x6ZnSwP5xFgJq
ZjER37Th08BxA/FHfnfjNosYMOlc+esYdcFmtwC59cfs3fK6yIRaYOq+M6RAJjhd
gx561OnS7wjnroBb3rCm2GA4zXE7CoP6FPA6nx2Kpix3n33fH5F9tUuKsmcPWugV
9xxJXt2y4UF/ExHpBLQk5yXGZZUa+W7DDd915O/HZPMmgfizPu9DbPbiTuW+VSMl
qFQG7fHAcKj5HxsVxfyUkjsgJFqt34fBOfm2jaipZkhk6J40kh8tMuQkAUIgsCL3
WK8H30RoRy5gDinDQi0z7iE8z1ppK0AEyI2pUmfxo5+zvB39OPpQ6mOdV2loaIfb
lXKm1rpbvF2tT+Y0vdJf0IbmSQs9itKk9UnzZXihkMbNLwcSDwHL7iAN0wU/zU28
cAX07GoCSc1IiDMV2KR5uYg1gGj4qkw86zv39gkhzN3dHb9u4wrQGZ1qpox3hoCl
qtZPhyZuXUms3H1J4+UjtEf5l5r8e890CqjIyeSuqcCQs7L7baKNU/l6ia8GY8HX
Dvn4m5okIq8N8it/A+Ok4bZ5eszRgDBrdEdvfdzYU1MmAnzrj8FsN/kWVH9bqenT
S9eiSi4rSpYA6Fyrq9xxKxMdy16Xe6N9fHhYmleTMu3xc1PjRoTdcBdsxSxweYo+
RVfN4cAl95N1BTf05fWulee2AqHSPYPsH5wnfJfIpopedYU4qKvBK1RMtuG4PVDx
cU9dOnmC4XwzOVc4niWD+hMAIg0wFlRiTmdTpqPEok6VXkKjcjvB7I/HMkt6+mSw
PBVggPGkjz4n3sW+LV1yrNyQyqTzZnqRpOtkI0WaPIBgWlgayTSCdsrfwrflwo4K
FPFaM5FuE3bpoelKFIm1cgmooQ/m5UKSInB/erQ4txgpRusDt/oBQ9Dkzl3uMFeu
fieThiLnm03NLGoNqzVj3y079r0NJVmWIzxCLyhDCq10nnk2Ojy3Qxjv8+HCu/oL
Z0JigazDpDyUEeeR5xfr07i8wMqUquWHzBEvhmEHuoRmDAzXoMQuKi5feYyYxxV8
zalS4YnCweo2JMCH/SCkB/GGynHDNp4KHVkCnC/ZNnM5SRtaR0bl8XJO9o7hxw5G
WxxEtXrhyrSdIrVQiR0UA2jR+dC7/4Ys9Zia0+NnfjTRLDqn1g/PvrSMync7r7Tp
gJyzieCYDEnQvIa/CJ8UC9ewSuE3C50s9tCVqc1ARAA+bWZtaR9sMfoqI6LId0mb
lJC3eZuERyuXUWiAr9A09XUnuGCAIjvBNVNqiENQEYkb6KuHLMHLqSpHEWpkfN7U
nlSEyu6dwtqxxLVh4fEk9UoeO5a7HhCF6ay0I2wPw7I7rizf+XsOUJ2N7Bx7hYb5
k25f0IcZLYAN/Sco+ECLl99E1yhxZ74a8BL7Ksk91uRSG3kSJayutSN9Rrcf4j5V
7eWSo+HBdng31omTLqbh/0WPMnRnseIgZ2ldKjmaf6XGdEy+S+oemMtXDKX/XXi2
K/ejqyJiKSdO2NngTa+CDYzt+Q3g67Pr1elf5etry/wFxnX1hKip7Z4sgabDEhph
WmPqgfD2c5EZTW83sTH4PD4cDDaLuUqCFjhAxNo7Eo9qPidbwdPSf0U6EEakVQag
IkHbCvK7OdFkpJ+yGKp4dCchd7W5/v+OkYwID5MFrLpRdPVmS/ap1SoFgH2oiCGu
oDqFnL4CODoXkdiYc93Nx7F7Hmr/Z6BwMSL6MF8rOjvgtIosFUKPWL1HPjhVtPnP
Fp8W7npxCQI0HmT7DYEMiu7tJGO89qkV/+XBH3TvfHEi+A8uZMQ7Nkspyz94MAFA
aDS9DmHctIgBiNBsX+V3YRjdBQCajzVxQQA2DNl6pVYMFa9SK91ifq9PqH8NSAhI
Pp4SdIOb8rvjYC118OXVWPRixE+RscqRTOgCariWJddQIIAdzsOK5IlXH6eQbNFQ
+AH/dPNMEriRt4xylzJ+PL1G/uR9/AKCVxA8qAHGIOEfOQnn1kGTTpAYwbv96T+W
JrnFfvYR5h5p3yxmQKFI5DgM6CAph1NWjf4QlfC0Q5vAISJbYDKD1Nd7QEuD69Jp
4+jSoZcQT5oNpVwWaGysyTr1ZWEIlxI2dULV9HASiRnfn1O0Q7kPf1maPjfyO/1J
9G0wYZuw6tRjHOvBhJXylETbTMIt+4V/CLftcMszvA64bnv/nHbfUAB6icJUKoDH
H4EOiBYa+Ih0k3vXlJIIIDtoC7Qn04WDnBYU3dAMJBYbll5xIspkKr42swi2MQBF
ZjckbsSDg/y5vBKXXrEAwfrVtVBgM0neUXaObYn9PinOz2ZCI8QJwUiA3Yw8/Jbm
d4158o3vLHlx7O6K9eekJrUZl2hYqQcU+uonaAdtJaKDzY9SQyQPigJhjLgsZL7G
UU/f7hQjo8Xl3/zoW/KTNA9DtA+v+eYzTI1FHlHGTQF4aPMMoivTS7XFT0Mt0Qdr
0Ii82QOr7GoOstyyEigglyCmWuCEIq8oWZQOrtJpJhjxDAYq6Hq3cpWncXjNSY2j
xsmwCJbqh61qS7hZHB3jhCAWyq9UFjoqaOBQQ/Z6cUezVlkGCw99Zw9g3Z+8D8iH
kBdBz5ItjjW9V4t/jSba9rz9SBE4szGz08ipfgzwCVqjJrZRyLXcfVZRuTCgUmvr
JrwkW39GVlCBBN9CwKsyqXijTR9S1NhZzGMU+K5F1EG6Tszbmbyp0AZGgWv5Dzzv
rrmaIUg6EHyDOYS2CluHJixLERjYdAE2ORYEGTnUyPBFE7SGN+o2HetG7xqdZej0
miNvYlRlCYkJMAedjFs1J6cdMZHOuFHjnvzodne3wEe2eTII0DyU52cxoBJNF14R
Zv6LCvLvqRKyu3MTzXsIh+RRAo1BAwhdyTLAGVH1mpj5sjuRBuAyRE1T2vAOLFpx
cfnalNAdCoffh3pkLU2lva7c6TGAbgh2YAZTGI+mvkGQ2ud0hJ/58uJDkpJsfdTD
gwJsp4xrCB0JAPBauA0wCsCIuUod7N2BP2fk6LnAVeoDsTyGCoz0NoJXqsmj/LlE
/RKGBVCewk0qsxpzGY3VdWp65yME9AEZ4mzor7WW/WaSE9GKcPe6OZupuAfsAQ7E
3AtYN00ZlcoEw2uz+kCl3fPgQTuVmH0u//wAVVFQenB96C6yGknpzn408xhP35gP
yEfhKDN2tWOQnl3J1G6ZHsDot58m8ZP8HPNHSJKMQsZdDhIOpziWrfM7k63Qdm3z
pPs5Q3i4ao1Ccuycp2cOpFY1kuTSadR4WOWB9+oTgCq2XwUWAKTvvobILUkw/Y2n
qF2SI7O2+SdFNf6bIyhQ0dV7wNn5eEBy5VAwl+Yue0q2wNSfb31zvDLIbk8ZE0pI
a2unNAdQV/P45HyfTUSESPnR8wS9PUNGmi1xRbBrQsn+pfk/tRzsW7ja0ttiNN+F
xT9TCOnPD8IQJ/DXQvwyShDP0hBvLkn+lSf4yub/EVUFEBM+BrcPlnJH5huQglW2
6+Un7XABuEtmPiRqYmb8ukKYP8/mQ/a523iFaKI87ufqFkkRoCv2HXLDVnoHHelR
m0/yj4Eypv7xhUgp3KPul/KDqqU/GyW6RS1VCgOLA6fRKK4W6ASdOoO4n1BWQpOV
6p6e9Ak/ky4RpYVBzDCGAyCRE/EEMqF/hM24tu/svFj89vmYKboS/iThUQWHPyAN
g9MPpH/E7ZG4SOhPlRg8ZyTUEoLWF3k4e5AYwhIEqisSf/HMSpjT74p0L7UnXTQT
pc6smJuMhU/zx2aePaqlyhlYo1oBk+A4UUceYBwWQIptzYuZQ8M0auYuOyNmjqfv
sl1pzguHmYqMgWd5X9nAWt+D8JZ/QUfGcfP4ODxZazOSuxtWBIIQHo3GJ8H0hZ5V
hGnCe963+SWj8WWk5dy4U5dGeu8Fxv5PZEnE3zjhSkPP7P/8po/nGRD0tZ2q4cMw
wTG6B6akouSU4XAkkIa6XQ6nqA5tX2FBpsstiWn0GuxYUOqdpyYAQEKjj4KsOaEf
8AZVk/oU+dGTamjqBhn9OspHXj1oTiSCzLc3cDb0cJ/kx/o4Ye2O6vdL9OOL1m+M
gQ1kNFBJLfXhGvXJTpg7nOjbLEaR8CDLId8R5WyiMCRZvHkv89oNyLRddKSq3iqT
xWeAtcwQuwYdCDXDY27n0hSy3vynyyg+On+pTBj/ADBw62Bn4qAYF/OAAygugBs3
Hyyjcvo0yZndriO+ihaEFX/9oPxpaLo4dw9nebZsRu7f9wnZNVsPjFwtnKmIR12n
5y5iLgvaszkE0Sw33ENLyUta86qkM6R2f3Wopv9UBBZURzvZMl/uNwohuB7YV8WZ
hhDbQKRX0YqMQFGqLsZoJTRqck5sXfo3eQU1xS49MICjBVPbuW5nML0arnilcqGH
bHDrL2SoSH9YKZtM6ssBHDzHmKw8soj56YdXm6p8bAWolFPw1qvqvwB08nFIjhUn
mmwrG3e/edXqbz6W0dL5ELL+d/EFx+y2PFuIy3JZSuucPS/6ypd1U6CqjvKXM6WZ
g1kf9usyoA0NooxyjRtYMiXta/XZfcRhCdMUbBq3Kko9cFvh9rQK6/GT/RQCHZRp
NFkQ5C0GJ+81mDrVjwvhh7gwQtGzZqc5TKMJo/tss9CmMq4If4ArzF6YvnNebuve
F6WYH9tNnCzi5KhC6hKXHpotBFFZRdTOwUnn54IjNEecFDUTSr9rdfjyR7Zxsaqw
PFF4R+/ZgObQEO4sOKe+yxxaZADxDMGVaINTCYrlzsj0fM+xdzCZjo0CszUl1sRu
cRWZq7ZN/o6XwNsGq/M5uxm8NEl51qRri4teaRb5onU9hEVnrxCmA6HSWLYGMrTZ
+J/ynzuS2GNQpjnMqi2ifDU8qGyb2IFG872MOvxnfrSlohFSjA/G0jJdBNn2qCdL
q6OghsDYAnSkU60I1hK6hkWS79FEW9jmPwurEmqv8awy0AFqMxVeTQLrIVOUIkVv
DjFMuiAuhtxrVHd0PLKzarcnKERZA104eIYmbu3GET5PJ90KmSNjfqClwlWzpBUf
ellSNNVeGUK1JeHmO0wTZ8FucKJLZm215JLC4tCogVPv+w4C00sr268jYIQq1Eak
I9NJD5uABRb1/5GktLL/2gzywLOWDuk/HhL+CpHdeder1Z9mb6NgeEHQslibNk0b
nl2oC3mDdzFxrR7aBGnZhkLecm3iZ//hrspt5BJsmxe13+/V2vGf2b6+ZD7f+GST
40o2hw6lX7NGces5XUrSeELxHXxnR8uNHBc9AZeMphvR3PPcebITq7QUdaAssISC
UFuOnyKLmrUbC2GzB9fx7teoD4/KUeDVSrRZu+SMr6xKUSq6FFwWWaJyaLaHZ0Ig
+fc4Cljx0ni7Pc9AKT1vyrZ2fuk9vmDGkF29GKYOUVWfSv1tOkzLbdAo7SD1cuud
zfwcKPciBaGHPzTxfA87yBdOCRMDr1BVYTfwHe62OLxGaEqURKoe7WNMEPjxcwEM
RjqQDTPFF4YMtosTDJ2atEiPVXOn9UcDSTkhripF74ZcefnyE0XbU/fvQwTJIeS8
NEhlmIyVFw3OEYAu1zutAcitNERCqNdcVonpRv7NV+lz04eaId6XFLLo5RuLPY2i
gFCKgMMAqVg6usOr7cH8PcltKlneHiaxLI/WwceDJvms5Qumgq/YCJG5rkxVz87+
m5f9IOAqIkGUctKvfDQRM5hU8/GQ+bGYf0/rYRNCMPRNdJG6bkgzdlLC7+4C5ycF
/Ge11ztqC+4S85Ccm6S5Z78g+8KKtnJWVnF7JHplHsO+D4g3Q87A8+/5LS4veCg0
EuS3YxL44YhCgbqfVV4CfYYdBKkTdXSTYrdAwoTY898dhZbAaAOVD225dVyEC893
uqlbtgpa5CHNvRAw6hHuMI3Is901ADcyzZAC63A6J+27nq58bpiAm7eqveGBIIaT
4Gn08nruzVdMkJyWVks1VhQNygSchy7avWGel6hCUp7g+N+aYI8QSGV7aC8R/CBO
ZfqVwiGP34Ppa9GkhbrlG80NoQ34hplfP8tn8ujuR4J30Klmv6iKFKC4grcnQ5Gu
2MqTv1MEB/nc/Z2I8cuNBPD+kbmfmjL9KB3wNmrAFSMneEANuZpKm7dUMj4rYHdf
DtUbpAxGPhlixiQV5k8hmm37+2OGILQkpM8QPfngyRiWPATVqg7+T+JuhzUfS5Sl
xjcssDNdZdHITDrqZxoQr4/Cj7OBeJ/H91TM1hZ1s4PSjNND1iskPvh+LkVlSZp4
EyC0ndcXS9OjwJSd/b2PsJ2oslEBtdGIfKM3R8TjLMb6D1RsvwekveXrDOvuChnW
F0194jh8zKb20LYxJK/0tw9N5pylXt3gHCM3E0W9UndyJUCyAaPCFMuxO6aNG04p
1wMDKmeVRInU7CSAjGdnYCsNosnzuGc2Hgk8MGQ1kQ8OioVUB0XIjyFIcFmpNAaA
jAU1gK/yNSMqMl8Ewn4HHf9Di4WmJfaTRRcW4jZjQgAtYwCSNE1TkiEiRSrIrwyI
jEr/EPOOuVRclRFtOQBdQW8JL9PYGCmCIUFH7Pqs03sXk3XLYnQ1HPNeAVplQjDS
hDuXYaLZJwwttkx/fr8rQfPXcPgU4u+tKNZ9wFLePnGThdwzcgg0hMNIxKNFAg35
z/UXsHe9Nb/y3HHtMZvUhHU9mvQgowlRGUyloE3Ji4Scigkw5rGCCSsrQ1TtnNx8
q8uAgyZZDcWQJoK/9sQnTt9OL17uQznhU+oCV7U5VvHjFH93Vf94VxGRRmQkVmkt
+fz6e5COgY8X/bC1Rw0Q3rlsYmnzZ6srjJnvHQz/xs+tFrX8Y+fusWvXv570dzhy
aJf+ZF2VdXZw7kaspeGx20A8hxnLnWa+EzCR6KU7SQMmkd8WQDKPRTAMUBQlgrlt
BkoKS1sCBu17PcJbCfP7k/iq41ZZlPjKTczSmVgVUKwIahNSE5+F4Pcdri/tZM65
V1eEKFVXYHv+/PK+oVpBtpK6DJbN3ZHALCcSYxZtHOS8Zdl2G+oNGH3xxWqyhCAt
k5ICa/k5ve6PNLiRtNuZBnW1h2JwEzKOmGENxlk6Me9DrBVgT/sg057nnlDigHL4
u5vkbWJk+2MH8/E/cVQlFDW/MU7EVefWTZRXZ01SYPDvRB380bP3q7pFonrn9HQy
I4QX/OWGCJETRICUNdS2zosDNqSHjFZFvOWVOQrsOt8Vxe3S3XABwGrtXL2FJ0sv
TnQp96925Uv1D6Hp/42G4UCMScGE2Gmx43hOZh+SYT7gtTQVLoos4Osj4ssDgIU+
7eqsPFQUDrzLRkdOGPPWKiJWzHKa8S/wgnLGdwf/d1wF+SAbXTNbuJ2rog3MzlkU
n/Ws7G0jjBp4DRzK4lqvMmUFzwGb01uWzkPatkEmw1rL9it0Ha83dqL2d/UU4H70
m19NKkYlzwmXK73ZMq1cKx6B42Zm0JyPSFE+XBPfwDjq+IFIBogELZ9Zng4wzi9S
BGYs9cUIWOmDPf5DODfKaX/3zCemvmJ6YSvDQV/ChX4Vpbn23fl/J23T6rdGBKgp
NJvIbWDT/WJ7wuwMz/0Gu9dJdtdqvBiSt5Sg4hoAW47vH5NZsQ0qmwGYsnHhd1N5
ZxAzg+XMZfpCthiugG0tSk6dCb97UXv5nYcYG200MPxO336oyG4xDzsCQ0WCT6m0
AqLHxyM8iLtMIVtPtkNAUK9ieeWPXwVEWloBcslCHPkL2Ul7ntNt3pjr7TeBaJ+l
LfkwnlpFJ8sm3dHjMy1UwEbHX6UL9qT0jpWIDTwg0GRRPSACZnlk0YDXoJi1bNPa
PuR2OVpLrwt+r+tSrypK2ulxUVTK/F5odjwjUCtTzgt6S120c7aHwYL0GzWW4MaL
ZQCWCaYsIC2N/UC4FCq1zJb3k5J5eb92IvIBGVmbE+weDCy36dGDycBKGwmQoVJI
6cHOA/MivrfcyeD2ZUq0xAYE+5rHtmCdTAvyacbSbTkCJdpWWhrPe25B1nPscb00
wFd/1gLkZpqGs6LrbMIKsj3YKmOTmJAYLf4toFWf3Uy9WgreYikQCC3E997T5DZP
D/ARE9ujCJzhG3iOsZpBSJL8TrDo8dUVQKCKz3z6IoX9t++VZagBsI/ZebzkpbXf
U282Rgajl6TmqeEiTczeto7fxDVkP6tUgM5W+8l3wQaDHoBuCj96CGFhTSck4zMt
gmZ7pvGzL3ErZC//Wi+6ykhM3ViZZxAqxyXv62dNCFQU+0UW4Xq4OyC3TvuwPLC/
CtAyZQB4eLKLB43pCBV/xZz012d4+x8BPlX7zgWa3sTkGSPxfeVM58v6hfrhhS/r
kreH83GK1LhO/W2VQn0ZsjWVeijeaFbBV1BS/qDI7lMsTmRm65ICsH1CMkWVw30+
8PDwRPHuHt+2pdSy8lBfTSuTvKlPc73jjarDipGEm8nvES4Lj14uJsYTZs4eBT79
jswBAcUWhAvunexQYiAWWvorG7edz6C5U+0emd6YVC/wafs8okquxiswwJl/eQ4x
YI8gtBiLz+6QQeHd59hN70F4RQrCf8xKitKwZgs/C1e6NPJ1UITe7wVCmq4hlgBW
OA3qARSJ8hALgKkRhTnc1Z2V4NEE4nV2IotQUCcaSb+U2peINuiqcPv4QfWUtEqf
CtfRGsQtgRBCN+vtQZ5DrLdFepZ2vSTUaLb5Cnny3UwbgNfzhR6CsuioeGZQ8eTO
l7bywAyOkFcwk5matg1CuJWostegZYFw2bGFbXhusX7WJ5muGWcOLav/pHfDK8ad
1dM8tJxes3r17XHj2J9qjOGvYHKtXl7Ze00ShGLqx4qYqbG+mu7ZuKkwQGBghj+N
ABJr9/f+9kGGnnO0PFFieydNe/ClUw4N+zxINegzASzQykh4zOlCkBZHIrHzjZ6p
2E2Zrl+PIrl75M5paeJf7tvFVJNtcS/rrCwKYBNLTaoVL5mHoh5xHPP5AoRJ1gEY
1nlPTHhGMPBrHj9Z53EhZS5VeQOjKhyEfIwwofee1klrMkCUmHuegvlFYd+wk/7B
zqa1HxBXSz3odqEna7ECpiHoT8aXTm0Ya3i/hseDRcYOZR9JIMU/IMkAIAKBCO1Q
kSn0oVqFamDFpH4doy0YU1ODFT3H8yayWKZZ9PKGdszMmVrh0fW7g0S7+iGll9zQ
Q37GDn6s5GkT8wqIoyY1hr7XpNYQ/lTriFgbe2dlQwBTlZmCo/KeRWsmHivb98gd
CU4LQ8tpJ/jufTpZ+o4yqc2UGsWtgyY9k/Y6PhAt1BJKKfHTmRN8jCK27t4tU91e
d8PYHr8jJgjTUx7gisluDZXGbHnaKh1kBclAlrRmZVdUQJsv7+pwlJd8kL5kmitR
3hGbVA+OXB0JcSnRxJGfyt55uqUywwaTQljbZVF+Qle24XdWzy0julP/wxKf2//L
ZGcwqRtNOEyNCsvc/TWZn2TrVuZUp/tqlFhpbCpFPo8RJM4wHAhib8cxNJnbrjxN
JQCNf3NT+26D46O2fMSBmwLbUfolxmnik8P7gHUCoMcDSue7ZNkuCQ0pUw3lnvD/
vbQFMjWLrQoYxfyBYgkgvFbOZAma/l2ha0ioKkNL47SXsObi3hpA6g+1JUz8nVVU
vwtvxPpbbn3w+wkXWf1iiS+OpyZGCgx+2VgPIm6anih30kPlKH2pX6aRJAZf2BBX
hnRiDbz68yQOVrrS0+Z9Ybw8rt1fNzFK/L1zLaYDrJZhjVVFBoFG4uOwEytw2rv6
BcgBAYtfV45pn5b77Nkyoc33/sU9/FQY7GksZa0hl72d4+ixOsI+LwGSYPb3kYx3
KCaWD89PqALIH43jlT9YTKFtgCAHJ7H/4DeKYziLFu6TzS9Ye4ckMldeLmBgej4y
vENShYb9sv/OHbTmZ/DA09v9sHw+/qykGyyF9kn7JZGjSHUyuFVHXQ0gMdyK7WxE
SbmtwJcf9u9TvLZOjntXGi7eWxPt/PLk/3bamJreufQxBUskBqF+Ld3UgrnKCgli
HgIjAKZo/EXLip7ZeVyMzJ3/hzS8ItWJ6gT0bW6qI+R3Gw7UxdxHTEInsEP9vT2p
RGUIMDo3xCtvGrRO1JCLlly/AVukZBAd90mQobM6McCcpg2TmtaZUvhH5NsKz4b3
xU29lmTW3mf9A8JZJ5kujPR0pgezi6kffvmvNDvSAy14l6Y/67tqtBDH7tXmolKH
Nvm5vE2RddU1d4L6/EHDIVgSEuJYErOLMNUp+aC5koJEq7unpGANhpJu803QwEvQ
PAnDu488mEQHY8NquccLsgnf/Z/1+ddby/kh3ZmIEtN0LXKT61hVlFMCy9F827u1
S9tpDDmJCDPV3QUoAt3T1+FsPhuAPryBlpXHS7SBHGnoWWHFP16apUpM/r7A0ANK
X1ZWb+9sj/2W5mCueMWYxADo1qVr+vF2Ehx+EogI03HlCXeviSDuS9Kj8xpjx4UB
Hx1dA3/PuOnD4XWFX9l1eqoiDBvSWVXT5lkndYB0G+Xfp32DkFz3C01Dbq+o8gIH
r0puNS3bgnVQM4siI9K4VFCKcshfPSYVmQIlpNSzJROTNCLl6Ymlbpy008p3/Pic
Bvkj+fVm7fBOo8eMVYooUuca7vplfIX9RmJ1EtTomnT4h/0CPgCyik4ML4RqWSC/
yqyW5406C0HwigWgafxiS1DKTdFazIjMFaWrsBLu5S2b3/gRwMcZ3wrxDBN/7oyy
7ZBqRAMZrdexT5Zh4kfUXYEn7AKsNioHXoJMtWRTRfNd79/mUGwxQSgSZs+qULtF
tt6IXT8Xsv8OXAkMWDNjerpHIXk+9kJkr45xC/4dhuEc0dt7XGGPCROEHZPodXMp
/0nCkK0O7GQ0L9wQ70He4bhPeEAMqgQPHP07kIDwPQ3lIdqrb75pzIzvk084LNbG
gmp/XrZSDS24vHOLKTYeHb7Ig7/H1aZTuzws7aR7pTkVUXnXRv3dW2k3faSdHGlD
e51cCFAG01I7Tl6mto2/GwXK0is5GlmUEQkCrhEozRppUFtskBb1dFpxxb4Td17Z
FDkgjn1lfnpRoBc5SeLBX44ne4BRfSxmq8QOazS17+W2o3uE7hIJmFmWhfHkm4p2
q6VQp6EpYDALiFtjUBwtNC+h3HPpgj9ApOp3eacj00PZZG6gnm7o0NWLKhxE3Ey1
bzudQUtU1DcHdnTpUfgTBH7fssYiIrRl34XNj5Ol1b3BJ2uZ1kVK4MWZx0SBBKVY
r4pEHCrkl/yrQwdkWMsbJk3jBN0rttXMkWTKjFANoEilIm1eF0ogwssOo2B2oMaN
upt9yGTEQj+31hxQGyvgeJGVsk0p9mLR9KczjKzmNKMUUZ1sKrqIK2tkmxXOQihF
WuzI+F1AMiyXO69vGaMML6jP4RWHT7vYgWyk43ClEm+5J+fV7gBmRG/Y6ngt/aSD
qlZSzMptMFDLyaI5GHwxA0Suw5VkEXQUWa+wnM8STHvC6x1Aq2ijropZHZvMwUrV
0GkGAf2aiIDbkO/VN4LixV3XXirCwpJKg7nJJER5/1aQSjEjru5h64RhUL689jrt
9NdtV3in1wENFSZveHaRw/c5rlfuAWwKFW2B5Nr5t8Hq3RCMdGmPb5+eq92dn7/9
wROh43HYuNZgl5oHychiMBb4IPvVFdmCGvjQKUHEUTUhMu7Owz8FwDwRlRhJMoo5
3PoELuYaWZwPy3hZ5lzCSUYPbty4dHPAM05wKNgC1ycoZHPDg9xgYMUXLIJvU3Gc
TAn8GtW2SY7RVqKTgTyS+clYIc/p4geJ8GNvE4CmMi91o2J7YRnNQ5NiGNTLUf8S
vvGfH/xHxCRQa8JB2aFYY/LTkPpxuj1KiOaQNwr5NXTJKb6yLrjQW4BTvzlwqNNs
v+5b6blpfvqyrEps4U/HIYj1LA7jRnayUyinkCrsqv3ufoqCk9EEjug4aMSs5uV3
vbvodBCdIo4fC8uAbl3FSNuUhfy8RO/mxFgdGcGdNmxzATFx8J/AmF+sXBQQAsGU
6m3OcoqATRkv+RCN53t22bGNRpuy9i8efl8JRMoJvYlbmgrynaBIdjXwa5HZzpJL
JprlDveeL64kpByejIX2LPXAfMRUC4RfU39wc81Z3AuKzuB9f83FrRUHF5S032VY
Qx8KLcS2J5G2bVYTktmiAsMC7cOWbX9zfZJbATv1pSiB+/XOGWnFuKz++V011PWY
VCdG4+DTGViwzo7Uyw3Rbi6XZVHOEUfBPZyWBaC03qPxsth9ZVMGxruGJJb5HtjR
1hZnHtqjKge07zaiPBZ1GyOi6pXH7dojNYe9Fvy5eeYx4GwpnO8clHnL01MCL//N
zSXMxflIlUCy9RYiEd3FlqrjQISGuFMflpge5oZ/t/xZx66LZj73lsV2SBq8ZUPw
oWh19Jv0xFMM/nnHaTA9VKeN/LDUEgxjYs9QungAB9SAIMhxLLdqJmc0rpg+sbZ/
xUJGqROilfu4jiKoe3XW/a23r1NqYWLzVl+gEzBWJKwjuTyFpdBLQO04mGCe42wN
0ha1BbbXy3633nTva1vX+02D26uRR4kSpau4YC95VgiZ0kVbrVPyuVyV7XXSS0D8
7QgFQJ3EdTS4Uu1cs9/cwu7sDtebpbI5AFvew8eCOcDXVDzg6Nt49LKstTgci8Fc
zIAXFigiw9Uz+3tzKMy3/FOptGlx7jmAQoGPBm8rF9LpVoGcbZyTuPmNDxh7WJle
PBLupaqGqOIEvW3KKePB/FkxMHMevExXgYXNGaDjiCpWq0LWpso5BJJSb0CjDeac
3zbmdWsaoxnbKaX1nXIWr/sYzw7nFRKae2cvJSjFWEGw8pnetJGV7YveAJMguA0t
rPYL7mgXspGuOFeyjwfkegssOBQ3mUsGEMbCgO7cR1io7LdHjC76kfTfIYmmoTCf
IrP9UHIpf5YU/4R7lv/fhaamfhtcOsNHmwVUSYrD3fQz0BUxVy94L8RSBJL1J2cz
TGniOI4Ebqq+Au+njK1eS/ivq6XlE+I6jHOGahc37pSTOxPKSf/yXGBLY8OBqDri
TFH8UjWDnUGSejt2aUvZikV48PCA8aGiSov9waBfOWd0fdo/ZJEIx0SuQk09X23o
qM5Xw6UFtkI22QUFUF/7xBgQKVKK2eVYK5X1zUHa0jtTN0Z04m5H5sheu4nrQPnF
Z+j4pmlZ0mu1+4fylUCiViyEKLGoDi+j2fduOi6TpX3BQuLH+ItMdsF/qDJoPyKS
Dj21vym18Wb6OB4wJkjtSChpkw6X5izBVqFf1fXlAJjTflrLfuHeFMT/WdR6EFV/
BfYCVWm60uLOLzbIB6b75/i/wYomhKZGF0Vd9gArZjTTqKY3LjUEFDZWihHGIkeU
VtbhwNDAOfIw4iLeuivSQfyE2i2DUB3cSPQKnw1RqbgBX8BNPDyv7CphZd9o/NCo
55HO4K5rG5aL1PrRwOtAXbnuo77Rs+wJmVT+Q/+fq3Ilg/DEngo1fv0UfDRJl1Q1
`protect END_PROTECTED
