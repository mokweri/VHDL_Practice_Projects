`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twi9B/gadGRd5zWWMh7CU9tycbT6b6T2eOe9AxVbA4qNC3/UGeEvP5vtcVmN+CJF
H/D9zOq4pnGTIjtaCvA9bds1zBiscyJ4KmR+7KMLcAi/KeU6p4HiNipzPuhw/NlB
n13Jp7at3DJrG/7CGffUkv3gQorCSFIOQmZkklEoGdusbZKewd86C/liYueOO0iC
aIZ7KIIc5luvzNrCxOaet8zWitgj0LHB64rhbB0PAgwXT+hc8q6b+WfKTd+Rn1kO
HLK3IDGSWu74UuCR1XFZhUehZBxcisst/1VeJy/jODMoU7InRLkrGDNrsexVY9R7
rBi0jqN9nbLEf/8PK1YAV+zN7Uxo4SU8aGdM7MoSp6W82uPY7kPd4WGb3qPfQAlC
`protect END_PROTECTED
