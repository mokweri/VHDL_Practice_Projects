`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efMnGt2DV31/zgFwohXJN/cY1T/AOo+4H+aeuPD9Eb9wAgA1ZUV+bBy9aeC1QX+5
VlaGyxue9/6DnoWOuZa7nRDpb9EUiRuC+WFJO0NRUCs9sUF0krBvNZbppJFkwehV
XfL1SQkZI4+gX/NfDwZEFXAPx3udrb0WgNW+ItR1oq+rt+IVAeaD98Xe/MSbmf7d
3uy9ueSPfUvzBGUzMPwOCfN73xVlSxHAfdSJVdavGWT95s3b+qcV441UPgBN1Nzq
EUqmtR0QDiHOXJBzjIThwDQEtBlb3Hp4A++AKJrF+FtuqWkyc7dsBocGuYaIglxo
gNRZAwkN4FPrGomCXdtwZVMgModziMzye19LmyPqtKBx26wZX8VupGj1bG9nwq0Y
hBSSdNIxsLNJ1y0RFiHG1TCawVlPuZWsLDf3QnZ9e3pLQz3xiRXhXEwEc9t8cipP
EWbcK7EfLL40QcpyRLqwQxwgVPiwcNvJLkNqABQCRZTw3RHlfyDeEqoDwpoyBhHd
xo15wNL/vPc/V/T+5fl74shmfnZMD8dPlObtX5p6djzhnwKWQbIKZr56RY9bAxYj
DIL47PgVa3tp5oLCCyo7MWeY1D1B+4ISQXuZ5u784ndyHYUFYXkOSLcKBM2GMCuE
BOv6F8ThszKMCKAmeXStSIeVU0COt9oexWKnn7oO0DoBKi1txTEZMbV/iPvOLMVz
4nV/DmtMT6bNeoAF3WoIcP2iwBrmKJ11WHrhia305N7vx5PPI9NYuPIGlYRm+4f7
ghmCbV8XbG3bE3j25h8QDMWgQxUAon2AdUJqfTTBx2A8TxoYMaTjt4FH12y0Ga2w
Srg8JSzo5OSGOYTRa/W/iJo0fW5cPG895pL8Q7OSEFBWPdvrl7vdUzjsUQdxOahH
HfvmUqy7TljeMov5EHK/fmdTZG/I6B+Ewc3jsONNV/kJP02e95GaBcfpCUOQGO0B
Z47u/fhi6g5eyrvqPLzCL4HHnlQCOaOr3fHdVPaPVY6Cg2cJswp7rTKaKWXR5D8E
pNmwZ2wjBuiFhYkUh6Ejge5vWncXHoHgHFciboRBTcfZdH7O+I+5ZCl2RTfW2cc5
RiYTnRMNGg7hbShLPHtEO83ksMPlCpEji2duUoF4Nk5fp/KlS5WTzl9ejXuIzzvX
IK/B5EjEhnkcXk1bylsebPE3ZNJEdBxOgbe9kJGoRomxPafnFhJCJS62VWNnbHb9
OWDrZD/EqfiiT8oLrraoPH9oWcyZX1L3j5vTlp1hkJznYtMm5/KTKZ47gUdVS0Ax
PAt8vR6iSxPfA6fRmRTWI+R4DRi3A0mUn8CFTkGic4NQD3+UL12i65YyJJ54U6Jq
1cPiaIrH15tACUAHQ+1xPNhEczRwf+NpHRkPxCk9S+L6HrUuFmVPVLh+bf7koSP9
AvpKgF0RjJ2rySLkqc9etwd9fjGIbY8iXvG/xAA+eL8=
`protect END_PROTECTED
