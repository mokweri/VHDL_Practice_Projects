`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tntAvljUS+J2oG77yht/AEISO0GWx+tzjWd/GvnCR5HKLCFZC/hNEeTew5aTU9rw
Re6Lk7GbvS0Rxue/jyucC/lznvpOCxnLtAcOmuasw8uBWXjDqKjonAjSOF6adRb5
2WI+pKRa9X5ww+V8Ho2IgjStygj2wLBL978IawX4TDaWdjGsDL/uRMD3+7LbgNrj
f8FpHGy60k7KS1HM9Gc4bSx3syw7O/eYI0x+JXZID3313qraB40Mawwf/W2wcJO4
6cnQtqbzifZIgHBlR6wgB7OqkkA7iLQ3Hn9RgXkHtknX0FI4GoTPResaw6wS4uW8
Hn+XsEUsKtINre2ZkA0xKqCxC6zA0+SQ5lsUyof2TOrP/ttGMePYUMeryeeHM3lu
bwlwOmL66Zzv3s/ieXdCxXDGSFp5j1s4DLmUfO1k/2mME/p7B45RVREs/djTMhkH
Vhe3EP5GZ+XBgWLR+cqpbz2LIRbB3nAfIzPRL8grOpynPrnaeXCaX0Wfz9lbxGrp
ot93Iw4ehz1nhl0iM6d6EVe0sSu2Ee4zE7VFs9wOYx3lZ03Ig14IDv6/wJFBzJ8y
HSSXU4VsXbPthCT/wWnGDnePawguijq6VT5Y25FBW33BDG+MpjUX7eVVFkxind0K
6rom8bnIC7ksN5QLa6/MwOrpCm0q9os93tSEqnuOOwTolDr3JLPsweg0pYkwDuW8
Kiifqf4StUz6bQpNyPmDBo/8eJU2sNqz0sbbEcjYf41Dw0DWU+LDndV8laaz6N22
334CEgzv050nZf15wdM0y9rAHGYTVu/o26AZ9tU25jLhxNR4isWBa1lT2RJi2xMP
UatSvfH7WylWA32H0L57lVsqsTAsDxKQ3lQCEtzhBViEOcrGl65KTnCwxH7knCZ1
GRQk7bJMS1tQ6c93DO0FMpDeGfYmOlr3BXCEmK2Ef5kzG5eQ4YEbupLpYfTwuFPr
Ofw0aim1U3gesXpRrtuL31pn0iMSSZvTuVDrRwq20PG6ccrFryT+2JJCC+duGIcK
9csAkc7N4306y0fYd1hhKfwFPNcf/sBP/r5uD9e5dZVEBRYNoP4HSSAEKUuUm7zq
YeCmR+HPRzOu8lWeS/nm7iM9JGIZRFpjLL/gtB9hsYmravr+8i6MUpSMgGCJDQgv
KeAwgkQ456MZKSjlMRLzMTObNs5OKKFTdU5nAVJd8cM9QpFYxgTUGqFNcHVFR9Qy
8U3BkreSmrfCoumz3OoWj9kA1UxcEdO+vS2xzTiu04sVA73RL9cOAVxCo4o4+Kge
Z/RqJNZ34GegurrN941QmomBLwHSgR6If2C5D/OhOK61PaCuQ71eswnzTPqtbYRG
lGIQ8qJ92Iru/aJPLWQeLPjf1NIwqKKSl7uyjoJisJJlvoBGS7/KSg2AYJr8oqGx
A+TIIKFpyfl3Af94Hm/PVpOy8G7l/yVaDYuqSCFs+2bka7Vo9nESqk6735v9i48l
FxxMbWWc1wCSwUEVNPQqmAbbrR0t/3vBXLSnt5huAQFDXqTGyZywoUlhJPFkc8LK
rSXNDaoeGz77nGacaKUhueoWGTHQXWRdGIc7xCZU8k2q5UwWW8DpEWJlTVUBY8We
spL2cNnAXtyCRSdv4qwX9xZux23NyX8tNdYTM4Q2dONV5Tu0LQHO14xGk8muSTZx
AwxqI1GUlW+C69kzOvg/2DkzgYZAOgPzOM6nhtxWoSjnY9jUfIxI3Aht5dBhq/9U
ygVRsTtbvyKMA/WZlOInSUHjJBMJ65tKVZjnB5PipWPjdZne5AiO1A4XzOTRZ3Vj
rETvG47W41bvUnp73aapziJzGcfZCjFCOg0fzmQcc2e9w0q7N6qmLNvWSW32EX99
QqUAGZOnT5ehGO2GUqe0xH1r3bzUhj789qmeaXe2ev9HDB0dIzN9qUN8BFzxmeu3
zQwSDnYtAhyDXm6oxPhRYQQ2bTqD/j6uVgLA8qlajdR35RaemFIH3cIWwDinp0cq
e9POp6OnE40HWwMqWI3k2L5TBaBtKTztY+/KAx/RDc8lzLVRHoGQFNFCv2qJIRX/
QJ/Ij/RvG6QS5hHLfNpjZD1scGuFGKLNGwRUCyBp7umodWQCWuuMQzp9xyEtkaU8
Kzg9q3NkyhgXD17KUih9cdZki/lW085zJeJyuwtnmaAQfRvf9gVFrCyLD/Vy31Ip
kWuj438v4/g1orR9Pi8mIJ6ajUWA+udKoWu3985Rjeni9LswQOxihUA4f6n5ZNt6
7JIXi+8qnO3DI/ZJ66c/a6R5zJdWWPKo/wVDAkMnn/QJy+iKfS8mRX94+I68GaGh
Mc66OsS2igMGpCSIjvQ/vRT7/YtZlhzkbSxS8T56xl7BVh66skGTyqt/OB2xYdp/
/DnlVjhcqvI9O8F9jRSGx7v8e6U/YPnoMZjt0IMAbDdm+gDTaZgkLNllcyjGxAxe
q+S0lsFeMK8UK6jZ0poTjj0x0rNyYZEjEPl5xnK7JnijTBIWAJM5f9BpNMeDokHY
UrCDEyh70zo3WELBdpfNZfxFiPpltt1r3T/2jhmmQ2HvlKlfm6Sq5uywIgQpTUYC
m6ip4JHqNXMBoL9+BVV/2Z4sU2qrchNeg3RYp9pNyjGbz87jnBxxgF19jzpn78Z2
meFvx1VjLsFOA5I2yNjc8Fhx0CLqm4IPGJNIjvRxsXAhzVWIXKbNgShQw+qWYrKO
HwprOaG3ZLyxu5g8A8utnrwRT6QYJAfp3t3O0tQYDWCbWoMz/3ogxDsqcQmKlXC+
lSIbXQh1RDBzhWkudoPAWz23QAYM4oOrlEdCtXaSrAY7djBbC8tpXlhdD0hRBwoe
ijSxweYpbTlXprZrBKssjHyu1zRRY9wmF92Be4KVIzzMiHl2LjVrGYDhLhWjAuiv
bRc7ygBM4Lo4GwIJMlh5k9z6He8dT7lx5f5e63rILSL0RCnkl1/Nna04J+6GmPUc
bhMZNuaCKngXWIdu0yxkmXIeTI+TN1xOkdbXdr6cCGhvjRFCfi4bmLfL8hVSB+Iq
xf6E4Em6NAlmMunbWhMD/gKPlBidvAgLF9FxnjmFUFOmiIN/7FSj8JHZaWjCVqeS
WrqwVYRLEHnTQfYxfCbC0qNNvLsnpSqpaPpw1z0Ejsks7oMosqk5HUdxxz42mHEp
i57Ci+BqSkRM7+/6PzmZOOs729h9MoEHgSs6fz2b9hjPbwN92A168NYfhZcOrxEw
xp4BOWzp0zxFnsQ2RnNvT7fBSy/jWb0t1j6q/RyB564ozS+Hcs8UwcxD2ey4xAor
2fBo5hn0UFseeC96XaSwxrtCwaGxsaK7Nh6LzzHfvuCmRPadONSfwXeH7hqbzxYE
tPtWTGw7tALTtLN+VucasSlKXr1SPoz7lq5r+H9Z5bCcCvL+sryCI+IG/QJ9NVW0
x0AQMaDpcDbU3cSOxYik8Tsx13KGnrB7Ltu5UNcr6ItJimNJdkn01NkT9IEFUeEK
s5Fcn+2yV1FQyDLzmQK6R2dQiEFyLRMjb7hvhrun+vuwZmWFjDTepSO67Z2wa7sd
rPz3c7OOPL5gOv8e6GWddli1D4+HlthFBE9oBUI9Bw58dfK13loRWPEk+qSoC+mx
7ds2NHx6nXBMMyqwqCC0VWWDrWGfx6gBiG38brcGA5ou5jUZnY77yiSF+OAE7NBe
tehB4ZDeOOUZ00vAxmv9s87GwKy6WOB56EBtXx18IjNYgohutJ6cxM4hCw5N7P+h
`protect END_PROTECTED
