`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
toBbPBfKma0AnztPO/oyOyW9KDgKhV929fRTJNmMjxT3GpGFrc7OxBh7v8GOxjtK
iUsVNP9Wo9c+ESqfWD1UcXWBKWen/ixDAQpO++OiG9QD9CQT06rHkHv8EMpoEkGO
jDjxq2QnbbJpKOtCXT764BgIcFuOXhIMDLCREaN4iEj9IcmDRAUot5NG0PUOHBDE
ugtQp64xIFQNz10Il0iifZjz6+GovfmNm/KCweuAX+iai6NK8eee0deMHhWlkkax
OZmnAeTR33pO5tg5Q5glgwvXQRkBSUbxLVsNUrHNebSyusA9Nco9NaaCqaPZDAww
9hX+2/gHWOtlwdYH5k/ixUSBy4Nc770C1PS4+ekACh3gZEX7bhuueEjjC40TKHvF
xdfqFc/4t5bdJxRvS8bzC///B+V8AhhfBMmVNRFcLA2M+xNO15TW4kIjYJPjzrux
WfaOX7XUN18GjEK4xK2eWuWJbu9/ZeIWs07VuIBMJh3UW0POD+hss4SpOFwjCXHR
NZExtHdDhG1NUmoANm+uj5ZtBheQ+cIaDYIX3I9GbCu7DiFsJTNk2kqMH327cFqH
n5jU+z7nwnWJnhuGeXOHdb1chqgXk3Z/SYoCKi9e/DfMcwQS7N9n0UtwDfGv0Qca
qOFdocGUTbewthjQ/PLxLBL/mQu8UZ4o/1vADqEaeIIJGibu6vu57lmbmNA7GgRZ
c9USA9I2os4NUij3NmmVGWWHHr6V843H3kFpwnPxRFVMglrt+G52RXUwnIugoI38
oXOfV+X7LjQUO8y0LiOCI1c7TkifXsEwBMb/xyoFxsH3eJKOuD6IxYKClfKZ70IS
d7XmZ2YkX2t12YjZlj1BDtdkzoyRtOmJuoDz78xRwFgbOKNm370llmNgO9wwqB5Z
s4vgq1aRMPhr3u0Tw0kJ8vQb9bwf4v3yIVHzKYaEccZH3UY8/MUBd5/ZUOyeE0L3
ykQ8xkVULGXKEJeGqkK/SeOfBvbUfukQygTJr+wbZFI+eDMRgYJo+j5NKMK9isJu
4BMnoiL1UFTIPKoDQxtmEw6LO1Ei1OLnKJLprSIm/EwNTFKxdGbuyqOaYCtk4X0N
NQs8isxivjMVWIRQ0fvQn9/154sWAdl7cYMth+DHOBGlU1LsszCk+F3TxJaARnh+
y2y/cboyr92tx6PRKJxgxgqp+yDwD+QcfVm/alKE2bWMz0LZaIpCXazrRQxgPs2E
xSonvM+nv354LgGe9/ECQGjEJNmZq5NywOSgNMJZRThhdjFICWXV6jg3NXuHZKQq
MlAwVjuxKQjiMzU6HhxiNa2dk5pgPwHHbqTSHKjHdaID9ENl+cByhex19n0EFs+D
rECKf270RKKBt2N16bfVWWKGsht/9fXBllSYyGrAY9bvUErBPDSc/VaJGui6vNyu
qsPUALuatTJQTfUapwDDK5Rc//xlqdzR/rwbBt1wAXRr+yfDPSz0m6VWlVMZ6tY/
ndk2NJOOrbhE8jp4Zj2H6SaEt5QvWuQWXLO/dxP9sPxLFfGT95z+W8zJ8WZ1tL+V
ieMKZY9dgICT/I2tuJVuwm6KzW22SdNGARLtNGYveZF8XP7KIc0h3JleTV1uNisq
VlLhNG813/0ggOy8zrxS3Yo79T13tqG08mihUm8/Zq9EYrD8swEMPrHSASfZlv3E
lrKO9szNgKqUdm+nrW8UbGo5NxcQI7yvlHndd7P302WL98L9yByAzy0FPRPaAD9z
Xbj/iNNDIPryIdS8e+bRSmWant1NRRKpR9MWSvPsCwRjj0O93gSmWiGxFtBemcP6
dnDvJ3mHPrsK38GB4tQBhAUqwghxNHCtrI/rCTKhFCrcxGvsyya8Y63g4YTsSAlL
VgaKiPYHsGqS1CVaEpTAv7eDZREEYWql8Z9UGrzD5vHj0LEovtepRZefls3CiEfK
XNii6XPs5MofRBk9LXauZJbboZdRuUwUcyO8tC4xsGMHZJ4iWAFKvk8c+sLT1C64
K5gJE00NEgUsxr5IFYYED3vIt3CPsqXZY6cbl3jNbQfgaHGCbkBKH3Yt/vNBOPEs
nOtxFtXRtpgieE35jzpEqVJQgEsrUGdBwZIsTr2D/1whB2M+3udrey74HeUQL8nk
p+4VmI+N5cYL+Y+l43dTJh2Y/jE/5pvR9RJNVky8jTS6dkFp+gNg34ErZxQPQIHe
ERojV+8JF34u0cdqeC8n9wEpYJ+HGceNlik89tnvdZ5fBKKBzPVKa3yuNfVSAdtl
ydTsoFORBNK6rzwiJoaLimZ6dfPl4UGIcTNZ43Odszum0hOWSAitAo8NZJyCPzcc
/aJU10Tu4gqFLJzYw5FSHMnvMyWU/SRlfuQfUjlJiX710tt2oRXuD07dAv3AhqJY
pSJQ9Wr+/Ly3lFTw2pYD4LRUyd0qtdV1ERAczRGAVwxFHwvVbe2TPV6a4VzRxMXf
WV6ZkrNMaTg8bJoEcvxeKpRHy+ug59ofP0yKWIhhO+mWC7ONUcJhhkwBpqUqDEYv
fGaWzcbaIUnYSf9j4N/Q4IYCpgshb6QnyeYhj/+d+kl8JShW37W0c7X7Szp5W6It
aERcjswRbvhtbjvDZSeAYrehISqriaWmh3o42hrJ9WtoMaHatzaqWqbGGp41u1nn
yB+L9RNWiQcGULKmqxLgjR/eWa9eGZRwxquoEDipUikSZZXTyXofeHLXH3m8bBFd
JrgEqr/+c16nNnIoyfdRKTSdxW4Wb3EBm9wOKzrO8NfB8i61nzlspYNKpbbwha4a
NfjFTJGYgI7miYCsnW/6b29oZ3/5jHdor6UyEC6k6HyC+sbyRTVx2ielygMiiNAl
ROL01yJ0bjVdOlpoq5pOBTykff68VVeHHV3q5o8ZsloVTKgkjPs/xwX07ZbbWEZp
6HhLhJgOw2BGFMAJKQQZSgZRmJWHdCFYxVkvQTJrv1jQP5lD6kVky/5eoF349z37
pue97tT9GOQaWBoQPOF6b1+Sh2cx7DFfJxtS+510oxtk30XuaO+msF4rgU7VRSz/
0TuF6MucKQvOnH5n9dqyw6sBJ0Q0YcOY3xTBvA1lDn/Ocl3YAM5cpVfe9l8pm32X
5iDIpJByhwVE8ARrzy1rLU7DcJ+sAPS0Kt7AxptkA+irl83LRI4QZj0s0wwNdWZ2
ST+ZokgTj4X2kIlXG+8aQMVM9eS66qPpKmlpWSQEMSFBghlLANm5H3bJUUWUzjya
Q9sVMstlhfrqoV04Pm9fng1VxvDFO8pjePAJXIqMdb7uG02UHqsQ/spRkH6g0+wy
lQGL77Yjo0LnPGqHUb3y+wW3pOd6AbRjdfsXrrVu98b+5dXZpxcQJZrHLsGPMnpw
E9WecMDFIMvueeHt+Zy2UtlNIxpcL6cJFink7zA9eo+OkroxPWuOLg0D2eqpm3lX
8x0V36LVHner4TSquhj0vvPiWuCYd0d7m6DaRk7cJZSqo8OE5/7ZYsvkZvBxlX7M
BG+m8hTCkMsHrF2Wv9SW9P5N1o8P28aslzUJ79K2n442NwQ0eRrqOcbQn4AIf2/D
q5e5mGbtpAC6AohOcF+VI8EPNl2ZxHtuAY7PkN/1Ae7WTJY4p+wEJ1T/nO1jegpO
KWfINtOzT2TEHrE9V7aLKk75a9ybpg1AQ4+0Vn/w1uSCHNX9wMOP25JTO1Lq3Vs1
GURGX0ldrw2PrXybccaxgXxUA9MeKpM2W7V6IwlpyxObJBszIgmxGnrTxv1SRfDb
i+3W5Z5V4FKZPsT9nxNEyw==
`protect END_PROTECTED
