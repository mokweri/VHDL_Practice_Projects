`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxjFigMZFrzz2fTQM66gwgaxEhQ7tKGfdbH52Oc+wvecL2wKfKLfdyMTAC2zsy8e
Rzm6yuQkENqQwCEuUYBjgaQqN2+55PTfS3AqwMTyZqkHhTUc97w9cTc+ZV2TBkQb
OXKnNR2W82Du07yRVn9sRIEYxrL88jbhbFQ/sMrNpkB3vz3tKkF9whWO45R46PME
O5jQk6Tujv6ii16L18LAckVoPXlKVNLgpwUr3tgADMUvyNu1lHvwDxT74kaxslY3
t0hY7hZagjFItM+Szr2KtkeYCADwNkovxi5Q6G/I+d29cXWxU38OAFevBEJTs22O
N6IOiw6Cv82Bl/iWbIevcQGPI2jWbEANEhhMxHNleNMentvriic7qunGDD+VoWKg
sD+ybMr2cojUgia77hiZtpkRk3VMSpw6BXIzPbcsoC/ChtUJJBiORMlAJtynmnKH
QqaIxkYCcBfs0ERGC0mc0gNV/8HFGYhxQk89Kb2iNPt9STDjygiz8bu9GZgRGgO+
V6B7Pnv5NtFU0woGcAw5mo3fokk/CaitWfC5wc7OJKqz04BBrO+EfHyT1llR/4rF
Mxgqcn+66g9zeOLVDGZWDlztGCnCYtq6ZW1FRg6mz/zykiIdy6Kf/VozbJCkMPEH
jNjVBv4zOwPx9IbtR0R8+YLDePxCGraJjMJ2pPyIndbsBtxBGVcvTddv0cQTtygV
3nnwrO1Oztivy2Psu8wkLhGZATUmizgiQfWJRxEU5nIPJMBquqZO8X+VkgIJBcrt
OvFOZe80u84V+Khw6JO8ge7NALFwbJ/INVR/SPQMqslUnVp8ODWeHoXl+sTOFmXk
J941SRhAch2VJeVpS5pipB4TPJ/hDmDgxVuJCAkFCls6p8l3DBz3jaV2tDr0N2be
HI7qCG/f+F7c9HwqZdrCZDotMgSQkgOM8uhgiJGBwKE+U8TOYlSI99Od72THIXKs
V8iQEpZumyeh6ueemjCuHlK0qhY2w+3aSc0F++xXlwkxaWZDjZL8CqgD5g4NQMNR
lBWJ8dcLIZAXKbP1HphqQuML56oJjlNmF2uPFW11G1sFQxbwN5pz/dsBSqXjx9ct
qe9zNgAr0+xoMenOQW1wbKBNUWTE5S1z/fSWDOi2wDFM1+X9f9e31HsfmUQFmQPf
KLROupA1/6ZYfh4cxsPRgBGUmVFcf/X8+i0w5JoSSa6nAH3sXPzLgd/V3wptty6V
pnHcV1C9lkmsH7FiavFu+fNBGuG+rXw5E/SO1dMYYfR17bCypH64fp95+PXA296l
CYqFAoTIK+oSqqswC3a5XdgWarC+8fk3RCwJ1svAzyV+NWe9qOdD/xxD/dj3S54I
84fDoKC3Z6y+evDxJ8BwrzGp2IJbPErq9uPzH67th4vUk+qrPHzqm1jwZ38xZ6R9
pKoxnAWxocyy/r7KyRBuuZ6xjh906ixPae1piUSqLcnuMGnwuez/zSH5vYpKZhF6
Wzqpmxp/hfTF0fMjxhjLmqWsxXmoZSngCf5EpBESZ53reNOM79xROqbWqfI6XcDw
0NTIE92QuZFuUNL1Cq77w6TXqlVrlTMcz1sk79Ebx0tihmJWzzKHvkowvWQFn1yx
14T9juS1cmc/sgL/eIO7Wd1xCF5Zy0Ah76IUCxioUkfp8eU33lhRJnlTFJMny/rd
J9+79qO0dQTi+paqHCZQjWxHAA5p9eh/L8qTDMrHa7LvBkuY+MJPb/HAib90Cfq6
2aGr0hSn0HgkF6sGvpwJska9aDppk5mT4jhnTICxVPYPTACa4H+RaJIwhTndKiOA
Qi7Q6NVvc0DP5l23vedad4qzn9cgcrZTEOLmC9t5ZYhR2ThdF8abqrCZS3YtO2XA
wrC+FxCgHqPASzj5kKLB/jxM4JA39J7t92BsrtRwJku3SHJ9nj6xHcpo+fn0+rTi
zmNSSglDEtaWRRSBKSbRRoB9fKBPkpLs5ijZ/Jh9hJ/7HC4C4gkW3W0EwUwY4g5q
LXt3+YHNbU1usgHLh+KRGaTWIBvIe343UUnWBWOmUfpkuWUQDfbxihtziN5CKeD7
ishkPVpQQd4FOkVPe2fOr16JfSAZA/iv+WoRSGec6YZzgoxX2B3tPmgFlKd5r6ZC
nFQH45+V2Akz/6CoGZepYRRxzLJaFpb5FV+RpPuzU86FzocibcxSzgw3N+Q8SFQb
pTEarakr1YKflsWfOSbcHoRG6XiZdzdOJq7xUjQilXf9iD1bdDbW9xjMUhNTDRTy
IWxIxV295EjV53HdcYByFlIT+OZfq5Hfz4o67VvYyxHIoTdzSc2/C4n37dTKtsTI
uoZKc5FJFDvDhtQsL/WBzReASioxaiEl/xiu9AG78/c4ktZoZbeK7tJiPHkNfZzg
0HVA3Y66rh6FuaBjKRJK7Hg2DuJXXG6lU63nNY5bPpEaoA2MWPOnVMJWLB+FR1wC
6Uog6O2L/BwMuUDzxZsk9AE3BtowcT8VZ7ERd5tlBx6ZTZqyfPHQ3N8VtLHF0pVq
w7oqw6SSma/qKlDPumsywqoWX7H7IyZYWMILKFveNXAJFLIwF/dVJcXddhhyVx7+
yEaUrtg3/sq5r3jxX5XGa5ZcfDBPZtrpUZ8pngqb/SgHA7a2uAiNQR+uOjjK+MhC
AkAQ6sItj4XMhqF2QF7bqFXk6GyWoe5IHaJ6DZAD7ktSGxUTiMtMEXluSQ4dXlb7
L+TISqgSrcLe2xg3HxRiWoK7oh8l/5ACLIpXcus27Vjqb2Z9ME/4GfMVB8kfCQJz
+PpqC8dTzenSDF/92zoPaUUFcRvemAZL4ojI1XgyjHBZH0j4cQT1HqFrI+zko6mK
rbMB5yVtti9mBEKuvaHYFBCazpnYbRfJKa9/bRxRKhBbA7y6iPg219qiNKE8PXvn
I3cQ6EKVrx2Dga/pAT7yHn8Deu5Ba5Kuswc2BkqY9JTRd3r/zWlupITXdBJLsvOf
++U79AsXvjn5SoMAYqLGpuaxwOAgIom0uDRXxQox7RwshJ79b1PsyUxh1Rt64Jln
rlRDVx25/lGVPfNh1ScLERJfBxwTcfSl8QTh04Z1p+PpswryOJQkoCuoY/V4gzBl
5XxHhakEbNWkSQ3yPDlOAuZyOIo+1jzNKQ8qNP0RXZfRmgUrWfdF8ogORiJMqgYS
LngNp4QZWQQrcV+WCSkQfubX76N5+btcnBo30s+Cp5W7/LdILOwe5STa6/28/ns5
QzGFxx0OQinXFPAWzLEfKLkr3CsKYsCk5sabqgPqazp7+g3ElVLiyE8v5KRjpf+H
f8bgUf7s9pze0Y4Vz/T2NJ6Cdu1Rsz7gi0ZxV3/QKw4=
`protect END_PROTECTED
