`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K4rPFjGe1/yOy6XM+a9R31sZGjJeSWKPkeDVcUh7XbFEWzEukqlVNQ//3qO/Hhop
nlNp00aR5gW6AeYik8GBbq9Q8DAYojrPTVh2MhYmhD/M4lMI4eAZM6SjIZJqXpbW
vw0b0TGj+Nrl3wybH/UlKcK0AeNHzu+brfazsfaUiniAVVociMeOckigqyY1xegT
MfLFEq1cHTo3Gkx2e9PUXX1wVZzEPgCziZqaoPuGS3bDn/PgRHUyeNmLBiSXAhAC
a2DpyTdf128ot/NUIPTW3VX4O+g+XfrDWIUoiT5ArcfryQR2BDPrScbk5v2M2ISS
Z1ShYgjtYFFnv6/x5p47w0TNjh4AugjkjEMgqOs8e3ZAwRWpWnRgsjQLHDWcdxk2
Ed8DTDlIBPado+D63pVE+KiBOZMVDA5zTFjKCSn+ciC5KwHrtiFkj0AfuWQ7cmTE
vwhgcBEgHLlRGT07QC4nHCq+kfegM4WnHq5MuuiWNCuazox5ZzxBIqiede9zQJdp
rt5+Apo07hrr2JF+w24cYBfiYIqg5x4qck9M6iZI6TUaYpmJpct7WbOQf5v/0IyJ
5WYD8q8C4mmXXpeMO2JkL22JKyqdVJkUPAYd8cqtnLz0DH0t929PYpn1keOxGh9b
m5qJX3aEbd7+/pRVEqQm6/+3tIGlmzJBVEcY7ITXBXXLxBuYcoMGsUOmc741R4nm
uOoeVwWeKoxGS+PwvWQtbMD9I8ly0t9Mx7N/hZsdzQX1KIxUioS/OJypNcDvVOSW
09YxhlhktBZ8iZ8+SgyQxCelHfRDpMIE3CH4H4HqzsLqV6s0FHB85etOHXfqlYc5
ofa9gRcbvz6IBaDrF5iqLCT0yqyUuZNCQf/a36zWER7ZfeK0yevZV3ipk7SrEkmI
Sx8qCcLlsnf2VmFFdvyxxP6J5y90/CyJuObX5wf8aALXxrDt9Alh9LTl7Tn7mFl7
wifoRqal58lqkg2uRyquHytBOtd1UAMq9vfyb5HAbbUt7JADDrB/xDf7cS0kodJ4
M+hKsbPqHlWwHcNOWkz25rZlhrNs5Ujb16kvravvr6WMQAKiRtY2O2MFFQkmtFla
Kgxd7tuSm2abLIi9K4ipmIy5dTGO0JT4+A3hn+VwTpuMUs5ZIshyMH5hmEU0q6ck
JISY4egTtcKj9MjMckSVF8G6t7v12oqx2PzYj844OhW6cY/a1ungW6tOr4ugv6T9
2aLcj7Ykkv150dVRmikJTiSx+7/z8zJJBEwGJsDWApPqyY5bt+SL4NnAnNtvmj/S
NbEfzoLQT0bi7njPO6AGs9fQ7F4eZ/tk5nwynWQ/N1Cn4V6c5CBjE8S+gM3JBjC2
qK2wMPhZOVP83WaOIJhYBsSW1e0x6jxSD4zAB6Zs3gLFrzdcJ3Blrb7HYuQLqtI7
LkFNDPKeJNYbzlWil+rFtAd4rZjpQi+OzkgMsxqe3lgBwYGoJ8mF45xOoqkJYEGG
DnAZ1k5Sv1Sgh1mf5mM+fV6leHLgxxQnoh0lv+7V8bnXBGh8l2dxNNt20jJqshcc
li/qr2p/nlVi+BP2+HjWFUnrG0AlAxgS8RMFMNulUUlPwhfPA2I01IzdFeqSE4aR
X8RJAyVMBffQZuFshbAUNIpYFLUv5gLJZKFkF1knwlnD2LFrEGznqEOkpOucd6/Q
mtXPaLJEG/fdEo3eZUIK57lET8wITy9jPf9wD4RHIVtlZGJmRfH0N6ANbjqGgPtl
fdVC6+crtvn6mcr8WaoqwRkfL9rNhhZ65BRFS/S7/5UI59T00MM5P/D7zPZgwhe3
ZE3kBtx9kMaAVbH0dmCLdPsK8ZprcJC/gffHXHB041DGCv3BkCamGLVgOmNlQhEa
w/4hCXDtA3F0n1XfVsmYP2HIJ3KazmV4SI12j0eMgYUyBBCuP1GEW1Jc2WxdTgKY
hIFBJcLRgY+Z1DyJ0svfyZ3rkVCnU00tLZulWC9EBj2ai3ZphShLSgP8E8wfpQOj
Hw/wnnjGc4n9QkIQDfbqGakGFMDaT65cfiZqg4F4hcSz3DpGLGtGAMHJu/hYS6nt
cOyvY0QJsOFniJUsugGQF94gEr1bOu3lwqlvsKBVt124QkhlwSLTxc3xAS1g1di1
KQ1T1NNMHLKY3Q3T7ccq6NysJk6+L74DD4tvik/b0hXHzoBl0f6r/ZeHB9JlMfMy
AxjphpTVhBQkCb/zfahjDn3iXH9q5KBL7JLSYjzWfBbL/EegBlnsepDhu3oLmJxC
saeMMUZUFK8wE4QhbRPzPK/jwwFGETneQsFeWABR/Ce+q4N+s5EX4GW25xwE+dr2
K4JE6zzHfXeurYprtaPnfVmauMGkE+xUIg1gULsYc163J0TvL9VKHMyF6Tfm2vbQ
G/4xDV2GuQbCxDMMcwssKEJ/5oUHLwyhChqckLca77a0E9b1uL4CaM+OSQIOqg4o
Z4Ccr41XKPj8uumnMzhbyuXOop/2FYWmy6sZZuB/Ns2MfPhI+n0lQYzzlJouMQA2
1lbWGO0MgTAf17XKmqvXcM2ijvO6xoW+08I6xl+xqF/VxEVFWZzzOWSiOCcqttMo
TDwb9zWsDbZlxo43j1sw7ZE/X6WIPCn3S/BqPqvAakI=
`protect END_PROTECTED
