`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dv5BjBAQVAWN437rHyPBfuN6X0geqMqLOaGJttxts9FPip4xvvbiqgg7bwhx8RyQ
vROLcg5Bkmtlgf7O1TYtigoKHNVTeoDb+wtJfwhqObd94qwFfugopCzilRP9gQIv
0oQ7u/0pPsnG9trQN27IOw82DNCqIwIfP0m7Z6SHIKHCoTVCt/3vRVaVXt/1XSum
ea7zh6tPco2SVU68m7BVZkw+oZbXSWJNZoFzQMZl+emOQ+F2QvB6AVD9fFvkpcvW
x1KpuT97CPLxQVACPq4d5eg1hvNEQWOIa/1mkoVYgJew2AT2QTzI7ZUQpc2SU8vR
WWF5llg1v1A200o+91Fx9P2bgTf43zCDgs7CYX8L54ZtKczkBW2FGNQpjYhlmuZx
lpqCsf+Y/oeKYaQ290vlVpH56/EQ7RXpUsvUaGbthziRvualGvLvmo04Rg1T9WjR
/n+dyTiUk4nvMsEfQskXdiUAW0umzMxmhvJEIVkZ1L0Cs4KZngs+j2v7dDfJIvl+
2h7+iMZCRaPNQiQTeKBTiaVCNdstT/4pqhaiW4VtFDKhn5RyEcxbmmpwsPgSB4jG
HoEu4pvIJVvZ4YcaCrnkJjL/Mc/GA3KZ+7EhQIQNJb4SyDDZUXSUS5/YXndT9Du8
pxlQk9bnzd+Qhb/LelN9gTHrdTF8OWrZU+3vSxwnQdOu6YVXyA4uI3ryfVPpHBAe
znqppvPl4JE9G2OGtQ4GiSIdrXOBrlBe2HUkn46S3wZG+dpbEmJrd7ajl+mzkBFL
Exqfarm0XzX8h6qjkk/hJ8tUnxunPY8VWsc3yvVzwLudoWAY7tqpvQ90LQqwo0tF
ledVqK0f1BlmxmnHLXuqUUto+Lv6dU6t73+/zOWSfcSVg25zb+dpPmWh9SiyCWeZ
q3yqm71eUsve4lK/fwjI4TyxrAHNRmG218TCHkmvms/XqIa/5fRqeKhzhs4bANt7
HrOnbTB0tIRlPSWWuCaIFQLs/6vk4WYPuh83J+1lrp9oLrI8AuO1frSrWBFb50h6
3svl0KWOIrmjLh85RYZpUwtabA9kKItIlZGFlr+b2TkvYeQgtgZ3SHSnpCMtLU03
fGZjyWe02V06INO2O7fxfT8ELg0ViYrVy6/qpAhOipChbFpInhW3zl5E5U0VER4h
EHHUbJGnMD4n0ac/KFU+U1h603BfxlvFQiyGP+pAsijlNo4TpKXgDSqXWSCGXczF
aOhiJZ1FEbdIRrXVE7ctWz/vAVhoeZqf4PMo5ZPPLmlUDto/LG1Mbh/WLjt3F1rE
LBtSBLpNzRYXzEALCmyJq5sISRvsUjVgvuImRvbEZjcKAVdotfkuWWwzfJei1EMy
wiOm7LtS6gZsKIMbDsonz0Lr5ZDe+Yx8WeycNGvjvnO1THKRQ7fVSsm+FE5/u+JR
LY6mOlSiGKlqKrbwrdeCJA==
`protect END_PROTECTED
