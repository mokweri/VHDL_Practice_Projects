`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y4PdO6t6DGvRTaKJCbdK1nMv3iZVrbcwGxUTT5WZv2LAge1ZbeCfBW8zHD4RzC+1
8r+iiQ+Sdi9E9W9ZHk89hqECQ2q7AGnoPI7lETgDojuJ0SYFLk0mmzfIplql7xl1
PqlUb0WCF+YxOu+wUeHFqbcimUiVs+asdNiQc4AOxKjXiRim3TKXP1E94CMHAQyt
vZ+Fu0SZVkkVzU30hF0Q5WeKnT86DU5h5wGvtmU+VPYtI5EJYoKVkuErGc8X6fEs
3LYy/5fpP7je226i+Krj/vr2UEyrbdl/T8hSFrWBcdx0MBY+5++QAMeERzBAWH5+
NAJBEexl+DJ2/xr8m+DTJhCtdnxNCJzyatggCyF44FC0EfrJyIWoUEeTQf9XEi+U
9Uq+d0Fz7UHo6NyFTlipIXw5hW0udJ2rznZVkedA9eKeKS7J2CPPKyeTC5cs+4x3
z06lBM5XXaMzTjO+j199Sh9p2bjXjgzTaZVE3OZZVeUAy4Ev4TIO/oBGgEd0tWSF
uNSBJXQIykw/Lr7Y1+9dfA7vQvyFH0bdE/Xb7JTDcE+M2bdz2+ZfpplpGc8fleCs
yi22JTGgK+lbSZRGO/uDlQ==
`protect END_PROTECTED
