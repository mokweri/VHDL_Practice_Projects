`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5J/mugOHG3fWHkuhQy5BxPeXqSH0kqYtGgoDixN+BGxkpk/FmmNiD7rPEv1zPVA
LMstUK+bunefGiILJX9DwkWky5erl1nGa1/OKuAKmcRkJ1m7xS/82K7+3/8tfLBF
LLsklnnZazfx2HkXT9RmqXB+LT2FP9YacrJbowGjsu41cuv5EanByjxJtjakjTNH
f5UVioJtFB9RbVbSVhMUttk8UHMlAILm3jbdQN7fnuzbLKQqs8Lg4UlSlFuJ7Mkv
HCoQld9o0CojZ9Yi6w3Q7wTQGXuSELM6WyeYAg6hc8vzFG3Lt7LltaxboNtyACnv
cDt55c1GsxICorHDFZHNCrK26a80gwh/SwPuwljI2lxUh1Y/0bkYfh4bMdPkCZVy
TmsiISTc5xm/KTWQebU4D/vB6ifuQtsyK4GmguTUKHHAv1Ad6audBNGPUVJ84eWO
MM1iPlcfjQpEdqVfXFzT3eOGu5eE379iOUjqEu4979mkNVSIvd1voEQyRakB7tJd
sKooZHlIfllE/UnrBZqWSMXbRvGhk/exdMFF+ww0R+mSXz4KSLesabwZDjTD/nMy
53QbRoRMFMNYyhABOwLae9s8FzXaeXNNzVFaWIIzA5PSgIob3oUzEpqPIMIzLo5B
EW+tEu15ar465KmlpbQ6JwjUUk3sU2ta6l2qez+R2c88yEab2FyaHoe+N7cHw5Kj
cIeWrbegIj5gv4dxdWgj4y2az9d5aRUYcHLjClZm+HTOjquNyYllZkFkJvdq4Sir
XhuoT1zAR5COhVTgPvri5iZnbFJVNnlKxUUsC4UHinGNS6CnARa3prOGOjEXIg2s
1Ede+EbD2Lsq5L6rElYeQu8gQnZF1THMBHMSqCIsYnKAwAKrqbBn9msFsK8KbE8c
2swazRZ+GHpPKEFwTor/NUyhUt6gVD5asXeoE0/8pTLbTRZZZSUi/rGHJQ+hVdnX
HR/iTdE5qSLEuMlh1IcptuW7+akT/YbsAUKXUiDhqQy3YKfxlpG+ur/qM4S6nlqz
eCleehqwp452bNGEhi0nu8p67F3EwbWFJWGYsb5n58EOwrolqGJUPwdb5BBanhAg
9uqSgUzo6nlVxWDYKTMOkNW7WaTO5fMIANuHHtPLe63r8ybkpCrrmimQjY8B+Ztr
fpFPW1Gu+fcXvyGuyBS0tMPsx4tFENdFyBGjzYkhH6A4a93rf/oArawuPAmlUkOB
4m7KVRfsSZtgjHeOwU8aa+B7acH65RSOhe+T4khXpHvkmkMXBEMOCEJtb8x2nK5h
o/6tYVDdgCswfErS+xvo7b30xErCnnRmUrXooA12rru8yNcXf8ydPZStNFIummTH
FLaOOu45DHhjtmYE3W2+wrC3GgXKrylCRbdvDRrY69xckklmcBjLTmrbbKzUTfIa
ZVWYs8Kxo2X/l3M3g0c4aLNKnemkqwN6VrVrDZoaXskjqXjPOwg6VEe/dzb8qM3q
Ioz0uvts2MArJSBJt5E7lrrgWMimgP2XtZQjwVpnJHA=
`protect END_PROTECTED
