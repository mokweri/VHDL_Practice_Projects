`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iOy6Sdn6puFFl25GINmSupHZp6OTm/xBhFrbB+5B98dKfnApp/022F/ynwuFyn30
UaiLKHUBZxb6Qif/93zcHRD6P8QjSiqOu5hsTSo1ZczHw+Cs6tO8wtQUdGIR2q0I
8wrtnhhqOt85yoFuPuZEFUcRvxdtc7SuT5k+Bpsn40WocqJbFhuXyorQrpc1Yy05
atVPBPYW1Gv1dcLggA/klJvOoS+l5IBIfA+nYjfIOfR5CFjzeZQvcXEjdIqlxMv9
FKO0RHrQhEGl2i5WP7ritulQyTKUeeLZulP4u8/rbv0vQODS+HQLM+CGm7pETwl7
Icl+OpIaK6nA1r3wGrYeiWaILzH/s7kLiOwfNLECHqrk+jr41zK89hUSqwHYGN4s
LAqnrckYEpvwGbYHxMrU73gKdlpni2ypKwDm8J+C2SnYKWX3usOusuXP5PGTfq+c
4KdDWKIlNd0q6UckCfslpOSXp/ADBZGybbjXeMpvg3AhDtWvC6ASmC7W0lSDLLpe
1ifCauDQ4ywcQNWrfk4pndG2CHJ/XYRXx0iCWq8+NzAS9UAO1d2hatiXvqEDez21
1Zg4UdKu1DqOmWPrfj0pCdnMDJRH+1xgTksYF1FffQgnlSx3CLzMNXGqeyS88p4Y
jfTyYGTJni0e5eeoXG41leBnh6/QGDMiCGafcyp2DxxooJjhf1o+JvZOkFD4jTtx
sAD9vW4IZ4FQDzvur18xhM2YcEDirbChq5JCjg0gEZjJr0EOWSJLn/yKj//KrUo0
QP/O0l+FgmC0UV889Py3o8jU28qftPoFGiKKDO4cq10lmTI3sSzfYv7Mj+PQHup+
o01firhYvWSPolcYTBNCyKlvMuEXW0HyY944SYPtbRCtEZufFvLso2tbOL51sQJf
tY+JxS3Q6i+ujtsNpeKSN9gKS16m6wPBuW2rv6n/0qOI5ITNfsV98kr7SM9OpTf0
36HOJfAeLZOo2xaU93OZiFRi8uze2Ux1/zNG0umcoCQJMqtx3e0JLq/+sEhmN9wu
MPqk1U5eFaAGu6aXwA8+NEYrhvU1iJnYiCuhqW+wh9n2h12sWjicQUavBq/ENNUF
UXBbObidAKQpzYqsP/9DTvK46eeqfY9ZlzTmsm2cqXmGvm+OiCIbZqhP7IN6G2FQ
BN2MNx/u7gJ7r3BkizL5C+eGRF53qa60syU1WNfIxGzyu5hpSKckP/3vgyja741i
9Vib1j35P1a/fIu2nsEIGTnvuZwM5bWGiX68IRSpNch4ARDJGJjZPn4+uYIuVG5d
LJCI+xkDFcFCfhUp+8rSc0mzgGspnZQ/uxdceK1K9wDlR2L4E37lXZDv7sbt6A3Y
5BHB37zlEQDxdH8bYBu+LizYVViL4l7yE89nyW5L4dQuttCXHTkQcTL1U2SEL+7H
KmpcWmf1m8C7AAD/s/aY53oD/FdxXbDh4qJehmll3mJsCFhKlnQtSQEwKhFnaBze
sZmkV88fRItvd5Ef/6vYwi7zOuid53YJXZfWKmm7EXSlsEZPZ4WE34V8gpYogquR
z8VB9efi1o9MOR7l5c6zMgNnqRUN/lVm34J2nRXMMNnZH1bN4/hKC5NXSfhWnkES
gByHTcKj7WkXaTQpQcBubv6jlLWD+RAva8qTev9vSOTDNfwpZOYTR40QkW153qxo
EPEZyNTqB2QnaDK1U7essnG0jqABfvgy48PXsvxx/Q/Xj1W2CpkebNGHgVclUin0
7nOqb2810+KW18N1SGpKRzVmO5hEFn7UFHeDGpscrTU8DNTneXnzbYd5VdLul+V5
a4d/4ChsChimGgtg+6PeTc+g3dMAhqadPkYghhKMXuQdvsf6IqQ9Qi54luXnKEcl
LqmVp130LhXDVDTUnR1deJ1GlysPmjJDYta6DqF7P/rLrqdL4I25TFFDdY/2Fdkr
lZIoIwtWpO4hEzM42BhcmU/NPMo+Af1mIXmZAcduYHPRe4ReiovDH69NVxYdVKJK
NtUjdWOSZHp/4x41Y28FUEjsif9c8csLtdpXOndWpn4ldPvNIXQOsH9yeLUm1LJY
YTLOWYSJXJovrI5uyFQLhEykj7Z6IyEhPb5GWmHsBJ70tblmJg6cTm/9/9mkFNqt
e8xNnqXl9X1VK5zo335aXDY267VJgChM2zsMzLnZJMqqKaBHbhd36YVZapEapQCo
Rv1Vpu6mvMe/69GVgfCZusYKBh60XHZBs07omWHd95TeaR5rIOq5X5hMYnF4YrQ1
LbeZfVN1UxaOQnMQ9KzjKFGwUVbnKhgA8iM8nqgxQ72NCLWfKGXt0fCCop5Ut59a
fozg98UZqbge9Xi/ZH3HLp1Sm24167yh+aehpGSUZbgvLx6GwnanBbTTa6keI+lt
5G+dpOCLn0TMFw6tWmg/ggyUOoSDgvC6aeAVD4f/GWc936Tm4K7chGCMvNL4+yWH
qA0EX6E/mUjN4qr9rPADFULF6iePD7S9N0CeGvSgX3CABIpb9jckccfn+ZPoRFm3
AoyVyrovKYXSQMTAjgSdwSDtKoUSDPTRPZaWVUIdItpv+ni/jFLfxyWkRJJLm/VD
NceHpORKdK2BSyeSvNb6IhbQ6Dpolbe9e8hIK9eJKZ1jYkpjbVHK4Xuo184mc4++
mOUlsojjQd/57nc5lZhdersvxGx7ACz0WTrzGhpc0SHmDZU/2onp+6s/tf+ZTShY
kWOT0fkAoq6z30UH7bdUVxXaEVMi6Ey/rXezyhUBAwKZzkKQ7SfUrWjdqzlwWEH1
MKYVmRtBUmnD9fMLzqUspRg3WCBFesbkfYqaqas3dv5TbvNkcVAcbPUtMwA4Uhe2
poWqPfxtV0STUfygzIcBTYWgxG9wmD3OiXd1v1kwgrVFlZOzAeH6hxIiELCho3SK
YYzzO3CiGMDCLxSgbZ42u7vjZKRqZySLbylfSkvadGpOanmtAlPT3I1U3mFCnMID
Xsfx1KXpqajVi1HDDBbmQOcGOfht9P+6kp3+KRcqSgRTeEelrJjrg8Fzc6YaTOUI
5p8vpKJuPNMH2K08O67bSuHPWIEooKzsW9SdoJ0fHgfc7NzloC5y14pvaQgVXeR/
Pm1ezqR6aKHyw/Jw4k5Rwa/gqVikCNV4bk1trS3qB9sn38FwzFQCHiRnLKYQ60Tm
AuB2QEjrgEj0bEXca/JXeDUBPlMB6TjTJt38VxRhnpdxm8rZ+QtsdrIMBO25+u12
ABLMIESffy4P2BOSpHATfWjg6PstOsh+g0gDJM3J85BVx+PsaVj6fT3Ot0cdM+d/
q80EuqYOY9qK5cTCOeuTMkbMsnECP+++ZflAeiRHKdAqbM8MSBAwfBE6adO1wADT
nxh2S0o+o7YG1k7RrRfjib91wD0w7SCCMCEZdQ+SSic8oSP+McCjqBNc1MEmIflv
J1VFWo3I6+bVn1hz4HQs+KS1zl7xf45XI1BON125YkdZHeCVdyYRuWxlzRp4VRW3
TYQEnOuRXzToZzBl0i/tKqmF4J9Vq1lftvnri8MWjlt8cFr6aKU/eI3pedSguSo3
evPM45rSD2WsyG/T6vMi0izJ04Qu34NFhP/lKxPxIBEEfQ3GLR4jn0a1Ru5x7EPP
pJJSNga4yTmsCRbeioDwdavcXjXpmnL5UfuMDmSedqtx0Twev/1D1WKe6DIUQ7OH
X6GEGdym3dYsiZMCBNGJ3i8S/egP8OHncl+Sm90POrJ9gKdLnmgDWzE5VQFpfCwE
DXSa5ROKcN4zFONltIHgiR8sZg/yrVbbAmAGY/KRnpnS1lL9X1AV11/JzbjQdwfj
4ZYTgLqxKdpU2G44gl2bAiq3Xptf6fs1xj+6WzYGOmMNQqmh8cKJnKLtnW0p4BNx
pS7OgUWRBdeDqLT/X1cMh/AFpq6TrWsIbA+bqlhxl4/u7itLxKoED0JoX9oqmOtx
tCjeaHC5N4r4IDdHxFUvA7UaXchoT9qFT7rDPtaqAHGYWq/fw9ndp2y0q1HpYqaO
KAO+yWYM3kza/3NGHc4I7W9pf0KcT9RuCjY5HBx4Ug0qx0L7JUKZRk9kcBNqrzRr
ZWgmFcGh7VhfLuoxYDnwvBLl/klX2W5hs0IZ+4NsCcOFVmPfNGtut5S1AUx9H9V8
HyysMET3SeO1VxehMTTHNRAJkVhKUZXvPpdGiqZvgiwEZgCf4nGXXtm9J7PjUEEO
IJWAHoSTQW/toyzplwxnK80gzvdNn8IezSBvAwc4OZJBZgUwwqw0/E6qTUkoDmVT
2/riGq51iMDNh7GNa12dysXautR/WHA0AABcrTbWGe0aEJjc+1dmR2cj3ESU6uTI
kgmWHIvgDtIaSJUW+L4ProARs17CLjJ1kAXfEcghv6wOmU06926l7+itDpsEXBrY
DVmnkN4+C+oXgy+aZAIzffbJbS1mcwdtnsh68UwwM7PChym1WSLHrXtmwrvNsRL4
njjwXdZ5WU68tTPLPgwgjsJ6WLO2/BB2fXg/yjbpHeQIk0nOf70HrdLvsKSCY9EN
FNYwOEYYLuzn8RZm61mJfwEMKWYUMknCnH8q21Y+Vaw0BW5fS/35xFdQMPInkyzs
715M8L6frZIzi2WVa671acOlXqRLGb58PvfOjv3IPrjgvHXQYo9snDocvyH6l++L
gCYrtkFlGvJqt5TpYh0Ay1H67dexSstx4rYOxWuJOgsdefZl8kd9lPTYFn15OjR6
BRyYNC0aBx3dURrUDo3RUh/3slcfZxfR+NqMkpLQXXJjKfhLWoAZHk3jKFF0BnzM
6TnNCEyoGL93KCX/ki7R6JJe5ApXSX3zOryVFRo4lqn/3EE0ssSqZzovn1e4qHIY
O0TxnBZWWxmneWz4EFRx0YTW9DIPENELNH6tViOroVKNbytu2m9/dPhKm8IWKOCE
jZhe8UFK+28lVB3vqnGg4pV+Qf7mREk4lPItXal/d/SsoR30by8sHfE96pHVBJsd
CgoDcA/PAy1pJkT3MMq+608reHg1U+0jrUP3HqrK9he0HalcR6E23H/9I1jgW+Yc
u3smytmdBqeIWLPSpYZPQ3bh+363Pt0Duud8UDFkjbUPMhhjCyesQeeAnCpkXArc
8YRIN9VgXfGs6OYNUn0bt7OZT3BBGXBd/Nx8C6LI5JvmERok1Xc7Lu4a5xupYFCs
1c8XgUnNwaEWWKY+ARcIrx3xXybszxrRz24KQoBCYDmYZmbR60RiS5Qrp0NJqKE1
7VQn9sjMpUGOJURoR7xMvKIALieLrCdO2++Cgloq3CAWN3+k8HjEik1NbSIiK8BM
u9F8nf7yhxVmA8YdUatmZrkQpCzytnyyAj8bcw+XZIVAqmchoPmwOa5Amnw3Wk7T
oPHormrjw59ZRWDlbcnlEw4w7Lnip3+FIz3T2NmDB0F2J7pjQ6MWypHyPG8+p8uq
7KGI4ZmdaBF9DPfarZsU0eYKQSwR+6CSmLFLr/0tp5Mq8O7HI8yN5HFZJOBdQ7cV
zTiP7enuuDwkpZHwJUazQWykP8JxNKHZn3Tga63jN9CFDf6UIv/f8Zh4pjEt9Qbm
FivbH5j4BAOTc1ZURUbab3uaMawZ8mQm6Xo7B4ps2tgLcCFCmUWGwce+EuON0qVU
ip8BGTq50WT9IZX8VA5cnf/BDyPbIhmMEB7ao+4JImbbwp3y+C4FowAo+0Booy5T
am0j4smBrg24Jwt264qc9X40SHnVxWSH4DPrQhnKViWf6arrxyiH20oL31R+jHKP
W2XQRoC3UW4ofoJZh+dfo4h+Y/DYfayGadPS5rysV5m4ylNS4dlldXWx9B50vEsT
x+CPYMUXEG3DGOrJpiCAEWYqgDGYzjrROfeFNNaN3HGvbUm9IWdlG3ZmbR3Q5z2a
Src8EHOBmNtnzYkMKgfng074scVYBs65SRIp2RGwk1fOCQYrLyZzpm2mUGUo3RRP
dSUmrRzU3YbhFNoOhSiJSaYnWma2V5CE4w7CpgwpvV4Jd7TUiWA4cTAs4P81fZZL
/ZEeyRYwisCn+SuFVh2RV63+2cyv4dXAIdSsPB743fbWzBScRGCBrLM4UYTvNUz2
gBQtKNjFJxVZOsMaf4jheS3F91RhMzit8ERdOFrEaGuXdoTZKryWp/VkKBsl74VU
iIAPaZHAsAY4TG2EUQNimrWtcV+mnMv2ROXTEigCHkMGF32VW6Ik8FCI7z3/Eh3l
grXi+3N830lRQWFlZyYjiZzF0Q9d5DT/+xSLLRoJ4o0JntUN7Qa35Mb8Po1Xt6Gn
LvVd3VsQUYUK1lJ5gDq6lHHwbAqPRJICHFxfzxHb7BVklghHS/xDKYVVAAf+ngwt
PL6Vq15Zk9g4bts89bkHoKYafnuy3ycSHbRzPlPRoWZaVH+zzhucqfesmKTT8nEf
uoej8S2jqiNEOYQ3UEbyRzY8HCMsa9mzZmMfXHK0/vrukqJewRNJeHBXvyct3Uo1
7M1d75DzpZtX4KXRzqBfUhGcI9jYukDnjdBQEGaobRqvsn1h5v2VI1rdogGRR4dk
rK07pU4NOUdW/6kLMRh0yL68IvCzcQQE3URvhwCAadGKaVZxtiCl0AFWXb/wpJqR
g7Kj+iSbA1yb3U7UIIu02ASEW3XJiUwChhPAiHpKOTSMPhNq7cY5ZESCVsXZcB5m
ZYFJXVoKHLc/r6XesvsW7MFm6UsYdjQlf043hnbD/sjfxXiucSMe5HGNieLygmlU
ufhrj+ynT1zbkSUuloCnmNZ99PWNlx1jM/1DkxEXhKT4CXYbaR54jvA9rQsP3yVz
7hFNvKqeMEZ1zvK4HRannn0WyiHbzekPlE/7LiunRHbxzQtZ6BbeTms9bQ/NPbAJ
l5djKtkjr4TvQCH5O6vgdl+7EA4ZV1OKWh6CoMIa2YqYbzynAusBBnI1J+/YOYi+
2Uz3w9XIYx0wMQg2TxhLxL3SA8yMVrK3Bhb3A8aWYdl1SRi/lMNiw6OjJose5G9k
ymQrGUG6XlMIhmxKPa/Q5UY0r88VZNABIIB642gKl2ZPvnQcWtqP9RAxXGeDglrf
zqxtiyjfM6dujcrNzOZt2ibZBzYPRwYkxaofHliUSZkEkKvlfa1WEd2h41g6W1Mi
7go3305PuhIOQw4ecWarmyofJkWuiL6FHThfIKdGpTJqpWRwWUXG1yWQbzw2yuuT
SI+gg0nF/pGrDaWO8BxwVQobJeWIMVe5V8J1xDb5tBHmnfx+A6TYmd5pr2UR0eys
UCPiwTO39WuD2u7E0JmGFepIjkp4x8nXIrP6/Z1NN1on9Ff7UbQVU/4hDHjsYjXD
jl5iBRRx9Hf1CP3lsUNlfaXtL6I9DML0jXrKxYDmhyP7xr0kxwUrs+0yTjJ8Gjnt
Q/a8JckXBs6hwncpEbtE4Yb7phPQQlbJ7kIveLlBgLFv1Rb5oCcbLUfUlMhW7wGe
zn0nsMD2mf7yQF+yr8d//hJnpPNgX2I9Ks/2lDn+MZM1+8t2kezCICOMxykKUMHT
oZ5DLrV7WF/7ob1oysAL9yHFUs/5Qs6EBgTCX9Cv1U6NeXjf4gQT1YmzVL4xOQ8G
Yle5x4YhqDTEpjFSAdFyvpAfQbFNNpM7L7XchpQmKtsi3evYdRbxgdJlEDZIZ+Dp
lioaRMP50fsREVGF6E/E7t8jstc20GW9AdByV4p/KTSgp2nLqRdO9FV+x8X8NuDD
iwqpTrYC9I63FXESc4T/85qE/n4IhUrTuha+axwnzdBXdvnJrbH7e4WnvEEP3jM5
yrToNHOf3nikCB2WBw5TsDfHDBR0j7q9oh6lYQKIGjzJp0pLuUvmccL7qYJgu/i0
JFq/hgvdAl7WN/01Rae+kusgQ6qSlPw4/l6ea98BeK93mHk9BjVOT/WKM53OG9qv
+S6jBhXoAR80OW5+mO6eQuGSg2P6FkHK+b2LmdYtr8XSDe/GyEwqaBP8VrI7AQKx
xciCL+h3XtQ9JfS0nxfofIHQ5xyXJyMUBJFFBglpWDaUVGGkNCejoz9kvBnvLVlE
t6FNHrEj+nWAzGpxMftKx++pdR1scrPb3SitrriLYST3yCzLcJTRrcIAh0SyRFR1
ZBbPUOmK4Q2uiZ3dXWFEUaZc02xy7eSW7ECSZ/kBZmaR4ty5vBYoZN2ngNeGtApA
8EnoRzItEphnBpUnaNcN3FXqvuhLfDI7XfQW9VeCmdnd9SX89o59yB6aCt5EydID
wHHG5xUWpuZfYIfhcN2dkbIF3OD/4yDHM/6QPU4HYjTKd/2zRam5I3OrT0mnb9c1
kBuD03PV+N81cu3gg+8cZtj99b0ngLM1ax+NIimcwxa0RD9NFOwnm4p0pMuJQJsd
Pk2L45yhFhG+xKu93QDPJ7Glp+ycYp+WuVs4ockdR4x88pPbIVHFC1soKuu67kmq
5xBq4MU2IumPG3AMNLWd+l4gxzv8JkYsE9KiHSpumxi1teYbAnMUitS+f4P2u6r3
Zbed3RFdSGJ+8jLsyUGsSSBUnP3I57IcKKHY3dpqHjrtiUi9hq3nGcyLqnJyOCnS
89+0K/tZn5R99p5CAwwB2nstoPqCtOfnZj6Gw42omQKjD/n+WuGhaqQ/Ucm/XpjI
vWG30iKhu2UsCExmzAttvXMtaenjlu8kV4Y3IUOU62dSd2koRVMw2pPZfzy6k3oM
rcQh6i9x1OYU/N/dmmPxKVDstehrdLs8TrWtKuEzWxYZ2auzXTpxmcofFhfOtRfW
m6uZCPiUT7axDwtiPM+jca+1YB10HQOT9sm2gszEoBdh+9mScRBelYAxDv/s0GgV
tP13mF1RGACymGXaI4He+JIUZ1jBrrCZkoDzHwvQROh223yLy7CMlr3kzY8Ultam
a+J32WAoBJq4uC8MDqjDdMvhcR3g7eeRaTzPkSubV1Hxmt1J0nW5qZTqmDDdrDNk
KniOPfKmLD/xzUAx4Z1XLcEkiYbWv/0T/4eHad3dKGcD1eT/70r+87odX+R59+zD
njPrSblBLIVMNBOY/ZpljiwXfDffrck8lmb3QxWouGOyubkrUsvGVOB5ZDCVeTcQ
/7Cz121+xlDBB/2l7NV+986sA4RF+IOSlYlBPeGSAJHtr+sBT/wQzNMWe9pCdFgI
dxv0C537QJtLHI90+T6WCy9do5BDnzfpee4iH9j768H1eXUMxCuicgweyj1g8PjF
62HqEOl8Ec/Js69z/gJeijFyJ2FfzX4GZvhzAut77Xl1DlVuRSv/SMeoSNEOpYOd
wzndjtw1O67kUu03zuktreZ4jvrtKZgVLgW+UlPDzA4L/Ct7GMDwquROMV5tYsYX
1p5iSG8s0kRSgCS9tNzxpztKvu5vqCIdaU0X3kM1w8vGZSC1ZGvohvqu4aBHDFbo
ccsqJJYGlkKiF9Q80LWCAIsrdtdzvsNGqYqJ175Q/w1m8jpuf0KVfVx+pWl0bjYj
cCcRiRv3rF6ULDvTb3j2f8S9VuXM+ngLNOYiNMKhKiQhKzOYwZenu6fYCM/i8mP4
J89KGunlbT6gppsMoC0CU332zSq3PEMmY6hGglbJO59TiyP/ZrJ/vmC5wZi8/gOO
5OeOU2PtuTDj3I0RCafZdqTC0qcXEv9bmdFKMFwA7Owx7VXnIHaVEazbdUDB7Pi5
NQxUWXLpBDb2fnNxGcrJA4pWAfXDs0ZsRMNJkAGvVerRwWov6QHhwvXCQuTTc15U
ONJCPPus9K0X1B3Zwc0cI07Vrn2i2vxBZqcbHxFGHc2Vn1+hdNAiqeIcdDJkVgWn
5sBhN9M2Gwh7bViShYTFcEH5eN0JV5qiR0rHAut4CrWKLteGG9P20JZQ3CJxYk07
yBFCptZ1ds+7dhaHAQdHsFPX+gfHUl3yIlakizSIBF7Oo5b3ErDSziQ/3GZXUtuo
3gv72tAgRWiOnULS06CGpqRawNcs5eLgtBvbcHz4cNsHDcv6bVyIyawLMGw8KNrc
UZkZaHi1jDXnQHQSctDwYnSTnC0GfXFJa67YAMRcnof635Un46ffAdNVxzoEOcaq
XrbOSuV2KMv1hIksNXYstnykpwhUo42idZBTwlVDHZawjy1ujdubi2K1tqa9ro88
HIHiifaJTX+Laaw7GuhzSRjtfwYxsdp1gDnbAEvc5jPoJZtEBCWqgl3o84IvuePI
pf3GT1kZrpiXSYvNZPc2KR3WViw2aSWWL6BqTv1b4TF450tgJEcpqVa9vktCQ293
Zz1XW6CxRmQyI/lFn94Y8KXFtwXCpHPQ3+ZEQPUB+3Gk48zsX1zjulZrSli+g6kq
BH3B3paLxu2uUSeFLTgwBMT+IVYIucbzRZNzFgtMjpJoQCHXwKJjgEjJbXPMKzgi
ovb+MsTDDOA8bOJXPAGP7clIM4R9fs3ZoGzsodMvsoziWdLx8wSFr1khwRmGLODM
NNTu/vKUFPnyGsRuovZB3VqMzmTPLLdZ4QWbEaMWhFOsmdk+urZDOlNHBS1B14uz
7CbsqyktSxpzh540NH2j6CuMuzH9n8DUdzZ6Ozi2WcbiV4Joh8T4SP7IVhM54CVS
3/F++JMHdzRZeSw/4EvM4flENaMn4f8UDutYBB2+DtoNGGxCbJhdYVQET1CTj3KX
cZhahYq+pyRbBrZ3oypQ548u8TCNAeyX/5VtmtUiBQ3kbVpGggtAZ3mLuwTbCn79
ruPlRwh3wqYc+2oojbLKyk7JG2AwLpCaS1TG2VuKdPRIfRTuJrned9cJz+uMnXeQ
fcBpwMPh5TTANM+h5R3re49TSup0pq4Z597/CzQcJI1GHA562p6Z7GhpnW1gl7eh
rCtIGg/fEUToJnYNYDWRVw3lvsIk96EMIDjhyMr18iAQm+konphBWkxUjdRD6tWe
QP3HTymXOrlGY+oJ5eGbiWlJQUBYSCAx4aBn6WXZ9jRnMcOpQ40XUlmAHWNufw6f
rZ8DkAHXADHta+n5YzG+xSwObyyUl+zAuog1ayVbTORGvdkSZT/AXO2akROFthXg
bWfkTU/jtfleIq08d/YIbkHn6FkgLDYq8W0qmIBShjmNOjz5FB24SquUYxeHVASn
JcWKYGAKlas9tocAUPPSRSm4Tl+JLNYH6i3U/cyxsmhY7bD3GWnLtB+DPmxfmqMG
CP/LFHyuzLGRqZ9pBsDvP6hmlyyC8QqV+erci7F0RZ+uhRWjIWQaTNG9F4stFhaR
gg20icD++ZBRBvf0u/w+fB7pl2ppu1avmaHQy3TZcVXgI49735zfCdF46oPuTVeK
K9moWbpG26OVT7FZ4+oyZOfqGyG4ZXJtN4BaqLICHQCqrato3EDWK+71H0JP5uTA
hR7W//Fyk5cLg+FA2nj4TG2l62GY/oGfiV2gIRTji0SW0l4L5ophJLv1kr6B+qya
LdCkqyruxWWe3y+K8kBQOPPEzMIUj2SvSY6yczckcUXcylL4BnRd8JqrpKUBqOV4
Nh5S7j4se72AeDILyj71px7178DZf1DP2G1Jb54Ug+P2CnzkMRvgqlCG7wpXSH+H
rfaUjbuTrQVjkKL2AhY6G9Wg4k1ZeOy2cEXF2gQAxpeO1rXJeBw85V+M43Ky2xNp
64jM0OlZcCD1vsXeb0Tb003YYvj0bsCJ5fJaixyZoCvMy3cQdmnkHEj6JXaTXx4e
esTx2Gh/dVw188QqgIw6Yz40EHQkzRUppY0MMq52nYsAK0cGdDsmrh0j0nqufL0a
sJP3oFKwr84Ek8Um4H2a9l6eABCeEQ7pkqaHC/f9Sw8CabI5r69LjEDaDGPUlyrL
O9QDuEMVu6AIzAA6Cyfpm0a9K5I+2Eb8mbZmxaFb5mA46KeQt4pfkA/K+UD56ADp
+ls64dnlZANrVoUcV5Xem4pMKdEthTmqdyDYkaVDHS+/Hy8Ij/Pgnl0b+aOQsKbR
IuNkJQ0+jm0p6eOws/FB2wnkRf+HPSPOQG2t4oyOykxdl4QikOhquuSxSM6UBcs/
sqXltpcdnkM/tJjC81vDFI3enqxsQ8BdgdeOhTz0cKVbGGNzE47tVhNkj2ybl/9R
y6j8IJ0WSemrh01arhNhwGua01lfcPWqckiKUaHqbI6tq3DzlI3Nb991ibh1urd4
LvOT1NGeFNQDVYWE7lqRDnNM8p34XbHyZZx67Ik92jaCjb0lKh6JY+kW/hWukmOm
dHEMfgv7N1R3UvFfgIEY+QlxHgsFNhveSPN6its+q9PF0kY9a58g28NXfU4F3Jt/
PZoc6m6/pr4tC5mpNnjPaRmlik07LINo9SRRGhth2tFzIEG3c9pAvfegYtv5fnoz
S0rQ+fCYhhDpYEnOYfN1IuRTI63/CgqPz59iyFcZao0Mew0DTIjxPFyHs4ItfDfy
0RS8dhk3xcnkQgJNeY5mIptp4xCvo2BfYH+GcgqurJOL46REsfpoMkzNXietWNnX
NA+fwmYAArXCjtqCgSRCBHh7KQkYb09WgJ3DMSJzU9bVvUDSrmVz/wLtVcRyMz5z
9WCW5EWepPE1AyOfuvH6gLr26KFJib9S8/jMW23O0T1fGMEDRLx1Aive/IuzLCef
qR3110qPRDNwsrMimlWvcQycCSbIXaDIq535Qki9b5YRk8l73K5r5K31WjOE7kjo
eR+XZjtIiEncvl9MbZNoEl1T+c8VbsQVbywbmnWW7F9bDJKn26pQzRv7QHw8PkoF
JMef+pPqZYbXd441obVToATqcyl95qIQpfve/nbvCa2qZpnHiMA199T5kDNGS5Vi
k7PCLS1/1Qy4b9ScOSumQaRDY5sAqISmlMqqM2ZgvfL5paGCINh5oUqiRcQbpJqw
Dg/aDLvJ/yRYC0XzH+yNvZ0V4PH38w8ofL0caUh+IhnfzZEkgOlm+bvprIlIKUif
yLp6hB6mK4dH1PDjBRBXIR+dFZuLxia1VN8n+E1/ADifntUcoShTBGpCU7PtBCBe
l1PUyc7hKzRZBPaXUXmxCBd8WDoBmH55ujQYp3crU7UAu1sWVuXPFgPU90/Woapn
PR8+lCMCOHY72w2sgCSdDb5DeywIBcpVwFgoVzWk/GpTy5K4al3V2EIsEsRYdcey
2OhzyV+w9UDfKbXDXtQy8uyoSvuyZ+r5B/WKBTLXGgLYQXb9RIbixtI1oBw8L9LW
36c6J//N+IaNwJ9Y+a0CYpW81fZj5hV9u8d8qCfqcuqaN5xodmmZ9wEEbcqi1zBZ
VeeQ/jIgoILego5lAEdq8crrg9XxYgafIqqVsXJ6n4MD+EkJrDKkDvPSkXshUm3A
y9b6FWnHVQqapQ+jZfgrFmzMLzjQgiNyo9CnKm409x+8U+aaI5Kc3hYkhdCy4r8b
XWsNUQ2u4ZqYme1248QZbiQTXblv20klUAdxvQy4K64=
`protect END_PROTECTED
