`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgfy67xhTelBh4qbFX/Zqt0IjFI/NnsuuhKOyKZC6+Xqg4UrnMlW8S1YaPWiIYRr
3YawRXriEDSWCbkQteoDN2Y58qDgo3y6mUq6y9yqnl+AYPPADPrJEA0DPn1SwpaC
vvNEMmPws2aA6jnm8gOVG7yaN0tMpL/1CZxF+Jv0lmjzzBdSPV/PjqVL4m/dUtnL
85HVgwKG8h52XzjMjD0R00jXV4o/bp0LG68nlnUbWWScCsnvlNwe9iOnqGpHO5/G
38zPUPNPxMmnqDB4xx6BYiopxYgYp6mvvfU2v1SnZcBnFLOm+2PQG9bvxspOcUm+
ET4vZG0YavANXQJvUyx8kh/bzk/wRdOb35eaWo8VgA8ZTeS+iR3HXr8fAS4apfWh
rV9/TBai8k+Dc44480yRQR38pWE7lCZs2MVsJSIDQK+wQgTQvaYj7b73MgVmoY4x
5uETew2hEoynNbh5a0R1BAmYuzIXSxXhgWFafrsYIDIR16XNp+g/QjbkazzDWS5/
knIcLJ2GWlo2sKDxdZfZGpvYGA7nUUws1sWayfA8DVZV2SoO2nSYajyLtnpRWwQZ
2mSa9RDUMr5r6JQu1b7scrvar0Gkq8g+qzsjNm1DrepeyRU8EcxIzWah5lfQI7JZ
Ij7Q6Jil8sNEaXCFkf3bmYe1mectTKDbvxyLI0BdMLm2FRDeMwOngfV0zgs8goMK
g/QbR7sHrGUspBG7mL+kvRVPtnW7vhx5/vMNOrk7122dz3yxsNqbXTmoJAYywJVk
wl5Zipvv8Sz4aohm2CHE64umYH+oVMD4t39d2r1dHNekuny1wlfuuX8KZS0nvuFh
LlMpKRCYCmjeiJZJKTF+qPGa8NWgaPW8JYCUxVVRw5J9HlrdQsqsIa4Bw7LnuUyl
UFm+8DJmbLz6wz6JZNiy8N4VOJ3Xl9L903zMlzaFV9lrqPPaBXu0J1oA25sQv+0n
TxEUbFzhk4ycQS3VIbTz46QqgQsfBUiREb29rHk7iJAypfVXZtlFTsarXmOMfV6C
n6xqUOLFH4g5qr9N/iljWfvVrOHe/lao/DUCdlO/c3Jt7pdABRyV1/NJ+7J8CDcZ
s5YizTR8IahkqLPZiRc3xm25WdUB+jq5KmGa326f6ZRfrYJ1E8sNN0zn9LBdE/2K
+A7KYU5aFbsN3L7aOR+6upOJsiHNH7CvwdtmKaaQLImkH3Hj0a6xg1K5ToWg8bX8
wbwaMKJvo72hqydBVMSxhBhkMkzhgFM3Pe3ETKjnqOLOVCFQRkC2weKTYOrkGFOM
MsO+Kn1HF9MheE+oXxZii9DokGeXL2UPnPAE+1EKWKsKf2tHLEa21lR7CCTQi2vp
FVOf1Q8vBIz/fBW4Qf4+GY+gfjj7FBF2fDthZJp+e5EV2X5i+tzSELi83/NW0OW+
+KIs8dMrGQsgsUdTrIyOi87Q/NyHiwRALGoje8MiwROtABV1RbFKa8LwV69CeehQ
HCDU+FDXkhQEaYOKEmUHNZa3ztBHNaYXVMiYMIR8gLLxf0nrCmyO8R9u/al7y4bD
R/k90gox1YKlEWbXo2RUCZL9rBvxdCH00wLFmjV6qV+H0nQ3uq7Kz2fP+5+ppR/S
D2IlAklc7II/uPVWVo4RCW6ReZo476cSZ0nGGCeATdoiYlrp/yquCQ6g6eIFj9TS
EoTe19GaW0LX3REinFYhFHvETg19+PJgVb0ZLsYsbwmPKbpEo2ArK/E6w+dZrgyN
yqvDJfjF4dAYGgwStsaaJNDQJ0N4KHBGJB3mABUpmIjkxH0LArZxm6dhM0ogNcpZ
deurQM7Elog/+qQP1JqckX4Ztzz5rXble5vqyhdXD/i8vGJu97nKnBSpd5hfzQez
u2nLaOpuzesbSKfRk2ZLJ/Ae/v98Czvsc5fesOSh9SHXQJ2BzN33flX1A3eoJm8Z
k1MPPA2oruHkSn2m9XekEHxIm/7lXy9Mgiq0f8YbFEQHXoiai3n5zoqmJ7upHnD4
QmdOsdYQp47aWO2VrmUVWsEPKlQdE6nLV3Qgoavyuw0tajvjH24WB55fhm0Ycx26
v+SQxOflLn0uzOnzThCdH1BdnG//xhptIvrfh9TEbGjU/THOw4ZAv0Hr8FkdLDsO
Jqb09AKL2p0iXUlUmNQVsSnNt88YzYsJYviRRTsSp96cppOp0K6kQmEbaR3fqK3q
hBFz6XJaY1qrFHu6ZX2TIjovu9idTXf3XJQumrBKhOMr64GsdWPwb6oOqBw6pISp
yZlwmE1a3PQ+HUGcDOO7GyPD74qz9b4ONEICTFZ0XH7QGsEetshpaVnJ7ZdVsAJJ
8g630+vu9ulkbYsTcuuE8oCxDMu0atGfmbTEY6JFxsnzXPB6gvar/8EZvYAOmbGL
QzoCX7aTSbciK9pY+VB+hHi2koqtql5BfiAuMbCQVqhpEtFmisgabdMQEa9HMVZU
xdaamfb/sHbgpIgiiTplArgGfTGgq9lJdVdC0a53f7rQxEskBopzxmg2BI42QcIO
jXS9e6JifsXhaAtoaOD7ZcxFfEnZUtaIwtQiP49qXtmiOvrn1i/NuMkhkAblyDny
uJTSD2lWpH+bMwMtR+Ea0I598kNObUXWEGqWostJq5JM0iBD424TWCfzsB4XCstF
ZOiBDoEb1LCRFMlvHT2HvLfGOunwooG1ipwUAFCQjyAsKfbIGxFTrBDrfWqmbXFO
Od4OvzqfuP65DDc7oyeAO7PKPGuqlrvhXbbyXjRVT6UDvY1gj0Bx272lWcjaA53b
YC4ANkDANBrpJauYcFZ9yEupWHUyk/sCe1cuXFvupMF70BffEjsJQ3rRzWF9/5nD
PdhDFZOwQ7w/IfTQ/ozsZpPgkVt/vwXDHT3a7FoZnZ4FN1/++A5Pxs3Tew5v5EX2
11qsc5rtd75blg1JykLiGXeGWQrLdBGxPLOQMnsshoCdA8uuIeoYcCrqg4u1+4te
n9l1tB4/e1C5UQzj5M553UaZOKRTTpSt52PHjqwwL1HzxNfZ6wDfe0JVJs2gvx/3
tRCheOzyPSQGUJzriWKcolhVrJEGblyruvzceKNVfEGqrClDGmP14sg7ZORN6DvG
fuGZmFX8UiF3i0bfXNojeb3oNZGZoJBxfzDjM+99jlnh6Qj2dujR8x2Rq71A0f7r
2h2jdIwixSu31RBf7lqnkRfHkCAPrqpcXHiYknPN8OQLrK9M5fcHRVHc/uvY8/Kr
QqfTW+Vq+ZQtb7jE+dS/OaOzrtiysJuV/y3cgeJ8ioYpuVmv7XDch3DAdSCBaWh9
coz3TBiP+/mlsB1TzaLma+8TfU2I7tQ/J6iw3DcqLkC69+26CsJj35q7axZRxW3K
`protect END_PROTECTED
