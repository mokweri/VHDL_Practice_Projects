`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbzkgWQRU3xU5l5Zs2WoIT+vSyjIkqqHyN52+zbw7gVxkbPlD9i2errChspYjB9v
ucJ3U0Hb8bo+XIGQeHjzk2C3LnVDfHzOoabWuU0xHpyXHx6zV4KAYC/R/9ymaqAt
zIwPndQ21ZURiEM1T4XhOyx0VoflTEODe7sJIqYiQCZswQqaXJedkukG/Y9JqgMD
HXTh+Upe116+wAsTQNDHhdSDhoVBJAeS4TLvgL2G4I3WMHrnXFozz8LAKQiVhnja
w0pxm1RThjvokyrpRlAdMZXOO8YTzMI4oqN6/IAods6XkD6VA3cO6wjnW1f3DqP5
el4eY/zmDqzsiA/2nN/nE6VzVQOSeyt0Y83fy3LpzPYfEkdyohHJxIiBW+62YfkK
cjVdR7kUg9w+l0dppIOqcAj5WfcdrCY6AakcTm0jmRaPTc7/po5gK5A+K897Alwl
qhxxWlVmogNjj7n3KNfPxV7sqpiQtOZh3bf/K4kyPQTb+wM/W02Z2g/hvDCD+/8t
csD9nzv9Ye3io23AvXXDcFbjDUhLsWryvYWHRO8oBPAdZeYrPVTkiWb2EIr3jizu
5M0ZUnvBEymcOv2uJRjDz8Ut5P/sg0v/RMStMR837eCT/ya2rTQg2UzfGI2CETys
9EKoDNXUc2pRPk8M8KSoDJwCXRDQafASw/aD9MuvSNXVatELwb/F24+uYs+Yt+DV
QMA7lm9xUbJWw7Noe1D3h9jrceLcJFYVuYhxOMGR+zUo7jP6mTErjJJ/V+z3Ud1x
MNnpxu/2Zh8kKdTSZCJzXG5oDWTrTkBpKTMjVzx/lp34wLSyuJyiHzCn1I1qND+1
6+t9a/V2wkLnBzFb6nhfM4gwjfHwr/yn0IYDnPS2+Bo=
`protect END_PROTECTED
