`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mp1slVB13KmKNEWFc5FeIfh0LXwHVBrwAN35vMDnfNDFhsK8tJwy68kuKNhs0/9n
sw8quZyxgOtfNSJnvZoTNTxuXZx8hSagAvvmY/CDiyReTk9+fkAmxKBT5gn/Ktph
MUarIIi9qX1mPozI6b4NCJ8Ho7lJv8QfMwnmefuihZym2dwnmFwQGH/QAXzl6PX1
ay9CgrAuFjQPE/wst5z1tRqAKVSDQO5DXQqDnWbTTPXgRf3X2Ezn5zYOS5pVzTnF
FpP2+OutTxiHATRxJBs3eQg+V+iwyhyJ+x+oErsNGAKtBq4wYsaM+N/azjeXah6/
YMSb8q7bEBzayQhvtDW08NWkIjJynl3NoIfi0LmbtNlyw78DfgUKFyRD9u/l8/rq
JaMtH94/diGm3YPxC7hMls/BTg1WmzaOrDv2nz2KabuleDsUmvT+AIbYIcawTtSz
M+0VEoKGrb/Cz//9xi8Iml02g93v0mZvli09jOIhfk9E76HTSCVpznmhrCuDd+pO
BFOEjuohAnGEjE7wE1I1QRXFIlLWzCMowSRj+wP5AoxFJ+tTneZ96OvKLpZ4Whm3
1RCig4DGLoTeJjq5irsGzxnXHXrCjbIv3mLnekKqqFGocRG8tnkPZXtvtVLY0CM0
X/eD/bmCktqdTYdAubfPaZ67uG45YrNzSDMta2eJuIS/nN8Qd2nz1AGRFg1hLNXa
lGz1i8YIFuKziD4yXU6F+gsKYoCxmTpjaN2Uc6upuetV5xvrhRhSNSXV48ECaJP4
IUg6frSm9m0rxHNbd6Kb7ja7MXLOFrPM5AnK8L+XKu1aVl7HIsSCJ+oHBblRnk5X
mHGAQEaQ5ioWYswpYkBjvW4Qhe1opNeww2Thz8ozEt1pKSpsT43JPnF4vwkiCaUt
mXJEzlxUIIWYD5xnuNqkWUTwB6YLomJD5STyZr9uzfZN+C3aHRxCU87Jo+3q9jw4
+naoC9ACMp55qa8wxtR2E5X158d6nLtKt6xb54O0omqVc5o+svCObRHiSi8xzLb8
8bMNKCyit9jAb44PO3UeXzFKdUFEvvmGulOGOLVZIcMYPMXQtwZRs2DKbxpi/5uG
dtBroAKvXfE6HZYx75lNqMQGvnmXbl2J4HCS+a7fGEJSqqnDz9ciyIOaoTpKBPoj
iNn9bCPGvlUBDE8YzP5nw2Y9imoK/zwBjymmA3Ou0wvHjIalRZMm0GhED/VPf+uV
0scM421C8tgOVuUbYNhY7xxJk5dpwUTC1Ba3wuX6G0SA5VoQSY9vsXTg9PcHnnsH
szQXSYxC3ThnFSpPKrsNOMky2IcTz+BYka3HEqATawnk1lHZkX3z7npNBuqdGgna
Ax0Tx4BpnvDgIHu9yitIaxxZrPyygBTqycrS9gQVhnUjp88mz/8gNXJpNDGVeqpM
U+TOcEvKMPgMfTamBOEgtuz7i9UnA5A4AVScFXq08NB8hY7g+R/MeEn9uylRs4se
xKaORlHdUqsx5v/zkYiPW2JX4iNJe1f4a/y76W+ERwXasRCSgNkOwI2GwQXHoiA4
CPt67bcHXxVWs8k1sa8sSsncKmQdwD0ZfTPnssyMd8BO3EK6SnS8dPXFqbCToUJG
gcekoX+sDl1AM2MJJfhKey5avrwk3fW+Jxa9/Poq+3yLSIgK56pTeGTwdx4Pmb5X
35rjVXYMoHLqoOpTr9OKiWO9dra466sPhEFtwcbImox887DkyGG+fGTJ19x0HhNF
TNEAEXUsmmo7uLAk/SZELITWdjKclz0k5r0h8F/elJrxPPsKYl/X2kfuDkZXBBc+
Q6NpnxkVaguJqZZtI9x4kT8xupafbstPXfVou+d+unM6SGLfhxMRAR/pHjo+Wuhj
oE7WG2CnvAAuGAywmutuqp4OzqsYziafwxK/UF0eGX5ZKLGeWANO9q1poDALSk0Z
uYXWXwFYDIU0pnsO9vuBkVXrvbSHe4J6skGLvQBZ/xLQ2UDQUzizLeCLWBgoI142
IDYPZ3fxDsDacBNW7rYwYS2FcddlRE3v1WJ3RL7M3t5BxdpFTEHapPCBKqxR1XHK
KaLNxYD7QyAsV/CVsgxJlfmvhuWioHlD0YZIknZt5F3B0XjqOSb1yurEg3u340sa
eu6LmxZRj4IVivEICrEMS3tqzWUY5fKY/XDfSCOI4GQWw4gHfbKbsAl6WHidC8Ot
a6eZn3gzEg/h1tFRBfEoF7XlncuBAL0VkLPLKM6S0g05YPiiFBnHxULfZLdUM86X
LeeZ7ZmJEj57Ew0oKHEfyZ+xBjKydS4mkUGJPpMu1+VA1IVIT1/TZ4TUytr3MDvZ
kN1mDJBsVXUv6XDMVaKE8bd9G1x6+HY7cIbJvzc5JP487092Qb/YFVe5rnukvQgz
AAAyqVs4H5tfkyNOmIJSvIsqhGsNbcCyUMLOIw5xV/pwdITTZsHQIK+oBqEZrhAC
TR9eYj/8XZQRAO8BI37iJ+qfUmVI12RU4CgnA8hZg1d50X1LqIdQMj4+LNUfiVRx
+K3Y+AqAcF2gOW0erfQqKcOghqWf4zZ2GWozei1IvylI6f6m0NN36CfAOxFpZrQq
G9iANs29AyXtKcUTCpiVaQRCtBpXjqRMBzrL80HJ6N/buANPFrew68T05c3MtLH3
OxEeSMa5gmqhdBsa5sVJ9SxbxxeD2DmcrR0JIEDDjmt6bSA1PCrIDA/mDbHQ7rQL
EsSpVnriuOanmaCvvdZQpB6M5GOmzmeIBhrdluD6+JpVKgWGEcg4TMoflyRPxIPu
xW5JdrfFFbsaJko2/M5zTqbFLdVk+k7gzROJpsayVD0+yLUdn/ZSBBuxi02rbCjj
i6qx7k2vdzgfjt4le57uDZ8+PGXILZ3n9C6iYw1w3AlQdBevoJNWmBMzT+m47f6H
yjtTWp9QEOOm5zlyzhXAHVVG1zr2IMYRscdxUlZTGBHaWm9MBT3PY0cBwo/rsSxk
jP3F9JunXp+1DSbS/Mqv2AVAQFxWcqQnwNXjjd51rQWgOV9XFSxhsX1YeRatQlUz
hntpOP+wGHs9KRbszrxCvLSHZj0uAatnLACs2SVEwn8XIFTI36Po2VAhOnhFuM87
f1Jw/3XlNEjUsEo52CJnwYPnlOqlmE5Qd6St7GncbaFTHbaVn9y903LY73FKSL2O
vZLUN4LKhsBRcIGfHq/7PxMBceDGCEsuI8/fyZLOszDsU24Dw8TARcsWbBa4mtqA
OL1drjH3VLijr4C0JSHFI32Ht/iUp23MtTxJ3nY9xNhIPIkvFdoH+UlrJcs4ySo/
hSWghVlP5Ypov9mi9Jb2lkjxEaPYNoF8Sxplife9bDYO48AF9feg4XZWq/d99bDb
sOGke1E3UOC2k2L4YwjDiujjbiT7PBzwy3ARrOp3NX9IKXfSDZba4LJpYmw3I+vV
J+Nejy3BKrq5m7og9A+QvS5dxQrt3al1VbRC2UABBnKkjGXDoH6huIA61JQ888uJ
/3HZgivNb+CswtoFcKZDVYnnSADMUEv3rnurDUX9boFqlYvZvyiw/jETgGyfIWuG
grH5w75VSaB8Bys1LawSi1oTbBtZ4T3jpKBKkUXhzXIo5WqZ93WbHCXZOP4upLP7
0C1tjZkA7ddH/8UvlPRQ0Q1VbhSDMq02x3PV7JkO77tRh6Xv5/RQxq50F1ERGe7b
KFd/dtb4Wt8GeId5gUeDfYJgM48B1SKZWxPMwqgQoobk2JMv5pzmOZl/kZ3r8J+h
8viMwj67saG1TnKao7HpPziVCvqhJFyJfXVtwCqYabuO938zgi5lD6NipdCC7Yjf
FQXODxQrLhPiOZL5hqY5zBi8WU3qMtwbWxcf/xZJilJqo/cX5oZdqSXApu3P8ImT
w8TrlbqLLT32UAh/4dc5uCi89Uqqr9+Wy5yYN1CmViOxp/gaxJ00btupBYLp4OYn
0bbOa/scc9OQkfz5HHcH8NVYPh8sVjTy/gd6/CgrWbY9w+6nnTFePb/L8rhAiXqH
IpsXK/vAWzMvUXQVKeyanBwPsxbi8MQDJShRJ/BMshg9T5qrKflbo6MNbAApBnTB
k4ZwiStVGCn3/KDeHaZHxNJRgnzFCY36fYO6BUOwnpf2PsWOddwK4Daao84w+T14
oMl9vjKS0l1JMdeh4MhCMcraIwFeftA+uOMxP508/XGCtiRiwqiPerGBXsSF/O5/
vNMVCgsajO+9qErla0bwtaL9UgEECLgjqRKvkh/A6pPSGyNceTnhfzHZ+M8Mo0hT
2s2pk7B0GpYbmmGcPdKeWrgEmKt30vwoe+PD6aTSb+B+mQosmk2sTsJyd7xznq4r
q+uZze/ehU2m0pZOlA7kGk0MTXzz21nuL4ERoLPlSPtRfxGi4+Qsy1yyu62uhImW
/0qki50yssrHij9QlSbdAzicW7UO8rgBHcOEhqNOGIUYOtC2emKABwXUen8F4S8y
XSL0yhomS3FWz1qzDsaOebn3AGPLb/CjLzm1NH/1gNpp+6BrDFIuwd7t1DY7f+ez
AchE975cSs8agQ/F1sY4mOCNVN9QPP5EMIpmbIgzBlec/MOnYxiWekjjIRb367oo
AMktWmheDrLStbML2ciZVdbQFCXO9NPoAqBMOVYsGq/YuoP0wqUG5rumB1InQtVs
D22szuZp9TG3Y5/AqHuUcpSX9TW52D9zWsG4fdJx/lHZ3kdU4mEe4G77egAxKY/b
TwMyGNeEz0qJdUk+nDTmPm3FXxGqxo7SUDFE2M6+4uelc+BKgWQryPTUwGT+Cmc+
SuBEcdeyVm1IWh0l2ScyOxOvNeTdzxGSh9nVH+vuPlhSw/mE0QIYzNPqWPWjWLaT
iW8p8yECRm1eduVHRf+U7BuQ44dopOm+kCDY7I5wjqM20b2CZllxymBWedx5OCGO
kU38rBL9pYx2j+h493ePjch/iSoPwSkjzgsZXb08j3VowUCwfdeAji7atRHVtSQA
mGcQmyI2gNx43+F/uIfteZJp/VoYhVOMcjD7I3Ad4IkADLHDxMS+obRufPyDhr6i
FHLJexpExix1yZHacmjpE66EAxeHnpyrF5n/1WtI/TD4iASh7Pk9SKrR3qEB5Jda
Cix9ciHawPO8uEE1qJkBisOwY0Eth4zRkpzV5hQklq3UmzzlWPrsYcDHrSAkO/ME
tITh1NK1/3mAS1ks1FrmLXk5mGnHQcb+NyqLaMNxDR1P5FNPvJccFAdbdM32At0I
In0kmUg6yXSsjdrm0B9+pxDMoctSCTaGrf6gGEwBHrcUlgk3nMAn2rDqxdtJiQaI
fzGaExvtGV7SV9BhZehSY8vTafmRf6Zu8g4eMG4cuzO9/7zZJdr5dKppc5SwZAGL
Z65B7/dbJfZB3XaGwDPBe3bVHUc2LqPga+fryloZeK3JOuGiC+WH6PfWldUjs1bb
lbHXFpVZZ2ejjj1jhr9HrINcv57C3NPmIf5r00Sj/EJCZS5GLnfNTClurYuopzr9
k9u7HRHkkEyR/ivuqXjbwUUx02upgdeJu2qh+zt9WRsnrc41rC8UC+uBfBoSj55X
bVtfjRsFyVWH9HdcW4zPMGOl36+rrkFcwTQ6DxzbmO69sSG5AEHVDK6bt+lNyZ/l
tlsIUU2lOenbZyAOi8vrsxJli0ILBz9jy9hYKNwHgI6EoaWBmS8+CLwOsgXdC+xk
WIDIasmuDA2ww8c6R6oAfq3CY5UBZEnaNhl/i503djqDxLxfwhxOXP9C2hlNJvtG
IezkUNDXu7nZv5BkcRyyn6mDuJ6tkpVD7zpkr1c3uoPgMU+CEPxLdFxOpu9Uo6R/
h7Z1ilZhBJQ4mN/NXZvbYDGRN7FqxgcEs9tlsYEMvJrndGWd8h7FsE/RgdFNyfbI
KfgrPKhsr2Qzl/CqlZiIOf/utRxTLvj1hL4oz/LUJEwRYFY60tX0h3xn+299H4Ia
TOWUoI3EkrHku7ayXLgpbNOT5dirX83pJfg7KwHa6MbCQiL283ZEaTq05nMqqRZV
q7D5Nv6ZUKiAEE+b40ZCchF7gkwPGmYJ1BKwKpHbGm9o5PC01bLF6g7eZLnVzyPi
ry837lXgKUY8OC8f7pq6HUM74DQtbF94fPixfEnVpok+kNEKbjFtBupGr+p3RdDw
1s1bfVg8k//XU2ahA+4Oh9zYnojioo7Ms3PbjU5uIYT+0F1GSb5f04jSJ5DNuchN
dLr3yifevgH8rO6HUaXvkPlhEEcq7dXWN8CYWMqTjGG3NFqmH15BIHsw6BICL9wb
u9wTo3I5xSNzulfVFf90IFNAOt9OKZXBpabHTY6Vsu1TcxVtt1yoSSQ6lFOv9zbO
jpDGR7WXx/EyMiCI1IPu1VHoiVFk1Qwz0DRfhAXkObsPaaz5MydJpcr3Vg0aTSEy
kQMaVupN4+5iEr8151k9si0/P2l4RSaWviVmr4qF6NEyyQYfDHVdHoLZaduCt03w
IvuNXj35l98RE5AjHFCDcM6kYgne2WVdsV08kMkDS5oAuUHZVoGkSLKzaktOD751
tmjYaNVlnzwtD+7RQc/qU1KTckIJDzJghjNpxUA/0gqd00xpTlG8K8wD8unvEeT1
oCEb2bmbtGMKs3NPPN1D+1QOsBh0wscnQNUwiRAPTBBbwFDQoKuewhAVuY/9wwB8
jQSxNhXGVLYV+wENLr1It+uBbb/u2mlVyQlrJdcp9k7Y84IVZAX/CQvOKLcnsAUn
v0lOHLo014u6ry5CL56MN20amYNuoNo+5vYt4D/4gMiiuzAE+N8qpTklqGC7YejR
RF9Z4dNJ2p9ESZs7csuPLUASLQa/gfBFxlCbJQ6u7GQpRViLH9Zw8qUe3Se9qR1d
vnTWwCSPs9W98DFQTPDcbGgbnXcFWWXstpho9Uz8gFh+RzVz68GXVUZl5o41L+PI
/8vNUmTGgbRz/LxAKZRrm4RWiYbYgjz42X75Qd68JuYgIm5qJenB4mZ7HsixvOIc
VxmEjZVuKuxGk6y9cCVW/MBsgpVhka3We+6Dq+sFzB3/abvl+9VD5fi5Le/DDBT0
T7uTmoG2oRCyxOSs46ALrnPrVxiOg50QezrDNNXz+ttfyIeKLd5rky4EE89lr9QE
Ytf5R24Xi06QQX4Rv1ZAM2MgYTO1LpYH2X4qg1dz3cSFZ1Ta+dS4WQmgNTpNFHU5
FCqjCXHAFOiItfPv0ol5nOn5qtF8vI+5C3HDHn8bR9KPPvtdubmmxCdSp517tqXo
3QtwGd27g2SVUpLJEDEPlcAp/ztSHeiPyGXSZDvLNKRnLVABX1FqYaFnysjUtfh/
W+GZ+VVWWoRJLEhsNlXwpBUU8dzBKp5gOcnBub8Jpi9gLqLt9pmXqsxOsLiqx4aE
8nSOmHgLGNp2/v7yHYhEWo2K0FJNoa6KlCEIwzj6eBWJltIVw3mvLy6VrDXjjjlU
aSgeJQyKxZJC1l/esws9A13i0JVd/TU6qh7+9oSWlLoOEkIUNqGa7YVirx4RUMN6
Xu8tWynbxGm84JjZiIv3FWFB27Yocuk+RqwLE5LbGerAAUSZBe0GcsKUVS7b86aj
/jPedt9/6t5k3K9VrbFZznB3VkgMXruMthEsdNzUTUKOuNpC+vKC4Mv/2py4hUIL
7XxDOxYlSZEY9tvFiyzshq4qxZ0Ppghu0DGKn1US7dm04yRZrTI6eNUJBsHlx37H
XkpBGuUrJJlE7vNzf1RfWqiZOpw9KMAMBToYaMXKO8czq7eBNPrMrfiEzHuDBFMx
AhGbJBHwdc6ztAKCUrjfjN6jF63p7Z2GiWSH93xXq19gAxjW1XqfgA9Nne7RhMHn
Rl6NrGVg1zrA+8nmD4cftR/eV1cZeGo6ed7C4dN9da4APB57pNvMSAReCRFumn3X
UKYcOd06uyUxRX7Z3Bjdb4tmNmVnKLWFeEIjWkoIAob8h78B4RRwKgYxOCQvyvC8
V4zVXx3yz+zLIsTOb/gaRiVQWvaiOgDAOxLLi6vNV0n471gI+Wz2juJeo3yKQmYK
TsNfPxZ1HNxPccZp/lOStkOj6TuIoCDxlryOog4PXk/pPEDDOap8NILCWz6JOhS5
2RHaJjtQ+yXK9sOiJSZJ5ewDXNDSmcmU81LxobB3mzqaLNDT1c9pK9QR43/gH/Lx
b4SUGAFgdWeCs2nRvXKtq4kdMARkq05cWu0FKtDKvw09eSnzIPTIrcJOL11EKfHa
mEtVZVblv5yeNx4CeZRWJK/PNN9jFaHWQaeSvOnKX6kiSkoZbFPjbv7aYlSYllee
kh2A15IQNnE3KDtYWUOxLlgDl6fjTzi26VnLEepBC3uEfwnQDoRJd+J3YtxqjCFi
yt/AJyW/4Y6B0mvbU2ncDaS1ci0iteHu20oGCBJB/rcfLcLS1bSDwKY+zwJIsRiP
SOMZAwdOAcSqjiACxAwDcEpVSLyNL1VyFFkqNIYg6fLR6OUnp74YGfz45WgZ5cBV
Iz+atIKH899CHaxqdQvhC0gPaSKmDElV8iuKfb+4+GovZw8BhUkBhXdNyCL2kPFm
pvB7EnZXFX0kKVB9hEh8+7xM3pQ/yQhQHQJFMDZhBjUGuvDno5At5OgVg2tnwqv7
vfIF/RjRhzWSyyz6IsEkbRC2QLcmp8hU/a2OJ5qCtlfvJCLbRw69Jtq/RH0aDOhU
w5QxiUxZ3Kqmtr21a1ZM/u/AdaSjjsyRB/xUR/WPuRSujeKtpdNssaUBFVAOR9x6
goZQNbVIy4+Ux3xjeZ/C8m9pQVG9S3C3GMMFc77Pb0NrdpBuX1ZZItqqsr8qZO9A
VqwhDav8wI73EPEe8Q6mGpUGeleYyXk/SLabGKy6uJ0ihbVO66jw7Yvktm4u/Kh+
u6UpMU3EUBATetKpqNWPvpxEvqBp6du2V7gNztKdPtpHxcb6oAXRvMdTaslesfCh
QqdnK+5I8ufXHfBi0B1TY/og6QQze2lCAkBvEB3DrxDX3lJ6pB4NjC2yRLbjFBO/
EvRhEj1loZV/RlUMlXe5y3btqT33RpkSSn8xQNm2UvneX/ZZUGz3oGoRFnMx8JxS
PruvD/m1dvIrVXrniJ5ZZCgttRLinVnMSbphH2OJD5++fhUmWj/J2kBtNOn7BRFI
VBfOAJ/NbCRffFeNfcbFjOXOjz82Rt8mSG/sp1/UMHexoTOhXd1F3d3/4pnmkfmV
1NAXsHb+bBrx56VcDJY30D5qAtV5mGKkkEu6g5fZQzmTMNfgFw7xQVkBa7n2aoC1
LcosTFvFgh3SQv59vKBUxpi2mgO4J410ZJBU7k8wGp1haNuRO47PfxroutgfX7I1
z0cpL5CqcTGbDaqX2iJRji0Wbli5p8xC1BZSr0WHDOxrsW2vTLDjkZX3KzulBwtQ
sZn1/OSWKI3lnpOztqB9EZoZ39Qgyo5XLq2JxcFNFwk7wuJ3Wt2MhCRsn3mdJbJ6
x9Km7pXnHV6y6xW0dWQPAkzoxvsE1fciaVjHKq+K5F5xqoQrUopv/rKa9H+yNuKA
RhHNZVq2/TabzJ4cSAt3z78SjIk9moLHHy3UDRxazqWft028U+HwK0gCv6h4n8ad
HnKTboew6iQ7QT21+8h7g+CF4votS7zAUy8W3hDHI/D20Vh0W7AP5cY9z5snRp9z
MdWaw38d5bh8UGY+nJ76KSDQ/seRT0abp71iRcYzl3QgDe0iOPWNyqTOPbE745wv
rURTmPeh/hv4saCLsHHWh2P4dRbomdPw+qc/ZOdaNtg7SSZgEFKRomIZ4EnwLgb9
t4TevjRsE4EHS76x+Ry2ye5t4qo5GgBxWm94TiLKofQ+URpcZg7BmLmw8Mylrpvj
S3I4PY79O+6QG9Wz3dDgobKh28g6/AIocEgY28SKnw9Hml5dojCeQCe4HL5TDG+L
he+NU6JOLAAVN/+9ngLDunqYyHK3smT0IKHPnXkSmo38PaMD/bssz7is8xLeO7/8
ibgQXSnXsiOMGHKarzeo8Sm+4txIousHlYMOETu/84pl6KnjFOYssixmzvACT8cP
ZplKFu+FJF8kyM1G+1KeSZP7iaevSu2CmdGrTYC8/CqYMYZ7bSIzQvQsDJ/jgkuZ
ZntxqQrQopCPOqlIt5ejJFJexRZQzQD3NyWbqjf0/VYhx71ZW4/sB4Nl0H8pi19O
M7YeIOfXUVBX0vlBHElqHL01XZFMZX+n6Zx942LG/7mwYFQAcL4etVrVBERJ931r
jBYzoEyBfHpiX1R7rjY+eC6hlDiWTnTXuSb45eto9Wc9La/7J+47sALgVb8XqFVQ
paBrw1JN5BIYWA1Y45av4JYr7OtXIR6QI4qKc5Nw7v6d6Md0phHqmUkwvfxV3xDh
juELvkcr09pWwsUKTiQRm4WTxiEhtJoZTbmzJWzkqHNLmyDdUBDWWCUNsJcIulfr
sFDOETiypUs8oZZ7tWPar6E0E7ZECrBgAHe1Oav5FEbkGaMxYY8X/CkVKp3HxTNK
jBzxjXfW9uPm9+iRBekRLqfwaoFo1EkLKgDizpKz0Y1OEzYGYGHaJFwTFmGQldyi
iKsFEhOv5cVNqU09f2U3z4HVc4rjjm/fRXtameqWEyd5WjiCHR47rXilGgd9bhdF
tkIl9lj+D2o2SeMVERK44F1M5703KyBmJP1GftjPqgiRaT5/fs5l5jMjRhI07qZx
8n6iwx4lrSiEbN9zy3mxVItplHIN7hHKi3P+vDFTIkPRSdl875Z74p7ihpIWQsZm
Hs4STzUN1DZMjR2ssrIYSNUYFqqv7A11Ykk49moleTT1AJXSOMSU2g+t7oL8G4nI
+k5W4p4tmiP28i2gs5LG9bcsV8hfx4H8KDghsFuhDqLHchcP5kUsj2B2qEsnagls
tsvbWk6t6IdcsnHAAnQffMvRVOcZJ+N8lOWtFyJtTlhYUPRIvAUgNbOfcaEGc+DR
6iYvyjkNJah7fUa+bfc6dwnNtLQcG6rzwHsuGdwFs+YMibNBoMLUhVf/8X1ypyMn
`protect END_PROTECTED
