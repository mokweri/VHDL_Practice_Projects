`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCO9fHtLSy0cvDtH/CB5XE7CAYFXDP2Hpokistv5LY8xa+2TqdV29XODudFQEakH
oIuxk8TvfrkJH/q8HonefZqFIE0cRSvKA4GtaIvKTtRBgrSxuq7P1UJTLZOjOyRe
TFJh3crBTuUIJ/xR6ETPjYVtrvXD5+srVdudP2xfsO+AK7+JMxCWiQ7rtJeKyKia
2iNx5JgGg4TjG97ZvfwFP84krdn50qTVErLxNYGnXIebs0P5rFvxh5HtW02GJ5z2
8C/YFXxx3hhmS1EIkVuMI5thm5HZfxzE23JC9livYiVHSYGMuhUd98AyMNVxR1Pq
XIV95edJuUEDWXnUKfba+X+0/IOzONlAMLqVMyicmQYEkGD2l1TPsPxnSQjehtZS
ggXFdoL4Ty2qmy0fhzJ5l3smQujLCmkMm0DLMDYrZ0MFA7uxtXFgCMkJZyWhl1r+
1tIWFU6xTADt1pN7oHL/hlaqYDq2SV1zVrg4WnreDPbHTM1qSSn8spxvPwr/7oHk
87ts0RrLvs7i1BTDZwTmJTSw87vRnsbvr7H548+XC54vLwHiX9ewmaCe1WUT1KeH
49P93Rlqjs3mOEqAIe8kHSXmz7dxFitMz/6kaTOoDIGgTDm/Ss+WeAoHMnOC/DcT
0MokgGr+rEapjus71/R8usustEZyPZiEMWPtNC4VlbJk9gcD3KIWl1UU4RqpALDb
hVhlQChcwjzBkjAKRIRGi84f6teS3CH9diUxU0UpWMt8qlwJrEzyjsJqp5HQS5XJ
sJlHtloZMO81G5qwvQrRqifRqhRMd+b8/r3f6MLK/tA/j9EEusQEjF54CoGN2cd5
KiC8LO7XNhkhVDgpP9Ld7xZPAm6I45lLCm3dsRkGSbNURf3hRv/351bkmdFMFTpp
ocap9tn1jsUWYXAkit8Hu9Eecy+92cW57qndkPxBWkA=
`protect END_PROTECTED
