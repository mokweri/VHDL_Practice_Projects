`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPbRCQgSBoNXOB7ufYx2vixcZJveze6Z8oLqAjD4gIaOph4GnGZHqOThNVQ3TMpL
RsQAHcCItGS0cUtbRKJYGCgncNQr17OY+IO551SOe+OF+gYhBipQ7Q5QANKwKNwd
wA31Cmt2djGtjqCfQeAGPREDGn4k42nvnDVndfwzKRiquF7rjqjgiJi4TNH62Qx3
gZVoWqTmlychw1z73MgsoSRQf5KSrj9Vk0tQpE6eKE9tWryqzGHMno5o2llbq5zp
askBildz9NqdEZri5TyiTSOL5iqpNZy4HUGsSuXG5lTJARi/KhONxEteGdHGff7n
lBwSslVLLFuo8wYmj+5S7NZN1zhwLV/4uqLj+wGygaNFPIlblrd5l2nxn/ifp0hJ
16czm9YQMq5GU+HijnC5vV3ME93oN/HpJXhndvgEsHjo/j1leG8HcqgZp5SvD987
2WtAXPQ++GZLmDpJFhpR3x3q9Xqp337bisouTPUIxRVCtL84WjIZ/b2m9JQaJ+eg
SXYMd8hWzUC1nxqvzs/1vvizjpBNpStXUKDw05c2bkE7x/E1Nb97M3HpbAeVhFwv
g+uDAd0YxD1XfuyT4wsrDrp3qMbBpTarjXY1OSVei+wI/1TfrCiAuc9yJWdrwfY7
wiquFOFhPZOSmH03Esd+T5l4MXZ98KveNguHsFkvDsmYGXROWb9ZHdKEic+0RXQJ
4FbPdHacH8fM9UKcn2lar8RTXBvW3dILftC/lwGZVRtStZgivoAqdgmNOOZSEGA7
IO6LyRpn4pbuTZitRH9Qlk/cQRBejDcCoXPkEhS9BBsxd5xGiiHSbz0x5SzBof7L
eCzmB04MmteHGLK+0DMcvTW6Wa/3Icf3yrui0hDO34Mh0HhHwerWjRfNDC+t3uS1
wJ7mvytsvkPujw0QOwH8KExgF0i+nUOq6gPM/bNbUkkx0xLGrDMn0e1tdAc6Dp/z
lXU/dob8s/2tJaWrRt/6MAjimT5XsiGptbeGz86kKT5Hmy3WWhImlmDd2ZCHumW2
3VwS+0uCbhYwrYlDLrP/CHVTJXPzskApEAPaQA2iabtldU2pT6MKpSxMqxUeSxRu
NiAs+0g3OT7SqimHAy3ZpYxXvM3LGJz4dWLMmKgsHjw1bIhi05dydFM7FZ96y22C
4Su5PBEHhNz/eRqdwS7QipalBCGdbfp2DJiVhtyaSmhrGb4l7C4J8RG8RRjTsoS1
MNMsbhN3kvoj3I9Xx2iN7CDT2sHFlhlzxdSx6i1sm2xdl13BCZlLKhatDL5E7Wpm
fUYRzkvN3kAJRe4LAnKIQA7P6XzDs8yNZC5/1CRPV3ExTrY/LmuH/uOkVo4MeODc
WDrqgRhhOoTqNezJ+qcbRvYr2tqlHOrau5a436vUy7lX1ZLwevIPOstO50zLWnXr
tzTTVyZzwNeOh1UD2q2AjIO/Fb52pI4nvSSwkUuiJtrTclb0LJMbMtmojsY0tM02
N8H0tCgMnQfAvpM9mp9f12t4rLev2Ey2OL2LazY5YRHjrkAD806yJ5dBTvM87QHZ
xGdV/l1utgXh9k4rX6ObCZFHHUsgpy8EdH8kbLTc9AfjQmIweDrgN4rIPtdsXD6z
9lCLnKUAc4nmlVSEtViZzQUJ50CV9oO7DfHlMLVh2bpMR+XmfbfcUR4hjSwt3v8R
wMSehm1xluLfCnac+mIFcZBsdfLZ+ujQYkr5+jUFLXovwwwul4iI4Iii9lN8mZ+q
Mg0VjyoblmNVGS8TI0JCItaI+0GAdR8h8p/kL1lcu7j3XxRHjkizULF0jZLFo+Xn
TTV0pNCbmid3et0mWSmUdLoUiVOI42J2F5j3brA3erNpWBgYfaka1NB0k8+Lgf+a
EcEPTDKCzvNN76Tv6WZ8lodAFm9HzGCgBmAIbhyP1Vbpqb/tUGwvAOa1NZ5Yv9+d
fewQg/4PpGXuwQPjw81879hFpMOUhUHCkYsaM0gDY2+IPMrTy38tlrEQiNOgZccj
eLM32hQKVMoM9/Kl+Rkwkv3g8EpeA92pzYEGQg54pecPhZJY0zk0T0QWS/ZjxP5h
/SeXlK57Z2C501TTDrxQ2+I2dpaYKw/IGlHxRFWhd8SdEFtFGbgk+2HwoBFrONtx
r1/djHnffDgpIzHS7RvzIfAc+JkIV7+UFme00PoZ2xpLL781ARdkVv98fUUQTMEO
7f2u23luqWY4eJOBJi9N7HU0Vsu9BvL1WxfE7nVNpZgG9sQqYFZoH7wclv1MjlUS
yr8YPMsn/z8GBa4+NEFFdt9auESf81Ob5DB+arWNnBrmFCz4o4R7UIeaOEnx1EYv
2+mVPYv/5qFw+NpYnOR2jlG+izSD/pWQUYy4Mof5EqlSnLoCeG2bjU4lPwCQfPGe
KmS4sfHngwozy9aDbYhXY7MSOSFuqVjEpaF2ybXZgHAt9bU8g8v0HCHBAoundzK/
5gJg5Z/YIM1qVL8uigNCZBjfphNZ5WB6AWD3zf/G3PWjKjGHgwZU385Ag2L1gHrF
oHPsSwSJuEDLXWV9Wm+DAXlG6j5RF2qUI1c5poa2Tm4zSekD6zrFlbSjPxZ4yiIX
82r0aFBOtCGAqaWD9VloCpQDRvV/XapWVGllUq1phXnrYzF51/nCf9KpbYoZ7s5p
ff5hsuUkkXfYl4xNyerqnM4cRkf4ZdN8TJgHJy8YfdkaXHoA4hehdBR2aEgOt75n
rI3gG/SjmE5ERbAfju2UWqiHJ649FDHp4DAPxb8On+Z5a63RqvTvwmp3BUjj5ckK
cuNtTvEy7/sJF+QIWJP/kb7Am3doyMaXV8PHJ4zzUtY9JcGrGM16Ih5sx5zYKIbC
jJk4WdOMoOIEMTWdrgs+Y0/Ht2p7GBsZBBMTshtcfG9n7Q0owsfcalzW+WsFLiIF
Vhf4VO4j5xHttLq6vrSN0OYg9R/VTTvNTz0wptUVaTryR5UFFAvPJ/ZhlokPQWy7
wthHWriiV72+MTo3RMZnscNIX1zWYmqW+WK72lduoE0O1XOK3bwBkbqh80phuET5
KZ4XABhi5oWnlAZW8/L/8HlbfQDuV/xbpTteU13RWHOJzO7/bdaGGynIHDbR7ae0
qF/u4n+Go9ZkSpyU2HfFQr1pYI/uYjnyUMtp+UvyhYwKQnaJhA4eLh3Tj0i6yzb/
bdIf6EDsGDFy4/7icqaWyDc6QjKL11zRqomQV0E7CGzaSVdGLlIxfNbLmsTrSUP7
aRvtIShWkOAHTAG29wpMjg/tof0aF6rfgt463t79tslisAroV75eJsPa9CG1yDEM
ZL+FQunARH24qkmqmUyskMvOx3CPu2TOSXLuI9eAupFE+QsV4D8N2vuQPZ/Tq50s
0GvBriHJx/ELOlRCcsekhXvGSFeSeejZA0RhJXhMvxFVSTaEmKISoAvSLIaMP5In
RfnIOqZwHOY/xV8TXMmKr/m3NK+zjjNGgcbFu8Y22INIBaZBubvOq0N+nOpqzX1z
IvR9AA+4UnSTyqA5ldDQm7SmEm1J8uUoKFXryjSkZkI7G5Y2LhqSoUekoLjRBp0M
AIFrFKRcq3wVH9FCBVaIctY7BOk9f9tR8mS2vBvUBUYS+0xpFwzJp8nMVlDaU9PR
SfZw2oZP0um0h1CqJzSk2osjs/5yvbiVs78C4CcUFxQiYM4/cGrUjixHRiQ8Be0v
/MfOcFB9i5rEsJVvlpQu6kopJFZKXJU0N07k5vuW+1TlqyCtXXc+WQlIM1F3ULO5
1vUjvi4M4NFzk/CKX1lLr3N9WOxnY8lq36VZNcdm0AOBL1MZ6bkWIPEzsKLtsED1
IH8MMGpAOqrHFW/FhbcoC2GeJ0A4YHDAPoBR3o2djYDc8wyIcseMuYbadv2OLmhv
Eul21JZs/PCDsdvl/9HBb8ZuEcqwKHvht760qOtnJcXIPoeGhNGnq6fpF5JZCV0T
2RpZpsge1+yJwkuvDQALLkxMHfvfev9Xfgn+ErOG+Vl01AVKzqwQPzbaibd1Xbpb
yHyEH+TJDftP5JIi/62sk+wfkJ82yf7sT7EcoQu+ODNP2FmEg7OJy2tzIEe3y8d+
5P+jpt2E/jo9sCwpBs32VQ==
`protect END_PROTECTED
