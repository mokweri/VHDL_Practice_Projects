`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OM63YOe1R0yLMMvFiOHZ7CXS0S8iP1+O64+kUVoadYJ6g3jHGpnInDM5iH2DWTls
hbtzsuQWc2KD/E6vRvA9vaiBV8fgMyaZr2dkvUH13zzXdSW8uIQmqxv6mH71xd5h
T85Ih+Kc3rGZ5jO8SU+UZU6AhsLStkaTM1Aj2UYw98++ArD6G5k/NfcDILic1afl
C7FJCx4zIzUa+Y8TPX+owxADTmGZSUJi6noM/mDekEUcCFLpnPo2wDkaOES8bEFA
gOWvnB+uXfn8+DHqcCB4VT0lttNBnU43lmY9jLNT7pXWC/EG6tfp+dwMbm1OrRq7
OvcB1nICoEJakSvVZZvivy9+eE6+ERimVod8vSsVXf5EUaASVm+SUnEiMwWuSbqC
Y+d9ex16id6fzQtvVpReAzTn7WoO9b4BVaCi0k3WMPcNYUvHU/dFnKQuOd1/9odv
/EZW5m205La1/T7RGpdS/Ghlb0xUMX1Jh3mqmYLiu4qrbIfBOSOSkWPMuAtb1bDo
JTBegHFbX9g3IhiOtn2tzovclVr5aTPb/rveo/fYU4u0WYVvqv1kr9hRvQJDbsj6
xkSdeRo9zkrkPsGgFJbutbuZzJgmZIFYEhccXvSO4u9zd5fCjtdB8GbRkExn0qjc
lTb2FtxXRsdEBke3WuYSj0HsS5BkyONQMGsORD4xKFvJikkcokHhbVFYWaZFeKII
NRmdFHEOLUVhj7F7hk1zOzKk8aoUaSgHHegm5c0yQBGGwedhJpHEBcn599k0Zz2a
d0LE3eq5fdmspY1jwMOqoJUuWlZAbqnQUR4rZmZTcKDiFvAdsGtRA20x9BqpuYV3
2gVTnqXYhwGGeu/3+ylGOPF7sGTtw3gWyabJBJI4Dnu3W62+oHHOtChAPNwgKvXL
+9z+bWe4roq/FZh5jq1ZCEJGaS9vrlpmzQtWVXa9uWYcxhYGZlKPW8jFcMcBaNe2
GKE5z16jkKlX08l36yo8xgGGV3kKEg5oFqTUZePOEGJOO503aWBsSY5K92yyiSB2
oqH6QPLznHZ1zdwgP5u1WDNBxlLCpEDc1pkX4z2wrYggoQqqBDWJXmo4G2WmqGYT
BRHN4fjFwoqAQ3Ta/illIfgT2LKTU1JU7LBYmeBBvjRfRw1L+GSzjgssVG3EBf8X
mHQNpx658Yo8VOo3vMyPl8AlhS87ZhtJNgsGfo3BSTcqorasVHoHNqmj8jAFwimi
ns8PU/Jk/JPeoGzwWdMSnT4EAMVK8vmBaQ/m1odhEPQ1EHbwgbYsZ6FxKjqplnXq
dnqbiTLHosz7lZmXw9yHp9t34RLzJiHu2dQZam+uYQI67xvMO0w1JWvZ4/K9cbzx
p0SWTnEFb3IgYeu7xeTBn9cFfBpaKrjT2ygNYVfhX1io/003QIWLfwSWhLPx9ZWd
QDzP2mT4wbzy52j4Jhxh7TqRff47O784dUoZjmnjVAY1H4qI8CyuclNHWjDCEwmx
hlulQzSe0B8Z3h6O/fLxAh9shQpVB6kj8MrM1LC9SPRuMwvExsspeHitZyAG0x6s
BjC2/FAKB9GANFTQR0fAwojAIHzBUF+27WFe/4taZViyBlTD3cP9gXTh7/xt3eiZ
NGJqcDuLzO5OnnD5MdcqD2cX7emsGvt2xfnqjl2vSzAia3aWTpJH8x9nsel3P7Ib
DnIQkl4hq/2TbonUTJu5zvssmG1RzDExuo4VsqIEUV+rSu4ClJ1Uk5kMCKpNCbge
6dSGeZ5cCGCzrQzxl+1QSqdQ5BfVLxb0xbM0mhIfRBec4iZ3/YwybsVngGp6ujg8
TCLl4dmPXzmYhoG4Ohl3tDj4LcQkbU3lPzGlzj0BUlYLzXBGL8vdShBaHkK/0hmX
6XhA6JFFlSNgMARYt4Evo9o2Qvnj6Qcb1fQayqnVhprH3jS0szPIIlplx2yhnWj5
+XgOU0DGt09I/SD8siq4q8KVwihWu4mYlX6xO7U9VDLhSFBR8qp1L1PtbabzwGn+
pBeyjW9zmfFG495lkemuenvkRDSbUEcjnC0kljCbtUHBysS+A/PAqEephRf7i/Ib
n7KQfOSaF8Nt9qbCE9CaCuyIMoDQs5scZQVaC7ZpcR62ucbg+aNuEIC5GqqqKnio
J4tW7YHtLYaj5G5eRSYdlUQGqhiQmcAowFwTKjQpXk4BZHYtURyj9xS/e2aE11HL
n1iSYLuinL0S87q3c9Enm5D8kBdpBuvIAwy97wkjmxeymPDxR/uRg8v/JFkHaeYN
tCbeGDytZtgNecUu78dU21ueJZyYmME2DJhrtIyLG+qV1Cmp/zRJhb4q5s9m+1Ys
InizVH3+nXNkLnycgVmgRevGzrFQnql3EV4X7PstUiGrMfrky/IJHz4gDDHpukXN
MI8Zg4O63bfCwOHp3mjvMnh0Xa4gos2w+LkyDrXKtrfwOILJeQOlr4AK+XxGTiRy
ReJyEdcJBRoP57XlHj7E4UVFDMXKHgTsWp3+NYJ69EQiVFrtla6REIVgt+j9lSAr
GJpJsSDMhX0fNqh6nERT5A==
`protect END_PROTECTED
