`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvlOqpG11m6ZlRGsd1wpRWc99pZLACcg8iGRbTdYaJpqTS4d85s7GUh/APkazLt5
7Xkh+jrN4izww9lkljmmnGZTZHrjnh/zg2iIadxzLuXXkqTYyPxsv7bnSH/s7BWD
LsYWON88fgG7iIfIZElli0bSmPE+1ygwpCzehA9joYT1ZQrgPGqd01XoVeFREvqT
vGlf21bWjTR6d3KqFA7H8taSJFFK3isnO46eHBh6WaWa2hEaQn0K/PWA5Xu2eL8x
uticy409O35jx4GWZZVDV0Z+WVUBjwPvp3LgmFjtfFu/gwb3LhHil3Um1bpeE/sM
o5nuOu5hMncqLvx8qZCWTRDzDl5wB3oGq62ZYOa8Rs3H7qsVdOe/5yguEgvi8HkU
K2qDhSoi9wlVoFmAh8onqchURkaTFlDLrKGt3fFMlDtqsq322zUbPCRB7/fAoBnY
pqG/zrdp6txega8meKzZDnomKLt1hbkCvOy3mdrphE9DAG0P4faTfCTMgZMiNxq3
/9CslkDRJbKIzl5BWy0Pc492fJHtnNHZBQj4dl/7wvyiOonSp5RFmqbGykdRXiiA
GVV8b6EF69f2cY9IqqNWDPvboQ81i9QMH9HJhKGW1qhvJKN4upaXQJfr2oAb+jcH
NtY+l2RBqPWd6j7e3OpULQ+dUX5scST8FKNVNtL+eSFHkKLRBOmZzsaTUhx4rL2O
mlmVZUwcSu2bZuTVsciOO9/kczoOGogddr9GXyBMF6TN4Cdneea+qHYKiZmJMEJN
T8EtouN7n4ZO3Euc423c65A3f4ugW9Va7WruJ0bGF/3KNR4ElTgDLIbPxXcMlDLE
xIz4grZjFAU4xVzuduGIv/8zModaj+flimHYBL79XBRBclrfYlTTYzbv4NrWO1vI
O1u0rxm61vwIIbs85QSKYAFyViMts215gce7T+kxHxfjPVyZQgKn4DVfjdOlEs/I
oRt5TvZ3EEJvpFFP2aEq+eQKLJMJ6xt70NfmjxR+4Ufpyp8o/X8n5A90/+5IQ04T
vkOfkn+yVUQU+hrIQm6zTDbOADr9gWg6Qcvi1sPqTFZGtRZrWTX91wlAXHGzZE/g
x65NaeHmJlf1IQUqy4WlCtlwxpNCMROSW4N2rScxKhc5sjzGChDIXtCaixsJ6HcE
mS2AV0+IQs4PVOwKZA/9YMLOvd0qernIQkiSdNES9NcA77Aoj2JNFlrUfTY6vRVH
4VPWooFPf0DWyGCjgtEzFw==
`protect END_PROTECTED
