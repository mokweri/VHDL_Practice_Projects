`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w7/OwCYYoxrgnq5kxLOqZ05fo7CDk3foGDNob+ghtStqVTTWB+AE9OsyWuLCIb5W
nCNiS5L37oFh/CIWT9kpj3WECwT6IkerFr/rTbU3M4dcaFrgcHrYdeZaz4HkBFaj
hCHsjpffMpGbwE0Q0wy/CUv/4x7lDJVOc0u4AvLi7qYlD5oR6r4v09yMqcn8t3u8
eZ7xlybpoU3dW3pKtHEXHC3k3YnYr0zM7UG2xfncng7gMg8hT0sC9e9F82AMilIT
FpBA6G+PxUnB8m6IfKBFYcGjirAPPh0KmzMLoZPHuAMXn5oQvM9VqtEd4NX4nPGH
NdJuA+JjGHIfbKxAY+D3SK1KfHoabN4pQAB6yYfTCvNpqGJwvrCVJkE9dJH893iG
kzvsIPIUlHtBtn3xFu5Uhwg0XAoMAAFePft6WpTLoLCeAWB11nddZyCL5E2+9iR/
HkVCV667pKGCbLz4V0Hd30bJ7271aphzQjQRA8HwgBlLTf8nZwYa5AbERsUfAq+8
qdpuv81aIUbii+pRc84OU4GP9vcxLHnyI6hAl+Xzz50v82+5Dj8GBCJ7uEhTW6MH
WEjFxnEPeLEd6YnzNIbai23fpzARFCVNlNYwAYv5zcZRp1ZHQmnMmsNGWsCHcHDV
QKkMVDfOVMDsN+meNWRJ8tjH9EwHLg+gfw7op9EMl3GSCd3i7wM5h1ia0DY0brqN
5bed3Ju6w3yGjsP4hM1ejCvnK+VTefw6k3t4E8C/DPm9zcfkSZgLt/qQPQh9jnh5
nldPeujpk8JJKxatgvmkWwNr5BSE1hDflxbMAVPy3qV5kWcnsW5bibJYlBRd+vKj
RSk1++nNqbiuGkows4dv0E74HDYAcfeGYOowXAG8//CHkq7LJUiEY7S9x3qkgdbV
atAsySL2xb5kexmgrtx10IA2mwb/6XLMPcBSSPcWB67cXDFt2MxVH8j7mNtjy7tX
L/CDDP9tTQcveBkhVkoslEKizW7lKY+Ina2g7SJbES+5T3LnBE2ywe+t/mRNcG/Q
9hhLQkkon/CouJa0BlCmXZpRUnS7rm6r8Uh3RAXkw/1Xr3frl1neFFkag8upFWL3
JTe/tf+Of49WIxvq/DjH8spBOfw4pfBFBhhFvO21HSnmX2EsypJJARlNSfAJhE63
4cgGnEU3T1i/sDHvoaIa3NkjQKAAqyUknVmD6a6FOJrlo/T+tYK5Lycl4tNTAMEu
RDRlHA7U+IW5Ggr48ARF6MpPBTvUYg7ASLAQF1HvTTh+zTM6BDL5WqObNo2teKKO
GCVvJndGcpvA4ERhP8bA6e9bXkZJgc+bjZrFLLaYuioKeBnW+7bhEiqfYgVOvJA6
WHY18ilGgMvaXzKoHGaUde3ylyuwtLQjExXoaM+k7QUvxgFkQ0zzOriqTfhgeCRE
NzN6kizW3nyLRiBMYZjckGXOdA2Hua2cvecMCeH0TuQuG6gsk7iiLb/U7R41U8Rn
6+rTU+KWGi3C8Qal+f0NjrbLTAyRk/aZqVZPwH8nR4H2dLSWUcvxv0DIFUePChn9
SyCQwZTX/N6HVnEbVuG+jMbLlzWBXjDK6cd/cIWWaoA19KKsV93L6vC+/FlXObws
Jh3M/O5r8CUq41ajW8xoPNrnj6DpmlC75X4jdg7NJLy6NC3EoGAqOXLAzLn0ulrO
AzS1JD/dgMNb3h/mjGoZY6gdoQozxYTIM3c10BA4gr/ourQAC+XKDKEow5g6H3Xq
Q4MS+MbDIvmagOkFHiJpkCMrVjMirgqMDFZ7zW9OD/o=
`protect END_PROTECTED
