`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONzxWCn5ZnXv0smYsrEEyc8gFj74oxuSJRB5xTjnLDAjw01X+CBegfrqA+qVC0oY
b814i2eqWz4X2IbDXOD/cEqYZqYM5LylUZum8Bv/PpOGCbJjqrXPn+2kYu/6T0N1
SKJWd5jOR7mH6vhvuEQnKXmj08CVyVmD6exffJOokbLd36pkbsjOQa7P0t6NmG6/
K7XnH8nKcSC+k7e2yEtWdVOYtotBr5gFFQObRNll2asdPzmtunA41mm9ot7WMN4i
Qxub2AnFMOqVXyLPl7rAxucJVeaITe+g3OtFd/vpydjMFIVpMQDrD9X5b3Zr2pEP
XgxxOy1LU6HNvn4pWYfxbt807KCCzZveIl0nvjovIy7gY7s1F7wx6tL8oa1GaWzq
wOBwG/XfKc/S20HzuLbhtoLRmnpUC6yNJBpI+0vitkydXsOPZoeHlKNONP1DjfGz
A5m+w7WYdYc1/bLZ00rjxXUhzWSjnlQh4kzjSDEx9qdoDlJmQ/0LHodUBCZp/17J
qjpHS853F/glaupymo82GZzFKVyGdlsZV9itai3q4FFHb9Y8bTjT5GeeTBB21yEm
/B+6M+4equaHlyP2Dc1SZAmcTVgvQHhM6wEgN+rbDAsV02FxfPjCnDRowH2dDIn9
ZGHknvrVN50lqhkkoO9IDu3uuD6wnDOcTsUhib+NInsAfPk16VqYWsKfYdkeYpHo
EYziGQ3sbJ6fYFS5z9iYun4vSCnXQAM8/QQL/uzaRkKgBMl3HafExCl93z1X1KRW
yyrSKObB7nGKpsGjdouzhtctCFlQke8MPEzM96782O6NePh1TxmlJRUf9mKRNjop
5j/0oqF1Qu16pE7QoNtCMcPHwXK9iBgxNHhBMPrINxEbbISTfomdUnCkD7On3US8
IWsRU6y4htJLos4f94Mm9x8L7B3apX3A4/XuswlG3lm5RCrgGIYKQUh2xIm+1dHb
UC9lK/iybdlQZV3Gx/lsZzs4azHydgU+DgU2xs18AAHYOXHl3xgeaWFO+9jCSjsb
b4f+Sz4mr+OBHhczGCE0il/prlnRM6IizmLlT0ZW95JT0wAR9t0ZzwNPl0wobSny
3fQGW3sZSe+fbz+bq+L8D7AUrsCskqyrccjigKpVAmX8Oq/DZaHAhhZTkrnCYjDF
tvoFYO47Kw3sm8exoVlt9A/RVdpn1yL/e1jDMtIIBiMG1MTZxf2IOkBiaQcxITbg
9j5pOUzqzgEM4xXQ0yZ5qZPjZZsOEB6DPCWIzYDITWUhK4oXAmpLQasUAJZTA2qW
`protect END_PROTECTED
