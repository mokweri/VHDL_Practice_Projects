`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ded9w0eC5fZjDlapPxzomICd7JIqu+YqfbIVHDHs99T5CiAQxq8YxOUg0kwhZMtg
hb9adqlj6n24ytt6DvSRvNMm06LnN0JkLUSvva8AbTErz4fLu88EJnwWvrvOEewb
8az8TnsIa9t0qcWHBQbe0PdiNLNNjArt7DYzV/r9UtNclLd+WUFs9xxotBFLiZuq
JahgloBaLozUxzMzCa986+FvH/IHaZas8AkIC8cMpPz+EU63uGJrk6g0PcSeGNyb
QRHu9UnY42JZ2swfKyIRm7Z7A1gk67xBmxRxX7HSQcfciVNC6U4HUUloHS+JQlC0
UzJqrhcd+og47hNX2pyU0itB0M2Iwe2dx2+L9Ohbn0lr7R+AqbaKGZfJ0hDdAnx4
`protect END_PROTECTED
