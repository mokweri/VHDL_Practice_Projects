`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDyttK0PoHv6g6tejg7n3zpU4RhYvdhlDKmgIRzOLGyZlVMMIdXl4+MJH0wDylpA
JElYTa9Gl6dC1lQl2xHlk+LPAJhCPeJ9VLgtpX7R+Fp91OGVpXi0s5yKuv77KifB
dF1gjLSeRC5Z6xp4gNVlGTcstiYIbo3MVDQ4IcfPYwxWJwvFTyHQdlmqQb9/Jhcz
moClR4O2a55PYhIp0h1+W3TTQHsQSxiPm3pwuoEYqVDRXp/Kv7qJIqXdoTrWaS0d
PxeH/4lY22ktynLz+yI2mfSHooie7U2e2BYmVPPCjM3ujsXzWVBX8jtT2EmQj8ln
XBHXch8DbjeimxAD9aMwPGH2vFgJPCWK6q0SzTDbXxEkjcvv1Y/Fy8BCY/aAyQqQ
IK3gJO5VWctzMwJQwgqsPOkstoKERS4uRYphdBojpQVzL1eQGf2upGqZnYtNjZjB
2ztJTwBsEoS/DafIoCnEj9CazzweN26wyFLT5GaoBpf2GoIlFSsr6Yd12S+rgndL
yfzqJjoG4J0i6875g757wsdCMXPHUanSKM42JFCrOF1TuVo/5sMwS0YvVIWAVIEe
rZN1IWNgUKCn80oZfq108c2eU4D1VhrHMzhdThsNgic/MaXGccOENMuw3TiHXK/u
hmsy42VPSmEgMfitH/2dNQi658Pv0rWx79WRvLgnNLo2itRK7h0K7ovGSUVGjWq3
faeCYvt1r8F4mNOEAbb7tF4BNkEJO7ErxwYd97zT+i7jgXWdEh/GbZ5m5P4gAVuG
X1zOMYZbW2W+qARBnn3gPA==
`protect END_PROTECTED
