`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhmFisUrsKfLqJrCJPp9SHHSq/kEFkfiXKRUerEedjF7pBlptNYSfpZjNFylmSpw
0ljwJK0rNetcmQzOKdbGe1mt4Mfxya4jel/wwXKH+hD123BjZeppjoqb/3fiVoCd
JgAK6XK7ggRqa40r+ZsjiZP+gtGeMLGGJPQfi0hknV9MI8KQtMBf0RAgMcFhMrgV
dTUXlXqDMx3ts4s/B0rwFEIkLjL/7NE4aUz2uj/0bPMwHoh8ncPjcX8exfMjEvk3
r2bu1CnttRTBJP4fWYdT+EpKty03vKS5ZylBMWOrpLmdBD0ASBcEQp6XevjDX7HN
t4I/cXi/Jl14mw8lxGYgCkXRnhChtU5q0FPRNf5JCMT+nHBb0ouVOaof0k0SP7/R
d1ip9HDdTjeVl3X7uvOIxHSuQhZFsXYltkor6uOSf2JRcWVdxnkaK3WCKoe9dk6G
z2gk/MqhLsjxsjlViON0yheRIn0q80L9hjxR3rcVyWRGc/XN7SLXCfekFR7xZtBm
T9bSe5DZA+ilot63Ngl+4XOxWk2cWQpIJmYWSUMSSaVbHFffXfVPm1Jyacoqk4sH
18F10qGe1l4za/GfZPAYlKNyzYx6hEyozor/y9sMrDw38vGi4z201q61qwvf4pi7
xlofWgOYEI4fdx92JZ4Fsynouq8mcWTZVrR+bPPbvywnzabjckPE0zWr2r2zc1uz
jhDCrSKl6dLdWQi5i/S2qYtfap/sI48kf2UoP8kgPZ2Hm+piUrFyCACnudCOK6C4
4xfFGfaiT71w1xIZJFBHXxBhCtAuwJ2j4Z44966yIt5Lv2uSNCXO2EsQMzdCm4nP
XswaPR+IL5yvd9z+oJ23fv6JW/KOwdOdqJvQMiYqwdf5qI9VS8oZZnIVz3tFDufo
5olhD0f74e8sGAUeKFG+9z0998+XBXyBBNJj6KYKeYnheQNRCiIRbdc+ZHM7j+GB
IwFVfMxcu1shoqXn1+h4smRdCbDjgDsLtvohl80zKAJiDyZ7Cu8q5bvYDZbm8poY
A7bTyPk79GOIXeBnc4HbRDSTYxXoOewsahOIIppE48K46GtHb/kbyFvSS5w88T34
32h+EGxQanelJ3o9boPinFfvRDrHyoWqeR/JPVYVM/VGeCcEBN2B71+lmCad213R
9Z2EZ4k/TX42bIUkNXfu1WZbPILuZp+hBS+xrpv7arf2wujBShDiTri92apSPZvB
Urv8ejuXvpIuqW94epDrCzs51xouybDnqtD5Lki7IiSdd73luKyOs2kchofy/3hT
f/JbyxqW0G6vrVQVEHgZuo1HuU9HoKA7iTZo8l3O9LjNXT+uiMRuS4Fp0R442YuP
in5JD2q8cjPzDQml4dWo5nvVjH88Qs4DbXhsz+v6cm8JzIhKX5gPBRn1z6iuPN16
n5ODwz51U5plMKEGbAD9rJ6lFG2LiO4AJgUfan31TKaCv0alNbFoa+fLa1WINwLZ
6WsmoSMdBdmJDymCbjhydfqKXfgJUOrdvYyrJtsiy11innjbZ8JD1brnNWnLfPsZ
UFCwG81KKezhvpXUvQPGcslT4HqUpI4+YpyzM0rkFVOJ7leJDZI0YvFW30Xi1A15
o+JGrKt1ZmFb4jRKFfOdFYe9gSbSR8S5zFWUdpgZkrGvbKeiGdbvUT8Fd6qvjnc1
U3jhZD954PWITBIZlbFFIr+BhMFIIOMV3UCTVi3hS7P9yOfXIFyWl+6fVLuYjSA4
zwsbpGDSKRn7KZRzIM2vBxdga5zgDnYqcGFjB1I+wjZhVkvJ2txveMpg1Zit8pb7
KnhRFKBc+2IYqn2haSY883SJ+zen9zJY7fHH98hYXiQcqQ+CFonf6LdbtfPe/u0h
6G6KZBquMi/NtkwFSlsEBNv7gcVaTfV68smHFcFJ3tRJS3X6dfLYzrR+Rrgnve2p
/VdceVOx5iIJ0PUChcA23A+trNjXsg40WFEZBYjh8DxHmEbtTxQJScp8paNOAhzc
QcmdwMF/HE5DNHbwaqvDrAKYwxLcYYXj630CUcEcIH7HXnxAUym+2G+NdUk93fjK
DCGGHi850IVV7HrtXg1AjpOEZjgDXSlK4theqTlEJbmRXekKHItHxd+pmnuA3/Wj
cKVfiwT3ravEzwtuILpRcBZbVYh95uHQmyt1bOBQAFHeyV3z79GfDqNgT8Z7jEOh
eclQN86rDIeMnKk0sX/HzyAY4FBocwJ68Kxxm72ashRAAv5PqUVKJ7FyWBFaxflI
VpC8tTBgtgY5J205HEhslh+ffAJb0LV+6cxxE+H49iwdfemvdW7ZJDUVMXjs88Tx
pc6duiWY0GRgNXg9EPDHu6VUoppTZaGfjX+n58WuhOXkillHw/GbHfErFHNn8agR
00SnSKbOYCumpTViqwchhmBuqWRVshyP9HXIctuGxOfIfEdfsMOs9GGbyksfcdgx
g4zvkeQ+AHIerelkrUwNkSAbC/mmTRA1juPwOGKMvh7PKNUwaiOmSjXAk+KZPH1L
CDaU/0+9NQhmM+FuuatraA3X4IVQPGu47NeI02uoh35MtiCSYM0nRQl/jZR02n+P
Tws7fWEi0YASuLd8jLwFr1zCbO3A8HSkVatffMxNd+/7o93M/pMHNScJ7SgjY/Kv
J0JRrhkeiBeKL6u4CH0R1ty0HjPMc05FIyJw27ZLGnsbrYL/ZdME2hkLcNsAdAQu
pXT60RK09eEGmdLm6fDO0gJcOkgsrTYW5DqSczoYbF6KtNCKALQaw1Cch150257t
YAMnwXSHxTF0eCuVIvz3BD15gevMqllvaO455wuiGfkCA1sMl3KqOOdo1DnmqaYb
LrGg8rDvXSa5fovNvB7BlEMqVp9wmGDPERb2dnzj0YhcajqIXZEOzmjf62YHKMxF
5mWU/NkXSNzF9vcNzrcF4vOT5bgvHJFK7Y7sTwevDtY9WrgdeP5Sj4C9zPkAGfXC
w2W6/qUWT5tiifHoX9KRe6K3KXHJZtpB+292cKlBvrVBHwhm47fgLbn/l3wj52rw
T+KmG2ZfP1FdgGwIj15eh0XzAt1VEBDuc+5ksaHBcegjUANR3CIhJEWXEb3Dj21y
I+aOj/Oun9QDMX9zguIqCGWhlBlC4qEkXVUTE+WjjvwaApcYcGYQtuVKzQWUHP1U
AtlsPkwWot1Fd9+qg289ESua65Z4hNsb0ZVZWS+HZLpQ9Z4bsUGnQ2WPnuM8QrCQ
UBAXw7CJ+opcRTqotyAziLJEuIseXpGesImpdGR5MlxpPI+4MIarXJnP0mCjdge7
o0sroJlXBBzCiKV9OqO2Wn6RheZZpNWQm6EbmLmPqdZQ+4PJ4EVj9DKIdDtMYuAU
tj46uYhXQOLC7PiZliAMN0/Go0PCNMp9hHql/0JLMNV/dNLALc7+T7uqHzV9sgX3
IgpdVrxby67RJ7CN9W6H4S8LMIgvDNwoLRcbrAyl9ripCazi9iRVAg3yhQuafiL7
alWaaX3GM/sy20BJI78R9OOJnZG5kdqFJyutdKfSp1K10j6JmfT2WWVzQAUmjgAo
ucx2123Eeisoc/XErOftJ0vgAzHYOviGS+ZREz50daKzguXVrXJzUP/hkBdgK9P1
oKVZPfO/9XpOlC4hx2KCwK2qTsjtfiA8qjfAiCqmfECttxRgCN+5KEnPJigi5N5Q
46WtiCbXtW9g95FaqZk53Ymx3n1f26AzWewp4JrEz9bliX1UMRAj+2qXnMcnXp5X
50WA78ogU+xkFytT9y5l6DYjcAD7Dbot4uPzXq98IvX85RC1MEHp0+3d+Ot6f+jL
BmcJ1mlsy+GT4vptMYl0hAtiZ1Zw0h8vQg7pzUlq2j0XsYlnrJdCqv+c15ssjSrQ
TeFTvkXUnozMMiGaiqxNAuEomOoGHLLWef4TMQsShSkJ2lAYLsfBzcaTznTWCUsa
MldYax48fdShH62TMm732+oErBIwuzvLvMVbCyK6eFlDEHb3ugQadUAiD9bFsp2z
UEEphfi+MrC3R8GBcwbsIdPWh5Qs7hq1ct26CYayJc/na60XR2VIXKq1E0JDHId3
UsrVjUAlPCqewgdkaIHBEgzNk7nvyYmAsyh8JgHOIx1oW+SnBCmKLAL7mMAmZ6NY
dBMsQoOVt6jasVzV8lOLVcPqtEwqMwQvoI4pkBmkqbRFRQ2Pr+DunLD7IzUeQ83o
8NagYJvnc8gnAhHGsGUcPdggQ+mNMcapeadXAIbX3E9g4uDHe1eixYWBqISJ6nsb
UgbfieQXX+B77XdZl3Yc455MGJGiNubTkJIib02d41zmDzfeeaPnl7FeQQ7QR5R5
moeaaZsfag+/95L74ppC8YBBRWA0f5DfNxJ6N2rnlJ6GHi8FfwiDRdGf4dH404Jq
3ZQOHdEqpcaRZUDNy8jZ7+k2lQG4HSoL3zJ0WXWVOC3U7Gj7Xwt3lqxqeTt2iwQ2
dnkV2H8s/KQsKjT4ifXb0tTekYHAFlrlWTgKB8f94Z0maePSid4pOqjh14Qrym+/
uL+/IeafmwayOy5aiD/An/9PR0hKzZCFEu5UpQo149pVP6rwtb1A4IE/EPpKIXSo
J35KXAn4aFIPRH2F1qSeQ68LqQSaJ/WzyHI3sFmiYbz5obWLBRe6r/jag42BWVxx
AbG9CmDEPRM23x5XiQ60ct1RC+ReS+Hm3ICRvEO9to9ULyqtNjHYASeOqc9BL+4S
VNmQF3RiaxW78E0JLhdrNYnoo/MCpcD9pJ2NgAGrsNlv0HLaMUcxhlO4119Spwrk
F97RBLvj9YR3QgDgto+xN9oLq5gWQFNA907LpTuT8slaiG5aXhPIWKUk0mEBW0bI
F1dLGjrFMv+7yR5gdj9DfXR8If1rmq+oCmoBjBdXvRHwrz0Ct0aYU413xY3QvUsd
VLnoxtVr3+53NvTFWrMD+cBC0SCWkPm361a7Og6JwbQNu7i/yaHErS/eUjDBgRq/
61pK4dkqLHlXw7Qwk27DGp7SM/V5PQ82hA1ryx5oIy1bwpSQFnTaw7zpBHE3in4K
kM81WsVxwl7U6UG2JguTH1ZUsBV1pjvnpLKVco4ZSSVotV1RyuzpxmPeZbPBKR/o
9vI2gENQz9ifnwuejQg79HeppDdiBIm5892zGd8Eo1Ob9OkRJzRWZUSLC1dqeIw7
Bz4nxXcOGKDbtUV4x/zu41L1cqNzMS9sCfdPK8V52HNq3s6ObLjAv/omZfm4y8EK
ah2iui70e3LWWQs0GW0+na9OqU63E0MoCwoMJFrepXE/2qNKLEcjtB/d0V6OOR6M
ECUQcOrr+nUTxepPhcutt+Wj07k2+xuGY9WJUMVyJ0eZES7kiKRtKA0ZoxdImdEh
SxJoTvygxBXDbtOeGJ4wnADBpgMLq8H8/SEEfgxLq7TwQqLHuMLjqIIHpe+Q93u3
ZPNhwabikKf1Yu9uRSySkQb9se5BZBFTf4kavJZPAH+zOyS2mZfMV5lRQHJVhtmc
srjhm5PWOuJoL5kuD55UDypVqpekqzzWTtsra8Q/RcZBbl6hmw3P6Xh/HHEXyfVa
XDjUIN0BxfPSHG/ly0CuM7yOrKaAAFPmt/qcGuSNZJeQYciHItcP54nauFBWz7QC
Uy/fVC7BP1YB9R5o8dlEEBVwbIyI1yGpBJvFSWwAIWsYM/mnQ+VwUDjBda8jDMTn
EUIqX2IwSugVXuUFGSWbJ1yHh3oKEHnXswKjv5TCMWRj4ahvyc4BVHz0Jw9QVfyB
WaPU8crUjWlVRRq6609NBJs2RWKwUpmleCkd8iq4yqKtuxB10dt7tTf+DhT+tFuH
i1TpwKap1ABwaxxwdZNJ19PO1aN68EYFkBF3icSV3P3wm6MIge5buzSt2aX5hlQU
dxfvQuZ5Ht9yR9m9kKorbgBNRmFSbNB1H3ZNmsqC9wtT6RIFHY6M5MhgqMu9CVWW
NahjRJkAj+d6W3SQacR8YM3bSXAr0fuGvikOluGN9X3p1vutTn3HyybX6YffQhrW
3Rhx8pd4Qhz9GnzXfsTGnqkmweYHQYwFU7bhMGesJ9osMokd0CQddbfeK9TzNXIf
fznU+F6Vuw5aNsIGn5xMKqspXL+FxNDhdu4UtK4DgzMRQpxMvcCmRv6MFndLAUQB
HCRpuyc4Ma+yK3dXZVlOj3BJkhb1/mbPhXO8CpB6pJHL2syVnKLz5kUbpjNJn5DO
+2ayyXe8w8geDnZJ5W8cs8E6F+0ZACZGMpOYYuXuRA5pCBB5NQoD9vljlviL7m9X
FYQ9q4ZXwCHUmrqwIdFUpRtpV5vkbxelvBIFz7n3/rha3aIBcSkS/Nc930uWsxUd
nXQuPztf6ldeW57ZwNMwW0/7XYUMgF/JfKg1ci+1dzqhhz/jpV5NrDnxiRepWi4b
V2BYxU37u+Exh3MySR9PJua5vy4t494kZIATMYpU/UcwgHaYxoFyLb+r3n9Wsrz1
2uplV3W8BpINfMbgkTZd3EfRoROOVKd0osQMpirthtpriG64X2Jg6Shys118xq3B
n3sNRgGzedSvVnqUprpls9yyY98DIh9PeSDTDxiRNQM6SzhA6zZKbwTptCT5xCba
2JtsbNmDlSoSXO7CMKaj0hZLdUoFeZuNMmlP8snEmvFbxtfdKuMQez3xoN//jDRu
z3bbSFe1s6yZlZDysBbDZaj0Ah9bto/nKuhcMEavc87XInWhMFPIh5DYPCSO/VO4
s4BdTzInQt4w0jVDR48R0t7/mzNNxaJbbBjYt+38tF/qHzbsu1RBZf+zyjkyRajn
Q6fFnlyOelxj+4LE+lexeNS7BbqM9CYc0TfHcALnI1aXgcEnhjtfAWV2549zi4ec
mUzdZR3P/1WK71Dup/xsihwC1Xjdhx/DIeX2H95qdNSs7jsQLyD9TUeTl+REY7Ky
gb/nQiR9/QtiLmr/hI1T7cTWfwtmdfB62soATKF2fOj96XqL2jJdmMsOSxVl3bmD
h0fhb+KH4V6vdjAO3fVsvzpIoii6xOV70KU7BKZ8z1GVRkghlEdcfnT9T8OeBNkH
qaYAsp5IEOpgdgyiQIOHVxk8MYVaF2pE7IpSom3IRV6YAlwcvbzahLnMSr9X2z65
CUDiyANKzMj1FNiChU2SRU8igCOkrTDZeQWb+zg9quOmYBTihgoNfiVkur5QEdKm
LqpgcyktXt3xWRyf+GDXLnqcz2fVjTphmTPabOdxcnpp4EOCRoYOXRvbg5xEPUmz
pjYRh5lvhcdVGxCr66Xzw802K9Z96WFUR4FujxdYKUJf+ufhcNn6mVGGHpnp5Uue
Iz+/PwZsdSseOy6mDhdMUfvUJ1xHgruRWNiKrSA5hMO4DWCsNqQrkVvcmahnZJ8A
IZJMe/6KmiJzCBK7MayCHEUJqcaWukeuYZpKMW7B0OKbcfFqEmdfw28kj7oIeGto
C/BvxOBRzklyG3v67hUOB2cqB/q05RpUB4jlesbwoWqpRSPPYIan1ATu6knn5jML
t/P3fODsZNFgK+of5SV6kDcmzldWDC47AOv3vs8Z3GCI+hnXc0CZXLcnmcKHW8vB
1RM6dzm9YvXNJMbm9A9oQuEChyJgyMtMYfm5R6TOMjCB+UztlSkG7AiuXVIJQtmc
o8zpYpWraXlysRUY1+EzMCtS9bckIvkvrAJQLMCG8WDeD8kO3+bcc0RGeXGiYkWM
61hTW6MR0DBr9zy7x10BO2o4W3Oy/og3zZmAL/x31D+WHCP9Bq90BsYhVJfpgg/h
r3p1cU7XgPzzt0vTkjW3acu3GRXav6Yp4BPuUA1c0kVx9aChKTPsa7vDwAfBXXQf
Py/SgRBx1ScJRijOQ6sLquYGDDjQVjhNi7p2n94QIgmZwjM/YP4ByP0hYhCFkeaF
mVtZYhkNo5XPMiS5e0wEB9UsTgB8qAFPEpX3tV3BRppM0u2YVfy2XZdIQqLnHuvF
U7D52Ie1NoavYajuFnFfDrZOvmENwKAsxU+0/n3NvyUwy1ZiKztEU78L92fpkWeh
eXdlaLku6Ny/cDeu95dLaFtF+OSFN+xYbToReeHOdAO3Oo5RV5fTuEmnWE81Rt8G
f9y4rU08fErTs2ZrZk9etDX4/pULatLh/i9WVCUa5FAhgybSoM86OUwQrSjbkU8s
dukbL88jgxds5t0YXNv4hYfUJQokGn2YYNA487sZwqi/npnSelCdXAGJcJIrd9D1
GOU4gY2t8sDzSKWIHdkmDPcosKJIkInpCMWJrkUZtjwq+x/9OIaqBrUZL2Yhs8oe
f6T3HJpZAU6lYLfjTHGBktu6zWIygI/Qa06S704Ekjg9R8V249I2+Su6OZa6lfGr
6H9HAWsIt8BbV7gIQcc6tG1nE9+q+XVp2KcVKWaygs27dAjOPyLrwYDGgrU5hTo4
lQOHzGu4KLi8irC0tp0dKqjy/qp4bS2TaEiafvicGKDX+XZ21A+OBPEJBgAN6yVi
7AQ2l9S5rI/kIdAsEWedStdJgQE8GqIBFV4WZfE0PtSKaSjhkKtsaZQxLhDNZQjQ
AQNxD8qqDzLIWgaxC5a1eiqcwMImFLK0hpBWNig3TQoSdQjMud6Rx26yx/btbA9j
JTLoYi2YcNpGV7/9WfeNr0HKmZjzzNsqm9obDLrOI7QTYm0w65JgFHqMTa3w/K54
bXFqIj5nw8OaE7NucIKcJ/pKqaCeDCKr67O3miBfeERtyJAZ1NL9IBf+qTAHE+3C
iFX10vxluWJTtA21p2gks7xj2FhAXkbOqLMvFiZ7Y3MvAkDABB3k/EFKnj8JzJpT
WOADCtzfFK43nty5FYTM2LNQ3CW/6h/dXqKXr8k/JTFLJGPogsSH1FEnPBZfXxxr
Y9yRoJ17fIelSiviFOMHgvYqyS38F8JxKl8UgTVW+Dnwto46fHShLn8KPJ1QYI3B
1CoPJbQJElI0jwjaf99m4PToaa6zBIT2m6EJZ4TlSwt++HCcChYdkFanNLjB9mxN
+X8kYXZ1D6QlYryL/aBBGOnu0VKlW9mp8tmjt3s55MhoTtIKnAK4p/L1/MWaoXQt
6rD+ElmQmCCSU/BJngVllOJPwociFoztkv/9skIPsbStxYqNXOQJe7cVAozWXVbJ
F2uh5beUljj0tX0Nx82Il2uQ8jc9R++QDI2B5yI5ZwaUVfay3osJn7Rfnd0AWwuJ
LAYkFXlVALoQPtblL2kimeaYJXDGudsurEQdPPp3k1aGjLFboTEWMbKTGEYtMfyw
f9xNze/hVwo8rKASONVVuYke1jjTtCuPAF7gCWpBJLOGibnUsqqKi9OXPW9mbHic
oe8cvcdEF3uRHqoFsCNvPUiWgrKCSHlwEZNuBhQGZuqy268BDlPyS5gJX7H2YSDc
00tBL/e3d2wVUs86HlkRTtCRVD4zBDWBCAjipcacn+MYeDkpmNi4lz1ZFW/6NOUw
OGn7kMCYbp7MtwhFsXQfBpvU0jmT4uuhxlm8x80GCG25JJy6wIody0p8ZXbqrfR9
UM3T3vRvBcwEnl/8dRyaLx5Vof053lY/j0IfUl5IfnizsoMm9HQnls0aOfXct27M
wWtM2Z/XAt8sFGOD80nXO4J6m4JQgiR+x+ongevr+YlUar5avgLzbqLXL7MiNQq+
mDW9Btugjmb1BmKXQzcJ87FxeoUvoxRploDa1FSH0KozW2cfMkAi44i4l49wyeeq
kGq34sH9IiSVRGkvrFKRotjjLEJzL6b3SM0zuALt1Z5i2M7NW6xVwEH80FyQCH4S
O2OXeqqsUatfMuUZmZVqwtlRJSXooA54h/yImGW3N2lFpgU3c8WCUf6v2X1mC/dP
sGGUAkfxhqvYhHphIpT33CipdSx4ntREd7DFUna/ao38PUN3JsGGVRsJGAEElFnS
wUL2gT8+YRP2a5rDKX450eQQ/kFEDUMdc5UTjeXbnoJMuVS5mYq/FHJ9y+zBsjay
YnYfopJWUpxpxYmxqbb0qsnnzDnpthYZhEgoV6Tt1z10jU+cnWdkdg3QI+wApuoS
+N+tBgN4pyZWxxh2j8hG0O5XMRcMEXmJBIMcdBN12flOFiVolfphL9WIXh/fUNWZ
DzXMhreXyycBKMHUgRSEK+VGZTnZx7EKwfQUr7PskTS51rfnEpi/u8qBWMzH/w9S
pilpFjWlidbfDHATojYoPy2QIyYo38YvZDxGVaxAfIy6xMhuvUnu3JsEf6L2zh4w
dFSGQqKPO9WCjscw9qPvE26JRHp49mUNUzaVIR9ZS63xKZFafqfNhHexjELN0C7x
Vk+GnuJbeo9/pRjLlt9Mpp4d3avq06yS+T7T75kAp/eezrLba4YkGhnQbC2SUZjF
jRX54RERSP0CGCzRE/CvgS2YdrRwmX8GjqY1A9uNV8kldfGZRCqn5HjM89qs1Nc+
yx8TSBj+PR9qVT+Bp4v85zzXrL4UCWicLxY+meXkj1TXU1TrakinIhG6gN9jpC1O
EjqDZhYfMglPzkimKcOFI5YHAbBqT5A7r4d56EKRuY8it/Up8KDaiuGCDoWqBMzB
G3CM3T8etTgm/7kytUxvVnUYWMzniyNgXnYBsoxJ/1KdYbpDeOscFRJwfD9rxWkd
i4HeSx7HHDELnb19nY96gxfLaqpNaS1AeCLwCj6cx9i7IZxz3Y4MKqbsy3lwYG7j
bnLb/9zR6GdrUiikF5uVVrxtChqvm/XXTF1/QWvqkNwztN2NUxMLRbptjGiMZT5c
S5QF/ePgBBJzH+rfD1b13iCxgok6PcJQyeL/pY9kD7cAdz+6Mz4z+Vye6EZw057v
1oZSmn5w45Ik/ATbuOByPxX/wSh1M/gGZlxmpr3o0048RtqmVmOKwyncyqpfYPmu
iUWqQIia0TzzY2ODXYmZG09qdN+Q1zIuixfFC7c2t3234otpIvZ9YBeCkJpkH592
fQMkJgFla/uij0cVqVRR5m0FBmLK/jniTxKJj6qCVoNZZPJL0pgWkP6tevX56ZGf
v7qGJyZW0z/cVYTfnNhH+f+SOgHzDftWwt9rtYswICDFp/xSXGmS+j2n4GtWXml1
rK6pDZH1O7DAxePpNnbZwb2xbhtaZknuVyB3fM0RLjXrVxaEojAdcsIEigqdVVeD
sipm2crGNAFmrBb+lyKAarBgTB0vKOYPB9fUeQFjvtU/FErsOGzwiv2KoyALpBgj
DNdjqb036AY6hPofvladINOjuoRquVKM20tgEpqqJDQ19fBiJ3Cr+yhU0WE+2Wir
byIQJ62QMoZRbO4P+pR14E/3O4NOvoBgWwCosV5B/qmQY2Tw7xgRp9JZ7gvqXR8R
+g6WS0LcaM73xFWNDo+ohru9cGta7izgmupxnGQmLtVv4G88FlLwN0c72aO2khx3
0sKir+pSZRLvHLAD09B5Oi4M7UwZJdxtMWKysHlyA9co19eXgG3pPrW4kUToDDFM
3qs1ym+wB2d+h1X+6jg5aR9PtryOdcsZ8Ia6qFf3SP9mjQbnGpoDjurvgrmYyuVT
vfc9tCdf3eezfKc6Fhez1mIzi11OM7fNg6QKS2ESC4iohIpFhRENyoH7uhdODLG/
if+qJ0Wolt+MLdDVYIOmSjTsm2V+5Xx0RZCGniluTaJD3OfkRWzN2HDiWyAOKRSS
ozCE0x4HHFurdRo3fp3vWPkbjUGnCz7Px/JmvNt1ftIt8P9l7G8iNI5MIE56kQVY
6fjSXBemNHrBuLLJ6KQmk51hn3n+MffWDL3WosD3HSndE7x7tjj/VIwR1ZwN4xZZ
KWvjuDdl1rVeeqI1uUZSegX4Hh/WfTe4tMOFRkO8jEgOcnJBWTCTdVhN49s7mD33
Udfwkbg31V9R9z/tcabWV9kvM3AO0a+ayNOg609H3Lg34A/ffMfS1Hl+1GAF5pZI
Njhn9cUlyz/JpYRscw529R+WfbyBnmnZJFHeVCUoGVo+OfTcteGo1QDMlrSlBZtv
4ICac5m0qqM8IPrAVVFGxwWThQia4CuJ4h1T+0zku9mNkjbB3Vt6sUN/gtwFh8Yb
i6TTOtWqDsTmt/c94xKGasItbjCRHYIzSKXeak419wvMmDOGN2sad5/Pc7oMouEe
vg1QI6o0+Q5tJieop3HOPuWb9gROA7QPZytbCJxcnfMW65tumCV4X/SzOQoAZt1s
1wyVrbD40deSan5YAaTXSdnjk9+C/DPKwK+QrvATHfrQRyxAPDgRMk5GrJycUS82
WhX/RC73F3CUz7+u03p90RbUW06zIfXt0YyiGEDLIQBuuQyiDjTvOJFXtd2ro7y0
tcofP91dFAIk/MQheaqFX9bEl0kgpjD/9aEn6rZIZ41Gt6TeMJF/ni4/AZTljug9
8SIA5c4qT6guoAF+y9ZKAcsoSlKR/Ub8cZ3VMULY3yH946iXopvnlg1JxpfMFLfg
E99So8KYwrZCSEUkRvin4FoRFu8p2zpJmcjNDplfcy8+Lhqi4gh+72CkmeLESa2n
yFPtuccHnTet+onL29Yzt9CPgx1TiKD+QSWQRPpwo2640GE4t4qxZHkTcRQDalZh
yiM5a2fdMSsoxm3BK9zr0VT8OMkzC8fLRJcqh/a3waFWwwCJWX7VwaHXBBs+JnJ5
fZH3Y0Z4MmUKMogn6fW5a4Y+HPxvBOhiv51PGvPj6aaVJjoYIRAV2kn7+VI9JKVj
T4flSsJG88O5f5rT5KdHyBg/FLke68kaRLh6D+HKT1SP1NZ0vxyge0B4VwOQWyaJ
6TpI0RK+LSLRXjvS/ztf/L/ANp1bYwhHSCk25fUHPaanMOEmStzgFVgLl2RPKeHj
4G018YPSI/c1R6JPZHDXvaOFGOrW2IKo2udNljSbHiU4nIJtKRUMqwUUym13Z2gE
a/Wb2ivvfVPiFnHOb/DOC71hBxLzmVyHugnXg18A/ehJL+ZrkzEasfsSS1CQ8YkD
/7u0l2LhSrbr2xtoiJiPynxgnlIWievq6trIYmZPpQcEWvHKB3c6PXPStH0VzGvO
MukL7FNEHXvzOdiwj0ROSMdAtAjMGaG1+O6ZEHVZi7P0vuc34o1IxxdPzCBW+weT
ryOeK42RXmoQW83UU4lASKTrjUkeQSvaZagt4ihRwWalQbhxYVYf8aQ51s0FKS9V
Q+9N8O08LFhGUeySq+xDgUlxa4p8WJkPDp4VJWM1GHsTqaD0aJWgF16PO04JswEN
lYo4TZ/JvuPqZqRmPwpmIwXuS0J/oHl2+F55S7gOvU0PwSxIXO+ULkNDnhZkMY6f
ytgiig/E9lI9hNXLb+/2qkNXTL81DjeSKP/t4fEEPgh1YingIZOHmmRw9bnUUYrH
P8V4MX7/PX5rwhL9Tu9EHXYxJphUJG30ZcMXaCzJvOUEXKqlfFEvUn7M/qexpZ+A
NwyxlzEMAFP8dP1skJ4s/2tgnGh5mUCt3GPH9Bevnsl6UucN0rrTA9o3uKh0HyHw
KX3QEdH0ZR+dc2hsljkJ5gop0HNPE3VYqVZq8wtuaW1Q75Q28c6iF1ZoWjUSYsz6
3yZaK6pvfvvcd0OVkmwD9QRtfE+aY6jM3fxaUz8jC1+4bqYqFKTq26toAflkrFXl
LVmOIBa0jmnBJysfC1U+sluAVxbpv5nfGfnDyddhzobjG7zmfQOFCuIem0vSP23h
z2YK9fWN8r8rhXygSFGDQ6gDMaq19a5TeYetzgu+eAppJ9scq5/IKH92Iuc0jJb3
tuoEku3Tw8LJPcVu/8xQhlLoXDLBf1I2gytfS8943yxvAWViV3yhS+y7qWK81irJ
/HMXpB4tVYNMQSGgZPk/+jiHmgT8B3VX3WRUC0qGZfPRQMB1qe1FGvGt9BuTE95V
kVTTEZS8wTDOYroAs2RznfRLxC3ppwtDuGHfJQYFZNnQd7ZsXCJuOJjnXG49VXE8
tx0RErLKbc8J6sn9fo4eL96kk5L0nCTrCHRYPl3BcnirdcM49U4ds0rZ7tbMTAkG
8rQfkTmwXaY12kzSnZ7D6UuvSfaUhIOb1zWyaGKKVK6BQGWyqIaEYs5xXXnQ/cmz
2U/YLrErIbk58E97V3Y4Hlyq7EhzR2E/UGbwkRdY8/qXDymJYG3sUEl569Zk7IPt
mRnHxQMgB3PzzfgYra4N/Ft2uV9h+2gPXZohpmdPAgR0Bxo/0Amdk1U8b+mG3GnY
AqEny41ZKDo6pn143nXwEp08vFSMtPKoCDqpLY1zpGKe/P+mnwR3ce+1zuDKJQNZ
zNCw3aQAL7s0oGP56Ll+BN7rgbqK4oJqUmUU4kEeDGsmUxamm9S4H87kQaQq/pJl
P26hHDTmyf6oGd9CRDqYC4KUpxP2Ga8qjgE2f3ACjieFptj3/p6/nUkK2YZ65Hya
A7EsTiQ6eUKroWvqx3TH5uJ6a7Mlrxk1PutoT9XABt/808ySPnPrDP42+7F/GjdT
WcCok2SnOiVXYriZBXR+WO6fCVYrrXSgT2wGQuFhRXW5gMsoTK2vcBecvYRnYrOd
wXvbfwEg7xIf3l3abMRqcHW1HN60kIFyzwXvug1+ikGy7pTawBuEV6d8By08r3Wh
lMomLlBlw7Ztt5CYpUaaDwFc9AWqe/3XdybG6NCD53jA7n5r0xrPhF6lm9RddSL/
4C/Gp76WiOQfjyVpVM9ZXjRp1y78yqlM5r5rTPs2I2Qrxwy6WnOA33eeIC1C21MV
H9IqARwq4+plNN1osNKtAcSTrsX0/nxQnocQglwt9RnOcrOjHLOj2yfxqgUgd2t5
d/m7si3NiwIrdx9AakwZ4NlxFVk54KQOxeh7S5sclmL5BMQDPLflUU9GAJ8EADE5
SN5DttLhLkaMTjbfyWNexCVME4OJPDATwE2utok4Cm1vSloCRuO4tNbuWYfaOpdg
W4k0Rp9J/jbCrQM9YvWhpN+Yfaqxjro/zLxVsEeytb9Unx7YCsFYa9IJDu5/KbXo
DIbbmJOalEsXPi8I6SXj6RnWJNOxC2DzFT2pjkyTPZ//WEE8i0T1xiywP1rD74iN
e++l8isscYDsuz/lmmxUeEcJfzjAvxGJzALwu5axIBeX5yUlhNUthX4vD0RhrTHj
i3+o9iCBvj74lUrIWYKMo5uzqvxxoeUNq3YErIKdUDTuBSck0U4FtYdiZfQ/qkE3
VvZ7JkOZfq0LxzqlDelB0V6IDwfPkwyI6dAKii/NXqq/N6010vjZdbCVKmvdB7Yb
dCkfGDKtuP1PonW6LvMadJGVXXmzns55ykV28x2XG+z+Okz/P/nFqA8AyJPUramo
E+4qks5/CaTgIrco4e1RcK49c+AFFhlTb1oTZ2Dv3qUTnDbBzaEqIHv29iU4rRkX
/4u3eg/Phb7+Z35XHRvfT/ukxzrxgx4GlA84KN3N3cYXkUHnZ02ce0ESJrbyDT6R
LwZMLFcLh+JmGQ8S0nXOCOOhxtvP+iF/uTeroq0owZioNeM6QYv5GgGwyceW7ztV
RcR5Jw0seHmNvln/LxxHaRqFWReVm3AAnJolIJsOq+0thjIl23S8f30J+8lvOZ2K
+a/XScc/yYyqMVaRCf8N4jzNqnyP0/1OjMuX1aPmTmaaDV8nixo3qTANQTgx+lF6
0e/1APRqFIxvp01O6FlAGg+DlQk3TqryOpaPpqI1IPoZxxU48+QE3wQyrceHCG2s
NhaNi68sbdnR1QBVU+9GoQVyXXj0gZcS0F0olSTE4OI=
`protect END_PROTECTED
