`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9TG7VuVXNZMQyYNpiLKK1OpIwZRkxB6SynNNN4WaQRLs2CCwIwc8hLGtkOmfigu
n20OuW3SobZEPBjvKO5nd1Nr3AayeHb6Oe72PObyDD6GWYuDgA6ZSfco8R1KMpe2
2IyiAutpXV7rDXg8nj9FSp54QjOqNBUEfQPvdpME0dEK6nMkAc75FYiuV6ZmvcAe
7RoWLRSqiTTZ8g48VGyE7vAwv8uWijAiQQBE5XNv+1c8DFSTKV+M8F+Q62vKt1EX
ZGeH0PJXqjyEXFoE02CUSSN2oe70EwfNKeOogMsMamU/D/K+IIRzSrb//XiDrQDb
Q2lVf3cj3O3XsPDG3rIzhNYrrMFkR+THPjGLSqre8UlNv9RrcgKJryTyCYMPWLIf
jQK9YHnAng/Xdp2WrHTt3s2+W23rwwWhYtGtI6TTWQ+xebcrvTYLp9FNNwduJ4K+
Y7mvdsLfxHM5jAADO2mA9DWf2boOIr/h9YR7oKTqj/6pDk+E6C6h2StUycQpxhaa
jSTBJ8fBAoQuSvsyJ5elwMXoLVkDkqYfUt2NmLNmczA8gUAAqJ96MnEF72TCMzE+
Z1ewNZaOofWh+QwkKgTTdlBdW1fdtowtgR3K+gIKQXPrTdFcUVpM4Ysnt8iExNMg
uueaM34+0+P3x6ZUjKAOozKTxSAa6XT4eSsT0kWQLcZGzLSdkLVxzIpDXW7palfD
4T03poQYqrnDilgAhY5CYQiusi/yweSS8HqBU4pfkunGcf8DsPzRtou18fd9kN3O
cSNZDH2Or+kqqWrAHa1rZTJVG3alXq9hfyzMZ/Lu3oCtmobu7OL8flNo7Bqgkyjb
E8pUXyplq1M7kt3vUNuXBZTljzr2Tzw9fCbFbcZnQPFELz0F8gTTj2jKcJOq95f6
ahz44bvpmuHWWaex9Dl71gUxDOzjodcY0DMpy6YNMt6xTUbK3g2HIUN/Pzxz+6qM
TaFtEwsibej+Udb/MYvh/1PCvczmpQpO3kpKdgndr0iiOPKYizIrpuxDsIxS/cih
6xEfxpBmGwwlFfmbEEui8EmZqvNldeYR4BGd4PXgbG7GGSmAEoi5iACserRun2/Y
+hByItHF4eXvd/8XzvZahVXZ6EB5nrytoi0vH7ZusZIq8Pq3+zJGVg8wLARz7wlF
htQQ6uQnRo18wK0jW5APBBOB3VXB3vK1X3lBgaksOx+TOctCGi9HfrGGxndgor7i
fn3GgBm3DDz2q8Dx7GeGP6QgFYAzWGklqV2nNLrQi5w8YMIWbjoiTEW/PR6WqIj6
ipKy8SkqrfWU7Dyat9DWtJNAhLxuONNK/yaIWq+a947NeiT/ZWJ9lne+yT2gbU3o
ao2Fr2tP/CZ7+LQqhSiN487PStcqTszfgZKtbqvy4AacMcedS0btRY2THL3bzBFH
khjg00jWYttWm/w1Lmm0S8FNNBUG+uoJ6WNq+zw2wshsvET/MRu3oCVY8eGfeIVn
LZkgUG/kgbmnfkdbfDejhxFesvOrgWtvZPUz5dXm7boMBe8RbtLp53llrmm5RGnX
5XzvhJJZrLspHv+EfF84vRorHFAtNqytMtPYnUjyU4iRr5QRVkW5I69uZ4Sej2ed
DMQaNl9S2rQJbfGZ+Zp0iW59BUU6jr9TMJ0WMZlME+BeBeGXuN6mtVKItRWgTE87
Zp5qzsC/tHxEWdpNHXbVyUm/MALaZUs+lBaownigjnU8M1fPrOHmDgWOgpMvL6hn
PMFMV2sZt+QCaiVb8xw3OeDfgmhvsNGQ/1Gsh0uY/fmmLXPSgXBPntqrnziHe5D2
DLRlO4KdNAGXc2tLCYDTJjQvXjr97tDhpsDHPyWT/OELPEs7f3b72BayXHW6qoss
amhuwbrBCzab87ZvDCqkgkAT35awfQzDVmc58Q18iEq2kkrFX9LPrpfgfR9USrMe
THg8Ekl8dOYgVwQYHn5HS0tVO1Uojo+gV4a1V3lesAtkB/EGpqAvpNKdTRwQ1iwZ
uXw6On0gHmK4Ahlsk5StEsI5c8TOE+DSxhxk0Pk3zDo+NMwxGNEE612LIvEziPIk
cd4V7L2BmCvz7iUHihvlKtl783gCZSPvnliI/gn706m4GZI81Er2WkO88CpC4AB4
+JnqJSOi72XVr5cV5zNB0tDOmoWICcagMS5OeE/8XvkU4a5pcLwO1wp3qRYmpWab
o9jsg5E9RiCMkw879pDKNxtFGu0/CbnQuvmJN+CbDlrD223JSGzYiysTTLHSO8Yr
4qQGK9mHcWaYTfuvyfjRANkPDsdvq/SDmyUKCofckfOi5uHQZ8mD9a+scz/lYV/6
Wh4T8STUXJIsdWYv8UruUNv+cfgTU/P9LFpnEvTM+yFcV7VR3PyIts2TmSkPJXo4
1FBtvbrBZI4wzgakDehEvHb0lzasqeNvuw/Epkn0OztTT4qkhGlWZaOdgb5xdWbj
VLkCwkoZAVRNdZdzotE7XzSuOdZLPSAPxzx4CVmE2mxF1CFVOzmYDm6MeTpMv1kU
+N8AenxhLiCNIujG6zENy1wTVkW8hRiVd5TQrYOsHSgaUfMGa4jiwdTAa8C3mTbM
ua207QJAKW2V6JM8FXPjVN6cjFuH5iOZl9GSSGVmnwrfivr8KcGWiNmCvda6grSE
VwcZBzc9c6fmKbIqYbYZaDJ/xDuGLHDvzIgRTMCTWeqFPQTKH7K+duAOD4fqrvYq
u+w7bDBdfN/y8DKdJk+U5RS5c6LP9SaNZ4ej29wRhW9jdVg9N/6R9uPOnvgoRLMm
2nRK+N2GICH+FSSsH7mkCf5HjT+oZ2DuwUvxpSVHcX566F2Kvir47jiRgOQHgDNS
sye7DC1hALfy3tDXrCGQ2OrkyMCbOVySuMiN28cSLqAzs2aRKXyXDYr2SHe7mxil
+/5q1AmD965vlyHAs0sy0Lq6/32HkuEKzdWUsluZvF2WTenTfglXMyOzBgUjXcYE
a8fo3hQojeiu5l2LEzt81MDP5LGBJ+Tz51nuPc+6qTGqDV6/D7c/YQuPgwDR9qTL
iFn9GOGV7Cj6BnG21m23hHtaKTmU3jPPPL7lTKUfnmZkbpoh4Fj35pUgCOje7Diw
9q33ZHOs1XE53jOkcMcfD6gOUxiFL6XaMX1exoOfT0EjjEKAIyg1xd9R3xX9mQOs
13KEXWdk8vvBM+FFcutGdf4Wwr7ZrJV66LnIuYNod5wncX3foyflh5q/Q74jNBdE
se686Fw4jPq8cfuinOEfMf03OOZZyzH2XpC8/xQUb5CD/YNMb9hhILoHrD5jMX3t
vnl/ZLDfwBF5YEwSWoq+lyM4P2WHP+CV8Oo2Wfh+71BI8lQzif9s4zTyI/hJSXD9
Rp6y1UJUbaq3nuwontxnP3VJKuNeXwHgnXC7aI4d8fnmDIqA53SdV1LstUaYjvn7
OOO9lxKirlirJyxxwI1FA8jYOxawb4NCOlvtVNrMk3YFiBmqM3J2As2d1AkWzjFr
K98zbHa4prZKU1RmamhtMP5rNlNpAmsz+Ph/koQ/589w1z5lt2uthOXl1SuTp8Rl
R2IlKsz6ZTRZMMfkD6ne3cyaqEKOc6HOHnBuQqUK3Zhdqb+E/fn6mWYodI09OqRV
54g0QDCnadSE+gMrIW8WDb+J0WFkngdaJxCp+WCSR3fRNmWDzomHf2MUnLv0izF9
UJt015vw0Bz7XSBy3uEfpIIbDpX7+pZ63F5wf7um5fyjOtSOxbi299HIql5bjqeu
vPBzbhHfCgYgQIJc0QjIxT1S8CUphQXilZpgTrbeeB5vrN9rEWvp/V6oyC/6ixZr
9A+KSHytYwoboqRskBxT0GoF47POPaBkh67mugLuXKvpNQQ4jXEnlmGbGAtEkEar
YyiSymoCUZuT5Syd8t5Ltgkh4AWhacIPPZ5C2lnpMYPdRPz2d5+RsZu81gNBbupr
SjST3xrTOGapqOI918YNR4pveqN0zjwNWacBXUdWt2EfUWkxbVDwIotBLdcMTJtw
FjpIdvuv2ZSLXlO4ZK1d/tBSpYmlGjCxPYkB32g+D5BXC/Psv3y7VTIuf8la1ewq
l2J7AbgvC6LfKAAmzsgVkC3j1zFt/UxrdBFs/NXSfqbloSUmVQcC+j8PNWapaS3W
Z3ecc1k1I6uxetfMhBli7Uw3WDxbngkY1/JrC9nctTztJhD2x8fI7KSPlLWz2prY
r/AU4woj7nuohD1hr+jU600KpwHFCzNH/EAqAUM/JT/txFaCPWkKab+2FnyAS9Vp
8lBWp3aSj8T54+ts10MVoZZS5CyrDEx3zaT0U3oUlnx6KgjOG1pm7FkNWmUdXOvw
jvWtnO9leK+nUf/y2a1nRHRDtXQ+lC06NIvqVcdVJiaT7+zopePXMVlVn6O2S/q2
yp5MymKgcsiRrf8Vy63AIyYRsYZ+/pYT6IyEWWVPUChibpsrn0Q/G7BC0V2E9R9a
b9fgqKZCdU8TE/tERap3LGxJzZ/aKh+dyRgLf8TbChy85ByX8wItd2it94NbzAXm
KIeM1GCWmDl45pDHhGyK+uWzabAd9Rw/qQxee3Tz/g/pBXexbceuFCZjQtpU+Kl2
RE6A6QF5FpjYc02/4oEMKORc+Imt//yukBi8ChDhJfefITAyuf1uKrbaWZIsAlH1
XAyXJO0+jlunwPJ4U4wBhMcu4Q4VDdpecST2YUN21hRx0xuvq9LiW2pQKLjCmnnb
EXP2CHlVQfdjl5YB4EZQBvMPt9aCz3ouWokzBcxz2x+MBBQ8XWYfcHh4vkMFH5cW
BYMkxGNBpCxbZAfGKXkqnS6/fOAONy/YqB1FZnMcfWp9DZKsBB+oJTIIch+ZqZqi
gmhKmaeKwla8YA8SmHToZBAbz68fSIYM65UZpKH9BTl8q4pWyezZyVkoO+jKIwCt
Wb/W72rjEXhwZNXMqqn+EZQOkFY/2idJDW1lLgLJAw2Q1UWl/J5e9M7qttQgMywZ
mGMUaGC6gxKCKLUKQ5ryG0Gko/gHLcqJsiI8SJ8Atg+I26eLZeh4M9H7PODelMk8
0GTm+5tiUySulh4eIc/KoBx3sbGPVXv10OVBKOOL4o9khd+ogX5JMRZ0bVs2yD8n
plmCFJJezdn2N12qFlhcuu93WG++Ri7Sx6QVDbBmBzGgB19GQnlPqAZVSepjdKmd
jCqIm6Y3iSbcQVYD+CkkBI7RKftHkSo/hP++buqcQW/r/Lb3zJSLNf8cinb25Z51
+0puDQNWQhW1nP06xz3W5DOcL4sICdKVCOV9ElS4zHLtnWJKa+8Ub+/gVxwNaEzs
Vc3qIMDbhOKqVCE2dmEZpehCcRu3rniQ5axPGQXAgNf0qpqebokbEriaN13DZp7Z
OhHbQOJHp+TK9IibqHIli2GJ4koDtO3oNBCxoXaYYwQTWLkiLw/4cZ9YRnZsceI/
oFo3N5JsUz1haiE4OuGceA9TNJTvr6pdobkRZ8QoY/OOWSTSsNhTlLZuC0MPxmsj
O6lTquoXVrhzcQ7t/Q9JEo3GhQHcYDUxDtyVCfopbraU1o4O2f6Qvq88RB3CRkRp
LP7riFvQzNwxiDhr3e+9BkWRMSyBZF7zRzvOcK7TQmtTLqUXpRMxqy6YHNZqZnGj
J7Sk9U1l8rTCgDqneEYCbbCF97Pcv1PaopEQAOfIZu3POMADTFw+U/atWxupYeqs
3p8119PlVkz1CWFKwNwAG+AumKmVY94gzG+zP7cCgFppqCDRJi0jrTiYftWJGlJ2
PBu6tkI4qSz5xYHAwsj7zVB9cXdxLgoiEWlhCA2X9kDbTfFoPPK1X9y/aPYbGZb2
c5JBR4HyzoyQlGAU7L9IG3aEQGL518yhBmGtwJjTVnIlWgj8g5jbqCqN+Kc0cKi1
5s+Ctpch8UFkn6yDJX76JLaw/Poc85Ep5JNuwbVzg4OmyTHT39RD7bCznbA/3fR0
Yoj3hPR0m1CdHADNOsWCZ6sSN8iwUQ0sjdZZr4WyPs/Ufa2RbLukfd84Yz5OhukC
LWLI0lgKXT6tuma0VIX39Odl1I+/I+QbBrhe6/X9M2lpz4F0U2jgr0y0yIL16Uhr
iRv9g20YCFGPwuvaoaBCj1rWV0tTTvTuunJCb9crN3pAuTcyWFnRxb75KZtSyOoO
XvmuPU8VnYwPSvBJUx/NthihZ4hP3HCyVVdygE0numD9JLr88228dX3q5XELfQ3A
9pfvfk++9miCCpiXbLgFjDk4nc0ENB5bYaNqfEiWjYKM72ULaTdX1gCZROOGtjZg
grQq5S7gnPnEtJvzDKKBqxKeK5klFMiS/l1mdtncLvv/gWhWOMBK3APPogk4cyIK
9hUj77CPDADUyXs2zcd3y72kdSTag+1WgB7EKSIxjCrg0Rmac81AkMfrN0ZV38vZ
cGfFOXu8yovumC0zf3tbiQGyv1z5kPwBh5dvDcYThJk8viR4i1kqG1DxrwaE8plt
HD2ccoQxmGrUcdmIyMI15ahO+Y2PS63noMTLFOtrx/jfXprIAwIo1bzyn909Uk+l
UiTJt8XnEVAr/xEXf5wsTawBNpsZlJez+0+ywWENX3gBReQnbXLPcBv78hTHfGJ8
Tt4vHb7iGPQDMt+7R4+ay7bQ/MhlZfv9j+AMXQevlF9HDj2ci2ATILu2n4hK52Js
r2fw65fJ5mTrm5lRAKsoC8b/vZFM6linZ4Hn4/EDkuCeZoEOJRH9qHvE6uvWCujO
uu8roZU8ckoXXgfFRHmkwNERDtTKJvcK4o4KIptcyH8p2yjqjLYtehsy61a2Z/ny
IEoQVl2izeM4CHs0+eFVoWiRIcUSDZm5beQun89XkTMWsHHX8ijrcxRw1KaVAdHB
DIIlKmprlRodV5S3sp83i8Ycccxt0oWjFk+yx7YD4lCwnKqBhO6wHEjGpoabKHnj
biXUxlSMVLH/LvMEm/JAH4rySveoNcNJPvVJicoEbqIPiLBupG5YH3JgV0tVy4Pd
OAe7sMALyog9iRk94AJtVWPRKaNhpWu85V5VGtJ0k/K4UPfm7D9ef+yU0S64MtRX
WamgSzkRxmdt7ehx8gfCl/v0JUN4FDcT1l9n6xg8rKutXhvEO0GNMbbi+YyY5mFM
d66tliwaGjW/30f6XFeXdbr8faCXNi99h/lZjeGWETQ1Q80cBMMUGBiAaeWpcRAb
xk4FwGi0H1IMaOp4FVXpvs7tp2KxXfpyKvtmMRzp7YBxaSoLFLiRdMfFIFGjvtib
xs0Na+mFT8JlT5p9F5OOL5ET0OHXSBKZXJaS3wT/11uC6wYnRieHEKcQAovF0fA2
TJrPZ772we18d9kx5EDyJ72/YYr/TOM6KFdjc0vOQKR7nqi1EyZGDpGBAy5ALmFc
8j37qRSBwv8gUH7mHobV+TMFSvVebYmU8wMPIMFSNFn7+I/ectVabbT6lcZZmBRe
UCJkmB8F+mwdvMKdRV9WYVNjsBK1P3ArO+ph+/ehvUiBf7zr8kTd4NtbgaFp8tkQ
JsWPg3Tc7cMhm8TiJnjB191dwUUdqEvQSvg2pYbr1uuwvTZfGTgimi1z5BdIkPmp
AK1Q8/ROweGCCwOhtJTzU48qATMdKRf42xhrt6INQc6/oceUW0Gf1Vv+zU2avbvR
f8JbN85eG2zj6hFz31L25U/hEipilIdAFuDTt9SlxgrRbKnPf8rw7yVZWI3NhhWg
9PS2AwQxEBUaTj0+uRNJc0Jj7T+A7WYbbEdWozY/nJs0eg++99Uzly9fLhQAcDhX
iCVnL2aMdGBCdGA5wzcIkcxpUCMrgzQgClq8EZ5x28toqcoaS4XsGQljNAgphFRl
qqZA/Mr+hWLTRY5AexPrgNWRdy9gxanZ4+tJkSfsDxWkuTUSx/pkad+uYyrNU0K3
xHAkyQqZjoIPFAqMBkNpKSPgRIFD23CgkVFs81vlWqJCiOi4u1rIngCWSWPWSuD1
9AsU8LU/4lowaHrFyVe23o90NoiitCGkz8Jy/UBvMFOrwS4bkwBBkr3JZhkrBxVp
aOvpVxDX3Ti2pbAp5S3VGhkCC2VER7u3zdhEXVcGWZlFRy2FET5OJF7SsN6lrQuP
FbmmY9mvuuzUVYRaJKcsyO9I2KHDmf5T0Cv2sUfPnCFGGCGH3L6NptPLa3riCsic
kdRAgZA4YaU+xejCqONFSZlSLA5ejtIzxVL2PzsXMrkupH5rUsWzxkYs8Zmlj/MO
SIdwu35k9HQYnf4vq/WIyqEuSwjRrGbcZoNuMFQKGSAHTpx3EPfWZm594ZkuQ9+U
XWR3DndNKKZ8Y86sqSyHaT9SpYzsvzEwI62+BTYe90dhLWQF6XL/Ew08Ow4VMjw0
dV5WDcxsR8X5ScI7fjni46n8rP58tPWvJgMKO3oQVtZPxT+P+Uc03U9FSgERO2VX
TwqNt4EI8Dx4VH/aBY5Kq5eK1ap2xCdc3nFdO13+zIhU6f8MjI86tr/nhPHMZC8w
aSrIEuwdGk5rAaeKNtzpKM7Ewder0HCX88rWYjcYsLf519D2RCp9FutOBGncqaKW
CB60lwc6P0x5aC+Ajn/a7QDNo7pTKcATPdeG6GRY/DNiYSHsWUCZPxly1GtO3ZQz
dTfIqZOlLvTIq90CnuKhZ+9e5E3MJlKfF6HDvwH2TszEENjyrgqxcyiDD/q77ZHe
+lwlKWy5O6T0le0vtmEOX6vZJNCDSfmP+FMeD+qqI+RmVZHdwecxXHftEr56SXWQ
ve8akezSf2RFTBPMD1BV2pbE117B/D0QXV8YhSv6XN1UPkHNO2DMG9+FBTG0KA4n
SqO64eTmNTbdoqvMWj7YrOANRmiOCKa1xlCSlpwq0ZLHtmIEgtWtMft+YE/ZaDPx
Wms+Lbk7HBKaDqgjNjzSA21pHiTzOnEtumYaS9x59P+/MJVYpG2r6H8uaEXlek4T
qAHMaU4e+iqX7pwlwePdXdAmCR5z3gNjRvVv32qNt5Ir+L3OUwZhrSKX7HcZCEPX
bFlccH+0bJ3ccaDASwUttg2/7IhhsJirQSwfPv9Yy4fmioHMDlfGHf2oA789A3u3
WDmUyFH0kcINkOBj04i4SXsssmLJ2yZLqBfRdkt0EnnZ3pGs5JuMtuYo3rbT7x2t
yeDt55+Odz690SgpX4sPJEnAgNm+gE3p+i5pjAy5F3RVdq2F98Gm5706h52wtgy3
PmWp7ls18qpz/QJZMbqdbx06KEgv9/ACOs0JvbNhV2dFdJ0qF8Tl2qcKq5405Hsy
Gjy3qgrp6XFp9wcxQa6OT2iYppGm4Q9eoDZeypu1hZ3nqpJuw4x8lrJw/5s0QLnW
bBEh/C2OfRKWQNJC+gj95cRcd89Y1VMMKqyzNqvTY6YEF4D2KuLdf0Ss2PRZfIRq
vPo0LM+G0Yg2JSS/23xg3EN0YxQYEiNWqOeS4S3g2e80XdTOFDEHIOOqDJel4H2P
5SD5MRJ2Qg8AtIiEJK9YOSVEtiFnjaOd5cA5rT4ZMixRDyc2mchH6j3QOqWYXGDd
7LWXNI1Tcz9Re2IduI+xKArfaXQEGWqVP2GYCzAjGYn9681DMYJeMQ0zzmw5lPpm
GiBrls2TPIGjjoGmFPYQMvt+ZRoMzwXvKzzrrtGS5McjgfxDSa7UXtgvC9UXmhXB
Jmm5qlDCH6ROJm/brWiNUjerkbw7/aMjwquoY3M7KwdpuiZ8XlCMJAGIBCD/e6+2
VCjKaFtmce2i7By2Tc4abLkFiHryhDMCpOzpFIZIySlqq1iHZsiiAS/8ZBj+aI0k
Tct5fZJmqWdML8egqO6mk9t5wlF7sXKn8/qLle0LtQPSENgF036U5tl52g5I3fw7
JB8NVTV9qyUtl8jyXH+5LvOSN4KZ30DOHGyR+dU1y84QhUrafbvgf/5Dj9kTaPGh
BrJzGDyT5mOypGDgOFAI0y9zAW3yFXew0r64aujyyINikM9IzRKfNVjegK0u8GVx
Nh5c9LxWO8htkotyMT3nD23Dn1LmsX+2Dqv8y6EZxtBd/4d2i+rl5HGx5STL8Uyt
6iVnGIQGHXi4HF5ZE2MPs+ZDnkUEVi6T0qZOjiihoEEDvRS9RiyH2DeNodPoF5rN
+uP1g2gtBZcI+znNiWJTBWwRwvIssvFlnchW7ptOJs4so3FKzqgfDGJ78WB1eF6y
//djfPdlYFSESdpHoCcuDhKufcwujNeQc1Ug0uJAcIDj6CBVOXsTvasB1pTOPOZ5
3N3zseiF92Z/S6f3OK2mEF6ENYRHs9mOfz5Yt6Lxm8vOuPWhnlyUodu14okhHbFc
3dti2U9JiRfQsbLrxZY849w5zQs2wZhCQHTL5omvRkYWWzMcLOFYGG7jS7jVlHv3
b2dbZCFIzwfr6ti2x6HOc7lYl1Ba0q1erl4vkDYDDFm/Yrd3Fo/MUz7iaI5VYc9W
sBrBppMk7kAYTWV3echUU2qrtX91b+JE9JHI0/seif5WHcMhhxi2DVSB1GW9SQmG
yiziPFsMDq4hVdG6vrpo6IHstTctbNOcFC8dzi6l6BpNl68IwAtvLcEuSX5ozclj
iW/ZdVaaO8mLV8aso2y/oCrUn9zZXoLqmQWHajXk9huQgkqpKG1eV1KE1FW0R7j6
rt2KxGv9llvQSETbO3KWB39hihBRq6cFK0C9NaVtBqXgvED+6SnyrdTdbA/Cqbu2
/GTXerIzdP6ozWh/j0Zpn187SLajhjDc6MVUWo9y+5hCRYV+Qdahhnp9O5CZS3sv
JIHF9rG5aF0WrtOP1PF68OCQ6+9ybbHkGXNxxemxko0b+yJqHKJlyKShlRqvHTOc
1W3VybUpXRsU0ScxE5NXh3dAjt6Nv4zFLHlRsO6omD0zLnNVFO36YHHi+AqieiS/
OkJui7RJg3KRLtGBrXRc8Pi/AkzRQjWgM63CYEjpouT/JQdVhkMjY3LxK+8AkoJ3
vMjDPdEKoL1i9aN5ZVEY7JXzwaIPCz/bq3tk+IU5GQkWRBlSC9Dmz9bQfgQZnoUw
Fh/dFeKPaiDN/ahhXk1JdD1dWznF07hNRRnaLHprsrrG0TDPEsglZudEDzn4/Obn
QNLsy1k22vamqr9qTLcQ4xEcc10w8q3RHVqO1RJYIaZuaMiykC7AmJlroMIYbECA
66Tv7DVF4B8XqhnX1w2L3RentG5ugFtTz+2oU/1J5MqWCXScbwGWh/e7ULxho8zj
byZo6kC80QG/8PLS2sfwtsd1kJAMI9INfsMr/z4PTrtyNaouNoaIhZqTbhk583mK
BZhakOq+5OwTWmN7CQxiVDJ/bDKNYNVrBPpXeh9LZ4zTU7//Qm9+8TjvUlx6jZRR
W++4IQBr0suC+cM2fAmz8QbXXRGHOjp/75bopGc4vXTEdZs4xOdjD2eOSnXl/umF
ZmtT+khpgw3hUOEQ54EGDpnEIkVZNitW+EU4XudmkRvzlvHrn08OQTKS0yRwosnh
IbOWnq5WFiyYmt9hnU6PvmyvA18CMnkxp+PPg+QrnBNuvBRT1mfP44NJ5DEqcJiS
ShP//CsIHMStjFhyVj1RgZtNLRjp90x/8ThBYOplljx9o8oSBGWo2DvVNz5DQOWR
iA+WqaEG27VMTqwFLDhgCQ/4FZTlkYb+UGRlAzbF3wxRD2z0C+8gEqpo33kAWdnk
jnuDifznz8YX8fGlZGji6kgXjGZxl0yBq+QsxQoTxrRGnWV/cv9rfMY/ZsF+Vay0
wtSOhOrI5zPaMd/v9Eaua0D/5aqyVLtBBU4gIaM88mSPzTVmAg4U6/oUIS2zi71c
9Lt9uV/f8ruI9jCxbNGLyeJAXjS7le83IF7JQqPk4W/L6QLPUq7VMeCCV1nbrh1S
IDR8TdGzd3f4u33ezVgi7OMoUva1tFhH+7Tj+uKa1jpSkat9rfq4xGh+ONWK9YHp
j1NZ2+bT0D/QGdi0skxs0P9yLSzi5VIfEIs9FV0eD0HUG3pOXESpgDwcbo4VjR0V
ydxuFi8z+/zYBIfvA4DghCHtOUjm7GHP7eueo9bH0i9+bxXCSYNe6Y/jKPoYPkDF
VY9Mf1rY3kGepAJlePm5AwBpwTNM+Veidz/jnn8ewDjeB4r2T/f5hk2abOO8pyzq
jyDH71hWhvoItQWVnrUfo7cXo0xodIsPJMbFugWyAlaiFU7NsU/sxpIB5uYr58KG
Uy1Bob2mgn5pU8lKh+HmDFayduOZ5+r6EAYJNwr6dxJ0rDfepO01NCANcFZGWCs7
+Ut7MF+/xd1QSo9Jbk/SzngZcXMvbCwGpVKC+Xy4K/Ee3kzm4L0DcL0kHffvMva1
/MPoXa/CxXcUXFaDXKKodjHVTiNjrfyA9N9b0f9+iYU6m1kiJuZjfh8s+FsPy3iF
eDg80Ovy2j8F/VWjwwM0ObcL0CKGJYh0Rdb0YCG+LseOSDfVf9trJjQcK5lyLtDU
NPyRf/b2M7AtNc+mvEXcOhTGN06BqmjcctFsNL5mBVobGeaqbtvs2upWghV7efCo
S4RhafOVKJjRE/ioTOLJsRu3qj0siqdJ710loBaPbSG/GXqzWKiTJhO4HCH7L5Sl
Vj3VsEhHW5cC7AAcwQfvLczQgy/qxIwqp5i7DfNg4n41zmeTKpKKAMhj8RzBDfoG
mW5xWjK6PxZXEVCRYpo4b/cCbChjs0yEXSIijMx8n+7u88qDnV49G0TDpDPj8hr4
T761PB25/k968jwcRXJskNGqtVIA9zzHOuBi8PdpnNegG4u1tOPQC0M49+4WkwqU
cHYkgJ3Zkbf5CmDaQifZJIcwzSZnEGJ2Ad5YSl6I2l1t9NnA09YHUXNcUjm3MqGb
nmleyKyFEsWHaVzYZgx8rzJ5Q8aM54jHwHUzo2wzm5QM6vUalMdwsaD1qet8axUU
VGd2xFztstduy4N/d3R9I2h1BAgjAXYPbkuuCLr5Vds9nbaP1EBGcSObMC4akzhl
Wc5+tqvcHduZaohjmRjm+G0XA56UqOommUEC9exWnie4+fGWCn2sVMl5+CQTamAo
z/Q5W6Na/2UDHIxEQo9sxERk3m6J6WHQ4GeduKOMTnjYxBWEnV2saBy2Ol+eMudW
BU8C4ri1xDsLa0g8VRRai0vxJ2UriOMyCVjmlvbv0ETLuOWf9XyR1t1VSmcUnTAT
j8jX8zuYTaZOgJUIx2wrLWLRSqs9+L0pmSj9qii+a5VscvGo0f2g3eilXhBoUKMq
giRNt9Fekx74lQ5JXxf2/GD0ehmRA7UoJbs8bxc+vnoQxSGL3GvISKn72Yg4PxGU
5s2zl3VK0Va6YuG5eeXdZ4ca8MG0Lx3LAChTwt6an2fW+1YjG2H0mALEqEu3E7rS
NeLuWf7eIutfaMmDmWk/P+O3ZzzeXNp3bhqmGTMa8hAxiBrYX1DInHy9aYyc8/yi
vQGd8u+RjqcorpX5qWen1YfNnUw5XWm/Qam07Tg7uH2Tcxss408S0PvgkScDwgHr
mY+2oLSbMIqJ9MGvvXfdj/ep139aZYQXbwiArIFQYtfSMxYfYw7zJYZqen/58BDg
3q6a/w41xsmVssBrrMqD/YBjt33wpUhnf5LIH6mbrxGH7R4LQE3r1f0iSUGTpO3j
cw8mBWQwu1T124q1+ErbsjqLSc1mOABEah9sAlxKw91AkbY4tx+Gcliafw0bbjOa
E2yCm/5R9sb9hxH7IZM/+eCKhtgABfsWNQmn7GQKU1CTJOLz9MAm0Dru9T1C/o0U
MZ0fM0y1YSHkDUDSF1MpUiv1PLUw4QmAt4HbJhKdJtB/qc2PBkPVfXvtsqqAhFr1
01nGp/8AFt9KAQkXlxtPqRhAhLIRatw/+tEM3/o/C8YnisnT+7rzlu2lgUm5ZDtt
U+fBD24hkkDbF/8kV5B4rr+kuYDfAEnfT6nzfjyZN0LKJ2yXDqPvhNsoYnBtMscI
K912+4AZQDmPlcaDUkoFm0tCeK3ym0pYqY5n+fEs6Jus6OIA0bxEuXljDvSWXbVI
nQRJzZrAXOFdqv5jpNiez1RDzQ8Ci6eYtoV8vwGpGqTZTYBxVXZV+VB8SniZs5TS
oWRbOGTnCyi96yswBZ0z5pKIS3FZH+YGnW65FqOfUHPsEcEVBsSzVoWALNgSBE2+
9gWVGTaRCKpcQ++AiniYY9K3gPa3xA22yZV4LDmkcgj2o9cdkuvUBmhjEWdMr4+x
3ibuSFgwT40I0HcbcjzmUVSvC6hvRh5gfxJOvUfFmq8LZq94SrYfWNtdl1AcFCQa
hzq+EUJD6iXLqT41yEXUkZz6TXgiQWoyPLY63Jr+Bws4ceTEaq6e7SruwMTsluLA
WewHtnOevUxuBxgUctpK9Kuhyn2jgDoAlTwpIp24nzLNes3hWUm6G7qYlzDdC4hq
y0y6C4EKKLCB8RR/p7xt65IsKHZ8D4OwNm/i1sjFwNpjbuyBdNgn6S62i0dqt97z
/4M5jihEcSfPCucTcwSbNr+UWl1FPLn+JkvW1b2E1aGsxvcYdtgJRA66MTTjRQjv
L/yTa0JXyCgWc98Iv2Vh5P27EHYnRncOPgN/hUsE+s/bG6zTjMpALmRpGx8H/bzX
q3wG0mRSNVLu2bcavZr0zU2uREpc8dA50n/L+u6x85iLZKJ+Zy2KqV40wB1ThCkw
vgNrzakqlmmSGHSqOqXle6+OdCod+PyhxnIEiixUk94j1YkOFAE3DisSocmceUUP
+n3dBKs4Saa7jhteWspyFF8+qp1JyyjfXpSkU8TkW63GrPJhn0l+V61d41VcLb9z
oJ2rUNdBEJ8cGJmoL21sadVMbuSX0GRNU4HoSpv+VA6AzbtCQbd/Izms6TBtatRK
92ea0eJyG9s6SExQXtuCujX2trf+ajuiLmq1lPW2KUhTGJtfblxUgFIqksbJ8qve
Tj7T+ZHKh0CJlN7N9v0tSJxL9S3fs/1rd6xOcB55AUgv+UGQPM6iPjznL5syTH17
be+TK9s9xuWgPuIHqUInBoR8laBgGSvaZVn3QFCi68od//wzhyLfL8/kewHTzCT3
Lg1bjd6z2sUY0nLQ5aLqlmgvnCEU7jyfsfasdROtzW2E4LSW9SgDHp1JQKbnye7d
wyb8AnNah+U4tY8mWIQFRtOwTVRWCaDpnqh9kY8OWg5N8Cgf9tyiIiyYvPS9vQEP
NEzSZykTgTloPROKZMEiEereFWGbkdvb3xlLp7McTh3VLgK+0+xfZbUS8XHDR19p
PgOdC6sSzJxMYqjhuzG+lJKKkqCuqtsgqUAhcrlN1bgGao4bhhGRItHVa0GFheWs
NVcov63rG8A/UxEstqI+mGGRdxD76kQ7RzOBBFXJgiuu4HYXQNNW9aZl6FwEjG8T
bcxFKutDXJwV1PrUWnEtdmyQvl6HDO81HxkZlHRSa1vMNOYkpajQUOjL/2BqWcUz
cUuPp6VSgXvzXDkIjBmy6YXeffFlwi/DHC91WBF6CxOyrTNxYm6eIXyDQxDPcD9J
vcZJBIm6Ig7Xlks9xbGd68Yi6w7EHXgU3mSeyosYM7E0DVJRgKzVnWQCSEJV7L1J
+lpvqdtad/RoiIeoxgK6jzOnPfHcjC6lTP6tkoUZ5xCqBkhrV9QeJ3KLtIzh1wpJ
UzlBbKliuyLqssXPbilPWnpyZp9Y/9aXYOV4sNCPlaAJkgboeIb/kOkEEBO1NnIJ
7FAZR6Jqa9k6RsdyLs4dsUKuFfa3p1HJHJPLtpZVGy72v4nhWNgpu5pg9OPy5Bwu
f6ieY38oopZvzx1fdGPm+xY1Yq0vxk85k2xcyNKJ93XKsDCtbiZ3xgOUYjdFU/k2
PqN10Xw0dF2duhm0oedHRe/UqU5FdPOfjPkx+dBk2lpgFwtb+9oJV0mYTBdELT66
CDOgcBFwpCmiJqon2qeOwFhupwMFTF4P0z6mtsoffXoj8ZuxyZnzubPSbXUEDVUf
MIHQtY/wYKFl53Uvcfg6mSVbhsCf9afgAcxnq4wKiI+Efs6zZ8yV35bEjPewaYCN
tvNYXr2mUm6w7fESF1eDFAZ+3Omw2wlcChkuMDOlXn39IWu54OHaemGEZkmN5JKj
mJJ9fL40/NHlAaTY004J1XoHp492U/A6DlInDXt1vHXCSv+Cq5H1p5HNT9og1jNS
rUYoB8PcCdkzU0EIMPFVCQ7IXkkUoClrdNpnUFaqQ7i9gMbKqtyAteqH3kRUegPh
/PAzcKF/EhdcTSOjL/Rh0re/HBdP3zpEEUhGrzDlAddHN1dEzGKJCZqNPfYeFhai
txx60GX5MIO/pNfjWBIzIJUTULlu8AhXk8GhEKCQWHDe+w+SWrhmcVQDZs9o7D8I
X3bkZKhYd9cBe6nxIwrb/GuQ+iZU9FqtvbNOiOo1ZND7vdFYRRZiS/VDxbB365/T
Ghuz/bsmfmd5ealnLyhMF2ralQp2HEKkKaJmyRmAthtn8IYb2v4Ekqqg2o7jrGdY
XWKiZQHTfPuQsMehJUxhfIg6LkNSaSGxXnDquKYfEJB1WrziFxa34BxroPfN4XHa
gIWqjXWKR+tPJ+Q3yFcq61iWgduQlDI5eZfDqxWe3tL0iOVmecscdHRYFpgWuhFt
jo1ZSwx6fLkXfs93QNIGQmCrMPHBp5brq4fCH8Ua8zLpN5QktRrB8eQR+wFCkSfB
B9Qssq00QA3BZ39TPVH0YhYkeJUA6mD7aMpGi2ovZEx8xC9b5bCkZCPkR2lwBSoV
rwjX4nCMjPSrMnI04B0iiDTwLOfIWatUL97SqxCTkBdaFZVfekUB6pqt6tzQdC67
4t+NlccCo8W2KWIDZa5WqhWUewkOmH4oWuX2UyXiR4W3EHxlBDRMbpykhU5exhrb
3dgSSPBFWMChhDkBHI53yEOAZ+mUQOB1sn6Ef4PHHNLV7avXocziC+9J5MjKRjzB
+IH4xJsZTU6Ng9YKUW8BA+5jw4EBDbIFT7mXGRYHLY6ITKZ76Ijl7aIt4DZsWgjU
asvScfjhNDXjDhSMY0L6T4bUyRKCOp24KK6ZvQcBKk0eR9aTldcsiuMp3VrDja3Q
bB7QKcy45rKhxxTPpJq31Cj+Mc7+86Up8FJmLnBP+rfuvCJTIBHw/KpjqA5/o8zY
L9uD1w6VBhQ7tqMtOwqzK21uNgKbU2J4whuuKGV1hqSuwE+4os8wMw1tKbyrS4rh
GCdExAUPuqob8pFY0MsDsskI2GsW2/P1T76VlKNGCsUMgNxkq7qMfwmJFUuVvIkF
JILBHJMFa5VAVsZWfky7G8KTYQXpwjwTxZ47xmgygIluPCj3JfyyHEyQgSg7QdUH
uIt0Y/VHin2chIenrooUpZj3jPkfgrlNoWQYa8B0QJhZEf+0U+fL7VWb42izYdj+
18qjG+EuP14n08ILZNnlssBzHOT4iMXZlah15vDMZnqXpOJsKddHGMj29pVi6aN0
0gtb48oSFqnj03taGv4utE4GJeX+3o9pOqKpblPN/jer7moDponI1QQTFozA9PEj
2y61sOVJcrCb1zAHGno54Gr1OFC9/zMwDj1bx0V1kllueatvCaVqLZBjEuVUnTRd
wfqN6IG174Ay0VP/DPJmT8PN2Bt2SdnsTSNSmdSa5Qspt2ktOX/V0xnZkaY6msbJ
oy4ruhghneOyAnoUMRF9Kp8vk+CF2mycgOWYZAdIObK0gB1v9iTUJ3qC12umDW1B
s4Vgytzj3Kca9wXrIY4eCoqCFkt8YZ5qwnlDDcSDKmBxXxKPYFWZnPIHlsnI+7HV
2VqgG4hCPTgKcCvU6sehsaF4FX2QFzkVIyleFd7Q8yAG4IFY4Fj4/vIe7Bn0p4pW
cxti9mWtcRgtEBCXL38YR3TfqjqtO8/4CbjUHrglNSKrvkNLxUzWeu2wzr6hyFLk
zWsjaAvsLes553FfVoRkSCwoQDhkzt/leNnV0NVZOd3mVQTO9v5pMEVegLOYZ/6i
K1Nx2cKOebj/jY2P50ihIZyCsHnj4DMXg0AzVFV/0IyoTYolQDFGvwjA5Hj8RZjY
5ucy5wvYiyh+lZtFbrSEGYarJuRVfeM5i0p+bq0a0TrlZSrSDK68zfTP7G+hFbox
WICPsJ/vYBeZugaZw+lTspSeT0mnxh4jyP++gAaw60+vGF9BsJBKZ3nPLs4mgsJL
GoBAYmwkDZeP65WX+rakzQQEpuZUnhhdxu0Q0VduUMnMdDfxzOnuMKFp8xrwLK1T
9ooTqSI96Sdxec+kaU9+2dYEAnaRL6eNi8wv39QdFBOMUum8TpN/Y7s4CtsLgSh2
xukesd+mGuu+sUPic1COaV7g/YSNYbMm651IgW650F7tVTbE+HrLEDTbgNjnvayP
g/BzX/Pn5rDcw1c3klaFfwFzFnhPc4v+UmKJ1up6W5B+rN7RycIAgLl6LGLKzWUo
JF/nX4ypUNIyioGc1fJ4cWAEtseXuX01BnO26VNle5kzm8l6BA1kompXaoO73tBq
0zmEKg9iAUhg3wpy+fM0aPblLFuSwyx0MuzLhl2QDb151pbnLyxYIdd/PEtQ0Qvk
HtNRkv8mQnxU1gbuJfFIuVOWQtE3lGAeRiyUeUpMX9X9k0hWqBCURCUSocfvZ16P
vKTIiLOmSdFpSK9h9XxcLQjcnw61RUR/4+WrIyyuu+mYwA2bSVte6OPS3eA7JWCM
F+5ShV20c8XbDKTdJTOxTDkYsELJuL4Co5KfRUUoQvLkDqpFTVzzZcffyvYuaM1W
f0V991RzKD17axduEPDoiDuG9E7WpXs9XeY8jlkAoPa9KdhiCiy6eGPHrLMnej37
aGEdEwY9fH3uHOGcKomsAmXHRUisExCzi1725VtmYWfVvMi5l3UrNK2NzZHz/ITe
iCobobaa0aQ/jCo8i+R1dy6W6ketkAMv9zN809Z17BzZH+yD/cOPDbIzsISWRtri
f5Ndd/9I43d8jZofd6TX6YH813eX0ZhM+a7tss0wCr5Lf/P15AeKOiIb/x7JTSTu
CXEwEys3ZHnQc4Z4MyRjmxY5lQvaNmikoDeHEENVuqbPjZ1gLxPziQ1G+4I2tZzR
29SnSBx/RCaG+2qrMaUhJtxHeU+lb+BuzQMTNetHZtApOs8k3QpkhYsIV3qUneVT
wJjW8pldlScMMZOA0FCZWXTyOaOCVAYr/m7BWdJTG0CWIh/A66PK4aQsXOVd4q74
kMgba/1zlKIyD/RzC5vN6fXM/pvtCvHr4LK3WbMrWxw1LooueKwFkaESI+69WLfV
FOBSCvZI7PghIT1gq7IOqbpKn3GwV2siCr0ZBy+tO0Zn5z5n6xzfSTD7vuAGw4z0
oi0tom033vw0J++TKs+i9Se37Q7PSHEnwUw/eFX1pHMfSyxo84Xn7aBR6pFa5Op9
25bZUkqlnkVFkuq47JbOSnM2Qg7/U98QUOBf+u9sqXp+SExhe4NLmIOg1hLEX0cr
+Utz6AnO08m9vhHVXiRmhGKK9XOZKdpoY1pN+CNtHMvrIt0r/S3jbC+Y5A7ljJW3
R+oC+zkgy9KwloWnzBbcCK/k5G+jaLTWBv5LK++JK0ejTypMsZmA+k+6ZNVBBwMZ
EyeawqHDXDprdoNPN2EhnkE+ntvcJ8wP4YqAf6Qg8je/BHqqd5Z9hoQR1xtcAMRk
cN5Dp5RASWJ1tROIdPJN37szB6SROQcCiatEpsJXswbhPnGfiiu1pIVcjDOOCPbj
/5edxzsdX81kYHonpsQ46n1lnJbt2gcRbH5zIR3GQ8Zsm9frtWWYvi3GtK3a4Dty
uN7snLENZn0A/XRN+zeOAuZW2OPstW8AQih6zWTbTIrqTPzpNrTMdHHI0VwAGTWK
sR8Ja77FTvOrgDuKfPHow2WP8NiucDtNBApk7GNHSApMR2bJDCz1c7MjZE6J4sQw
e9I7evRdBzgFeYX3vWrAJWSit1CHaJwtd03GN0aWJzJb0K/tSeH4Ni6Ux2+dCk9A
4sEQk6DI2quJ2JGjpqSPtyO8/Yed13MDWaJx4EcvxMfISujmUxOWLPEZ/Z+M/ufG
oY5VLJDsTNFSODQaJaiMSY8O+x9mA9zt8ECwVNNMntP6iZ6cMasuL6GJ4riqnr9D
y4PDW2iPom/Cv2CpvZve23vUI5D0xY4xdlr4H4Yw8Y3Jl5AwAF1/zVSFxvlhzT9Z
2+6lHs2Atd0kyFa/bzCcf90XYKyRNchFhHWBP9sUeZOt3rg7sktmF0NVD/AXtfLp
IcMPZckGm41ni1NQX5SJF5vr6Xx2nVoz5bimpdGWpjzzDZZaqBhZyX3CaLo/jJsL
0rAbx/BuufVK+tymKKVHjBmjgfAlt1O025TBqENsykHtgJhLabr3SJAu0cfu402c
pNiVhV68H2zedzXLvBBuSfmUn33t7N1Xpnbb4U80FIR7dIdZlP+lXJNrhlID1n6F
nEi8nDih4ZPt2Ep5Obk0qShOrs1kKh7mYJk3pfAG+btIQGCHgrebEZsGk8JHFlY0
GwCHiHNjAi11VX3buEmAEvfMr51vMvk+YpOCbZHn2RWWQnAb4X0nd1qlK6V/mbBs
kjUwwt72qV3dGhaLJz2aK2lqoN/ohxHh6/zaGVW96/w+ZxGJYZudOFE5/6JcFWWq
Y+TQrsA34nYp6Pcwo9+q3u3aZqYIV66hB1D7aN80s33vd2OceyZUSZxcE4p44c/P
5gLPYJeIkZ3I/VcJGuFwoq+Jo3vWEBPIN5X/rW1xgDYqhoqtfi0u+BbT83hkT5JU
kmn14wVnt9T1EfRj57QtUsTHiolB9736aSvfH3QAmQucOG0WKoVCmU3Dy5ZSDL52
P4D2gB8UsKn1VOYXtj7nwmLXJwZX94RLBHsMN/vUjtn6bBLpZGiXPk7Ru4Y3otDq
hZFNHOtKFfXlVWe+g1jBGwvWNNyvWBwPsfvtrvlc0+csfretedZ/nGpIgTW+8f33
SHn74x0Uacqw9YI1/N6+Kf2l9cR37z7DPsOTtLnFgtcsDgfBRZKhzqfvemFYe17a
kixKNUToPnyi9ow2wAScLWct1RVT1V9nR4CsiOiuoz6S4me9WSHOcw2WDzKnEDD+
MDjhI6J+rx96X73hJj45tkW6DLuXxhkXYhHuFXpic3hBiOrQGoG1+bxanDDlkYy6
AopunGGweiDAgB53y9YvSapfdVY9jc6vV51oRiqf94nNembj8k0ICPTrA5cpNQdC
czO3I6XerQnFwDYakyFyFaidhGJgzISOvuPFj4RPP/PH7Zbb8aufCWO+HWCCZqGb
JuehmZ3QFXcSOkiYzyX+UksvBBXVKvZFa0eFkQ6fWXia1xYpS/NDiW3qGnKhU9r5
RGwcFhy0PUR29yCmoPdY5nlv4wMtT0EpUG0Cwl0f+YDUPG874obLnHA7sJkF/HWM
eh2t9VX18sIfYR2dVrycSqO0XUCs5jk3sImHL1S0TU1VMqO4zdtPbNQggFXx814N
R+vz//RapfBKOnGnDE/ZO7KXnQGI0VvdcCw9jN/IFTPZDmq6YV0+r+Q5SoYKRBdc
9FuxfSSjkP7RQaFPLGeflZRd9wd7KSe4R2/PCJPx9c6Yt66oovJc+QFdRgDPFxrq
3snXEgG6uzcTWYxT+Dul7E+Ul8ZNVZItsVsgSyJP3Mmr8c4LiQ6vF2A2CpUEBYIV
8uL1Z0I/1CB8ErcUMO3yrpkW0Aj9NOOgU9gdCYh4L6al98+45ob66yfxikSiq/Ys
mFuBDc+xxjvAEi4tGk/b2t9V0rYodcy1oBithPS2dUWVMluFEdoyDO7lfoidCUgv
3MgdGP5pMYGbF7ZnxAROHxIh+McHA4w/gXGv1m8kVcl1mWAhCwaIuTEcwE1J+J5F
Pg8kRihTBbrznkdtfXWJ1Sbjotg9VDILNcIeZWGVoX136GIjAUyWa7rp22xQupC0
0UiSivrN2m6r2LEHDNqSk7AzeaqVHo5EFCsTiG+E9xa9I/28l/R3cUYk551vvdi6
W2caJdUWPcuszb2/7fCPEQ7fwkxLUouo31hW+g0/mPSRf/AhbGjFCy02ZnU+wXGo
JXGCoWlQKAetfKlHkRpVlkj8nM/R8JiifUNa9yE/6YaLpULYNB+c2Y7LRmmP0y8/
JVa90jKX7FSiqHh5Vn+xpFQztHWaIxvpbjP3ZOlM+YOjiPO1Dph0FvsLj7+gAzQi
6jn1TzXAvg42hwKS1BIUNvEJzLDhtAAbtouVDk1BfPfatUjuvH+QnnFPjnjKPcl7
KZJVneqj/1YSZ3Rm6G6B+nSzNWRbJM9Wx2QXONMlCYK8S9a8YBE1hXMRyiUgBoPN
4YY3NDNG52P2sMdFGXKMK18aS1my9imAwweeWtWuaf0Xn0p8DriKyI7BLZnpKTgB
sHya1rII7c/ebdXHlIyzwfkVh1Z4/M9Ga0eravh9OYsX2NiU9fVqUGA7i2LZkcan
kCP9VVzbqU6YO5y2j0thPOy6gYVV8031E1V6T5VkDxL8Yw4gMiLSR592mV1pl5Zz
zoqq1+Ak+pscutDaGASIwDMU37TLvdCOJsP83fnxDONs9hAaUiwBRvPRH9BLOCpO
+9FHv44DM+EJpECt57zZIrt31b8ucM+hDwg9NPAvh+VL/P0nkemArkqEEMYTGSTO
fiESZ8ShhbZyfbr9pgvwYnvldqX5gGwv9NCpCiPDx7RtwSWOm1+YenLCweBRMm6N
UrAjY1VOLX0ZsWBnUZQkCfBF6OwR07R/yyhEVZcC4dYrOZo0VzvM9rsxU89b0Td3
3so1/1q4b8411VXTNz+XuA/N+WoXNu49k8PU/0rvfsQaTpeZCC5mjSHG1MZXRiK3
MzP+5lhCFGcohsNjMTpXddflwzxVZfIEPsDFVWou1buDnX2Ht8+2++szS5OIeLbi
3dl1S3E1kbSzczzIYcvVm8RYNUOe8ZyvM8VXaLVLOS8Jy/OY6GEA8N+dMNyWsVVi
EXmHZ2PJFik5uULJiCiNKDKzAkz4Tc3KAr/U4bZftZUUIA27g86t9Ay42qylzPwB
H4t0b5OxTmkyKk1xmiE4ynOKDeahrWnY70DDsSLZ46xNEr9/Wa2JCiDN6u/8nL2b
CkbRdenYUUbIicKlCHfZGZhqFzA+iPzizj7KZ9nzjTFWon+8lqm4N/Oq9iSaPHBd
AwdVc34PsurChVh6LZqWQ9QO1LcOiQFPSIxIXDzPcpxW5E1pdFISTMDaeOCJMopG
LQfbx58Iec2NQfWtiKa9pJm+lAcuqNJhKj/Lsri+NF9mw9YNTZrnFA3ehcDd3TRC
yCPJBO1KRnvcshA67M1zCDtcv8OLccSbeTns75lYzS3RztCDbZSO7nczqST1p1vr
2L5IgN2Q0MWHpAqmwuMG1gzAytWc9357/JtKk5DRuvXmKQu7tUVH0LSy3PQoJVy+
kG44+rZVKWeX/C2Nwzus9IEMNISlfWufV50OWEIzZwBRbr5+Om57bJfoVhA6/HiK
sFVvtP2Txi9TVamsjY10VJ4hE76hfB2UvKz0edTzbX9wF9Wo6H2Q7C4jdAiX9K5M
uhC2Iyo6ypRThI7xXgMzsER1lYzJxB8/r5zNIue/uldvaWElyi49YmyIgpfMktIS
SM69gbQBshpnRxhyYtRuvccTQRjAygdy6/KodtH5LdDpxYW0l/XHp670CoTomCH7
GBQ7pP4U4U+GPcWsTIc6yF4iWWJ1bdd5iCJGiKOWTZb6FKKAlyLxGwgqM8PdQyTA
3lzIkwd2ZtInfEzEd0WM2/gxA5KPclKkUyIH1sXq17NAcHVuuD3IOVLBT4WfY+Ay
cwj/Tr+ardC0g+LnaNiOolnaLdS6JTZl17b9hoYpVom6FDaDfNwa28V227mByd6B
Q3+h3VE35JtoMHMl1SrqOPufLg1+/DkDuFq8Mk3HuTYIDS9+C087kkC6jrnO8yvq
N04hNOqNH9xfwRaxaWSRj3U6yeZneQzocsnBmbEWGoTr9JSOVEjvgI4HK8FPZ06v
Q2SqJXMnnJXJaNieBn1FD5Gp1qBKwN9qLIS4ok+0TubD6M9i6ehHiNdPsHMPagtG
cfdCkyHEaI7aBjnY9wjfbIv7g/395bWKbr5LbDGTNc6hadFOz+6If6jkdpKAp6HO
Tma2pkMQotzbFmAqr6/1pLkGq22qx/9djcXwUfM6VtFEFCOV3GS+J/qmZ3kyTsMJ
ZrjhnJa8E+URRdAqRW5tqAxnonqOCqrkoyVhw64iYGg0MWNCZI2ECuLp32Pwes4q
wYy3d0aio0lCiD3VgNSnl/fANvBU1yzA+aDEGjtwCPTUXVTgpW1g9pyJKF6QxiJb
Ki3KbdvZcjsL/szCVmiHlGBxigM3E6LPrk/uq3OD57GNE0cPR/Rh+uL3QqXbKSOm
tdU46YWFNFrUY1NLDAm8NzH4pKpYNimW+nYdHuw6xwi0ka5R+Dmtx/sJVaRVzE0J
Eot+3rCFc7PvlxRUvy43wermFtLsJnxE40czSDA9YPMc82BpRGdevXBNEEAxrbty
iAHL9bRKT3j2t/d19GJnWXiIPzmgUzLg3jq1joZzToc0+tUEillgWeiKbdLHbsre
IebuPgcXaF9TPEjGGjgpS4oS9sU5FxO6Pnx3YPmWPDutVJ59nafc7SxtvgobRmhi
YZL7dzzRxfukKkzYdZZfCHSg2ogyngMZyXRSKv7rEVaPE7SGoJ1pJdqVS/w1j+18
GO00zPf8MugN0jwRz9IBHylfivh2sSZv5MqkLVwjQYR/T2gi6Lnkv7ko5Ja7VmTB
b7B2IM7zUPxczLlFQT81YJPsXqueuF4eZwQL5cLPIyJJpXGjZYX9vyaGTPvBnEu8
eiBMJgFIewe2qAkK40LfNYlcf0LTtKLB67QZ5aXzzmhzIcP4ihL4FQWzmQS2poWk
ZbMiInnrit+2iBFM6sj+RC0/b3kRB6ji+7ldd0szFVgyHf+r1BGMNj5M8UKGE7mr
9BrFANjRn0fEQBKxkwwAH+chUD5ErRoYNRMjeZOyQfxoOfv7h5P1X/Q4vNS/LAMZ
AdVOab/ENKZ6eCqKZymCwyIr289l/aL7NkNLmhh2d2fFtFpO0WZ4bdN643ctu0aB
PvV+JT+/DOPk/PJc3M560KWyXgZyhJwf/tNDfIqtL4nejQ9Jd0iKAcaAPFOUrqYX
x8TGJo/w6PktMXgBcvY17c5fempqKeCs3yu6SmzamU/kFSEz65twpPHvQAgo73dQ
lTc2yMLGIy3ygTrYxd6Vo+kJVFiRjzGieYRV9wQjANwk84UTK5YdUoH3Du0EyseY
gXvAl9H7kWBLRuhvQbb5LgGXnYVT3TliZ5lz1bJGP60hXWfzxFqNtMwk1nkWplIj
7FEdcWedrFhLg8OLUfbL85N+ujeBEQ11uic/vhgrJJvfcSlBRmOkZ5elrU/Pqfuk
t3LLfr2Ol3KFfhIvgvIsYJ/mEahVrgkVYg5c1zY03vOmeQaLZTUi02FcCe+1QfvZ
HuYK/WzkGNKztxuBtYocy2OA5ihLD142UqL8ag/V9vjU5HY3ZhCwEuoFmgleqrnZ
5TI2dVAF5opqKSm2rL/zU8fX80xBFJ4fyrpd2kxwzsprnBpJGfoDD2TTC6Ib1/zQ
+06ZjvwhfmBBT/el17jOd2LPjOVgDD6YO0WNoaivWhiDVmcqa8SneQ9YuFOg3LlA
YEAoUKA5VoM/B4TIO32hzDjDG6rkls0aE8rKhX9RRfhxaGg0aS68LE3xVPbkDRPp
uh7DsFGyOQKg0X8MjMWzz5/QKzSmMYGdLyDiNchgW4EHVm174HnOHUy1UOtk8icE
oVY4uqoakM9ZHj2yJ06AkmO02UsYv6hHbX4jjLr8TepBMEGnCh/qK3LIdmk0nud5
0yEZ/dUjV16hqMd8zlEeZW2r/5Myq/vOnp44213vGMhLWAGYzkvZRUoBszmh3whH
KTdozH39K6jfPjBHdW4Y0bgu1d5NfH0AGKGePRHOEW9o6f4ie4uJddllbmxb9H26
RRhg1lHna4kZXwTyf2ptt7flOjxEDG7qzM1pzgGeNShoBaS2MWbNADVc0244j253
YU6gWsEqxPJ2Qo8VeNsHx8dwdJjHvY8C0vZlm4s0qW2ir0F4sn4ynlmBDN+jBfFY
MyezFGU0q/GVXT4dtuscxFNiCUKBM9CUpcdMpDOHhj0ZI7EOFI1VvawIaHEtzFVI
3h3LKFC8Mk7uG1Ae9aNKoO1DipT5JsBpppVAMiH0SOruocVb0sEZMHqsC5Ng+ZT8
/g861u63PDS9dGcmcf+Z3UdsYFUywr8LVdMh+7ZCxk7vfs6Bhun1LgB0+KRCXziq
6j3ZRbvKR1SRyVSEH8yhAu9eXviDZ5Qk4nQWf/C+WiEiatyPw8THDDeLNT7A0MJ3
h5xhyjT08kkYMF+ROKw6LpdCSk96UR5xGQn3z6fn0pm+nRtVcobeYIZPnZfMvwFg
hEcMd/JvbRqkxNnrVnFPws1llMmDpaQGSxCY+g68igQNQ1GUGS31SFgxsvIrdNaL
51J/EN+fFeM8r0qA2KzU34GnlAin1Wfb1rBnDRYkEZUoKyGln1hVw5F7Gif0jKVU
o0c/TcaDRr6H7/+5q4brrPF5B0fYZVXXOdxhNVU9/XMlCKv3omrRANDMooLhN9s8
20ygIBr6MAa4FgfGfduxf1qAZKhmu3JCSPlX6bxYwL6LJj4dM5UdQPwoZ33gyHEQ
FsWjq8ej8JMUZVYzuA29J8j6A0Bdpkibsle18osDctMf/h1DKEKWtA2Hm98t5NsD
GkqX26Z3hH6w+xir7rfpv8CMjp7laAHyzEYcd5FSsNKQrinpQOLZZ5Efg7SIAn/U
7MSoCy63ZGkppbIUyAtQ22lXQa3dteDg8rOxmt6Tb3uoL6W60HGJDQSh4+gOgCdp
Es+VRiifNDAZkS1kMWIVjhsxz1fdHDHDSVtByWVq7FLvR6Bk1VsoVuzCJtCjoxyK
vQ3FGDQDs+D07NCKNGsrkgjfUUECucIIEYhWt9vdiJzgNu+5rf5N8tqMRhMnr4j6
6XANj6RVAeRIoibl0prE+3m0vV9X1hJpN5gD/s4PH2P7VFkBBsJfIwq/CpN0El6V
PRaipGA2tiaj1byXv9ltm8B8ylMmfnn+HzxJEoxoEA+5BDhfljBSU5CDVlzkO1UU
aJ4klhe+CebIExdLhLguVdqcqJtyzrFyv3kpmDkJHRvhrGh42Cymxyv15hgZ+tvS
c9PjdhAy2mRrzGjzsdKVklhukstlBHpSQFFGs7OrilujP5sMG860BtoHfbEEtJ6F
p+df14z4sja6Hvfd+JlGZLJuVUYzd4YO448Y+M/R1m2uXvp3sjnYjRUtBVR4JDzO
92bthJ3YLeODKplWmiHfW0t61NzJmkxAlrJAMIaLOXlWyFyO69HGXuFyjUHqSsIM
29C07TvoGGWhEx1W0ioszfF8gG0pz8+S5itzlnjm9bwu3ChBht+F7iuhLv4uTuyr
o0M3EmBVIwyBKlh5mV2yg2/qcEljc92wkX+eXHowzcjHDwPSlZLHoZoL5BjlvGF7
GwCVuX7pc/x8dlPsb3Z3XbzfOAUOeADzu7TzkKQVfMD8czhqPZWH6yXUps80jVjD
eHDbs9dyY2gTtuaIRzaDYuYNpjxlA+5FtS8lDAF++e4mcg+AfuZkKZKASZNLK0af
6wTfIpDlik7IWGpdLN3AlNOA8JpGWHoxLESdfIGUSuPko0mQga2Ywc3LoLky3py0
RjDenXpMqx1K9zmJ/o+H1y8QW+xQdvzZL9dJoi5zGHrgUkaMI3dee6okoUjvnqeo
QSBXM1YgETgQjmKD+2dUXibXSstnrWUnyJpr9NrLWJg+w2N+o+vzdC9FWW3rhTJn
BR9nFJ0XgHS3aYRDxYCd5h8CPunpFN/10sT/o727PDI2t0NFuaRHFSnh82oTtVJU
FsSXVk/BU6Ol94i4hncKKsaniLrPtzrqX5kZ+CBE0VIidZAliVGy6+PP4xv/czEp
PQzGsjZDYBrt7kA+ML/k+nyzaI2M+AhYaeuWOknwR+PMIbGZPXZmjWV2DlshLdQ6
yDDUWiqJfrmVJAGzzrpr0bS5rffN9gAWNsgPJwBzpFYrzSuNrw4lEEfvupwFH3+d
hLVZHJhB7r1JEbYdoBedFziz1jv62/qm6VrwZJ8ko9uDq9Ej5WRZpEbHtyypOOBI
1muo8hs0hcNres2xSqeJsOHlUbGzDFveTXxTvTMouXGxcNimhDQDogAgOadVoQkd
ZSmPGAsFDHHOmujMIYbrAjcIwlM4gDGyF8TuCN2W+VA3WOw3ZhyEzSlgAzwULXnl
WDbPDoDyWwoAmVSxg0xsIb3265koSDM42SOj2lSTHrZlLkNYq0jF8h2m1q+k38Zt
6S+/oMFX7g1U+mFwkUguNjdlBDwGWC8pCGm2LiBkD5yL5ZD0OP46RFjk5W/QLO00
/78fw6NKCS1ijpBuaCSaGbkobgmH7H4mVczHAb1kVl5/5busK8EdscmhuCVEuVTc
nds9wgjlDES3dalNdbEUjLA8fwmtNaA4HrzRk2OGs6KDVNswFwVVw3Lq7YIwOOwC
8CMCb2DVHG6DkmgENhGTLAg2t8uDMDYcmR1MaFDpWy+tOW1mMR5K7onFjEGhqjm2
96ZuihEzLDiRZZmoxvDTMEtpGPJTCosrAbRpKfPCHFD2MGiS6YZ+tX4ZTFO9uw3V
cS16X+ZQAvratZNYv5GKxGO7tcR+N37ariVIr2fl1Pgdx6VpOBL6DrTfDfStcgnS
z5fL1p8E5hb/CgPfj19u8ZgWp1lQwalFKRGusWR1flb673xxXXeLcmhMv3CI42V3
PoFWw2nzyuYbreKn/zC9gPXj5IedOeLFYQc1a6IQCJoYQNwJcx9pjNKniRiHGJ32
Vu5sXV53oc918BX6J8W1dB7ap2FcHZcvpytyzGbdFSMbJL3w3JAEVcNAu2BD11Ez
emtqCI9RQFEjXz3k8G9o/17xck+Hf6pscgO3KGCckmKQNkQyPId6i5ZdHPRe49E+
vMrPpRdEdk89jF5s+wWb4F7n18Fosu1DbaDcGnuaKLxFYPbNR6Xi87sM/WyHEgFI
sv2gLnfSqHcB/Ay6RHNCF7I+MGUz/yjhmGECfDxREnOEY+yknP16D0m92ax48yTN
AukWGPG/U43c84LOYhFLj3bv7ofZIZqwfMZw5UuJQxaZGxeRg+KJYnTVBAbeUyLd
ANjp7wak4PcG6MmRYUs/4XJhXleXdBhIGcHmDKHHOekJ6zHaegqNx9J1M46MqXkD
udvG7nDBXCrKRhWHUUBc1m6B/EiSHUW7I7n8sYDIJW8JChh4YGUoHnBl/JHlc9+B
1prw8Im+mnA7CTFDf895xWInWRCY51zaCxBPHQwa48Qb/657ZKS70S2G0+cPDnk5
zRzOPSlK6YU7YGVmmflnO2C+Is9dgS2RCLZqcTkRdMNF8eCy+I6dCkP3ZuBRDb/3
QS0KM8BWZacrlX4/KoSp9h4+7+sgjq8hHsbLmU/CQIz+cA1mP5hftFDPud083GvP
+7V9ybMHwZ4ER6PvJSBTtA4g4c38hvJF2JFPi++R99sEU5XqNE4JY2LNxZJ70425
I6AkuZMsh5nJa9UwaGLS9N3DvXo0RjdRm+n0tAGc8Dt5pJQSH5Iwg30vxs6RQau0
MnVnLNbdrPKI6bJeWQ7HQkeF+J3q9yXzYrC2xfP1R+uwe7lTkv3vJySJ2WdM4d3X
4MUJ5G6DIGIvv06tOR8Cx3ZTCAQJVxeiwI/45pzYtqJxHZ1T/LKOyDeP6jEA33w6
idZ0rqw9+LvLgF7DmQqA1dCqepUkWaLfA621nx/7vtQpvRjk0KdThpwL7DgVvBxo
JmhxBYsteMzmEGaa+LQju+YWC4pJBnqjLCj2fHFKX/rQPsj4pM26jmvoGBbXG+HU
Lb+2q2/ncqYz3W/YTDHA787i3Db3gf611Iu4A96rVexDhrlHNhpcYMzPNLT53eoU
dMa0AIjsXJ7SW/8yDpdA/CPRuivwxDYY/1jJ0/Kzd84vzY6k3IW6d6CvY/NlriPv
GQGMxqb+c9Kfe4Pwz1exa6WYefDu0FOidHOGMUiMHMC9Aet+HRGpXfngvLH+T6EJ
IBsPL8mGyinYfEMBfFuUIRD1uDWFrBMO6FkQdK32DmSqGlMcFrscaQAUbGIoIGy9
V2DEz+OmYFwpssjbyhTsGGcTU/c5cRfqCdk7ZgbUT4Tw3u1efLhqVmkGrzNxx7Tv
Y1UDQonyGjsNf1zdeXmLScwzvj2iZTNZO+FMTQZqhZJv0OPegftO0t+cPz9TR4i/
7RkA7udhUufYI7nrV44tINcGqTT9PPNLY3mj7G4I1mTPq0XbxQAUrbkjPb3/6o3H
xG8KC11wSuEH0Bl4MbK0nqa+ym98b5eYvJMQm3WqUgoyw+xJrI5mfuS0IFmrd7B8
EIQxlqxQURRPt6sgzH+1ppzNyausZm5GdwZmrL9QtlJ907KGltC5I8tXQ/Ie8B95
RFIU2ZuLQCxB/XPYLue8iaKPX3Gng9uzkVrZyqkOFlwJIZuWpN/jtzyIK8dKvpO2
hQnzSiIqHF58JQ/9uT9dqLhfqlJI3OWIa2F9R9ijzytuo8bVh0ZQI2egMdPO/fKF
t5aE3cY5MbBk9fMEFLktnWWHaIV8rnsjF8Se2gfo7KwKUCHbkO/WNm4Cg1hqBnYS
Xiupo0sKEWf2vpBOFG6ZdPfPatbR4JNOUB454+QNR8beMjWruDSTYvEk2DHlujyH
CvslSt/XHGhcVTbUPvxdipfbicDkTdkOjvhkhL/p9M8Mww+e2z88lRQtdrnS525X
9OIB1WEYVmZsWhM8JfLv/CNE3sW4/D0VsIhcL7BtLfwBD4y4I3yR4AJKVENKH7KX
TABaGpxrQittTZKZSw1juySpGoJD7GBVbwZ6QtxwnzGQcAEHAOwKWLcPUxtccEWd
eH4ZP3i6LBz/9p8/TUShr7/0M6Q/h3fsKoAuZqeH753qaAgLcyQKfIV36PaCXp1Y
2cHlphFJD25HExvR0JCCcYBV7RqfK4+BdKx0TOQ48uhegGWlzDp0P24u9yibUqWV
C+VyI2vg89jvS6bvV4EF2QzCYa2Q99brfwRD3Shixd3Wafrc0XEkcVI6D/Bv2AV+
v4fzvCorDzkoERVCdA3eWpuLbAyaONrzrfaXVgkT9IseLDNfW8Iv5o3R55JRiGQf
DaEjaDvPEsBee2z7MHIgWNYiGFQd0b4j2vuQojPUrpuNWHcdjnW+I4MhaCysAzjs
ggmszmqhRiL5sodTSAAGvQLBq849ie7F8XV85NqMZ/1JA4rLdNc4J0tWyD19sDDG
XOB8CsesO4Csqb/R1WmiujO94v6vgvpAIGY9m/3skKOVAVIthUB0hpeG6VYaUXwR
YY10h5J6DWI6XpD6+ZYlhkVBHMiopD/MgCRt9vmyI1UTQEgYYRVcaVzJ0YhRkYKU
/icbKrQANkDjpc9gRnWD8SGgoPtMJwyBAravs8xjN+3aTMhi3oRt5azQqysTV64J
tgCDwKVT4xglT8lYWpcNkVll0EQa2dIZR8uAkbL30vLIjZZHzAqv1Owrafb6+/yf
FfHjUnMFAude/oY8sTz08yZg2CuHQzsWj+veimHqxRBlK2S3np1j2P7pfFHII+p0
pGV9P1OhKeMNtMePLOVJj6XnIbG30XeB+inad49iCIBgBfpZUTt3AaRf4mUn7MGI
AMTmAFt+E27MJXPCmN+HLmdlHQEa0qGP8EN/3s0/5Sqftt18rlYbG2PKn/Vg+/X/
jggdn6eXVcg6dLTCELcwLOxAJP0RfC0BHmYvk6OBw7NOMXAyeelcfmoFMeyT2HvF
gSe6+ueeJjUyUyZgc/tadr0YPwx9Us/1wzslkk5WSF0YWOzZh3XluK8EHGneN6MJ
O9Y4xc9rJWicAr9hQdYjSfTZgKTGzRUNRwb2VjBsbXin+Vxw5AJqQcVBV2Oad/yO
Mu/VdgxLq0DKr/+SNEfmxxjntfnfexBCtqhlWOwuS5metHb8qPgwVDlV7IECmRW/
IvSKLSAlFAJuisKI7RHGaQNssB2c4V3x1d45ZfCk6AoErxwsQ0QmoBRmE6AO3PRR
VVUpBc2ItKqVAdAd7cLXFOXwRWr6O60A83Y6dJLRspzszCEVekN4nHgrrbPamZ8d
EikOkpGkF9x7bhFfeJCTPSA16MRbZPN8q/htMK25O0910r64KDeZ2EY8AwaksTQH
PSf5UQmS33WeBP/QOQDLW8cF8PXWnnz6nESM5pFeVNM=
`protect END_PROTECTED
