`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iYtABsR+ccnhmU3zdtxmSCwmsXk4tu3saYWvQIid5FsmhC0tJxtif1pQGkVTaTTc
KV/V2AtXoEg9kdX79OHC0z7NJCqusUergsckQ+ujjiXfNfKVSOSh4BuFo3EovwnL
WRP9qJKDR0ZlCsACh2LBmpAf5Lq6itM+6aqNWYs3yqB8XOL/UT+2YzuWNsAPW+Xn
MfBo66AOfoSkLnJTW82LUy/swx8GKB9aoWr1QudY+mgF8ImgTolueugrk9pkATEy
sOwA2J48NgONW5HkwFia/SROx6af/hpalIlKDXkr/MWEuyZAqDddxHoYMuxC69/I
tpGKFmABegUMiTVHY5s/0001kysJTQsyBIhKiVQG30FZkUfgGmeNhEpMQJTlq/Ue
W0GbPLnxywDiZnmxTE243jQHqj4P+fkbOeg5DqUYDG/AbXyjCjsrCK6HKcLbqumi
A+xsj9k8r2gfM7lCboZ2ra3S54xOzR0vCmWPLNZjXYM2eXWHUOY9U9eBQw7VXskC
NlLV6GpGRbWbjlBDW47djIO6u1xQ0ObDG+/ebsgfifGImUpLP0L4Nux+KLo9Q5uA
VLIcfUIzb7RT34qxdD2hkURvGwB+kjd01+rJF7SbLJF1STxETEiQ4nN4IJzOc1kQ
tdHqDlOhaLdGsYj5M/+nr9D7Q+M34xQ6sZu+QsRnImRIjguF7jMqU44SK2vzy3Ih
nxHTZUEXWiKybsh+zP+aRMx/StNEXVFfKhv2r5l6QeBTDV+EDegv0NvoZPl1RrKZ
q/Gwf9FvNow0hPIELHhxdAMKELUBgSgEz2Jf93UB3PFeLMEFEVd2TUHp8cyG4EJ9
xlzQ6GNtz9nVajPQ2cRxkqtkNvv9CnSzDWSjJg7E3F8rkdLWOZ9JQEe0HIIqcsp2
`protect END_PROTECTED
