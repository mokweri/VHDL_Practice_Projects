`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8gEsHro6JpyQVhI3ZDGCtw8fO262FYR4TDRpbR9G84Xksz0lcy1uAVxcJ+lZSMA
GOvaz6ngIUBZVoEA2DNobMxO8W1pUK97uqbSiccxMPwBkOCaKABF1GIWIKJI5FYs
vlfqSibVR3pdb/5PjFqL8rC8lid/6BvmjPwiEdKyLo8rw//AIQn8NFZ2eNETVa7k
bTtIt7aMA8pGWJFciLqaG9IFGSUxL0f8BrprviefQ8KDeSBFGjavm/ZNXn5EX/U1
blYr0LE49uHrSnvdZOd9cP33W/1civ04yJrY5HNnqNyYLIpOK0OaUHmmnGZi/HmC
suG8pSLaqQ6yAqcLrDoko1os6h6Fmhqag/ZR/HrUXOiBPwPEV4nmjjIHbbLhibnc
ZWY8+xXw1rg4D9mlJB6vYPbdomAOEsOzBvrOb4SW50s1eA7PsHSHmEZtMLnS/g7x
Obrltope1/Svb7Hw47iM6w2aKsXVYdgSf58sEOGTCqOwViT9gviOopdUk4J5sY6C
SqlwVGg7OtgLT2Icc0Mw7du/4I7SqoHPqz0Q31tSG0Is01LjJnIfKIo6UX0qFqh6
gLHqYdbAh3gmVOfsj73A+LYFeg6zJrnoxiEE9qELrjeJEcWk7wAwEmcElBxH1Sdz
s0HegmcY4N0vGyjsBdfY48J95BN/HYZBa6DkecJai0SBmpTI1/4xHt+aZAhAlIwu
NtY9bIzgp0vpDI1eU9l7ekOYUaZsXlfgFzgh2HnX3BudWHRh3E/cv43D3P1VcFPG
SIgv2GCRRONnWhKvIeNjUKtr51rIcvl+UskCzhQVjwb+v48INJwmHLbdHsUMQlvl
He/bbY0EBabcDhit85UX3/Govv1qp7w0xMdaQrn8svx4InJiOSY3kgC9udQlJ4s7
1pVUc2YNilxRMSMAt5E+YR5KgkA57qAHcIYsxJNEeyloVCEH3YV91adJacQHfT64
E3FCRMIG1APtPeTN1WbopIrlOtjkO2D35RVJ4S3VmVem+K86GNO6MiUMHElF2dFB
5MDnoyehcV2bEFBYmi53tiRIPbOFbK00keatrE3NbKJ/gYdqieUMlnt7IaY9TM3w
ALAX3aGvp84naJmujmgNBcUgnm21G1o+MzX5Pe3pOs1kh1eoSsizpW6X48yr+Quq
bsPcqjXfS37+LNBLKQQ2+HWFJyoDnAaJqxA2qbxfW1wbGvzyHFH7tQP212hT7jDQ
uTZ8CFirGmkWHhWxcNEw4HiS0N7x3nekXZxvAOjI44G+BvDId5k5O1wzBMcomNp0
UoQNOOkbnJi8XyFLjo8nFicZn9rK1gf63prXFskHfjPQ2q4X71UwhCRXJN9ayGCD
6SX2txMr2CjgdvVzk24ysdJOEUv5XB/q6rifIYTQBdOVvbFqO2w9tPPbQ0kpci7G
yfqyDtf/y9Fx0Qes+jFj3TVLlTpb91TCUF6PtT81DtgjZ4qXQNnaDJnikFETemf0
fjXpfon3PGiXk34KIJM058RWzqqg9CpwImKpmty9a6yb9ZyVHuJ+T8ZXJ519NxoH
hOixvOyOj0CzxMTdRFad68qtbu87R9uJofUi6g9BtClxujM8rS7xdLW0ttNa3wKn
VjkRlklvisr56o3MUDroCMYcBl2VtGfDzSuTDoWqjXHaHQnLQiwxMP/e8yaKmTnk
9cHt90snZKW47M7rI5ndgDXx83IJVK1S48citrd/d/Axjp5kMQwxg3Oc0OhRg6oD
kw3Lp968aU37gAhoRbu40vjE0r9nk6CYL5urR0gihVYz2TS+hsdy4XElrkL/6Y7q
wGxb0ciipqULXZ133lbym+74kjs/lmLLgMXvXkvrslOLMV6HTOmlEFm8xEFP+WUS
UqMqpB8q9eaeuge+9a7WrtSAjhNC1n8LMCqysKIyp6QCQhqxaJo+Djk4MNkjMfAa
XaIkvgWJ3i+QJe44b5XInHSzLB7C+RUWkLeDiOBV8AZF2iy3p1alw+w3v/+XW+Ny
PwAKFiLYYP55HGZR729APMAry41W0ry2LlY070LKR6XHCGLP+w+7f81QJ/OEwlZp
iYZJ3eEnML+dGqabBZZ6nxvlAQ05N7i91RdaYxxGpJn0QeYRp0dlk0DamF200Omy
r/B9wUbZEU00dbj53irJNfiZyF0JWf1ESeteM7cb2+qRDh5XIQdslBfxRRpA+MG/
VCi+QxTqd1BdPh/+9k460/xjTSda7wjcc88/KWKPb1dZIaJwNiw/aHBs0eU31abE
bOn9kPKrx9Pn739L9iFUBuBFc+9PnRCacFUo2zU3ib+vH8X7pxyY45+Z1UxPNJpz
QJlZGGYilkat00M5xr5I8m/7k2iNHBfa/vHdr86mVb+Ka/ROEGUfWe2LkVp4seqn
qbbiNKBTvq6LcTtdOHT5vvj5vLq6Wr/6AJcrANdbiITw0ywWpUGPxYkw5EV8j1c1
`protect END_PROTECTED
