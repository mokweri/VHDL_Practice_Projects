`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcpJT8ex5mmTSS852KF4uUoo3b3CTxnA+mvd7cOzoU2ZLySowTgtAJ0DkjeLwE2+
jxPHs57zyq/KBMPp3FHOXvHp95nO42cyPP4rRJFibaJewuEKN9DyqEZShMyHMnLH
IBy5LytLpoGtpK1g19kROsLdself+W8Fe/WyX3V5+8fYbignfijOp0EnFk37RGl8
DSYXTuQ6s0jA8rDGcMcMRUq9lXgl3UeFvsbcICI2dGnc/vrgHJoUcRanZknG0tF9
V71JEfFP+c8Xn+Xzyw0pwdycAeL7U3Plk8uPlhlZRyYaVMKyXVvZ4r+a0CzaK2aW
gnPfa/tNt7k3sj7nN9czJ97X8mIS/8Auh02mHM6dJww3r+j5GkMxPlZWZqxNKNDp
K/NFuWBibZCcRoSoXF8HCaCeMnjG3JvlLFHRwBknx/T7DdqkB2UMf6fuf/lUiEfA
NfD1W/gXZ13XYkXAwOV/VHstQSMqCm1q0EE/uaHfoss0G+ljKciZkUrdTKVSy9hm
RSjcT8v43lAunOgD+MwOxLMmq66d35ppHe3Axe1lcGFBKLgZ3wqHV5Xtz8f2mYKE
cbhlCcOj8UE0Vn32VJMg8khJn/jU4RkEMD4TPRstqxOgTvWZQd6llemgIsDHsM5u
SxaHcSWodZu2vYOuPTecGbknq2LQ0K+HcJjN0r5AA2zUvZ9ue54/eZ5tx6qnUP1K
OdAhoYEjAgJTWMYerq7cFpqJTb1K2YZyvUUUGfUWF5dAUmL1HtEnYT1oJ2ttMsiK
QmKEJ3sih+h9FW7Kzug57Y1fI24a+E2XTH/Z5CiQfkwICMjVNv3uq3lDSdQ6mx3c
7Q1AOAQ37a16aOmM1l+/kkd7X33/SmqvGIq+vleeFlccq62YyybTDbyrNwXHtxW5
BIj5P9ptwfvweo6MWLVV3fdMIsXWHkeJ8uYFya4lNUa8yNhNbs3i0l+t+g86Idir
/sQ3+hVesUun+6ayimqmmCy/ao1XsY9YTRwL5ZVYsJZKCEqaGNJA9HclbF2b80Lc
UCJpY/H8HXLtUkiyWWtIQTWLbY0X0yMC3l2K2uI3c1MIOoAFw9Fr1VYjPv7aRPCN
MeBVggkNw27dvvDyOZQoFu7WACbG971jaXO+/6nCRNqbgaU9vHuVnhnIgMdwHN5X
UNJKENq9beHlpSLhcl7++fQ7SfPb3xy5ZTQn+1sTrnQzhKZzEzTM3Au/n5js7Yd8
PS0fime97/lqI2PQ5Ssb7kZDVAWypRv+AdE3mOE1XBx2NixlV8CYVXOEjN2SREVb
UN686G+fc2lf8j1AH8CA/s/6kJuJcE5Jq0gWx/7MgjO8KFSeQIJJTVhtJu8nkq9c
WawO9kCcTcRceAWpJr0GY0x03PRNySyLlDpgZPwxqD1+fmhBxiJUoPNRiRQwDhES
3UJ0u+PN490eOFucONuiifUK6JM+zYjoQIPT8Jvjh1nJTw/Dec4ADONfJnSGU6e/
FJRSe0OoksVwn/605xo7fMuiBSIVI6LrQLxrZ1Q0SnohpBmFoCpTUXpOAUoZEu02
GF51FVOHaYmvoEikd6t/YhhjiU+/3pvALJovSkrnRbkm7VJmynskguRukiLBQyIu
dV/D2a6MmJre+Lz5aad5qa4GMTHBjH6zp5y6JpeMW9A68PziMC80zzUwCNz+FES0
GsDfiX4URJZ6GgiGFne+Sbl4q7fCSgynLkrN8h+A6HjHzt55fq/uzs5OptdTQzZt
uNsbYHrIawQlvVIiqyuvstvT1zfh9DeoxIfUmi2xPFlik4HFt6qim7YRh6Qswpx8
ShpMN3X71u7pP3euOkcu5oY18f+c7G9hzKFZBrv9kRfT8PfYQKpKxc1CAO7R81H6
AdT5EZCf17LdS/HLvLfxQlpRumDPD43t3sRL//O8JhCl0Wr2UiQaetwf3ly8CbO9
0DqE8kZkzhYOzttTSZZxts4JV3Qm98jbaNw+XTANHDXuhJi42USHIVOU5ZHLcpCW
PKZUxUuEV9OTxf7z0zGrKbUDLUXtb96XEcuuKqRSboRyVynYqZ0bNNrSSM8+b01B
jHHpW3J06+C6++MQaM+fEmksDURbfgIp+3zES7inGedKWYYOFCDBxll3stQ6eluZ
0isdizlljqlSRxOQKRlUFZLUD0o3TM5R1Sbq9v1Qc2hDHfrcezRUcfP1yBr0gd7h
FAoah3GVMvc7QCFXQvjmo/D/EGzFf5vJkc12wDYJvxBuCgdvp/ZVbt3ss4GinImu
sOdVAl3b4WUMZr+QFXLmQtQrN3gtq0/yXEdGsENKZm3qe4U4cSslZJ0GH3SWdSWK
eqetmfAinJbJmnfGz0SqxvwH/jwFaCVl9hWJ4MUiYF0v2nHS7vPyPygvyv71Y9Wa
8AC2OzfA6rsnwwxXz0apDoqVvAcw0LhWRlpJn5/SYPzKeG5cyx4MHNB1SPVCrKxi
2rniWEK23ry/Redl77eAFk958yyt9WDEIXvP8Ge/8fZ8Dub3IUexzPZZl5wdgwBb
d1EE38upZvmYKAjWcguL8q+hxzazXtQU2plygyikEOPimrcYRSwRcDykys4KaIgo
AOXNRNhV6N0Cmaa4K7IJK4Kv/x0F+x6fb6KPLLhVRNbW/Fn+LLDim8Jx3hY3H+XU
VbRNicYzBIFpIeE80QKFB6m3F3KxO57rDQRE8N3H6oaVDvrnT3h5cdeY91Q3dZd2
RO+EPgRsDrsPB5mHucMmqw==
`protect END_PROTECTED
