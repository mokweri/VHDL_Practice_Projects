`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eGvmDNd2E62ib3+x5HTttSomNliOZr26OVx8I3pGGrI+J8z8WXTgGFzDJ4bVR8r8
zkp7b4rxyvvTG5yWuA97t2YS/lArC88A1E8qmbgYczo2MCfZtwLjAAQi1l7b6vaK
H3QTGy+0w9RgrSr3Nrqw7D7fTd7VcIBLIgfzxWa3t9VVWELdB87zBZqLmoFUT3bY
fTS/iGxJtJw31LdkS2lU2cdqL42zE04XLBcVeAKwzVf6x530c9qOz/dBG4jTej21
FfJOEU9DH8Skc959Idc9C3lao6et5Y0BpLPVmclj+NTpezM4zIux0D/hO3Dl8oAO
Kw3uJ8jlYMXRsAZSVfbSI8NnZufhmPvBVz3sRn3CJnFEvu97CqmUA54F4S3Jh21K
SBFMT7PBEjBMhJ8BzxHTSSWjL9ejEY+RuC+hrIrvjZqx775vmobgNJIgsSXbPXMh
Q6z12f3Kd1r4w+fLXM0zfBozc/lMMVlFo/D7BBD2+LLJZj/tK2aU4BHhdx3IUpSR
HP1VKr9Cn1+/bNvIOIh48o5GiAPNhsquPZ0FMkyS6rVYgO0+IRlBkmSkl6bzqdcA
KBhryiTrVyxV3z9wTSewHbMUxeVv4kGh31ZQR4qxJselhW1M28nF/pfBL5kRPE81
ejC/Iq2iYcdZurxNphBunI9FHitLKfjUTVyYQB9MxC8aIem6ke5QCysZFxtCHtQv
mBKDHlG9JRX7zua9b9qokVshvYk1FnceY/VSSQSgvrFDj9nP7h7Zak7TPPpLgJce
XrSteKUAX56IR2W0X+0O5vN3P62wAdTF0g2xCjV6juBI/lVD83vM0Y2hWR9piKvl
hlLqaandnCIzSM5JzCX4/FROVjEpJQDKr/kQ+FmBCUXnRRI6aYZbrxvKsUoWlDZv
6IOwbpxrjVVqOdz+X9QYCpa3B2+QtRSMqpjmHeFnxZmEz0crtVfoIndyHXcaGmr9
4kKbOAcPpkgvK4nJ8Lk5tEFxBMdDNNBtm47F9vTUfy5MsYK33/xzIyS25Mw9dvwi
b+b/bQZHWHCX1jn5exYLix8JrfmtAGMPpclz7xXBKLTLcIA4VVu7kQTkOkGeh/7j
vHI9BbEuxTsKDFXyU1IWKUbCJ/Hdj8JEZyFyk6pFsFuBSRgZIYkrsLvIfQYpuNz/
RGpjnQ382ry5FScXIMceeORs6VjKUFCs9kTu1XawYuqX7tNuD4w69AmVgjhEXrLu
zMuRtWP+M5wh3CSRf/Fqxwh/5LyW7cPJSLCMW4k768QFbxUsCtICELPuHbs4xQiJ
xQhZqalHKrPAbBq1Dq4aCmADyDMrpb8gs/O2vy86sIEjQSxOpMsHzptdsS9Vrm5l
vK7vnSdKO0C728Hvrb+khJep3MoBHYGJ6RsjZX3EdqFrOcaH/byhZIr41tO0XQL/
/4CcVvHH0kl91hIx1cS+BaxjgXF2oZyFEUGePFM0yvQcJlt479YpJ0oU1TzeNs8R
O8+ycbp3X/rshBgbGLI4TveHC7itGp52XbtxFE1cMd+ixQB7X5tcsWnljYB3RIJC
jA5R4OrA/+zwvovMeGFCM9tBWFprabPOJZDVm0Tc9hHaYVC8k4zQY4PByEZYLLGl
AnE/6erSLCaS3sBqsJg8fXLdY+upYy2JWLB+U4QN1gePP0fN6MTof+u46u6juXrU
HOLhRokX+UP3uSb8WChcRqC9ZPpzxZ+cDLfV5MkbgvR9pyJW+SzOjI95g6w9Q8hk
W8rn+vHTXHAf4aoTpc6j+aqkAoK4V71TEfBb33RfWv3+Fkn96g6OG8PwHXoQPPKe
m1EY2eJ41AjGgQ6PF7SaHHOWjcLnXNkhhRrXDTnUex43HBfne0TVUFwootk2nZ14
1V/xQeHlxdLunI0ll6Vmj9xzQvOj9sYxaLg4dlGnitpT/R7FQSitPA0eKELbMD4v
5JEQRb4hD6PjJOIM3cDZpJa/Uf2L1QdB7wh3gBSby8Y3q0REE2b+OWfLzfjJQJaQ
gg/Oq2IA2D9qUlmTpH7RdiST3oYjf/s0G8GOGH5wD71/QuKqsLAUevBiGewcZ3r7
ZsPjYmvTNjkDHnFJhAQuJMWU2ZieT6As7X+wD88dbLhdRU2n3umda3HPKiHl2vRa
6YY2qVg+fQ6yqoJwK0oFzllXcITlnZRnnXvnPPSiNWc9mxeKP4A2U11hMl5Y2mD+
WwFAHFD+iEJihNz+B+CV7oUQESEQTZFnGjeUd9jKncGFuHEURtvBLBXKro63wOUX
GxVwWO3xoQ1n1M6yurHUN35XZhtd5bcpxicmU7Wqb9tAcmJVkrH28PVR6HZ9jBm0
nbburKfNuEUg4b8VFfF+HOPaGRX+qg5Hb9GBAiljOzfyJkzzy3o4YqAvvJzJda1b
tpnpEhaeOlCOeVGeDFseYGAyPoBL4ZwZSw/oZZj6Y2lBZ2XdEdOcGZG/17lI5zJ2
2LmiiczVcqrM3eN73X/rl8OmmIVkEVL9Vd+7Pmfo7k5dB4s28uGAccaumXa8ObwJ
XPBNsBz55NsVbFBr2E41JCYrnSpSUtLWyXNL5hadhNaZV6UcstL7I141wC7i865Y
rJNrQZSBS9wQqTEzYnt5q+989Olc6xQzB/o6iBTPKdk2szgcuCCQsL0XMCMhcsbw
WLTDZAiw1XU8JUvkcFfe2kQL+h7kOJt3ICxIyqiVDO7CDzDazb9pMMihxrm+q4qX
YciU2lFpWtfv/ncBot7ADfF9iKaPmTH8QXm5TOjQZ3KqXEqcGj9eGgDEGx3A54UI
MwXrZTMWdSkLfXO51goRriI/xMXT3pDjtDqD20kCTpQclzOtLbgZ3TZpXaVBkLeP
c2beR5GYdku/p5tQ3hp9PFwvaIDy01SWphLZ0SF1/4/O3FFrDc+y6QZBJNpyfSIk
suLXjpRbCst7YYPVwOuEbxjSv934p/hPyuTkplUBddBHahm0Wt04zuyAMvISk8in
MIhy943JEuo3M4OLriK57ZKqzQTBsGzi4yVsOUlKFaq0ip0l1niF9ZE+KMYqsJdU
I1RuvWkK18bOXMYL/8YC9hgZFDsU39gY7K3T6BiFF0gzzupJKNQZ3Qnn/bdRBlUi
WMkz9b8BoX4qvnB+A1IA7VHcVdjqu8zS0C8XhTZVHLWFdrMA2MMtH/5Nx71JllAh
AO9ZjHluaubqvXOAdlA0r7dUn1KLVG9bRQTecZmUzuzVTcuWWxBNoaMEhTGRbxfZ
JYennplf8U9OuYemgjlayOhyMw5xKBFb2j2nuuX+YPrfPRj0broA7/tlTXgpKf3N
BwYAB80XJ9lQ6wmW2XWOGVyEj+pjSWb2tcg+B/bgh7Hyb5HGM8THphTsuDS8vGHt
nTjqHteCrNxq5HDcxAF8OuCchipV/ByGKMOw5G+5fIxC7G/4AU0adE+RH73O+ez3
cArnvopPCoOE2JluIT6iygP+wreGeNwm0EhQc4IgAVIxwxHbLYFE+VtfzDzdAEcj
UsWBsKnk0NnOXfHCu18oI9w5Iz03YYJYfPf5lE2gthHWOWah5bCmMD/xNZsngD/i
+hxhFXZyp52leLxMjJRkXjjli13MDB7uF76K/4jWSzmWST0xSKjQBscuMtdGHv2f
HYYqK9SdgO5d0faHvjNQirtu46soVg2iWlR+HhM9B9AQqIzdYfbKhPfDc4+tf106
M4tmopkzx2PMba2aWmGnmBh7oRSussRuGuwnPzplP63E7LY3mS7JPAUJOnGCiqUF
2swsqgWaV1ygmFbWpbobCTzjMg3fYrn0MVVtVUD4vlBa4cmc5E5/e441g1iD/8dc
4dnGBFobalFQgF2fpthK9swz0oofQO16siAQP/VvomAHDOgG23AjPlahpeG/F9tS
8qSBAJ6BATV3+VxjPrhNfib6EF7fDGCabw8+zqMDfxWbR6itLwdpEBvg79A/MAFs
oDT2ULFhTmNS+U7i5WaO2WQL6iXsFYVU+nHcjHkzRfQyCJcNfUbWIR3+r98QqVCM
obr6k4QnFTPF0OuYL6jUoQN3kR213vZAmq8uLdosiIGw3wuuwExdD2WXezKNPc7Y
M0Z1xf66Pg/zKNEjrQ596N0QVOGC8wU/6XCV1aaTw/1UIc85Xhc/SfpUJ8Dli2eu
zxm1saNB7H+aYzaE8VYSFKWlvEiwbDA+UuBZcA052BHjcxrHbm0c4Wk9rufvyeiK
zY3KK+Pi52Xrx8M40V6GPKg6FLJ421AQOv8D8EHIA3T3rdmF3vfWYyveLGMw1xVs
WXJLFWrawuw9eh09bYxvzE5bl5D8/BMZbtoaVOfdnLxpCb+HO3z0fIADSp5N0a0t
yaE+9+0CLYdnmcCvmrmlCzq/W8kuJN2C584i24EN63E8oJpBsWl2B/xaQUDHSShA
GCjVTt/86lNj/mmhBsxvii7zMjYCoFhCswv/1z2ropGQGoDSyAxaqvYVjE6pN7c/
O7T6oj+6xkns5W9pNuG0rza2Mp6a5zliW+z2jz86IqG9+ykza576P0tsqfZs2Pzz
WP4Gp+jiJP/m9KbaY8Z7lDGxtXBd/GMJD8Z46Q5WKqBSmHJd2qeTiASpJnZ279i0
874K8t2nLGaP3reKNhNhQP+uVjZEgw1tHQWCCNyxQPNWhdT7ynq+D6PqVMVeUZvF
Uza19FLcvAdODJO/Gsz8Kw==
`protect END_PROTECTED
