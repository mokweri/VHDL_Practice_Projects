`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3r8/mp15MjWrjOYyetKSQWjveqTi3bqn+3uQROKx/AsUREUxv4iXSDMkQtXSbzR
dGlFQFN3vkqnOqeYCZgMSsmPHHmZ2UbET4FTJs2WV06GLQYRx++qrElWe9A+yY4s
vPvyG26Ux4KdQlktVU/GAPcrne3MtgwKlk3IFHOJeGuUN5J9d3AWSbxdHH9DtzCV
GlL2svfp6u2RvGexUV6taFi0BluiTYeCoH4Q8qq+evxqYEq8nMtxMtpJ+rsfxl5X
rJyu5j7CUZnYAfdOkGhYx0WRmq8EsR/oPMQgY0AW5h4DhtzUjZAQPy6p4JZ6voDN
tDLz5g3EZu63FVRtKsWcvikA9zuxrKMcxu3c5raoNnik8thzqrLQ3RVbU54FtcvA
Gj+PtjXJ4TO3lCG8BYUHRecjPhEsQg7D3JNUANKseaixhW0zH2r8v3NWUBu1LDZG
PFC/2VKqxdnniGpPvbm0FDWSklwPNmy+FidtO4AVQPI=
`protect END_PROTECTED
