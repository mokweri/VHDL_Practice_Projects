`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ikw8ioYPyC2k4k2bFq7V4cZLxp0xdpUJ1RE0EbfX5lzarzK23kIfkWfeNur/v85C
v0LxTEWKsDbeGZlii/8gUaQPjCPIVFoLn3gHvScZCOfaskAmYo1j+Jl+02KZSOsF
9C7QkTkAko1brfMxFI7GhJ5/zCvNLb6bk24btLvJBviG6GMNnCGpMGiSArePcz25
Uh20/ziXgoHXa+Mu8H6n7Iln8F5uspSh5aOCFsrIGTi3Z2Z6wok5d6+tVHrx1bCZ
pr9zb+4SrPlyCUxKXw14h0FYnuPLx3/4+agLRKe2533WLCjQ2AM5Pc6txx7TK515
Ai9YZ9fpjNn5P4ucpcC+pPSuBWcu89eVX6R2SQ3evvA+g6oEUpqpz/RIvUmDfjer
aSqVBc6ot865M/jHoC3IFB2BDn/t9i5vCrTSGJqqlRLYFq7jFmUCgMVpQ/rlmPxG
3pBT1K/lSljL09KUMrnW2yjNc8Rlk0S/RdJ0Ri/WPJEXUSZrywLWmuFCw0xyKNRb
bl1PHlE0GBfRVE08x5VL68w6wkVaKJxirD/ygVlc0xZr/ZuwNvVLtONN5CVk5LvO
0o2cC3+FaavsWLc2FzgFEzibd1MR5Q543hXzOIZLDwbcsUG3Xmm2N39NDiTFeOKu
ahEGabUqL7PS+kFTj9kN0pvv46tLLYoGfMWhMrcTuIjkqJ90LLtmPh6Z7AYs3D1d
XpuNJYO55dn0XBbF9NyI+ogfj1ya956eddvheUyB/9TioyjG4vRlA5it51dY5Gtk
ACxABDLiFxGFzT6rSkGqtS4O7rz5+TJmQT0WLKzEGryFkhnToObzrroCc99Df3YN
5by/qovGFKID4H18MTR1lIILsPyZLhXE16LnsoqsHTUC3ktBrSCfqVikOu+ZWUyn
/hJbHa2D1N8vGWU7Ctu97id1+2bdakgI1B0gRf2eHMZCpoGMFBlaQiLBeu1Ii5nz
MtZDzCkqLH9SMZX66BjWn+Qklk0yWESQ9QEHDtWyiEZHcLUpKuqa64Yd0z5w2VQK
vZTQ4sG4lr9DYeQodOBGY1kwsgY5eY0I7Yg9BVuB9YBbZ0IYWKyEmDhN55sYzYAU
5S7vsFhVma9an2nSL2x2Q+CDsHwEIu4SZbxYrlc/VluA4tzEpNopyOYh/irgYC6J
dI+oibu1cHul8cHhxNs0HTHwiT4XU7nkFH5ckg9A9eSTEozJCDlBMLw2jsXzMedI
OcBp2sYWy1D8443c2j6rFwobdRSq6d7tEHCYiE5/uVnJtR0ZFcJgUDYuGbPIPqWq
SJqjFv26vHb00D4Shmc3jPMnWBmk7s22Gx7uIAMzvX3KakrA1iezNlGIF5+Usjpf
DJlDOAPFHZJjojBdT8NnVQCctUmkom8Kzcz+uHvPhSFsm8pZAnCVXCB1drNdk3+7
yVu2Z+bldC2x96DvOYX6HT8zuk+akEtUhpSjqD2wTtjmyE9jnEkM+1fKFCruJPXP
MDfTbL7LIGq9NpqMmzAWbBV8vGAJ/lQ9J9NCmHFRd2TNevZ3DV0YK07LW/6IHJsr
mUxmlY+NhYnhIQScH/JOk+xKnLxKumB34Gor3cV267I9HOAUb1qIbqiyc+gQ6+Uv
VVYderKdMgnStRdW1WReG6f37dCZxJPmi5wLryEDzWR5+v6FMP9UXHyyOyYWQbSY
OzfJzLrz5MuDhbIKIx9BhmmQSuR3qq6gvpjr8m5nzH8YcVONgS7ZILa5XUkugRbn
V3ps7txC4zkZKXO5uVN+VeTI7cZcb2B1AiTy7VVumGSasWYlrCA9FQw5VYcxdh6+
9p9jkGjf+gnLtJUX9wcmxQ+IbCQsDPYTxevyYDX7yZKiseZ+91JVpPv8Cf0lZS7a
muVIR+XEVLZ3Jt5elDnfWKCBgC7KA9RQVTLDBtWlvbOlzKXKTM6QQmfdSVIW8oNt
LLYe9rfEVPpWw5UGsG/LVaLQ2T1NaIPrhZZJZ/vaAJKysU61zfKg5fbtCrvP10am
nAh8Zkk1UrWr0n9Mobc6Qsr6sZv1TLvgC5xZ09onEeEYutxkiBT88qjY5ULQUpwS
mpIEF92zYjw0pN8XAzYCnOwgPtNwkdo5mYf3sdAduJg+bJeNR8bnh+to3ZE3h5Lx
UV0owqM7BEsyHNfK6tuV4+OIN6cjhimHK6jYtJml6ByuMazm5HD/zEPao1/O0uWG
vAv6PNhhCgtF09WAL6092VY93GNf5Tz9IHPgNqek4iO5tJejJx3EmVajhegGNOEX
tkPIDwJ1hXwZcgYhuafzE7JWjJAvZBHiphTDTiOfhE/VSv6Ac1gvd+/h5fuzS4xG
VbQgT3nUWZASZy3fEuZODg==
`protect END_PROTECTED
