`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1pkpSMKvmwy/Nmg5iiUZUMcEcz/Je2bldptICfDq/23rbt0a7FeINb49H4KcJPFN
aKZcBvmuK7I46YNjJicYEYI2zKWA2+cXlGKcDfd3hhjBag5pbxMW5zutjlo4tSYk
z+qynIHT2aBvgR91neE9DpxFU8yrBVN8cKXg+f3N8vPQ7ukO+w0tgNsv+mTGkUlK
lW8l5fLB6tog7jjZTUbBGiZRNrk25mf48RdiCSUDHhY3glu2E7j38ZnA/lilxjeu
jPIsQGEeFS9xTPl4wuWCRLtng77sRtTF4MHvp9AhVVz22kFUtubmSjPAU38xeHtE
nuYj52Wd0U7lD7eI6MvGeQwvw00pEUD5CQ9PZDWsYV1c/GVPYFmRdjIAnuBqMcPB
JpH9ehzYt2GJMML0b/ynPxt239BCpYQrU7pGT18GhV3Ce3gu1YkoHNV3YaO+9Gr9
QqaB54+BA8SX/le9mNo6WnlQ1HGcEll5huNE4Vlp2Aq0c59Nr8AQchBdeaunpqo2
noRPcu+fkiJPMZVZZyMqgl1hJXdlPmZH4y6bvJLzdBeznyWKUPxxzSMLBt1k3FSF
btEQ9KxC6c9Ydl4knUxCQq2um9eNLpj7CID8R1lZsYF+U8RHcxHxEin/j3OkHx24
F86PZR9IyXRr6Zcse5P+SGSLqZE6c2StpE3KHngHt4txzsUT2o/WeabsiugbDp33
r4Y2RM6yhOnInmzhuVoQkZmZDjZAaVPfBbTiLNLu4IQvDnYUir0kxd0uk9pn4c0F
HoiSZ/BPWuFqlfUdKWnS25DV3EQebRldd//xbexFm4cctrpdtd5SoWHjgbgMBs9S
Sq63y3jxBLNyrjFjVdqBGR5mIjyXE1U02+3h7TFMRxSWqkGBStBURtG9jBF8YlqL
kOYxCwLrokBCZjuEVVmq56l4fsNCTMoBJte6txJT3RxhiKgMOhlUVvy1NEyeoWhw
DM14a8wnUK064ImaE1O0MvJ7O4xTkPD110pMwDAveYnUBeBFVAD5B4un0vpt1YXv
Nk8xxt2HOrYJIUPH/kz3ZIkvxSQvYM6YcGdPhAf8BysXMyoSECK8PKcdJCBA0MIk
Em/gH5376HVb7NM0TlKNvrs+0fz1Hss77bc6hFr2Sz2EBW2OddpPVk0HKFHkz64w
E5LDOa7uqnyfOyeO9fFb9AL8RL9/mUV1MObiYWx/1k4w1PwBPuLE5fM8dbNDzhFq
6l1HPncygWo92AenVJt8VIzYL7LJH0sx14svkWFSZdckg5ZXIvnXrjhVvqrfqcus
CY2tNg8jQUhFuYLVYZ2Bq2hw8KnUX6WftpEFd70SzMj0qab7otuQ7jvr9Yq6txqS
ErPyoQQ4cWEAEfwnSAL7f2JG345fMPXqWaQUvY8f6nUtTLx7e+0oBh3c6LX6fyho
74amsmIb39xCBMH80PkIxMridIYDlwCiyuigknDE3vXwwlBbLSR8sO/sWcW1Rf7A
`protect END_PROTECTED
