`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QsocQGVu3FruO9LIQcFYwM6YsaiDQG8T/SP01q4z0fQWtG6GQwjzyLTulbKDWiyU
gHGQyjL22etDqo3qaWTcQiB8vcFKYrr9EuE784/UDLxpfJRs5ROuBJnZMx/vUA92
fiszXTrNKL1Oy1jVDjMaHlxVOxmCq1YZqKjlRay8d6oQgQ5Fiu/LqmxiGhs2rZ56
hyJ5Vnh2u+8j5oNAGebpPRXMO2zRnfRGu4Ws/PRm4vFaTkt5cFkwBj+cQBx8u3r3
GAPXEBrTWt1s6o4xwfFyXJaqZ/2gPdIGzc9iFzdjOcwSASS7EpXc5SRdulZStDq2
9NPiLKCxi3vQZ57YWNp7jWhO5hTpf9XicJwESSAXLS67IYy/bO9CwYRi5FDMiQlJ
/ViSaaLE005278sWi2aAD0XBpCEMTWWRfAYDey9u9JFtBuP7KiPfSRBbaI/q8Klm
Cx7XLv/qBqS3o+PSMEUivhWbZk8klIiUE0N6CDiqRx8vtfajWDVAoX0pFWd/FXzs
ezvl7si3Z9xK4iyswESYWIsHQsc44qgn2ZBIODMIjEbYDe3TkfP0AwgaRgJJ4QjQ
LNA+aQrYk6+aI/anG92QPSa+V+XriF/9rkG+KnmkALpn7Q7IhBT8rjjrgnfPbv17
IJq52A16yFSolr7huhByxzB7SqsHftGcaM6WRAqqzNkZxKU1CBko6cZG3+hjGc+u
1nSdnHJBYyDaXk2WQ707GU5lhrweqwlgpHEEq6sk/To9pAjqFAyjM9ROZc1AWiFX
0r2yuDqPIcNNdxHmbB4zdjiWs+X6JZqo+6P8v8L8yq+VwtqTuLB/Hkkk6C9zok68
vWIboYw/o/LRujA97yVY7GhFVYrvkEHuvwgKN8cNyWjcoFgYWVve0uqxWBV2I2Og
KwuseGi3JXFVfOL7VCltGkRzYtf66fziZzOgx1wxtDZRU1yVAEWa1huwAOBha8q/
rn/NaQBjris7l0zEM3VausEle+ywyLYK+Sq0o8AXaD4GBhBop/h4PnHT1uY3676a
MIVeHAs0BRA/p7nXiW7HEI71qc4UqxhxHmiB0PICTjlXjZUvJgk+V+sUivv3Q4be
PCkvRKovpurKxRZ7RRTHXvPI+2lbbT/ndF/jMDFB96beR875xloA4Mx+X0lLH6HS
QOiHTUX9WoEquySOwzkGVFvHFXWiG0GOqERqIpYeTx0TTO4NEFwec1Wy2Izi1hLb
syAfRYRGgTeNiqZ6mv99GguY7J4Fyoo3xNPTxxUfGpGblz8gnhWHKZmeNGF49TNd
eRcsI63JQFesKZuWTp5rq+EN7skh/KELeUpih5rqRF0M24sc/BGZAzxVJdtgd/i8
BWWkt9KasVawKoXe+uQachVBU4hv0MAkchnwBsnG+SRsuBSeD5R9EUkQmo+DBrJz
fMeCuRnJFTqKoa4JeiV5rR4MNHbDtTabkh+EKcMRewxDtCb0FRaKBQ6k7Ru2mBXO
x9WMBTxOM1BLqUtCJUMhhRZfL229J8Wa1P6w8ODC62S16T/VTq1xUo0F87WTBxhf
+3TKnzz/MLEXg+RUZEJ6hPqDQQmPLzQ3VTPzHdtzrehersebyLgrAcpu+eQUBt+f
HJJW+eSe2Neoj6hqTBxsIyBBQQOc9d5uRtMPGUlLiyrnttYVjaW8al2DJ9df2k7i
AnOR7HsTq0umYcehJEHmeqGJzgjxxtuTtwREK5UDz/4QkmpFe+iE8nufdJalzZgV
6eS4EMncfu7KCISkbwAecg9i9/ZqmBnZ9kV8ZzCiocw07vR8b2DDFApS1IrCS2gB
y2P+4sf+pfRRUHvnBdsvEFNR0Fw9Su4bmO+kor7zWSfFhhIl4wAPBENFMzKj7jkU
Zt9L6TBgQU4dj20VghZic0qo0jnyhO+tGz3QPbJrijzKz93HSzJmq6537sY1ce6L
tEhJ6/qv4jgwLNnx+5NLBRvREVbrj1/xeDXYahSLmJ+EAleitp3lC+PW+nBWXR/H
G1d6LPxwnA1FGV3wMGNwMmXb0Fy9dq0WLa+xtJubQlhsTxbRYJzlQkmrFe5GAJ0V
L/pfxx8bdcwDIEvlPmrdOS10YZkxa1VIZJzYhQO8kq32bfT/mh6OjctweCDf4JM/
QTa8FQgH9TFji6BKyVEYlsXaFmNRq/8IZqMI31dIkwA/dFeAnz8Npxvr+pEHcm7q
QNe+bl9Cg7TTUb/ESjZwSp5sLFD+14H06Qt83tm3wNIsHYPiPPj3VStlSxNfhuuh
qg+JmBbfF4isuNE9lwJuq/Cv7T6dSYVEzmJS/Sn5lhpNrRD0UZVuznnNznfR1p4h
mCWlccxwoq0+XsjBDrwC5Gh3+8lF4a1A3sc8u+AixBLZay3EGEiKtTHiQPBTA6dh
4zaGYUvutENSlUpoH/kwUfeDgs9S9uGrZVzKpLt0jX4F6RjGMFataf2bRO83o3cZ
hkVoRa0muEa5f09RK6+gkXRPO83FOy+rOuP6yVmhyklrm00xKQGJWlD4Dpm09K8M
w5kWLjmdBad48XzGmeuc0IvlnfBYfXBSk0BeSlCFAYpO18xuHWlGtfpSkGMlDXrf
7ZOc+KC3cDHqbWqjazmc7DudJymHVlqfBOqwktjIt3vJghWnFqLS6GctlU36Njsi
CcZGo0KIPUQC4Lu6fkwOrSd3nEK9q8Ub7wXaCc8SMCdP33yG9IPJ4fi6aaJheewd
qTtIFKK20Bt8N6Iev29z0CKFlG3e2WckoiIYDGv2pjL93r0Hc3ktdHRkdCwlwNAv
0/4jxj+KoFtZ0go38akz/Dya5YQXHOpkZr/Dj9rPsUKe/sIYukfPR6U8fBygDKfF
v06QbN0A0wKHXqF/srUml0GerCtpHIcR2u99sfA05xsg3y7AESu07/4alekI3lTN
4wi2vKbVlwA/12g1YsXr5zF7ZL686/vvXT68B78+teKyx4zVV4eRFglOkApDdAnr
Ew9LtaT5jctrEwLaMskspmQd7Qj6DR8/juFPMeCGd8GorZhUCgpTcGZ5KZkQNIkx
LmGg75Obq3CWwvVLJlZO3tLV+f4Ic3zW5j/U1o1TAQzNCk6xdHkF1Qe6dEtUfKh6
wJzRIPDvgse6ZOcwHv5WtnGOPAswbQFh/BtCEy4AqGIdP75jMrvvTgfYEoIhcx/o
yTJI9Gj/BgZUZ03CtXJUKfQXS70zeo+8frgTGPoN7L0qbaifQ2nWY/9MqT8M+fYx
w0gEDmpLW8GwrYzCxyHhtvGYrridmWVNiSHjpy9kYLmlibobKT4XxJcfB4BZzPFG
HOL+3BSB8BgLXEMek7udwa0zE8yWHjnq8n/JI5H6d3y6qivWB+X/zPPBT4hGc9A7
02mHcVbHKsBTBCgpylgq/81VoCXv5n7ZxoEX0l7Rbx01s/NYHJY8C5PUdYsIdM/l
RwH2DBDde39tLYedWhBFXqNAQz+rxxpJISqIcpilf/2wL4ZLgJkkUgYKzwdGQCYP
xmSzYxqWjlEZT7FpCjnlu2Kc6zZ7wua3qizdBoBQu+EsLqP/aY12P2zbPcmABnu7
JZ3FY1w6w4BPrCPz+HtRkYbc/AxG1C1p0axdpSsR3KKWfS38WN2zjffT5ziBoAUM
CO9dOe8Las5Virl+ttOPggx6mGtaA8lTMKK7D1POV3LghqyvxwfQDU7UOtS6TKgW
zVpg9uNcm11LY5X+7jDT6gV1QzrbnTFB1OigRPumF4qqT/er9Wxic7ljk4m6TYPe
VsA1Ww2Q+WI8ggBt1GWwo3AR2XSyP5hAFTwu7ngXLtC1tjdfHIwPfiRb/wpWJ+mt
U+envPEGh1Y4QW/JbwhGRIhkBKZg+IxEzalZ3U4ZXMRZPDZiJFXN4VopKG9Ry5AF
z1hTSFf0lR5v9k0J8ufMC4V1jP38uIZJbqFqq2Y55PXRg15iN0qvYAB+af7oZAY8
+19y5ydifGmeVObgU1w3/bjEFUHWCdaFQ4OQysj1SeV+3t/zYHSy51l7u+HkuM5R
0R8MF92vrrO4tTvJO32Gc7AqSWZKE450xgX9dpSBsGGBFbggYTbToZULx8uD4Hxx
fEAJh5W8NhkUp3xqiKTVHAvzV7g9gIVtY0J6L2lhNy/7LhrZ/+8ufL3tv2JzEmcc
6WUV20w5/fUltZsH89jt0lnsHrgtvB3Lq7MGUh/cilq/kKPolFdd6/uS4RbJwL/6
HB7svQqwcuMFS0w+a6pJ4Z+9xPUYhC+ADITRV9dp3Y41G2sd/WgwEygliY4KM1d6
xMhhdEY0aAaQJoMDkUYQBgXhpk8i99ZLbD4n4XKMIMitbZgA33JZkvOx2JcDsb//
NPczN8/ICkbCrX8YmizcQp4QGETqBkveAqoj6col3AG6d/TkvUyGWAxD+OTucdur
QbbMHT4wCQrP5wfgOaDXmtppuNm2MqmhwMPUln6U7hdrfWeRp/U3GnbgPnPSNNWw
yaWfFpbSW4ewzSQWVMX2ULVrxNNploXldvAMotvr86mYNK/uCG0QbtmL0RkGtFFa
ogyXGnOwtK8I68KXoyI21srKW0Q+67z2mVDHT0C7I+/ASPNSuIc5RoyQ6tXNChlw
uUl/2HOBebpjMHFujW86rrAUH1TlhcAtwr21URe4fBpTZHMclRDj3bVKwyKhP6f+
lXBPQkPMdWxRcZpM39YTVArhbh6Wj8TkPEs51V3RYdIs0qxXnwTEzRaLBQvxRtQw
1VOW7eNBITimAADj+n4jam5vrmoEGuO7AGuVnMMSgHPOaDzp2fVEUqRuIQeLDYFh
ZJcfKhPVgypRufIkwMAX2q3nfFkFtH8BR05+JUqz3eCjncKjOZ7OvefaifSSVVDz
LHOIkA2eevNj7fzAoRGrX3j2pS85Hq4PCWMeY4McwrHfXQvdqDicbtaM3/6K59Rr
3MHN44QiSZ9IO4L3Z3HRVim1h5y1tU+HtV61DqDCoe438U1R8BblaIjpHRO/w0y2
eZgjFD9c23GjXpXIHPZVgs9m9kidZbQBt4g4UV0xsVueo7h7U8RfCbdrRTyo/Zx7
GormFNhsiIgdWr9RoKJGd56vt7HooD3p5A5Gvyip8msl3DFw6+NqUy759XgkZks+
SZw523XOSY0FxeUOUSx6j+SG+uXRKuqzyd+x0kjXF9jcDxjoRCv8Iycm2vxchcj/
l5xXO3kYEWzSHMn0l5TSxfQT3m6fWJB699MWBAToVK9Apejz02SrqLe6wOTQKqwt
TXvXzpE5iTboGyCC0+picTmz0Q4rnwjAT+QdCvIoZ8U06QoYZNkynpwAzanvQ9Nu
2cDbU3wTDDZSm2PdBsvO6hUxpGnEKTn3hIyHna1aNJuQTt6E4XVPgQLTUBZ0Ksbi
gb4La10TAifz5JWRP1asMLoQ2T8L5yEfLmmx+UjOfcJ5IKI/MK5Bg3knSDvUb2zh
PW6jmQ+sAy7QuQxJ+M4Dh/ucIvOM+/2ZnRs8A9wtlrRUxfs7NdXbSHXb6B5+Oga/
Dlw0g8WyewddC9eoswPueHQTdLAWSoFZodkUYtDXb+6sUfBGLf6e3FOi//KnD1xE
M1od2ZtSMm0fAJCpEV19+CHDMdqHHcFTQ2neRkfhxdBhkZyb052+VW6nrIqP0+HH
3pyE3mcd56F5k3M6ouoYTwROcUte+hHWDhS5RL5b72MV59Gj8gQm0gzd0XGCveBo
Xbw3bI4rrkkcrJgeOC6Wdw==
`protect END_PROTECTED
