`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/RAVE8RD4FNjisI71beeuy37+RuKTvhqWvcDQC2CTY7671qn9mdsUL8MVwTbLvB
6dUeFejSHqPhSxuWovc4NqcYQ2p3ci2ls+zKr9Zs6VfHqLmQ/uW3ugn3tM2QN3gW
s6DuKM8pOiZJe9TUV1TPIK0bG5JxLamZ4eSSbId1bLPOEG8olLD5TlqGdoKtQW4B
N0fvoH0lLomK2XDMvEKN0AtryD7lLymj24x6mB4bmKT1qBETR8qpjzvSomdbarBr
2A1iUJ8kLqSDDr2+TXEsmj0SiW4HNDpUE4w2LyoUpvR6qNH2Fx5bhUDUIO5kZ8h/
SECK/1AXwJWS2F/cMOi+nhAsIIAVsnx5bFhoJY+3opLvtNWUCczgWRCIFLOzwqrn
C5UA3DpkvY8VfOqR1VgR/W9l7xVUvwibj7CcXyTTtdh4ANq6xhEW7A09qqFm0FzH
Y0QbzqhovYHvE+Gllj6x/m9M55Xpv7jWsbKOHHwQvTGHQ66CRbwWKKZ0UfPokzbe
qhHWwrANOm9sP/w6gwbvbM/ReTmA2BsP2BgEZBH52fwtIPqZfT8kZ6/O2DtzUeho
Z4FdlOQEgzi+UKamUaJBoMn4i8IkexDgVpd1FyVbTQFbOJaBLox32bmFQAmILor5
eUHWHHoqfqq+WXT/k6WG0Z8ALTQMPA7RYatX7k81tVN8Buup3IRImXaIgZ6T5m+R
4MiCl4JtzGvp87oHstruPUNhKeMsCtJ4BU7CYIDIKqWXAUVngR/FvOL6EYjbwYDe
oPlChDuVqxyTv4m4MUVZP7sSZAisv8EUK0Yc9ZxDaCLLZi+/6sK5r5gCz0l/73zf
CoQwKHUA2NHh7h8DMdM5B5+Fb3MnEXqo2Mqyhqlma9OY5f85SV5vxTDxjnqhi/d9
wcm+c+IaSqw9NP+rlFmiQ7o8HPtwNFfToq9OfIOIuPTXgeznLfwmpeRH3UB7M+ic
O0lfl1t5hFhVIaqXn2GAIGO1mRG5iaJwpWYu7MD5BGOq+r0pSwUJsaLMpvdw7+Kz
jgPFZVY4dLbMlgefS8PDTeTxnfJOtVGhq/nDdT1snxthW2k6pRl+YJ+RG8Ot+B7/
AYlEVFSMI3ySV7IqHN8C4ZO5NlxBS+yJo3v6rUC7A4UO2G4XxF2g0UuMTQE1/9YF
aUYu8y3DcLZX+ZI1HpESOi0ADK44dfS/9t/KAclcWAOJY65pPRL8S4GaTlER+GDS
rP84gtthJ7PuPRIwYPsBCFJgtjDJKG7/n+hxOcF1zp3pof2+5TuuIk09AtFaqRyq
ZSWBslEoiYhFsjum6lmSPXxkAsL0fR+KAdkySee+2C82dcQSIdzbMlQYOc9CqKBD
/W7HW3fZnyRIbQctaPkVUIk8ZBr9ELXkPY7F9P281xYSC92lHkN0rsvUBIhOxe3N
zx+bGXKYyshIdipeWE4IRryFkv3PRD5qY1b97uox6mPWGEDga0SToqyVBXxVZtJW
ZtAyrP7//7sxyqbi6EyYWc0jbQh+53FlCv4/jYJlM2OIe/dMp2CoQGQ+6VhsHfkh
LgZnzPQeLNhSR15qL/IKvEY+JT3OjaJ5wda/8zR3AIX74uIsZ3fJMnC1tIT1PRd3
koAmSx9mtyBemGTLA+xd0eIjH7jDcyeF9tj+dSqtLVhM4d/n3Tzqf4EFr4HCM7bD
xCxEmz2AXatAH2hZPItOTqiwdv0R5+e9mKC5W+hlehU=
`protect END_PROTECTED
