`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdC/SheE9/XusahMAvR3ADTsjQHDaPptxqzBggW/4mmj7/5kBinXjbgT76l5/+Xc
SVM/GzwGiOJ4/d0xSh2fDEZMD+8WwZofdeGjBTYX20PXRW/hJ5szTb/aYQkN9voW
sIqeA54CSW4WLPTE7xKTGIYpyQPx23KGHvltTwgOReuRsnGCiJFDfmN1e1Pn/twz
2IGDBT3zeiL7ee4B636JMJp7jKQ50idhSj8G+JPBiAEHwnDgmdSwmcRNhMcCKc9C
dgExWlBiS5jIclSXDhwaC8yfqKwkrol3ko8bYeE7zq0YC3joiF+AhoRREtrZbHs4
zbjssjTGl1ZIZTsT57a2Er7JHX0iqT+UTd7QKRbCxsoAK6kIOMiOhsVzjjJw5oD3
PZ/aesK4QT4iD2AZa7iDCxL95407QcqeMuQR/viQb6fDJISdH2pP+5o3ff9gxHJJ
qPjn+1t6ApyQrEHkTut5Cjf+PddJjC3tc8qg4QfaxtlLGtykBkRYeojigL/BPjWl
Y5jQ6yQ4kpMuXyiCgGeHWqbl8ROvZztupq6FrFHT3x+9BWwwZIheegz+06W3/p1m
uf+ynONWHxrvsAVHCVSQ3dS/Ll12ekPJO98T+4o1ZDpawKp2FkDs5pLsnZ8ddAZq
NNd2vMSfqMyfEkc80plOPWb2YakS5L/J7hsdoEKEM9F9hKmasLx4WPk9GHlNb9SU
xXt+k1JvTZI88wBYl8vqu4+9fRPSEeCjRO5XofJhl65QI3B12HG9/VoaBXPetlic
IBYyhFpigvG3sIe9AzhytDeudoiUxENK0LFVWqPN+hUHAo0Xsk/0c2BNEb6JVcAN
s22xR9dWHULttqIa1+KpebP+hUhclp2StBFJgA2kmNV3M+LKkhMV7KpAPO1lGmhO
lEz2wuJfyY339FeTHWE410Ow/tMYsHXRHYIEpJd0/rDdIRwpNwzBWWA8+eU+Ze/Y
hgHF8IEAI1cXM6q7h5SviENDYCnCyR3fbjoN6jZdclLIXkGYZNKuWX3IADZ86mHP
wFkjBjPh267BzL0uquPUWv7C6NzJu03EzbLN1DJCOD/vupfHm0f5QB8WvG6/ynjc
1C9SL7SIVk8qjGsMzj4l297rG6BUrLsdoi55qRl14whdEry4E4+xAfunhDAfGx+d
3KGI5biQ3QXwlhjmaKlUbIxW26mPnsc25TTpmNgbt2igz1lQlRYCsaQAvuT4+ADE
VOmyW/Cy8Jdzg/iB8zjJRly4iXgywEGtfxTIIV1wpPu2HY8XjZn3GL9p1K5bxTS9
ut13yS9PkrVoKrxjfiaA06D5YYmkaLZ1tPJu6rTrmme9HyJ1GKCeDCVMdyT2W8KZ
jCH3jE/UvyqjV0u4lIQh/ljmsEaf11Ow8WUdKED0NGOblQygB0B2DbqDtBDNnxrQ
285abVVugORKktUE2Z7QV1V58ZpV2FKdFtsRdbvXtudiF3KAdJz7PQKJNgNxSHJb
pg4Bi2NXlO7jINPArsfop6ttUvQpqeQ0xmgSvJcpGQn7OR4raJ63eS6mdo8RFXD5
UxO+Qk4HFCrwERIlC2542tt01SAVtb92gNm5DZiuOQZkGAnguf+NQwnLddizncJ0
GApcDFW3yagvEf4HqS/QQGGop9HQ+5OBxuBhEF+UnE9d8jQhW+bjxymGjbPJucU8
CtxOf1ZB7JENSOUJbbDWRsekykiGp75ua9jHGyQGAuLKIWKjBESffM3buCIE82c1
69TjXXKt0pbAYnFNJkKFgRDGjUCbW1xgdzECwoRgMJAPplklrMN1Ky8iZKaqia+w
N1NWFdfFDV9wu7ia6pYTijkFrXOG0B1tOYEPyLLm+DJXEnakYyyviq3TAXaTEvMc
faCHkt2bJugOVqOiYE5427bumSfLz8TeoA+FpP/kBr7UytNE1zOiFMf655xXHkGr
P48pXXGAOUkAnsS8/p60uoGJXNl/aG7SR6tcJgSdoHcixgiwU32JItwJm77HX9Fy
AwWRzEaP8I6kQMPvphc9jGmv3K68D42A80sj3DP1C8ukOHiiVCRdFkMdb4EqjiJu
52+aJqZAeJKGTZWpuO6AeFKv6KjKXL9x+KryKB0SkX+yRkaHb2hAbvui9pXCKoym
vVkiAmCA/M22h18BZlgUHk3AX9SQ6B5tHsSbr9vcmvX9PAY2f0iHlqsLIMFa8gLm
lgJL2D1bba08cZYAn+zvgFxbwS16GdyliJFBUD9XQc+3EiasxZsNZNeK0bK34MP8
MzXW7bO/T/58PIhRP6B/tlTAztps/765yn7hCu+Gs4zBiCJmav9/yIy6NC/cYoHt
5Mdeb2ajV0rV6uQCxx2eCBUEYzkMi/yp/FQBEQgaI+2hITbpcVTEePkySvWS7Ja6
GjHu1oHwFriupSt9nNdl/7v5xiYkgPfWGTxRn7i+xG4V/3rVs1ISlX/xZScGHB90
q9Y7Z36ZRxXdQcYGAhnfJD4cPAwwoZuZWR/3adYAAOOxynEnc28+Vd6NoOND+U38
1iq4Hh/85bpgA4pL0LVz1Icaakff1Nu2fpcGsLJCoonyqJPuQqhscXEbi2dgxa1G
ilLc/bSLrKRg0UYMyaq5vmnk7sBZ1ZZg/AU1sR8HtvOPege7FnY5h++nDGjP99Oo
jz4WpdOkU9fUA/4TqRbln4j6LYFeFaAaqbvrFXHHqKIrHYG/cSWkvlY1kwTbno//
YFisTpCwBqSIydYpjXFH5bwNDHNK+sU/MkM1ih8NSghEvRICT8F5b1WRMjvjcAix
EuUl2Vgzm5WTTFef61ii3QONS/CQq9PYT1yxOdEeQdy22KkY0qWa6OwcDjp4v0JP
nRWzy+1q6suJcXNdv/pR4ARehAuQq+KXWE8ggQt6iXOUwZdFxEHVw4r+58sOuBgl
/BkM40Ja8CS3rVhIFhhAOBOanxlm5D1B4RDbG2zY2OeDW3Xarf4nZ7RvrbGxElQl
GTVPHb77IvTyj2eZOVY2KGH72FuveRXu8KTwBI55hYyQa6Y5B6fFBqiafLqNiwws
rx/bw6iAZmbluDEz1ZfmLqv/jQDpOOdv6nVfZSZfRe7bx1QA98jVh3CvLPNKmj7X
U1vl0+lYBl1epdzs9jZUVcZdoiI1D8bGc3zHQ7s5dfQdmWA8gimHu5MBsZRhg7MA
9cy8DeNJB8kJNFSndszdOCOUZTw5vsE6x3498Keh7ANDF9YeFvVytEsF1oHG+ZKs
aYdDiJiJyGHsmo0Z+uopUk3Okk3Gds+a6UrpvKlKLknaKdWFBierKjMG7nvzQ61h
hYTe6y5kSb122FElcpUryIO8x6A5jiwgo7E+LDdUhjfGAfURPtDKLIEMldacWT1E
EgWcmm0eP232Ze08ybht0lTE/WifmBEkwq9LsgnwgW5PtMITQAHAjhyePJgOjrEN
71JTwK57SJinl28JwH9zIEULX+07YmNem61scVl3IPj50pNwpODeKpp10zLer8hA
uK3IGgOpsW7lMsYZjJHaCqaWM8dYGtGR/CueH2hc/RY=
`protect END_PROTECTED
