`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lIVlkK5DlPanEbE5EujKRuqpwMDZrXJLPXU+ZAWOxXdoux65jK82oqN04DhzSiFf
33yFFzfGRiJU6qcHFDsD9t6bk6ne3UPzO/BK7E8lVs1+BIrZzB+yPNlfCdbclTkS
E03CoAzRh86JWRQNAsfhXoznJipiIZfkDkkB2hk+N3o+qWG/XtG9VcEziTdv14Pb
RVtL4O3jnDMRUs9PyMMt0rb2Z6dSDLkK7eDy+S042KPaHxn56Ty+xdmBEJZ0zxzf
PsBqRW+BSy+vpNuxsj1MYsij7hsGOoZypSrCpHS7u+MRmsppWAm8jZH9M5rDFTxG
XSQN9NW4ulib7L64kQa5IcKMSk5k1dmQ4wxFsanadXSiSqlZjf2pKkHvcNJxiXUg
sD1Mdv2r0aKbOfeYUcCBHybPfVFUZx9vwkLWbnl+t2U=
`protect END_PROTECTED
