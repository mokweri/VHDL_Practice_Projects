`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ON/cax3zR4RHa1BtB5AvHn9/RXpUG8XxszV8BVl7luPJUnQs4LxF+oVsKQZSuwB1
AhmKNyXW9mK8Mj2u7YEIqYNFhECADObBp1nxJikxTuB4tWfGB9Sf0cCHS+5j37tP
o0jc8vz5X5xynwtlP/HnmjsyDM0CV8JfWnyMn5o+Rdm3UBdYMOVny2p8UMr3Qo2t
OHiX22UG3N2FnJrgm4m9hdUS4zTP2PcA+Duejoy+qeD/ftQI0DM2SXGDtuB5nT8v
6KjbfKI5cAqx/Ma7l4vJrzxsowzU/I3ZtFW6mCv/2DylwbovUesCYjjbZxoO74qM
7R3+hQ2h9k29EmgrcO1E58zLqrVVOAzRlj7k1ULjxngt+gE3/JabdGg1JySuzbfZ
fsT37I+5Yng4Ivf1bEx37pmldLL3ScAkaq2U/ykXh0/MvIfEXiHOikGdCUh9x/q6
w88QtWA1beYfx5ZWX1iyBMle1Tq9Dqjyf9Qp+QGQqj+NQfUtxI+A4ysc3BloJ2nE
JrAXSZ7WU3UqHNaLCV6lHtI/IEjwhgLycE+ak2Bnb/iEI7hI/4wleQGOGWArQj21
56s9IQ4CInaErO6biYGnHE+/gUtULjvAad07buVyztBw1MJaSaRdwNLjwRZokqbt
tymEM//xh+RNonzv9AP0fWsfS4N7YeTopHEE8SxtOwSzo9zq3FLV140K+xkeOBfq
SSuHPmwmpVuhFm90rKuxQrVh/obAenvooZQH8vTL1f4CdydPktymsLL7061fgZbE
JZi1V5dyfMrX2pCqujAk1V7jDuJ/EC4b8P1/rHgqoUMOqwc+TCkMzgmw83C5MgIU
PZkGkevvS68urngMkoUx/91pOgnRBwq8WVRjqNxFZJLtYgx0hZ/uqtPi6E8Ro3K1
OFAXrMhvjmRrM9qHabJzPBwhDgq0D/MVxm6XsZK+gxG0rLYalk948hQ8Yi8uOquR
DyOkfnx6ClyU17j2DJxD+jxFdccxnCwgqH6vfphyRusuvoZfu3pfwVuI/Lkhmewx
gXloNEbrckq9+Q8PA9RFBvArWWLh5iSwQqhVFI92tob3YHapUEsDeM0hXGNuoJye
vp9tvfNa7lZ4y+QbHeJH46Nld9LDiMMHnW9X/LWoXOzQVsXVOtj+IinIuWuXyFhK
mx71ie2UL3ni7L6ZW+b7s3ciNb/jHGLQId3WKQj3AP+SK8xvxo8MhDaXzcxZ1Jgd
Rc4usUfMylMn08TEzAKHNWswmfro5EuZhReobQr32z6GsXDXI33Qmf85vKE+81BL
g3vZ8sR9RrasIvMSAIyg2WjojUbNE9elzn4JSrxwwFfnV43zjupDCYrmu7/ws6Su
b+ACmYkzkLEaHAxfTEdBYBULEI8kcXP/4gOJG01dX+Lzkt8LmvnIa3RvBzmm+FPq
FuNUjHP0r/wjvpE2YBka1SxAo0fz1rkRmNfSadJCksUR0ugDcpRN9LckvSJPWL3G
eGaRtg3gmb400311s3xFLmf2RDfPqVDHlUyzKnFlw/t2d9q4/AlDU2Wni53bSAoK
uJ57j+ALU03zjRzXWmCWB6Plvw8rc/I1fCU+yQYauyt6b7/hshYkWm8ZKUKeLqiv
XCi/DdaHFeXws4kMdxXF4ofyozl/EQdSh41RVkS4T+31qyUZcxdFktdrEO4+qrFB
rHmFrp6ykktFWEHywoU0IsQlb46YIwo73iEGeFbYtFp31y7M77CQDgmH70bU3RkC
WBlcfdnpnUzFBzkEStq31G5LenAT1GroI/yPtm8i0LZvUAqur1DgYuutBT2Yoqap
UFE9TJ7iRl/DXOiyYGQ8ype3+M0poW0oEmnubuMnPKNEz0kpzzgHKsLGEhHW4pJJ
A0I24bZI0hxEEoItcBsEHTIr4WKNLoOtGbGfjcKCOmNo8G/z4t0WKX7AL1qaaS3l
hxn9IGXow+ERXdhmXpw0lkff5GQiD7A+ggPObpkEtomfHBBFM/5ATbYlv/wcc28n
WXdhYYDKToD6lEIZiumuNJEHq/xZpgN6N+VJ3+piq3U8nyCKgXP1oCzZ2HoyQ/MA
NIQzG6GuhAYKDW8LXfbHZreTB4mK5wmwdyUxcGr7wgyUpJCtaAOgYDM01uy0zKrb
d1Zs3E8E4S54OsKiRms0Fpi43Lxzoi4tG0LmbFanceUvmyaHVO9mXksNizbuCVSV
9d6CMFyjx+ocPQiH1/NQkaTuH6yH6H95L6KfAa0iqi21OB9G8mp9rnD/MyvIHt1v
Cyt43u4HrbPwWk9/4yH5ebstyzoN9dJP4f9WKcdb65rkUqUxUinG/PEUnVD4fMHU
4QPI+42vIM9AzTWsLE3GTPI3QHJGAiEfUq1/HrEbxdXfa/RERoQtQ3C6AzD4npYW
Pk2c1nd7BUVSx4qbeD/DaZBtOoWAt6nAS4dMTe8eF8AKgmC0wq3W5Xy0uyEIXEnA
x/iq2juT35d1kDgACH0D+gpmOrn8YycAeY4g0WTsYP4ZD2ojPjyQ8iih8Ax7VvT/
BLhLm3IyYBBFsAHfpu9vG2Kal1qL1LTpvRpZoctD2eLBGJwG5/oXMMIOBABq/EjH
YVeSB4fjtPFz7kOfZJ+7JOpSxZnQ0B+LRhAN39W9uzMKlXuLu2VODWPkD3cJr+Th
EeAJLUfnEMyj2oYIDhSQDf1uYTbkdMddoGAzt6FdisS8JxkGPJ3DHUotJnTJI4oS
PuEmcagtPBKuGZgvUQRbXE2bZwNoYIzohASOCAcavKEHar/aJPQMcaC4wPwlQXQO
9i6ABhaQKCJsjkLEMvAE8BGrUImiyB4uSComciQnvdQCAQjLZx/IDsACq+Dkqntp
6sAsngYBxLjD4ixpYkOvnOLNtktpbOLjmieHvgGaFSlK0+d4Ca8YKuQZ0Hw1SXMo
9Ekp8rXN9sIidvywK1VtUb8/iktw85evzcD0l7LjfDFWjl858wZRWerxGUUOJ9qI
lPDLyHV0A+wu5V35U5mt2dV9tVFgv0Y/8YnyN+XMRqIH9lHBcDoJz4l2UZzRsKWc
lVurKM3oZZQPJbGIoyXF+1nVQYUbw9h2bQ6HC/v7raEyUYkpvdWPjwyMfRcjk+LL
puEYBrFdtGpvkzgOZIORiX25fUQ9kFQC6DEVGBwoAuLNLWmjDhXY2HAfO20EdOEV
qPfwPay8f52O6keUDFsJzcuhF0Ist3nE3SFRqZkoyajdnyYzNP4sYD3JZbGE29Mi
uJf0Q90XwVa8bA9yKqjM2WuZMrxBv0e1jupIbJ+AEXeKtOH/oHSVvdW1KpFTimjp
DhD1b8OkO5GmnH6/t52rq1eOai1VGp86Y12MBTIpYBsfDI9kqh/6gf1vW/J4lj70
7WBWoEMbUKHKbhO6UjRSs70/+PfpJVBCV78Lcwi4uEoH8p4rvUM1K1AeZRrJVLgz
XFXxZHAuVSyh6gXT5/GhXOBmIl0YIbRYQFFzGV8wdpbXWaUgDot7uVff2oDexEIN
0u4VHbV6L5TZxBcfA2Ti7neBETyjmN/bqGODuq0JTlefuaY5QdU8ETfX8fyG0lR/
GWCB2eOOn5+vKkN5yCe60IODpS9EKLgb15e4wmjFxkOcZxe+suB/DWskZ8h7k1/d
H2SAp8brkSWNaq0X7HGFa3+6Y80+rnheA0QAuLHhkqnhg6AOrxH44VKlgUYuU3cK
H0gP2e0Y6MkKmFfuJAZQZN2168n+Q/4s9Fx5858NESlRKpcn4a2saS6m6po2+bUb
cmwgbV6rDvilN9Per18qvQ==
`protect END_PROTECTED
