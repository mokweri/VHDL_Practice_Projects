`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OaXklq2x1II7fVF1aUJGew1J7bwe2aIE682QH36bg7hV0tr9coUVGNAGcqXFGmLp
YvpiExLxKSZuQD7sOkMSmj4750y5iWw5vWDBSLFIeDtpCG/S0tVhiLOUqOOUzJ6A
aPoIcs5DEpTlpiewrQZXqDHa3BFtHD2cRUyPZxmnv/W1Gv9+unre4P77ASTQmsPl
gHfHo0481LboCqn07jiSVbBjYY1exsOoetgsHv2P9YZgqP1QtWBmTyn/Jj947MVd
SVuUZDKeulaILLc7qx4RvZM8JEwLIIW6IdVtuCMr1tUGyGn9WMvD9PCHgdfpUkjj
1utLcESc2QN7rBjHTCUycWTNENRcijvZvlUjkvgKB8jI4a5RXamWxaQaylJ9/Mcv
YlXmWbqZe0KAwhBIGjP5QUuSBP2JqJ8UesSoF7zKAIf1r7dum0VilJlRplKnSHh2
J33QW+C2OiFBo9atCOuPTLhTeMIPatcCjnnamle00n4L4l5eeygCs54SXhUL3lUw
awGFt3Mx9BbJwVjHMtz9F5gokYDl5OTx887x+oSwkd2Nc6gf0+ypE2vJs9MYwMIv
xUeY28blNMyubW+2KUrXxJ+q2XzWzKsu2aJau8fIs6pu5itU0B+UuXguxjCJ/KLw
Kw0BzDHbfSO42Kxv7oAG5WLCi7RjUuOuk00EXvzGe2B8MY3wTdLg9IBPXFIcJB0e
Ixw6vVj3/ix9Kc9kQ0ODT165kTKYLzuejHVfqdHjjxhkZc2cQeMHnJFmHVWZZgb+
98FYUiBx7k1EWjS19wOmo961D4nxoa+mgkoTVsqWGo9MyKEnN0bZ53cnh+rqQvFx
EFoE6Tr6JJSHPlAEbDUjrK3MRfbhwTVIOAhyKDhNJYVRIZfFaorJwMzncXR2wAF+
A9Ef8ydbQhY6jsgZDzk1DWOyGuHaX1HzfBeav0OXiISadzNAlcEqEVINRipnLB+1
1/q1o7ISfZlYjm9NgOUttdO7Hwy5vsJxa7OWSAe0Q4fDx73C1kekh4AsjMK60jc5
Vs52yuI563nCADd9w3472ifdRPyt7R0TZsLVYabE0iLTpDnNSx2yORa/GvtxKVs0
Lcq59eU7QUEOQAa3AhzLnLwRnBcbaTijEZm0B1+kK2sBQLQ+xuSk++ybVaXF6ZPo
F1wIcAu8FBXFKZaY907o9kNNnF4V+tLffXnnduoOBda5j54B6cZgbsWANFhV5Mi/
FR1SAXYfjHvhXuX2qV6ob8hZnIUpPkbdQquQv5Km4BCeekvgTNF9GGbrOS5KqXvH
v9nVXdDguanF/wTwL0PORU9EEEec9O4HIpiKLyY5nQLS5b/hFpMw4FIBHXHi8jJl
jet5agNx0Mhcki+Q5Gtk2d/B4asa39j8pzjLjWFO6FASP+0twewd97cDGpEq1mF5
oSOp1ex+apU53TiovkMD78qQBsvT9sfWM3euwQ2H5fz6URFLIl0kKfnmndj6J2lF
jcWXW1Docm7BSfCRtJUCZMtljLaye9QuFnilaULlz9k5m6TGmfcvoNd2fGk+AvNr
YkbYTSTqqNqYmgFOWrerYy4bWAfMMk4iA7SfWupm3FA3j7ifKuuBuKCNcV6BSwws
6JIl1mjeJluK03uyfm8FDLPqmgLGU/JKxAE57FjdJweveOFY+Opgxao+UTD6IV2K
tCw/6+6pjU2BCNjR/Ffu0PXHb32pBoxD39Y9AUqM2lfWVUmAsU7Ts5K+6ygj6nfJ
96oPpPmq+LqmDCLkC9c1OZIVTSVHIhnMqB6sKQX7hytg8ql9fU4iSa6fqWwVV006
s1MlgZTTWB2ZJdLBkXjfP7+angqosyvyG/8LCVrgt3M2rv30WWWZNBxlIs+KEc7w
v7VpoTtezhlxlI3QXW0+6Cb990/0wQDmldYfXhmXl5xK9d/GOpgzJMq4lrqfXj02
RYmQvJjvs8YCoyH+mu+7N6YsRDZvEF7zykb9cPtqldusYWNUAltqMwdya5GELLGi
br9cjP9ONWfc6MYqJzdOMbfAl56jhmvHXDPDr/wTWzzdM+k0c90kPptOK6cYqX/r
GANj660k5Yb4Ks9X3V9NiSd5vha1JlLuH58M6iU3BxSJCARE1Dj6qRZQbQMm7Wr/
2777iPUU/Vo9EEJnv5CRkufGl0NCiVcm/wug+E9X1HJF67GsqG2eV01LzEohOrUC
DcBwUQ6aSiXaYR/EAc1KsbtvIRTOB9FfgIiDOyLXI7Il4xDPZ1nK83fcicfxH4Jp
GQ//qHhy1IADMu9HWQ0wMn0EHbEcq0CZbrJG+CvljZYYdrOh3D8RdHwufyGcWA0u
5izDIKLqbM5jefDrsCebeZKUyFcu5kB8DHeS6qNxaBi5IJXaUTiN7mxv9n3NEvIf
HjeT916uD1FeUaqoltV5EIl7HFFCTV/7I3yDwJw/tu+gJKlurzvS8ODUBLszwJht
TPD6eIg+rdOCAIPedVbCfYc0flZPVyew9OJAbo3PKyOUpK2W5zWGzAQIXBtnKo19
rWYDjq4RRbrlTTh1NZ70OBq+7akRIk+OmW3GvV831qt3uwC3uwrumHCZ6/sXFHvg
SYjpgoj1VdvZ+3ln21ZWh2iJIzaxPTG3IcsntBb76XPnNuy3kaAao38AF5f0FTcc
XJ+iUKZWILIW4f0dqFhvARAudg/RujLsbMhl2/4HBJd3cTT5sktMn5zZaFfWC2CO
0CuQw6tS4UQQr+dRDyd8YkfqiDrN+6U64dAj4mkTkzg7oGgmHuYFzJVeMGWfubF/
lhmF6lvhm6jZftdwitumSdtNKvSiypOHX5NdJHcKX/tPW7ZDNXMyjYOL0pQud4Ru
gNP3ZS1U2K6epKJOXxLRIX6/1ZmW51rgyh7X3Uq1DevvrxFZrCcZ9wNoeMJ0Xcvj
b69xOTvCFrKVMcRpcmgigFrBVuSdiZEoWOMpMk7misAWZnHQGwSwioU1nmFa4VxZ
w8El+oaA8ueDpal0wh9Fmi3nhaBulCxTuRfeK9tqKpIg7ezdqvrSkXvwXAVHT37l
C8lv0S5AreHif4CEX+Yg4ekgmHgCUxURzfnnNfDNv15miF88YPDxavnQCaf5Kf0Y
H/AjYFUeFrz97ZFkU76+4wmXANCyAMWN0ZgwtQ2XfXBaUSDAASRYFvJfhQgJg5te
3KkZ937pjDLDPwaU8iZIW7juBYR55KKEzgzbk2dXnYPCjFSuFSo88B2HOqgFaaCQ
VOUA7Ziu666yKs0AWnsm09U9IWWuAnjBlDkWvYAKAU6kmcFz0xDwSWRDC7xMRa6u
4g9xDgr9RhOX/2Mx4mjNNZs0LlBjE6MrhpKXP/GIvEscmo3k+l7BX//Rme2Qbml7
JYCM3bO2WplD5UHjoPo3UbXmR5PFcLtko+I7YMQopi3hi5PpHUFQzRDQdrK/lJow
gn0xPQfBWipUJVz7lw1R+BORmDI1hwMPb4nYBZsw85St2vbp9TflWut87lv6+9zR
FjipPL723zQHxJEN5/ICaOi+iLq12aFi3T9FBS7V+EaVZMcPZAyVu4al+oacnGXk
jMpr4Vw5pdLdtb9F9o0UmLbcgU7+Oktk0DmvHqaAwCzs17mlyzjZVc3BlXx54Qy8
iH/gBBo+RvlyUuj4VBEToeasrcfGZniCxFCyw6k+5uRwZ3F/+TsVKGKjPcDAPmeq
Wn7KlHe80kSTuuCqw8oXBNz7BlKDT8EF8tH2rC1tIECons6GjW7tdJbMxPaM2cH2
wRLfDOxTc8KyEPigHIwAncfB0fSgKKVVUrncbCIevJlKtImb1wOOXCtO65oT4CR2
rH3amuqn4JE5MIDAk5JMuNMQZ/FkIgXtIZaKAJREmBBBW/rYUwTtU0wHfnEgdWX+
ICB+maRSfhQhVvDDvJvGpPi/X3l7H0ALigxcv8pgry68HUscsMciOaBiIUfs1/Pu
1gZgH67k3M7dqytMLtCQXNthEGf2yh4I/15Kqs+zNASlDsUsoHcTQzdSJFKy+KM0
DQZXGfHBzbLdgCG8CETGOtiZL7O4lpZBJ7UhWGO774QTxSYFHk1bjSuGr9Xq6mMd
QBO6Jge+1QRd/QlrhzTfGUKaSyTgM5cI2VBHKpHZT26/imEt4N/Ul8cdjJ75b3LK
8pG1USIWGLwwGSxpAkS0WUVhX7bdwdKaiAYGaGsnIf81UqpQQBH56rqVTE7KnF6F
O4YiAYPTCrIa0+i+RP2iuC312GxBAr1V4ZW5rXCnlNW5R/7GjdjN4zh5ml+MWG5D
b9p1qyR0WlF/RJrkn2D5HnnhXRvBEK3/jtIbuljQ5GGPpbY3zdM4e0xYZJqNJ19g
jGPY9b6ueZ7QWeTMIOrbRaa88xU+miQK3nDAUP765y0V5zX75x8NfYY2hazCW4M/
nFP4PIG8PC03PQSfOnwJrpoc6nXmMqpP2Ics7sEotMDE23ywsOp+2XC4voaDW2+t
Fr+Cifh+WHvMLkgaDRW88ji03T7febwCVkCqoGwW3Zb2Qu9sIxY2ikHgqteUQ0Ia
lLHIKACRBZPV+jjC9ZGlJ2V3MvbJ7dqrqm/JD6cdprIDLAXQBq2LgY8PhuqzS9+v
32nTiG2pzIgRyXRSs5wcTv0oPDU2pSqQ3D5f1i4ZK1qcHYWVpkMuBAoGDCiBM7rP
e0VdoLzKjku8L9YTg3r/DNCM8Wg2Z+xXub//lK9fyH9KhbNo4Z13IjmJA+ThggOM
98PlFEWasxzvkJwtn8DAlqrr5BMTFh06v+Ca4burmaB58piX6d7qcC9Ex3xzE5lN
Wm3dsYZGnKcDFkXqX0Os3dlL4SCzb7wd9uYg8aU69uGrRAi2Ckpdp3Gvv8PBCspy
K4GsnQebNLdLBqdp4g1poi2gJwLzue1l9JfAHVR406gKy0/MTtWRRexf81nJJa1Y
iJl32AGqeTNJp85Lb97pfcDmnilL7FFZthCO3aMpqG3JnXqV9OKEAk9Zi84O/art
HK5S+FaMQOLc138Gz6UfDGB7va1XzehfvfTFVOwhlKTO2n06jEUCtHf0yRvSVB+9
JEhWELQoLrxYp3GvKAxhj2azbkAFQEcXEJ3VSVgY8hhMmFclrRb2KqV/ReTPEUQG
PiT7S0kCzxocZQBhuE5YQggTfZ05bKk/sg46nPK4kMvgkLdpmCdRWy7A0Q0FBa6F
2B668O09ZNVLWVs6kE7VgSFuCqgKNWqD6Tb8oiqdLnuHyWHlHyGrmpc6nricN2Z2
21HxSgdfOkdEEIEgYA7zwDsXzPbsOChBzrYXla7K8dbDp3lKDyX6hpSJdktb6pwR
ezxhUInZoE8CImYMRtHD7nu1krJTsV4KEnVTO7zCXetJ10dlFpcfuhW0OfqNLoCm
NYsjD+HYWQxBTWScjwEYdTHSqyTuujXpYQwf61hBQi4SPJsXc7LLV/UBgQhiCBl3
3nxLcs5hZwh3BZeafvN2BqhYbtrXZvSf9hK6/6Tm/YazZ9jIUgrNseeb4b24MUcD
PKSTRLUt31qxpI2Zer+nhHhsQ5Ho6bVIBWBEL1qU2ExgGbJX7wg2P1DY7yAhztxJ
LwD734sFKUGxKBbq2qb3gTQAk8FCILsqN0ExX553Ll1E3/s6ZaFb70eMSnYIrHtN
b1Jmxy+gBVJE+UPqGi+ybLdkYMr1c2eE9Ek9mkIzOyaBwE/ielwU+oAs4V1lliwy
BJ7TdZbUT2uUS6M6CzIQxCOJjxxtQLYjHgLFDkbiwxKVoU7fRWtiI+kenoUOEPOz
Roy2L/WffQ6RuuByVzZTg0sJAx2TVAmWFEePiukhnQ4sO+Do8jINgF72AOkmKoo/
M0zU8YHo2sLnAoEjzTzTZpfr66EfFyp5Zclt9ttqJFlH5s/WhSWy0X6uVrK3NPIY
M+gWVXQzK3VgorU/cRlquS/DMww7mQ22EYlt/hOx1o0/PE+aDJAv3McG0bq+qnKI
0dJv5gvv/Z3+B5mFeuczOPFpGeRPSzqcBHtQEJq6d4mAFj0Un3PE/UykQMQa0d/I
MEVZA+KckR8bZZ5LuTd27azwQZIe0jC12+9zex4xYLaVqOgnMyPiZryCajd3E120
YTKX8ZLg9hch9zWaS+4pudlaUSLEoL+JREcHnJd3af3kPqUhdbAc58yFpQW7Ncyu
2kN33ZsVD8mThFZWmA//9MEJrQ4TtSnzUxkqpvZk1ommSPlwtNcj+0P2jEqfSANB
9snLer9UtiEguXEpa7KviqB4Dgwbv/cBQbWPRwsqZKDYku70XmlKt1/lzNvuEa7g
zgfHOsljzDkUnKah9xijWTMAfkQrl6PwNKolFIEKCc00192ZASBSqcf4frwjWA6Z
GuDXTeWLBlkGW9/jeAquMyxLI2G3DHxPpVdBEWb7Abt319tc8orKHDr9uFrKahZh
y5i1LQocYaTSuh+MfXum2f/Cvn+OUHcU79sYxfgoJ4NjFuYJfKlYBSfdXMf+eRWy
VYnsWJmU/CNti545AjxlGmL2gc67uJfsU321+mrcKcQOs+TDIiFAgH3XYfH+TOrF
gxrBz88jNlI6NvGEqnqc6DBan4FQ/Y1puTAD4Jum3fhBuZ+WP/JBcSwSXPiubzU8
C5lWbEA81FtdJebrWHgjz1fcThH8xP47DfC65W4EfUmTA+Tk9//KxFNzJBPcPD1i
NDolsdPOaZTNsTXp9VudVqJW8tZ5s11GUBySitBzta0gUtdCCcf/THRWYofKDuHE
AnG1jBJqy20Yeb1Wtpt0qpUSCvMTJki5Xi9ari8EwgRXNHMvceSwRgo+cH3sqkL6
WTr6vHTdPsKpy53jofthG3g+bJW2zRJD+vfe8xbiOvh1SfPtHSOnenJumnZKZwM/
tX/Nl1ZqaFGrtfnFRAsOFjzDGMqB2TYxIX9DdKNOUdzuTP6u/FGA4TvJWI5te2T0
2buRNs4PyHHbgz9iUcuF+BA9675nVjua96JDHdfHwUJ5nG36/pIV/lxcS26nM8of
s7vj5EhsJsA97/RR0CEMmqar59DHyrhySl+U7kdlUNJerY5DpAXC9RmH2VeytMow
ocGBN4gYdQLWnCaRBhrewvzgoIoPH+D1NC8YhZ0ZMeKjo8UzQyaYSNor2MXhT4+H
7AsMzDjJhZj84jQEGgIALCoGDqDzOLeTnFwNMjTLusbZyY/sHOnP6MKNMN9ArHJM
B/Y7Aa1o38KGrcRapYlu9kD91oU/l6BAxRgCyKajgxHYhmyEeQ1Fbc9aTgXSGcLW
l2e71r/YVDaQ2sC0gFY5QBsin3pNLmD24K4nLSfUH44dvyy7Uymipk4YHzLFeVWv
hzZE0oTo7/6zBy5C1UeG8AmhE+7kyoX+4cC1YXrSIUgReZMdmXzLYiVu8pO1egO2
+DwAtDSXHHE2uFYp4JxihRchjvGbxkgffNZp9vey/0vzz9itN0rlnoFNAtkBNyko
rNORE1FebUhmtwZCik0brKunOdC0xD4NaB659UEx0pDdgHZDM7kZrCGR1qbEQLtb
0fJJqoJpML7xqRPI6Hfl4ojdi9QU9aONIISIuNPbQIS2i8kZiG0lLXmZPrw9hG3G
AeitB+0xAmoEETYw/8ymca5q6O1N1TvdDLglHbWKObG83p91wW+fFSN50cG35nQX
HcqK9lEoibLvqOz2l+sTgw0R3RFTkUS4GXerT8qgdapUikqL+zVvhSMyq8a2TCoT
YGmUqtttytko35N2Ov1jwziioqgfOYxI4Yhegr810kMp0I32dZdpf7nRiRY3tUF6
BzpymXqML1o6tOXczDkkTo69eBUkGe5N08FXTBwOrnETC/77mcaXti/nPlatE2f4
xuTI3EPxa6N2LdlHtG6zpDv7QF+FCuenA7oRtG+K6XvFGNdjR5AZbBaJwLqlGRaY
6dFeBrppoB+yg3lZ6VGbUhIPYrAP7+iAKc3FqMeWe52nv4XgNDRrQhXGlGg8Zw4u
rbUfYoGafujgCyCJ/96thHC5XKXARpvtmfoeDIhSO657c0JC8/ZJ5e1N/icfNP+U
N9EilBpqJrHdYijiYPYdKg1O0K1WgUQhZkYQlncGpN8LLZ6hXzQm/lsAdeJ9a8NS
zNJXFJ/vVx8AGFVJdVNdgFoO9Jt/8v3G3Imdc2hy0YI=
`protect END_PROTECTED
