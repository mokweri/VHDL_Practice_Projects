`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iGc4zwimXbRdhdV+Y+QHS5YU5gVY8LSzVR/HZaqzSKqxAaKXzidSpxUIV0u8lJNI
jgnfxNv0QvxEp14YYUzfPkoL3eAPaXQops3hGZwfo0G4azTS2C5o1WopanIRgOiq
1RSfHhcqUXsBPLSVpaLUOvc5d0K/hmVtmv7JUw1GAfVmQH3QgYvAYZqBaO0+ny65
vvPxifvPmAs8XN5i0WUAWmVrXFHp4G0owqzeyAgE3slX3qLt633yzQwVyfb+k8oN
iqpQncgFFObzT615LtHkxr2idhLFHPdF0EEMLm+Q03GPF1aK0W7h6Ilcnrg5QnT+
0iJmW+nuuDogdwSE4952its4Bxr0cdM9Qt/NEbhoOmkWJWeVGt/9ovObCm1Pz2TE
qcSOcbZ5dasoXWWGmvVEdJuDnh3aJoezkTATw1f1EFryIpBQXMl+8DJgjQVdwo6L
LGOA/VtRj/V5lHSAxQGeW7qIRJqwZHcMLBSwOPDKzJI=
`protect END_PROTECTED
