`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4va7c/s6bWq3q+XmEXqpKbESJDre85qCMSIzmDK7nXcqO8+B5aaLM/j9Lh3S3rbz
xkM2901dvNX4JocCdOtNayA0l3DN/JhaCQPttx5zPKEnyhn18lmbm8WFVRJnRhrJ
6RlUNwH12wKYCrqZvcbpOwbzejMGp+9ki2211NlUOhSXjwL+FDI5D0t5tjXvlxrG
IYMIVWZtdqUhb/nhefgRUefp15/A6W3Hbnzkbmuxs4VztlgYJDDtGJOxTJyyuJcB
j3BY1Z99rIORKHPk0vQnn3QmslqFi8WQ7aWHR0I9Zvx7NMXK+2rC1zIvpPascMT7
zOrkZWN3YaIDN/zEBz1E28grqAKAbu8G7liCJn9YhNFQDcmOnFhczeWjdK7yibq4
+OItOuiXzcYMEIofbAxOZhWlf839XuSyagKcR7qqgOEqk0yURVi1HaZ/1Wc+kyzO
ZCUGF81hJx9w4v48Kx3bFjUcwI9vlsL/PA6PukZXCCNZlohy36Zi/OzS3Qvspyv2
cp0p4CRyU3P/BgLtgaHQE7tMXcxsJA+YtxOYnVUp5Ob+3/KfR2J1GOZA2e+EwUuv
jyKEeykVGxMnSSDZ40nmIiVGWGownL5fQ8S2frKzYKkCybTJbgticPHqj71bpTp5
zVRbGj+EtCvSToMvGlYfZZequ10PyrIOUnHKGd90Cxo744GNw7j0cLC3MGCHwp7m
TQ5FLIDH+O+N7Coh1fgI9ZFC4rPyekkmFf5CfR1H/XtA7tq1JU5mLt4RPkn49B0N
91R0zUMHobYE2Qa6FrqRvbPX3nLPaUnJSAqcw5qW1C8WXsetqTIBX+/L4XsBbf/O
QPcDeCyP7siIvL4cvnvmq0as+rNwUwO8542zdzW8185CtLE3gGFJvmV7bk5YTHht
7mC/OsQMrl7KdNFVfn0godFCTUC037HgEFv3dQIglH2Xg/TTElt7zlgjXaux3tk2
Pl6i/dEptkdZzYubYvOq6PldhIXhVWVq9e/QwlEAWPbVES1S3u4BtAdaqgJX7VJ9
K6wGq7XjKNWCyOb7AMq+0dbiDSL66NjK+3vXrGuXBmdE+jXAsQbIYqRmEOKMUEpl
URHF5jyKkYwCHjGwl2b426zMCX4Crw2RBQR2rDXIQQc9tKXoAGLzsbiL5WYoB5aM
tk9yQZ4eUBB5h4QCO4SThj53LZmR+UlCaRntfIJr4KDHWbsQa8bN/3S/+CK+/rt5
tuS46jYl1G7hpmO2w7U/SOT1FKIfEszZ5Jl+cExGXku5agQ4UjXI8KU8AXSi1XyK
jOaoI5GM+0hY6EMTqBW/XrpNu0GxahFNc2Q6hKX1/pYrbUrr/b0Z0HJNF60uMePy
Prvh6GzQZYnmY8Pdde7GIdrmFCYw8R+ZPkZp2esrdxE8acIXU2+QOeCMPwQ6ElGD
A0/iHURsrLezNCKsTMNbmfxLWptCPndfgvF4NpWbOPzABSwzde9BDyyEHcdk46/z
9jxTa9/Pop4IzvPFriP1RU6Qdmme5cv3UhgJir+u8YQMz8zUa8+3Im5/706ycnWT
ql7MIaKm01lMiLEs9M5WNh2BD96B/0UIDHIJqlL/oZ0fFKYySYs14dQtIeMVPTp6
rMmLqMhafxC84kJqOeeZGHVnBD38qwHoxP5Kr/RxqOUZeSjbE6U6ToBweoYEsuYR
J3hvv2u7K2vvjnQZPfaLXk8z8xfRkqaQ0xt7WEmjyG8hug/tRVX04zvnsofMSrkL
W3WG7N6QqrJ1tfar5NUNyQtHpeo3uTeABMOr8UyXj8jC/CJerNUydwHh32qDTAyf
ZIT7oeHRZCLMcTMLcPVIi/4AVj32ZGoEbeQRU7ej8f9DZNriR92Yoi99c3bAux2U
VxyMQiizlGj1eXVGYCvTw+W5ckEuRIwq1MWwNQt0Ps6Q1SdqbI2wGqy+4jdN5DtA
sPZx7QBAI9/vINnl/nDPMTiNrb6qCJHvVguVUBu4nwz/rwUpFHgCOpL+IgkBAFhz
`protect END_PROTECTED
