`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONk43kPJHmRStkGEsEncNLoEAYhj8ZR5QgmPofWWOqEMCE4TilHb0H3U1oSn+JlS
95Zu9r4Qk4v1NrAuRnVj4BdCnPn8hl/JjcTNXfPRHbZRm2PO5WspjybWhfbNK+fC
WlaWZtXPOmunXS+k+zYcp6pXVdsUyCrWZDjAKQqmVW7i4K7PGmPVI3iXmCgmRXNB
5wAC0rrkL2gM+rNRt6RU/4H2Sl507JLq29q0YuIXeqvqAWjbcafzynsQml/8ZMoU
Hklfph2UI3I3Vs/XB3xPFwHVFzgPNBXlBByZ/pv8h/yaSRTDmgNtXjdlNpNd4nHD
GNpSsxVpjm4L8Jf3v+gk2CE054z4CF/NL6ogGexah2Are7VD8n6XKwHyjTjRHoB6
N26T7u/lcer04PYsRoxNlVRrNDOZn5WbwmgmeCvPcTEGu30d4BVBLMkDGI2ws74Q
MgBIvmmy17X3+EN874uRqeVjjLaSit8tuXKyhTKSh48NZQSYkBR2cXyW53dqiJGE
S8NmQeP8X77ibx86u6CnOVVya5glapS433TwP+f/8L8yfIi6rV+mkFS3cB8613tw
SFA4cseliDHQ66iMNl/eEitymdTos/8lvINQtWyZxJVpbapCujWl8b/eU3OfF/5D
DEmgsiXsD2lPoYcyVElZAnmm6V+DVYKNCUjqWmC8uIPYo2EL8wwZ4Z5zfJ5pAnfj
LmALVPil7LKoZje9S2nQicC+MGvqN+rAsenTAAs6DVYJtSPPf0n/yZFTWT5pd2iQ
c0f4dgQTzfDOAj5pThn3mTydgxdz5IO7BbG46I0vPcpm+hi/qt6Nm7ZQfQ0qhHA9
KxgX+/bR5J8l9n4u4vllmfCmLleMD82H0F9WHfYmOuddD2O2TiiVkwH61l1AUSQO
1HmHApCn/HWJyNKwdHrFk7HcXvciUUndj/DWdfRUjvXJVWLoi0YsflvDk/tuqis8
F/glOXSN1DsMBP/WA7/0LieRNcgHOHwjISP9ZG6YC08W5N4Tsicx6xYT38oinc3S
WtAZAAqpeoGxL8jokFah6Hly5f3YQVXp2BvrydcgbXaRkcFO2CXmeO0uubhrE3LN
TtZiLUcwq5KAzJdIlwN0b9m+QdXhLcSzS7RDPvlxBOD1C4hMcksyQX9nfL78pEtq
GrYOmXEudVGwyzrsCAUfrQ==
`protect END_PROTECTED
