`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4WK6HdwfJGJRcvBL2fjZNDWpCtEFHfVq5EQKhtoyDTgS3weBQRQIRPUdWWECnfj
6ZrEK+ncxsufdIN81wynWeMyDaqd2EC3/YdKSvrIYMLgCNurN2Y1KbqzS0L0UO+f
cHIdUxu/LNunWc998WulgUz4EwC1VfqIWxqaVrihd8paqDdNcR5H0cGQR0N4boOS
eA/VpmdNJtecdqYeoBC147p7JreSE0Xn7mJSsCFf58UYYd6LqeWoyVCw8WacIg6n
V2VUM6oAlMYYMV1hoy23kP4pmKvhOPoiGMOQ3zxvaTsQ0HhyITLdEUD1u15BSL17
zgLUABQcbBOI7iFGU0w8iX0w4lEPPbTTUXywe3h8eTjOVndzn7BBpGUsrDFuNaVx
i3BcurreNt78RG7VCs2Qv1R38jrMmD5jNxcVhr+UXLcFYfYeMmiVn+vmh2ukxgdS
dJHidJGZCg5Q1Jq34aN0SIxvMdh+N+ZhfbGHvRlxyxpUyWkj7YniTfUEGjmnSaYK
Uq7UdC0K34iykoZIl4zhzz79QFvjtRpxyP/+nFDy5FzADgq04Pdk+0Rom99GcSag
vTD9i/xuP/c056w9OR29qnxuJt3Zi/E4A7GebzI4dEI2xig71oIIYnUOZzaEYva4
suogzuNOrbxnUNyM083rOfWtzxJPtAsJ68XwBHJ82o3cnTc5hd4828JvGx2V+7Q3
ByrayKEiH6xN8WpX+WwL5FV90r35S+CFn7ImvZboz/p6t/9RC45GHiAd0cA03Gin
KJgrR/zmltMRJdjDLkPEgpXWxn4q+++E4tWZl30Y3pwi70LmAUYUgl3SFinqHpDv
F3XhQb+DkBfy/Mbfd4PjEK6w8h4F6ZqOrKiJfnHSRAdNi/8JyD5Vdhog2KbltoWP
D2sHEqLHT8bnR0PNj/RRVbRG5t/Sm5h5khJQ01EL2yAfVGxGzl7oEq6akDty0gvp
z9SeLSNits44BjC5Sh0ib8nO5sxD4z7ZTF29CL7MQLroVubHIVyFJxl32SQTUbVI
f9itkVoC1jWZQdcZ87H9TEMjNijwtcmSdH2lBclQv5jELMP/oHIBlmZBKoeQdlTx
PpbB6nwEWua2VgBSdq3m+vr4xLLgyC2nBc68xi2COHi+bNPqsZ+OGpmSKqt687l/
mJnzOqjf2IYnoqgkfyFlQ2NPZ7fD5gqAvDJuQPDMVMXkZpanINCqel4vNtQjS9cX
1/JCho9ogG8IucdmqGeyvatuxnocXooT99uwKDKtZpyDCBKwznNMMWAr9QOSKpN2
ewCYf8UxuOp1Io8s+jMUf03tQBRLp9Qtz8Z1Od9IFZ+S+Ff5+QtYp4VEbSNkTNv8
wyT6YqP4MoH7JUJPRY5+jJBA+afyItLe/t3nUoJ2lX+QRQUi8MVE7996N6uCQlE3
Vg4tCUPPmqPpwmJq7iHVkbAaWLjxDm6UZ6k8wRFHc334rZnEepC39W6WTStovlNj
D2UnlEOkUC11nSwn1TYppiH73NebxTyNUFBxK501m5fnUc803jOLT5lBiKo9heOR
J8qFMvDn6hI38Bju75L0DOqZr/FY4InlIPz97QXflJVp1F+U6AzmJe0cS2l6uM3V
z0txQIMypU3KE8Y2fpQtrMRz5Kh0AplV2sxob3+J7//GqvckAtECH8X3pUDwk1Nz
k92Wm9F35V9cNb8wwdHSKlzsqCeR77nYv4A7SPKLf76uxMOxfahDeOoFTMvIJgbo
cSGpMhTS5ISw1AsNnwQX+fufh1h5YVGb+0T8gC4fdzMB923f8Z7auLKOqpyJC3/u
rkGHmZ1+2IdToi4aOsvk3Wqi6JzV7QY02YuIIPa3n3Bico27SkJxWHQh5htji+Qw
z36Iek7nJnllc97rpro4NnDwotcGoXyIfsgx9bgudoms4zLaA8TWMpegvfffZviG
KdPo6q4yjkbse1G9CJ8W9V3LJKRAF3rSW7GrvdWLy/hxNzccOQDFfXdrZKojt9cN
RhBzQ+FFXnUfv159031vyGjj3stkQJc/If8r74KSnBmtT78DLb+FEY3zJL9d3EnY
vAr7DWg0iezj+05X/h7WCRLIWSKLwLB6YWDROdHe3xh/AcB+rM3kKD5QY0DINkga
8vStSIP4bUI2n91xAZmHwyEQdDJhFsUJmM7k6xbFhOmU02WWdGTZ7wtedjseE6Bh
+jec0AfShFDCjid2/uRnmQkWLv6NPhD+oxo6zgNLqPo15hb8QYy0UT9VkLFmnIv7
vshUh8zBpB1Bwe8x+3CNlGGi4dkiTgZXmNbfQBLbatv77Mm7Znd/AEGEKiiqzJFP
oQG6DN0sVRQkjfr2uH5MKlm470YsSDHx1lESwUcwnZXNhiS5VvziUCCaBsHHOAQX
vI/plb0XEYuOuzL4GfZthAnI5Kc/pIF5PpsVDgdY+90uHtqB6lBj0QZU8YkKBZ8q
VJN6ELakXl+AhG4bpv7R7aGqB4ZE8p5iyx33ogVgBu779BugFd7BwVaViFWwLU9K
bgyMHFXy8fjn8q99JS60P1r/K+IMcqs0TSyhgLMNrfw1yuB5JNEstKdUq759DyM9
yaaflWlGKokVfC/Yb83y+7naIPPxjHDAehqBvHoYOwZ0mUOxg7f3vZL8xX66kZzs
7Z6fiCaZWWF4WMr9/oe6Jv3z3M4tJelEDDyBwQ+7aylHZD0lQ+exwh6+jm77cNP9
p+ux1v2p+D84HrOLDqUMdxx7pBPwdjublGhy8yD4ALwpFXkSIVIDjygCybtUdUjY
uEkppa1hL8PAZLzRw4nw1OXXVzcye1zTUqvjG1h4UosC+jMpyrt4JotcRHRUZLfm
J3XGy+3Ydmmq3Aqodon8QdUyfiNNjHJkUTnvC1h+g1wIqqDnYboisFazhPA6MZW4
VnP7iYU8HTvQi9+HXmlVzFAt4M+XURqxi9wr+TqfFsMouxgD/iAOYNP94CDVVhq2
VdcSdQlfnycOnu86MofH41O4iy5vBGmVw7Jb17ysxJzyAYj3gYlbnJya8/ITO/OW
h7yELz6tG7GQCru4Dw6xfZ3ECRZ5Fqy8ddrg4QlqlPOJfvc1Dpwq+TmshWHqFISl
xEVyzMGg6Jj95uAU0OakOUQRq5LhI2zf/R8FLrnllzJ/MR6XZlPkL+I98npzC0hR
rQyyztVCY48kk88svKLGCqHdYaygnfgv2lVN9LPRobVyvRwzbyuYKpDV6+nnpMuT
wCtTsTqHfo2vDrfWzGs+Od+boVdjU7XJjIMKmvNZhnBRcwaBsnvCguvztBm+GoeH
v/IQXLHuD2HsUMys06KLe9gYn5/sIy6k6hI0tGRzf6eA+vHdzJIuQEg/mpDoKiQB
J61M7rMmiGpcSF/EQcy5Z1I9MTLwmldjH1UKZ8l7Qyj+obVqmHN6zzrICRvymYHb
MKOtBQMigTQ363e4BzOOT2G6cZM83zdQJ84PB83VIssK5cP8JiAVnZlyP3vdrsLc
2sPGefosh2H5gtqeDlkwN4PzdqfEoFcFhEBWxBtG2JYTMeo5KVBgHegyohsMnEId
a6yRjCN0vRcXO3enWWbHwnsaqqMRyHNvEIj22efUYSBtoojBaMLq3E37j1d2CGj0
OPPqEBaHKbv+Yd7Z/hUfIpTuGss61iwLGE1sHlHqDB8rueiLZAX+DrRdSNgEpxCO
59RDxakn/wTOGMaJnKVP/Lul92bTI8IGLnxts9tHPuUT5uCASp8aC0jAFSwBZK6o
C1ZrYn2lLVSKR0q7dmTQC1zkAokV5syx4OlXAen9yp0HE1QG3YsHpmSzmLg2Jmi1
giCtzjZdd2BmyWT/XurTGqcLOy7WakFYseLK6Vd4lCxpNGCerKH58shrHTlImNrR
MI3mmX3Oal4+3LHeXxn3U2+eGtJc04oPv29Zen/H+y2PJY2etsyCQzX+5tNz0YPm
e5D+gjCrLPLtZe00F7+lf7uYgSYEefPBYkzQWcW/WL/pn9t2/y0kJDtVu1wNPYjb
41kUmhmBo85gY3n3pvZOcviz66f1YxE4SlYJnxstzsBsZccMCAKaoQb9OWWA9u44
AoMIbtk+AKMk1zG4gB7TVfEPWt5Mjs5DwNavkhANre1roUGyzi9zkotPVmUOdJ8y
AVsau/0zllLZsSq4p2i3ZgXx+yhHcOV8dLkUjblDPM/u4sFce5ulqakupjU7VoHE
ulOMLm2kthxO510Ldns9AdGgGscAJuuY9580pV219uw3n1VnyeVn5GHeveLRL5HT
0xPIPbJpb0UDLnJ48ROFO6gLg/JAytbQHY9oxSL3/p+Ankcy4KxVx2METV/wqked
kNtvqh3/YOKE7adBBIeRUEhMQBq9ibyY1aZP5kRRYXQKZQkqsWnM2lnieiXZrVII
8DgCnX5peDgAc89RAt8J7Yk5IR3NqDQiruUo+VuEQEyKO7FTd8chvZ7edCLw7opo
m4AfhnykIJtuewcntf62uBcXLnjRNkSdbqfhaLhi2pDfPhnMZHk9vXn5pPbZ1i8s
hN+hS7r5S3Id0OidY0GDF1GotJCdgTe91SdWYasltSZ3PbtSKpNl83uV7Stm878W
cLdrchaWB/mkv5LZnUe2R9RIASeMhtRUk2o/aHNTPC7Ybw30KhE2g7nDJFTNl/gp
ITB45exNzE25bsA6/81UbBvae7L1TTc4+1YiBE3OBdNRAjOd/yaeiHFDxNizcE9u
c8Pzt6hygJNx8cVh4lNOKGajN+zTKt8AbA8Zx8NS2eNAR8XplVHN+1BgnLLBKjLZ
39TbRb0F7R6kq2/UfXT9GHJPdxxugAMhqV+x4OOuam19amwYKDtSXHHZLM2ThDkY
y3ZbsYCdKESu4r1RQ8Tp6NQnPf97sQqZngwb0obS3q6J1l/Cg63MkXTHYu78vsM8
wwAklUsJ5njLxDb7xAar65T4Pr6h7305k6ORxR7NwZF7XQB4WvOJzuy7kX08fMy/
hr1YjAx4Xfpi8urEkm51x2aq2KIjl9dvZjxB1NN/zKB9/E3rBEs3S4iiv1fohzPd
QAsAXFtoU74efbkf+jdU7i+wUksrmGNzLVUK1y3odSbs6mhIVaFFwiXK5Egb4zfp
EuTrHaK8fcTah+ZwcB0vFl22PPp/AUzZZMLlbBy+j8pZ6PH79hurIrZU93XeNPOe
yNnMxiwvHoR1CJsNuv8x3GzRfkqL8Gf8HBgnatJN3FYBbOj4aU5jC1/VorlpPh6l
rrhXoYhgXWe8VCriu7H7TRWPwcVEpuS7oYuuK7s/dsmrI5TXf7hysrdQFFz5beHX
pYj9zA4OzinRc+Qvq2sBvgIhCUXNq+4U4P3utDuZxBvlKZGFLyYcs2D9+ylqTyd6
AK51EAmhnHX8CjwWvuVDjel0kuGK5bRZVEhFKXav+np97WfzDa9eUzGhnoy61Ipg
Y+c9JXe34FxmHu1GthSK9isFm7/pC5iLXvIPnxk6p8XlgOMx9DB5fDBTi50vS1I5
ykOg1w8FlRT/ZrLluhczt3Hh1yScNO9XpIzAgtCV4+Q/sUkn4DPpHWr3MpX6AtG9
ETv0N+ZkITCnPRAF3pCCRFoyyylLW2GnQfpD4UbpQcc6hKv/YEOG+oBdGPzbU7R4
LxosvnOZnj1fIWsTG/gCtJfUqvGRiPawjIXVk9/R7zv6DmaM8YpEOtpR1o9Qiytv
ZJnPZlmMQfxCTZ0DnqUXU7CoVeod0iS1afXmZnNOeKxpK9L1psT1pXYg9/UhyRMj
2opSsG2blzthIV8le0WRWLQVrrkyr5pMRLvl5HJUNYwF0ij+J5+eTCRJjE3JJX0E
C8XKCbzKwQ57DvsD57BmHiw6r45VX+Jd8oQPDMNReM2tYaQApeIJvbWgPsJKudvq
qGFIF6cwiIvK/PoIu5qLO91n2QElb97gnGGZYeW0UILMr5giZdUNGfWIZM12MD8Z
vrl4nWE3Xdxh+NC5ZNdrEXS2VQ+QXlz2dGXX+oJAajmn01wLMpIXuKFpUJCDkTRa
pNPXNFIsDpnX99yoIQ/T4phZhaQOP+2bST6Ebt9/44SyJEGNNagywpn8ta6cMJV5
17zRTJ8/MPXKg8e5PKrnlno+UNTrDPNhYaj0D/cqRuJitAleRUT1iy+2vFg6oCgz
NpD3lHkQNLOoQLsMvLhRT1CCsAOVlne1fNEjIMAnN+3RiTcgjPwmQBAGbf3pbxeR
We3B3YmEb7oC0VWTsZHrFhRpppVzd11N+C51UvEiZhklRzQsAs5ENLoKKxoQgsP1
8Lrf1GZ+lXLxz3Gs4+6hWQp3cAr1nhYivT/iRJs49E1U7jydz2NeDQcX0DjRDfaK
IozaChcaXu28VV8mBSzmwehMOaLq2iBpfNtCLDxPLbpcp860sia0g26TU8qI1ZLY
WFKx6iLU6Vh0No5hh3WG6r9dryoUJos197pc7w/e+Sm4XJozTL/HZMvnLb8eeRNA
oBPrHgRHbdbgoF52ERY+hfjccze3v/eviPeCYePWZtjGTsV/rE8KKKmdM7cCa171
2dTmhLdugMb8ioWGDiNaZbWORkf6ZsYd45maIm+Ek28JZNx4SdhDPb6+rKXa+Nze
E2Bo6gqNbL47FAT5RqIWiZZpwrcSXH9i0AnGLyfpn2DDizaD8tRHmYLvatEJeXeO
sw41WKoMGpfX8+nOiGjhiPu7z1LeHFISaJ7UeT2oHZvOLTExK+PVRNyAewRZgFbA
g/dipvYf6vV2EFBlOTokQrcYe4ntbtYGrxT0vJZ1H4/mXt9/7cOqiixYdrOGUfPG
80Ck45uOvJuGFDJOAdC+4F32uv/Hmbl0T9noC93rQg+zm33nCQwdItdhrRpChfEk
73/GFbdfDCq+whsFT6RlXGprWE9RS1mjjH/QYwgJ3VG0sZ2hH9f3ILHqDE0Kg3Fx
mmoLKRMxQM/7L2kbLzW8RKcc8GLIa6Ekxn6ue3iHYAhmBkC+FN70+pmrbAgCY9jY
aCpMDnPtleP9SWHWS/TcGgosrzwI6QJrbRPyU8hxDi+xRlxvmaMGrG+jSOzS6PlJ
uDnoKC7a6rMODEBNKTl4O+t+Va2/Z2Js2/9ls1CDf/SIdkoGjHRgiU7P6ElbSF6Z
QrHLfH49mcjlcOVcDEotmZ9mWkEG/CJ9UkaiD4qI5H7YFrOxUCiwnoCFXURVBx07
4vuLuvIK4PxYUOYunhgr1ntW3d2Y+nuNPdd5HAQP8czXGm+ZSS82VcWPIT44Lrvo
9S2BfKbvTfPbWcll2DEvBe8pOIIpD4N/h7pz9BwTbbVbWXv5dZlbvaQXpXThbj9e
qRr8Q88cg3gLS8aVzwsOkIUs6+o7yYbZ2VD3jvYODdOjX3xiLfVyqq4DXF4QG2ZM
9lEBTWWO+BjbJfh4xyzJZw==
`protect END_PROTECTED
