`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYwlnOM19Py6jeK6P9Jr2ytbDNAxawwVNVkftVL7b/8KAiBauhQHSZeK+8oVTtdT
37BEj+32MtbMKwCaPDAJWX62N5gsGJNjDN594Hm7hOzfbQksar5gG34e55rdb8Ad
qHs30vCLyxq71urUB+4Z6IRfnVxtwPoS430OXQUP/qYvUJbpoBdSoQMykSvQwTnr
UGjjcmqBqO+qFGfAOg1vZguBUtIrm88caBAn3tLLb7+FInIdRvFFsEGOv7NvIPzH
LQ89OHZngtEoDzL8z+/FeVJYa3J60WQZZJ4D+Tmlx8K2pMjo/YohAJEJf2UAEeE9
TG9KQ7deIjUHAMgnOR9aB8ARhEWXkTuMQvly6Gt9lLHI3vKrm0hk/3aSdlR2fFke
OteyUtbKTBvTYr5Jja9gsxi/x/LqJgU94P/kBRIaApcCpd542Qj+QsGGKM5iMLG4
fhs7rPRBWpY7OY5hyqivf/2cBox2/bJkTPx4WWu0wyMKUGyWf5ryOYnwEvOGfOoh
rAP9BbtRvQNaE669sgINOPlR2ewb3Ljoed7f0enZGtNddSFXAKXZaefk2ONHnojV
2WucaQVQCVSzIF8HqJp36A==
`protect END_PROTECTED
