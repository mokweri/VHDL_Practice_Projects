`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qlKU9Gz0lRSYhx9DvwcHyOXbB973VOWWx0IIBPeAOhOSzYWBNBx1fJc/6YrxQCD7
CGKHY872YaFbId6FDbz5bpO7usOAJWdw0JnCPuAVFgJfo/8nZyvVw/306h1peVeB
pQE85LDmJHaYcE/eUVTNBMplp9Pf5Nt1ySqf5zgIFjx3D6AMErh/QVr/aIrwak/H
WArJQX6yIQfMtPLuEpzFqhHMg0/iu2kanCqQh4na3RGiTcQCjxHY03iNKOAp77HL
DySidZUtMnCNhBGqwepJcEooIeThUzuIrpymWO9ZhMid2SIUEA3d/IVih/HAtY9N
v0rjtpWTDpRNhABuhr0era5l4Pn+8MkPzlUppyyrkuB6xfo5UqOiKIo37VI3Dr87
iygQUidIGyyfMcvcpXK/X64MoR0rVQHFfA4bvEUytkzYnNQeaPwayz94c+0nELAD
4ZCM0HYKMa4SEfm2QIQA6xky6iVhuzcnLljm6Lgvf2kZx8NAfDXZgAwH0pNO+mmr
H6GVWDyxUa8UpNapemeTRbv+gj59M17aqqfUgzOw8uCo9/CG8UwDZG4OApjKl/Ff
dsP1M+OLw7y/wqVviwqdYPQEIs7tyN4llssteXpL+tgHKH0Gl77O++mEYDHxIjhW
k5rwBfNilIvf1NfsbIqOakbmaxG6me8WA2kczJ2XH+UYVYjx1sRLNhl/AM9nPU5E
nKn1kilUbAFtRHC9n71Frgcs4HAaoImlAUzxhNlNoqapZyYNxpb0vafeYS/ho6ET
dMqptCL7UAIFwP3zuqIT4zfnWS25Lbx26PeqsJS7rcd/GixC72Up3P4h59YLFdLX
2LSPO4eeFxQBoSl3dEedoNFIKcHMV2hLdoaXFbo2S32PNJqkdb9p5r3ccmvuJKy4
h+aFn90CN+5HLwDlyX1v4EJwyAq5iOFb6otVAKEbJYCrtkPsi1QCCA1ZuCmpB4tJ
CANC3CEVRiDJkQqOfPyHZx+zsuEcQKBCYbruN4IkXQGKu+VNkoNnXXjjFdoh7RGB
G5rDLkVUFHk40b5HKdPGiENbENS2F57kdEx/Pa4KfriylIa8BNBto/FFhmVl+/5d
2d2FzZhFckM1cB+hH+XHu+m/z/cXImQfcAFZMz5b81cgEUG6gC3FrxN6AU6LUkuK
8CreNuVWrk0obcQolcTs112/ovtSdl617AWVUuUVFIXoKki/7QvWsBtQkxHkfkEi
hieZj2UPtEN3hgqpVsKJGDj49RuXg8tyBrFyx5T8Qmim3mVL7qp3A4p1qPl4jmO0
`protect END_PROTECTED
