`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XvW2BTT2r0AqkVdv1e5iAVvJoONTwH+D645Nq0ebLkaW2K49CVnTVs3zx5LX7iek
vT3nndF6DITRrKhxEVHFexHAc+617ky1gY/Z5zdwwywXVH/gWrxogPkXVmLIT6EC
unXrIcIDPrAJho3uiL3XKQh04+xC1qzwdQOoGu63mmtdO/509Rb90QiM9CC5eD6H
yQMxTTKO34WboQbrIcb00ODTfu5NCPTQGtRqnNSbZBSX3NsxsguteWgzUJ9ykH+r
nFa3WBlYycd8deV7IlSHh3pcERT5oXgPCwE5QAa2T3XzJ4ifgij6y7IvwyIfHAQB
twS4XBbz3WSkOz34JCeB1ZE0khmANHBObNiZA2iLEV98KgGgiy6PJSElimWICBe5
nk4XCYt7v72pA0LlTK3pdzv027JHxDbyLkY34+GZF32QTusAHnY+Jvs/pdFZRQMz
6L4IV5Y24ULlz+VBBMKICFE7dloK8YDPdQ742ypo6BJhgh8EGJw9nCrhjKbKqDry
qvcduewXWgz4R50BjxKFxFu3Ukix+M7bmo6v2kgGBjp7NkkxeSNJqcQITeab97aJ
gIfUsyd3yJFRlsO7FM9ozu79pum5sYvdTt8+O1rz2Fa/WjjXuiVZwb4XcHRXwe/8
lzfp9STR9HKf8fa6fubG0uIhkeHG40GoRKQL3h7nQvtmDbw1s3B2u3UNVopitg4j
ENMvNgHoo0PpRfzE31CzUh5y1aMoWowkKOjoCygb+L/57QC27TqXYcFdBnUXx4Qv
oHw3Tg89MhMVPjDVIgkGPaP0I7AA3gMZFCdwLn7NT7fQgwoFyVI75qOiEqOnKNL0
lf1f7VAW+KrH5YINku1NJhj2eLq76KN0LCsdt8gYcjHO98Wche9LkYVSmLTdZCJi
0l5a2geDMheom/X+znMr75Gw3O+GV/3KjAhcDzedtka2Bs2Ko87hdcg35TYz43Nx
2viu+gFKTAiYvhjguQ2TVe11FfrNwMtQzekoJU4Y6ZaA4vOXvakx2T0/zc9/AmJU
XbnycRL8FWIqQIo23IdRrN4QhEMK3UeoAcv2On+cLWRfrko7K9R5zf21Crpg4/y8
gG19/SfuIdpub3eaazpkpYBnXTQPs975LVSrmqjr289Kflb71GhDReeYDT9H0PBN
sNanO87jq03FRO+uL2Cap2BTbzCobFZBjVNeYMpTCNtMx+dz9C0MgT5xZ4cAmYZj
2OcKbgCd7Y7rmaOlr5xW+j+smZNbsE+l1gGba6LXPTpw1wUZEFFPgE0VlDW0V6Vo
uSCh81HAvYThJF8I4+RMhMMxt46HkxPlbUoGs5AMyg3bMdNPr7+JjOGxeRqFvFsp
7HWHAZosl6GujWQi6f2XPAx2j+sRI+Grj6i07406J+Qeoxcg36MkqbA9yUWEf0L1
xGNJACOje1VDoVqz60MqFYXGVlhCCT/KInQZN8OdxuqolP0kirRgJCd/fgfWxROQ
cWofa//6LNCkQhXPRCTtj0SQlZ1YyGPzyzdTdy3Pekkqqp/TYqhnW6oFfyc4TtDZ
I5fhm/bp/DnHlVYEJSSdVrHmLtMYrJj983wkdYT4yS0UWE8zBQoiTKtsMFwaJfWh
j0k8B0wmrnT2isVXQY9hLwJSBeC8uBbT/4gfwM8wx08/efnA/y5BHC1y4LssgiH6
nXtXYmAT1pR1VBPYSLW1LafGnMhWKL72xEyNpiQ6PlVinNkoCQ57xaoAM3+G+Uqz
cH261DutcszSGjNtcRwi0Ffp0Mk7UsCZBK8pmLAJY698qbSBBMFMHAb9tDACfyJJ
naq/HuR1ioPxjH2telnUHwoJZ6T3ZIN0q8w3RENosg8/+IefOmrVtNiE15ThXrWc
9jgQSFUMUdN/ASTdFlt7j4z51cPxdosYH73rgPUfY43eGDVVXDACBu6WfD2V2ANP
ylBFmvgCoIXkOsj3uf9UTA==
`protect END_PROTECTED
