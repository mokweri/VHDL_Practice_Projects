`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFl4cXfizh9GCJdC7dTvd6T8DfKTwQ3sy/SCPoF/FcVhjtroXVLWJ1QX+Iyf6hXc
ATGLEaCJvgT0Fk6GGFSBwdlbkRlPBsmFkO7xhmgjFRILqgIPj0782QXXhwv8Bt1w
xtN/ePyFVo0naU6Afzo0tB/PetO8Knezk9l8G78Z3gJtl24b3MHQxtpcEbJ0Opru
gFhNcUVD5cmiI3goCaGMEaLOOxD3ubFT9Ab2JmSOh/WHpAeHwhwQyqM610EcHi19
QIueLIftTksquw1o89kaz5OaLZJMt8wtfjRY4iHaVIBMC/0jIoHwUWT+z2gIRliJ
3GKevL9/O418Zo8eU0i4d2OaWd1oLHVsQCvtSUZkCZpnDQeDiZvHDSV2AP+KrAMb
h+V+CwGMtqrjlHivH9oXgiN+kPGzG2C7P7OHYpEd5VhSvg0gJ100n1N2MphSkQhj
ssae/PNh6avMyy8YrJHaVS1liw2thcVCfMM03equJjfmLazY8RAWP83HXwtLsa/y
XpTrbNevLC4WydA2AU5UYJ25iV3zsIJ8BJUY3s3a8HL6AnaKrmzfuuvYWOnyeflZ
ipI4gu3YbCcU8msHkHW6RoGGZn6oE9whx00klmgcyLTuaA49xhSBZUN1dWcHLDJm
urOZ7BYiAUarLpCUXt8PwBh6qPudiYe8TiY/47gvZ7lo8zloSacCrBIQzfG4ZbvN
wUqLnFRpSg9I1o3zAnwfy0Opo5Io0yklhoKeMQpwu7HNMPbctBIb0CR26cMCu6h7
d2E/PskKB0Gokf7UzXHeHg==
`protect END_PROTECTED
