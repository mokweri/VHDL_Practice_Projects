`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQ7+S7fQ1zPyq61pefM9+0qY+Xh8eYX9Y3tp9+PiEHotm2k12UAOC5F7W3XoykD1
p1L9XzyNhgTT9OmLbFVMzRlTyd+I32x99uMaA7k78+hA4lVMGhdMQ1tlOInDXlZ6
sHLXZ5NESaOGSrcP7Y4u3XjP+cMYEMIJczhDHPxjh+xX/MkHiwacsy8rciuNqne+
OvlTe/NkwHtxt6GXMYkQ74/dbFQKxIXAZaRglZD1q2avYdBy149qLMYxU4aoRCJy
m3z8Vsrv7qX8iFKKY5dSZedLC+811C0tzQjE6pI6wku7mI2kSUQo9iOPdwz7Z/Tp
NILjL5rgEkIby68BESGzrR4PZ8JCKJqo5zFtNwi7pwI8BcKnJWSHiGTN8I3blQbg
SY2XfADsMatzlQW/cdZnGSWyUE+BuOXj5WAOfTRxEY7pFGJbXXFRtMo4sJKSBS1r
dhYYtQMLGhL7n9pCyGOJ1loAfteSyvcU3OJSJPEtbke88k2v5sThf8cphl2pCTwP
GDWR2otdKF6ID3aJogtvTICnqPck7rc0oy8bDWd7+iGZ3LniCfQl5nSb24KWrfxF
T4v9IAlexiow9P+hLFCR0jW0OlfMRyJumgo2y8c6lRusIxqteCm3qYPRuObcBmj2
fCROm27zIrlAPbJPFcOdZstbpu3BMiI4VhhkfQvPQ9uHX0slnFTLMzRmNzrT1FS5
SthDfAwBbv4zFzf4ko0c79PDPjks24fivjJyA/cggItypYdtOZ/s1Z4YDg6ZneP2
M6ZQr/rY6cWmcD74UmqGieV+CYWy3a8x7yl9dkwcFV+4tUdjngMC620XitUOLGhQ
apDGrpYuCnw4JOdCRSXdLbAjp+gevBL7HD/l3Mnpg38iZ0X7IYVV69YlPtrphkxO
/xCvbyRd+IJWjdeXQd9yRjNE6orYvgUGlr5e5GPueHNxkHxaInYM3aNnkmDQuY2s
niw19v/I6yf2UDaU8r3b2eUijoHnWf+/pEksnbWcnT/oGfBcQgizP5nfva43yu8W
0y1xrqBFDdiEteB3kqh7EvZt3mMVa2SlPpsR5W/EUPnWJFD/uFpQt359rgateNOu
W/bnWRbtM8EV8bjovGEN5x2OjrGQkjTAF6sZFZfrwwjc3y4YZ74smQiLUfQIXwz+
M9FPDvZPPK/MZreEkCS3ux2OuXseuhJhkpJAzPXZZZcaotFR8lxJrBAZ0gziGNl4
P6ikfaNfLZrQtk7MxiddfhiCOHHyG7tYEBik7TI3WQltHRyEMHyVwq66y7+wvSLF
3xrshlMnGQByWRG5v13YtJOHyj584vvARQxr+uEXMNfxWR6WmNE+9qnPK2Lso8OL
21ACWMvNzxv9HgTBoAnDWU4rfFPWw2TDTJdpybVdGnvoO+hGjfvQFNTjVn730ywH
Pm5szig0QUdsGoAAk8XhCOauZ5a9kSehda+HdZsbrNuQTZX9d+qbLMt3wcxL4mp3
Un8Yo/pmF3lhLQTSvGEiGA1I5InwU4EVAvH1G4wlS5DlB2UNN8gCTjWttV00/XAc
wLXdEZlO19F0GSKxpZUvoLkYGxFrHZe7s4rxqGgiO3Go6LLSiJOGWN3w9PBmcNeA
VjlQK0eF22sLd8wdxIWdWMLgPCiNrVypebvirmFaoc34IZ/Tm9+rdECgw81ZoLJU
Xw7FN1DSmkN5749fss9bskmNjAushr5PzsmkLrBl8TfTC5V3gQvC7OKeDWWob0a6
qQYR8PVJHpC7RPm+LgnYpNUDy6TgpsePkNstxpGL9eAllSKBTAbbaSBwuLu0WAE9
GbZmP7jyiWEgr2TlSEOmbZkBtmvJ71oDKjWkaUf2k8yiCADtWbZoiJyMBrZ1KgTN
xiaRigHFLO9wQpEtIQhfOFHtZ/sYPITrR+VEWbh6ATQM6eB+Z2TtQsRA69GOIGr7
WCf+Si2GY1KNHLT33b0/gSKENOjOzUocjJqep+4gbroE14cIdffAawvofZ4YcZUz
n24SHmNm7P8tUrPoAkw6inLkXA0NimWC98ZoOxI95Mrwdy38bqx8ZfcdTOY07KqP
eeyrsURvP/cH2HgujQTcHUANbtQ1ZEFm3NFvh+cDDaYU2cBnfJqSGlGDYYXJp8e6
NS+UR2kZDe9KlN/RbuVXeEHzNfQiTNBlXWmZ7e+TpAHQtAZc8R50IgLHeczBYAXP
50IghcirMVQIJBALN3byoLrPSSJh1azOo0wqezRv3U7lI5mIYFREhq5HdhK0uqgx
5koUEf11B8jYFnDK17rhOUH9cl8ixB7H1ADjoi89OtzDKUaTMUTQafBWrbAvvJVv
IA4rYKI/ucaLHIpsZwgLs413SAfjOQJ+0a5VfN1iXtBfv13bR30fHOfo8wBtBBYs
LamrxGRaUl5csKXWhrK0yKQAIRNojDmPcRgB01McClpII47gLq1o4bw4CX6n3qrP
HF6/3m9tHimBlCUrRimfkF6RGn5ktbbgODdUuuL4PrY9al6bsA3r+sfjLBohXBDB
f66pe8Kxz4fCKOwSKsNO4Bcy/kkyioPNS8Z40uqUcgoDKaEyCF7cxn3USCUiMZHt
ILcRYHZtE0RFCfmahuqaoyYPYUa92dxE+1jszxFcnI0jXQG6pNjKN69MyTqwKbQD
ex3CjVeOi3qKbNwHWHhKZd+jbb/nAIcfssGJ6Mr3mW4zICuvCqks5zI8zBiNLOjo
WhYw+IWalUwL8SGYiM8jzFwEUjUdeSA50CWkVrUBcUlqLG4RwkFl19wd/3IneEAp
28bSPlkwv/lm3cabra6z8QDHX4bV+uw+7RM1au8+eihEwD4xQ+hl465HuH1Y9tuX
ggytLbpQtkJ13dJPeKIFHSwu3+ASq3YWlc+DjuQNYaOGpOVDW314JuY+Ud1Psq7m
5hltmenWICkGrnoMF5GZydTd5HniCTgSaE3an1T+nPIWl3yh8eyNGU+gB9WQHE10
xBc4SbOIEmePaGg2S8hTAi1WEnpoejYLSCWomQMy57sVXpkxwovSav5KqY8AkmbA
4YL7NzAbJ6vL5UXkj73dDxbmCw1W22EO5+Eei1p7G0OGp7PHaUxkxTYFC5H5F+SZ
hp8raFsLJZOt9E1ljXUPzGcGFaNBPQp/RVszX7enqLbQKS2V+r1czRCkRpRs54U1
NPlyaryU/a+NzKbeyrBbjevWhgR6FC3TfJpOMZ5GRwaBauJbgTSb7+7Jlo3ex80F
l+jbWZZ9hpXhT3LVNVq/GfyYbdE5EW8bKSt2gbxu7tsgAPwz28hUL9DT14mogYOo
uQMQ81GYzDd9iu6OEcBRpyiCKq+TZOSSL5a/g6YV4AM62ypCfe7H4pBYYNT+KfZu
ltOtuxvXqiD4+0VK0XslMdqKzKc2OpuH9w2whWGIA38qpYlKfMln3cmMGHNvZCDS
iuV6vHulAN43CId5as3gvVhUOx6ze14OYsQQD3UjyXzdMWfnIMbPIZI7b80wYVHb
5EFBv7cA8DtG76/dgjxKZO/4GPeXCGDHRp7Rv08TiAJHonD/dQvHkLVV12teWQ8y
WM3QnFMAzQDTqziWz7l7wotH6eq0luiMcLZAonLRAFZ2D642Phk8VJ9AtuCqjCtZ
6d/W5PB+P+h0IkUtjBWcFY1SkxC0M5yTfg9zS+cdX6+wwJ6fznx66F4kBo0u1L+G
y/776dUCm5jYgNTBEJEcAMV/+U8OzOqlqKPePdABqvolsgfPyRp+i2imQbYuP+pf
VzrCRDIRw5q67gYAlrfdIbY2eC0f4JIzjSfwSFtXGmDcI0SBQrzd/o+IFsL5s/8k
ktAu6LHMj6Br2yeq5JV5L7a8Ff+0ScIKa2lQ8DQ12i/0OzAZa9Xg5FN4akaen+2t
MQbXYpDhZwIOHQzJP8fFl+Pf1EMZ2sRvMmEzT74K8ut+Kyd5ZTZMoJHpsqCCX1k9
Vd4DJxsH81CfmkIHMOb0Cvqyr2UyZ5wGJ6+5wmFK6QpELr96avOw1/jQBhOCG4CR
tCW3A07DC4MKrGVP3V1frGFzXAwDCUlWUIkIM8ElbrhwXHSbIkKTjJDfYIthiNJM
Hx6Mv5UFD2EbykuhLsaT8C/MHzctpPyGf5JQ4lvXj++p81csHW0lO+uxctmyUudh
6FCnYgItymM5ofCpBPq2Xcqd7XTQsNQz0ULE0vpaZVf8vsyLO3PDw5eEQrzPiS+3
E0mqk9z+CPa8tBNLxThW2PNfn4J6STNeXOITwxvs2H15bHlcOp3x0eYCzlYJo6dE
xyxyH1sqDm5jbCoSB0CIQiqSkpCepIdryQ+RwMhBbUN/sHsloGTz3ZMwrI9lx3vM
84dArnrsp3x6o9yvUTYuDkYTro64esZEWBsMPBAEq5bsjqF6sUfwXJ8jSVHe2sdD
VZ9P1SQgwtKiwcBaFDL+FbUyEcWmohLkAsbFTdGaS1ro4VlgWlmOJbp1e7tSnxhS
3LitsgChQEroTge9TbovZA21HCMR+HalSVoe/OmNgF8i1zTVXwDuyKqjfHIctP5n
cmONeYvtcE52UFKA2jG4T+dVoFeP2HaXP9CCYt57wSIM4ebsqYsDZreCPQNRUTcV
WXIpTuLGWPF497BwaoBy+0TADLdPOr88ggC331LpShws1+NqIQ0/82rc/jpvf3CJ
krEyDm0kE0nmwsI23ti9mU8LlzVAC4RgzCH+W5vuxObws7ru9au385axQ8+d4GTz
OcXdjjuCXE4cE5VfkOYxjEH3J+sygei1t6iN1L3FfSRpNTNRgTf0sdNkDYS7357C
oDmGK9Sgpdh74x6uAq/gi1pf/ocpJHbt/4jf6VirOQ/3pskva2nvm7hBHa89vSXh
iSG4ECzeLXXgzS4XKssJnUuCbMMbvDqPZvPW5QMMALYmaQaZdxi6u80IYIv94jZa
KcY/ssQCHF7vP9r5t27j77Jb/lhn5DfAac+faUQkhd9TYihgcela8fxJnOWscTOH
//ZPHQ4oWYXt+5YTaSLWDE0xNueCs5TGNXcVkqeN0qg3EGf1Lu/uK8ZnN2eWNqZ1
ENlE6ygPkhMbfuD5poNQ9/Kl3YHYHINJAyHBCMevu1GXpZzhiM2RJUv8Rr37z/Bv
SWf4pqjfXGYb773P/xc50wk/VSdQT3F4fimK5NvyTRj5mJnJ/lWX0nHqZTqaLve2
jINYWBcJM4Dy8lFHE5wevRfYSsFS9Xk8CwP3oPlrWigHJwwZ/OYmK4xrQc7NTwGh
WLTDOoWvpB2+7dbU85FGzS0q0CC0K9FYh3fc0xXd+Q4CPWE7hq39P1frL/e3n9OU
lP38/mjU48IVG1755d0z6t6QH9BO1RChqnvVl27+0gVDnSikQGMtWcYpCb2w8eVW
QuXKmaVw/0+l7bK4L2aYP+5XwCRsS9xqFGTVvF9dR2cK/rAwb/BTwBAO1QUF8vzd
E0lz6Zx5mWrOYFxnPHWeUk9+8zDQWKzmn0TF0qwuDy6sqlhTujDoq5grJlEz5+Ax
GTZqNZ8Qm5WICiiuxJbb85OQ7NuLVMRTIIcagBVAH3EpZteQ37QOSE1H2NDKCYEk
/ADVuOcipRLFq+2G5KcYJ3hOEHZOnB30EdHLtQIDKPDDc4SOvhp+HEM7LIfofNsJ
w7P61nOilRcoBr0pll4mKu75PpmiZ4tlZRd4NMGTx7iC6ncaGdK6xeNVHH7X34iv
K/1AikqY6xTn7Aj63Utu4g==
`protect END_PROTECTED
