`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iZjDYpJNj68XZsAcM9kBLQghqPpKNT/sQVhkuL0ppSUoyGHPqtNeeJBmBtSklNW8
pscSgrIBQLEuqT/LOSLiM626yTAgPfsI01cQAud7ayQZrVIpp5R6bsOlKzhOnFcB
dw0nKJYLU/cEFe16xcuZkSJqO+oaOyINkNnfvgNpmkKMut1ZR4/YP8DI50PY4d3P
f40GNdRh8V0dpoitWR/ceSqctXsilouRkj3e8cDwwevn/kCOZzmWnaqzKXtC2pXz
At+5riN4wgAlsd+P+14GqcMkufSV/N1rCWFHHNxeCCcppah+ewIgLGTae4vo4S47
eAOZ5Q23VqW5L4VFHelI7kkp4EBm81SWV71GkUhK5AjzQGJwB9OKf+cm1zGUvMlT
Wtwpx/PFwFkuPzOermsMhQN3AbHcwt6SCRzy2zCSFyT7iCVaJtj9rSKPJnmjdgD1
9C1BCroft/gpFoC9ekBl7MXdHv6M5QQADo0fWjRN+PocMZKdPLP2MsTrqlaTeS3i
UKcIQ4NlaKUhJTnYqiw86mQinydEYOuR5OxOpfhMXxH952N+Zkh+tiYs+WfWswDv
tSyz6wKrAUKpS3/bwnBu+Ziye7eN33/YNxa1A2RgdouBVgaQkDbCHgzJKvifRkzs
9X1AT/D7dDI6G1+TRH5QQho2Ues186aOspuyUurPQTTxUEZwcfRTIgTLs+sFRDHI
fXzB49Ya5lyfuptdm0HmSrq5s+rbNkkzeJiukt6qKMM2TR+G4VWDozAA8uwtL2Rs
0E4evVYa7ZjmtP9xITdYGhFFSNP9Xrkr5rA1itdp1cG0a+fzvOD5PIA26nVg3480
kcQ9M3ZLj/4MlbhilOutb/yJO8NIRBJ9Cbi3wOipxjN6Pa3TP5AJTDirzNHJ7YB4
rMDdHrQHaxZ3BiGPHeBULFrFif+lta9CX/N0nWi7AkUonpvSlcp5gE7JbmKJ1ibB
sb7m7Vao+A7mZ2gRi7SnacjHLnltCvgKoJFfhcCGIiNyLcX6h1uuQAonBJSyL2T9
e3Jub3/hzeTBDtas728pOi1HSh1TxrBHcB2Y3qxV4JyaFkJidkT0WmoJ7aBz/BD1
GIl5EPTEW/jy2JkZdbA05LsOF7eXNPt9L5VIwJ4IuGyAJR/iwgQLQyM9Nm0koXm1
jLFsMqrT0/wP06mhzMMbyyVCnwphtFHKVBg8yynTr8DbVOx/ZNnDSMbLxFWTPQ0L
WajPmfkMBZmHXVP/nqXhzjMB17IQmB7oyoeNZTqgUbdwXQCsXeLXL8RguOxdssm/
jn8pZjaCt+fXvrRVuAeSNmB1v1M7Ho/l8G78Mq+5wSQMJR9AJU/s8WqVjk2teaB2
wpFMtQex3rF5KPADtX3EDZqJNqEPXuLffBDdVWQyzsBmjt1IN9zqHNSlfUF/Qi3c
1lxGugkKepncpvMCuwZGV5TK2maU58I9h2Dc6jv6DG+1AYr/Kuj610RPXw6dhkTd
CgZJ8juE5TfAsrVQrzA6fH5DqTkFbzG7R5vJwmBjq7qsQWwB2VuKZG/dLlL9zBc+
PIVtaAWOxH5x2LKD5XDVf4Ltun96Q+SG0rUUxaoBTNeZyW4NLhmgg6anmmVNgOKA
a1gj2wuLsNj4yNskbUq6Lmd3q3v3Dyj3oZ1y9IDxzYMT4mWM1g/CugQRIzJ86w26
EtGJtYw/OHq6cGWjj7FXufku0q4zFRMVunq9CNw88+kvbkth9P/y0IqB+cJ5ePD8
zkiTlKO3JEJik3qA82kr/R5OTVMW3ghbyaTA10ORT3y6isKbe+K51rfhBccf7J/4
jfe662L5nJx7iwOBouFsOHngxyESv4MFozWfPqhjPNEpikCo6+H5xpViZuchPYmI
R0JzmNMggoZZeKr8cNXvFnoxULmcz5m3bKGvqdnm2Wnofk/jFJH8FQgQ1fx9mN3t
AEWjNqu8kfXrN57yknvchCuwJrKgcxsgw5RuJhbqD/vwDwgwRah5YPpoo0ge8bq2
lxDiIA5gQ+rdm/sthX+It7lqfu78leDlMeEYPqZSBNUbpn1GsMiho48E60v1QGJC
9tlQwvxzb+slipk2wgIYwIqH5vxX9OalsrZOfcLr3leZJeHrKwJddULdgYA594CD
olRU2m131SjC4gmmyrVD7aZx0a6Y4yW313nKkpeB4Jwo8JJlYUGRbm/zGN7LIC/Q
AxQb33VfZfFOEnJEKRNSy/Sff17XcVf81xE66Q+q95/BzLX6epmWB9woU7dMjJy1
r5drkn7rCrIohe/ePj7okTbcKos0s2xFg32teyK5PiVkziAsIbfO1dNwDou4P2zv
uAS8eLXfLuu9Ug1/HrCd4qTAwD7Em3iBNyqKmqEe2L0MolsnbtWknl1RaA5rAux0
hqCgRwqaj48GlptJp0iu3rY7pFigyLVSy/eckUSnr237EYY6O/NsAmSpC1gTyJDo
wdOLq+Usc6mXmV3ZyNeuzN5UxVCgouR3XpVom+06vR46NZwDCOQ/e6MJzUpeqkOq
PjWR/HPmtR9TKhuDSYj5OO6SAJBRBiCcruFdsLVexMjnW/wjG9b7W1kK8BlEckv1
8MHq5QKy8/n2dnaBKYGpW20sbVDJvpEfvZZ0EjRE+JVwl+EEjidbWnGvzMtIM7Y0
KAkeLUMhFeHPOtDmkkvXk7RMqLADjW4MlrqoXbyikHNnWO3rgsb9O1nRnoxWG8JO
fUPrMwKXJnoHHxJS+CpdZHXdtHKQKBudT2C+dG+zaNjjai/yOIL6Q7dUdUB8aNLc
TqUsjSuz1DYaS6oZT78+6zJekIE2ewVbf1q0DeXijuNlgL4EjbQNbEgrzxX+zWg7
VpJW3ZwllCPV1ljZsIaIXcRb6TclSs+QQaoG+HdgTlxikKW5Y3Ha5twKqIVa1WSs
0ROGGVqfASVglWBiWTQLHwwLzwrdxiwKelBVpFLa4msO0yMTmZIMgyYw/TRk4zAb
k6J60+q0NPZweRhkt9CLViyVClfBWI1bzglXPlhJMHbELicposphJC72jyWJtj3s
yC50uEDKtmHYjsGmy3MrPBJswQ1W9svYNsKAy+DEfB+5WXG+9ybjTbp7Olq8ap5E
ZP2x2nSVu0nZ35WPA4Cj/U+bVD8mr/0d9otQSDQXJGcQPqJUKZ+6/jM9Y3qrIkg3
p/bbMRh5yB16i7JbnCM3U+dvsZ2yvpe4xcq+V2NohBHGMYPXfmn3fPbLG1rB/hVm
XJDUjgpiKH7TwHX21GkAi/TzL/HkeM8yhsv8ZpWfoItM7SrPBNM98WRdcaneT+2Z
gX/z+BMHOP7DGoKcLAFYvXvcgJmDU5aOmTP+r4G7Ooownm89GmQYjqXCIqTYUxVv
uBWAiHPpBHzL9+aDP1kqBSwaV+EcV9fin6VpKZ3QlPXo1PZhCziLkw5zxIzjiMTz
f+ZTt/NTL3nPBx1VGtbLKshmXf4lY8bdlv4aw5ukzmyqeD5zPe4pN3Vca0sTLoVs
bbEGugy2CyPjevghuIWXUuyu8RTSOxYDCThPgsEwi8AuGlt6HTjTkfbEnLd/toSZ
4IaUJTXWMlNnyRjLA3r2ZNc18Q7NZZTGWli5nEymvTj/PZe6iNLt+FLMnVfRPvpU
/jelnC/byty4+MbxmhNOmlSo4aJ7sBR2cXp0MAQRyPExG9i7WI2Mzy/aHEzuV1DU
OSvy57as+dZ/ggVlFTjJsEH7Rfwl4LNrA/Dv6odZqU1G3/bQ1H3hv38TfXGWspqi
t4oiM5Um+R0I8dXAyInmjk35DCypzcMNKO3mDOrkLlGe8NH8Y5XTPheGPWpzAm4R
+uQKziFHE4vUn1/4/OGM1vQoZeaugIE5SMlNEa3LgAadlpPlGUX4U7+p5aINprM+
2T2xVcWSuaFOnXVM9Vk4joyRhcdcVmGBCkpvwjj9VLUiVF6Bq0Ei5a+gQpCEN/fH
7XpfaKG2JIxWOdLSytYWG7N7mcBZ3RZ7pUHFlzPw09PZLxUk/ncfJq42604z1svr
9DfT6NyI+QUBNGDd+jHaw4LfdLJatiqhTlSMZb9ZOzOxdrCqHfeZfwjw0vKDxZM8
AreZX10CrVXRoQ44qmmtRle1+r9p5j3s3SI6PmGIgPWmCFa5LpwStHwD4qCo6KGi
eeM/hXQ47XTg7mfSjzK+EA4b71xfd5KnGyUOUgn/W6hT+qygpqXCnR24nRi19fNu
CfWeIyVqHNBZ7Q8uuJj7EYKMIBNFyoLcQhPloLN2l6wKMqarOR5BTFx/erk//fpC
fosCMvU0frSS0VSLEG3QWI0F6blzGeWy6Wf7wn2sqAZkK5CkjhVx9OJRAygvi7ki
x+I2IVk36goT3kFnhXH+YtAPuTHvE7jv7ZfbzezUdNYCIJxjR7JqnUP8pKNwNiV8
UEHzdRLmBRdx6RR1WM+hnIZas3j2N1Y6QE+nWzuzHRTYJrS4Eb9wCxKMvBK5U/IZ
yJX66ZT1YFfOiQNmnXAczdUf93EsOE5/m/JbF5jcKtW0QZLE4C30h3NRQb5f5o0Y
6hbQruiOgKxay7SsDK57if53b49YhHe/jBFxaiUJsoC4B/nojdRrEDfWnGHrFGqr
ujmgwPLkir7NSDq8U4qqSyevRJzZwwt9IU3cLSd3Zt9d1psspzPGNntn4M8Bu4oh
Bi/QTFAmWUHV3LXEp/7fe5kV82FhEyGy1OrhGGJvdzZFlPFlXAwalfz7cjLcir6b
HmmzVSs3ri/kWBjuhInZd238Uu9O+q049r7mQw4hEpnsIdtqx9RkukMxvwM5pCW7
8a6qtbA5pCGzlJmwS3QEi0KwGiFYptGBuKHwQt/x6HdoJD2aHUUMC3RCpUxfI5c7
5kzf7ABzLg6KXyRX/nMfXMvJDIhmNZnRjMxVWEIB/nHiFhYPlpSaDyFauq2KvQNc
GDEkdxizQ23bVUu4EuVk/sW9gkb8z3cOo3zVtf13xdeXBkGOYMcfS//PubR46Kfi
UKCcSZqkFHSjKP5b9pQNlIfSjMT3pyZTcdeh7WNo/i+OKJhvURkGbKoZmXSkVsiV
Nfb4jybBIMBUWkfu0PfY0jX/g1tZl+ck4p5vD5ICGPW5UolPtin6K9efszhq2XNH
VzHpMld1dImV/SY0vs+7B6HVCTzzkKvLL3rqzEBQymY5AkghRWXzNJ5Iz/xizwt9
hv7CaEF63xTRLmuF5UY8xIahPo3pl2kpgWvPCAFn7twpnYOJWVrqoZfS9ZjdCeQr
6F/EpIWfZXrjzdIqfyasYOy4/U5eEHe9BLlsmdPI/fZk4pL7j5OuI122+Cg8JK3I
G2eSGxmvA3f3RC7RTJFgMnnfajw5CkPeotpXykw+YC0v3OxAp9cmLal/BSyxh0cm
5JJFKHNaUMk7i/gkKqogvsWXv98LKPHc3v3dgy9eT6elRBQR61tdxJ955wYLtTCK
JdFh9nG/cp9NF6/xzF5V7r+CYHbNQvUwWiX78TkFCOXwvzhpjiH8h6np2sxkLTz0
5vHly34y9yV2WV2iKIVC+67sU9kPaqK2bCxLXNvavr6SrMwXtMjzBX+v+Tp3fsGj
gLClQIPMyH+uaOTDd/WWjCnoOFuLLPwa2yl4p9LS2y6VjXBKlUXXqO+sz37bKW8T
SKXoJMx323LgbquiK/PTF5+vEEkmoKu2nwyKSOyiWluG4gxk2FCsQppRrXopQFn+
fz4+52CirCt1QzQGszJtnAmW0wdwe4pik5oVx1VtDQv1/Ad+9HXNZSAGlhKkrGZj
Voy/NQ+hAMHlSSHsdRduPHWIgtcFg3IzpUpfOOOBLxvPZ2djIMEXBaWyaOTI+tHS
yXv8vXW4WMH3PyRcc3KOMG8mO9Up7SqAh70anTxDTwHWIAItp/u0B8I5FgaTSHBO
ZC+q94mH8rS0zJ8SSFNQTYbANSHKE/Bm/ucf4xr9u5wIb44vvKxQmu5qktEHXt3A
Tm8UOIh2e77M2z778sL9l5zdcPk/4C9dUhgxjUcOkaZ2p1qmUZqkBsmW7AqHT3Yx
PNW+pIfob+PaqX+Uehja5kWPZepmXdK4qZzcNGe+VpBqJKe7Ebi6G3fe8q0OKkuh
x3cIBXRZMtWJno9kzgOaFviVr2zBL2I2zxcAqnAC9WMwiPg9eXvUNzg/Chb7hbkJ
R8r6hQGQYMvyum1QbPQcHnkZDu4ljHW2xtkDJH+kD41VWIMot/8pZKcftuWbE+Vg
VMCyUrbK3EeWY3Wm1aW/qQPkh9r9pn4wZOHCFZa+VNpznzXZuClFK3bQFCYnYkh7
4pGjyR9BMw/excUZBJzc/6vS+lELNr9V8DOAXoJAs1O1CK1pUMn+umDTR2inyzzn
CZWl9xOPRMie3CpNRvUF7AAZX4uu93p/07RuC28N7GqqR/Qwmv7ymqIOqyk3PGTn
NgWL1U4Om8lUH4WggrwnbSi9gO2TLIKq59NldpP+xiR6HmhpTTAf4g907ZF7Jj6o
/zfcBVqm5jz759tkPgpKD03WUjhvdB/f1/puAOU0Fbx0o1ufSZE7fygeGniRs2gc
GjQHQ4o1nDnaKslxz0ssd6xzIyq2E6drjA1+Vr9hO2mxW7xqhoi2a9eLJC5UUznw
dQrwAr5B1xJoXaH18lplg3q2qOrmyAxVTiWYlazXApNb0n+a/mcvw83hVdzXFtr4
rW6RC5by1ENagv9v+6/cmYDSNgBLyG9gzvyr5tH60tkyM+SI2u0oKhcpyLKdo12c
o7jigbkw32pPHpKAABHOCBqKIi8l22oMVW5exhhujSUVe/YV+oWY8FB3GAQfA5zF
/Th+2O9/NbkSN84aEdxkStCSGkiYgc1hTboeSIdoiD6jKk2wLqsGC6V+t82H+MHb
HKgIJvwqm5bxaZb4VCpt6ZxyRQ4og1Dp9oQkWBLsywkfPOYrGXY1Nxbo85OiXpVP
`protect END_PROTECTED
