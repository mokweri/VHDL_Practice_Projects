`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0BiKRMpIktoF2tDwtouPdqKCMsxIKhDY4zBT3CvYes8ANs6fZ2bCL7c20p96DfF
7kwhq3FHw6y59lGRTifl2oJ/4LOK5YFpWtOonTxJvGXz9jhEelvSr4+Kr+1TOm0b
RGq53r3qNN5jHSxzOb9bqMeVWgfHY+rhidmqUGQVgsKyUxwHEg9F7WjCX+R37wCB
vBiqcGgPawc74F1ZN7d4P6oTCsnTFAXIrzdHMsmDDb8AesYgGbXz6veIcRbQNSPt
GmNlm1M1kVg9VLjLNuGvRvXLJeyYtEDSVgd3SXOCFBTiVLqzCe3ztjXKAoqV+RZW
HxGhnKQ4XWABSCfon+igSublbG82RRo2nD5yHWHaXeMua50yuzvVEwOqatQ5TcII
RxrAXP/U8kSZsQq5zxMP5EZPp6kp0xequURfbu3pNgzo+cvXP0O4n7hTK5Riq4UN
qTt2wBL79feTqssbILp3Yk0tkWq7rXCj+oaYGj3uhx+0i1+GMj4tllN8Bt1PB7Oo
zeNEwjedt8AjfuJAgdKZ5WAtxj4CIt0BBQRs9+cY6S0nIthpfnYYsy3bE90Wp80k
hxOCN9lTDufEh6yxTrnCqmxPBh05Xy7fr4Tkb8Oeu7//SHtf7qOdvYaIFS9/mMca
yReTNbqVsA3FTtf46PYWGy8tfMV0btqVh5syo3VcHTWdv3rnmAruDnps/xPf1fc8
9m5MTDAINTJ2bbf2Erd3rGTJLE53nuD1Plbglcy0GyPZcE8sCDGOFwiCVgp2hxyU
eLCsH9WGPVkirDKrkyZaAgNAe9c285rig7dAj9efvV6kj4MqQ8mjFeKTx5mNd4yG
gykig7/MF0aHAg1RStqISZqkHi113tEHURBE4X9cyqAdSvZx8KdULH2wvJd2TS3J
MgSlcFbvA5rbrjDOaC9wc79jBV2T8f8u4Er50TCB/sk1x/xQpJEnXjzhUpCbnCH4
CXMd0MgLIAYDkl4nZEPhR58peoZF6bZgKovtBSm0hHzE0YK7fL1+Qx4eAl+N0HDZ
yKiFoBIzJHZxDOsqFZk++fXky8hlcCdAEjgi/FAj1uEZZrcm7e4e9W9NlRHqnOVE
ZdAbTNkLVK2af2KLM6ORDHjD7ujATsIU2MEh9ingGGG6S/m8S/3EKmG0N/SJFYqt
0ElIUF2PwQreTEJeIP4ct6qVsfj+JtznFD69WDK/DEYzTCRuiWVMYr8ZMYVc1HUU
YW2eHwniLWz/U8/dsXrP4kgryUkFaWHtKii6cJW40tuKQXrin95uTXuvZS+SA5Dk
MGoE9lwTQuiBHch3rtA3gIoqidpvWTRU0IVU0A1F8AYcRbHg6QfcucKX1ceuQ3bj
icf8ZCJRm8nnahfJNADbQWB2+ZIB7ubUWTCHKUni6hKbDGNph6e3ZleGOM4uSXCg
/L9MX+cYWtoZ7jFShBVjrk2zWacLkpCsDcZA7DRiRhIT+zd06Ibr2Rg83LyUnURP
DAdykOfkbNmQagPy7id5ncYGxch5YfeF9kaXwWqZRr+nubf7AK3A2ERUjdhON0UN
1fPJkMghKZVQ/qY3idvc6T9xOhKuVfUr/gKCTT5pno8is2qR0OVLEi/DWzlRERAq
dtsovgSP8h/gLmd4f6Fw7gfxceI1USpKqdEa6r/hqaEb6OOR4zU782mzFYHOz/2D
dytGOUSKQA9XGC1IlRlAAI1j1z+nw4NNhuEjEzSiFApEE6ZqyRUDln+P3Ru6Eo0c
wxvXXHii80T3x7G9fw1jZZ/S8DOxixZ6skRk0gAECG+nASHicu221nFjKALRoLrq
`protect END_PROTECTED
