`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7b5KllH2uuamcmZxwMSX80057/KiVeEMxrfMQb+dDP/DK9ACZxH3Flu3GDgcfDAP
28EM1NQA92xGIohyxZAHdEYAl7N6ebMJxPad7O8VrckTlvmYfTuUfr83RCDJl0Wd
RSJHiQbsXSDDNluxOhFED4HfY2gYHNJ0ulZbprmHiKlQsB4zd6s2Q7xvdM0K+MQ6
D9Im6x29bOvy0+PD6WGr1BAs48t6T4e2U4fGFQc6QYA6wMX1IlhwnDpAsCcoYtwV
E2strBp7jm46BliTvcT7bKPo0Kfpj6NA8AHxdHyOE2/VjGdDtqjwzz2/v1hvoKdk
NiTXFk9bImzslBRRamlh5HPhh+bkUO9JcomuC2pIqbhX0MeaalfKR02eAnFnJRsB
FdEhx4vt/V6CzBPRkAChQnPC/5gzsZryKAOoD1zKPX8wjvjB7LvH6mo5gKR3u301
0dJUmyC0Bt6kF2JlawlkGziVuibiewbPk+vlk5JKp49TaKT/zGiloXd+30wFjDbh
ozAIsC/Gf/bEu677necB+eT16gIyxVyWpKMHkGHDlVIEObL3/1hcqhFTdyW00kIa
WO2rdtv3Wy4Nji8e5aZNkZXJOwXwc78g2QTBqAN/w+NmXsj3487wahdoUviPa7K6
fEHIvE9KeJtnZw+EVxiKFsgBMFrckho57sGO6zPuJC3chYhihJyCGMhmZi8XNRDw
E+/+Yb6qu9EKDWqKH7AhfoSFWjsoRb2/OhWQYDldIv/1JDeOaGEDVFElt7vkNb9p
JEaED3HRlddVtJbnBjksQoQ6jhPKgTKl+HfdV4z0JZJWYE+t9ewO8E0xT27QNCGe
j4KmjqASqtT8M/1xQxim10OmciKkctCTkvmKmRP25+w4TQbKrpKgHVHxScnPdBEZ
Y1X24tEIuqvkUMnVkjAmwuGH/UZuF4O+weNFnAyiqbuQAhn5kWEEdNoXm7wZ5sI2
sezSRggpjqXr81n8HUvJzud89blsvIPIJX5laNiCOQIMqjs3aY/SojrrRnef7vCU
bl65KmNc8PmzFkPIh299jO05JwU3ITSkwuhDz+UvgadsV+/qZbzzHaSqXadAtTTr
zkxUttfUZJyRU7N89I/pihF+/nXE4wNIjv4VbyWw5BOXvBvZZgOGa8iGRQ2lBpRD
oBjxauoh3rILC1uXDxMm2bKXy3CetH3mORcsQCj9FnLaUIcFKHpewnG7TN7y8eNv
yUvp+H5tWhYNF0+PFBTuFSXRB8KZFtL1vIgqF6j4wjuL0ALcuObDuuC6oGNpKJhN
EUgjvZGQbCfy9T2SCDOq9UBb1B8kZdY+ghtqxQ6rn0zKDBUJTS1+P8YTue9rbMzq
1d4WnrJJXG1C7CBwdK8CSUmhqFPRSJmBpVOEionCLpsisg6AylfymlWC5z/5SMCU
kTgec33rLAKuu3lIEu1l1cWH0QDDdZUZ9eGuJSN4l1/2SSNRboDqBlwtSqZEjSF2
6a/Ni/qnVWu2TW1fkLowX6HX/1acnZ3Xh53EnnUvTyXpktgMjt/QkNzuOg+UYoQf
431QYF1DpARM1dgqpcANHc+wYHqAbM86LDFM8piJdXz0h3pJeeMdvEJB352sY/rz
n7bcWU61n/rkzT8qOKI2kcrfT6hGs9fq7XeoSWZRSWxbiDsVXQvzCetF8PHnOgQy
vCxFrknrr3aOKDQCFbrGpivK2ES+XeRNkYFsH9/bsNjiSiNq19GtL3WaSvimIKD1
GnvxaBcAgIIn+C4cppYwlvBwdoD8OuIQSslsf5dZBAWdu2HEw5t8B94U4Mo35vjY
qbJJDPLuaU0JNPr9PQyS/nmLiJG84fzJ6l3ZLTjBpVL5AcwhzNHH116GV0B2GPEI
cT0fcetphCK2cT9PTysQcTt1PwTxEeYS9vooJgHuZ8xLKyrPs1KdBjyhqnLmgVRs
kiGhuWHAXWcdUZbNFQhUPgw92HcVePl62JmVl6YexHfLkUeyHrbJvI/NYfD5Uj6g
BRPW7UJqDA7JaZIjnUpwtExzU89c4lVnP0SAtdKRseX1VOmzTif+8TlMG3P4ugvp
OTirZ6UKFQ5Jp/k7giLvP9pfVOrWuMIQOLvE4a4aFqo87zZuzKg8E07YKBhQy/BI
G9fW6809U1L5Vc7Jv/gEuPUwHwqxfE6z540F2AJCI9EvA2o732IqkgUAfpMoQ03q
d+zdeN3CcYTLiRwU46Hwvt+EKNxYZi3lplBIZ/Ix0GZy8H0p3jE90gAzcl5j7ACH
eUBneDqQYU/zAiinvtGI7/g1nlhewdW0nE+sCBzvvXKe3068eVwmfmdHAU7LpLCM
BLOKoidTG6uRDXX9mCMT9Yx+eiiBQpYSPK5sl4JtD1QGH1ArQKnGPgKZP226iiCr
4Y1Is2S840g+PCSu2wWJNA6LQPw7saIv+K6dO+dQurdbN6qbDj6lGpmcS8JQHWXF
tZLInKboWcj0LmxlU4qNr3J7Zp70uEt0XKOrdyNHxbIoo64LsJ+pWBJcgH3qjPwg
sIvj38jMcAhogfE6aNpyw5JPv8v6/PeIhZahEDLRrdnhknDg7i2x8g8iNfK+NsGX
7KG9VAk/UqnCCKStOZh6sqbgpI1yoDoaJd4qqopKU1zkUc4u+z1nqjKQyjqgJ+eF
SsE1nsumtyYZzq1rmUdl915YDIe1H6PSZFbJmde4lW19Mk9FohTdz0Te74pYf0/9
r44hGqDN5B2CWGfpxtwI9OXKlpxUMJLjvWCngsr27I+gdLqO8AUXPypkARoMgKuF
sUmx0kEatjZd/GP5mEOrkJ10BRfnPkg87a4dJYhJQgqZzptuPMELXWcie1/bM7eu
WEVmBrz6P7wqOIbaknui8eVl/1aXg7pkrfnkEj5TIDodYUGNlczqOp090iQ5iDS0
JvJ+luHeQVuiIfMl9wuDqTVw70NbB5B1SYkynwPGdcbG7Ar1CdZklEceb/uwwx0g
9xRe9dH/awBY3TxYjrgCZXVTSuPLVzWgqCo4Z7NLFnqAJmaW5vOiegZVX5FYwI2/
Px72AGzZISDm9k7xalTF7S1K+jLK/1037f+drlvuLyRym0neiUwTTxNFOi3lFLkS
A+vUrFyVxlepbIca0yfWSgrYQ95ALW5h9UxBcdZ7EW6CgDUnu9cPg9o1jlrLoUJH
JQZLxfU/yvGYuXrQDbHnqzPNP58JIWhuf/uM7pz5kJqjB4qjQK8+uWMsw7XerPTp
X3/1iF8a9fPdumXNpcHgLGam3xwzM7m4rPJGiXJaMUBdLvEZ72VjopnWBy2V2ce4
FoYxXcPHI4wmmZlEdU7BEH95fG1SyCif3s+R2Puz5xXjJUb1cSiHQXex8frJu/jA
CYkGePCz1RXWlOixO1j7sAqfilv78bh9X4sMmfZeYYDEMHfLJx7LLO3HkoxG1n53
xlaEvq14KkqntyqfyWz3IskTHy/Ln+pvBBtj2iU5EaGSUwrgWh4k8LLx8vNKZF5Z
l6pOMr1x8ybXxyo9RS9DedbBwpWJFZRd4qvuntQWbKX6KQbe29yc1vgIoGiJBi0O
7eoRXefY5UmgHre6qeo24JVYoqGS5ttmYkev1bpr2TIAXSMMjpjC5cUUaKx3WSQQ
XWd7UIGqaIyvhSSpB+ayYax2//9I6wI3OFUe3/2T9Yu4ZUmUpbB8106tvOdWWsRg
bxmAncVQvjCevWWcoSORbSht427LxPVZYdJW1JAlXBSfqKdqzgjK54D9K97brGV1
2QcD4dK6qEWV+79wr3ZMhsw6An4RWRehN2yVcoQ7+DE2WPmRe2dDuIk6xOuBoZWU
ez2KEcuCsXehTYFRFEi0N+vrGFhXrs4JNOvCnzrTC3/Ctd64rP5rMDBYq7Bk9V/5
YI/pPoB9TusRRiCnufjdMxsFKdODHPBTkAThpYTFUJ9XsiLQKx8XAnpOTJibb870
H1XWaLARWi4DaDa+xoHloPhItkwMJUhdZYOKl+3P9A4bDZGZvh04GqJtRlJzUEX/
dZzsgY8xTo/QIkOJHrtHkwPrBSEC3vRt/Q9OFxRV8lMz7N0jO4zFUC496cTK1IaP
h7VmICipZUzgdyiYp41HS6upalul8K3z4Hqg9uwFrBY2QnsSpnDX1amsNITOiHpy
wF6p0bv9f2wNkUAJUwnl2/ap1Mcrz1dAJfGC43OKdu787QinhCiUppC93QBZA6r8
wNSAxhH/kGgW/wl96NYvmhKxndmPsvZYzB+gmL267x2hLmEFTlH3x8ruRSMR+E/Y
ow+lwxTteZamyz15dOng0nbksSTENZq1XC0ug0F21LODqxwZpn5tFPCTuIPmykZp
5cjpVzMnOQBJrdZtg1uYLU7A0ja804G+48vQ0VsPO+NnF0/RqXwpOMqb0wgEEMbm
nl8f0GqH4Skwfb4o92Q9N5djB8OBPzRxZHnQVJEvq/gnkmYJlTPVjEAUGcfy3H7C
k9ZpKXVCy7wTJVNHGdA6JBaMTiPEuNU7hSZZaX7Xx4IaR0MCiOZgFaWR+7O10he5
rg6o5mulo3kEiBwHJSKLcIPP3ZKy+T8AImeZ1U921Rjbb/IMn7Q7b0quES7LqsHc
joUHulyqWdGpnqxrYvduNNZv8yP5a/Lz/DEy9ULluY2YXRxPzVU1UiikFwFqe5Wx
gjGJvC4vnqS2i/KC8PNZ3VlGATqFYI1Tdc/VNn+ISDozsc5Uzo1pJgzbdAdHvR2b
7xwpZ2mvhbtc+FQCqJ6S1XKhdS2T+oPEz9p2+b9A1CCZNB/cBgE1z40SPRIqT45i
M9AASYez1nbxTw736ZYJtejBdMxZs7XVRKLADHHzw+h53YcUXCSDL3nhVYpKIPb6
ob7w44BGRpbP1kmdZTlpPdFGfqdP1I1p5Od239CGTBoxvAY2fDnJaLD2KAt9XbwI
itmZlLDh+4e29w4+5BZELbOHLs0FK3i5U2QijqHygihcsygUIzsrP5VlMPCBAkGz
oqwUkcL14ShcmyA/bSoLhcolVF6G1F2xVqvMatNjf/En55R1GW8tm0U5ko+cu+Xb
q37uh8zptOAfg4VVQFKj56G4QaKOvOt0jSPsU1piXn7gPOH2RlAChJcqohPZYbm8
QfsSQt0s+eGdhF4erIzceJfwkNSk3U2NtTS5SzKkSOdSpiufpZrUCzo3isomq30V
J3c3Xv6VgJo8U2pZf9MkV+5nb7cg4g3Q9p6ahGvolACUD9c1TSRoMGig4AvFrP6/
l9JAOsttfCwXzpExdwvVP8u/ALQzFLYMzEZnQJesHTJJ6djLu09Hkdrckpf13e/c
ln6VtPIdKr5E0hKnXvfWbGXd6gGo725xDWsCd0Z4nuYtxmN1Xx5koREVirwfk9AE
LtcFIK+OOPmHd8gYJg+P1LO5ZGqLGMh/77MyPW4EijSPH6mrvFuTSEvlvnWZLCXi
DFz3KHRSzu9nicHUnPulslXw9PgdDJMpAguZS7EW9McHy15Zt+aqXsnHD+S/pEH7
H1LIeXcYZptqwjeHQI0oUxoG0FIzVY0PcZM2vdb/U+liSac0pqcWLVb91xtA4gEg
26PPHF2f76J2jLBQOLd/HJvvrLdYM70oSID1jDcoQ6RslNjjV398AR55SwgC+emH
Pr88MqexqOLVe6o71OUBetdlPUlb3unjHWTeFl/fDg2//RUVuuOoAfiMpbVqX89h
Ykh2UDqjoY3YjLqv4j0vtX7+eexpdjHwVl9ABXcqbDkduPGGf9H39WjQQtRkNKS/
i3DoA66vtbCs/Kze+PV070XMVv5u3OfHoJiqY464aKEbuOwYvk6hR2hGkUdtmqpf
LNCkwYW2qdL4t92H/7CakpIJaUhvo+weHLxSURtQx9t1bB9DldwDySM7978t9zp5
AL13hrLzKhxZuxMvg0jpV2RF4B24VmUAr0jjTyDjXYWxwhV2lQeEx2h7m8aPKMRr
5D3MceXhbSx3QLrYI09oRRppHZKRrCCU+shcJg5vBdCimEarZP1gG3dkK6TRVlF6
I0xrGou3G48pszm/f4LhNLZp3iCzwXv0NRAy5/UfqAuNWQVnZzcZSsC8fvmhgnBS
U+LWHgvTX+ItQ1AbOLL2EVQSJ1oeqxS3IZgLNmnijLHppgTw0j2r3SaOhiuen3D0
awm4GKY4zj8GK4tWhEtzjWqr8uQZ0vh33t3HHRDi3aWkkFWfOukKmvvkEaxCTl7N
olKA/ljWDA6WrK2+SlOtBY68fS+gBuTuGL6VLpzyV60aNcLR9+f05Ggpbwz2gLcS
NE6XcZ3/JgtsBVAWLRr59VCuLLANd2j8TnMC3x8a84YvpCIvRbUGOvcJQgn/MORN
P/iDfzKZaSZdcGTmhcVGDC1PUvdorpYDCU0a2j1+QZOT8vZ9a3cPjaIIfX+JIVyc
8Ew93CzcwNXxfuXzMm7QKRf/UHrZNkE1CoP7UX8kaWU35nuP1CNm8PTmENTzI8Cu
CXqXbydvZsKzwDYAk23H9ZYgMlUWSZB3yzIwU7kDsQkO0N7ZFop5ojCEyuofHnF9
eetO0S4iSCHdCF8nVpDkwBx13TjhQ8+wpDQ6RyFKr7/NuS3FzdblY6Pglv2kMUeV
uhYkvUreqU5DuFNak0o8TMvcTa5cuv8H/ZscuiFDmrhpsNJacAR4GkVH+B70vR47
rKjxyLJEXSHsFG/QKcv5T5DUtUFJMFz9Qsdw/ifRlyzoTLip2yV7imHBJ3+2W4k+
`protect END_PROTECTED
