`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFGI075utY/rCEs5VhXPjlq+qsYZ8+3CYpLKGRJHifuWUSP3htnSJclr5ZdD1VC9
Sim85EvL6pKNUh2hgru6Wax7ceMVaiyWAMkhUoBHjpgRdgsw2wMrfZ793fx4YBT8
lTzCNIt/RtxgTPnmXcZPbTAdMj7uzH60gHg1x2/m6DEL4qOpfHJ89ZkIhL2JP7YW
eqzlvbI+ELJf190YX0N7mEPAl38GZzI5NEbgLmJb134YbFSpe7DIbUNaMvdDr193
WMj7lj1TQ+QlA4u4oXkDPKU6w70wCHLA1sHSZFOUceZxjPQeEYa92fKvr4HvH4ZA
xw9ibCAi0QgMCyYoV1FN2K+azZut3pi+K2vqpeyBwlRCn1ZadWuW/WSD3uKrQXdI
NCavkQAugwEuljoU8X0rEC9sjT9HNZeE2l/G5kFLgWhUf+ODZ7yLl0mAbF2ZHOYN
nVUUbQE+0GEM6lqbsL4LgrNXFu8qv8U3T3JxQvxTc2v6/468Td5x85Jq1rplGhj5
GQxCxLpsAzqDLbkf0CgurAZfhoPlzvZRX4CV9ddzx4f3tWPk0x06CGINEZ72M53l
tkChGaq/auaEb5snOO3yQcUwefRVIycWbutCoGKEHHC1TdpbQlOUwbfGIQnidwLx
`protect END_PROTECTED
