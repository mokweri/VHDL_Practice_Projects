`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VOyFC2GwUTmbuNmI+puKOFHsuk3lGgMWT7gnxzOmODOafupq2THFes+LB2S6mf1u
fIz5ouo7yTehaF8EwRP9Ml0JOLw04vJNWt+136KRR5iQ/qsvEKhGruLPuFQ1SBeK
tLWF/eo/5teoefqKpHxpM3jwETkQgwX/K5lINgESNUeZ5r9Jl52R5YjwBo+9h5cD
yisYe2Jz9594Ku4KiWn1GK8bsujLSFV+2rWaVZdhdJqItw0zllnAWn/Ao3YN0vLA
mVyMiOjoPOF1n2yy1TfE8i5M95Njh3ndcb2ewjyjsbf+YZs4hKc4FmNgdBiwMW0/
07bglk49QHCgNmI0bHe0++bs6JI4iTl5Ms4nFaKYYYU/2VekwvCrjPiEa7iqZBhk
wxz1Tq49oa1MqHIGAoXYO+7u8g7uK0HX9RLQGU03X/QsKRJnQoqWI248nXxxoKWZ
imGiqu8F1KR3A2qA3l3nYh1Vs08wukCmMOxNPDJfNV2j7ngx2PzQ8Jls7AOBeHks
RDJ/jyyFJaJ9/B7YOix2UJgiE43hq5JbW/joT36OLHijgnC1gnEuh4FUb1rBFqhD
MGxOycsXl1VTZUUvdHZkKU7Ratzpy7WzRgTnFTb9DCuJ3hdYYz3f2RicDRXbf2am
3HusnmdN82M3dMw15ioT4Q==
`protect END_PROTECTED
