`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRNQNH8qcxWn3JCYLaEwy6VgQmvLjYsY394rcDPox0HKXQFCokkG38kIZCKJSqIN
GSbNm1/XxLfiDiNa60nXy9SV5wIn25pWPxUzVM5CMuhmyluumpMskfZ3qWj/40ub
cSB4AJVIkMf/JqUIZP5ipbUczA9CL59zkSR0xF30SVNKykZHnTTib5zE3H98K9lh
Q0tBlpHs7N/xknWQF0nDRMTXtPyDy55CpSk9PT9MesbTYm5ZqN9QpRLgjURW3ytB
5YKzGPWBiffMpNQQQFVlI+T0c7mjAE2v+QoG4tlwXRlTjZdjSSYZqmvgu1b4nclc
4mFjYcMaAB2mP9Z5g7MH6ix2Hjot4aYhiNVdI3GwGtRjMBwqKUgNaQwpe8aEUuJn
usj2qtXFumPh4FeUycWX4BDxb3eRoDjJOyow9tMuvYEWftPhSp70ADfb2hSl9yy3
0qOC+501D0Go2cYYoAbII4rmHD0RCDtAxd+ADmEF2w2XEbedtAscKylveCrzGxtG
IgUxyrawVK24IH0vS5AW74ysAMLIQ6sdN5/qn0EL4M+AdpC2uzu6+GOUqDtZwaIP
rrc4R+lg7eiJg9vDl0v6LBkR+0NhyGk2E/znxlR/xJUmI2pnqOsrnejIA405i/Qo
Y7vut3HoFcVRzxRwhAj8jEMWfeCJvDugBKmuW6aaaUnmqONujME9M5jGjUbb3dxG
ObQ3SkyzbQ5PaZRkCm4KOxBh0qxj8/+Bi90AwC8fmJM0FP9+emdkHwX8lHwaatvE
1Frk3q7c8Mm74TuuX1grCn1kyGig2jdHLoutlDLHSxp5UM8L3RLIxWEBcc8fD4T0
Pkn1Pn6JiAx2lB6PDeHaR/0x3ZSPpCQErCIiHsK6Ne+ttIhwGIn364dMZoNEP5ZH
ggzm71jxeA1Q74J8Yp3AHCnPDPwNtye03vRmV3M6a0FVZ9AjXA0JYHykY+Wg+XVE
TXZTrY/CgEPpzDrCL1J6yI3soPXhqPoLktUHCiDmLQXPLhSUPWWkD+E0Y1PeEqOY
FAcF1530I69Gj8NND1R3odj7JjAOiaDYhMcJhH+fUnT3DdWyKzXg1fVtN0K9WoYR
97IJ515s0x720fU6cvkliGqXmGbb8JypeH12uY8j6lPa1pdtlTYFWLJ0cWfbS4aJ
l0g52Bd+3m4fh6w8ErWpwA==
`protect END_PROTECTED
