`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vs7PbDJ/CTfgnqxtCgfIWjV2A31pNSXpCQqAOBAZ1ah4VxMZr4hAU/Gf9S2nL4q6
oLcOnkZFhbTfBJsxm6F2eMTjRSZg+g5+AUUEv4VIsnydWsHx/coieFaCXINms/vk
hGnbb3tmsUT+UWELuHtrkF4cwjczSzdedY1eR4xcEx/Yz3t95wtwZZaowzU+iNal
ErXmtN86pgrsvHVHUISe4HdleFgGZIQzxIJ7ULU+uhzOVS4qIhBhWUJmd6MeVz45
kxn8KlfL/UEus3vSQA9v6SZB+AB7rztspYTWM0mlZsoY7zTdCDbSsCZIHbfhmg27
JnmdnBgDo9ejvtYfm9NMUDx8vWlJ+qwJfOfOJh52mr+q28Cte/H3Yd03feds9qO2
XiEI6Prk+3jjyMNxOV5QxnfwROqySvy/N4V8FbJoze84D5rzBHRpV7RGUy0CEDbp
aS4x6IEdySNtfZ9vHS5v9L6bVjStJsEEqWn3JEz7sfk=
`protect END_PROTECTED
