`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5ojSAXABTxMtidpWzBGnc5ItWl/l8vCY7nvjilSqJtneg8OdHpvz3dxKot68nGp
ercejCLO/1vUw3+0X0htKGw4pB7yczNZcj7U65xdv10Pp+6iN0wSchBR9nST3Se+
eRgOQbLFMgSM0T3ydcT3SJOKtB/wHJgYkIznTA8u/+ySLgbe6n3lIicR9wEeiMlw
vEZ1KR2mQ/sC8riKCx1YvjeBTL5CNLydLuIP0VpAKEKnsP7DppVESRc4PW5Ix8So
VyZ32voYUAIBh3TFboOeVqhyEEN2dN3Qgr9ghT9E8mFWbHn39Lah79fDn9w28Fqf
t7uGYCkmD8UkQmLGqSYpUPshuCsgoVuY2ajUALDaw8sKOlmMt9YYhEkmr+3UvWOs
dltFlPOpQ1L/JjQETLUyydYbPDcKN/h30Z2b1LNb+XdLVd70GtiXZyiByUI6C7th
brUvq/sOovqLpieV11hHhtg35mYzqCKURMWcqKYcw8X6PIH6Q2ukvfWN+DqGbq1a
a1E49IVsRiMSop/cKL9+iJtH8+UuOVgXfqBp1LZg4gdY8NUGFc9PPaScBLa9+7fX
`protect END_PROTECTED
