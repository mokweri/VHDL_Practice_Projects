`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N3ZDK3TOjUlepieypSS/6xiKzQUe4UlLJXhtGcKNNMipu8x+IJg8bHXIA6OIUTJ6
EQcb2/hnF7deC5b+8H8DAGUCA3OMo163NgJL3X6kmWBuleJln/mdMA42Y5A7gkY4
9n/YFMLjKoS87rSPqBtbpFC37huWSmYV+NDBtjAbh+pgTnycO7AG7cyOhQ/gcZT8
nodVUyngHwUh8ARwb3gtyBG/Xpo47xX5JVgG+IPPeFZeNIAgOfqGdnYPrtLdC3Y0
LtI1GCOkp237d9kaJHBS64HVQ0sD7dm/Wyo1PQj88jg8ecyLRdGZg58b7FqV2z5r
C5mPSVatBRiUw4Kb5Vv2VZE/ZtBl2t7tEJXFgut8byO6879MH5NKD2NaKAEM6efF
KQg/W1GDEeNJHLj1hEId8EGjk1u2KtloaoOWmFHUsUb9a1SFWZl91sdP2tpofFxi
O4T+WMKA6I30bsp0yVUAbRLBEsO3VNHmlOAxJDLlfc4kwc+1Rxgp5q94khwGnG2z
7qfgKcKwdX7cagrRbWPXmIT0BBc134p4noRaXZdfoQ9rW0vrUmFcXITz0fGsJtX5
iwCS0wQfwzdR+G7F/BQWlqkS/ZL726v6pYu3BsM+416dHCuF24XoLnSSWqtnP6HB
jL9EpDxC7UqfyN1UdR0Sws5d3T3trA1p/mJoTwcqL+0gvu+s8CVRmklTL2WxNWeF
aBORy/kpChXe/1bpWCHwDxDX3/S9s6E8DFShgIxPb5oyLWcmW/CS+ZCpA+0YGUXX
F9fKoxKgysVQZ8jNTz14tUqYIgYgVi5idQLrao4Ps6azWVpV+xRJi0o/GnZpI8Xp
FqqEurRuAwaf74Hkpltpu5EPHkRe45YFnoSmJZIdpZz94ILmztInhWZ/lQzzVjFN
4IfnTjjJ/qFL/xgKOpasayXO59FKwO6Z98/Aw7SxVz6xQu7rFDFvbweC5dm6Di7i
/kdt9JgA4uf25A7V13hiP4dnaTAPjimQScEl0IwNjsYHGh0/pB9qyjihk39NM9GB
tNHZbgIobzgg8GcHRfDa00yGgi4R+EbXAnAqSjMapN1aGQRiuONsqHvp/Cxx8q9e
dXQ2OiJKwIyVsn4rnJaPLJRgmGL5VLJmADrjHNYkjLxQ+p+Dn9jUxv7EWA7eOArs
prrewjto3GWl2/+Jzi8dPF7S8dHQQYtfMMHMkAdxPRSbhS0NKaVYe9owhsV1y1u2
rIqzSJ59ksxhHEzzGFqx2Snxq8WvPbRd7CuUQTGCpgjbsjGvnC1nh4ypUwQzeR2V
Ctlz9iswU8T1wPDKU+X7HCIEfFYfo0MTSoY865hEapEsOqJ4jZdd6NW07+6qT8Eu
hZYLvy1IWT/shAXs4ILDKo76Ur+4vzzbLSZykRVE0O8FkM/hWssFkNoEprtTu335
jlzxoRCmQl0kWoJbF5u73dSMA8FL8tW9hYqdeDommDxdjngNhbMWznGNNIAtfyGg
iUdljl8dKSsQPA/+3XMrYadnM07xRuACAzTqEEFVcsGeDw2PNBIvvkj9b9JZjxea
ElDs8PVycMBITou3fjHQfzzEqwGMvKz6rO8Isdwy8phtbTE+3kA7yuNLQEb7wlvE
7b2hrfAd9ojzTqazXF8OLP4smcG0csL+/hdMKD3DienPYw1ExR8tqJoWHcW3bHqE
OlXTJvcMUyLGWedCv28Acm+VryUvunyssBmx9RcvdE6vIIeGfxG1Nz+wqACreNxP
cxLNb1MBd9Sxydt8/bTK0M/UGo88dALJDSaBX7jkl3LPTWqGomKVDtj1lECXCZK9
qafnI8aTWwWIAaASow3Qt8/yI2hGXyuJwA5Bq6KVTlSUHLJADQEthjzoxc1h9t7s
pUQ1Wbo1ej6J3op9sxXyHW8kmnCyLn6zk/XQGq1M+YVgqJjk73KPbU/hv+5ChIUh
dKmdxSjupb4gKnHOJ12e3JHXiHtW1M4VBEdFclvk/Zu0JSXNVyu+bkD9y1LXz5Nz
U2TPTTVkvohNM1FcpYOEDLM9rDKG7pN2v0jOL3HbDqLjWsGF49p6DrbCWm/SP6Z2
TG2tzWXFQSNBQw0FeJ+FJ4fCKnmcSjHh1BDb+BI26pKCIxEjnU934DyalmcxUuMP
vWDsXJGmAnOpAca3LUuyuwIRF0zxCKi1D44CKTx27lnY8M2x5uJBrYpuHzxHlPpQ
lllQkZvxkfqRDXxBlY2IqonE5yfjh5H2V4aP3GkGIchiS2DhQNfWeK0CyvT/W8io
6/2EN1hCiAw+Yco2aQS8m5uzFmpLiy50XoiS/YX/VedkSQm0fiETstgFJnDaCTdt
zKLHEfb5aAlTw+dsS02UyiUgOwrqr/G2rpU8OKOGGRy0tnVamqoHln0yUzwg30cR
u2MHI+koTHNrzUCuhrJBc7v3I+Hm4hFM6jL3glz26kRoKqOwh8IW/hFQtbVzKuJR
V93EGH1YqFn2I1/uZj+GfCjnxYwcSLmc1q+liQ88RmnuVEp80RKapHAmVs6XbogV
Iw3N3my9QIbb540NpVw0RYl6wJ8kRJcilGqfNFlPtWtATpIlVg1URrUnMml/alCc
EAwSCXkL76ioTAxsP8ltDsCwXmMP8gqPhOHNTqiZlcbKmQ3dzrJgV5SMPDdumfCw
9yoSqxnejb0wPUgyxkIifXfxEt9MjSIWer4khpjGrQVk6cz4s3VhVrFrFk56B2JJ
OFRp5LQmbl8wr49qJQqQA8Pmm/fgZXexwU+SjXcw47zp/+TlOfi7cy+9Qi7hFXCM
nUtDvMGPHPcG+WcPHgIKOAaJoiQFdAF0tGai40N/UxOzs1oPj4ACagTAtzPk8wcI
8NSvyI18uwo09SIfTRrBeI4x6e8WFZq1MoUqAMe3LokVmJWhXc7k3M164f4fBl/8
dgBC/ZwWzUPTTgmUTRcVHqiZM1PnpGUgKzqlKniH3qIxFu0JSPLAPapQkTq6iv1U
2fuBdtWOZ3oG2WwClsk8WpgsR+GAbF52c+8uZE4dAfithJ76hlN9VHgSoNxurMc7
0n1AiBc/oZFTW0ti+7MU9TnWGK4QL1zv2RoH1vL4sOyuowyKybgqjP2nQlmA9WlL
mXw0FkrLWPDQk+dZWM8sxTxMbduu8HY+djYiHZZi5H+JnRKyLCZFtXy+Zdo24T9H
DyheRLt5PwGblceT0WxHu4xlaz/+CBqO30JZ+N7x/T/2WAMphSrF0cVodxVf6ILL
O2+av8Qi60GZPl2bXHmnRU8DBr618us+XSRjB/FRhon08Iur0o+lXfE+bMF5SxQ0
SDXolfhNoW5AKq8nH3xXlfjBvbU72m79PsfU7E6VhsUwQlU6r1DbRgcga3kjXgNq
xxfhaKi1Jx/hjq8bMI4olGkPwOg1D/4o7AoxFt27LBwWddE4ZftFD8CfG7DJ7jiT
`protect END_PROTECTED
