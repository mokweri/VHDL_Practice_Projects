`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MJbpvqcRyi3Q0gig/V1o++txEGjy6xuJpdA8CVGeHkbkm10O3iw2vkgej4vFVPX1
Ug/Dxiu+NFUK9SOzxABeg4Ky8e74IF/lemItlmpXULjr/KZhOK5BGVacLu1WeYyt
/Guea2XkGUVacoCkuOgt4HFvwJKXHrnllPLnVoZ6RFdiNIDKrlea3HWEKkM7yS0u
UGM8sRcXfWKt7+y+gp+1UAdKbE3+5cqZvAp8sbmaYehPv6At7wfLtm3CaSGJkCVx
R9umVrJgWuwOCwSaK9QZxwgJeE5saUpmSTXhipAYMB+URmMB45JLb5rJFHqbExZd
J4nHoGlF0dONvjT1ryOiKUqoXZz1TEBfbIzrlnN9aOCrUhPXs6Euhsb4xkjT4ZMj
tE2mnAjIai2xxnfPygnlyG7HYC8p51RggsqAmI2ysFzLXp0VcN2Rzb1JFgxAWeTp
x56GCyVBHuuP0djBY6vQsDd+WAFL0BT3AAPMNfhFAVI72gzW2FKhs5NVrGZ+C7J2
y3M9tnuw0N/fmIKlecxJpZbibgkKXmCNvrcmBv7vM4gh3f9tZc61tepiW6cCTwfO
RoiYCg+3kxKtlJ3q198hnFw9g86VEiZR1X3llb6CQ22WH7F8dULIkkX1wjn3TmoF
NzxCYqmi7FRLmOTVYjsxd94mMUzMVbagynwW6CH49DNJigdokDZbrCxlcBbdQ3lY
fOAt02+29EOE90J23jNbp5BHwNb8g1V4C+roXDpSQwy6B4FHlzRsgqgijms3Q2Wo
GpHCYVdKb1ZRnXdVqWOVPFdgbYKOrnbQH412cMazRj+FjMSvuTJYgAWNcNWPzJ9+
wVEwBzR8WI6fgK8c3iHCD8CA5IQL0Hbwe6oufExdv95TfeUVBgOXBUT0bOGYodro
TGlwb9Zah+rAdbP/SvEj5MlKzLaQfDRCjrggDnvlsqXtXDQMMQ7g6sJVIanvQz24
PbHF6mJbRmMGJfwWKfKuCSAiEZaj1fBqlt1LtPVC92gyhSMJEby9x57Og957CWUe
A9gBvWzgkyhYbFJjHmdjJDBb4J+X2rjptCObfT4QLGvuUeBafRkF5AoKgWsBJ3Cy
/asa/IWPAWQt7NUXhUankq9tOJ6Ed2s4JIDOixTK7xNoTjsxTHMwX8Q01p2xaM1g
qwo5wB512LwggbsXdtBJOkrkIMwNe3KqS7BRwwigzNujTuPl77DBN3Vw0Qd0EhAP
OFtJZGt04yqYq9Ngs1JovK+VUOURpRo4pKnUT+MpHX50pes/EwWba/v14Ue4R39q
ue0VB0aRs4JFM5XITzZpvE0s4dXgfP6H1qdh4rOSuL1ZcHwg1DB7TVh+vMeBT5Wu
pVxwDfFzRbWeCq/8GThmNPYL2q2hWROZGJ+9rcGdqr8mvLuZmfO2P43JNvDxqLFl
X389l8FUc2vn3bMYcibaI/44ISyZeLVvgtPGKIB0/UWRaR1d/s6SYY7SKbfzlZ9f
HBZJX1VwES4XFsRP+LVfYXJ081mJ/wbenH6PYGRKQmGFqIczxRM2g6ovqTc+sGOJ
4yv8SSmCfaizUpCICTu1kmk2Syasl8IqueGqUpiagyP8aKJIR/Czw5szlPbhylIn
PBrwGzI/6m+UVPCAtezOCtPGln/adDf4ck9CWcp2/aBrYMtYcRtZVbzMFkf5G+sc
CxvVG0XNfdtecdbCznu9FWog95j50uV3lQKKE5q3SmRfJ//QhkuOhoqujgx0HTla
69B/YSmooBEmUd0f/tLlcSMtMb0kzr9YuYCcq2c1l1jhvi9ma/45Pd3o22KzLUwo
ZVLdU2sbmaiRMM4HpnGOL6AxeWjuBWEdbP4LDYfsUd6RdAJ3cXaDDpzu+Ic6xpqL
yz9qIADEzbM3OCGk+A4sEfwIGdiWSouMZrsyuUAVYLSeXTCBrjFu/ZlWI1VeLcdX
XRYI9HeM/+rGbXsfqcDTK5yu4P86g0JfdioHcv676WojtUTeK/ySxPpX1HYFIxh/
aSHoraktVdsvx6hTMZa8bR/eu62X6hFPLGlwS4pd94JqCWTTnxWySu73uFacBCQ/
fWcmuFpf8D8hyl0wlZ4oDl1D1SE74r0pKgagw+9mlKTU57jk9+oW3pLGfyXd5uIU
Dz8aPIurGRQZEn8tGkV/PlDxzGi0FKq6z+roHVg/4bYgE6Uo0HfO8LT5ImmLtII8
qn5XiIy6I0Tf09ZebQqZb/HFXLrw+9rbk+5YVZv3ZD1D56eQVUnYITrPdzEqupU/
6pKU7+IX0jz7mFhHxwkE8+rH/uQxl76maKiFgRzDMo67RNO+XY2+4oxiS8fUrU5c
9i4fFI/GG1nk4XmmQBEJBt2gfLW4Tuu879CShtqXa/uxJZ9GE3wS35GAIheUsK3v
rCsotx83BHZEyHyEX7T180WRkCx4zq5CX1ylHqmBL+FAAQB0ydD9OatmwQqEG6bi
WgnsYtT2J3QIR6a120aYEEFVMXFdSOk1sWZZmzDKjGLzmGOgvXbDWjmn3QH4Wlb2
NwYgDJlxEWhrt3MFo43K4b+ohC008J4V33r2zPltfZCwG14QcJTgqQWYol2JBy4F
D5ly6LSxeHwVjlWKAQygIZRyTALp7pm2AvIPh0Q93HjlDWIPg5OaDGYDOZO6jBmU
5gP9kYSux4VxDIBzEhRpz8K/ruQTQb+xDNwcesYLrZNUXARunEQOY21+9dsRQHRJ
v/g1hGjpYnxhZTgxI/prj6MFPmWUUtb8aOjEmvmBw3cJfTpsBMNKM1honbBbVEaM
yJ3/rR5ZUq2v+QD7styspCa5LCmaEZldlPesl/ckoukm4upUaNkGnV7lnTmh/TMl
Vowg9P+3E4T7BuoQbow9Z8iBJPLClf082Wn14Zy9AIKMsGXAkUjBsVvNP7ZkvCWC
j6IJeheSUg7wM+qE+JM4AM+Mpa2ZEIi4k2ImymGzNxT009YK92pcuCPIrbHXmUBZ
/zMXuRR1mtukg5DvzFqlhOTNasmWm4179wD58ioGL/cE9bXmwLbr88PqcgxJaf65
y1KJH2FhjNl79QWOadxZ4ntc3Wems7thicJiDMVWdnMRa7UxqAHTDou7m6Ud53eu
d2BM0LNLjALSFgg2/iQxazLz8WT8qQ4RiZmadZA/JWeWVF+7GvDjTCug7IU4/GUJ
XQcfTFdeIsWLbgvjYMEk+2fE81AXQ+IYlEydTiwsIHaWjE4S9/6yojtOX7KMZTwN
mo/7U0B4IXo11tejn77WRUuevJeb/N/MKYgUMgSJPNJVPWtCdAV0E6uh+UsHiKA8
z+AHQIowHzo0tXa6HPG/lFFLeu50pj1LV1rrgOQ4id5eW8gebDubiVUUEcgE+lmU
IM28EY5jLLSrj3RwlOowPYVXTlw3NuQXSZaLz/QqFYonPiF+dVFR7rrzJLIyctQk
Fk6r25aUvmkP/D43iLimdTbmpfS92kczENgZwI+VyeShss41Ik9nyx4U654m2YFg
9tmjxYqv2F58FtOgFgpcpZWYlrR517MwTECdQjT1mJkDMk4nYEpVTak7S2nPj1Pp
7eaaWZAcFiV7HiZe6LwNdYx/iLB9/NVfyRo8jCrqaY5rutdYjKwE1NfuSMAXOy5F
7ZkgzZ6my0BfQh6tzTOLfAbBiWio5gTOR/hvx6q7YPxas7O322TTfZVMsLsrwKaO
pYA7Gr+8trt2lyduGQs3Kz3GKYqF+LWvb/V42/KezC7o53TaKUAoAfPFaS5lFkWf
Mpmadnnz59GD2RHYBwSqT1Kh3gIgt+MrQGhIz/pVa1rmUbZjPYQjRe2iXvktd+E4
tcASDtYBsAaNBl+MPjYW7SvIRSudGj+PbrVrKldura9vXE+wRlNTIvjN34JYWWA6
Oc+kzMxZX+YzUTsAVhp1WcN6d2Sr2fOtAFeVRaGe8UCBFTmYRVPBPen/ksoRHg/l
qrfYrexZca0PmVFAwR5y5/6jj/0tlaFoJ/0ULu1NFIY+R//NnN8b11Tk1WhRwYCq
o2Wgjrz90q8SOPnMz/UciLMCDmN5WZeETCFMOXSa1cKjdVx86eDhtbULyKoR5nWw
J/CzrQVOCi/xRy8Duu2kceDM1V3dYou52BOl6UTPkLlpzrzxKvLZ6/JGnltNR7Xn
jxIgYbZCZlmdf4smyro75ynZWez4dHce7+vOxJo+oad5/d6xTTYu4qneNvfpQk4H
3GTRVNOFC4m4p9jPIiP4O2mo4wQeLZxAZ+8ASJcBqGiN5kadESWjqStvRRQ7zme9
YGyKrMSMYEiVgARhqadLP8FRxEUopIhP1XdtFS4EHjhUZ7M7/eaK4gXTgVHDE+JH
46BkHS4Xbzv9J3w4zO0nDnhzs9A5+9dIqvng5G9MP/yAB/8Yj/02taBroiyeT5C3
3b0/jbjT3xUccLgzvXM3uevLKUewzG8slekQhzhMdrJ7nXN1xNiu/pLR6Wejihys
vSLFOAzRtSocdR9ZHYxeug/GfND/Uun4Y2Vj3GpJscK0eFANyiMUrqhsYkwgc26H
ZopEkcU9At07FtEUyxAEReaOVNDonCEhakE0BQaz6tYIxyPoNcBZjXf4k9EJYKQS
1pEBVK0DryJiBAGE08BAFrMg0d+5u4qV4mEwV5L0nbx1FePVPZSG68FP5EETul2H
OmPm+eYrPuODxlWAXYc7rH1ybvwlA9Eu8+cOZWvGCtQfSM2rXHgXABA3AbEW9IDX
3zFD6Bythyu5dLqVeG8MyfEn1olAhmJeHx62jkDXpWxHgjVQDHv2TMU+YRCY7ouH
TRI7fS/JM2LoVeCe71g78jwo4kkX/VbLIyG2ZR5/x4ALpBAC87/YcX4xpMhPQCr6
t374AuwtQdSyAmuG2PVMGcCDPVZ5aMAAZdeK8LamSJFhYg0S9oYpJmwQIhToX4AE
Ycmqkwt+PDdjlEUmn4A1y/14WDDiTZ/lp5vjKfPEXeaXgiA/+SYYedj8kTJvYgE5
jS0aNS9qBPt8Y5ybw1duBd4VAX5Ixk0k0fZ2vgTjYQERxUBUUP7J5iN4l4nQnghm
BIrM53NzzeFRBej8eaEMuJYj4MB8ygbv8zTBl7IjYV39trxTkJtQEqTqlEuGW4pg
AqjQilkwx0JQO6u9XotTaQcH4tKTWt8kwRk5oFPBuTus8atuoPZSwyyWnG+89Fij
LHRJT95WGzFO8cS/YxDXBGeaRuookL7hHQQPSf50CUmrmpryhdg0iLQQKNJAD7x2
vH4TGhVqYdEAdH23sHYNSfsFHn0vikNaPkovub0Ph852EKESbrXcxDvuFiTXIkko
21VUY4yPRVQHgWymAgM1wwOmMaZyDzGancSGW0SU5I/V3rME7sTgqEBVuPqRalbg
SYs9Xd5gFQyofUwjlTjYnbquTMfjjPg9b5zBPlfvrE37h6B4rSVYsEETSwdqNekl
zpCI1X3Qp2UmlFfiKSolJUd75ScrA952006YMdl1Ac0L9xJi1NoejY+gPfr6zW18
g2vmgNlx+P5zFDqEkeFGkWBqL92xvubxGp3Unjwm7IdvZA6Lf38Kjr+bJ0fHiB9Q
PWNKyDLA2mCykz3jRDME9eH0mxsLcrbT8VcblcHstY1HAr263H/MsjuLiLFVSd9d
0j9q8xCOHO5GcCPh/HE/jhSMmOvbWLYd1LfJzqsl8ThYA4zwJQsLF5ywjZ+XBFMM
4FTqEtp7ngr+GXsO2o+gU9qS2/ISNZN4s2rbOpea35RSo7drOg1cxo1SKHOKRRoE
wMGD7WftB998L3++X9vOh9ZOAKl2C9mz1ylRBWeRTsith1VPLglgQpSYINw7jSDF
xXIiuWJTKkf5PNxQPRzZ+8vQgdqmZfhGkQEHOQM24zPna36hYATXg7sYJcc8wdIa
6OU7zwUKtdJYau33osa892kz10z6xKR5ohaYFUreD2Mr7wgHWsccerkcnNvGrwdz
yxz5M74WMhKQhQV7bylRHR+L7mb1T0s05QiyHsAgmDEMphbcUqseZ3iKReJoZcHD
oiwdZrSK+gcaug0v1Ew0MremfH2gqTVEwTVdMiI/cLMsKPjfIG8NgGt5JSMx44Rz
eTY/QRZR2z1AAdbHQjNINmP2C/dIQxoPUWFqa2RAFeTKY6hfmsmM2x7phk87+ml/
gOuRALKRArp2G6xP1r672IT1u0V6OWy5Rd6JkYO3ymyM8bX2q9KYOB/R9PcYokK0
QK9pwHMEudkKEafiupG4zn4F+Vib06igjcshCIe1IuQp4O0x7ki+AOFKxDuxhOLD
n0rBryoL46iwo48ol9648oe0Hz5b6spKa8Idy1tdymvBt9/M1bp8CEN0p68QoVep
2d4/zwYWVrzOmF6WC9MizEHuUkEiYoslINJKMH6lxau4qwnxms15c9uYf44UIjBV
yNRNYTQ5YW21SDMGozvDqm0kGTJs6Z8kiYgQ9X3nLD0ixfwnyxlfB06U6QP9Sjvx
prRvFCuRiyWAor5/mxxKnmaIzXrc1VEO0B2QHH8ia9G6/InxUOE9ZKU17ZGPb14f
e5rusmGoAGnCXv82X/WEsaBC/urzty4dvt+9EUD9BTScAOiDQtB8aMGeQ8S2QQpK
EJDh2IWtepVl0TbkeuBAzeSAQ1JymzEpQq9st12zSxVMkZabTgBH2d80Pl1oeVhB
atrhZekWbsCZB6gseVk5n6+W9jB8tZR3CbSlHMXCKQ+edcMeJjBSrTGl6weOfTg9
KQaWWiLbYU6omcLo3pmqh3+s2XiKpKMexCT46LOnGVKLeM2BcMzLYsbdlrcfDxGu
V/5rTx1przFhzAJjBg9AYa+WFW0RTHz46OyhlzLq5EMnNUYysxSxfP6HCPZnOiNY
lu8t8m34GT5JjH1FP9KBav1G3mmSW7gK389NMCUL/y3xgLCeM0ABuNe8d/qWMIwF
5WG7YWBiI1pjSe+Gr6HjURerK542MOlKKOZVLw0y9M2yKZMVFfy5Zax4C3wCPjEx
PlqSdhuUCJlZ+5dpdJxDtCwPLXTjIy89AFoQwoy1gKOzrBijW5BiMz72XVja2TwL
yBcH8rmTtze8BWxxpdEY61VlIQhAzgk2IB42AlePHA5MO54NXvkgN4JzKltD7tUb
npfwzptgzePJbsOAEdtQXoEmaMJj8IhKBv0uCdTT+1yEd4JScR404zdXU0kb9Oag
gEdyhcgfvty84cCbVOmO0fa74E3IJm0UiWqfSZWoHukn9UrVVgi2eoDD16nkhpd3
gMiDFbCXo5FzNL12By/L81IyZ2ShPazWf+sQBSnSpiPuHOY5ryQvBC33z1dRh8Ab
vV57yntxEaYK/LTM/aFKHxQNiYIR1tvmrfjDQYwVrwOnDv8dRkFYbBIGUGCFydTE
b11kkhIhvWmyUNlZKafhO0LVmNbfq2SFf7F3/730N7gQJvpXsy+/JXphoawrx0y/
+GSkzEOdC7FPCTYanQdXKX+sQ+0wDxSVCQYAlxEKPT3APh7U3wnceZiFz3lO+qqC
gra4IvRSAPFaH3eROhQO5IfRcTHdipbUllN7T8PVyxqC+ypn05kil7l6k37f1iZw
/fNyKbhtOwkLnrlqq9g3LQs57KwDt1NrmLYHgs023hAe3bxuvllC1tccoDq8qIwb
OzdbOuPck0GeKNnAqQKg4MqksdbWjDzwPcRy2+Nc81rSNLcCQ/dKwgLLsp9TOxt7
6DtXf6tieI1U8IEHshctGNAzebPY1dXkFKNXHwEaKXbT0hV9Q0yF2gFhPKG8Xkrp
mJl+U1YdL5/ZmOgzGWdYQetWMB2qd4Gp6j9SJZKDtzFqGHk4NI677eVcgsufIx+m
OHJ1p3Jpy27FmzyGpXh2ZYtpQdsdRxmUeRNviOh3Fs3Kg+fSyTgvX627Zeek3ezQ
AL/kx5rUhMi9GUJm6hk4rjYYeoP4G+wK+ARLvy5cwMSBKS9/AWBsexm28tqlK3L8
GYEt/mkILbjzegZo51Hryp8z5A5lqhE62V8M0fipU13mkfsdMc4yfQU8r/mB+G3A
Uyngmh0onezTaZ9rNl+75WmODOFZILVJwgNxzAnjPnprNWZNqsL4cDU1SDX5ReFW
rt5FoZOqTIiSdKyBzPjuOBnq7DQzZ/YrljY+qQZPHdAoo8fVhR7g+nY/51cqiG3E
yT3Fb+U5aGpfZdqp7FWz3fRok/6fygR/+XTqD5xmvjZtFD1Li+07FNC2RL8dhLiK
N5C8wrJBqmNLiTEWi886BhsvoeAL16lCNHecWGqIFuObXD2Ro0hlWih8CTg2B9BB
YgdieMuYVKBjZZa8rKVf0Fcx6dRyaJPiB1CTbQdWb0Dd39OBaR+mna9NCp8h1VFQ
Oa57bN0QXDfykf1i3wobE0+mQVBGeHWdb/9O1Rs7jIHsho81teua3JfLdqfZ2cWW
WSy9JnhQ7D9hZl0w8XOe+0A1BALqLECzsXhm9dmbNw1/Xnc4OB5NlplPMncx6ZDN
+SCcKHGTjtaGZXgyBgonpi0hY/KUyY9V0NWLIKeaLzP1B0ihicx7MdjqeZwWawBA
VyE+1kPr8vOesZveU3D2d1uJiR8c/0YDtyRkTYJD/Tu8byx4ihGw1J9nX/mMMzZf
k7nL28hHKflKnNi3L68ZQUiaGQ/RHUSm6mw1BpanJyNwraZZlcfHzM5et37/lH/p
lXGv1iey+harlo8dzrlu2JGyfFbLl4JJG1JWPOMCrK3XFiKZ1bDE/ccu+8H+HP8K
49E2RNal7fk3iUZtz20qTlhRXeoNSnWLPUVOeHCqxlusQkIN8ofCyid+ReD5P4P6
T4xBxtgX8m+2S3m7pn+vPT/Ua4gJpL+Ck7w00s4FGjeDFKxz4nI/O5mlxK3a9acf
3ed4Rfzvayu8fmtE7e4xInqTDvRR+IHw9r1Mj/fATR4sYfTn7WXjJ5G3t5Ckec6a
xQw6sRKxd/DuCrmAAQ9daLccsgLPPg8Y3im0ZclL+yqY3grZwgWPUlwEJ4y7xp04
em8fiueRe0oQecDGQ5KHFgS0BGr6D4MeE1eibon3yvIEsXwET1B9NiCz8E/YWqME
SXCoHtLC/WnlH9NMbRi2zTozKCLoFEVKmstAJzQYI79/SO3hs1hCMozAuJcXCvdv
U4jdrm8hx/L/QdTf5pzTCInGpQP4WHQK2y4Bm/tfCH2jdVWJynIcE9nAcx7uqaeP
cc8CLQVPSo8sjA4UdhCThAdOwV95DlZXhUCpzSirxZ/XIaejakLORjARkR0XdThL
TcPJaglF7kWLoWdpb+ycP4qFrGO/vnWpPoZ7YaSf+d84q3XKTwHA91QJT1HSK21l
LtBRLkgwXm74X7plUaZ9kTno42rO0rNz2S8t219SiW+78pMG6XG0nwsE+bHLkOTG
4C96ZPLTcHX/JrPCeaC8mzoSAabsgH7OSrY92HMDBTe+N18GDF7tp5Galdsdi+P1
0K+GDygXXHXsuY8IOxYhx6fIO+0XTrqx+XPVDQ8kYjM0DPFEw6TVLaKNVtKs+8m2
hQJ+XVkfkSD5pRBZ60sC75ts0JQyQW8ybH8+OKXXg76/QMK4VwChGT8d7H01unZS
uKSUTFygKKyI8vftlzQacx3W1VLxT3vFmqtkkbva3oEmpiI7ZOR2QkJP2QxDA7cd
AnJ03trrExBtT8GKgssvRoEHL8v2XeHZV3ulGUCKhW7DdDi0oEcBCqJq6hSejliD
9ka53ug+NxNph9z0PZEi64e5IlobWr4NkjFAa9Bg0xp1aFqOYNiuChvucMF1a3wq
DPYCOtIFuQT9jFFzMp7/TTxADJVV2tSd+EqphOnSqUZXtL2hM5Nwx3DzaVLFrWV1
x8Pjhs9MIWzcztkon4FcN1KcfPdCEGi7PgpQryUHD7PIoH3zO3C66l7glOkuylSE
VlFbmRi7z4zhcgkdc0B4UCDOJU4XAx2Kr29oNCgjrWo9gCxJGa2tX0CQXmIWC8I2
UNqGMwypWFTqRbS6jrqDPVntVc8ENLMeSu6RQ8OXixoHK0zn2IBq9ZWXWyGxdYSz
meoOA+5hS+C0qDsqoS3GXrwddUct7EIwwU8dr9irkcTVC9WmwjVKICXXo0JfEXn+
M5t7kmHWzR3Rbe0N/UpMfgopoGbQ8wmb9rVd3fiSdg9kbsgQ2l5MJTpdsmcoqOVt
uOIhgrQfr02+j9UReB2vM8OHk6WlcCXMRoA+ghkBUkq+8YgckXzRsvZaiGQ8HQpr
CeoFmwG9E2YCkKiBbpoGUv+Yi+59zIPXUCWpEEfaUY/VSlMdAusEsBAfAzCnnuDg
1JMANF5xEQoUSkZH4H98T9T09GJgwNwAYpULR/HZVplCgFB6HxxZJD5yAtuIiSCB
Gp7v6nJmW+2tIY7z94O5wi+57cS5ONNMKZ6o8prWjH9NrYkLJPqu5UuhHMqn7aQ0
9d+lfNNd/4HyRfE2VDGYCNu/ihll1nmYng+e2duQ+S17bDRFCzz+b1Q+Yx2dxPzt
8eFfi7ZDoM/qVvxsnWbynrZkYxNa4WEwVkZMtQdyMWOehpdWHKuUqZB7w7oSndrq
oHR8Jx9YMxuW5H0EIM+IZvGQ9+3FFkcqHIe5Ax2Is8r0iFoLqaeQ9+XkW3khsEZR
jxRMV7UIfLqnUBQrbQ5cSRbGe6aPKnIlkoJ+STlnwgYXBtdgyDfZI6vxuta7UL3i
9REX4QKWlP9J5OJLY/pRguJ1PfnEDOin/80E+fkdQ5UEzCmczBPprA/9qbEDzzNH
PkAgyzRJsUsmDpqPM8ZfHt5sKpo89gJefRlmTl6tS/pWqfXLDInx7fAzarI5O+Qe
YXjfHAYNO1q9idSxcwbCNg==
`protect END_PROTECTED
