`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AopD0WorYKdAB1QutAM2BHsn09+XK/tVnt1rZ3LkESQ91BvsrmWiMQsJ7swVGQZb
mObiTvvCxmrcsR/I23Rija7GdN6dA8feFDVo9hoVD37kXYQZ0kKXRX4NBT00x48x
6zFl0QooZ1BFqEC2AMN0ZEHK+e6TL577FE2dobPLanMuva4fGfoRXDAriBQfYifQ
6tWELs4pQZOwmo3M3NKfVw==
`protect END_PROTECTED
