`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
469jsmkyPlcwo7H7bukLbTUjrI+PIOvS393amQPyJbEW+LAJCXBgLZcV+KPo18y0
CS7K+NVkiChAq3vvhZmVTGFz5Gk2x/i1e1rhzi4WKfTKG7VSYhlLn+ufYzmGGbXT
4rYNxfAcbsY5DG62APCCu/gvAH44fKwmOsFYDP3eWnY3NOjXpetRwruE/whS6YMr
OsKEbO+Xn1Pfn38JudMurQWUQn7GMHcUs/YyZ8frLjv7OwYk55U2Aq0hJHcfWMOf
BHyZsVrFU+TBfrCSXGyzzhihZyuQ9ZtRXrt8BQd4ujby+6zq7tnBxQsY4PC5Js2r
mLp8eyxG6WPtne5J3kNein4hATubxLMYysGOI9wdzcXUzisxHiyMgphus7BKLG7L
vsWzaM6WwxZek2ym2Ri6yxywX+P4XZFNrTVtcehTejDBqItjN2ueVIFYkvDXp4X/
LTj+zxBDW8EVVQobZtr9UgdfmqovK/BaQssOO1YJit0Y5j7rZR8MikalX7USuW2p
ks6SMgTz7ogexuZXyhKHC6YLsLhES22PZwn77TxrFhCGWTZfjb0sZTcKsi99gqUd
VSYbSnVcToBB5uqoIVOJgB4lLy6TR66NI33Joo33Lm1DkeYmqy/ZhS8rdaCTITDP
1EqsvkayYp8gTftbtYhSFpN0EnYk5VrKsV7mpRHZEBigZBInlh3SmM/WO4Fk8E02
nIK9Z2upCXQQH2myMY1tgfwCIP9lmY1FeMh8O+jEUsD1nnidooSWMhNsYjOmrkFL
ENY+foBWSTW8Cd8v+8MAavBqB6iH42XPiquhvKdv4HsvQvm3C+gSImz0iHLg0H7M
E+rCVcKfQKinohaUF1nl34kIuXoAVLSR7yLiboVFpnxLQEqkHlGn/cmsWYuzfWAU
0n1mJVGFw9MxvYz1z8EnrrWQP+GbXnc/AjBHZUOcicKGqXKxwSvu5QHF+1tdUQwk
6Y1DsHeEuW6HWMTWbPf8yP3U3cFAbyj+F/AcLfg1xWHidGKe4JdWcaZofh80oiXS
6OWqFzzK5lQ7xxCnpavW2jO6e0LAnB6sNHzgLXRchzJyQIuUvxPI47JAx5BGCXvg
gQeQKzoOSWLVjqzzoJyUgdEsLvtfKfeac5E5c8qZQvKWXJfmmMnmobRB2brA621G
ayNwhn5Z6BNMshJHqrWGIA+MoQcHoa53mqivfBWF4kFXgnTuDswMVyko9ceSBumq
`protect END_PROTECTED
