`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyFjXW1piAb+BsrxtKM5iwmffFlLietAuEKYt7HYP6rnUdTKzzMShCeTUPydgVRy
CZtEBeYIveNjK+B337reW23yskzgkw/fTMKM/CS70jbKULa7p5fAVgRHwIDz1oYG
q3+qm+lwz2JKjK+/jqHQ9CEF6cLyczAf3VO3DF5BJTuaR5jpDKnkKZJ8+eU7iUrI
dD/fHv5p/DRxTJtQO68QfQ2yWbMVCmu6bZb80m7ixG5mblhmWwGH6NVwxpT1R0Rs
zVJRzF9rvYA6wm3jBnFHqWciXVX1kyVYRUBjWuib4SBtXGx5HVOd2VMg4Im/ZWHp
T8JgLvU2y8qlys7gd0ziTanphm8JuXDzs13QI/Rq7sw5c2YhZNI/Ns9sfl2wGY92
V2Na5d9nltCkB7xDRDmZl7Jf5j20OIcvrnGvYH1Q2VNRMebsaTErPmcajWfGf/Tq
9xZ3qHpSchPboAbZJj9rITgNYr1+/VuIUZgcxiBmNiNX1JhYBjnoJMFRVpt82bsq
nkDgGfQi5WNyOZN36LIwdGEBvRECyDcvihDqDDfFDHhB5b+wf9O7eM8hEDvY0hgn
3byjik+7WPZDRO1RVb20vUb4uW03vyb4GGfzDHVXXvmll6q6AM4Fa2ajOGrAHD4u
WBo/GQifImSaN695r94Ahytsd6grOweuZhZZPbOY7uKvtZTDM9+W7BAEUjOMKu3w
NWQ+CNfTJQmFUYrdL/O5dZVKyVN/X9EeTgzKGLxIEDgHN5z6OQcBTlFspCGNt3BS
4eYmHFJVSAPc3AzhxHnGESVolrhn3+6jLLBzLzoJ+snUnz1+WCbsh46p2LASf8/T
5LrvkAPCSey/qpawgWz718kxR9go1WlogUR9l2U/OEPOHJxtO89sLNsYknkDNio7
7wUHToQNa/ZN8YK5pIE4g+Aqir2JZpAOhKX4h+hX1jrrmeZE9hC/eh93+yWwdZB0
1q8S5P6gQ9K7BRlZ80fuYUa/LCgLRq4S7GQJfa8zsOOSMkLxMhFj2mhMZq1crNCk
8dVs/nFJoueNfUY7n3aZmdUOFMkuDaK06Dk+B87YIc9Oa0I06sPc8/wrHaChCtpM
bLsiF4Dbw0QBiPnyvQLR8IP9MA+ZZnSuo+teaA2EtNUd92kG1wzD95wUdHi91Tho
cAzyBKIh34/16tOUIwJg5t3TuOCIh0Ny0vxVzeQCU5hchqfjD8abAUUtQ/kN3sT6
Bt6Xo435WKLSxaOeezITVafBsOCS1JU6HMicfzxkvLSApGS620z7Xp8SiPYAgw72
Z2ccvLKamf2w0D09wrU7J5l54yHQe8IiO+V0uv1iHv0KX1tiCZTP1Z70g3TuQxkk
uKbqvWJO/fz5uQkwlWIw8Ywm6Kw4zCtgoAqY1TGlz8DoBTIKYXr74fLoiu3ym7u/
r6f+2utTzHUXGbR7cogaTnHjk7uz7ag/9v9EjOWnTm0uuTlcyb2SXA7PEP9bv4t5
gcVu08YFr8SbEj7RXmsvYWSI6uhxMopZA/tFqYwD5H971UJr4vDsZEgFvY4GS/zB
LgRTNSsfVtUebSUbcOlrPyjEwl8r7hMD8FSmhykwzj5YMFB2kkJkZWJwnNKweLmN
dUCj6m4GQcg1tjNgxnvHbMc6DCWnb54zPq/ErEQ1I+G0VKuGXqJNjNRmGyhowI1a
3OZQ7YrutFIHq7P+E73bIaZtWcOjgFEEdpW4f4E+YMwKRBtZTe1U3juCPZTakhDe
pWyyYBaZ1KpeFhYArrVmL8ekcWk9NZw1lHuaR2YQVHHZL6hqVtW82TAafx4WWFX+
xRKha9AwekeTQrRxQRWKb5RzVRV2WcQda3cddMS42zd2k0g2F4RDjANA6o3Auln5
SpUTFEzdHnqHcP6PA77IFiOJYAW2qKBfxfH61nhGf2L2e2MWXC6rzqS40TAogYoK
Py10TNAFzjtWDG48j1V0+ZXxNXllSI8FsHBeHqVsrMYWEW73hzdPMV5SrU1EJIv+
baL0S8BNfDHWY66NX44thlDxRNEzZXbGNEhgwiSHRnc/hBMTJCyqAA5pXiT45wt5
4fHzvwHQdzAMsSwmum/eOhSDK6jbefMsBT0kgfg24iEvqBoy6To5BrkCXrnh5M6Z
0fKRpKsWoPqNT+1eWvIbQPdPMNCWUnq0PBG1LVGt4dE=
`protect END_PROTECTED
