`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+gZTwt+Yqo1Z3AWhX4lq2zu8hU30MXXVxPkOW6MCN6tlJnPD4g6ilcrWlroNca9P
m4tlT3HqnvUQuriD17BTeUW+z+RW94APHVn7tBxFdOYSSyoXDvyfG5KatLhWjEEA
y4Ic7GDr3KZHFVtQZ5mV75L6Mx+fx1mblOvqBQ01fvUuavP6G2EunD8rUZ9jf/3J
E4JRfRczJ78rcmTNZ/Qx6KXxnpITpvFitMwKFhnKkme0llluBFRtvkhvcIF6lerX
/ykvmq7NF/+SogN9CB20P7fGWz0+j6PgLMoexXo1++qj/LjP7vCyefpuDfTmoydq
hoLpiyhvqm7rzT20cEnJW1HCjQQdmUdW1GtK1ZrXHbkArw7gbegshBB2YOsIvntA
8eTwlA+wP2mNTR9I6PPS/STAkgCghWblDvnxGbyDECXxjV9+x2SEjExoisPMLgrE
ss4yFTAuNjYl6lJIWFzM+eFmzZ0RmRzTn6U/JEfsXUM0IoV8g6c+fB6MnDNRFMko
bdKi/YfFgdHj+VuDYpDvxh0MN+QNFJwd1Bkjg7luTWrOlkL8ZW0PZNlB539SoI/2
QLFN8HXz3TPKwnQy8I7omLhgkYPEEGb1nkZosQs6HSD1MrknEcrBpICOCvhiwz65
bGfxyPvSJg+m/Ca825vcvsuta/7iAwLUkiHgXRNkym9uUA2r6aiAlNaPzUy1HM0+
cyxmyVvHzAFUGzkFJf399jGyJfiQAKm9bjhqzPweC/DRSW6+VigSkMqJAI/6r6sW
Y5Jh0mm/PFYj+ZL5nE43DBKnWbE/L2crwJxRk1hCi1zlYgFdfXQv4ES5Nnhp8ymA
02yMnnTbhUoj4yNFc+5/9cF/L9Zc5kfDg1VqqcDeH6eSL9ak/pVvNZyd1icpyHoh
n2oiI1U09Io2TlCYCyXdCrjyeKK5eYVXqLtH66zdbKrI4gWs1OsEGG52zMW+v+4A
mb2lDZqUaetA/VwlLN8KwN8X8nnxuabTmyKp7JMwjJckLJCVmShQI7k1IrEZolUf
DU3qQjA8ytRLZANjC1Q9aElrKwuGQyytw+wo7DnTiM5y76hgB9QtbVFp1JVcH8zm
yIvt+68fJJLXdLw0LMX8IUbHQO/9+YCKlT6mknOAqT1xn3ROrL2hU2bZ3PCcZaWj
4+k13gt9W09/ZRUoQ/RDXcwaRAowxP5Zaowm1f004SRhqdIeAj75LPNs9A7E82Qy
xnjQ/sUGeJ3kSQry+SrB1qRgU4SIfcmfM2bxMaq2MFcSARcJtj5In2uJakDmFyOU
mIgaTI3GDawGYgFUMLIaClk952kHR4YZKwkxJpRY/6W2xLptkoaPOIU8FiZG3Hs8
ETFcnUZ9RppxBaG6xga4ggXz5+oOT75rY5+NwSauwLk8iuP/in1R8z8Yl09d7XoF
187Yuj3LIw2JI3c27yFYNua6l0GKmTqeq+GzCTZVz6DpuCIcXDNN6BNK3qHtwFlv
qM3L0p+8W4Ze8NzDV7PStWNmvCE9jdmaTTMOsNa9Ktpxbb9pjmth23vNqBMXlo5A
wU5ModwH/oVcAl+i3ouVTcQvGv0wY3p+ZtBB4ACmrMJ9vlaSUMk4I7jNGlXKhypw
qJ4EUUS/36+FMRLyUd28X0+RY4FBWPN58/ahRtZlfj5hIRZcnaWQ46seFkXbtEYp
KJk0jOgBoJRE2QzIm9VKvJ8b+erVq9oCzp2UMq40lxACUdhWk/s0QDaaCDSG4cAy
0sQ9ssmkmq6t2uprubB5CwQGGCo4vodABo5HSmmkQdwklwEqP5AahZTBxo03pnRr
C+n+wfZWOdc/GYca/54IO6Ws/03cjfV/LxS4RULq6o9KQNlFwBk4rYDoKb/slCZU
yq8JETyzmG43s0xnjAXDJBjHmtoU56g+xFmm4s1l6s87PlnBUmmqoqFia6GR/9vs
eonUeJYCKVZ5waxK7TtS1Bt1XX/R7xnqoww6QuCBbAOcjl4bSkt8ZkTxNtlBW4Gu
V/cRCZwv/nq8urso2/GSKauVRuKN9Wzku9Gw/CtCbyklWacWePwPHx+0aNJbTNdN
UDOmzW+md8FB31acYUSdbN+1su1TtaEkzk7ZEFGbNWun+L+BJA+zxvsirK6gUO/b
Nn+9pgqqIcH04FnSf/OWCuEFqYT6EUF3XJWfpfsq7+f4Buar/UQSha7b//iAPQOe
E6UVEhmwcOQMo9oBo9J0FVOK3K4hQqYhgHBfLErsBUfDCdJaagmlxzxvwZ1t48+8
lg8rAQZH+ptXu7O0fcjqd+c/56kT2vDXRD/xEAv3Ma2SI5nxTPYvtmjoX/jUX8xe
Awl/BoZtCCbLqsDJ8wPTJap/rkzNRqe01zoKh+e+8d/QYc+zCIK/Z8LcHZMF8QOp
WHOMi9GQvqct0NI4fGJ3NpqVJ751boJ2uS4UDBCwVyw/4Rx3N5Ofs2UUhAvwC3it
wcSN0q0EyUKq48P6t5ZSadf2S5GVi44MeHz2FqbpUI/pF0eEapnYKlccVItWCpPH
j/uhtlgTK3djee+ggH6x9iZpbT1Hmg9z5pBbHMCyJ4RQufB/4wBz7HJWLiN2KC1i
1G6lHGWClMXC21go01vL2TZUofN+5mNucGFFthGOGMtL6ZE3EH6KULuxCvvFNj7Q
2QD+lts99GJTb7JDq0j6XXKM1sJaROKhSZIbYL4DggzEh1ZGeap1kRAkZxNt/UsP
xOMigcmKSRqF8BK8Ux2dPaxjjEdLtVw2rsvPJXlfq0+MP1HgCFMAEHHu7k3mDZPY
EP9Tv1Iww0s550xegQgyibW63OlgfqSPcPbRVhP1dDAjHwMhzEuj++AO1uOiNlX+
KAuUkX5mDZxI+VxsYpa8dyWvfqBw+4lIVSet0jlJkxp7CeX6yV7tPo3p4gXjHpCw
glsommZ+Gru3Aw10hSYGq4OqynWejxfX6NwJIIT9hTwhqLEhvKwoO2RTAvXBFk9z
YBJp04358+m7NbMwx9ANUj49n6gnbHyIwQ4XiORYRS/G5xV30vWKjIBtVHUqdXpb
GdiXzg/t2aVLbMhV3aFqmosy4cOi7z6awm5lNl89KlOfNeyzCSH2RWXhVDkoZ+5r
T/Qc58Crwl68xjX9gzcic8k5xlOY/igK/HlZmAd4taK+2hBmTNdPxcHUFWxF3ieO
jFGY5Wu038IPXXqx64bdMWfH9XEkRYBucbF3vxHnxLdWd+o8r6USJN4MhbkOdHma
M6fSZ9KyG4NheJUcThq/VnCGwwD9HHLt2JCIzULMXSLYPpAHSkB1A1VoosS6FHvX
qyg8I4x8H54ASkREB/digJGGvDZP//VHlXdJWYczKqUCWyLWV5+3vb9JjDfrUTfS
r1XwACwQpcK0S3lyASji+CsS0MmzGuXBfhAX9CM/37GWMwo9IbphA0SSEHFoqbK8
tAl6Zr7j0jvbw29mzk2b5tgr6lm8QE8c1muzJC8eJ7x0eM2RJVYxjvDzjVkt8QJd
BJKixNQX4k1SJGIPj+7mIPssi/0ht1xJKLGx/zFk06WzZJvH+BSG9aD7K8lBwl9F
kOg/r+b9v1ZU+H6W+ac9+FD4YqJ9wiKm0uXAEKd8LWPSzDKa29Uaamp1yaTBP2Iq
YkWKNorA3bnHvWbQhlkwMHDQh/1NRgpaaUZaUH8rjfj+HVjDXqhqFKJRuraA2yMK
nE8SFFx3soREKnETbhuEtPoFby/vQAh09s2AOrqjd1NBFmIC6O1TcJkjgWznX/v4
old/f8IfU7PMnmdUsS1rAjBSx7vWtotV/yrFTIyRAaMba0zynaZCeiU0TUZscX6t
1JrFx6DJ9D2SSBbk8TCKZZcaItyXNIqDCvgpG+uNfvYTKVlOkrKkZ/YkMq4JRA/a
AbNS8jsOrr3Ugk2g8PBiU+rgc2sKdvZXIomKyWRVHDZ3U38HcJwYtFbpHVzyWhJf
sIkFmGSjfhgn7GaYpZ7txMeWP6iAhxEnBcRtGPhTk6Yq7PL+mSKsgnp/iOFHPJoM
Lo5JzTaPjfhWrJKJwBwTX2uWdVOEPqTMNNbxRog7YIootjoCgtGdr1nvxw2fKYIQ
IDhbBLS9aOa+Sp54OMEpf/HDotfhhBA3t3maMVByUNGF1X29XdI+Mk3pNrUpRVOe
BdWd/J1HXcye2N9ghmwvs1THniAuiFj+lZ5sS7ijQAOeQXHAorqNPVOopxlgJTJ5
3eL/WwOC+EB7hxobSbKDCd2RpKjgfKiAUdl2kheTAswrBkw8HYdD0qk34IKO1GHZ
M4t57n2muO0CappD6twoe9Er09eGveg6l94oIXtiCVCBJQXbE3CGanVAu1a2zVSM
6jaHj6p9VmcJAS/XmUoxMcjyOXdXc5vHyfqMBb6vlwqu3NgDnuVaZ3MKqwAX+KFO
G6+05NUXfcfuHo3adPzHUwUDIC+6EAr9YhboPZJWzxAaqW/u/dh2ndgf+iOYtyKJ
2TOa/wOMDoWkkJ3lj4dlyNgRFdmh4dtiq2RAbZk4Kr45yUGpNuX9xjwgwE4F4MpK
s8zNmM8DbLRIORb8jXXo4R1dt+iDQvs9DFuFQILYi8XjAH3desXCNI951XqJ7A88
W+3PDPKHYUOVnzzxTCimqPTb8PPHKQTxrgg/D7JqbEpiOOn0GHk/7ovYdi47oxmQ
85X/DlxdIbiAcGIXtm9zcCc+DmSL3tykhdwTwgISFUqkkYk7tTRgB/My1qNI6L4v
ACmPDmdhAVcX7ZeqOsJfqSBgj+ASkji77BaNiSzNn9tU2CTaYpyB5IjQJ3BFHLDg
Nl3EFVNzFy+I9vOD5eHSx9AXVYpwWOGHTZVcUkkmPczMGO1YQTs6LYLXcDlxKN2z
yFWEyPZqx78g685o3Aez1nJeeFICJwMCXFvkQQ+2nSWuDr5oHVhxtgSHgJmzER5F
1h44ljb7QJnEyL/q69L7JvpnhKMdFWu8KS1wWGy6pNFroCQelzCyVwg1mtTAGLTY
hPzgsy2wHy1XQhs6xFOY4+/WdBtOOF1XEj/TkC4dnaOj3MYffKb+vf5Dd5hEl+zj
WXLY7jMkUk8bDxsSZxspZgAg2NzoFKMGDBcvZKcy5F1h4lhIzYiLJdx7dgNwE90K
u8E7yV9GDnh3jG754Z9W92WVJbz2Uq6HdDdSM+p8Q/I+mIIdniOgHkItNpVv28AL
3UlNHlRBngC/r8B7VJCzpjhLYF/DspMbp4NRMzmu26QG2C/0wkYez1xb+kaYGYSb
LGu7Ql9KrQ+KNL3QcYJ2w/oEgp7IkWw7GOlsORs7n1Rrzj0U7QsFLrj2jO3X2fr5
jM/9G+mNOXs7Il3hZRFyWBcL+6dBDc5Dz+qThRpfVjeaLrJjnY2TL699RxN6A8PZ
0o3DxQTAO7SioLF/Wa8lCSop5UKHoRiwzlNSpy8SWVSEzYCMnsi996/5wCPxF97j
rjJ2ifEzzEgAq7PezFcYz3xdExSB2X2bP9YyvRNiUcxZU9PyDbcnryLrYrGCN1Ya
2xLUvR2izM4gaby4oD/icUVD1nhCOYRJ7SILrnaoC1Z0/Pv6aInT1lodY758UAMo
IlH5xEyHMyB7/m5Wz47NDiSXNbBG10qdtWPPbeTZ34qOZzO4X0kumHFZ+nSPW4Bn
3vK1aguqw55Lplw7ZQbXpWn3XRPopM7Fs4lVubL7NSAgMItYYzXkf0oj1WJbu8Cl
FiaHUP4DqpPqFW8cB/dE1BiK2EvBZjkfy2b1FDgiRsRGrvYFetEvcXyiGgXujbqY
56qoVKEp608ksujM2bvX2zf3cp7+PTZfbbeJaR+5wqXaaWEGn1FrFXp30DJAs5RK
g3VndZseCeUJkOSlGDFVNXhAMMgeKPabaKPYuKKDMMoIDKzy0D8XMGcCbtcVcKYd
Y0qQD+fpzsKwqztYuI+i4DfJn6VeWIMkb/XoWHJd4WySeozlc5cWclz91nFGbC+P
A/4MkMnjs0dlsLv1zAX6H6pQyrO2Gt+0DyLkmUOtC43y7EdK5iMhanjixXtyESTd
9c43xDtspnk+aQ5qVch8fI02m27Znw3PuQwflKukO8NburzGqYsWaPpInk5uHxMc
OSP612rud21oslqO2dXjo9AakdpYoKGDicbiXYdAAdT7/j/Cfw1ecAJcrKtzGOrJ
+IU0TLXRVXc9H6UiQ1qohDXGbrp54Fb9bBehZpj8sqkTPTub9VkqL6D6zltjMf3/
b/+DastaxakJVLQyh6Suiw==
`protect END_PROTECTED
