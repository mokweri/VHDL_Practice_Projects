`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCYf6SZ4cuiaxa4m/soNa0f5vroXOZeH996UmJurOEOSwgBAI6+8EiVy2Ug4V1t9
nzwW41p/YiPYEmOdK9/KpcOQ45imZBXkJLQrxgXDTmFOpLLLRSFR0cWr5uLKPEK4
actJMTzvLNtPeyxM5FlFGLGNlYCDEplXNs01TN9hjub4cOBimatDC0fViwjJgDT0
CAjN1vZlCbn9MTLC4o5+5Ggr1wQnmYQ05E0vpIkBglU+gdQMWfKAcad4seKAr342
uOTb85CRIIYpi7awRdGm//gN3VX/3hpQoY527CDkx7mHbX5dg3wiB18hZMT/vCRv
QnTIYMjc1Be+WKCsExNJbBtcYPIenutvJOEkyGuwwBztne/TLQFfExnaoxeg/SxQ
WLA2OYD0RiEMziDqPk8Ohfls71IZd9G8cT4FpAJKw8g+ohZdYRqVy2vbbA+IyJeF
1CVGcFx78X/4kvZoFNQReEdKWrSDSsoY9U/1O3+5ka0QGJRoLB/C6x/WICWl/WQz
xnMFvrpBFG+gpRc5Q8bd9o6ygIUeBh0E0Ock+Hvmqo1hVNqLR62FWEagMrsMPbKs
5rzT++K18Oy7Mi4ABEN/LCwcTp184aJOKll7zjOJYzK7rfL8PNTMZI69WNcsrNZq
Snhf4+ErQRnRouH/fq15yVIHtfs1434wlOJNA5gsx8SLjVtlMv31Dt/tILZSKGTO
RcltR3g+2iwj33nm9NAPcR9LpbGQW9pcmu/cpVmzVIs=
`protect END_PROTECTED
