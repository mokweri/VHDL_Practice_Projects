`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldDIh/Yqh9jNyVppvwcSoj4ONH1OsJrTEvp1YCBk4oCLUEr0KsNwjSlfhSgdmj5s
frqHZp2k2v8PQ6HIg2suCBjZNxcp6T1xL0DM6pSmZH1ETPFgA/4nB916s5Dql1xc
WkDhRakJqG0RyBhhtTvyAOUsYLhFtIoTQSQbPcZmLwSAm/NlFkGUd5/HuZ6BnCQe
oezJPZXL8GFhR42jNtfgtxVj0cX++8Ofk3efwqVX2b1086BRWXY4NIYBkEIMQAFc
lkvsBAnbgZx+pD0kEi0rsX6RX33eNu0zXEwM74jEoL6xFH+JGRpExrRCRwz6mwMK
Ayrds1+9ZB3oPjLtYnm3AvKXfkeKG+huzXtPe6yAJoGJBVxT34F59ki5SKO+JEy9
wy8DyOzbAKUb23k33fQRdE5R66QIIlFo1p70Z7HarhFz0XWKHpthuXrb9fCN7SBB
JGanwLTg2SH3FmF+EySET5C4YyRw6Uq1l1hs+0gHROtYnUOWm1OjP//C1telO//T
grsfsbXP0RZwIXmry1F+mdGqmhFx+d3Ja5sG5mjvu63uA8iwiuTZuN7yroilyN01
J0js/jznmh+emVFPWTy7yemeeuZTD8X96q6rKwhFfFiBbljt4P4eSfjgKP/JJiMl
DCZEEAFTJML44Ig11ecJfURZHk8wDVKw98Weq03/BKENqn/tR4YCmj6d4Tih7sWX
N5KMsMzNKzdpR/iiv5sKoYQ0Rooz8xw7P34EnOGZh2OyVWfcJt/x/FuogMecLlcE
H1KNycXctX5x+wKy0TsKCklhYh7ZtCryEEs6XIGKmiaQfMwqrnlJaqdXot1R//dH
KCX0LFFGaAXfrbgy4yRM2NcsBEZa5+PLnBUvcAgausd6jg+1CvZ6kUaLTUf03xBL
olR1NqdmlWqffBtHLOtkDtOj8w5ioAW29OsP169PPaRHQcqwIpbZNRzYvS61mASH
WJCO1B7E6CcYk0284dI3uWJ61VDZcXn9hWPw1d8xztXPamVOZvandnnIMoazkaVD
Mx5uN0i3+RGRsCJXp/5DxxVZnPo0bNpnCZXFOVybR4PJj/dVIIh0yZNieCJqULzs
yEt97SO1y6YJBuPZbD/avGXYlvOCri4gkWe4+l9uDHhKZW8e4wYbfn9JUw4nWw5h
RoOmogF9ODp/w1KSOpa0BZaf7fI6BFVOWMihOC/xH2i3AHZqqvfubQz48tr8b/i7
cS5562SqL7g5QNT/vZDQ6CKBAEsnLV/+2KVym4Q+4WFsnN+yH3GgqpJc6xlnGKxH
JguybwUzNN8YSEuADGzJH00g50h2XznkK990gIZfB1LrV5PR3gFxOEZFOHWu6ENV
5CBo6PfdzkAy3dgnFGPIVnH5N0v1pt2g2bfV3LRh1uWbZrM15Y+hSY9aq7OKRYr7
FIpLZhOn46ubvKzRGqHyIhx68ssT7qAWNoPJrkVIdrJjn/QWBMSPXxklH9hbmGzz
8Y0KVEJTy5AGydvBRU4M7UGrYwUrvr5ebVA9nLwUccO85mO56qcYrStZeRpIAA/c
d0je/meyvDPpNHejkWPXF/dC4W4R4vYw6wXDvYokqgMOqBoWTJlVv7T2x38e1BR/
HVc/hu8BNHO6kSlS/pMIg9VQfCacxI9dlAk9ppw873KCu8l54eIdq2uGNPV4hNdE
Sekmi53mshIYwbCzoNNL+0Q8s9D559lJLGTOpH07x9XFjD8elqV8eT1q5nvKCd7E
`protect END_PROTECTED
