`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nz95Cfb8Kza2zQUkCdC3qmoH4I2Foi6Bmw5vTkHko5bn/P5gph5JsKjTUxgzmYEO
m8RjH2GmBMN0kyhCh0KqS0j3R9G9N9t5sLLOr56u/jFsX54VX6e9o3dC74YiLmcb
qXu6Ldmbjc2W74pFnMcY3XocR82v1St/8RxABibzWjQencb/Czp86rbnieSH0lkl
INIdVorHutxIz5bL52k67IO7j8Wzzv8QpiwusSo8Kt9nYESQxpwi4vfUMx3GIr+d
MSbxdEdGsKX3C2Zfyyu+T9oPR9PrjdbTWp4U9FXE8zNBsDZ7D+RugGOEiMfGQKsW
yAf1Ud+GYvA5b3t4AVXDqMXixUMRoxz9Aca16I+Fs2LOOPQ9J2yh2DKQyYD3aiWJ
jlvNZ/wcT+kiHjWiHjwzdhX1M4BluwW+Ej+v2wG0ral3yO2rNWLT3IlXA/a1Lc92
dbKyaDVCBO66oQYSIIUQw5Uj9bktkNv+Z55abKnpzzf0aY0rlqdt+7UTmnQSoU7q
9OKaiV8995ZJDLbyizCIfPktWJO9m5F7jc02St8jtnmCn30ngmAyBD76qj5i5BMS
Ie5Fo7NZFPQHfPNCZRQVcA3BEStKucWa2fWQ7WiI0Gf1DDh73OZdD1V6H+KKnCDH
27/IUao7hdT4W408mXZ68E3H4FI5OVnsVkGBadzEj4yXrFnlsOiU2rUO8mHTLuG0
q6FIzvRl4ThMASZ8zsQBHJZIFrlBD1tEkVb8pPAuetm+bo4VUup5HMxFyl1c0iGr
XI+GICm+dJu9rBrrN9rAlUKAVboAWspk33fRt/ECYgqemv3Wo60zfZWQxH1F44da
Y/GqbnKBsn4nsZN9+LuBsjPKKqISG0pf8LDFD8I5ksh/WHEI+NBBN2/+UdycBt64
LJIXHkZax7QI48Z7+yKyO9TQ3KfB/oeSFDRVdO6W8tsvJpwQI/IkGF6UNqzpkRhf
Rd2Etj/fK2YU1plEA3VdS4dpe0RNinEUbfpTsK4jPOM6T/oROYraNnVPMTvsQlYo
6xge3fz3RGyBXNil2+H0bM41XrTYsxi7F+nu4psRfEjVez1boRcM5G8svqWVBit8
OOwb1Akk+MEf+fdCokTnPCbVxL31+VkT1VYj/dT+6ThVqtgNVhdrfQf4lkmrw9dY
Jrsp1ApmlKQxXcbdXPGyM4AW6jWVgXjIKN83aI/qTx6GPjJWMQuS9lzwhEK5Ly1J
MnGtaWx3ku+UvPFWSyMMKp4v57N0/rpQa9tIfTDc33Xn5P8ENLHFZXH5dQWJz+k1
DaaxLeCm+nNl5CXI3cclmBEdooCR9ld2+qR/jReAyTjPL4QmW6Hh8F+oif9KCZ4v
hVz2yDdwIft5UF9mLDsH9MwqyenOxa7zK3KYhMe7vgcUv1DfD/n5wHPwXp17Xz2b
F3hrbS0dNAaehUXHy78bH/U3wCQbvwEFNSndVYi2efXP7g50P0JT0U3ni7MzyAIH
4fHPf1Mk8TLn/bmIkEn5umRpV/mAMRbfSPTcs0FiYag0oxETaFikIvkXW8nkDXPS
Rf05jcNslE7SmlRTQxURv2jG4NJKb8ramAG7VIoDViIWJiN+AZkQoF4B+lhg9vdZ
`protect END_PROTECTED
