`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkdzdPGQmQxHiKHYGwKElRx37HDlGt2sXu6lY4xUQWTATPramlINHMjcF8pwQq8I
MVFRU0xoYWSW2OI9H3utU45KS/tDMwdGQaae+GrYb70h7KVr1oCJVXQK8BQMoZk2
kmiX0M/8rkJcvBd+LYpuNze59ynnAowc1gcGas5VGaSztPZqiQgzU1xmq8w28AeJ
tRUkrr2i8jbbu37OSmLwD6MYYncyBF2MVqaM524oS+tPKF1VwWAc5CM9JjuexWFq
Sti1jjNtlvfFQjFyrbTdiq0j2b+ly4Dl2QW1VH54KM6ByzPlwZJ7bL1+hQxK+TWm
kk3D9hasIkQC5SuBKehP/ciZGuOnq65P8jJRDbuz/VKRYyLOzgvMvBsXeWi1kJlj
2bCx1HnO1JfdZg29EDBGV8l5kk0BgyVTHTi2znli2N+TnzrHWR00sMicfya3N8pt
xLbWPyozEc+/N1GLULQ79dBPvBE4RpGPg5xuvA3l8fEPRZ5GmofFWA6SaPFDiCP8
2l24PjuUyxzrGXh+6r1TkwAAffxjFz9o5+bqz78t3UbcMBoeRQCiovdwuHl+N6lv
jR8/etwcnn3dQmU3Hx2JvctSUmAjuzLPoajvYbNkXAhjmLb1+iYq6pbfppIyNL54
MSclsqfwSsT0CB2EdbgjWMkHyNMrA5BSUif5Hc4rLPrSV4G4X2UxAgRDPYiDNKct
3BX2zpqO98zfYVJdLtPShKZ4RhQhZW91bHvqpqdk3Miczh2TkfyAaSbmp0vDAZve
8qGkvTKc1hKT6JYDR4pBrZjQF2q+Q4sB9gW1l6WKlM4xilXDD07N67FwegPTVEp2
Cu98UmnzzwU5mc2lrfN4UAVGij3VtA5JPQQWBUPFtANL/Rq4oqjOpmHLlcdH9CoP
5KBibdWtAIUdptTZ7a+Fz+TJOVfYAO1N65+R9FBIhTD9AAQtJPc7grsaDxnMeHfP
jycb0KlfTq+fnier9XD/J5h8Fc6kTaqhjc54GSO/tFu20U0uT3eqPTOOlg0brgbj
FrhqcVdHus0tfwc98e0e7vqLf0zc4YMpTT6JsYALH4ShcqWtlYgEdaFbS1ZakSFF
Ls5rIEBJZArxyYLDtbQzP8Wu1B1WgAVL/g6DH6jzBZcspmumZhEk4HufB1made4Y
7JNG6ISPGDmUCZiNdcjy8LEnq3miFBxdrPNjCfVNE7PdKvWfjfQzBAefweb0/kzH
1a1eDOse2K3Ik0B1Su9qaoXzHaQ/wHBswaZtGcZB73qnOX6fTE3qUYCq2+npLUks
MoHPk7VTXrf7Dg5Nu8yQS1sbVs9r6c866pBm6b9wYF69vENXx4ek/mxA/E2kLAZh
TaaZrnmEoIJ+Y7xmDPJZaHpdz5LuN35ru12e90rHl8s1ppXDQqjeASweo6TUm1hH
lXotU12wWPmbmlaik3anHKpvb1tQhnSBrEBYWxZ2Vdt4ZzowNtvGwazjrzcXvW1L
Yh79JxOCFA/Tv5HPh72m33HGwuix3Mn2k/rrhvKkoVVI6xM8jmSs7Z7nBPaFAQEa
LL1Sd4peA1094wbviby6sAdJPlh+mtL13qlO5LbjBxz1vio7s5P1mOh0t8mM8T7D
DJ0FiA+GeV3YQUCYLbCGMOCCHd8/cLYl7ecKRfio0a0taCX1akQpn6HK1ExqdTMI
IE1O+WGSr3MzMLEdfvgs+7MJVBr5au48G3bjYcz7GfEoBQNUGJuYP+RoYz6j9t/p
Z2eQToi5zlZAQfcAGdBjDJrouGI5nEZOgkaubf/OsGtPfluLN3gEUTvuRpc3y7GN
XmD42l/JSjb9YV0u0Djqz0FNcq6GuVJLdAFJH6UOr7b5prmyjErf9/x6YSfGLlN5
4GidfWkhIuJEdunipe/A7P9XtH9/RURVm9QknQJwfI2dV1q1HTAAU94X+gWptgJh
S8WKuOP3I8c6n3VX+WleYaziaM/4ohhKSL4xVKQd7b8k9ejg+ZF5Y0zU//fhsI0L
ZKXkzRgSFS0md0REvUYCwtwChnZSp1Y2ieNefQoUQXV84iDHADJXzVUX1nLTmuCa
z75qo3XSDgL7DAfoZ9nh5LTkS7yRDvsuyVct13vxvAqiKcSC28cBPxAPE/5IrAtH
7vPEr8X+LTC+qw9u9pulgg1bNwYbbnXSGPPOGw0t7QTnTtrJvUEaDazajwqCkHqD
0KgmZ3KMtAA17pNNCj5y2O3DYLuD7aZ07NIC091CwWs10BDNf3RPhoDq8AxOP6de
WIQoObiScW8p89k+cpCDiUpKXvzXLf+8r4bQbHPY+jueUqbpPGOui4ouKKpZ3gOU
hQIiffBogfjjgw8SoRAFIqe6qqu8Sgb5aRkHkvX4NMfGLybAgthO5XeRQNzRcoUI
kl0sTIvvJJCQxlvDXuJ93/w9L4vMsAud/ItgleHEYknLr6lRzMlLZGPT8B5su3CT
/owqQhZb9iytYBnfZox6s0jDKRvah1Sy0YkYQJOFBs21rOpvuNKeD/rtX13dpvru
RaYOp82CZtV4zwemk5rvuhKKVzSUIWWgT5XCoEuwNJs=
`protect END_PROTECTED
