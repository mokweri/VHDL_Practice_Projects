`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+o1mGeq86flj0C9C5RJbM7cP1cF87licYlQNz+cYrPmI8I1NCdi6D3dJjm4POFm
yyIpopxFjQKABkle35EomRQgl8pJzbFgHGphT4402SpS3o6Hne0FX+Znsyi7VIk7
CIKz9LxNkGJ6KSIYpJDba7ZW+YgQn1gtOsa1ofmDGve46o5h53LdcGUWel/2cB9U
goZXhhvPX4DZiZurN4hdgG+DuIE5NufIUEn9hjqot2h9jGUPQSxAKamMKRaYIEuw
UYvsio0JkSc9vRDa6I3/rkKBAkx3A7z23qvZQYS0jkvFPa9zAIDuw8gm0CrANkZX
sHobQtfz8GZWXtuQdEiXZDJZdODE3mcDmQADB1pIcK2aP7NxiyXC+uKEK2mRC0dj
V+WenR4SiJZMuqlQ1Btq6u/LEOyT/u41gddjsny6HAccQ68mIShRylnHU8+pmMAT
XUMXbSI42ZnaMwQccnD7F0yyJyOVoaE26i73u/ZU7R16jJw+tsmfAr0XFte1Uixq
m5HRzqr0R7tjyvZaVReYFT9+BA9Th8CnqLEobR3EF1I=
`protect END_PROTECTED
