`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BLXBUpu63r1nhaLRqjl/XGi3wonx+4zdlwFjwIv8inqWn49ruAZKZTT1yNPdWSHU
3J2czUhAf8QsnB/HIJ6FdnTIObVNmnl0OPhKpQCDEDuQ9NoqJvEvAF8Ljm4cy/q5
iJnldSyvZ23ctQh6LcY3/OAHrDcKDOp1tBkiZ5wH3pIW5/Pt1z16bsLSVvAPqD+f
QeJYS7KldlZ8RQtHfe65o+CFpgdbsSF6Zh7W7S2zIBADjeyT6/W/aduI9o5UBCae
NwQH6JXvOFSeUKh3FLRkm2TK+0lACunj7rojjxLmb4ArwLk23X95BZx4yue6xZPX
JlNj/3Uv4ysxQttXLMnyKIHDswoD9oYEHbFiz5PNPiLKa7MWZK7VM72HC8/FjcjW
Dxji7/ADyHrD+mYjXyqJlQ/88gt+hQueboIJ5xd5D5BOKzRDjp3ZeqnzpxyPrZGU
kq2UkB0xoqWTusxk/Th55v+DEK6tocPuUOyy5qUmYz20N2Z6y2o6Ps8/17MrgXyx
kDc9Q6ty7ZhxeOVEw9MV+lxFdIDmOSIQb1zDy9834NtjiQXUg9uYTLOqL0hVNWpn
Qwzk6Rw39/LGcz8d+cEQHzCzaEk2rGy3aq2ueRQgcTwoylgfsgVFTZgfXSXQjKmd
lJaUmJRrDEIilPCrcx5ip9Ifp23UmTHtEzJzT61pV/XNaHa0Iq2MD/hqVSPGx3xV
6HzH2TThpiFEdPsezHEKUSMGByuNaVSoUQRyoUWRr2anZG1Y0IMCAKLgU/G8/JKC
uFe7FpKrIWniTw5SJ1Jr5iq+/pzXmSg5NB5YCGL7QXi9Ewuj1gE+DA6NOJvzgRnK
7vM9vX4s/L+p1DV0C+sAIrTH43iP/y7g6TVYkcz2UsyjVzRdNCHMF3OhlkuVyBzt
Zg1q3swv9mJWoMD4Y575WgGJPgnV9ml05/I6GUZgUtsVdIC/D4ZJGoFpc2L6EyoP
rFbQ2o9ITwFnh2o/tZMrfsh7SbFWct9lFoEqSLE0m1MxrciEFQKG1mdYPdFldqN5
DwtJIsiEnhbwT/9hEwnQ95iwRaNNx/yIg3vEC2gtfah0CkktXfjWwL7OcIgxdq3N
DmfOzchp3uCLDS9IUDFxErkaJgoJxyU8hBDdgIZjueSW+HCb/NZ+BEv1Eqc0wTX+
u29tPNu5R2EfORY34uPdA/gYmr3VsqYqhlM0XHf4u7duIjn5q4AzIwh60djRtV7o
l2etyU8Rtiom6PI6KDP3+scr6KnMC36pERl1OZIHZ1FZRYi13PpPoa8zc86GkJVT
Q1BTcPykFLwtckWvq1uUs3GSgYtrLT3zPKh1maFF9jmgHnvqvjR/aB97vQK1GwFc
seGmRj1y+NlO830UV7QPHO8j7KWuzCwmSWz6weLiNwFhDskr+NLXSgqnFoGTYVTN
bUiYY2fEnJ5HHn8jtoIJFzCipF4kCCgMgOju5MbbzdD8zSScAj4IJb3T0Z0ptJw4
T5XQ8GAe0grmTrwSwAq8sEhMEmrMOh53GhRERoev8GZmW3sOZbQapZ46KK0WmmDL
P/e9LZzjxaFVcRw7xSZfLreU8zfeoWqwEuRYgCesrOSq0nbTrKO4Rsx40Rb7zKOL
JFskmiHR8ynZ6WusXIPdEcAfS3pQqvrx0eCa7fOqzXlWoN0Livuc+4EjTxeSljvX
E8RZDDBc6Jlm0q+16f9OQuxhRgQYdae4yD6yMb7Ct5NJu+N5BFoR39nABG8XLgZA
OcLcn0tXPQTxp2Mo/H5URe/WPRTkT5Xi18Oni5LyLq9WmQpgXvMdk7cfkQK9e0Gt
WJOVIrKcsnjXRvSMcMq+9c0TQetE95gOA6yNa97rDTiUjZlGyPc1IwK7tv5Y1eTy
CPhCdIHKhLuL6rku+Tod+UwKVUefklwSiWT3qG/UcFl/BhfqyjfwuCCIxmyRNDy5
g5uUKPQ909W+AmVnl/7LzmMZKJz/BMvtaTOlbbj0vl+uL9BEpZIaQ3MLzrbEpVUn
pYTy9zJGdgGz0t97sZEHHEWUSUvjlQGoJRcNSdXIsnT8XS96Gz7dVwo+w42vKhWJ
oCiZx26oNnrFkHf3ElP8Owjnr+tIDmkoyspBERkPwErzxjlARLZ+LNoKiNTi6Sb9
BBoh85xIgpdJTTkAFzu4KBu6VbI9y65C6G0lsiWU80zk48gMgnwwCer2zqvn/e6G
HHPM2SgGuvyHSWO1C/DWm8MvCDwsJAGo4jgZ+bqnQ9EGhAxMVhc4xYAR4+kgA3zp
dA1zwwt/P2e5+uCkd3wMmR2nGLN2twG/ndVijpyiyU7rEDe4vNQQvkNdydX1nWMe
L0zs0krMmzO376795LCiP1HuJVko5HFxYoPXKdIgSFZOAbNN7BhldRrvJgnxFKfp
qkR6LyxUUm8SrviX6HqqlNk5uiswzYClVBvfqVTadnuttze+b1xpfrF1p5vNZnUL
QSehraYTrRFyHDtxHrRmOL4A8o63PoIS0DFm0i/EYVIQPGB4wVLoJmZfWHUUf0XW
Bpw57WyOREwQpFWazjB+f9O+n60385TzXwU8rUOqRwF9c4mgaCr7UkR2C77voxFL
5e/iCHeyN31N0PY7erdh+RzMsZ1Rm/MQo9MvDJQbtyMsNV8cFCBgG6wzo4AVi27U
+N3U0MSioiEqOrXUH46fvPehUF7sE7GBG8nW9f+1Vrm1Lfj5dCmGfp9aR8KNjFfg
1nXuQiq4uqgvJ3APLfYSr09WBFo1S6qBFe0KZIrnEoppln/OPjpCSwYW167utw43
wMTbj0BuiODpvy6VWvzZ5yUYyC953OE7p79CYwfVJv/fEeXM51d2gZKp4hXDZS7n
La/gwahdob/DuAn2XA/PVHUQIIpAy0OGpBfLxN42/jugwtFTduqOtti1L3ukYaQx
K/T5pumcCz17fWjj9X8GL4iktRlXc3J8xSPX4a23v29tOUmbuUaOZfC7NuH0OdnV
BvFL+mCu32YsD83aOhUyu/MVGsx+XgZctb/024lVAYwMyMQx+TUDtlMLGlUKD4tm
7GUHCJa721lTufqKIfK19nW4IcAwPJfuKumhF/rQB4qP/ypmPFcHFQ2mwykwMVyw
YR5DGIcfiqdpe+TKtE2/fEExagV0OzNsDpgDZd9SvkQ/Tj9wXtzvou2/mjtIPbhK
DY42u98hCe5LVfmhzyVKhIOyHAn1xNeqKESNz4agG27OhdZGmu4qHczdR5wXatMG
STkFskRkEybNkVrBbFtjfCQdQx0CmzNHuo2kw5z11WUKubd0mw7XwPDlCKn+itA8
TJWht121Y7pCKUaN1mNJkc1cO+dAU+GF6y5ZQjGwI/REsOZLeoew9iY9Ob48rosj
DJwM/o5Eo3sbbQL1RFz1t4fcCT4hwA3WB8GHX6SLqIy9XLeeB1cZYDKx9JL329mY
1U3g4gUO6DN6M8Wg5Lz2tZzRZ1tmjaHOxsM5nBpbN271+g0DoGS4g8oiJNb2jgXE
7adEjQXb+jfU2t16uxaiir2H2d1FiG8JKlSAq4MNUhXRcfTM/fx/x1x93dpXQkN/
G0BA7TUZzjLdKMpB9YuJvdOd1F+3FL9yI+5Rg8dzffYDZfsuQFG+r+Z2guue6NrU
eAyRwIXfJaX2DR58HdjLx/jKUerwr368N2U30raN7x8v/4Y+3D4YSfks1/YfACw8
EsHmbn1zfWDvnIgqFvrE5U4/vjmW0v2cCYwEC9Mbgy3qbXBl2xbiA0UUdHiI4rm3
d/5XSHJaVS/BKSAc4I83Lih5L/wa/vPSy48gUWDL5C0SXld+73M55HLYclpGCh7+
1epRlllcLvNkDD35nrCO/ToCvN4MGkkN/0QRdBAFjbgU+aNVsGLCkYZOO/U+G+qL
D2IyAjvTaXp1h/Hly1WctVfLuIYzeKetjGsuMWtdIFYklMqIPnYNYi5Kdx6Ta+z6
btI+qhuz9nJF27q/h8F0vRFR39xu4lFFK/uSQoQHI3zo9acH90+Inpblqb1gS5od
VOo4X4mGHa7AgrWgCfBUrO+91Ge5NjuGK8swc5RDZoMA+iHBei+KdHCYpo/JzQ61
eWsciVY4wwzi6SVB4yOPPZmVS2WSv+LgtIDBrmrlHw4hT9zC3EhUVxRBKaga4k49
esnFyDIH6ujgcfSRUvsugDmI3SVg40J5T2InO6U9+zT26xXkcDpUAISmhutk22sK
jxlVg9cz6dTQ6WsQW39rvcJuAIyQH+OPiPA70+KqzKgz0IIOFVHoflj0DWG5nktv
Ea2OS0BPr0xMIQS7X8qDr22AmhL1Ab/tNBZGiODnD8UiQ0S2pV083Ew2VwPY3ked
2ZMS2H8yevmUVJw8KJjOF7G+Ble8dXYBJnAyb9CPYIS9KbTudXpgOKxVfkTruCQg
MONxPMqk+OG+sQPxPtMyplySMvYEuPu1/M74xP8DBfIVaTivpCVz9kGvkSt5KxMR
LJiwQ2f0ilodMJBo+2HMRi0T7aorzX8T9V8lfTIZYkbA1dywItIkkMjJ7cYzaycQ
FvsDpZuoSdBj0pEsX/XqzFhD0Ofnl3xVXbg1RK9h9tLoNEabXcsKW2bsGfScvUJT
eyZVWAAhgigBsUwYPm5f/GVqsw/IZOrsWUxdMBb0j4DyQWOlvzRkJE43f3ntuC98
Ri4n7eIZbKzMGSue5ZPli82QzXR2gGXg1I1eMMznH3+abKqiAFvifpg9I4+JBuGf
ZX48Z2ar420kSSGPW8uJAQd/4fYUnZewG1i6U988jncnAxxmPNPxqoVHCNjt4YKY
22lViTrGc5q+zwfbRnFVAxGDw3aFHeBaaTyQ/kRiB5lpLTVUJuOX7iruogaksqNE
kIOhj/YS1NASNrHhZ7rRFAZgW+8lvjqrMd7opvEo6G2z3KaLiN7A4W1eE9CPUBBu
ADgdOzht9ctmf1bj1oEoMZT7lCcrcuXfJh0j9grsNOG2ZYX8gaSpmQXU1392d7qa
8cg1rUO03ou6PGMZUYa+XmSsHGp55XDcMJtq7GOPKBtXk0IgIdUMGQYkwvjlS7O3
j8+Q8grGw9tXMCc4yeUc9bAfQkZ6WJzRcEADkkf1XPi2uVlOHCtIIqXMFlH0WTMR
Spe+ZXiHpgE9vVMigAgtdslXwRUEHGfDEImink3XR4twlFvXHN61eL2UVdI8tcvT
s7vY9U335Liyc/briUHMjxvd/o+8YSXUmpK1MK4hlNP/9+MmZMBILPyZUDY21RCB
FR4XxLnpELBc++N8nnlitGq0e9pBacKKDVRR/6Ykj2ZCXn99Ebk9oglSoWxyTrkr
uRtqF/jrBmEhphncZKazC+0ggCp/ZWXnZnhMKrw3cerXp/x3TnAdejI9+u6BfOL6
4iG+YT44tG5HmyhEv0NhNa4OiIhah3XxcORkwDnxpAvxnUi2Duob2jBIlXY2oVg2
j8fqHPJ3Rvxe8tuHQQgQIE045d0AxnhSzQREkBF+Gm0pHtdjVempX+pYIEH27BR3
Jv7whSvdoGZrvWg0olmnpk1hxV77BtsQLxL/1LX54E5uIHi9tPQnUbOr6W1ZP2pr
srhU2nz6ThRCUm/CxGzRPf1Byo55t8OSmvVEjYYWcNTn0O/8JYd0me1SZ5zH+gc1
Lus8I+UD5f3DHJJ3HWR5doO17KcDBkb+KKN+zFNnWfaUi4eX28jwWAcsEKo8pvvY
VUJqMNjt3owukqMkciBFX9WNBf+xLRYm30TrP+RTvydvk/QipyDTrIP3LunIPZkc
iuj0zgF5HPrAHpC2/S0IsSwltVtSFCsFcewiqVSbcnHqPnv/vvocBN57TlzxOqab
mlLkOqc0zhgX3JXS7I1nLzQymXinuV3fU2Dc/cMiiY4CKYOOfTuFXyuFhiWmR9RL
n/I7xgWoCrqh1kqnY5yCz8sEMLn0Eof2JOc/tnUmBNx0H2UTHtXM5x/cLrTaE4F6
8Y5Kz4EvBw6qgiF7djCj/GW9RJrrJoEo4NZ6XCnfG4lSgzfVeLfE9axVkpbqkQbe
YDoTK/O6yb1RSAkLpE6orsiD/Qqgb/V8RKK/yqYTbvBY1YWyJdF6WMqLvjSrbFrM
2prK6s1wBLcjh25MvOabRR64xibhmTr7p2Cajk7t6EBiSylGsR5QMbAIQCsd3Arl
tvzZ2U4IaN9rjvshACcBhrdkuGYUdraIT9gGiaWaf2Ismj45H8/N4lraQdTSLxac
CS63xoMDnDhwXlUlOKPSzgPDknudQxplAK2UcifMJHxXLpIBQSJqP0InjuJG0lU4
4O/epJHw8cmMoO8dbwa4kfSV/uGnDBeeZVONpUr4bx+JfS95WoQ7trsrIe10c+x2
bHmTUpbDyv/wy9GACDbj/rr7abmoWPiHDrnqqrWjL59iBzdQsPucP5W5QNAF5Egi
KockXXhyiPX/0bDvmUaknIViIiQwnYS+Z9D8C/3Q22AzChTNRQtjaBnUFqWVzjKi
ZXFvNW5gA7Dl6eqKkkYJPGVCz0lIIHeR/R0pOux5YiP+Tod7ZSulqVUfF3Cz84tR
fJ6sVEZEBOHNO9qqjPktZ3lXrs3RrR78WtGd6CsbwzSlIeqIeDC68i3LvJurZfQ7
AEcdYx7Ljm8I5TXIKDu/1eKqDhwyT6Ry36s1uirlTaZd/kIubwr6SwF7oKJLk1F4
/em/I0JWSf0s6Dcj5nqITtb3aFebCnNOE0QUfV+Q4JQ6hYOVUj9L3jUMnZmKi0QO
Qzxbk2p9MqCQTTYG2lOmxA91DerTgVmF4ElEgdxUgA5IZuI0tPbMeimfJOsoJxP1
x34dbG49etnfhRG/csu6BXnQbzIZ6q/KI05eQ92wKG8L4fvSL8gEPBHrF74cgkV7
CLqpmx1FHYKyOAbGljpk5QPPYvxpRgxl/iz/GCScj9G2E/20UkQk4eBSPlLJ0fge
ai0rCbEmoyrgHLkZSVwQAx6zmGdl/Ykn+hL6jpl8ZeqC2ype6ik7HIXO65HEedNC
rM+dLKDjrittPOb9h7bqTX3OarPbcWr/apvW1ZsXJVWLIdy+cbhjvceCNTo+6lrC
HMuU+Uxeoz3hMzksPhRIhJtmqdQakzEq6smkZjReDYUdBExfJtbvYO9FSfM8Nk0y
W+vbSnJvLkUBjlTFBJZqyETm8fTCUm+ygAGrtvvFI3ZepFmGh8iHceR6YxOnxjaN
nC7j4pro8QM3bhNOMjNzVf+IXSZGK6dxyi5AaEAkKZbdoe3TNigbxAL/xFdvRU4J
Z6HBwhbJhiT36Cw9lHGBhCh/bTecy99XChF7taYwUpz3UJpVgHqkgAiAMm97EUIK
EI1PRZr9nbp/U1VZEAs21d9jhkx6LhIrUghIaCd0Fm9+4E6ecWFAtRJpEpv/v1P2
c5czbtKyP7jAhY0MbmX/dOzx4DQyPgLrYeuSYh0AxBVfQvhDs+7NrtBb9OhbVH1y
1h84K+jwgy0IajmROexNuIhu+ukj8PHyqCGLprYUFHiJVIx9iItn5Wz+06x7vLD+
0glMSaWWZFAic+7QDBmWkoLEO4fg1KgobBlIjkJIA3/I6Abqv3+6O2oWqsyJafEm
kEzcjkZ96IO4n6cKjIpquCAwyXuKCt55n3zHD7GDWo0n4Rb60YzUHYnPm1LIPiYM
8EuRXFISXyGiAkU73BiekNg7YPf/7HZVFxcPYv17zUXtWloPue9r0L8iL1Dx/PPn
eNAeC8iqfXATisUdTA3L1X6erpztuPMilcUCkZEPyqFsg2jem/DDfJypaAtynGDT
Uk01AGdNmiQVtO5bSaQf3ESatGH03kLvr4wMEtgBeYEFGR3UFmuZ711DOr0cPxlC
PhY3Ew9jXbX7s5EBrA60R/pKCyFU8v5VtOgazg/MmEKh+FAdGuYGjO+BA96KS+mI
egpf6yxQ1oV2DldE9je8VBlZlB3pqoP4z0m51mhyqmK+/ihjUOjL+AOvrIoE/Vl5
E0iDk67ki0QrSsq03ZH5PH/qiHqSilg6fUxSas5jmS9zNfxG8lbJNZhyoYw2PA0s
WerVJLrK+SAcvRtCeOZYeiyTsWB5/XBcdjqr17KmRMJ1L9cDLs0BXL1jUNuCkKUs
o5dygr1U2YQpkUn4VZTkWq3ikxsMHDTMLjbuBxAZUDP/U1MWOgcpSy8BKIWWA8Eu
M+CYXsc1b4f+Xu2u/s8xsx0deQMhOdbOWiRom3zNgLuQBrjLS0pTT8xAbgVfqM/G
jOx+zuo0qKItIIrGQCp4NULOF550kGk8YAQgSupf4hDX+Jd+xpO1OyBERROLmHtx
MBd0JXq61AI44EEPMIoASCdAz+r8vdrdmAvA1wA3kRQfbcaGltwF2LCX6IUFzdZb
veI/LQ3fUS0J5QmbxZwfboivqDRLco5eN68i/NioLNAes2DkDC2RUYwTFPKFAQNW
TrkzIc+1NcLEExk8732iXtyGIdFLv0GPcijLfkhw2EViTES9vr9aCArQDroe7TVn
Wbk2y6WYC3pYmIcVIdXe7Yq1SM+Rc1O4SxfpGxpWuDcK651aI5AN/MVPGV8fgwT8
7eGL3kwhJSc4lHzYHH1a5LmbVvYIAFo+bIUjhPUxGnT5EBM2UVXErH7D2RFBIINz
1k9nhDSxdYpOooUu7hIVPFdMi+2ElQcZtT+8kOVYdHvVf2+V0uBeHg+kI1vHtvLx
CNoOPo9sp5WeQ1h66xChPfMjuLhd8ZT71nBzRE1u5OHN50pURkhdc9Emnq0/HEco
V8y9NY7IgwhxhX8t1/wKOF3Htf/i99cWkz1zhaAMZWr/VoKAdjpL49sHeOmboK2w
Jru1GRxg2uVaJS95CWwHCM+RX4teI2jaGT3lbgEl/gtict+q3unxZRJAJtPZ52uN
HCihDYv3RdsVVnZbbtUlhcJCeys95F0dvYfK1USXDbiYQJKLARJ+icTlZK8AEZRP
6SSqvrDGnTz5iUISfzOXnjiua0kLxm5pjncnis2iO2XhnzCmumvE7+ZrjEjSfFWw
AQ5RrJO7yohcmrgzpWukPgZQ7myPUtYuShvLJ/RrOM1T86DXLRjiyLdorilPdYhB
t3iVL67e0Bk7m7pqArwE9jbHgLV71UURrOnBEBkCMI5dRC62eEV1PMsPWLzYFLns
O989MsnZpX/6fOf5gScHLdzJdjbeROjbH94AYTFuR0t3xst9IOs24drypraXNDG/
wUYhheR89MRCrfQKythc8PdmliSqg31UA1WuAamVkQ82NKyOOvvObVO4npc1qEDE
10kXYAt2OnTri84CeTnA49fkOK1uoUrynSQ3DCD0vw2S/zf03lP+UXRSV/lyKqnx
ss+O/qao5/wAVvtTgKwyb/OtqqBV+/OW/R47HC0Cy1iCFsLi4vVifB0L1ebF6iie
P+Mj2x/7B7Cd7wNmJGRTx/rEGVf2aOVNFOQun0vnBwy7gpS51YoXdMuJ7svv9njv
5rtlKnefwzHyqC2aZcUZfUiGPY9Fakc+i5uEmfQ4D57z0WPpIep4SAQNFy9lbRqR
GNSb/m4WSv/8B0KaCa+RdfD3rYAI0YEu04M/He97BaVPuqNVQIc+L/MQ9vjMPZet
MwREUVdCi6c8rB+FF+ba3O+Ra/pJ9dMBVIdeXNPc/00ROGZcpXK/+oEf+SoAmbTB
PyIRQdUNdit6s9n9g0aQTwYLx98mOgCpQJaImaNUUYma8qnIbYaU8uPT6/JRbIff
4sw6TQf0gJ70jNnPZDG5FFsYetNyYQPBTEKeHr/H4+QzQWymb+5KD1HDvtl1+ogg
BBMH8eSvFCvg07GKEf6IPT3sgedLvNsQ4yPfH7C3hz+R35i0Z/WfEeALxYkaiZqr
1bQ+8tKRN8kMIEZRlAgrjvJgqvkYU1pkkwrOB3lxRPmJNvHNnHyM91Nds3TI3NeZ
Bjo0BFS+NG78a/4P5vGujODgwykAOE16/+d3Eyz3s971JoKOSvUi+tIzf/CeOtYD
H5Joo/RnIltCJl0AYmmRRGVnHD3bOF4gEt4T1XSFwJJjgyY7L0lfPINJipnIHDYe
xJKQsqPd8f8xxdi4E4DBvpLqLEvzZ7nC2UYbRndoxdUmDE/ek/bIEuTRuOUFx9G8
eQq/kFFkh5iY0W/8VVFlEyHAXJwTQIXgPHQ5C0S+AeKTelAjVjYkjGTUTHmxqiz/
aHvxkvHx1NHVouwsrmPcbAdLhecuXLC7ZBV9Rp8q2z+vHdNePLeo29lCHImsAlxq
9+Fr2Ne8Ql0/aI/GVDENgCldkbP6l92HidSeIlV1ULhL7feju6z17Ez81geuG3nG
LMd2GgF0NEiR36ZUtE6BAVOghvV3P+8evgerREdbX07lONPqO+gtbDrzOmwB7VsS
LXOfMQCYsXrwl880jTkEP1tqqcdQhY0NcQAWfBfB0JDPTN83uyo1R2jN06/pX2cb
VIHkqFcWWQfRxpKjPmYPp7OL5AQAn0PhQROWfBeVcmCkt+AM78LVYGhzDMwFpNp1
4VMPXA5iCA/RW+a5LxU+6RRfnCXActNTHWPV0aIV8WadqtMoXFYb0sIZOCM91c5j
YkA2macRpSG0EIStMruSo1lt3PZcZxgSFC3HGO4iiFYSOYfGuI/2gJ0ViN+fZQuR
JrEk1dNo/6kQ6dR8VcT2ae6tLXgUcYss3WDLgn/24gphdt1XZQMdYIVGs4E1zi8g
5B0j5a/sJY7DQggMwaMHmQ1DVaJ2rOTqwHPnbAQyoxdOFhnsJxiSJCOOlJBk3BJD
A+YiGMPSu59aHOPRpWNia0IoWLrYwCCtSXgmw5IkcOJfInXdA/7Y6pd05E78g3Qa
uZarK2seTTiqfa0hOKr+uB8X9spmCTgQteOmDfk3X+x8VKreczkXrghcVa11rFZT
rsP3D/T6EFBZwVXK/qtavlwZrywLMpK1V9486LOp17+LzfxafLrzlyKbngTrXjJN
C7kS30dYA/nZanvmgCSRf3s1maVqOt8SqaJrAFvDNRMVUY3CEfU6hf1nIFR4AHqb
Bv2u6NegwZpqX6IXbs3HH0xqGKc72F5o544FbuKgMT5cQLEXuD2w58W1G55IWwPB
KFRJhfwXeozqn2H/Blz1hNjQM1OYADw8/NxgtcpkBL7El4bXW9/1MUK1mUDcQRNI
Pp2+5yoz9BiXbC1z3FwQwSdodl3WYBFOO8/GTMFdQYeMc1CCGhSn48r1RNQRZ+t7
RmEOinRAejbybJrrhubns3QMGr4XO98xLiLMd79z/rqd0WflfXZpQOcjydiyMdRs
OHh+zbJKq4UTXTw1NIzW6tnxf0VAACnXtG7ieq4ImRw91d1fctXUgiO9196U7vOt
YZq/JSwVCP0sVOjmz00Bb8TU3hQmNb0XffF+nfxeywl5SqJbDoHmHx46peW+9fwn
4spZzGqegX/TpOs+xzKLpFnk5vigm0O1xCZG0OKcky7Y/WUzCXnMjWzey9SnAUFY
vSGRFYSJEsUXQopMhvaAkxkfujdLUQZsUmVcPHvAjfqW8g+KrUKN5YGgQaRjn11g
8RXWZE71gBzc7FfaJNHKjUqAkG5hFeMNbxKhnwVFZjkbCsVhoX2dr5HGDUQyhoz3
enH79IwmIt6tSt+wwyPHmikVbM0W6K+49x/L785HZ1GFZAcpY3lmGhNOhtOR2PEI
M06KMHjR5gDnMzXNJ3BnnNHMWWE91P3j4il60l3bwPM+ZIR8tMHQhAlla9/Cr1d9
RcEIW3JGLBa0pY1e4lL81d6aQ/AH6TebuKbFGwmQ1ZuEJlVjRqv+dH8Nr0TXirjp
tPSaMZepZsy+WhUIqNk4rnBD8v553LpoA22M7uGf88lh5ZPYihVA3zD9fsFASnZk
hqnUn708ETsKjWhsR9uPBVg9UKG9ziUPjBG0S//CMiuCL0dZhtx6auyknbXMaBR0
u9PE+B3xbevtr9MAq9i7gkPFZplwQNwcGHifn/3g27YtVtXAoYWVRAtPwds/VHNA
DogXr4M10w+u2TB4X+DztUqqihJiNUlIZh/Ldz0763kWL8r+mxuV0YGI5Ax8vhdK
Poh+th2WsRwm01cFbq7X/R31n7VZ9GyxrQFI+APEyf0onmIwmEjynYxUTNYkNTLe
Jx1MjhUgWnYQg8a5+Y7Ya8Vl45dnt/LwkG1ipAdd29xp1Xo66HJUEGOTWWz7t1A1
o4Y1CpF98YRrOfSxruunaGennZoeUreshReU3PQtLupoj4nzZnppK3pUom4I5oKE
l34dT+8v5S3GLd5AyQDGMVfFJ6y4sauOWUTc+0YD9KmMfK2/C6GDs0YeCNkgBNkG
DZqmlVCnV1AjIpUAh1ZHbJMv5KWD2sn+qgmXorei6xmj6oO82BEH6ArG15/ULc3h
eEltyXAgXumTa6LgNm6UwEmVXsM5Cq+F/FWahvnJEWh3cDc+IE17U+6ppCGU9daP
LXawrzhSWK8Aa0dEZMgPFM2vP72+XN3B2F7pSZqhdVX6gdMJzn5j4mlTHfS+2wXV
raYa5Y+P2Q2TMV/xR4eYayedyarKIP4Yzx7dd0yMhHv1YacPVDXIATf/CbeaecaM
CqDD+Uv3fbzwt1IepYEXchqofiWyn5qBpapqSRIbB2mPH5u7x6BpCnkdyKdho2Bq
X+IY2zTMHWfqNlaJwGtlHWO0sbeBmoWp1Qylsfdk5BEB7aJRG803cRS39+bG/qRu
5z9XeRV4lMKtG9Ibi4M/W0vog+9gZDPM9KtUTEzW1gauk2dyTJi5saGM7sGZtH9z
J4IFGJdSs9ouMsKJ8f8feVKUPs7A/2hz34Ogz+aLFwwH3lD8NdUVzAsPkq2TsPpE
wXu4kvxQgDQb4X78b8uidGXM1D0jVcaan6Cb6fl+CzHTNCjrV/ZhcdhN5ENaN+Ar
FPuM205J6lZOSKU9jGGGfTcPy2XkcF6sGRLo9aeju2PYnMAPtQa0GheQgu0yq91q
rBZzU/KxzHlDWGNSREkK4p0YJs8bpOnEOBt3MteKVdxGbdZGxTsreaJ43tqgMebY
78GXM8m1/vTvMr3gE1tQ0vtNKsBZqjHjZeEVcnjc4WabI1JRzMAk9wgtVy0CuE0b
R5b1gcmiETqBiWmbbSBTWNUHVWvH3LdcepkiEovc/Vv7WEAVlAGh8h0hhB/TgdR3
brS4nU/sOQzNGh/jwh6VSwaxwZtJNVheQzJgw3Tma9q3ByTDwMKf6Ol09toiSMBU
44SgshalCQ+XTizLutgESOxSm3cU2NwjxXjwOFRr+DbUfGIEqoSbXUE8pDxnbLgh
XWKDIhQYXQlK4ItQCILT9kl54saLpQSRhCsLJukTLWBRUn81zS8dpyY1oWrtNq+R
vXstNAR9ngMh3uJY46JPbEVxkkadif0PWyogR2jg3H7jZLXlrcb5HVt1Ql2/kerr
F7kfJKglPPMfN204TpukyeTqRt0PDO9O3GCtCxujAfxcvFnOJNFeL4WauQt6aW/D
/KhJNoxYdMAfEHSHStYoxcFEQApx/W/XCK9Og7/RPIjcQEjhv3QtRyWH2S4hhaaS
OCrYcfLMn7Uv+6jlNHtoHoxqLweXErMUUWefRAlxW8jOtvhKWX8cIyCZbyivCysy
tVxBxO1lzTArAGZ3Ac3ZCjyk5pjH+n+JEWP3kRYiOBSs6BvpVtDBq8Oq4zUK/MMS
zwRmQHFzLGU9U0cZstDXkrt7LZyD2fMjpeshowIYjir3hAiXULav5vGMxdHYmt09
We87FZmu5dX+pXUS+Z0GvwdjSswnoTJh8nF6j7y40NbvvTf6HKFAKU3mRN1FL+pN
ynJG970aPmupyjgqZJmm6p/PStcGWEzSUF7L0JRBAPGtbCSkYrHNLe2iIKki6MV+
3UA0LznTe23utIAt66YSVDg++Lr062g4XID9+l/jlfhmu91VHeAKfRLfh4+nXpXW
OagbRU4OJSIVqCgOnTsWk6gRO6ao1gkla08mYoHAmCfTF7W+WWszIkUNy8vj843X
X0smIIYAR7H6atxR5M0nGO4yUpukzWk8Gb8e674VQ0WOa9PMDpaEC2OH6Fii1Ud7
TUsguleMKNg250YaW9DdUe02gwc6KbiuOgKjlZBwytl9saqxW9Hq7Gb8mOX14r+F
lComho30QF6R3enx48RmJ1HGhrN8WjGnwQmGU9tKimyE/iepVTb5zI1K51DMh/dr
OpPJGlWsGgtCUV/nvGOaWQit8KkB8lwLnjlyueEpq4QbskOrtWF/92IWsW0tXyLj
ni27Z+w+jEXIkmbllI8zARtx/KG8fyQ3pr5oM+DVr98UTjNIbUQGM54moirIcbZ2
Z4hsnIA5mEF2j+PVNJfl0AVx5nTYsUbj+Kmqa4T44m4B5LWEZrERf7wtjm39n1RS
KkNgBK1O27aku/cQyrs+yB//b7culOnXkCE2MaTHBczUvR+JCt3iiQjarHUsrtjx
X22jmgYvIFi1zgR8Ggz6j5EpP0p6eI7Sy3qqaXadTftJ3eznI2/+cgCJ59pm39A3
d8yq2fpIx4BWH5+vp+uLaunyZ0RWGbvBjSkLj03pirlyF9nuJlBQQp9rOnnTr7Fn
smPeRv1zOp4+CbJJywMskHTnGKJP/XwfRFNWQjvv1vkYR7rthJ2/FdtgunaoMYPV
F4afDwgXMsiNfihYLTD5QZZkndmOOXM3LTOfMgh4gFoIN27VTDsFK+jj56Prq8qZ
cdlu7JwiXJSgTOSy33aRhLNYVF78qwqgmmOR7MvcSh6nEeYkIE844kCG98sQNGjs
FItLuAsSinLM2SRud/6Ed4LhnMqZgLIAPvQOmklOWXuXv1B7gk8J4cZB4PNNgCoz
Ee7Ip+YiJfgC8QO8HlBhGAzO1RsKS9oZtoA5FvB6heqM2lrNdTDGOW2IuWOg2eWv
5k/KEzpIrgx8bUvs2qOWUQcShZaRfQxB45ZEoJqRKYxtcUUy3xnkjL0Va0CNhffD
Ajo3J9NOyyH1lwPLVbLJns5J9AntIK2smCCuPOQwdruMRNdNVYmVhLCeoxVf2rRE
QIQcK8qGlgLVazsismS7qQSh/t3z7Yshz5VXIq9uOMOVIZeZO3B6OMC6zbpzRIh6
gVlc6DsZXx7nc+o6DsgiwgJY14fAT2e5z133DKjk8/ttJHHsphJ/O7+MIawdxvgu
HSzHq6r8V/LhzS6zoRo5CRd0sD4f4ux3uRYLOWX2JGoknLSVPBTT8iVAwEKoAuUR
LRLbWLq+9Hm8EnQDPs5stPxPTwzLpBSh3MU2eTql3bRjndUBb3/J9WUgFjhaNhc/
l9j5h1Fuc+gvZN9egVMb9G/sKDoG5jS0OO/06LLwm/w4NJVVBs2hyxZ3NLMXMsak
J3+4zy04zIzoCQgS1YAUhzKLgX5nu6mFUPr+5aJr4OZaS7Ezm6IECPbs5tX8rEa+
V/IUaORmu0VBPNOY/jjWkGMdw4g6VGLN+++sMBWOyjkZUhScUP4kWsqDZKDgMWnA
otnW3pq4iU82/qHD6oHK8bq+pJtbkk4vnqP/5VArPWQxZfFOXf0h1muUqTLflRr7
oqJ8AlPpcRoSk/2zqznA5+WcTk+pHKVjLuDIWfZYTu/v8dEqki7ObKmKujb1UL+x
qDLjE0dviWluJ8mQhQHsbpQxRfxLcZsliibDGE88bCja7tR7DTFh4vHME/JyJyV4
bbJraHel17+TLbtcIs+mVrlNks2hoxgkHmXfnMERmSnCA/AGOb/hh2p3kFYDMDuX
lW3X4XqrywKkWNTD2jwIEMkaJ40hkFcKFjPMZWAOoTQddLVEvtgy3L6RL/nCJd1b
tKdR3WaW2GJKYIHCY/TineKbV3WukV766827bVGuKadadKxFYhlkOeZ7L3b3NjSE
fB+KCj5R4uj8qiA8AK18VimUnn9x6g30Djlyj4FEg0i/RKu+R1lJSTEZ8UuVuRdc
gNfImIMlGlH71ZnH5byR6BIbEMPoezxQRmuUKoaXg+L9Z6HnBuZKp1+QbKq3jpB6
Mc1v8jxAquyEr6wfmM8BlzRSzDyar0oSpZgxwytyMROxXArF7NCq9XTxmaX4zPCS
9ZWFZnm24x2dLvSLvOSDYE0tZ3sX87Gc6d1QVN/vWNa/sAjVyhOshZKXwuMQ4L1Z
QyelGb7oFKVJG9h3TioPeRrnbujhkbiqUzCwlCh32T0B89a5yBwBA6lroeykU0uj
Cqn/FwkkCKkL+OmHBN/4lkW3vs/E/k1at9vjsta/GMz76C9HNiEN3KsNc2So2knM
eI59G0t1140pndHVWb42rX3usdoWbbYIrWUYI3zsDCriEx87DRXBdZW6AYeyNMvn
EDSWd3Qi8TdL6YlvdOzeJitceCC80RQhSTneBqyKX5CSSLbsd9w5X8eowZCR4DjB
NcPdoUDVBJXwdP97HWmE8/eq5wF2XB3Q3iCzCYsna/zKMNER4xyEUEeN0OaGjQ6Q
CZ/ASy4ANLtizXTrUMkb0ysFf/4chJXgt3H6NAc/VZ9n9keYw/fWjZea3698dUkk
5M7QchaA4cgDX1WWmdJnuqBszn7CJRc62glkIeviiK/Bf3knJmoB+REolx1IC9Oe
ktVXCaBmtAWSjvXZwy+I7BDrbFquD5SPTvpoCKnk8oJoRXN8t8Lir6OgSDygc978
xLGNbaiaI+A34oGiAOquYreJ1ci712yPP9CfMaN91z9KWYMEKtsKELJT4KBlbmhV
KyiTOOMpO6y9Kz2uNNw1iwsYFjOr2UIxgGstcAgcosBdv9i47DTLdfJqxeJzcbIc
ZSyiiSxhwP6yq5RItEvHjfc2yosNboBNuYYPHXpH+DCqDm1qjv5czurW6WhR7Af5
K/FzGXDD2jmXgrLl01GDggxA2Ss+h3vO7/tlBXoJtGTvQWqfciHc39SM1n5grUq2
kpID5ZNH9VSo9bIBfOlH6wQPA0beZ81sF7D1oX3NUtUrA+B5VzHOqXi2+1ZaIBKt
vCCzYBJTMgqRfxqmTw9VAF7M6yHysMmZQDcUni9NZC+hE05ky7fcgmoSrh6uVuZa
14bxpPJ+/oZVIvM8CbfkjGBWkGY9o2QMXMHCKNKn+NWmHhgf1FqOP31We9KUvmhf
ZHREH8IavE4Cm9jFgv3K6oKBklGFsBBTwU4OwELeWxMvrHviW3XHrdxrwStFwV54
SUrR7TUZEeJqBOBSsFoqsZ/GIQ3RcvF4sxOuQ/Di6ZttS3EuaddGNBm+yokjYvEk
wQuePe009sug5+TN619OO0P0X5reWjA8J9B9ftnI9XNrIzti3zQxHL8Dv3a+P5/T
9pI9ZxuI1aJIS3cq7M1FhLDtUp1nfQFs6fXEdbaJtm2fh1aRkd3JdNsKreWY4XqS
ffw7ZXxuONq9qcKEy0+T30gWILGl4h/3VR0tHbSbArog0OX0kbkh/f1SVkTpGGpi
fWLU3NdKrljkur27KmPAQUl/vJ+8myptiGViWTlw3cmlEojHclmmT4mks/pk/ogc
PIVrXs6IYlcosIV1FUod7DW7uOpxYcO4rAtf0+SoHFTBRrb/5LPzNVC7C6VIMlTH
tQVjwDsgmk5CPDnucXOLU+e7gNnLXr2/ur7wz9cZAfTEhXw5faR23kh/5A5YgWnb
EG1gjb2+etA53pUDNH8DqPEODzhzM4XcNg/IBLUHcDKFRLPgmihGZr1pL6f7YTZm
BNv77eWvec6scey24PSSlK+p8kx984PNrBSgjZhYkJtjXkz93aGNziUoV97jLEp7
wxMZz9FvoodZQOYHhc/utdAHjRrGKYnu2GBNc9D1LcpFpjzxDAsuD1h8QW3iDE2c
FjLV3Gtr5Bewx1U3L9el50CMuSVPjgXsrFvMX5ubgraZ5iIaG1yK/kEtDO/C1mpQ
fOg4iXi7kUcPY9WfWZAf3HpYlECpUkjRsZ3Dc8A7du+ZsqZY6yoqnxvSsw5rABI9
5gKL2938hXYRtBnhejrbKYxaLbYgWufmtXkAZH54PVZLfx+aKbRaJN96kaNrA/hC
e2KyCP8MmVUl/jiTRIDktWf945C04BqzoN4G3OuwMo+ttyv7q/nKtQQDLCKX3ace
8V2RHLOOEGolBmmyd5g557XXcTZ2qRq1vHxZE6eiS6OPXuvQ4yjYZPM+fxEzeyQc
3JDLhk/xFwkyuPJe2ICaiFNy41ZEaTNPvisW3G+5M1UlQ50WwGTSM0fgT84jpJZY
FAC3vF3b3m1powT6B0mNQt5p7uFxlWSc5Hix/xS4FAVYQ7q5KlSJR9HLq8Wi5GvW
LhdzmPQIDA9x5tURHM62yISha79TnofkvlGlLdg7BC0pq+m2k+q+UJ8iuVIvSfOd
px6DxShYNmGKRNzTnTneKp2IjTjzc9IBomnx232NPjDundgNQIiZnIMioqjWKJnW
oCG1E3tM1v5DdcHKpH5SW/wD/ZUEZPQsnP74pg4ssHOLvscwv18x5YzCjUpnkD9i
DCOuamdXvmUnsQfo/N/vqPIXi06fedaUvVv0D/SZTxTFhAVQ0J4sLDW8ID/FKxHY
53o6Gv3kSxiAOfNCja8C1kudj/L+wPpLRcwM0hgKJHthF8hXgeMJ/DFJCA1mUF8S
ICotUJxLGeRkBFXg46F2AicUwuqXiG08C0hNHApmsMB9lypPZRCjR3SP1kPQvTnQ
VQXGQZGvRdJSFXOJ6ehws0cQs23qfIW7EdNormbkw561QeTrM5pwIo56axz4yYyj
pbu+nkXWkQ8eClJrt1mtCt4mHvlVmS8F7fUEjYZ27AyorgkDHmhhFnbikMnXq6IS
+p131+3JYRoYmoRwcz2zJDgPyQJMAF/db0OBt44WuSPC1FVZCzBXgWv/tNo+kLwN
XZ6y/6gptdxd4RQDnFZ9o2e+ftQxVt215uARG+IMCImYld7NhOUE9VX6L6lSwdI9
XXtFG0jUEZAgkLQwp8SepQ+sesqACNTh08ifR2pgwlLAxjYQCNFQ0KJowfbQZxhm
FkHVjRnm33fsz6mk7bDOT07vjfcBf5YT4p1MuS+cxE0l+iZsWdCPaiy8lLDfU5D0
d6/QyRtCnr4NHZNXwADq6RpP6hXo4jLW/nPTBi2Snek5r55iPzB+Ery6X1fCLyz1
aJCKZKNBR72nIch5vojKYuqnUbtS2QH2gtgZZEWNakmioUJUGWyr3lvnY20zbF8m
qANnel1HwWf350eBonbYyvD3l1JnYcYhrU0J5qwD5F2v6PyOvRQXZlyJWlS1FDwh
vkT1DkErZn1b/yyMjjw9REZxGp7XzUYfVSUulgY03NXUtzcRaGFvaE0M+nG9mIby
C/sYBYIqSOlLJLqy+k53r3w7DGGIGDJ3EKv5l6ayzi8SgDNubcxAugQMTd5afB4N
cZks1M3ft9p9Y9ycDIDqX2cv8y7ELyA2HMHB3e4h0blfqsU0Qg5WUEMbnfOk5lCj
gjIKbmmenwI4V3tcxNuZcikuT7vSd7aFz4gkewCfBvIR0VM1tTME1C6pJvRLV0aV
fAxXvns2mBEZNtdse7aKHSIUM2xKRCoSjiYqe9XLJjq0NwF39QYLTMFLGNnpJW5+
5WasY977n0E3IzGbYxOV2UOqacTgiq9ysZ/DFZDx+Do6gNlQ995SlcJv1M6zEfpA
1X8t8AtPHl+O5H9mA3jqYoMlMKPnEOFmCrcPyCkp3CXypHMtJwJWOGhMgU0e1A1R
DliuPwkkPfyQ4gAj7Y22Hgikhet4k5CTmoDOr8TZFM0Kk3P/+kkKm0V5FuDFq3+0
/sr8RrOYk3CFUYJuGXUI+QhVHrnXuiViKhAczxf0qJF8StcahFzApaxDnOMV4Cym
Ib0R/SzKyyV+zABlywGQkjk5qhb3zgyomYYiJy6ITYNQ5nIC/FC+E1AFy9l6fotU
MXIwfA6POkQM+1pudGgThhuk/STGdDoAb94xn2XqGYlkJ484lEa8aGQwbe7hRe7J
vWBTKHUA8i4FU8qvfAZIVHx99H3rZ9mtXh2uuqXSF0BpbS/UlvehKj4oYePskOLF
CsR745tfX4W7IWk9m5kVuWv9U6EwZipexK+YMPtiXcmmiRSXPlnJoIJ63eNH4Nj5
GWT1WsBou1lASfedekY6k9NAP9+FxxXu5LScuHVqbLYn5JneplttbY95yYhwyZar
1KUcbtFQOjbbd+uXCBfvDBFulTp0XW5fHLd3o38FV1qo8syJLqGWa7ixfU+46jwG
wVuf5VoGL2xNHb3t0CJj6tIqHZjhG2jX5vi183QFhD+a0Rhnx3lIBT2X3FN6Nh/6
Gh3WtGao2YQ1Oktk+W1NJ7fRTvVv2StHIA7I4DiZkHQq97KoDpsHXt/0RHTVvkx9
bniOhhzsdwU3cM478ond+Ns+ME/o6NMTsCem9/hXIxGlboAW4S53LgMwVJRBF9M3
u3tXuqVD/Bms0Mj9UaxxXzimcRVYIaib6VfBudLT+gJ4+6OeHAbX50sDDZ6azhJW
QWGru+uQiotBvhhB94m5KYgJmWDVVqifJ2apjD4f7ARZr9skEEgAAan0QBMvU0+z
nVlDDqqCh8ZlbpFB4Mn/BoMuXkTgir8bMthlfVuYyAMqyEXuJLQaSeyWelUtvOAH
aoHPi1GjO33ovDuVbbPmcXVse0EPhH72YVhfrNj5BjuBC5dRVCcBxj+O0XTg2esr
9rYdImqHGXzy27ma+I8VI720S3uQQFEoNDeZ4lVMJdnkK81XxyHzgQXDoE34UHN0
Ztr1YKGak5+R6ho/ims/WffivDJSb/BTfvKhk6D9IHbGKV4KL825vjp11E2QzIT+
Q5OaZwx2OQj0xv/Wwl8z7gXYFnItguij9GdwhzDW6UOsVpc4ER11PdbkZIz3rX0d
7zu4TFXrweGhTD93dtzWPIZd1yL9fHxE+Tp8GcjTxm4BB0rjSbdsMh68gIuqXlA/
fhvj2l2a2PUUtxVN8JE/CxRG+mtOOkgrpjJWNU5JJ0NP3TC2zaTFZB1J1OIntbxa
tksq6ksqfKuroAu0bO0/B7s8ZdNIKLzrbesXQ/akXWe1iWrDF/PeeysBi7cpotGs
VfL2EMJrV2j/5JJWBAZDCsupzms+XDqnILZNam4BDt0BsL3mu22h5upw/vFdRYsD
Jj9aeeIf8c+WCp+0AE3wSXAn4EbAjX0ehEof/y+gxNXNA8prOhcAHCNrT+h96T8F
yDmF//h6STZmAyk7DccHVBc76K1ExjgpHGjiUszncmlPEFxh8cWLJk3dYgfPr4X5
9DwKy+GwxT36YyG+on+4jOp/16Rlxu6HCLy+nHkfK4m0k1F5KjWvA/sI+nZYKzyH
KWHfNvsW+4RGCENfFy9YlJ1qzH2l+wWIdYWkaT1kAeoEAo/qphXbLWUoKhgRBeaD
S1nMxZJbluGYLfhXFbuitKLAYsgxx0rlNN8XaSILF1UkHzba/n/aSjCmYMmu3nnF
9778n7m0el/Bw6sl1nSo+H+lwc7a1c/3xW6E0TPkZoHvxaG7xm2OHopfoFnpvVBW
xZPd1HWXKVtzLmxm0BuiYntxlFjeRETJyndZ5OL7cfqhfqh6nsURGZHiC9Wu96YP
Zt36W+bNjqJrXUq24j8pWWzwI9G1KJN9JFGxcoaOx3md5A6XIRgHjqyRzytkU2R8
epM+1piKVmiyDsLgQK73iuVOAv3Z4TxRzoMR9BobNYw7Rqd0ljZHjhOZbCqp5MhH
4tw4FcNcHUGm6cqrvCP/Znx4EOHOBJrHWaLVyS6WKJHQN/45QuPrPIdPqChGYujy
CwhqNopXuVhFJQgA/mRNjvsdXvi4YS+kdBh3kBIbffMvhKy58DxWbt5Ogf/0aTLJ
0+f2yeUb1KwwJ37Rzp69J56fZ5PyUwAZK+2eStsENaPHdr3wFshkbPsurJUUtiWS
5Ujw1ZoShDKME3rreRhB5JCVk5NnDf34ZUriv3lG6DKgIBmYNSiZYLWHkv2pV8+E
X/MAUjutxIpYfGy2fuDElGloY914mmeEjOM2VmvsKwLanlwHbkoIa3gFEbbLsX1D
eidmb2zGW+Ct2wXK6z39sOyryQxQX3uyCn3QK6lMLgxJMlvAH3s1slIU2PA78jT5
qbX5STUMrSOhJ66D9EUSH7ZQaXG52Sp8loPrvbFyftyPTmqmkS06C5x4IZRrmtnL
3gYc/Waw1XsXVuZLdOr1mgofA1GyRHFK29CoQYiwqVF4bfvZ+COOGm7tAKhHSCoe
XRavsXZ5RX7jXHA7+8727TED+dyUqEWnFGVW6E1OvxWtINgwu+PI8NcDO4q1DA4r
fgbnwEqQ4ODcj2gg3Xew/ZPjZR5u1CtP9s5akFErrdoa6KIjL3TsrKUDNN95vkgF
RmrzJcsYIucAQqiaO+AJT266ZOwRgNm2l786EMrzqny8XY/QMJX6GAb5XyvQcvlf
7WLUp5CNBu13jgYfkh5qtm8qdwfgdENxRw+s9zeZcgH3/cTkDJ065fKrNh03uEvH
Pne6bSmPHGohsIF6oJNt+hGXTUdKib/MnTbOkGHvsox8wE71p8AZiXodjMy59I4Q
HCT9CGiq25MMFT5OLpSBHZsXS8vVKjslC255SOOXQJtHuY95MI319ah+IZTpm0Nu
oe3Q8Iwaowg9hzmQQGk2ofzS4FCCRRVak9t/0Mf/GkCjT+oqyiRuXXwv2R4e2pgF
1ewxBPzKqko2hbf9Gq0KHjrOo9omq4sS/P3leOXXOxafLhiV7yhYsETxlvOL+Toe
+0GCIjDX3DeGTLUilr9b7keLKLUN2dWpq0OnsOo7hBxwFRSrEUqK0G0YQzreNJ5g
lRxrJRFDT+tqhnlneN5moBQZ92nfWhbu9C+Da7Dk/d7uBYytFJ1lvH4M35HJM11o
W93zRTX+Utac51T7myb8Pool6V7tifD98h4A3HeHQg5nXSl36sZW65D/X4Zn3Tr9
frdWrz5o4By6tYkTt0FbcERHhfzWykhUfPWy1j3aDPeBQ9SVrIv2XjwT3K+NeNXG
BId5gBVO/Q8CXNl5wr31pvULlLKptftvXrwizJwssL+LMtsZU1MifRogm9eClhyP
AAjgYTGjtH86E6Zz429QjdxOZ1637CLMPibndZhRgCSOcJgBhj7rEtT16QuKKN89
zHyRLmG2K+oeuzm349n2MpyMUtsApBG1Jo+LKBhC7b2cX70WsL1pDRaS4yUxjTDH
deZLd2sKWz8xR8oZ57EzhsHDKAajlqYGOXrRyueOh8X/bMUzJxQBPTMx4LQJqlzZ
sqthPUvEn9+f/3l/bGzPyfQZ5+hICmTl4B9pKaOwdeQsSSPvnuKXpohjyEsj2GP8
4PhugLpmWaOesP9rZnKNhf+OW84jEl1FN/jjVL5QvBVDR9p/FPEsqLZ+VX0Fv8Ct
3VmxubW1Ovhgo+Ms4tYwrqjEmgLELXgp0LSMaZ7sDVOHicjLVe59I/lm3Rpt1jFn
5gjlItMqjEz9dlgNdktawHsls0woZ2cfFtd2GJ3cKtefZCPXGEqremzemFUrTEsG
5Ed4KjXjAGDD6w3NrjOSWvE2azDkggjlUGjW3OInQewrFLctRBkzmU3Tawp8KHbS
gHsAU2onCR0ozJ7RIGrUmKltWA9pTlXg2/uM2eSpY/Dy2jWlIS3O+Fl77z2pzu1X
GmMf2+YgD1k7EBreorQXXkK2W4SwUC/icQtKTYLvmhi5agwG+p9UfzkYzaAbGNTz
XAFsS5xMG6avPQsBj0jhm8Ht4Q7uTDvpDXR+5VPaYSAJSFLjWWo0tfgFa3BmIwRY
spE0nhgyz57Jxbb8/aISmUFfc+3E03j3MOI6bm7dIcilxZY1e6OmdGtK+N+QLIq3
B3cQBq5tdXEX7a7/4U6jLOxzu3pP3wb1bFdaH+bhrCkLsF6+Ae5L0PA05RtdCfM9
1GoBGnjXhVAajXtbCX02KN9sE6/33v993SXPY9LMbFCoI9mDWkn3d5+G7Lj7T6VE
XqQRhlPkug7F1Pj3BNWjHYszex4vsvv0E6LzHYURPfjc8xaUHcPJZIO/R4Y/7+WL
h9FlwnZeHcmaxi1IDxXGeTHcCo0ypYDLeOHPqD+Uw6tE4lbifHh0qv6Io7GwMP3A
pW/54/DTHwu3a3yEl8pFgocdtRHhBVM/PyQIcV1jUAVy64T4MG8+bJ18+FSiph5p
cLgJDlbUWbKhDW1Pntse1BEPm0yg5MjjZi567mew7o6sI02pDhysRTsvaGLZ1yMS
oDYx6S9ryYT6aLMz4wYnDNbE04P9XTI1i/A+yOebkdfsNUjtM1LYZG312/DiGBMf
LsXVzRI5akMetHeV/0xOZne59B5f43A2wbD3MhB6dDKTTB1iORjZkxWauXBSjnhu
6KR+Vt3lmCKxVKInRIKDNyWGtPedB3eYayNgRrhfJGoIuGLDxGWOpgKjne0M5Zo5
j/w12LGKpWGyaPHTLENT+GVlG2KwpiIyMlNb8iILPOkz0jlb+moksU3Xf7ZcsWuA
8rzzsn4EMt/99ItR89iOaUdLGoTR0465mLQfg5jiPLKozF2glglABJXEoPFTcFGp
i8Zk3/TPHmaLkQD7GmfdcQwPZJIOWhjD86ojHV3+BMSDDLE5MJqIcyBskdUs6SKt
Oy48Y/VgcNEOfc+tCXehpoUdBYNYxmcX2rR3Y2TSwWSRIfHvEfGPPNuuZSFKzaVi
mD1ar5a10H64G86e0zEIN0+L+eQtLsODD1wgBpZ24gEV5lTqkHaexz3Km26jZFfX
7dS+z5jOjmksB88uTFxny21P1zHW7/JsPIylEhTxE/bc6ejZ0zYxjTVhY7EbF4j/
oQ9777qM2p84tWcH+3BebPkKdOkoHe5SzzCpeLiPqhxg0PZbHB8pYAEfHqQGPL0g
nQOZh4HwlWHxLDo2zamwQsg8P5SMRnmBahkxy8lt5k/iAATZrYWOMyxi31pcyvN6
bGKjAHAyXhnLaNogpBtkS2lh3Q12mkwAhlaVt/BwmmW0AQLoFupWsxf2FwDRrfKS
bQpPETc+YCsl74kyz03dS8HFfJkx7WBANRxjcUZyIMHvqC6bQkg7K25/9AnP3D2I
5oO+NdV6nLw1o8D08ZWnjQ7YAEt1fVWERnOOmUrTsuWez6JCEsPnsvTlVswkcYiz
bjq6OARIc7WcZ32OOX89L3GBmpP5PwXzJnzk5qsJLAtuWNe98DA2NOcbVjb137E3
6aeTmlWV5Kjo67Tfhzq0JfxMR2AX0wwIM89XYE9H+3yDIqbA8h6HmmfKJ9sCK1oO
YvXI4QTZxwGLNzC83nuJwRSpmXVeTPH0mPoReRQi2CM3TtVlLfnOJHrVxV4OoQLQ
rEt2PhGAt9OqYoWElF3xr4ZvRXCvPAqrNlQ8qYnN069EbRMDH9y0zWwThC5f/1OT
W7a88JCb3XZERf4BXt+0DIMGs/xRlgIPQsgakfkzdsAG/v+Vv4NoQtbitRE0MKfQ
0L8oFh2OMZKAQwQLNthpL/6ZOBJZUPSboLkkEeDYKmpVkjvc67kf9Ejp1y5XQmGr
7pwlJt0slbJVoRoFP1Np2M+Vc59kD8YZH+Z6hVJ8G23+c5z+4Rr8wn3jwE/S+cG2
lzZUZWDAQpKWkn6DA06se35r/Tl+2NfQ7H+eDrdzBKXBq1TMDvvnj43cSNY6QbbG
FjgcI4lIZ4exWdKr90OV1eW8hF2AEgODXhsJ1Vc4mNwoAPOklBEbAl6Ng3CVxpjP
iPUkHiubdIfP00PZVxwONo6ZL9tehnKp/kh0/IQkfky3OXI6qhD4VUsdaa56BA5z
zuOX4JxiroWFOo3ic75u9Pgj9WxT0tffeynNLe1870tpXjT7rudxbhrKH6MrLUGF
8TrqckGSW0KpCCvHSSijudEN4MXs8H5wZR0qTmdRrRdXP9HKMx7ScalpQNaTTh5P
sIbvXST/xHkBjEAOY1EERJ8FxNZC/1Y3fOAHW9f37aCWI2m0HONFBVMutgF2yWHt
X5nHfqebiKIA2nO7Nol4LulPkSFS9M3J5V1dM38MlkWcIZf2iHienotiezYJT6LW
IVo6EpjABWm2Z85/xN1EqqRahKLxsvT08uR5TrFR2L/hJT7gt6M6bavSCpoTEKWc
6TWdYzWF+HdCduaa251a+1hbsEW1EXwUgSRjYkJXar/PEBxfVerH2SbA0fBt4sa+
/Pd6SSwFxZhJ78HS4RBNn1lHTft+ia8J7rBz5fFn0aOCoYuoCrlyMcjYzlL7V1cB
NZxWcrZGHfEm3Q+WWL/a6KJYWx+b4AB8g2ZAOgifH4jv1fhO343s8FyR9eTooY7t
bZVLR0miDxw126z2kihZUj8hyw576U8woLWnW7usW3/dzaZKiyhN9fLdONq0gx1R
wda1DNH/e9gn1lvehUxoe7JT+8R2UB0cIGJiuAaYgEIXdhm2whqkuGBejAjbESPe
m2WDLZvRDVvh3jmd99kSRpgTyaHzYqqCoCkRBediLcnL9pTgabM15xTiq2SF9ITR
LoBsP6dMxaEG8bcuDhG4kzw98cbAp2BpLk7xWg7Md+XXq2asIBfpMHgk0Ablwqvj
pcYVQfKME9shx/QvvZs/cTRaNkBjzvxa76h3OkLsT/s0kjoQAY2VJjlogendBjDr
u4mahco9TJZvy8yV7AQGWcMGBnbOgMxjLnRmO5+dUHdovZbav9QNj+pbAvMcCnyp
0zDTXw+Ie4KYIczWc/GUWzNefSk3siqv8Mhkq6I/gZPmXFuDzXiiU5mBnmo6QcDN
y53hTAbVJHuY8s+3W9B+xmedjDgpGG2iSe5EP28F5Yta1YP4jNhg4pxDlCKLUBbc
+7pEUxjLXsLcuXUmYkLRIhSZYJ9Gz9+FH+g82Pfwj4duwKpAEugSfR19vO8uar3i
0pI7a84TQzT8xPm+QO71T/xGH9mDkK698mCseFkOD2hLbZ8H2Pl25DS+zX3Mx4U9
FX/Op04f33aS+eV2TfaY2PR9psJpPbqFAzHx5Mn2TpZ7U50tZgIHFGTw5kPJxFnT
U/G4jiiCIyUb8wV7i+6iqmw4aPSO+9etER5yJuYX3vZ7jNy0reMT04pq+DDzK6Hr
estkR6agT5Ig/4YzRcN9+RoWVufqdb0l3b0KyevDaIqg1f2QBdDNAvIXol4vZY/J
2AUe53LtATr0+WKp7gA5dQiVnzI96gVNZ25Kz4gMoXJUEx8whEvqf303C0q87/MR
d02exWJEq8aFbW5IuujKPjt4nbtIGNHCo3pBfCpNFtjYwTDJ//jkkKJaSVbqeyNB
Rg+gN7kTRJkOi8NotDFUmMLIMWmL/k0QYP2bL2AuFQd7KrLg0i/z8rjo8wuRmAid
dzssPdMzRBxILl19wMzkKAf3VxJSXIKwrWYw1mEoMN1Kth1YMqM7f9ZWP1UaBNdp
mLhZ9atpv4ThbOBXZ0qx/GHP/EnN6lGr7TKSddtP7jp1Lymwmnlbfu4hnHqxCNSA
umtEFM7k0hV6SVS0IXN3hpArsFDusAZ4LVhYJGMfspCQPkzIE+WibIhrdjhZQmEg
263XQk9w4MeZ9ZpiURZTKhz/nmTGB7xPJsgIKCT12zVicaOPttvf6tK9WLTCoq9w
r8EtydfzDDEgPZ9dKSRSo3naEtkNcxLc6xGeSjtHhgETfNGH3aHWBEmzbneNTLSA
QSiNfICILX/yziymKDxQsWrWeIV+JCELtua+u66FAkmAEINAEl8pOY+ITA/eWcUy
ir3LXoLQpI8MIKrsWgELunsTuPTmnxpOo5w75fkW7u5aZE5+TsX09k9V88pZDjFE
hse/OJg9qUXSDyesLyu4KKMiVlg1T4ll+08Xrg7WIWyhikZnGhGCNBF1WgiSH4uj
mOrbudsN81iXs9ZOKN3elbLo45OYp/z3mPWjfhlXUwCaNo8Sao4O0d3WXvDhvw56
vpA/dJUPRTz1bvJFuwwWfKQnmItmWUFSbg3NOrTbDlcE7R74AAAsa5fDvAcGJ1PW
MFP0K1QKoy4tuHmg1KIYKaAqa46lNjSK38m1t/2d8ExK4G2Nh0oGn+RQsTx2bSNu
kiP5a4MqYlJS+Uu1bXTX6+scyomlLuE0YvqU6P3lYd4kfkxssvCCSLYrLPQNc4AN
f7uic5ru1pJyNCuGpR/ELUysrkRv3cDrpAPEuDspAtwwKpJIgbdaqwjHCwU9AfnG
L1cUtgQ36JlWm3BtmpdjG5qk8QGpvSNqKIuP4bvYCOY7mLL6JIY9p+/9sZDkXHQM
VVi8tC9OUGUFUgmnmYP6kjI7loshwJTW7FRzC30F4zWe2iAu2OhrMECgjMHcG6sV
3UMeP5Ux/RFyJurdlE4cSr2Pk9RjyaqCmN8oY2qdNjVXC3NL1CmZVm2FCOl2fWCC
qAU8Y5JQNmaZYwCWG6K2HEcW9MD90nGYmPVhV49MaYAe0c24UUL8/5lFLQkIqKmQ
zJ3nIb39Wc2hlQoqk0NdV0+MH6AkdUQMHjhdHByNNKLl6L9WqtqGI7zyQPV95G8o
y3jwCe7tHasz9krBLgmCcXBMJ2h2TvcfqbPtQc7C3BY8kG7KclUWHwcT2Q4PV8IW
CqOpyLorf+/3F8Q00rrsqomwmcwPeGLXSYLy+xyMTmozrpd6mVbqEx4NNe5X2Zb0
60YBuwhBNIXYhUKMC24McVIEnjUKDtas26lrTguBKh3NL1+mckNE1UnP89Z3BA1C
v7KgywHI2M5bkoWHBYWseasrk4QOcjPaZL3ZVk9BP0R+JBDqhduPpr/CUA5L7Xo5
6O2OUmP+Bp98GXNhY1+8XdZZEC6mPuei/zOws2wxaToofv3KLQttoF7WdGXdNnL7
IQv53Ysi1lcZtED2dlkP1VgkPusGeEkCmLktg0vkYpAInOArrP7fG+8WGoBmiEPy
v50OOwr5kE5KJZC4xWPXq7jIbt2bfv8yLAFeQyYKjRCdo0nDSY1lKd/o2gU7w4DP
bHlCfZmhS/ZDK08nQz8H5DhUyfFKtrnVyCUEF3M0MHyT12q/atETACntcM9vRPUw
W3eLZBpeI627Cd+TR9Y+RpFr50tXnL0BWLpv7G5DZ8X59KLNzAeN8J0rlx5vxpj/
IPFgb6GH9bh1waIBQf1mluRT3G8ZJnhpsYH+2o6WJgGR95ZGvcet1VKw4PDfj0MH
NI7d0rVOieiH8XDQkBCD2UXzxDq/iVIqzQx/WLiOf9wX0dkSf14q+ENZEC0z0J61
oQGKpC2+n3NwudHybxadAM2bqB/8V1XULeLN8mQ6FHXES9EG61w08trKXe3Y+fFw
A8w3ROz/oRWsHYZTIXLI34ltlhMe/CcDbKR0Vc4fGDEB3y+dSrFpOLfpyq5uLj/c
aVW9//QZJe7wBJpUw04FAnqyc2UdQr+Nja1QMMPygGl0SXpnyxoxQldAXIUk3T14
r9gsFP+4O3pvuiJH5RqW6Gbf1FiiiQQZo6I4mUmvcmiyuTJe5666DkhUN4w4KmTq
MSF9ANVFcuL9WcMmQIH/r2J1hCFAwuZ774eeyGKMdPIN8j0fmDlJw4GhKmrXJbjT
heU2rgyyvC/mks3kci4mfyp4ttMRfjdz3Vv8hyRZf26YAlpcDTNOwaIcpGJFIcWl
2tUZq3X5GKJrc111aIfKuf4sP4Pj7NibmmgI85MwdvoXsjpJQkyAEejovqR2EMlH
0xMrGRzBlWsKm7AZ4/wCJtoZeN7EA6uJFLGkjth9abroZ2bL6KwKNKdb/GZOkV9k
mP1KLjh3M8fMGr7rBMuqkmMqGFGjeII01Gi6JQQtT1jY8B1fskZDqTVTrroqB0nP
LFGF7fOLxFdXDQm7wIWsUvZsXqRwj+hA2lNDAR4PFpPsKqDs2DD3OVEP7M62OKLl
BH6cjbXWgAIWC/XKOjvoWXpCN98wwJPR1WShOdX8jrGeiNHK4UG2KvUm36D3Ktp7
yk9/4rtaTm1qku2Onc5xdUdfHxvJLC6P4T0b6XSzieqaOHrhtPPzh/cav5tVCzAY
klpUQpodKvRkZ98X3dwTE9n59barORqiiu5CeC1B6ISFqwpdl8OIoX7MxxLrASAY
DXS1ocneU0SJ60ynpB8VXTTcVOKhFh8TPKOEsNETU8/tRAbvl8w0GFFfaoQs1KGh
U6aaWtZKjQuWJMryp4bcTUhCPBjf2NkBg5EcOYekx2EIcQnAEjwnvH12R5YbQDPi
TbUPvA8jzHVKiZcqoSf8JStW6H9yVr8kVNsQKPlqLooKnAuUadUaliMptKUERx5I
O9WWaLCvGJjR5al4GusonWoIFJgvT6kLp9c/f5Js0dD3CUs7nnzdKlgn1Tx6DSCK
74Ik2G7Hhzo+Kj1PzYZqhC9sC+ogONcPpotDJDjmlK88cKDFS8ZIka7tNn0wYol1
93U/QeqK+k57QZ+h625V1ikbWHXhrrxb5/qeC1weGiqNzBK+7X5OT811MPRmeuSp
K0nrpXfILtZmmbDZ7cDVc9ZBqmQAIqp4xmyCD4qM+bLwJBndlVS/LhqKbUzHYkDm
JOb8htlIGp2jjIa55dtjP1f8+3TdDH0tIQXMNSp0x9SCWu0EacC4WOJvAoJiKrRt
QLjsePaI5ysvDvnWtazdha3XUaqiS3xE4azspMYTWT4p+RRNSJoXKvEtGHGAsR0H
l2iNGUE1UKciekiMKHCPD/oWDULruIFbIFIV62JAZuRUA+OiYhs8/hcQ0dx/KIQN
89KYs9K3oFb2gYicrzT5TqDiT1NE8NxjB1mxLY9rJHWYEu//MIAWjvgeYCOBkroB
iuI1m0KUfYQF2uuPrJDcsgU66Pb+FtWYUTXbb0VnM/MhhDcZUONe3tGlQHlyoYWW
o9jN83lirJXaP0hU+kEEyZshLVuSTWHcIwIrF/I/R/PX1j2IH6iA4zksctRuYAzw
9tYLigBUDVDebObNeQStaFrperbtzlnHKDR44qYBx6OqciBgE+Yvgm+SkY7ZcD4N
sAOTNiJXj57+bmXxAcDQX70O7eYkkisbf6SDjlUmhSILHpmJ0Jeyu3KI4mUg09nq
mWh7/XxDToxuNurShgNm8Z8+biTQlC7vO7XBMVaG0CSl4ENMH2o3k6HEro57Dy8J
351gQ6kKfTBIdwZ5tWcqSDGeIIWNtzLBuBVUbYICUMLBkzoA3KeQzlFGmvGTmK3m
O1RInTnlxHnhz855erVH009OdKw9/VcFT4JvkFVWxCk8ZjaLdLPCxDcYGcHMVgQv
sMrdUq/jSFIjVLvt7KdcV4fu/3931+CN5HO/IZo/nII9F7B6c4smLteLmQd9fCMT
abBBiXb+yi0DKtLRzZoZewREJF6cexmVD+WlI5NzQkL36bsXhFzhLQA4BMu8+uU2
SYfWoFP84jG1pGcjr+IpgdprDJHTtDeUtel78/KaasYBnWyiLppyx5qz4Io07dED
VikpoGupx9EfySm6ps4Klccdrya1iJsSMM6FjQsHeh5A6hXhjk9cN7gBOeP3qtQx
itO0Palvcpzvc4fWqF/SiVXh9H7Nmz45Jnhq3sK6x+eFaN10793V+vhYKF7Gx/4j
wRmPTRPvDiedl2WS+Xp3pY0WnGgoqaHQAeI4p2sigQEIylDQb0bl4Dm+f1TieXYz
LsQcUWpZSibX1m5R+drEzUzicMlQ9u5Q3keMoi0R/NcN2pPjjhj5bvisnIan1CWj
cXxZ3ixhituF3gtkfDPjxmyeobDnu+ZAxjVfp+zF/S3+PH11nOfMWhrIxHhtKUll
C8Nk7n1tFCJJpvt5a7D6BSaeW6/9jmgF9esblAKWoViisT3V8rmtlguDMsPf5Xfb
BlUFKa9jS8NUn3d20qRxv+if+fsYCaCT6/JfOFDdzjWtM7U0ozCz/Y9Wl0P1a9T3
Bv97F6M2YfQqNlM56XE8g7RjOjNV8WUDUZzcrgi2RFn/49yX+HLQz2czWI4d4LQy
UOUS7cPEUXqPhhAT3ahKIg4csXQgl5Sz5dYBPxIcx+TYAM5fynjCSbHLWWB/a0zc
vtisF0xuEHxiPywyrANgWkMpfnyv0zEHqePgl7/an0F/O0MeM9kMIvxuSf4vLL2F
cSoKmmuS5RVqsawn4ui0+dYPa2tN7VD4G4BPsbrHzgLgKLCh9hlnAm9o6sobp7A/
B1f3O2nH/AbSt48xpHQLelBmVJqUdlZxznLYlyfKaxINP7imbGopy+QMiqAYa1dV
jD59wBfkhJ4FNaGvvPISrwEEdgXMrVh63ScsoB9U9UL0UCg70IITMgeg7SA0XgNc
lUOlkQNqHgMeSYdqdCeJIgFpeiY+iK0F78I1zshjGNnQb0+6M2n4jZaZUyduTl2u
WLYUB9SYGhGs+LHa2P0NQ3GBI2F05c+SXRNhwdLETGcRv+9MH/vIC3UkSgXsKpX5
Ikk8c4UsXZ+U6czpwslJp0m5Oe8xoW5cV1eY3LEROP1RKAc5BXpG9y2mAckk+lq9
9LrLjwHVTKXMRag8IM6EVnClSngtGSwdBUGCrwtrikclBa9Ld+wuR1riyEYcsutS
9jf1znt60UDV9YA6GYZx3TbxOGoSLKzVPkV178nwkxlIjbsky3pSTDJ/hrzJE5P7
7rrNBxfe1Klk/wXI6IysciCeNYiipPijDr7d5eHfvzwWHjdlLwyoziXByNL16hoS
292ZgUGVE8wWXv4NwIlh67Zvi/nIcrdrTEQ5MpttaGGC/NKAaUzfBVPm9PfCEua2
v6zJ5RQTM41nwbFlDaNTZWUzj4+smHg6Au6VLH4Phf8dcdId27rp+rHlCsoJ2iD/
AlzdCa7xyt7AQbHoh1pRG6I+tgPGJ5RfwSofuUSPjJnA/bYVJhbDZX1Sjiq37Cty
aSX5RaJpXBbl477HDnrAbXesbOGBRukjIv9BeeRQLTXbwdhMhD8gcolJDdkyTpG5
z+3e/SnO2Q5OG2AuQOJdllkLp2QBw8SSdB6joTA9TcMgFtrECww+wnMLEOGovtTD
fdjmZV6vi3C/Dt9qxu8K079LY5sHSAwJ1b8LosqHsR5p4mJK8zWzr8aAgNp68ruc
Z48Ju1QylYokK3Hye6tDHz2PmbF2KzuZhvoToWJZjZFze2XtOTrVsgupeJQfyqd1
OFVZL/5pjxTBDwU4MAG2TuFGl3+HElQV3kpLwtXrAgrIjtugpZXv9VIXb0InX1R9
BnUGoots/Nz0sdoUiZyAPk46VFa6G6AvNnKhJUTxjKHzKZDNFApH2TmO8LLeRee5
WUOqcESHawekEiVM4JbQE3gjaOQdiSpsPkZRsEfX/Em09xTq8IeiQLWocvYh8F8i
IORSNuKQ1LiTTxsfmCOOIaAgAbTjBQ+4lwBQAdUctf689qQrc4cKepp97x3W+utX
tbkU8G781ihTqDbL5Dfd2yoNJX0xqB0pObuY6pPyNvtTEcqYJiT3N2E2fVfY755t
RibV2Euffjc/YgFHaWajIJrnbheA2PzGFLMQjV8u0DLmRZ2BoIiH5K7m5/y0Eynt
+xkBe6mCYCnd32mwE9rUL5mYutZpmEUqkUI9TsYu0jdtvm4WAz3KLBOC6I8h7PoN
NLLXx0mMPVfrrmyoG/2AmFNUO3fZ7/m4eGWgo3o5pCoAAAf8Z08GXN0uhQIPyfXU
WuVLn4n+KIrXI1M96aBLud6iEmxwaBGU0FYgjeMjq0w1iwNSIXVmHHLZpEe906Mo
hs0KkQzxASvqXXMuWrbk6Nn7rDwd8trEl7qX6wES8GRLn9tTuoT1rj5cUA0pLBq4
8K+wY0mMlCxmTTKF+W0f8ty5lzJiwnkLVKmWuemFnrPJWr3m5L/fc8BRv5IgGvTH
kDsiZS4Y6IEoVsgM86tB5HVg8RRgl2Gw5b3NMwJrjZKhW27TeUl4FpY8uFCPkk7t
RN39tTJTgHgnEsxgx48YW3kqGH9JcDOlpEiiAW66BlHv+Qm3ahl2Ux5bPAXzDzXH
jd3u0hpRqY7W5Vum+ZGXl1AwTXOdjm8TAqBY58OQ57g4xa11c4pfWlhgZlAyHZU5
nGW7mu4YUYYBY+4ogK2MXUAT9Llkx1VGjm9WqMMEmnDxw6pZBv1kqbXLgLWnLiKR
f39OSTVJMwDfUh3EEZCXyKA+m8ATqGboZ585Ad9acImNrFInX/GoTNK7vSRFyftY
9RxGUdy6YGuaBV02RVGicBOtrHOgugTWiDab5LXFqHmFAoWjDWqru9P963piy8Fv
88wi5rEuJP338A3DeNENzwHl3pniYTD6MlSg8OEjY6v+8SFpxnTAI/MQVoKOCIS/
GL8ouM6yp40ilJlg5UCUJRrolkL5y067WPKFCQxNqEuzSSBlZF0hhSKrxbt/A/VD
6LrP09oMMox5NQD96AGVAYitOGKKBsAX5lONKkoUCFVKgFOiqQFTCWcFelMZqSZj
Ju4QyVTsK65002a4Q1kUOo1fqmcZHAywGHoABNJ3rEsFuOz0r1QRj8DFkWkhMwlK
a7C6vTYkzV/qxfyIy50JY2a6bZku1x4555ru9klRYk+wn1xA3LtUSjlY50KG7GmJ
Na7sF4b/MCLcbrVqNIGGdtSfDY8KrnUiRGLwYalG34BdKEVDWnrfFYzluPn+C3vU
sL+x0/m6qvkV1cmdig2WrBF2wK70oJaBH1n1YkUd3gZVleETelF9EneRlt8twumx
pg1upGLfeoS6ggKrxUO0G6DOC/p152tBzpFXSWQBy3jWsG5UEm+tO9v1sWsoernw
r8kDXymGFSSZdUtnCLF1umVj0NgRW4i5e/dYJxziZ9x3G1YV6ORt2eSF/rVsAt8x
1/Jxb5qY+aGbKpVhhj1gecdzo34N6t7r3BZVn+HcOBnuyXs42zLNuTc13B0NR+1a
KkCII1IxoOwH9BUe/zDzcU2qXghEUKIzJJq4W6UZRzVm3Qx3y9ngt9h/aUmt3glx
6lmKu1SM1cSXjbGrQr/MtPr2kQdGm8uYLG2R7wLF0HnjUzyPf3q64YAojFj8QjcV
L/M0xuQfMAVHK3n5eJLkIksf4JyaS47c03wqc/3nwwYdl8bJDi9R4YLtRN+8IhKw
K4F75QE2NAea6xGORVFygi8nsS7Vsoyt9AibyPfVa3PNfPA69dTp0a44F+1OMGx/
I8Z/hqONkNE+IgMe+HqaA4nrlKhhNry+3hbHA7cNwgXdGG6TLREs6iPGpz+tuu5/
1sjFSwupz7Cbus5i1bUOiSGIDCjLcrAarJEGcS9GxVmxXlBlg7k7DQVAIMQw3O1t
+WpQKupChJRZb0qDEN1vQEm/YsSxs5uu9qV0k8ionMXVZrWnN2EJZWr98GOOkhM8
p8H0gHLh/IVsAfsvXr0+1X8Cyvce0TESBxEnLLV//7SE6SMXyDsb5o0C4hots9Yj
e1oyhnw3M7N1RNoOXd0CMuzfz2S8J7fxrTEAymVLExfx6FecL99RS7ayF5GSLviX
p6y6nV5EJn785vkNO5JN3ImLKVy/FR5Ba+GO/L4cEcpdsIU/N+s/URVWz3WRZG/f
pf8bUVwuUMyaiKVszvwG3UZ9eMxAoIdwctsg7c7gQtl46ayMJ+ukuEvT9T7QM/DW
7/eiy0yPSYOnbeabssE4r0XP2cx5RZjhxZMcdWgN1Mpm03ZQBYg47drzkgj9+Znw
LowU7N8fKiEMTOPUqi3M0+BP3rXHWYuHrwmPb6IJxfX8NFoB/FFcxQY9BnirCu9I
SjfpMCxXuOUwkKYJImt/HoCQmbB0+gGfqCkbLtcoPK2ltLSu8dsWS08qwponMsQO
yDomRLpIw0gB8q6EW2ne8jghjUkjWM/ly5YoJA5dTj8zhzPy9eVZ8+btLBbanTVz
0PdXSH0wqM0I8PTDGvlhN8pb4ByjurQ16TrPX5dbz0UWXqPYefUOdrRiKyczUo+E
IEwE2/AAASM+RGSP4RM/QKkFAYbHLRnCFC/f9Yp2MynIPU1Tj/DYc0ZPBLGPmeYs
4dCY+EfUT1S9UHI2zkYYbohqQ9FQJs55yyMy12i9dE+YjQY5XCujotEEGxAZSj1z
VMlLnDEHU3W3bRgHjdH8zLTkpfdfsUmyh3lZenbmSUvcs9mCH/N+YTJUfsLZ6JtE
BQ06huXsvYI7v4cW7nFKQKr038yOqBz5FldoB3wE8s38pPMFOMY7taPQXyfBDGWN
fGvgYRMXqvMOs1h1GprFfYqCtftEtwu9fgkzNbYc1nGqBtZf2AhgOjL1FdHLJhHh
9CX/l/mLvYIsCbgiE2cbBMrSPbIeHOUdHLEYLVgRgazLnz5PdlJM6BAM2QYvds2L
FDLUTty6BIW0YAQxd81Aa/jr8IsC9LsgqFSIu9pJweDVi+pTbWWkXjR53d//AFlm
I+tP63NDpzptkQ9uEyZ43UF9SuEQBDCMBpr4hdovU9a5uoDXo5uKXP30jtRHBVsT
3YOoT09JywAHv0AHPzDNwZaQZR670AvSI/Jog4ms8g4FqaoBRTg5CZK7NgDnExVI
m4NDfARaCs9RRwKC3d4hhJLhR6chZRbGvIw4TEg6dqIdMBwQWtvpssXWVEeyIiuq
+JvKTrEEIoquRCXinAkWr+jm5hVlZ8ji+INoikC0ISNC4Q2jGB9V68K9af8VI5YV
p2tvXXn0HuttmEMQ/DE2Iyhge5n6ogUJlkuRKFBEMeI/uO6xoSvBcowlBdit7djn
lZH9B2O4h/DBhqKX4djostVAhEcDBRTvw3M3SWSBIyFIHX38dW9paVcP2RRZXmhs
6IKj2Hgk5u5wjJvqLnr9wJUk/0YWva8yIkLTWTG0aQ7V0t8Fc01eABBdXnYSFHpM
zDIJlrytCn4OKmIV1S9RRJeXYftSgzsHThd8Ry1TcsPw1/JQDjY9WI7OcbSHyIdr
gUiZqfUgQtNT0rFnW0GEaUe0lCFc9QWE0vD2kkMgGnqnA91Y5g7HZT+uOyF+l3L/
nnnSJfFoDY0UH9ZoP8uxb3HA/WpHuxHjODrGtI7ZYagftf282pJetoWP2pHhEW/q
4LEVdVWchXYcQPc9trqTo9Fw0BRZSL7dQbX0d+pkQxldP8mnM9cbPpXr9CvwZuhK
5nKdqON0/Kn/m0v1AUrJAn5hlHa2+KuVHk0EVb9pzuGZtmPfkjU1GEu9c2RvsNG2
frsclxaDq0yY6gRhTx/88t32zFJ2EJAUXEiIRuq+yN4QLJbnZqY1f9PJPWCNz8v7
5c2mIjQSXuZ+uai+nQX6hB6FW/ZusfuB8OWLvuo5Ga1K2rAUn4NqI2wGNGXDUd60
O6WGJeBhDvQ5a+RqDWP/V2FcNchyDzFwtOWdl4T5Sn2kNozgbjDh3eC3jkMrnbrv
3wt9jjNMXVFRMMCl9H5k3Zzwl07Y4vKYiubpoPXctuj7H+tCyKrRVr+hNqHrk4x8
b9W19OcL/BLo/xODOrCrlIzPqeXSVkIlBXf7duH4OmLx/awjOFuaamTyDMbZHc3H
nn8qCUhnKfEWZw3QeaTW3fv/JxrMQdS4T4NS3ePZM2nqu7P4796TVteZhxGcNXyx
s7VA+MpDDvyulhzud2Sqv8XRv9avPlFvUFNJS7/pE6b50qOYjkBmS9YQV1rlqgzT
PdnnSiV+kcxyMuYTsmlqE7yQX1b2QdOsECS6EoWrmJtbmiIsMEjCbnP9FKfdp8t4
9MXv+uDvqYP3iwa6dJAJcD0zOsFGlv1lduzQJz7R44InmfhWjc5ob6LBxZ64I/mp
gZqHPiVNjNtqWI8sQ9l1xRR5Sq+koeCPbjYieWzV/6iIoM6D7C9kVYiEoC3yqc+3
qj5L/+WWuhkZpXN6ODL9mW7Rujy39B2xe1f9MhCFN5AJTu+Sj/vyCzotuuLmOe5v
ve7E4J7fWaf+C+yUPXZ2ergs21F8jacvBEsjdUT4TKKFv+te5RHEdmJfXY+Zqmnh
ls54sa8/NJXYsNNWCieM1iSRwFH5+92sJqAwyGU6sH70wXS+vALIwiUWbYu3SwFt
IaRwkikiCk0fV+32HL/+4g3Fjyw1Og7vrHvs3gcI3Vt5DPryvsIQmektks/5bSez
/iwS/JJYUqy0RnE24csjPt5UtdNFIfhl2z8AA8grekS8iyThMdjh4YqMroxpjNU6
gs2Zi8Wid8b7Wc9THS0fTX97WjDAtzycbdtu7LAaUCGt5tIZK5o47insu0eWqtfz
jLDqit9u1HMHPv6+NcyrWzq/HNMVvmCO9Gr0ynjAjL/eTe9dfDg+339leonVeY6c
iZuyK52t8yMSsiOhNQeXXeybEXK0oD0pJ3OM899aF17B0IqWKCsWMmkI6OUd7VXI
/LCAMb+W+YkO1Q9RP4j1JsBolTRVLBf4UU8l11QiPhGH+QCCUoWIu6BlUlr24ZqZ
M5c8P1LrySo7ZisJtD2nOgpfdc+SIUGNeT2/Avca8yoroVyXc8LiX2BfoVtYv8v5
eNlsag0gYtDFVkcKNHPsQDNxZ+50kwJPyYz87zB/sTUjaTmVCPGAVrF4EOEx0TUt
7wfTtUfM8b9/kEFmj+za9RD2AW/gHyBvdvAz2ZyT3xQQJbBMAbkzJkoQ+3ksv7El
0SSIZGyiuN5dhqhHXbJud/wacsPDtaAXtXM2V3M3akAiVRgK2PvMFTMDZsX4b/j/
ciXk7y6G4M3krN0evuiqeMygyLBPwXiRnKdhBqhzwhBhmLa8jEkY/yIcuI5nTtH3
zYnKHj5e5ED+47Tk3XvxnTIJLCTB6IfRVkgwTEQy2hjgL0u/MojGLQ/8dh5lMw40
zVP3Dee5LzQ2pJv+cmn3GvEVanMgNQGpgORA9r/83sTg5dUmAQV5UEzbvRrvnA+9
M/U5ehdsnFN02+oSugoHD/1YsnnyeWChcBOgfjVCiWMuj0K+GQaby0RU/wfrqFI5
RbjMmpxxoISvPmv/V7cA4EbHOBvEfdXRRIZ1yNBLJ0+qidHJ/MDRA/cc460srSDr
by4SVoGaLvyqhoCLOGWHIFJAThUy7mx9o3PdwRI8sBi2kJg4HQHNcjJSkVmN/awd
x0uVX+0Ruzzbl8on4jcxupaLQlMPEn/+qPlVYTl0tlYYXi/99IAnMnzG3dc5B2fs
GSWmjI9axYivNKvoOawdE9aGQDVzEZdqxm7HLcrYu0NRPpHIDEMH/845dUlkj74d
QZnCepzAC6sENqAvNnAX8RLbCXQSDwpYgrTgrX/1Ab5jAclidyBbGzd1iSCzjE/Q
ipgsKJoE10dbyvm5UDL46w/YaqhyKAJ7ySzd/kFMqNSsKoNqMMHnqhKuuYBuDKn2
OkOJdb2BCDz3KrPHlwNon2bESSns+XI/TXeFKfK7TRA2epAoo/u2vQ4s/S1YrSdq
F9KGpDHwAST0KtXvKqFlhgPI+5oSGeZTW0iD04LPTxsIziPH3Zadlkry2xgnkeR3
umYJIq7o217KU51tea9RLKgPI8ZxG6iinL9OMz6FhdRJiNliJl7PmdOMUGrPfLMe
7rCHzI/0KdJDchm/F0npCjiP8Al7lhMphetpsMV9jh1unFgDF94fgXsezEER2Q3b
ITdhxEnCMXCLZi8kPVjHLy1g8xdTh5I8rKvelBUlL5lJt0GI5S8bJGxOVVh3+UDV
Oq/m8GacViHC/5Ike3j+1jGkFxuDrCaKNXC4R1Rsb66XEXUXRfWrj0Nd8YoJtqFh
tgkMW/YEsriljO+qQxrPbmtXctV3R0qL/FCLIE2b9tEzu9SzAlCgXcc/MAABzhhP
mMY4Z3h2bxX8zfgLap4FdkCeRENN+MF/FLJq/CNuevR1fOtrfaP0iVYAGTs9NWEB
2fBjL4zgJD8lVpX+hbmst9ArnYztI1dyxApbXnbVP8Nv/RuIGK1VGnIHX4TiTqbt
CU9VLj77JgY1sfpwRAC8hmyHK/6MH+AJZSgg0SBgdgDcfreyukqcyl7fx99oxnUD
URWCpk0WIKmTkYR5UMLdwEG3bbUgdXxVZGxZt0nxHkGem8CY5gw3MovIw/CiqREP
hZ0gXZsjUs7xZBsG7xCjDr+l5PMOE8sqZf+OL4OBDkF1Iha/6kkRL/YXh8ljC7Mx
DwW/aOE2Ki4fGAfiwhCJwzsid3Issm37RNl6DS+k5jypzN9de9HsM+ws3iT381PH
Jo9qrVP2kwk2cqtlq46NYN8B1p4a16ArN4LVd4f9Z2Duh7hYa7FY2ZeboXQQ3+j+
zz40tNrfTYvD5oxYVJB9TJY7m1w9sxTm7yHoktXLj5cfwDdGNuowU/ygnnAPmAq/
FlMjuQ7BLOzC3K7ELPAyqJBDh6wVhr7AQlgZL+wSDA37HaRZyXVKMhvYv0UAL3RQ
dXOVKTQzODgs170cJjISr8bvWVzk4kX4a32CmNhmw8ZxXZPHXAp8Skob7AvHarda
7mkn33kVm9phG5ZB4T+35HqCa8nhhQFvNl4lN+tJFemEzqGl9wXrSn9Ia+Nxa3yB
3Sf2sre1sr1WWyDsuSYboAEpDalo88SeLDiBkPnFaJlauHPRGn6CZpOl8WMUKpx7
+JopHSdX21f3bUsv6wsyHpcTLrVOSIvZ6UM6NQ2j+5vqaT7bakDqVbZkmOTv3qfc
wMCy/KDwMtyNKI7kraaNYzvT4LtY/HPHZht29+pPuRsmfkV13dpcOd9whjJIDAqK
8roDa0hvyEcV1EfgFT8R08WM592gEgixNrof24F9tGEuL1CRX6APIitcCeGhuH+f
fTKbcC/5cDw8Y59UoPHYd2ghDK6b4LO5Eh7YBSDY6yDwxSC7/knPXL9L93oPMNiz
EwWxXCYGZ6YUCa3F65HxooQ4nA3VkadMiMeCIdYmShLmB1+/rVWoW2UvBr518jA4
STr1027uwhmTP5GZ2DRNumUFv5C61/SkqY6ODnStU0qMCsNWuvw9UXrH939CQy/3
7GI5L2SXPFpIArwp1FdqVcfCMKSNW8hNhwYkl917/eN4sTa+m4dmAB0PCjOW0mdN
GgFqODqWcSUle6eJZOI2qohSehrCwEqbZ2SHO5jTm+kTztdsZluv9CXkmm/jb694
K0CZ3pUUTxmmq9IaWnfbpi/PLScj7NCZSXiwsZ2xcKAX76CgmXNjSYDFmqw8gRs3
ryXPiWqcDJToRPFFUfJ82uQqiGErB40w+ABJ47srMxsMNVBbIVNNM/qhDBlL0AeE
ZTRl80Q0J6LC+IrlErgXB+kpQh4g6pv19C/vm22cH7Q1cAF92FE0XMF/FYy7lS25
sbQQ9h/qlxInpP9VlrN8T9l5TY68pd7zLiCnTM3gqzArZReERkQcmxK3PIOM+WAw
0SKyq0yNWAZpo+zmeyBTmX/0u2JbibqH66w6uhtkcY/7Ehw9g6FD9Ypy07/hwG8k
htWP8WchoH9ecruvpdH8xVUctyjjWlNQIhnkaru9UzZeuB9gDxSjXBjWX10c4h6f
vjxYIkiUM1FC5MBFfaDLe6U0NdOK33XzsPX/d0btH8NmCcyKiglYQAJC0PA3nb/e
PhKLBspNnJW/R8caTu8nr9Lo3b2Fl2xbhMdl0NEJnEb7+Yox7iIv+LpEHvS7tkh6
qB2Ml4gk1nCb7lZoYFZfwzynkn6UCTgjMb9OOMEqRR6XwgU6xj34FTez80qtXZDc
0Vd/VVDZMSqOm1T5tNYxu1A1XmZ7xozLuO8ht4Q+oHwsoy+CfViEBfjeUs01WQAr
wsDS71G2XsTqPTuqElSJilq9ZuaSY+X0rIATNr3HXIkfT8VKGVqVTNZ5YfzPe5S7
RQEzR6y99IIfxlrdxs2CuTLCGzEC5cYuSm6GPmgp/j//iwsyNIYE4RPViWh2RwKb
ectWXsh3u3FkIYg8cJn2YijDuPsNokhDlDSPig4V1+c+wNkRnFzGyCCrQzZP5EI4
F6MDl57qKt6cdLYozKoeeQsy0T7Oa1zlbXa84qTOpSCi2MDRQYQt0aWP6AJJ3UNE
xw9TAgh5FO+0Xe3sw7wYRQdUYOfWi5fqxuw795GImICC5C5aRHcVxV0OlbX5BqE5
RQOogmaVyBU+cvcTyUz4zxDBBX7Xb527Cgv7tZVp4KFrixiT4sTLKayg87xVjBcT
DRa8KHr9UKK687HdyTM9zT8FxsQh3mTxpae6fCmxNNGWuYs7L4l/xWyaw0/+XpyT
o/qLylh22A0DKUwguouz/mYRZNeq3nWQK07TcKopPZXfNTAhBxDSIjGd3pIcG3ND
vn2DVwAzR0/rPDEhm3zREZ8aEiXkP4UovTGg6Nn6jAJDKkNGJCoFXmI3BkfsImpk
+I+sqnumvxmLvF/dpik1SFicQf0kO2l6BmUfpFtcIsu6ew0rN8Z9xlZoPqEntqDl
I5jMr9vl8QBEzhrBXv1ldYRmGrkzDS7exg6jZy8IqA1Zxm3MHQ58qZuKWCbDavLg
TYFyNlXBMhcxb+rIpotvLU+FxewGpImx8/66ccpipJUD7aALHqoq6/+GKwR+SAZt
fF3Q91XOLNS9crJHGCo7l3Z0EyG0gCyBgbCbT98s1Qz9Hy/wOMyMX8wacgmL87no
S8rJ8Z3zWubXdmOLD4xct9BelocYid8kFe5NpY2jY9uu40/MvkIRaCeJDqCAuErR
Q3N3Rxy+bGQfbTbdfiRft2uNLdbvQPQuQqfLziBLh7IL0IjBfZNs22JPoIteJfkO
Z3vdiNsj1WRSr0VJ2VCcM2eHOF+vSkI69FKGsmANZxbRDrrnH415fxkm4/2WM53s
+0Dc7WVGpPedQHN9Mo9xn2AiKJOM4XyfM1ucpLK7nDn3uqFcLbcCS5+Ufj+OFiJg
k6ckg2jKLypoIi1A08d/TVBJQbOnkQ/rBCAUbx87dqJOhc+nAyt0wP4SfqcZrGM4
Oa/GLA2f2A9e81dYo29osV6mymBNbP4DArTFEURo/g2amFdAiQubDID7OXJNM0K5
fDFhS62M4R4y0b8EWr/KmHLG3OEZI93IivUEHo5VXhIe0gwF4NMBD3/+khYosN5S
HIvP8G6bb26vW1qVT7Y43bjJB8CDxCPJ+sAWrS2ERmY7xfHEWs1EpkOxKplJ1zq0
6Ry+jAMPQZkw5X2NfxztXAEIF3OdXtVwYzZEHoAhZWikWrdPBT5MA1zeI5VKvMRu
L0+j9UJ7lgOySAV8yuuOPZScKe0Nm7Ko0S0dmPe2sHQliYTfOPxnCTqOgDBRQ1Z7
hfARCXcymchWDKgh/yZiPUz4RvQ+1YriL/qL4ci21FwA2JBDTG7lOYIPqOzdP2Na
qmGVJZKbLfmIGR9AvQzl2um85vERncS6lfYF6P2wzGBLbNHn2w8kQYCHlZEFfYbU
9fk8G6fkDFolg7AjDxuz2Zt1i+2m+qS1itLk8jbTrUFxqJ7W0Eu7pJPa6BhyVEho
8CHeN8x5sDxzECART7dVvf6YnTVfnEcO21phvrNSe4qgJM2mNzwFnfjIykDxdrp6
cSqxn5Xsk9UCeyjdKtyxvoMXBjzH41nerXJXWkrzDcX0DXBWNIPhdeivtvTvMl80
Kvzl56gqR5lrdlveMAHiWedp/vM36UBKca+mbuyKlfKtFtpOZijwiBCUez817/+W
ssMvj/HBlX03o5zmeitdEl55/bhaY4vduOpNlEsLGDF/ggxQy3LU5Dv9iWb7ahHO
EE6iKnJI8WordBtrC18IIu3bMbyYq16dyEhNBhn5/dvPkPpIz2w7ibRF77VbICfP
9k1q5s94A4kk9PyNkpYpJ6a10djF7jvxcl5Sk/Ul20ASUO37ZGqyAAuS1m3my6KL
SEGd92gsfrkW5JwalDLfEoOY6bfOgTimhUqePlZO4Y3pMxlSygu6lVH8G+mMY8U9
WhlMZHT3aZZnQy7wIhTGIj26/FLqNy/YOeh0J03jZYZispUwCGGfKuy1wsVC4eN1
UK9p6UrNXpA1Km/yohQ1742J2PeeezfGvFhxhdrSp/ioIQCNOvmRNJfMjzhA/0Va
V9/2dEcfisuAGjaJ8aO7/4xcZWVJUipoRmzfzq43xldGZXvO2UWTFmOyc1bP7HBO
LQgzSGO/p5T4Y3FnZ+lSa4+zpwQSpQaTkwn8vP2irU5iAqvW2Yhppx78UDJPJsuT
TFHfzZn1KqLtopyFuyZR5ekTwPhQOXLTtKud9L4tRe9yg4x7/U42jZa3E9moTkop
/JVMFG/ffszpVOAJ27gTltCbDnRVIMgvBRbk3VWa65QxHl25k7k/K36K/yPnFySN
nVXmBRgEmWdcH3o++7KHWzN1Bj88Q42NpRdSUfB/NkFdHrIy3BbGuJt0GfKu096r
mts8nni39GwHqln2aSX4eOXiPUtsazPmFXOUTb/3G+GeNQE5HJ1BWs8swfO/LkHl
POAY0sNA29e2ycgX3/goLhATbAwBTvUY++EsgESu431CyeuIWDEYZTiBAduU95UB
95q2SU6MovBZCzkTBdZhlRz+j+vdLxKkqX+jaYKI4q3NOeShrBN0+7n+XKzqnpeJ
iSdNgGTeNC+nXt+xguV9Mk6t4ASeUYJx7axl6Oh9pJ/L5My8KiEQzr7X8l/Ct/YA
zohKT2o2ma/AndfaSoJM3mQ9FZi03Ktca0+3KSHOreISxTJN8ZM9J4+/s+Jak+aj
cmdcFAqCY1BZI0JFqoZn9VddlE0ONdDeWBG7GaIrLYtSUqeJZCmnbVGWxDs6uNgS
Gfsj55cuFYxjuwGOZKGXtbX4f4AiZjrMBpIvQ0cGiJeuO/5Bug3rJpw1D5VvVatB
CzrEcmYVHfgwabpE8UBmIj9xpNhCC0lyHhakdPq5LFp3dm2FI9w7WBbZ3mKzpKxa
5HGX/NXgnU2eoXOUeYGxYb22p0HR6iW9iFScZ4kgP7UPOzzOSGGoy4bdh2Uz7icr
tMCxNdUkEl6vZB/r2SlyAHbmmOA9eATxMhjAlHMABSxreljHJxLlWvotSUcabBV5
wxfpuur3mi6LmDlfGEQ9Eug0cuZXCSyy/zpO6fWCk/6OuL+0dFPkBkp2J/Qs6hpr
WfetdTL7MIX+Ag/qQo9aLX683sSTeBD20Aj3SwrWnXyfeR4ziSSvFqr4W+wHmt3v
e3Gaw1KNHEa+pF+lWh4D8RaAOL4f9cWyL4Jc/Hi52QCTZkv9IcpwyLH9FY5POP9c
WFewGn5Du3HnBjt/BKA5k8tXxyFyzG+NaNkMB/BQqGAcfwMraM4HOzMrAjFz6Ww6
+/mz4qxI9j/5S4B9ZgQGnIVXcXFVkCVMi4KNeYjJqabhf5u2YQ0UXmGVvdl8Zc3q
v8ExiKbuakwnCnUZW8uo8KzQyP/9rnQHfMO0X0Qi3ihC0hSapCozxNV4Yq83Heqv
lUgDYQEZhiVQIc3+1a60cENdStm8mmJWkGqvoF0Hms/pUhMzC9aRRxJ8OrAQN3Zq
qI16W830UTiIuwH3W1JNwohLMRqdvZdXGLT0STeIsO9Uvqh0I7ekwvQYRD/p1qCA
9CAtwIjKqdzuGHRLCXMV/HOrANr246JQ6aOsKI3sG4QanD5JiLg89iQSIiT2t/yx
2j5QuK5G5PUv7IqZJPLwaFSS0sd7hm1NNr3fdQXryaUGIdawhzEjNSkgxKsM+PWp
YruKhES6MKn7n6qiEugJzgRRRAnRoMQig+qlgcj9qjZXtesnD+S/VbqkkXNgjKlU
pTUyD7HotcJXIspJcXEoRaOQCbt0j0PFEft4rxrVQxx6s2ppaStx3K7bvldmYQRE
yqsknWi8wl0DLx8oHtmJB9zjjiHPqpzbGW0a11IrrvmxO5UIH0p7Ut00p2um2i9n
qJnzXqsgFe/1yLa6hnbw/+m4R212KccVEHOyJFcRNGKNakHOMqlHkWbnx0YDmD+h
uhs2KZOZso1w7Y9o+leWKECUx2YefXvA4AzkpPgeZ7QE1+M3KLnM6NTGk7DTNHse
CFqYjopWqroa9YklAmML8rWRScuUttfF1w4IQx/inByOME2cfgSZjZF/si7XjITh
XrurAIQaWOWBO6wSHpHS7/+m64ahe/HqOItWo0nD2xwKnR1r2fJAaXE+ihuW4Fuh
FP97Cfc+MgzYFtNWtrTx72wnL037Zsv5zVelvuYD7OC/QlwvhXwAJ2jx6aIUQePS
L+SYLdqGrH2ONRZzcE9JtPjL1WxQ/t13QiaOEBJ1cYnO3P0kQwpcMt5kOJ72lMIx
TTahFVDzkeEy10aa0Exbd9MqtoVTaHoaDAjxyYoAriyas6HP116VNo9hOq6t3WFY
8VAhzi9ymN23yW3rRE8tCzeGWFaE+BpqriQ+YZEZlxWPPnLyaAzErS92s4gLvZ0s
IxaDSqSESk4eW7fVXDePqJET+VAVahwcSyziL6i/GXd4cXOUQ+vodtCT9N9j2+49
pK/nvUqPxhbg9bK1MDruexb+hjbBQDyJiWIHwDchxiIBWMX//DjwEZmPJZAJnr6D
kxr/hHiVRiJq653yndlYINZG04jYRhhL59jKvRH98cyMN9BKmKrQl8mSed/BWRwD
//3EHF4iEY10F8XCt0TGrHJQyZ/YSMrbaYC/91giVPzYZig29apYV2Dhmdv3JQxC
UYxG+PBs+GrMn3Vi3LjMKvClSVxDsJA03lzQbAWzWWt4oeGlvpcGpqKTXC/mzUdb
u26D5Ke7QOs7VdCwLLNy9qwfA2ok/zOBi2D034g4Dv3VrjhAyqAis9IAxLqdfB0m
4GLvWG4iD8cBZdCI5aYaSQnK0RN7X2N/WSLQh2tMgx6vt+TBNvmO4nmcGQ+fLFes
AZNFTBsz2MpI/TW8RUKS57L3pBhjemTAj3BS3U8pFBz056LEDB+Fa/S/h3TzVm3A
Ri+fhQex67Nd3ywWb7D04RWqQAYFNhzvU7mlUHEoKlw4un5RniVgJgP9G8bMCJzS
9Vl1bfqAw/pNEmFD92SPFr5lGNLfylW5WjMsTARJXvdkBJdWo3io/7x/Kf2lWfAb
1FsRguDkzN2EU2ohzOgChDbq8ODkyUJxV2tbmim5vp8L2MAdq9gEYriKRL5iDnUS
SvJzCGSrKCe39V29UX9tmAjgIgmsusdSp1lh7ErMts7O6rfEM8mLyhB9aqWjfbq1
oNDt8Um8ZUj1BuzgMWccuFJQelMqcKC+0K/2DlyqICO3To6Hry1IaFSU0WWKo3IC
pGUlt4cntZdWQ/WDa0xJymFmDsOSiDaz1WiV7cFl7RYFTd0YxjGqKTpWZHRBfGFX
SNoEmvM6PciVYEDYSG+LHBiukBgVXRWAarJtFXQiIjdYsSbD9z6rr/Ewyw7ksTV4
FKmoRcamLMKpRA4h/7HqaVDV7hyXR3S54vT6ZiTcF2Io9/5PlSNBFbp1erRmCD+1
oW539VinWKgeNM8uVapqcqdNMNvLRdDWLbslWCJQc0wiTqIPn4QgmVuVt8SNp75c
aeSuvfNTPezvwOY5waERjE/y4JQ7f8ZQ41k0IPg7u3Za7nsfVWeZajoHSBytKdHE
b0+JilnvH5jugoUWnuc+ZLcq3QpjAkfFkh/fBnwVg7nRrrl/KFB9ZMROTRgnXSGf
WPzTw3m49QHAICt99LYdx6FjaDn+Pi5aI/6dA9VG20YqnApVZD3RyDMpfTKS1fod
YyKFKhyrs/eQG08LwHd1/7GziGjxuZZzleehvA+eNbFRjTnEJqhpPxBqCK7friCs
2cGPLv45z7UKTE5EUC7MHDVXspQ28bBTXV2C0rDre3IWlEJt2nNP78MlcZFtfTg6
jMBwZz0HKdzDjMgT970AOWBySj9hSQtf8Z0RBkH8zWHs2vLjOw9bEnirV71HYLDU
nswdJ+jh58whjdqal9+9EbZjT1XyvJHZQVfQ8GOfPdpugXL20B8yoPvmKX3DloqQ
snyQqrb8xwtlLVT94ksaIiPfG18h18c+MCKhz4BbU04+s1PwE5VslKtEptRqSayF
BkkGHnzWcOPAl+axcZLr8s+DZSMrRBrr4O7W+GmlpaRSVJ7bLEyEtYBVTyfd/iCc
Tk9SOlBnZdp1rce0jJ9/HAdynWLaiuPTtT8HaAqtVSzs6HGGTdxx7l0xWF9r6GC7
5KJKOX4NRTFdCfRHGSuoAuzpkRmJFSh008Hr6l+DhbIgn8gQobqlnJKoKR4Bmi/B
QSFNqK3ZyPV2euFhmKRgVgz273n0HPBy///LxXrnbwUlJ7eGfbLnE+csQf37QBom
ZBZVj2+uSpTizWnxMpS9ZPFB1csEhnwNgNiCj713/LOefKhlp990UxyFsOpl5r+V
Ox9rleGGKyGRUSeu4bn5GBfbVG8wzQ8GYB/7QcgnWJRe0H/yM8HuRujkXtLKq9Lw
w4lzzCAIHLun6zGNtTXxga8mJqxNBYw9AGougrfblCwieDbI9QaaBhSzes0ekJ+B
qjHmxusJowZH+oaWAFrs7XQySwC2Zg7L/UB2NZJScfqk4ePbLv3bu22EQKcWsDss
r3XVvcYNmsZuEADIe0SYs+OaC1R9flxjyE54isAbEmXD+WvXroPg3Eby2UF5dM69
AJqRLAik2rXwkAPDnuc/LfFFpZlB87XgEA5WaGjBi53Jk6/HjO1fhqBw4vGlFj/9
LsptJMgLswQ43FJ/hPybfMlpTYB3QKolqYIapZde02D4n+nIk9jZZqcETN1YC0EK
aaWHvj+Jb8iCJakUF4gVMPCTSWeKvQ7RHG7PLYvOvYzK8wPcZ5iCciXp6eDE3pLv
L8I8wm+8czzwdATsMiWrWtUKayr+qCqzBp/3ML41bYBRrLF0NpzP7kLp3QEgZ8ZR
QG8T9mi/a+kEnM3eHjXyvDX28gHFjAl/EvJc6yolOesfG37ktDXMz7iGLUduZ4UO
q7zYuBJRGLSu/I9qeclADzSJ+pMUh3sJorIHmV07aEqclyFT8vpwZ5GjNvaMytth
gsy48uLc4A+6jIWLqX1Uosag7oVcRJEB66mRmz9e0+dYlravcOa26hbDCEo7H43X
zrZqtJZ17ArTdC8ewpea1ECa1sgUw6UZnENYt02KDNyaQpdIhkyWF3M5lTjQCDH9
9J+H4m1RRv1DTafuVXmS94J/V/74f9u8qLRkYYxYtpuzsW0jT27d52uZbZsC1Ujz
GgjWnhodxEtxdHDtaZBFBgIFp1Wqys4JgmjymRRT419nqhO0eDgfpNHPagLOnVSQ
YLeP7ShJwq2DGQoKNIZTJ+V5Nadx/Zass/VxkrrGX2HhcRGt1EdongCLxVeOFPEI
SjaYm9ja0rKLZi6kLMOzXkND8G/gNVQzWEaJxVN7YDpL4+KMFj/t8kximspONoOG
37v0c44VLcLtLnTMdG+H25Nqp5bevWw0LbG07I12opF35i4xCdS6mCfP/KU6p/Yh
c4iFwMfXOF1hYTq9lrgcIFwRSFhKMT227i+EYsYGEC1Nns37yhOqd3sRrl26CKBa
vEp0FgTwTlUUxjBj676flG5DTMHg7rhx9OoCS/KfDg/Le6hmywJUldpEW4NjjAeY
R7ROHJOyqFMPE1edTNRecKPbAS+s/hXAedrrsBF8gKUAAVicyi/TOOgy8B0XTo8D
UQdoZZroy4YvVP94INy7/Qm7xFtm04wETUCUcVyknDF/6ttNOLVyB3JVelo5JrvY
bOy3rR6diFRPJHu1GchudGp0meJB0T9rkwuoxPU1q5ReSwlCOhaVPON4zImSiIxD
3jm4+LyXmFlPE5dVqvbzZ3xpLa7un7YotjIlMYrgW5QresUM1Xn3jwo+lYJHSHsW
Y/ooSsVNSXUWOGduCyXKSODoBWIvf/eVhdjtFH+7AGNGfznXduKHZcSesQsezlwe
2N5HmBj0DTB2+kDmqteSEpagUXJE15/noGjwuWtD1Bd4ON76DtyuFXZ3Qx/RWFNP
Evi8RO/d5MddjFKZAjTxbpdbyawrQvgrrYf3wmaNr8eiZEBippYTxpT0ouKtF9RT
hIemeeiP0K6Djb+Kz//lv0eAoQTtW/phlDxP3go57oDUzBeNLThtX0Kp4rNdaqlm
J6eYrZ4J4tbzby8S2vytLRfgj8V4yPooGMTiCUTq1fVko7Uy2aaOghWK+Dks0qn7
Fhbdc/ns35imb+dDIkx9fKun9CLwdr1cez3GjFnrP7uUSOWkn6rcyGUVGzQWIU+h
Sq7If3eLkcvasOqI6C2ssfgzAwO2sTUf7kKpi1497ipgdXtwOgTsjnGUU24/8YXq
CfW6jot8MpeR7BQYAlCVIU2JnfElVdyWlxT8zL37qcO5NpyUygGRdJhShMuj+rXG
VbRsbBVn0tIk4sSRZiizrYSubj5pgozbp3Wf0xfNje50hjBCTfWsIU/vqqo0G5Sq
VK3f7VwbXH9d8AKWaIIbCt8oiEKc+isg4Ir0uhZONHr5u6dggtiAg6oIROy2U+Z6
VEZ9kv6SCnEqRSVcWyf6n/GHqLJQ0YZfYbt+Wndg+tMR+BNTusp0bxONy8sKDUEt
xyWoxtdmKiVpCNFeArSJn5RTYF7WTPoENbEdmEYTb3w5JkLmy//IuYML2ov8iLsB
3i2cWecRBngYRzlOSn+LdqOfwL+GD3cL3Mxe3yZqAPCjxQdeVq4P90+pwH0oiBE+
W2VKyWSmSkkUYx1TZpBDMmPkJmmkQqd93U8h5bDuo1uLIgQ0/08PQV31xrHiX8XF
GKxRKsW6ti1zvYmkNC2TV4KKhPfKLRoJzP7inTgsiqD0m6VKdErlpmXX7TyoOOOI
EvO4uGNeQw+LjXKzxshdrhG+cJfXVArT5Kxk8fyIsVcR1hdwB4faRBJkHknRi49O
dzww7VMqFmgOhJriSw36+1bcVS1qYR/l/WSJ/WL40gDzUpA0N93IDjqzN6VcCT5O
1VbIdcnuvDGUgwTEVV9dfe2APFe3ZCK9OADS2fsBwLVbwnaevhe5EWR49DG/rVpu
CEK/FuTI/vQrcG7BclPU8zEmnPtXCZCd2EGbmuD3D+skZBN6Y6Zf97X3hkLBkjPu
O0HOcrrPL0Xt0QFy7KVkQukC3Fjt01pHZirFPf6AcbaJPjJjYiNwkE9Rr1RtjQDx
Mw0N4kANj+ogOQTFlddRgijKVVhtYlVTXgGZyoLYV2mHYH0oJbMMSeOunrS1C8md
srGJ9qPjKZY1yabs5paqUGbm1Mx5ANYGJ5iXy0B4CVcl60pidbCAHTrzCtCxvG3u
68wgvBWpq5e95LsVaiQo5oFRf5WgzQAPBuuYURgCP1RznFAdAOOWVSKcfg0anm08
BoEcusngqdpFwls9lqep5WgKS7NlvSengeppI6AvQuaTEPSEfCF/RUeaztJRMAEh
icKfhIW18sBGHb+cN5kHtnnICwWTyXvMKbQ5fosqCn6lXjO+39Z1zxqewo5oeel6
L90prCw3gR+PZNXF5sLt0mEBbphf74iESxZ+y5s+F1wOalLnE8Kxrg+/FwCNu6a1
EdfOAaDFw39+taTo4pLEFAzqjHYe5ns/14Y7LvFL0EebP71e/PonFqKGZwj8+NdE
RQ4dYkOVRbCUnzpduwp4fmcJOu8V/wIScnvQjYLUy7otjJJZmkO6td0JF6dFuNN4
zh/8vVHvl+JCGvhKNMklcrNPfgcKmmGT3iix+fwBog+2IMXA3z+U3BONqOlGDQXR
GVflIUC4tJwlmZzvUzQ+AUeGtf5J/dsoCxq5jfNV8rEZYKUEhe4IsGOClwn2sKcd
6A9zMpW9sIVNfsrea1AQ/c0IZ+kCbcfbTL/s5+71/8FEzNLN8QAAmqdYUBJjiXEP
e7WSYwlgGhhRiA6MO1HG6UEuIzJPLNsTA085wDF4/mL41ZteD26MhPkNhU+UE+r6
ynUI6zz3zsjDgRriUNYvParrq6edzgB6FLiGiPQz4OipRPR3o+tlNwL1+lZ07EGr
qu6kOL300uBVU8BZb9u7qgN5AaffY92lYoMO6vLxWa5/DpOu48c/FTX4u0a8Ec10
olCckdezgi/O+7h+cAatmEbw/Nz7gHPjRlOd2RokICWjZU3C5cRHv/2/zWelZKJc
qXYVbikwbNTugeoRaLYbM6j1WIZ8Pl9GDTgpQUbZQCF52yOiZA5y3L+QMZnVGdNi
O/cGO3wKUjn+44YEOiyEpLEiieLQAGKyTtrKbvHC2oBeCq4lDds+ioVzzQ6AnVNn
of/G0+FX1PmTd3d6PIpgnHvmlTZCAjV1lBkriBkDw+S7srEP/un+QYulJbv3OT2+
CEvPcObYA6K8BSiMYD4dwKBHSlPjJbrBbSUc/lOkPaRNmtpeoHqKCG8nR3itwSn3
8zou9hfez9HcnD3CtUpN6s5J/XSMozrGj0/qrrJbn9VMDq0OFELt+BzXqkXDR2bN
mOUruDnMK7f4C1MPCzBKETwPzZW6BP2PreXOG4VbQ/3GaSMtd/zIQT7gO8N9ubGg
ZQyPE44bO/LcLj/ISWtu6cXN8+8W9hR3qSseRkLsuWaMznCs1NI4QXSPYop+RES/
jMT1yus8gP/JFGTxo5VK/gU+Q+jBR0xzsCMf3WJvXMspu5XrOAQiS1d98n0R4uK+
qgFYfT5Z1/9ifPiTV4x/ihH6YJd2PJpJES/CAodgH341g04yH2sk4/UzjCgynrqV
htsXS7DoOnhlFvq3lQdI6GJuLqZjEEe/mtPPYBLHSi1UEbmtVYsimxIOSWDcX534
Misugh98NisESvq3ENzqp05WkDpzEa7acQBoC146K9s+oP/nGij596MloD6njIYX
Bg1IpCJfTyfkgFsnWA5yJySpkxmnSUN0E1QTZf7ELjAGSbXRHkpdS45JXa58REU4
HhPtLUkpKHajccVIGoBH/BHbRFJMlacg2WKHeVpx4ZqUON7gEzIeJc8ILAXYL9L1
gtsmhuWltgPtTBnx/Ts0lddVuX/sl8ENxG7d9Op+XvpdpKHKWB4WDObEm2JuIkVK
xCTQMhE8NFKN+85QEoPe4zJkfY8CDIr9StHoKm38+7zLkk0JTDN3IQ8DL2lxuyzs
BPVfvy2uSAtSGocV32lKczsAUilOr7o5w/F9m4AlA0sxFmR7RUfQgTPl1drHBtM6
5CJPFVImQM78S3q+LKHWz/zitqnKfhfvmJCRjOwn+qgxrv3rUJlD/lPB+SgusN2P
KRD3ojIus4zLXCAh9sXVKzZFqIB6c+KSK6fa/4wqb3ggQh23SM+eYi74S4vH2Pur
RGWWn4iN282vuvXMmDpeYthDv78wtm44fqx35kbBk17k8Usx3w+ecfP+2CQNTqHt
j3wvP/NhZmE1ik9QfZ+63p6mmdbnFT4/ABYdnUinwVpZDkwcCrdG2FZj9b4EkYRx
G0x9rOsvVbJ1jaV+PwxwevmOvOcJccY8X9aUlOrMuUnHZdDGPMwdMUUl8WA7oqyD
uPE2rfjUuCsLoaXbqaUUd3+/2HHHXhKEgGgpUMaF6lAX7bxDyMEV2nZpIiAdzKEl
vZNj6vANYAOGHo7XRD5O40Bl/qElK3brAF2ndkUTGw6Z3LdPc50nqfHZC9Q60jzL
EvdzY270a/eo9Llmy9waxuViZ7j4d6cUGuf1IoLM/sEaSs1dtkxzUABjpT9I+bCD
82saFVHYTPsMjI7XMHT19PzJps63fHvLU4Ekz9JjWNzyFRmb5Kt1ZnoWwulebZYm
6JyKvMMbLw5EuvfALqTC5KWcEe3NARhGN8mONvcGWFBA4i8MWwLf5ypmyNk+FzPl
H+ZKi2eFY2nyzoUrOIrX8E7Y4XR1bNM1DnnXQnY6MUYIxXAeJXaQpP/LYZpcSE29
V4oYPkMs+S7eQ66JiCOoi9NHPuJzgu/vSzL1uH2XrBtiC2WIfOstMduIogDypbfz
cRyKow1/4LXcZIw3S3Uwl2Mqqm9luBtaZvLaRgcazioqEdvo5Gg2uwEK1GcVEnY/
J0aEFMk5ILmL9rzhBHOqrAF7rvt3JGBK4ZK5lKsMrU+KukQKrfydAXl4CHhxxZSi
lFhRbET0MY5RVy2279ZAamf3E77x2YyipGa7JSoVW93ARpplLInPsuLeUi5h/66S
0xujDKf+R2DooiTxBcUHAa4uWyR/O/Za3usyNvRs8W6JNeCEOVMxmEWsN0F7w4Il
ddsTLSURWJ4EcEmL0EOqpIICUrv347SpS7RpDMmJbabiR3LmD0m0qTVoesPQr+dn
uvQgc9uWKzVcKsr2zKFVNsIBPkCcQEpGxGu07BUaabi1QJsUxciWKhF9tmzIxolZ
DyaqYF6a2pII/skmRywUal+agD5fvcQdvA/kU88QOGsrZZL0ByxpQNqw0riEmtcd
PCGFdDN6BGKdw8yOwNyU5DoYrT4QffLD2ak8iA86iTjKKjKrnxyVtDWt1E9d378q
6dlsd3wTQeb4y1rtLk8u5syn6iHeaM6OnrdJpb6Y0V5+JFAVekQTTgBtaonHhUwD
my7xHggmSIIHnkjPFLcBRjJlK/urglRsu6NMgSBShX8PWLM6vYGNvvE94CDQnIwv
4J4I0Rf2Q6TsIGIEGzKD4vbszaVg2HaY3vsRgmFQkdgo3uNXr7ADGKrcUWnXoESG
4g/MN6qMiO/I/+TWTpUPdeIUNFBQe4RSOWOs+1v082g9dFVPeu8pHsbe/9R2k6L7
9lVmbhCxJ73llgVrRU2FJ6d4A18+F+ABnTN9ZxvxuNM5fEHcd4DbW38rgxHCSnbD
TgA9wWjKCxGWMSq4+Ot1nQa2rn3LL1oV1D9GooMqKTThC/kZ0GpRN7EsjhSPPWAV
WZu95GjGO0Sj5EnOwW4YTtr7FI6XZjDACsXQGYuqzQJy2+y+XQz6lKtZIwfaAzbl
bCqKucI7wvjYTMceCxlNsLuZxd7d5ZVr/z6XlnEiycJ/LRICUyI5f1o5KTbjiTDs
pRtChm/zVeaD1VD3LWseS57ZAuETrz4AmmS1fTdIBb/lNqdshnYp5I0vEOGdnWgL
LTNA5CvUjiwRIrA/jf528QFfj3ksHLwq9B4kmNEb/Uz60z728OkEZSP8UZduA6It
BQFfFxhf+817rts5EE38LwiPSDXw2/9u0HPfpMTUvNC3UtfHLyjxihQ4ZY5eQiVL
DTtJuVdLjdsVOthd8qOobqsVXH3yS3TC+W9A0Sdy4Vkp8glsgCvlI78RbHIKaRAS
oLf+HAVjkOqqSFS5AgCASwaOHUFNbrn0v91lnycvSLdcE2E8bNjRZy6sARt5xWXi
EFwiUMaChGCnQdKZIErWkfk4ia8rttPHWzwLuuycGQeDWUxXcvIxKMg9NLTnIAZo
9Z/Lrkm5ksNERZwgEW5hPjQvj+jiOgpwjGOrx0kTzU5CBClQq6+fylTGXNRAB6kS
IOhlVKxXxy8xsB1onQOF+40D8QFWjqreIPLB3zCwxiGyQcrzJFl57ajT3Ip9yju+
oc+kiOAlHFcePulrudONX4j7tdmZHv+924FjHBiC/pgcY2PvDy3wMVrrAqFF7ogl
uQTeAtcn7prMEDsJQRmFvgXZaq5AOR/DEUltR4CUgUmxep2IkFQ56onjqy5c6bjk
Jc59PSQG4MlQHP2Hcn3jjCmOe8A0ea4JR0jUWEOsjIL3pxlmMwgZp3JSjGpmeN6O
PwY/FhD+keeboY9/wqSOhuDJRpEc4O7v5BGJbPdJkvv6ans3JwJxX+Vi56sE8myy
bOqgztHiiZLKVWhOB0hqyNZ1PhBcaK/1DkiNhiWhiqHnkYrxffxATLHImX/genSD
x6Nft9zdDWA+AwN8XViVPW6YotcDjIZ/rj+dYRxC/wfoP6Npga0ah4vClaaeDYcf
xDyceaITIqV6BFAKi+hQjB1Nb89CPlVtiuoecC3E1G49OXz2zxlIQNBxOxSiFKXH
WSdAmlxFhMVNIKJor1eoYyR4s+KiBjl6CpURJXXzbUMlfC+VshhzolPSBmShM7g6
X5PjBvcaX/KrxucLSw2GrUI12gSm43maAh98RkOygqCLheYhexH0zvOsAcmu5WSR
vj2nKGOPlfzWEnvxk8zp6heo2aBATlQLSzYk68ViWve78pCrVaEDT3rEX5UfaHHb
QzF9jkBBKCv5AGM5xYGKB33KSiW3nr9seGNY1sPZ9wzO1123oDyN4fBVWbCPBGo4
7HEhd+YTRR0868tAObbN1yT8bU1NL2b6uQSBH+4+4KBPzX1YO7q6biwEwelopKiv
SWs9kFG5v186LNdHP5T7J4WzKRPijz9aiqJsWFaIAInArJuKIWjT0dDPOKYZypTV
qRCzBs1D18N5XUunsifw1+mcloZ8HhN+28U9uA50Rkg/akfT9/fi8vzMPKu/sv9H
IZPn2vF+uxQLZNze1vohIdaqG0zQz2gYjiAb8OmX6GbHd7HELFQRZV4UOoUiUJF3
3UIWVY5+DvHJUmgwbLyAR8qMlJkzbyTY2+OXRrTcYBBXFToV3OiwKkbI/hAdOFaW
bazvCO3hJ4sVZlR2ethbg9+2GYNVfhTRu+sbZfMK8yVhcKO6vVUqSkn6Vx9p1nFG
/3ofLO00wGHFqsIW3p3Qk7+BM3T3oCxwiu2KerRLtePTI2wI4tatbSjTgHeekE6s
5QHq9XvrDiTL53+kspjLxlTQu0+bCEZuVMBZa2zLimKZt/ihZTi0Mavh5WG9oqI6
6UO8T25EUC4BmKF3AnTQnu1Ub081L7L55cSThZ0ZsnmTk0jZaL6GHX5MEliLHmIg
ERXcDj9IyDDIc8Zr0RAFKp2SSGCKRibtFVE1B7mUrPNoqeVYlDowoE68/bQ2Vndc
zbHMnr052SJ9baEX5b8YSbZpfUNcuNF89PwCzrQBOM9EzByF5polUmo/h5Swo9n8
Vh+uT/gDC9VgdENWJ80KZEWp0Cb7iMM9PeXdz1R3T7+5LiMKaNx537dU8vWzeSJE
Mgh+PO5Mu2j7aFA8llZN7jg8JOZcsFcLagTp7T2To90CSVOtwdkhdJMN+jHuukhE
J/ZYBNiFqWygD/kUB8RNzZgGzR2yEbrEFhqd97zrV4F7OOJpAPvHegPQyAEDdygj
SH7d5XgYLj+XctCtKemFLuIT8XI9EcyWLPom377pLcIuvRXbcpMurzS24rjOSpfH
u28FqGiKkibS2sC5Bdxh/YMxEXvlB67TJTdC3IbxHH9RCKrp0SbiccRxMJ1Qae/C
vo7NkRLKwAsN/uHLmatngQscIblbizhALO8HBAjDN8+aE7oNE971g4Hje7BwIDef
rPRMovBqQ4tTKWVSTIDj7H7fL0BwkBs0Q6kaTNE3l3bKQ+BYGuBmNR+kMB6bk5v1
o+bXcHxJDVC3KxhXNW9KtKf8tUOTcMLVoveGEnKdaAi4chD4irDanSmQ8csVWcjE
tVzFte8enc/TyKVWpDtLy+9f/+TMkIcKLuvTkzrxmRtwAdq0glMa6qCdasD6+P/d
6azRP1McEEMZoILmfcpFZuBdjabdWJ76GA0XLWBSmUXQcmk396wP61fPrRs6JMcr
Gi1Pgb+gAkK5WoBwAnF8DdMZ1FmIVkzImkxY3O7xt3MAAopTIn5D/IKXRnvYzSgP
z/ZpVuK8guD2miB5AcNdDl7iNEx0AZ2nwWzjZyWlGDic5xbVvkQD/w+Qv1/RAJ6p
OdXjRP7khQEJ7ZZs1ElI+bIJd9pshtEH8U3P4Ynw2niNU+I+2zqziQJgRrUcgREW
91LxUq7hUhaG9qwApSZOJBpVN0LyhLEFBBVIqTP4QwcaHOvSmdSXTJauDKilvjT/
zBErb1Dx8dTbI1k9Id9vjeRy6qnpjCGnj1Nn7PEN7G6XAPnYiK4+bCHI2t7POYWx
Rya5jcG4/b1RxrQiJd7miDo8Jcgc2WZplkhs1HFMJkm8pWXZqeKlQCutSIpTmVVb
Qdj86dNDEOO0cfWYKUY31XhUgt5Au/feJW3lxnwFBrmXK0dc9mmkCB2uNdAVWt99
ZF5FxmRBPjtqxS88b2wPL7t//CfLtc7xkL5REwzitV1mH/FuG4Fn+75A2vPecO68
2seRFdnfn4skyhYZLJY+UtycsBEwzTBF32nhlNmw69FFE/Z1Q1HQzQMQyW5pUi3x
9PL9NBzJJecPqPFILYohNeGjhO71Ry43WKbaqZ5vDWB9UkbNUQNtH5IU44IZ0sfy
FbXdoj4tqKrhA7QUAbkDej0V8JQJ91tn7Vrfyvr7poxVNl7f+D5Nzr5h23Y+oqYg
PtyVMmyBeFYYGWlVK92J4Px/LOqoboQmeUixFmMJJvKEnv/M+hZJQ1vSU7hge/TU
d/iUx5LveiVBIIkCRTEYFTnHmF2n3sIVunsgoS2SaU7Sah4V3H2u+0dONtzLp3Og
tg64AoFccLa6yV16VWrcEm0YxISPr4w2N4/JL6MOcLYmgMklWGia9LFjmso0XOo5
Kp9b7uecCqk2VwmtkCQfnNEpaps9ptyA3wgs2KRzY61aa3MXr7Ln9u4gKVOM07PV
XcpKSsd7C6n9GjML23g9FP19L2oL4/h3ELkHXlTKig0r9eCEZCmcyCntvPk5Zgwz
CCrE6jCJ2WIHUe18vt8Epp4t8OKjM3L0jBG/Y5lCyH8rVraxf5sP8nQ2JHunkSkH
SO+lUlsAnFr2xOXcg1z2hvtF7PwH/GeputB3qOuJoV98l1s31Rl+hpwE9bEDEpbO
zKXh2MmsTwpfhKaP495sMMsZCQB/j57Ls6DrAc+Mmp2e3sjJzYCW20BEOTrDh5pS
s+tkyY23JdirvPaF68WIkxNpoMkaPWrxlYyVoT1axt6MQJ5xJXMWwprgRkhqbK0f
eWCvREN9Of2KdYMN2NcV8bMGCn9i61a+CLQz31TUt4gqGajKTK5nxskQ9XCI7jpZ
VaBzHLMDlveMtPkw4Zk1GqVLwQ/EA6eFYCNNJWt5C26b6qu8Hmf3CcWwNpn7i9b8
cEgCwdFDZFP2RLXqpsLG28jrDlZ+44qcYqYu91v4GJwYQRsVXvfmVVIZSw4d8d06
9LLM15/JWqbxcyjF7JOecZdLTQcq5aPBDcP/Qv7KfHHKxF52pwjsDObvrFYer8zN
IUmAyaifGvl6s9eWDWBIoxvX7t+L3XxfCNzPnXhsN1GyEZPv5ZfOHAMvtgOQLQVF
v7BFzg3IKYTWQ/AvJNBexbAP5gQlcNI5wvWLI56aRpRALFacmHaLtsmFWaQGWqYF
454drCVpcbRJd1/xy2mk0RLmN5w3bV+bPql3W87PPM6+0w3QFzN1WPe5jy+/7eYi
GCl7BgSHOcrzLLi2lr56Uj99JYCB7e3+xJmZcmS6bdcU1dGFrpb3wFplbXL/wmkb
nNvQu3pZxX3JTZazL5p+an3WDpaGF6L7Jy9vRjoG0Bo8BV+qxkB8Eqduwa9GlVSq
462G7dZFlMTH/DDa9ywezaXny+RUB/d/aL0a0kxQdfyZTUaLQkOX7AyBm4Fo0yMc
E4s7znVW/59Uzi0z0Gb9L9Tw8XpJ6Z3D7yWB2JC6NYJhkFeKOkdQJeXecvI9w2zl
pGGr9FynwFaPYt/a/uefeajY6geENd3Z7uOyFcxVuFdHCfos8gxR43W5BLKqPLb3
oo0xFUXxjzAGXPJzjGhpOWpUAOtZpU+gj2nn3VBf/E+R8pJBiy9bm5/syZf+LCsv
afk9QO7tuAHyStIsrYkM4KzAK1BVJGlmMWnjOe1numA4Ljx/Sm8UjydoBwKqT30e
CYAMGA4DWgR+nwT+1lMrSHRbFI0unaPDWRidIOleekBrZgxCPqo/B1WRYyrxX0eF
b7Ymqyv/uGGaTzTCU7P7s83FQt6UqLYoUtCCjCeB1mv/KXVgQEgmhm5LsqZaxKoa
3rsyXOODCKJC5RZ2mUs0a+EVZO10Zu4kqleLHyriqvxS4C8CsZg/1BKJcuuqqhN8
BMtGCR5UYDafIU0KuRnFHixcw18Z3e1/50KQS1bGSdM1cHlsf3/J+Z9EFj+uu54L
KRzYXth8eAXOA4goTHTj5owcsB9UEhIZc2KKa5f9mEDT3077AB5hiYXBhEby2oml
i4Ld+FqvW7Mguu7BSw+bD7WA7lK6RoiAbm6lsVDh82Url6FiGRcJhB4HqD2nS4N5
oajep93lqf+5zi/I86JYB61JiBBQr+M5fE1FnuwlPsgohHH/Ev6UHeHVDbBh6V2w
XK2FDyHsAxh6hUga3U2/vVazyrdejIxJBZGO3Vzub46ruzQc0Sz6jA1xJIJ0Kk5z
kOJticluSt/lgBUNEWyT1BXaNUDONusbfd+7mB9oPtXbezwRgzANWeP1MBq3jQRW
LL5T950ojamoyQg5vi0BdPtEy9z3XI2dmS5Hu66MsQlDAmCZDjqiN0Hyeb7CrPYI
kTu//sTQu/Ksz+Bf61VnRWUzICNe7F9BAOgk93ijhU+Nl+/FvJr8MN10HaJa/SCt
uigpnrUXvAtHOvfvLEV2C4WnlAvNU7srNB7nkPjOF4d5HAR3kiISumcO1VN13mn1
e+g+vOujs/IGGR7hMkJO63LhZFsiNVI5kZ5jcpoO4MQUCIpGIp4pR5G168iLRqNb
8XxSzUvO3bUwMtCCcLeyWXBvyHZYLQ0G6EVSXgfPS0YF7z+4tHafh/HCIe7VWXUT
9egTAMHG5oMWiIHx7B87gB9F2aOffogA0VNytyjF0kUWTzIFBWfQ2YJJ8cylR++S
zg0TRBS8XsbFhtJ5wzwZtYei5S1bklXbI3TStVTwm68PO6el1eTwEw23XnIalUSZ
Xg7i7sXhlwlE7Ux1Wwt+tlsUM4O/YBTXc6+7NPUyLypODDSqkSgLMIDPFYKcQQib
Gy2K9UefJVt5VRVybEMp2/TjFiNyv7TWWpmYfzoLpXQD8U2kmke1tNauItks3MHl
ezJB41TQdBv/ZV1wthKokJzThDswafg5+HeLasvDkxObfG2TSYO7jFT0PutYGECz
XGFCHCycN2dinlwWMXvae85vE7k0qxB/CMVu14JxZ/za6oGaYa8M9/MmEQqSdZZo
1hnoWTNtqrdchyTBOI/bcvHFYd5CMPVxPGwWl7BMJF6GtHyevIqGAsRT4KpnPWP3
DMENv8zRbKRi3FZ+Rt9y3jysXA9hPvrf10Ye49iyjjWhiTKUBNLQeDNRE5GiqilD
6TGrP6bvNK9iX4sJFcKD8ODRKQrdLVtnsbyGgM4ne+clZWaRj3+Mgy3l4zpbikwT
sztti6NGo4FtDZpMB5GDUVRUricxS3bQYC4Ve4mWfuDvZ/hv6uL60ghaetxvDgv1
4C9paU4WiFowGq5QmFR/gfcsMPTr19ZsIjq5fmPjVhevY5UCzjpx2ylRSUSkqmnZ
KllyPN8m8Mbb0ndQjYRGt5Xb5bS6vwuqMYbhpNCFIT5lIXPBGlwQ1qdTlYTgNGFf
cqQH0gZEEKniFNQKNYsEYgvgasNreZkiQW8F6PcFmP+LaF4jdAcrtg2FGWBrFfWu
kaHOuKDEgpzGpy/KGWUH6UDBg9oesYyfpSaA57szQNENQzs25q2ThhD407trYxYp
mCBlIA+SsCa1pf0gdTMdUG4sNVJd4iXIfxe/TbuvKc+sWPMH1pTAG+1wxQ9qVUwI
TMAst+x4aYALLyWOB/AWb5Ji8DvTyYdx20s4QvGrow3s+PlB8VqCrXpOLWqjwley
a06b3Pru8TVW7uhZbd+l/csQRjGayBohkxQ9RUbdkofTv7yswZzwVe+2UiWvvro6
ORn4Oit7vHIGFplvvp6PTQ3MC3seCQr+8ljtlJZNiUxTc2kOs7b7jB/Ai2llRpri
VKUZDDVaVTxllWhRLhHz3zuDKN7X9JP2HKUZFN4osUCIZHEwC4tRjU9R/LP2MzC1
NiKPXAAtYA2xjWJaxwak1ssiqTtOJ0vH+YgnbofU4usLki1ZiMQDOVMNaKuF/vOq
IJf0MHfOV3gkO80mWetC0a+/x3VTjPOYN+U5ttkW4RZ5GsPO3ru0kJrsBQPxVAyX
IXmXJrEmo34xBwa/QIYNUiFAiKqrZU2bPk/UILYwN/rYowWs45tIWskUkXLlFugy
HfwtRQ//yxbXa9HFLtoqc/GLL8iDv0qWGClHqZvTzTpiSvQkVr6s8Y5lblVeYHF3
QO3T1UrbtH+0ndzoBb1SWQRu6A5XdXIo+MctbasRr3DIhEB0MKZPsxjlddHybJwj
6bsWJ6zwI36UIO0mZ8VEwiWse2SQM27mX4mtTh+61nGuJi3vnLl+C+mup8xfpw96
hdYsdM/wqnsK8voTVnCGgToY5U8ydXnUqL7Lboyn/PP2OBN5CopO6f65WvVuTBTs
2cGXnS7CwZrbI3yxgR3CzqeVRsh8csNhqGaws2CnJH8C6Ns9+s+mt4o3s37Ql2a/
cb75LqncY4T6COoESPCsNt96jMBkSAdvisHmdGU7xSjgnYKGq/teqX8cgDE+mlbw
QtZcCuwVt2l0tqzo810wdJPl2MNiyCWG1yrMKTZs5sPiK2MNfknYIuozO2u7CmkB
NTs5RN2zj2Opm1MYiSmRkuo9h4vqAn+0BSfNS5VjIL8gt3hMxTfpV6A2FfiODKq8
+xkIhT51k2ARRaxJUjfKWXU7bkI1AroFr2F2zg3h9MFrk4EoSZHPHqfr/2vmflWl
7qy3i4+/+xZVGID46o5KcOeWHGhJBkpXJvEtCEZR9dgZGEJHMil3ZOI3aKvyrnWz
NUoYf7qdU8LjeGbjFmtloyrpvkAfPoMGFDQKr8StDZF53xtxMuPuBWu26+BpYI+N
txPQvogiDqnT0rLzIEFWJtH/QulSP7zZ4ac1i1BDgv0/RBAYr6DGDLFHPazeDrSc
IxLegB0zOuXKE6orbtqzW+Fh3TyhvfsVpOQsLrZs7a49zk/lREhlKcN3R28abV6h
ULndMWaNtGWwB97WRnmUGQKyYwNw/368oG+F+hlCxHvvRxHzYfMZYoluklXDwdJW
0jfHpxh1DLBhpbQ4tuTU23pLyezYaKIgYB8UUyOHA90uqUOtpXE6b15WHfdBWZZw
QJVbrspYa9fErcqeWfvH8DGbcUWZPT046fs9POlPIOdx1wtOvH8Uw5tcfJvRtxGP
/Mf+fcP7MBUHSBuhg2NoXLIQYTbqk2XuGt6ofUWODeJth6dLG2QyM5hnhKWPHVxd
PRGjLgm2W4qp9fjGl3iBUJlQY0QHmaDTrT1zpx4YA3/J106ykr9f7vkpBjHQn9ZH
nKcEWWhX7k/62o+s0gjOR/hayqErBnWQudCJgtjBg5Js05O5m9NWSC9HVHEsQyVV
91uVApY1SanSLouI8r1FAOWGabIdi4KEwBfc/HzgrY4mXoRP+T35/+RDSLJtZptL
WxMaixEvVNISkESvqWtj/y/hOS3ejQuZtJ8C1GhLSDTfTiY+HAtwKJeDT0zjbr2a
qoD275ljL1rXOHT2+CDD5sCgP60bDBIgtHg2tEK+xVXKFv4vFnCQdq2GX2DBr4pU
g7fe4LQjGIN0KSULGOExmHYLrRkv2CYzhyh3MKwUG8zkF79cJN2DcE3PiGxIPjUA
df8TSARF2Y8UpurQQlTp1XAk1nOghF5i4icAY3lltCZ5L+qmfwdzwLpQ4WGOdUgZ
oW6EQnBpvgoJmInN59uJKWHvEBGpxo84OaQZbKFNbAQTXEpFeVee370ruH94p692
yBEa3uJqxHzO9fwo+k2JN/tNw6yQ0NIq7EIdeKRxlce/v/G5eYV/5k1tuYwVzIpo
Lv3c1dCszB25bYwHYbgHIrAegaDedS9nE4C5lBJnaNnjMr69ksj5bLVV1dd6brjY
sh2v+zIsENy84r712y7Xt1z4DqSFU78Hd/r8JO9MrTqOMCoj0BooCbZUy+K86tBU
LF/TcIwe6lt5hTzM4N5RCY9KoSAXBmi7mt8+HP+faXyWl9OTR9x5pb9pwWO8fehn
+REQbFRRu9JZDY785M/r+zvib49G1KbUfWqeZUkdc1uNRoJHPiExBJW6nmO69SPh
mHjdzySzx8QsaO3mocXEsn5i7yIBkVIRCtM0sd+Dcp+28NCx28p3Bh51Mem4GSeL
G1Ahj6CVFARP6+P+7zC7bh5nme8oeYL0G+aGUPaopoMMtJJG1lKwpTOpC/aYdAN+
4yF/1yB4Ds6MXDaX7O5CUsDkNCj4GegxdmehTn4IFo+t6o2B3uCyE8TnkzDJRifw
fGQ4vGwi91hD74leI+r9bskaZBdKajPI33pr5DMpJ4B1/O7G3PTvntRcqSnfdRb5
/8HYnka/jMcx8SQIs776du37TgtouJVhz1XyZ8MWb/W2S97SOw/VH0MNC3cqeOJk
aeqwIalpGQX36a8rWY+HKjiYfPapWHtwMl9HlhlrV49fczmTJVcAZtZWP5aGlSoq
73Rr+srtck8rXRpivpUNpNIApZ234xZRZ77NOHBDJMR9sVQv0oyP0AUcoJl80Fzk
jvB3MZ9oWyvcGBWPbi1x2IEJfbG7IoYtmCyXrP8/FKy1JGexe/4kJf9QYIDNcm4q
/rvsrMBTiyFE2cV2nkSY1lfmF3WvrG4aJEevVhyLSJCAWnQPDdeqWRxrwQa0/+Tc
Rmtkj+tWJyUzcTsTqVs+0LzZeDtB2EqI9rQ5z2MA+6itvmk9ixD6HPL7hCz/5eFv
MXK+nJPOXA1EWwJ+Xi9VB6rArRPdYf5IRyhy87lz57wlxUEI8uLFYqJLBiMnXXLd
Je560UIiqmHqYcU3Sh7gaG1RIb7aj+Xm74t685xwmEwawYnUUSscwVKv+Mttwsha
n0Ar88fXK0Ex4J08GV7OzcvkXUHq+R6A/vHlBmUni3nIJy8Dk5/sUxf3RT4JcbRH
VA0JeLlVSR5G/gI6QJOOFlG3j8+mxKy/qUwmwNHdl2YnsxfeIkDoBFoWYklhuqAZ
YbwXOj1ZBZf50oWIhVDc0FNOxajCb067xRZJq+hotUAPlZv2jm0u942/Eaw5Kb3F
fk1cO7pv5lLinnI/Y56s0z8I/LPW5O5/ELIE5+8dz9e7FZ1LiaEKNgUcw3ptP6KI
gutZKrZ7eMz4PHDD3JB33rQ/4FBNlkSR9nQLBtviPpSeKwHqXWjlkH5FzDtut+OX
EToamdvRgWticaDzPq3uDavZKNMwJZNZ/3fRVmJ2iGhiyeffKIv262LFvKuxTOSE
UFrHT/NbVqp2VDIwLP2yE44h9fjYywlBFq3Ihkx/FpsRcsD3NtmkYBGWlxsHaZO3
ZJvLV39MuDMaYqcmwFRV6QqVmlI128YuQ6t8MCKtgJpbvWcFK3fqcV1pBa/9H7Tb
sD1SdC8AZgZfXT3pQSuCzz9G6EbrkiIA09l0vmA/QV055Q9La1hjDoUU5osylKwq
hRCnbSLcHfCMIjYoXq6mZXSC+4Oupi8+JvTk9h+Hrn0hRpp3ASldBB1cnAwJFFsr
4P7vnlrET5UsZ4m1wvgEXt5KbW1SquO95wuSpw6/V0kxC7leRUXQPwWDKATDW0mG
hLZYq+lgnlkftk9WC35rXuMLzyy+boo/o06HBDkr1CYEzMLgGKny58V/bXLcgD0K
8D4PlWP6IK0K51UdRgtFXeFlds4K30KYKM8RziEd9lZ4Mth7rtOyXHaLG3tFKk24
bVySjCHe2lTpH5260qimaA+EUKH69qZF0xlByv9o/n+35OHnU60pWGyrAOqvIzbx
G/+UduH/qRur5oMCwtCTWUYrRM1KVGYm3/Jak+LKHmIMEkz8W4hfE3fHJHAeuu05
XAOVkx03e0BtKHBRLr+h2/d+7ofu1ZyTBwiPPvoNffxohns0xMSB0lZfjOJMCxLq
OOT6MAxD/7sLF4KOao6owvLGbbA402Ov2ceIJ73L0fwfWytz+JRsSGkvqfbBzdgg
Et7fhabb0A1EcAPzPSmlRQmKjQQg9wlETcTz9ymdxgPwMF0749Cgextgi+kKLaMJ
MpuoEx9dalavx3vtdENz4qLbw3OE8w0MGvf55kTkpPeWBq6x/9CTWob67MTE4k2s
H7GJXzTMocrwp5lat4Kdm8cvFcP05BPmhjBDOFpGsALfJfnTxM9HdS2NZrim24WW
INWOinuBTM1BjwobcpVjEmjOU54CCLLd4sAqcP9SiKhVlgzCO7r0REIIoN3/NzaO
s12s1udAESkWH4Fq1Pb24VlK2blRz2eGjrpraHGtn/HxQ81tTDXV59h00fd7l9JY
AJxnpqgoE4Kdmv+DJzio2kF6hNawmHRh/v+Zr0wpmrdRm/gbFlIL3jK5wH9OrStu
iBq5TkFCHu/Uce6m9Tw6gQIihsoZIFDbP9ihEJhJW+QYdpz6fP+4SKAqvJDdHdds
vBI/q+ffSUkuShhpZq9ii1bMwo8thMcp8ObNnORsOcrrUXyHlebFsxfgBcuIn0UT
oi3UUfDotpLoI8oteaMvPFJUoGfrioej7eSDPS7LLlySKCBsQ146jl0vCWbdlW8C
J8i4tKGVVmPlD9xtBef47K8gi7yMcudQ3sojkOaCLeIakp58l+v5QEFtCG7PJhmf
RIS3ukuHbCKX1ZIqV/YocDY+9QS9Bomv6Xv/Lb8bdIbL+XHQi4GM4EtjNT86OJWH
coYK+IYV+Zs0naepOVxE2pk2g7AkawY6OAb55voxCHamFBrkuf0937ObtVoX9pB2
Vm+jGH5J+11D8KHN9u3pslG2Gg3vP373fOeEDRDbzW5iu1Hf/99IUcPiECuPdIIj
NSo4CaZHdaeWAIfI1prIyw18b1aQjGLT1yTVRwD/LpvHS05J38VsMyFUk8YBjiKw
z2VIvMXH+oLeymND3c7gGP75nBmD7ND8CnIk9lz69AwUcrA1a0Pm0Kj09QJzyHdI
UAEOtIQ1jEyME9+mJorsVZ5lf+sEfcK6J8Arc4RnCB6uQy/U+qOFN34jg1phMlOo
833TOaqvz7XWkjm+oIZsWSU+XAGeLScijiCB/8T62gc2T+V9FCpMCVuI9ngiKIbA
2M6aH9hkiWYmrDDgEuUjunBvXwgZu0whv9ZTPCFf91ye0aKCsMPef36Y4s6JB9Q0
t91Ek6/NDPIGub865CO55/fUBgZPLq2vdq5YqoJAfUnxYUuxpxAFDujeJjMvg6Zl
xJC8ho4r5lspgM6UhrUQC/KbICprpLm1O41oXDEWgUmzGLLbcQEaIWsKFI6vRbpo
gd6Ylsi2/M0T3HGzRMItu0mMGWEZKZyWnRtLtYEO243oeYd3SVNTezxLfY+DgxxC
aoTt4kYUm3eIpXnZlZ22sAk85BJ9j07u/EX8EzDvdNVBTiqZPrmnHCvyMIahe49/
TWIInOF146qh0SI3ydz46g/j9ivdsxmM1ZMITaoKNxPE2p21vrlboomndT9p9DGy
7xxvNXq7tJ2UVQTEau9nxetw8q/9Sx6m0H9MtdM1yjBnUSoxuBGeyJpgAXCUC1Q8
pQ+Vtx+o6rhTEqjXphDlvjCn5iQNzpQFhTaZpVw0AIHTa1ivNH4d5/LdmT7aP0dG
H/aS1eaD3VycEIsXh6VIOG0PqcNvVTO5LYD5OS/rhf3FAogHl2//qV1VUtT27R00
M63VPH3jwm3nY02QnAqu/P3BlD1reHAF+87yzVwkuUWMCQ/m5i0q3A3itUnSHYZd
qn8Wo57Gwx05R8gdel1xAiCImWpGHVD9GTZGt/jpczcRVphmvnC9SacP5qn6n0SV
/kBg+TmJ5iZgPZFx/Eboiuht6wSHz4qUTKHhW9sI446zy+qlQ1zwTQPGIRZLeCvb
COX2NuqKl1stOBBZMftHc90r+ZnA6vOiG3c/XYcmjKmirMxz9j152sJNpD4GebJI
V3Tet864t4TQzB85eSqY+DS82GTZerLphUIZ8JEQEiH0skc55SCez7hjsdr3qznT
aSGg1DItQPtdCXf8iXrn5oOdzkNi2rDj7szALSV4wFIUrzXAxtIjy/uKSF0gEbnt
Jd9A8++azicuVFYqz7u/clJa9DVRBcIi0QCbXpQZS753Fp8SOwhJDwnf57fsX/Xh
aEb17xonqjdYjVagq8mZO8TC/2c7rHx03jQV/IeRjFh2jtOYpSGwhM1iMa5SYqR3
iUKiu3afOF0DPVWu0KY8ZMKXzdb4YWGPxGVzDrSN0sZfXJ0PJPTpADF6pEGHO0K+
vF/v6Zbgutz3Tt/BjnVbx+4ZY6ywn6LxXVlJhjM2Q1+i2xZ6A17j7/3zN+xFpiRL
MllF8ZQ9q3tspj/rz89+wieQB392NPxDIiUN80gDhkSlPNplnk27QsFrNI5W+ogr
P7wRDFaXIfoZ0qgmNtqWD8XmAIeujIRnQ4OipY4p9QLSh8S2wEu8cIq2+Q3A9+Lp
UNTadSUlvccJ835eLPw58AC0ze98CZyPJbOxHDnBE++T+fP7iDPFj7nHcrc//24P
+N1zr4vKEwkM/gbaf5IPAoT6pKhAQ8GPqvzk+G+40lBSfvValCSjTwVOnE+YrfPC
NI+Fr8oieBkZKQh27QVVkYNxiIu+ll1Zedw5cCrBuPVNZWVFtxWvATCGp0QX8EcH
4c0OhNhyoJR7OTu1QoBZ8LktEsTVLlLGiK6FvSTeNLP/hebdWvbyETIkokgnoqPp
n3Urgln8OjryBcw+4Z5k3r66xAW6PBF1c93MVsUJ+n9y2rlh4ERJPyqMm8fDnJ9Z
ofWrwqe1QrUcnZ29UCBe8VpaRQI7YdsFyVvIQ5Sy3xiLojSxSA5dxDb4NHYaqCpL
F0dOJt8GuJ26gCFPmjSMYI6ThRJakGdz8YM/YuyMxtd1mdGVOHzF5Z7fYkayMTbk
IfHS4dZJbYZXov3Su73AJIX2GTlljkpHMfbG4KiLIU9KfQhEPtxuIHlNmOJrlgbJ
2tC/45sY+8yOk+cG18r8qYcPWX6zp2QeBKZEBOvqrPM0AFfAqmkZAkk5s8M9EEFe
/ymXEd1YhgLOsU6hAFcuaO8RtN3CMV8UebayxzPtPOtNnsBt2HXsEAOMxvjLFTpf
V80KaK2lc9DoNdg+XavMLHqF0g2WK1LKQp6+7KmDYELuSt6r55GotEE7kE2I3cWs
WoRWAHQ/Dxm6ZOMxbU4MDwa+iWUdSEqTYh4DdVvIHZ39MVMqqD5981nLEBH4zpVx
L2KLKcoZQ3Vmzyv8vRuYuJHeeTVv4sOyGPBUaAOpTNTMXpe545l16AhEE8K3cD2l
0zQxLHJjqYxD+K/pl+IHs5SiEGoPXKu0DRlE8JKYdeG+iquRkMUQNEco7E2Xgop4
HMlJ4vSimEBoHTexr9D5mamcsNBWViz+v18Ng5Mz6ewMPE5xTzEktsYrL98jUpJ8
wvgTVStDy8P8TnM4NGArdk2lg/na2nQwhFXYVxmEfylxfDVDiTMRK0Logj2GiuAj
ifqVIKpsiw41G27E5wvsvxJZND+obJ15TVvlCAewDtiOBS4S1hxgF30hOwL/u0y9
3NU/5vXjIJRFE9u3MHB5bQg0sJQu8ECTNKmQoJ5r1bH/I4uAXAuVh/6+sF6gAb/W
9UEwpKymsBF2VZF+cT8V3iAmymRhdl0odEcsupII1afDK9JGluMbUhyaGbKEKbG4
bIoE1mQ4fmawfacdmDmxB2MsCpBt7A0UrUUY40EbXFgB85kSOe+zxRO1y/kq4sKG
IC23+KU6YAfg58LHgQOnhfBA0hWN8Ci1eRuxPlgSnWv8/sju29xejS0R7I7TUJhh
lnelzyDcE5xpUJdyIfD0SBSgN2lBSisSmjf3zKS2nIKC2mV3OzP9S+eJ0cZAFzGJ
/hBbA+vewe7TUQFYM80KVUDavBq9OYht7SwJZ4R723jOeDgumM2bU707tiu3zrwG
SUpAdcJafd8Ymqm7F5JR/RuN0Z85Y5AsfAuXUC04q2CXwgxpXgXnCuoOxeoRdWZ/
p/MnESDkihVhbt2Q3FJOz7kjp46uLSne8LaldNTE3VcMsl3u2B0dp6tEuxCJriKl
0wzUobyY+DUrp58rN1KUNiZJNofCamRMrbCbj8+BwWfl+9sobbVIwTxsxkGovwq3
BDPot3nEsapXxBtI+KLwpE2bJL/weZFZj7Gaum2mGPmJKCNRXvFCMWM9AGmDTbpd
UIKMGIAVuC4AD/7Z493GNmkRyTW0xlW+v4R8WVrp/L7Kc05ccLr/+a9hmEN8fAPo
hlk/vziorjNaAKXIo1zeTGyHdIXBy37VthzePbodPUxn/HTvAqWmGJHYQEhibVYk
dPh2gcEnx9kUgeUwivtoKHo8oUFvG4BjPkz/gmo6RtB3a/heCRTIsItJyHFY0Wme
0CRF+DWtzMy4tdJEQZ6X9dT+3hFPNzFiGWPexijxURA7Z2/7LzT1c15cZUpDgJYm
VztiAHAI51Va5xP2NoE6hBIrCWKmOvjVRXaItk2OSDpyxBnjodsHxyfy3Is6y4eo
AWQjSlh7Eui0+tYwv75Vmpn+Iy91xDePiN2ZGFWrePowZujdz5wq6+76J8TIrbHa
e1TcMz4NzgYlojMw0AluvXv5/jqsX8ZK15y9oCxYg2CuRCSZIUKs95O/iphugMNR
wLMzzx6mEyAd+BqMR26GUc7wOu5sdoGEZXAd13p1X81sAAucFHOSM7wQIcgUlL5a
gQnwKoxSdS1utp2gOqy+XDttFAmbWOURr0MuJ4cXrivYRxW0boYIOshzlqsWZC09
AQRt5G+J/lsFY2ogjGykqYWIVwOtfNyQmoWS7MBAXZp4Zzvbdwy8Sg1ZOzn7nc/D
fqzT0tG33xc3sj9syNZEuXF2PIfa6g8KvDrkWlohhQ6+SqJvR/+SbLMPtj7dsln8
tPKn6Cr+WHuedhTroSTt+U/CinXSwsQcmxN6uyCMCZNPnTMNuUpHv6N7e/QNpD3C
f6Gs937ylA68ucnO9tcCDei0NzQlGAjyhRjkmJb2A0Hnj0SwQTqUDfKZK3wzxDOo
RsuwqEtXFzQF0VpVJXyib1cKw2Kd3K4/NsX25zcnwYR94Sh3NsYyEtg+6sWDVyTo
6wLEfMu2pF/gtL8sLguYi2z8qd2tMcBAbWIZSLmggD5c29YlF21T9469h/tGZ0xP
AaplxCaSweoRBF81RKt2ffmbQG+n7XOmgn8PYlNUNDlTmEb/rEcVlJBAVvYrSpLo
muOx9FjkzbUpXeAKELe1KNdINdYZRhYc7opr/G991HEJaV/2Mdw5jabQ2DmDBZMg
PcpLsw4cbpBZuL4A00QfWRvV7/qPbq83Tu/pq3rbgjBE0aUiNJOoUxrAvTA3hQ/z
RceWmiIUGfzNDJ29vbAfz+UiiprB5VpxBZqdXfiEwkJ3vEm+7HocMYVe0OOOzjJz
zu/U2pB2MRaEDVEVHm/iEqMLpGj0OQFcExCPQV0xJND6iBVCcn0d0xoMW9DtbJWB
dqHLjwF2k77PA5zDDHE0ZhEDYnCQPFV5++ucibbUu7b6pvMInCBpAFfdTs51/tqw
PLcF9bohnymr0zp3BkZnbZpey2/dffnGZFiShlECMG794cBqc/+fzXZH5e/hFu+N
SpFb4g08v5aE5W755IYi1CKK+MKQvIimo34/g1keXCewGG7HCKNYf9LvifjjLj37
fD9paQ4d0eA57zDMwv5inonYz41+V3rcOWH1bPmWCxzdR6ru3mxzzFMnXyLQCZAM
ilJxMy0ZXWRJXkvAtwjT8S1sFXwjk1VHZQ9g33JVA5QSuDXGGLkowWwCMqB5GvvJ
gqMhd7H/F6jzBMewwCWwLRamdVz3ygywKdXniL9WnE/+EKXx5bLrdkOdbyso2RgS
7jHbaxBpwnLY1a24llA2+ffMcBzbyOyMHbOQONJjfBcqT2NfPojpjTLh2VUYnJYd
o+St3iJIbh3TmAIen91y6zH+OZ2qFKdl1gE53s2fbinIElW3Lmpngrn0VgCHnQlG
EMKFOerkoc9+qyJngsmJuLbR3QAhRWGsiUPE4mQM5w5vfSIqRL+hIfMhm9Sp7ndW
8wmt+/94FNbyGbd5t2mjDgokDHEePUsuhwRxpN6HajMVB2hnw36ztndKOFfpSJN4
zLM7FxtBhjErPJxiUPX3MP1NcFakCfpxlvBWsWt46N5mR0kseYAw7T016XGRh9XE
odSUOd5S6ylOsRcou/FPg2QJlBHe+i2OHvpm/GOaIty45+znoPkeJF3gy0jl489l
vqu7kOPWSSw0n3TGT2jqFg/lGytimO7wpL8WtoHNaGB5suGAmKJjsR3l69aIHYCF
MMGtJACwIidolMvVVkfqoYu4YNalJjyXEKQCqIv80n9MKqoApe37F2CwsaoqnPnL
glTxz+oZbRtpDUxE/rDRO8BMCMmae01thbcr9p74sfAjuoLe9OoINCk7hO1sKUhR
933xBqCrTGUAQRicQC2J6abBycZVpZpzIxu/vOBMQ7Ds+/ABW6FfIe6OvvHV2N/W
s/26TShBn/z2AzB67nQGyQw64ISJ2XmOPoBkCXhICuwDvLJabTRUHdceeaETidzz
2QqTBCEzYJ+RIxtI37L0kLWaTd9BR8qCUhT/vu3nD6D7k9LO2wK4rNz7hQVHqX5x
EDv77UvcxKruw/wxKwDR3cy9m+LU36YZIwx4ICuIJkni+dAFkKJV864RPuoc2sta
6Ld4zWr4B2JrPQ9vVJ0MWH+IDlXUtHjcOQLjYT9lt/QzG1x6ncxSW//wp6vHUGVg
75aLzhO6QqZntjr8gzwu9ku76jvbMk6YWawKVqa/3LHCJyTKtgq5wwnIhblabxU5
fc5nOCEinEQUBmkblytiLvdpvAqfO2/jhN9Rhhj8fXMkTutdv7gjU6z76ySEQ9Vn
GRu8akJcnGTiuoZhR34uj4K9j0AZQ6JtV5UZgkLNArTxXwnrnPmN5tEUiTXGOwp4
tsN0K5Urwpx39eQ3d3FaZcxIv3GilNHYhPXogyVH+U1vkyPtZnqIxzB8EAYE3i+3
jp5rXQmJmHrRrhoKrlt06jH0PMj+TaWGuFLddeZOPLonTxf0uz8LDJY1q5v5KY/g
tV6J4JiCBYbx3CQqnRyrpCf1tgEZqv3UABB2KopS2He4Ung++YylHq+ZdjCSioyw
QH5dBsS3AXP/fcjXSD3cA/7tvBJWPRUbNDE+GYFZ8WzUk5jmyx56xkESUa0Gw1vY
BLnjjX43J2Dg46Tq0Rel+X8S3fzkbCdStwb7kKIJX2wRNIB7i3eDh8ooJ6h9GL3t
3aPrDMFkxhLTRVYCTblDs/xvrcHQN53p6AkLkcEJDBr0gMWIl99UJBJqMf6zdF3b
O1tv72Oqx9cEMCBpfMJodwslYHV8sXRJ8OlkY33cw98ClEaMPycUvJ0mL/1a29kW
agwYOS5r7MKl2eB0MO95fiZw3YH6/YAgfswHyocmMBQDZyTLAIAyglw7O4FFevoe
wPtWbxIJ287p1TNP4Cq+dM6kVB91ZWWmRLSV6qrt0ezPrNc0sqa19O1nJpCZP1UW
d3RSgflfjRsPs45PsQ3U2sYrAbGc7z7yYO9lNCxkmhyVDhdSvRJJT9kNGT7FT6wq
asUlxniX3+hetZhD5EQJ1Ysgov5F96YqSb1RrXUBzrf0XCPoGPYgdEDQdsim+zdD
GxjlWhpMNZs0Z3p+1BN2WVJFGEX43beonAW8tgjrKkaAG1GdYvz3z/CEVRQ6STH3
5tQSqq2kME83kItMxYXWJDtz+DNWAF467LfYKog4ztEEvoobdC1Y0k4IoIPrqKLO
9Y6bnWB1Z9I+raJFokBpN0fAwbw/RyzWBG+TrxZUeQ8YcbwmsVcOM+FK2KDJOXK4
veFlHfny0+wKWAz/+NmRGC2Gx4p1Zrjg8Vq7p9+hPs97Tk9UXF9ZAaGTQvfPy3/1
MSP1uTAgM9tV1c/gsAa1y1Wis9A2PrR5UNNc4eGXhZ7bVYOy4rc47QvZXWMNKbOs
Wdls4COE6xjBNzxjp8wawJ0tscd00wbApdRDjGJThR2fYCp8crrXelFtBmWHXknM
cWHYGez1mT92XUdrqBmZ7F5iZdJ1zNjDlYzKhS34V/NsA/bQfu0BxeFA2xGiE9Pi
b1Adv66e782JfuHkiShnaHc0UJ5B+wMZcSIguQgtyhM0gkB0Vq4iCTUqA5ysqSQe
UctckQokSpoq0lb2s50fK7Z53ic3qUtOKqR4VLmgfbkT7uyMLo5YGVktxPrLCfBu
TuZyeOrZ+f/QtxiZSMpL76sKHPTawB0/wCXJm4Y/l8GqG32uYKa+QitVytfTnbO1
xRLZs2Y2/op7/ChorjN9uTG+HYC8qBpKMS4gSbb7gFGkWvFOobVt6Q21+J+dwrra
sup71/w99UPCIjxFaJTA0wHshnFEBgxHH/EY29Wfhen02Lpt59sgCAYBjar7IuAa
ZCAU5LXuKf8nzgHbwFLduYguemwHmRtJg39EBfaBwC8vbsQCPpDn8sjccMAHCkyA
rfJIGeGcpmiOcrtm2l/cYYDhxVcrhyc7zHrCimF/dsE/tNHa8ylcVyl2ciyXbnYF
Spyq5i5efOF21hPesJyWOj+tEdBxmY7cNsL83vMV/nryP9Q/X6OWI5P7bINg7xLt
Ye6mz+k41b4k9i/ZWGhmD57zBG+uxw58aq06EkmeLZdDLdWhg6QdjJjOAGTy+/AT
rg5Zx4NRQcBPo5UKSjJiAYwkU4wRaxFpvi1v4f+cClhMA603+VZaliQvQn03AwTw
q5tB1irf9adcNaC7zpIR7cqRb3isS53/G+xoUSOJ8Wx2f2aVtcdfgxYaohMzP9Mk
8dax+iuNyJsXaaE26BZLtgJimEGFh5Fwp6m/8sqf4E7V+xCae0eyrnetkIUEUpK8
X0iLHGWsNaHJltFngyV/L2NJxnpHIlODTR4u/UACIjgXiWOTp21XzYSqzEKWNur2
pMyGT2616aLlIoAzKn8lByuT4OH7pFIO22zPSGfHm2uZmjNt8qop7THNf8dcf20m
AFklIEb2Geev/m5U2rswmiF2/D88DDs3DG4lwSzCc6K+38PnAV+ZHAbkEVvplZnw
UCDtR0Mcuz1AqRcMpWy7htaX2UUp5H0oFBFZflrgor5yqx26LJtPfRjh4RtClUgf
vYTWQCOvwC7QyoIOlC+FTYTXtV93tHeqwSRzl6lQL8/fXaZOI/2f9r8diOZ14Hx8
A9vIg6mAtPGPN1bTwxSMzxRD/Ffw+TCoecFFa0AtR/jxBqJ42panX2DFY8hLriL9
+7ej3mSbEVsfSWziAyZD80hCp9iOeg4+zTv6K5KQdLKcovQAFTzd5n+DTdHH3mSm
is8VFDVMGQS6OFDgZWUXuaW+rnP5Z6EuQ/wXfDwi8qzFIaZ/PC28zKytXAEOy8NS
RI9Zz6201tAv8i+Sl067m9DWP6P1RElxH6xEKIt8BMuXqXiTgIgibAB1GeVURLl8
Hcke7fE1mwvGz9BidIpRvit8f8CmIK8lVfVb4XGuPPmgRZ7WY4Jw+gVa1+41/K91
mW1IN3clgVibqFxfTMoXlNoIzWSHeQaTxuOz1dh4XoAYfpfZK76RAQoPFmd87Kdd
012fSqWAjwNUniEonC/FZG66k0yIR307PFDe4OIBpyNVZYWhn/kpowfre/KeOPuG
bLtD0Awefvsst5UZItmFR/Gtk7L/FughLIbop+gLX3TriPfsyUd0yUEXTnAo1DGx
ONAhJ1CXEITMJY0cUXoLje0LuwOy/InAOpduPpkH2HNP0Yg9aeEInzr1cyzCLLz/
xb4zLoYLBFn+7IUP5GBYtL653UHMg4BWJ/0IyPGEZw2YX/Dy/fgTthQB12N/BU/a
MHk4+pXYty1Q2DBQi6xRecco8jYnDTphykw0BzadgOmGt9QMXEf1oSVjYNw/sxWa
kkPhJr2St68kIksJ0eoZZY9HQ64ljrPUBc6HyBKn/FbnKb/5UqdNVtlUbh1u6Q1N
JjtNJ/0RuacdFXpMjW0oJzujMWV3vHMotPMWGxPVS1wBsH6y1FR145wLa0SIhhzW
w7Up4FLR76jl63QWileX+p+zuDj6SzaggDBVgMY7uuFZuz48RH02V/Vr5BpT5jrA
IpSSZFkrnTdANEve9oVCdapjr1clhQV+1BAU42aMEiOanmQlnqOSLm+ISzyPE8sL
yy55k68VlpeGmD8vEImaqipd3alEDOwhbIqbagYeCNviYpLUzt/8Ncvz6Kbpv4uM
jT0JNWU6oNmm/9dPcOn5tdYNHIxhTyQ3XgtmWn3RxwqberKZWw1fDBVa09Y4+Uy+
lYJIpbuoizoCo+l3ZF7xkU6cBGgraoFfhMyPi1OnKfWyzucrzRGa264CzXau/Vjj
ENbmAf8WAQx8bPWILhuKBNnLKyOp0Le0ccANh6yYkYb1l3uLYENxwjIiIdRMJOM3
M9H/qlg6r+kBcWyHKDg5IszqcbZ1BrfQUGRh+ZNHuZhutjR2CTIQaMo7YJLvrEpm
He+F0YPqKwLPCPKaxPVgaENGwgBlZkREP9MbNziUgoGu3luNRItnIM8+QLUkSZir
P9rTIU75RiwVjPQcU0DH84tfeVGRDdsh/GMGIWENlW2D+0BGplWrfyxnxRNa2OvV
9W8cFVktsO7TAE+mLkGACZxIO5/Uzh6NUBJZry2iE7hNPYe99Hv2LMh8+mZ8GSBQ
WH533TWsEaw5BA64IrOX3vGEdhEGLXlgEZYfKHPPiurDemsp90bb5u07+y5B4A3p
t8Qnz19atHciYaIbjThnq2fUdfOqxWjn2EaAftFgyoKUaD4JzAW9+wfkIYnaPnmi
th2L0/R3oe8uqeTjDyFNgufKuhkwOzAVwvGj2kgzY5u6FvkD7IAACX64muaTCiim
OZGSRHQzgGvlBnyVqAiJ5bc6CYV7nAhBrvmvDP9pqXG9ptRAB0iKPJh2+5nhh3J7
l8s3ZlRgTFg4tuARA1DREqup42UIp0Rkfgw5xSQ4vOKhhR1Objp/IBhXnd8x2Coi
+7r5D3Ob8oc+eg52MXw87xlDIg24z5kCKuarNf8uPCUq+AA+GZSgIFG+rWOEEynr
XpElmGzNL0gM3Yc6dfDdOy/dP+mPx+XyzUken0HgTtx5xfGfYvq67DVzjnKA4by+
fy+LrypjVv17J8qHtxM801YBIVMJahkrj6CBMRBMfXAKNeeTC/ni/mLHXJKEIpAL
byMVHhKk5bBN2ut54owW7u5NE8+EP67+1oGS+XQlsaTvyN43oB8dE+wnxW1lChl9
Ts8CpVLRK8/l2Uj46qpl8gQ/K+ytCXZnqpWs2JqnG1CD/4GEhS7sKbATGHc/A1S9
rwMltrMgzC7wR+Hs288RNQw7rY+7yDJ7zQYTrpWH13gte6XPSJuascWXiOFPfFEc
w50780D5yMSdd+lvXcvqTg9RhyCUAS52pIPT+RRuil+sciKr0Nc8PgPHMMJx28Eq
MVJdA7FsVxpmNbOVNp+5GTah4CCaUcbsTSRVNY+u5oBytUOfU1iz4zA7zdPKkvEY
cc4ez41WhhoFL4Vxd5x5ifD8FNRp6njwd2UmnZq/J+OOUhnWWtAvVM7KwRCzUqgN
BW//+i/gnjtKZcQg99XNQ1EmV+pbbDFujVZUuY4NtA5Hw6RzB9AQF6bJaa906C0R
JR3aUwz5iLi+OBPDK72aviVdktJ/08Wa+YQ5xSYiQk5q7yIyyk1piHOIh/xSBacG
EHobPQ9qy6HVlVcphQru357yJW1WcI+uCjvy4C0F+etKIVi/xmaQUHSI+MMQko60
gkdHIosH1LQfB/wCPHZoTMeidYyahMxUQnXTukIl9OnsRRj79rN0KSht15LiTCn3
3K8t9GYBgZ4xpDOKc9LQoa8X/tWozwWW+nCcfxnfCEkmqoq1qXbOPiRJTENUpLej
5pnbppK+hO0LQtZkAPmNkuAEgSnb2aHaPMs+ZwF76wAsdAhQTnRhJnuudAbuibiZ
fNIR2L9UCvpwXsJ6+ZZZBo59HmP9em/aO4e8HKUbnTRwSj9o3F1Y6/ZvSR7/5Fak
WPNFYBMW1NMWga/SJegztvtvOxCyxF4x8KYBkJ0QTuJKPM8lw4a2DLNR7Rq74wjD
dhb4ElWcD1j1vnHcW8LpRGUuWlVW0/ntQRmt7n66IqgrE1BK18tpba0tI/R8tcGU
dCwytmQAsL83ztAHzyMdHIzhGqhkbUq1XsDsyegyqGbwKe4Y05sF0HRgY4yDV63z
SYOr7x5noMttZ04JirOFCcAYlGSgZAMmi6J/KVEZeWTfWbad4E885QV4ytxKjtGd
vk9Ha7cyU88S+vXM8Bhjd8hf7hg+6Nu4NohD5QH9xtdtV52hfD0ryeFMeD/ZMlbD
2mmuocN+I3+Km0IYyXgCENqJSpFmLvjy7wWMovHUc4zuJEYHmr4/7O+qnwwimy6Z
1Euhd1/6wbBuAiPw7K2hLede2r+ezFgjhC/OglAMFXPvZ8cJ44U9Pw1Akuoh09cb
5R/KrrK/0kBcm1YX9tl9NJ5fUGVEwl3fY3VF8yrtaGxcMGMk1dbBxFlpRnnV5IQb
ZBjX9RUi5SOVk7Ej9ned0tq0UaDdl+xEOLOd/B+7hmPgtP2wC9+pyFTYIBX2h8q4
TmM3LV+BsDb3e2zzf/ubPSaP4nFWoAafeC02zoi7zK3GJBREhLu+RLH6ReNP8Wwg
dXozdvsPePSP2rERR/4yhm117zT0MRRRiU1z6ZoSnbwxh4xgDc8gsA/FekyBhtc3
Tf9MQ8f/Hyx+wcZ2/JFNqdwAXcnV5740q6Na97q02nBPHVZOFis/TRpymjXMJ1SF
aowENsIuoNu7tllZnNITTxW6z8ACO/P9WVO2zFkruzKGss/jNHF3ffeaP5TqqZ+9
Nms4ek3nYCLeM/X5kiu+TcEmg20Zy12+GAX89s7Q8eR56e7uJrJhqT5arH1hHy8T
fzeC0d95VVXs4RC8irFM121+JTYkKCQhF06c7hlzaOdPG6LbMjjXkSeZYVzIdOaI
svioT2M8u9XL4AmykbbHc22pJ7YwxhggP7WHGRpHfB04yJGqj61U1y7yl9mciqan
1wnWy3PzZcIE+ND+WUXPxVLzCzfpnS9iTySR3lqSn+tLGbI5P417/45419lHV3qs
2/fCSU07EtU0XqsR2cRcfRv6BQyVXLyvIbqvcX9l7bLwJesOB/uHrrWu9tZLcvxo
KE8g+fu78U42jTJAupDLCU7M4D3LmpDU8io/AdmVWNzzEm0E3JpQk5V93ql8+n9j
ibhk55y3cEoW0lTHD4wWMbG7J49TpBlkIXSn9jOziJ87ekShJc/MXZREMlyX9K7T
4hSZRxtjOc8ruXzKB8xVAVoUaU1V7TaQp1l6lwc7DvmERkix6boUBi7hm/Dkxgbf
soHVW0YKrluCgMa7FDvnfqwcFwUGoY4Sg+c3nVQlG+wCXujmVts/+P0lw6bsCoHZ
8HQXQfMCwCfvIUsdzXWB5rZC01Fo+TGA8KW5QPsYCAVH5Kis0/oL2NrSTgewUWk0
7QZ3/o4jUhxfC71CECICvUM/0Lxq5fevBB5ubPZ7FABFj1SDNZTWPZ+Sfz6eqJta
Nz+N+6B/qiTjj5dRz8OyLqQSQFYM16aMlINHHk5k2Pz+7j+Qf8jlVo85z+Ekz9N7
uSzrxnsPx3XTvhpkrj0Wvrq0wP07aqyaCIk9U5MynWIenzst2U8wOpR1YdLZT5ef
tM9go4NfpGNmqWk5ZYkzWBz0t+9ay8IPKK/KkBxAm5Vm3NrGl8a/M7jRJKB79ci0
UXizYcA58QvZrTuPltJmOoRsqwfdTIB7yO9NAOSeBPyZEyLhV5XTJkviQwWNDuep
4E8TYyBM5+A1xNJOQuJ7PejxEw7+s7+EgE4tLPmd6cEevhcNPTvPUhU1ue9iWffw
97CiW/9dxul+QE9zDQ07ugIIUvmkUgDAv5/vwhcY1mZUWbugIYOjww71fzv053kW
zhWLqv0ayL5SdcRK5vCIU9GyT9zqyzkY6Sd+blVpq2laIVfrJNdqzBzb1D8pkOme
ifBRPg1oN6W1FBw+IqG3kOL67i9YXmkW9cWxUApHjOdNv0KzPeWdHXYuTlfwuYp0
ZdBZpeES3O99GNR5xY2JNatLGYf2/3J47PTYP191pPCIx8BWZM+RiCtJGDnzSbdK
WagaCdCfO+Aym7V7ufI5R8l6ZhYAAD4d1QI69W2gREsN3DSc1YuPl3Pmz0itGD4M
cWYAUE8AZbWXi5W8ExyZy0+AT+KWfp/U1xAFC4TkXeaMskq/BhT+qZB+t0zYgxSW
2Gaj+CI+S5487B8lgExBzgu3+fxi0d4/Yna3AEfXpYXg6tG3JICJ1SAhj1ywjO1m
/tgz840sb1zb/pAt0gwBW1n7u4SlMsjK5Z1YNnfIyh+lMUtZLxJDoxpAFr0Gbhb3
RCe64l+tJ0jWDrnAQKttL+9ZB/aF5TG5liH1zXVoUJgsM077oOTkNWQidmhI7k9A
Rz5PLZMhJv2VmvDsNa4p1eaP0L/4b2j34Wc5S4yF1DL57Nv7E7ZZeZlHrg8wPDmY
1ocoEXecPAkdww9KjGjMQFQdfc9vIkBWhF/Y++Y4N/65T5D2aJ5tPp+vL5Zmqx0D
ViSpPMNP2J6dfJsBdfvi3mmJawpmX9zgwzMmMb9HZDu1MCFrxQ7S12KCaFAiUQWy
/2pt6cTE3Z5JccwRcj62k5ldpydrP03PZQODz0S4fEI7SDmfh2TXH1gBF0YMrSFC
w3+2K4TYD4lzRnUfH30U1fhtql7vKjHOzNMvv5DSvOdegYd3XcVoObaLvtQ2g+Bz
FsnhPcAmGd18Gzl4uzJ6zQ+Hw6zmvZ0tyqt45dxVjiO2e+mi60OgkxT8hpOYDKXO
P/NaN3LpfC4yx2OmTdv/9fbviL509jhjT29XLK6b5fMAl5QjI4YtbSeEbq5/8Ief
WdDntndG3r/BOAYL+4u88m/HRrvNgI2SYzfZQhRKw91ySHAilg92UlvIVHrzYPz4
O3DebS3zqRBNZxup4FM4t3xnG+2B5Qk6gON6cZquVmyvSU51wToPueg4QtyjiQEF
PnpzYhljD6+GKPDKJGzAS6SviJT3TFRKbWFUmLp4J0zQcabiHxPxZa/GQ1Spxgrs
MIRkt6ZXJPYeXWfnJOKcTlTV2N0UUUKwhOM0oJyUhME8mfYLI4CBtrHDnfRGbM/z
m2CkP+7iyqINQrduqjGgNPF1pmpq48bVYjq09rFP9daSn4X65lKciRVWX4erxqVV
Kd3cOi9Mxs8gGMeOlINnlzX4NcQ1/em3SdFVrziU9sdPTr7NyBcOAz56on55R87l
LS84P8pWYdJz1XxG6XkV1n80/IvlCJI3+KuxOI9Vj/+yyPhstFq8OPQefYE2FyU6
u3lSVISv5hgZ84WpUj4UATIeKBpS/V3JwSPU9ivDiefw8R0VyEGtd3R04FHae9uF
EQYZwOGvjeLLwqbrqKLdO5Gqbevosg/ft0d1QdAyDU8+6fsWjqBbbK8RdLgjEQwj
oJnjb6HMivf2MxRNF0KCfopdy3ZBR8u+5grcHsu90sUbtqTQyGwz2AqB5dPOptnH
RmPEon8QRHzHuI6FOM2TxLDMY5gg3CDX4Dt5bKM+lANEHfVjyhiOCPWJsKfL/n+0
mY3xAs5lQ2/sVAI+m/niw7pfdF0jOx/hd4X+NBgrcWWpvThZGNs827WfdGvipo6V
LeTn+0eDF2mPTOHvkvBeTN6C7T10QQN9K485teWiWgnH9jpk2p3uUK+GwvAwu54e
7OKE+KpRZ/vgC9NhYGZ+V1UCVxzniffS4Yzf+nSlqu2c+vyoFQjoPEjG6uhKsuxP
EEwXLxLNj4WWFBSMTDOn1LVUdunywbrwOtuimVYw+chpP7+NqG72foHViiyxrxO1
98cc3ErIkJiDMhhmDiNUueAEBPR7j/wWg7UQHVqvc/EdRdwrcW7zspn0hVdORwa0
GOnkxJGbvJCS/m0nag2vPhevuzu+wfliJLv88g7uhWzZcddI+HgLMCmPi0QXgPu9
gPoD2PqhTZOSsIj0ptLRsuUX0H6A7dfwBFQSQeBzMbAXKlEwH3ZsMxJKVSoe5GKf
z78XKF8vZXZovRbD8FWGz3diOWavk/l3BKR6DraeSDMJI01z1YdWCj+9mfLwpPyP
duPVAnXqyfeUtKMKdkvSjQPlXdTcpremVxkijteBI3wHzPq39K3yUYngnhJNCQXT
8F760m/zlLB26FEpUp6WxHG691rnKl5nffKfiAnTyuSIaGIv/i7B1VpxflGLmlC7
kAmXUa6/o5ikvPxdXa/t1aXg6v73RLCFO2c3UnshbayxnGO6FFfJpUale936QdjW
baClhrMN7KTSEtOZ2NpX4qOvuWBiQe189nxAlWTcRmFGQiwNDG5HkkExq4ayQs1m
xeqvNYnp/5AQ3oI/igHdZURjlil1ToYDGuaFjHL7eQyyjTyI4VDcFCQpNSgG/6YG
dc3lHZdb9j8ShT7n1sZKV2vd4kt94BSegLCywHy3LD2PuVyoT+JdCmqOlyiA0Gem
5TDD8rrRzWMnLkin+dpgCLAzVdl1aa0Z59XmvNFN2fsZ4TJiQygWPcawuXqOAPCH
x3GfKiqOIJUuEkAhWw3jBbbX2q3crurcEAZ7CO4kbACplx7/ybv1FUTOazkATwL1
EXg82RePibjWEzt8J1sIUps+7Mc2ArvBgCDs4apk6WRopHj67149NJcnPYbH2LNV
Mfo4WnAcyqChXTpDFOuki0h+lNX5KqtY1T4R+jFf3IM6JPcsV1eC2uljIQgh8onR
v5xAXHMBzVGY4jiR6qvvJ9NDu2BRVB+VA541M7AUGqhrR9rx5lLyCWOj/nw1kcE4
14hR7AwMcuginKymuI1FvqmyT9H2yBE4awn1mlqu2UY1KeXLdjBgmODxcLpAdaMZ
rx1QvR5BA2uRm6uiom5hxd7s4jS7TUyO1Yd8B7WNt9VCu8cFxowoKPRKBN2/l39u
roIJOzymfTW07dtgvQfTtev8ufbuKBjGhWCpthEQl4R9YINLlEegmDH9fGabaCCN
6LVL1rFgg2UY4nwN75uMK2eWO7raphOmcBX0GQVPBMXBcHZn7G6Oxii1XDSeJYyi
bCneqpYfE5wV5a+g8qeUmOPgwKJabIlZrIEnOA7pkGeWJCTLprOpxIPDTm+ceL8i
SNwCNcUpMXPJG4fxnP0+lMuwZE2OTUJZEDoybKIegMJeUWOUWal+SlB0XGqHkpOJ
wW0purSdl8OrhI+J6RUcrLDwtkxSK54ij2d8s4A1GyMxLsgaHg/4ue+wQY8sy9bQ
3d6AdWDDiL9Bx+aBSMhSrIU/kPC4obwLYwL7YNWeHhQ+aLiKD7O8Lu7+uBjHRdrY
RALIWEIoK2xl3n4ihcVISeu0Gxc9hsY9cV7lLvq6z3wrqTgY0MCRkIWMt+hKVM9i
RZ0+4s4QDtIrLS+PLK7FOSsokW+ok2sbkbg7YDiM+9HggPMfWt7Qdg8w8W0PU62/
3p6SQ8Yw12cmeUjYIhb+MqAaVFpWMAUkfADAy+IFLdz1xRWNiSWrPI6BsNFiAXZm
O0LAQ0XJoGfrDaUt2WTmAAx5EQv6W2h9KqUKktlzFnQ0Xz66VW+FekH8bgjcwFZq
W2CmimgAE10+HxfINbi9UqPiUIHeCjR/n4gjMYZWTv+lqJTy3I+CmaUXPbBJBId2
GAo97BGb1x4OZSbkfYT84QJPJpCJApdsG/NpTJtXGbBrW+CB2CWvIgQ81oVTM+by
UfxxnegybsdkCL/ufUdBCEk+NZclgOFFqNK7V3uqQ9VmCKjxi9P22N1lanwE6w46
ddk62PeOaQgai7s16jxSDcPliXLC2rhGC2SMic21eeig1JFOVNeEVHxF4ihsjGMY
1G7uCAoWIiEHu5bcdCffbmMY5BQHA2/l86j17b6oVVMAtTMmKpm3HyeQ58u6NfnL
wl5FIle2qAI8/+giBdUPP3p0sWDht6cSpobhkBGEGPL4wt5XNxjNiuZ/qtHPKM0y
e6rXqxJ74oPvUkAop+eBz/kcS2hCa2DxLO6BJjbFDLp3MD00RAbZTMoymhJ48TlO
eZe7VNbjetR1E/SWyLEtIrRwBfogNRcENaJuO0h4Uwqe+r8zM/PkrAUdv3PBVxqB
dRrSPC54odO7Sw+lHHKEDlKXpyr7i/gjNKXNNc10x2JMJlo1MExdSjLRl0JhRBur
qXPWDRNxlK8RojIvK0EfTI/uImgVZjw911qGedco9/huNcrgzMpMYg8G/3+Z50JI
7MYgAw9x8uA8xYgFJXVYl231pAnDgZM7KwaLOCs5zlNgVi0MOoLm2lJU1sJPo0ea
MAH79S3oupxr5ujgUPvLSUtwWZ9T+e17Z7V9ubw7O0EtX6i1aMIsmCZqHrbLA9XF
CKVeWcesID6wtRGLwQgA2P+Devws8a4ZdyRbTNwcA0teIjC7zdirv8fAljo+NnKF
V7r2jlC6TkISSjM99h5UdFDO7YGRoSdNly7PDsDB6i8bNZpHrIgflt8U5blh1zH8
8prLz5mDMXvPWkMckoR5umZ8WV9ESTi9yBHcsDVeKX+XZ5X74v4LrX1ZYglCNzL9
/CgZ445vVdWsAwFEC93oNH6h2iscpOp/i0u2LVkCZ/8SXbxRNmv0uceQlbNpSQJ2
uCkw0xpIr8SHLE7sE9guy0Vl3xF6Gmjbaz9M4lMgdfs7lrqPtWTNjEFJrAIcFp/x
xI+Yv/ZoM+AgySIpDYwMb7MBt+OU1U0jonNyNBlpH7/rjkpRAb5ve6a3iNwj/KeK
vegQ+um8ryQvXn62zw8wPT8tJvy5K/s8h5KSM5oi6ObT68Irhu5P7WYqWOdTHMKt
fFOr3orayItD7NLBwaard2hbmotkE7I3n2mb6R+UAOxLIM3su2rvfeqA4Z4RlEJS
Ek+tvNN2FIgLCO5tQAgk/LP4H500KkM4C2OkexIpBxxWzijCBNpPtKQepvNIVz0d
Lb4zMTyUmK6U5zsJ0y9cYHbqiELh1rGCyVO34XCYKHxmgg3cYUiQp4sB4jm/rU6Y
qLWWEAob8HLUXcQviHH55S2ioNjIpwZuNUVZLsoFKjJbqiYsQlFzns0uRapdYakw
mBnR00S9YToEBhJYX4GC/TB8k9y5jaqpPLiLqqYKa61qq0fvBwubcRh0T0PtRfBA
OgmsbKPFoiU+TuC8NchAIFOzxacY0lsbpz8xB4f4rIzhX4gpPukmmGQIv9xP63KM
WqjAOS9FVEXbZ0vyNoaQaTrfWRlE3jByq3hD0sf0a6YWDnRES2Ct7Ot39LNkUWiC
FnT215XP0Llq1MjtvUftZm3+39C6rcdI14KCZr/Pf3Mr1j1Tc+q+BlcJtM3NInnu
kZ/odaorZXPldhzPWCphRl6iJRPPQLzYmbhfw42jreKqq9Kd1kLJYqVZXsNjk3Wn
2xanjh6pGRgnRfSxqHApg4S9/Fzrydw+ODvFw0cJFUqHsJrY0J1HegeUyjkxuaYk
t3A4dH1NyuilYuPXLUlv2N883GFmekm0oT4NtnAtMUSdMNbiKjbJ1QWmo/vAbn8v
w7aEdQg9luVEfUnyRO6kiyflDAm7ZRPiaVzUy1v1qIo4Oo0MTU8kpw/gIQkmhSLK
mv0gC2CfBxCqcX087AK9kQ/94MuudCx/A1mjJlSgcT/Xb4FUquZRLAEmf8t1iXWz
dsFsxKjDJjooFfRxv0zCO88AdKsAP+CKGRyUhn1mBgri71wufZy8VkjR2svw5Vzw
YPNdtlfY1oP9cTgG2N6yARoGzF5Z3LwMzWgGN1u54V7SfvhwYRClVePazaUyJVyC
mU7Bz0R6yHycxXdh3a1qQcrZ1gNytBcw0y8TD8T527X2O+k/Ynr+1eMsMj8Ifucg
sRQ7szNNldS6iZAXR3GtKJA+LWdIS5vERFvitHe33KJ7l/z1wPhvXwbEtYGUgeI1
mCxCx1OsS6kA6VRnAnzreeaLvvM4ltTLLLdkqKrgTSPbVy2lUQZtLioKAnCz3BMT
AOBSb/ysRXCpBgbANgOtzbhlEUVE60yRmUtNrkz4x+nQ0EG+8iYOatHZP+opKufT
usS9efUht/wai5b2qjeXL2CChQ4JUZXlyg6d6jqJzYfhGRawwP/tuWL07HJTsUA1
h2ZSQ2OgLprazJreZWWCjh0pEAovWXVui4rZLEtXBrED+W7XA3Omz9AP0HGhildu
iM6Xz5OYShwuewbhiFCUeWnqYUiokJJQLpUd90hldwaE731CQe8Z9W2/0f7oEVsF
CDHDSlynMuuVjKl5SCquR24ux/w96LqsICkFfE0InstU3WnWZdHN834LzOIB8Tqk
PKIDtZ7NNVVy+P4hyJpsGPZcpTC0Yj8BgTe77CRct6xRCoEXlVRxU4v+J813bv20
S3rYILzEKWXw4PYXm5mJdIvohTDHCVcnq3U8HiCtJ3FDoEm7CQPLHYyf40S7TolC
nVBQJlecenuDWLpamEcbR0EEypxp2Q3Ug5ZO5LnD4zV8/TU8lFMutE6uAKydH2sj
0mgRxqyMWGCRT7bzDQInHJVgCkL++7aH+H1jAJ9rV8EPfA5q8N1cgPxM5KjcQ5SX
VHIWUr6wftStgOywWjq7nXsmII07auULY/WelKziplnliqhNreFRRPDNHoIELyVV
Nb2g5Qg4RLe6Zxr5aZuZLLD6ri9xrp/nzgUzlZJKYH3wYWqlc25RylNxguzHYVv/
i4Eo7atS4sJld/KQBJUKu0Cq5CjRwA9HH1TQjOqk7KJJtcTSWWJb+AZHgs/Xn35B
LY0Al+KTBvn5tavMh68WaCWgpSIKvu77YjZ36MBvULaUgMJ8o4kH1mxPwzHwS7WA
1spWcfcudJDyyh7OCNGGF1PiwtTsKj4a9ZBwe8n0vz2EtA7PHrJwNn8smoh8zPPZ
ynSkZjp5D6OKceMRP35Wy6o3wlggYi8rXgtsT6mueXtwjszzFdpxlxTAkhExAw/7
k5n+3ZWh4NTCjpQ5YuPjkPYRv/8XaQOepoyc5Fj7gbZEb36wEtVSivkAvWca3/of
wtUwzl7DL1nn4bqiX5yZN8Bvrq8FVcz045kJKIkDJo0XvEdqHWxEmGVCUDIM1JYR
MsDyaRZi+qhGW0pzKyNvKuyQNF6qcFe8rdBjzD5IzmHc5HwWGia0XUJhjgcKjvE9
xCK1LPe/oMVfZl/9Qcg60jQmKRR4PpoermhYW+8Ea2DHb7b3XjSVg1OPegZTTmQB
Kj1wB8HjHe8SxbS3ylAltt24WWx8xOXszFM8M9GWJIFF0DsmblpWCMv3KA+MUDC9
nvwsfiQ+bth6tiQV/ejrDHudmmp6IAB+tTsxKXeA/veT1ZlhqAn1jDnvq6/C/W8s
9OxcBGhf/cK7FdIYn4GjxQNFAm1bwgD86lo9f3DZxEbpDXeg/FD+BYsBG4bCIa+h
ZxQzjtaJQ9ITmH5o0T6c8PonbAxs4Lqt0hW+1aXZWarykI5E9mP5OrSPA9jfPM+e
UQU8GbYzNGQ6hh8lwA0Q0gktpeuEh3VxecI83D72aX8MabsRAj2zvMURydYKdSqu
N9kkHa2UuDvTBLdwklVRY9vHeXoMlWbO1lYCPC/JAU9itXdAy/1zXKJsYCYuk3pz
J0RH3NnWNwuj4NsPTHP7O9hsXrkN+dq1Njl4bDrPQk8WJkYKyocqGN/7QgVk+gJr
A1stTYfeQjnZ86vQeBNKp2OenSW5GidVOfEd9Hdg8y0WWejUFLEwYMobMjmiloB+
H+ZyD4+5ecpbpArJK35UppvGVlOndMHEhcQgEl2ewNVrI6knlD08Cu0UILgt9pkB
2E7U1PWIx0rV2XGPT6NMQiUG0T+Kw9XO9Zi23L2Ms9cuGtjQ+ErnS/o09LiaZPcT
VYwAwcNcyeqyWC7DFHlxoWfzDNpig+gpR/IkGTr0PxaaD0tm76dhoWKXL+yRRKZ6
3rrg6DV18qUHC+Mndw/amBfUhF+Ywi57YOSJK79tcHgh1sB/6IRkg6lidQ3hUDJx
EdOaZN04AwkCJc6mf51czPltFMC2DvV/EPeNx9Q/PqYvW/vm75kNDT8GRjVdG3sW
LNrkIFKNR1mnarfhlO37hu2WFls8G/W8BWmCZQGBSLGLPGLPu2VUUP8bPIBTdZOl
OTEemBxigMkPbBFIeOao2dyVeeXlDarTN7nmPmVX46x3IhDDPFu2HFAmQj+4RGtg
tvpM+tPCpq8ghW4S2v7XF8iXYysV1NudBuW+vyW1as49Z+7FH32FbDIJR2Fiiz0u
SQUlGuT40Q+tS6w9hHb1ztU2/nBVzgdCuCLZl9MxM3iKD4XRwfcHu1PqpS9u2tv8
56O2NURj8+TorTX0IS+ANrboJYaq2NRQwVl7LsCeqPGFBDKrtr8INIT3GwO5CtDm
V31dGeSjVOlOi+4zSWAf5Bu1EHcNWGD54/kUuxlrQZ3tLqq2tijPn0/6HXMk+jU/
UHliTd8IYzgLo7ot+dOEoyUjcrDfY+tKCUxfaMSdF30w2yn53f/Obq/0YkmQjzcs
Zvmucc/OJsdItktZlYAAVHluiOu5GYWBfzxKf+w5EXApYfaVPzyPr8kvmh6ady6o
fyEDXEAF8F/siYCBO5NO5UbrZHaFmiJtgE2tfUKONJye7nD2H46vYDxVqEq25iLT
vjQTo/cenxWesJaDfxmG1WXXcg79S6NTI839nX8639ClIpDqvhlW7PoMGYnpieg5
wQdHVEn3C8E8QQ1cROi5d/s1nQA0+ioAra5AWUZfRuhDvkpKhw2VdckwRgrcChc+
0ftGmB5W7HJB8E3v07dJoA3sp/fAVB2bCLWpbEvMQGQejnfQFEVG0WH4nf5Su4L4
6+M1bed+lGaKB3qSrHYrZ7Fh0hjXk3tsrqWqc1j8sUPIOXTwj6k7zvxbRl65h1Dj
sTxgpNTEkxf+n+EOtKOhCqN2jKv2FWmuVHIjtb2tr5FodQEfEKbIiISLvHzJvt77
UGWAHDJhdTcZpvk/PybBBzoDzFvcjop3B7j6FvoRuiCRcC6KHGM8+gLTtj7UjC/3
lNr520HFQYOaAlF+IBFxUSnJN5Vs/4z8sX0A0EZ7sYVPOCzZ23EOQOkSF3gk3yFT
bdeML7CU15DcHNKos2PhpI2sVbQvSKVitmLTp0MG/2yybJDcgb1tl6DLJPWJBDEL
SYlAbsx9yQ3IDsS1oY3hPQ/4iqOU3umWGjxdXacPHBZKTZ6D2ez0sFXzWcYiwDNv
igYh+PmKcmgQ57tw7XiMBMueb0VwlsCG+NEBz/K/MDo3wmP/mvcz6rOvOUkZdWgC
d54ZrtrW7bIWwrrljjGWTSrsgqE+ayzEHF10hhhnSQplkbEqiK1dZ0h0+pjGbJyg
cVr/6drTleiH85mIbLkZ0zMFEOnqPVXhUTUgvwgjiepuZaUZhpv1EpZhWXHFvUcO
IZFqu660Wfod4pF52UrHbwLCsH3r9/Sv1HYbS9kg4IDRGeEN9Xkqrz+haoO1tnls
xiEPvbHgqbmhnTdWNnDqq/ZTNN1gAptHLFJBO1H+wQvEHzIeRXf/frfUmoD0bcfE
Sjr6PwVMRvA1qwGVsiqOR8H6PxWIT4gJhBHuRGHqys+gxRClvOGb2fBNoqJtItsY
L035GyWPekOMRy2oYQrIj2D+xD0jbLU4PgzaNOQztqhkn98W3/NTiDAEmncY40Ou
nj2aizTXsJm0qO4yh7Zga3AsRjOUILj96M4ntPQO+wPEK5h02T6AgHB0HsdZwU1o
F7XjVp7EN4d9n0wslzQVwr2SzJddZ8d9TrNmHXgNTjlFX1Nd6ZEv3o6sk9EgP8M8
5hHjenuQh/A0eAUh5LQ3540L0W4XnjzDbEP6XFdRGcSs3T1XpkX2foyp27Y5onj8
Ry/+m6XarabN+uuoKk21YszqG9CIXpLp4DghG+zvqI61Lo++6Kw3loGGjeF5e9xG
bLCUjzfD0e7fUtnneyGd948R8qW4E5rdrIIGYw5e1QYdiLszNzRD3oJartHhHOXX
okgQQxwhgoxTc/Qx2GuuTCdiN5VIpQt6iU5bkEIrvJXQBNwUfJsQwTKO+Fd0676Y
HfACSsb2yrr7qSd0EbdWHO5CTFIF8GJfFIonGEkVHfZxBvpkmQYBdrdHSSu3SAIJ
lkSo0ByvR+IagsTgNdUzn2g+z0/uAaBuekHWZ06Y8+sfcck58vy+rBGybwetb+HP
W5p1z6AU1zeULI8vZFk1xtpRaf3cgewSEHA5HovNyBDqWBYHbPC6S7td4JkJh+UX
gmTz+R5EFMhymLbClxJCHqw7HCCS83320tHUw58+l3MXsaFt7kKosG5XMvbGyEaB
Mn8hcQEAT4MWD8x6XNARBF2jQEhi4lBmek48cDHwqySGqEYNCamtBhEE8jOJQw0n
3UPrtKBadRAFk+PJC/WskJADjav6GhmAzi1K8XGoMl6lvaK3tZQTXY7YgwQSAYhP
XS5Tiw5hjq17FPLtljvO11TENgiInHEz3JDpq4v8tTH5jy7aBkgRWFChJWANL/zx
ZXV8PtzS+6x/0X55rmbHsjpV6RUEiFMWiV92tfB+QHb62MHn3gp4ZsNQb/P11bPa
ESVPjFwIuReY2zOZfL3anZnsv7pabLbWpSL1gE5cm4suXDZgD4iGuZRg3JoGOD6T
Y9uTVHbqjjakbPD3+gO3WUhqm6A3SI/O9KtFA6U8ZpmUukEE+QXrmpKnZogl6qJ6
1OlKDcP3kEc0vtxsmjQOk3VLgHNMVGbbAOoyVbf3n3Fb9YtGZbxc0cU8iAObdyfT
jbb6MnCSUXM2we7Hg1y6BcOie3C2THCqYHJpCJmuHBVPDiGzgSZUNzif3iE2KMe3
rRZBy7k8NRWCyiyeiw3A2P4L8GaZQxbxsBaPIeNGLONmY2h7tengVsQV8q8E9B6I
qpzdjZwfxracoOkEEXg4MbL1oW93YLZOhr2Uam0jruy/5tP3+Ev9qoQmdLGKV7si
HnXeqNjvEp2BQ+vPNnbyi9qARnn0SMtFHlfgQplqWVGN7oBoSpuX2o4DmYdKIozS
uEaxeEd2Ajk4Gsxu0/s1bWytChYZ39Fwwh4smlwfso8msmvSjm2uaYDZAC7lYjSk
JAn4zZ9O1uzzWlaQu6vDOi+0iF1D5SY9HHcZkV+cvrLLtn/J+Zh9lOOL+XI2+8Pr
5Q7wfb4zmRFvxkowjgtc+bOMor1UW6mWgpF0Fx8C1uqk8EnouUUq8X298pYn1Tzr
Y+BUAbPCjWVY41zQh1HWPwhjwhMW6zmUQ5cvoiWfDItv8PyLoeRMlYPHwraQjcjJ
kavKu+Y+Suz+63Oh5qc2gXv6V4NAli5hRrwYLRSqvY4Qdv1RyY7f+ywk7qfC5kE1
vL7rSyqYGjqcZoC85igL5GIhQXGTk1COGftVzaMfKdl+Z4X/0nb121ElNgYZI70r
+TlK5yyQeSt/Z8BUHuxkB/r7mj3Bp6JydiEjVSihdV5YyyGIJHwOPHZDQfVi9fb4
FtqyDnWgTsAGYKdojy9/lS3sjPaA/UMDTde+kyQQ3nKj3iBUxYXR65VzUjOUG+0c
aPdvgY2/YJBVIP6pUJ46nQ2+4xoWKqOy+A5jzKTDn0CVCEd5XjqHM5Qvv/MSbh0G
z8nDDzcb2UzQpTyyAcMNzjyI9CV0IEUA7ad6LxxrRsr7gi7EBOOU58IGsKRnZw0U
GHLaLWPAHSdANPqyir0BYvhkTPIMqxd3T/5xkkHoLy4vqaYzwbyS1JoZXaKsp2Rw
OR46wj2W5OqA9AVvJsLfjhb3tTviQRsQy3LuUEvqSJU5Ga6MelPOI50rkTdefMaP
BWHEnxWwKWdE/IJUaMpFTGPQWrhB008xY7U+iuB9JyLeR7dWiKaTTgGwQelzS32s
VpWdmhBYsyGPwE4doT89+E25HvXT9Ttgr1Hm3xFPtrU/9MqKlDcqeS3emfxAxAPy
nnsY69c0cMA3GiAuHp2ucpf9ZFtO3HvEs8JUfCbQja/P8S6lT+SPkN1usy9Kyht9
x8b0/QEyXTuuXKJqLFWwUbwClIxVIt2cAsG1zaIIf0dKrdCT9eYNLc0dlBNJT1nw
VZdixRjGtSWU8QvvJTtyphWHEe9iH72pTHJLai3zpn7RrGb1Rhq0CKvv3AquPBD+
4IyuY0qB4/fJCtf6HO+0dgUGqUiqZge0TpXG1SXJl2UNTschPIsYxrkaEhSLdDlJ
XYlO6pt15KiQpbRrwKkADf6KOO+d8Xr+BwTOpjV9qm7w575XBT1zr36AbqBpr22v
reO7m/rapLB02+mtLX/AnwZQugtG9KwSJymGbbw29vA6aIsKjvR2kUATREk/nfeN
ZCT8DyatVE1JTdGaQjq5FEI8m43QmBL0iyGDbkwEau1NngizzY4w8elED1JgQ3yi
ENIGCI7iWZHPoOM+Y2BjrpjSN2ZbYHoU5vg5frDlZWUzsz4KEAi8XmmDrxmzpM66
XpHYSIyGEr2aBpihRT9Bh5d6hzwEkn21Aax54AH3eX9dfIYbSiaWHlpgq5S6NGem
UlxBu19Du2a+36GgIRDhh17N6GP8UxaacjjEyU1ct5wD7xEauxkhEbtbAZFetbZ5
xEpHASYVZ3D1svqyPvh2yKU9LQPJ+QmCQEQzB8BLMbk0q/R51cpXgr1YIaVUEXvP
NRedsjYhznlE6lhdqcfgSMuCFaR3xCxcx2C0ea6PXZ642x1A+4Xkp3JvxhJ3Fw2W
ye/W6i+Yl3lDvXsqWgFZCGULELtN69B0hyyVd4Ns5XIvEMg6H42gNZ1mtOveggGT
2UK2l9vnxZTKeyKGJtjbiqPuhhxugRBxW4u/1Vk9I8dfDNv85NmuTdgT4KN2LYMW
yCE8x6zX3GWq889cG0FAbDykjlz85LCv01xzdsn+bJQ5llNM/xqWlThrsF3ziDMk
yZk9IsFINS0uc1yjmLnq/McCjrc/gPyhNIJZ7e9tfQce4tCpvN4sZ/FKdLVURHTn
75CrSGK1h4hCGbzQ0PYloq/g4xERkwQ5orudzPdt4fnJWFAExbcw9QKmwqccjR87
mlGH4kZLJLU+axx5f1ErjfSBUOtsAekkTTOEeyZ8PGhhd1X0JfJC9sTztPoWQZjP
Ri3mDtLYeLC3v8CZ3cvfzAnr/UIrI7DYfaRl3Anju22stOhbWOwphngd7g2PhvmH
ax9MuGLZNdyOuil35e8pR6TtB+vb2TtHQ9LQ4epKWNAELvZqV9DTVRd0gHY/oRWi
COxyEXwGxtiprW7+RKOXQ+FoRNEXR2GBv5PVqu0KsgVdWw4zV1lhxlxc+b3TQr+o
gANiHiU2wZpGgntiuMi33EJYcwSzIXME/158zLAh/qfkeoqqwLs9cx4Xymusd3aU
5qqRRp6qjTfdgLGRLPXZKhTKkF2SEwrXwXJLA5xl05WRE3XXEN/9+FusXMcHkBk7
1fwAbGUiKMJNi0GhYECLNUmvyzDY1ThK6eZ7HqX2EmsDp/u9iu3iveVVCcbUlok1
ikbxiPhD8LeUrj7gOMTl4W/iBfNRcuZJ9OegSlu9Z1YbAchHJ7ZT/vajBUEpCiNG
1A5IXTyJ1wFWcRCZ5o/2oeeZDzizmp+cy8uQspxgcU5WlWusJe1ieAja2UCCT/Pu
QEkIiaCvABN6A3AL/RaSF3ijjykQ9B90ZT06xUZOU6z8kRq+4d40ExY7iRr7wxyF
WamVSRGK+KMCR2YIeO6XGpn1CWB3nw/0zgxTs7u2Th1w8gFw7rXMuvt19Cm4jsHj
EvPgswb0P6GZlqvmYTVStM3Y98g8VLKllO8Nfpk1V2VEL3lY29gi8Mk16gP/KaTj
9Tp//sxI1GapA9Ug8MFimK1Vqb5vKfp6AqYHCIfI2c05M4CDND3Yujr94W9oGKM7
xd0hf0XlwQwzOVfdNcryJ9/jmQ3+O3+Szl2mnvEmyr+K4rnATErABoCRvwN3QP8n
wBuS7K75uaaPbRDC1NzyXxPUruACjo58LnsXEbUNAw3kT3krW9EIjO20GTjvbgDs
XYPCHXhaVcZl/0TwYIPPUoShkGgMGL7ha7M+DQ0LdBU608tz4gR9x54iccTqfPx5
8auGVGp9FDBcWxAx8GTzqCHWrdBhSo/U3SJp2uttpudaOPj/turjEAt04su6drcR
0uqkS8WSY1pOisURAjSxYeKPrcFIqD8uRfW2o1p4z2SWgonTfnYPrJ7rbNr9kIzI
xCJQWeVO3pmovp3FCfwxmkTihATffy7wH32I3F5zO7n211xF1UE31+I5J7XJnZtA
absY9NP4FmSpJZdBw++5abALoBmrDyPnalax11di9JiBgCfANGx5uvTXg3f+P86/
DTXIhoeGybFhgiix+vZvIS+CNg3yTvqSk4hHoUtpgazVzvUCAahOH37Bmm8zaGRa
gHmyAqlMvyOiWP6NJqWtt5PgeDAjj6MTxnOT8qxNpXjpOXqIzwsKbViQfFJ053Cu
VlElYA5IHoe8vhg4QxofCudP36jE0hRsV0b6vhcK/wC/xLqEl3pVbwHa1YAdbx6r
auHvlsCxRAP703q5hRJyAKwMixurkyAF7wkRqe11XXzwArAYMntJ5q1jlvLLrPaJ
AmnRkSlfxVc7Fx6DgtVVNm6UZ9z7DoYAVF/+aojTN6/UyfSjYoKO/brLG2MRsINR
ETPx98292Azv7H8XgAYVUs8RXj9IRr+DD9G6msohzYmvcSo8a9ZSbuhnGVABP5Pd
zTu/DLBQc0j0+vL8FY6nktqcnwwD6ymwDHx5WI/UB00gadh3KRUDOnXUpSK2dxFD
6ezBjOBNqmMAA/eZtwsFEwbdCK5sKmSAx0YkvAh7SzF5MG6oNq5onlx8Gc1zaN5p
MkP2sck+JIwU8bRLF63MIMUKkZmbMlP8WcgNnJ5k+dhtJlHloThJWGmrxGZ+QO9V
L+U2ErJkrQfRwaEmLMERpid4/U40ADJgKLNL8TVKOG3Gsr0Pg2SFBL/qvGGHqrLm
`protect END_PROTECTED
