`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GAZgyVP1SDLV6beX/H+FnTWeeubM0EqbEdWRRV5KSMsr87kg4todzh1WPcRe+ZxP
caiEdIUpa+Fa/qKqcsTe7T5tywGXM1MW79Yy/VvnDOXxYQgbJV0iA3KJSPrvrYut
GwfghMacZIFq0Y+Me8g2ovI6HEmp+c3i/2KHGhmevUDMvmuAxBweLZpYk7atzSOy
EbWLuXRMKNn2jIfRsHXyAAG5+AhUEld4tUQgts/kol/pY67kmRlxTmg2lhzyDF2T
tXicxC2IOcbpIAmaRNZKDBhKCJInjSsZesNhwF33xY/y3BfPjVrhpsieIaogsUIK
Oo2Ao7WzCrqcnYmObG+7QBTeyu+4JmvzCwq3VwdAcy8MasA/lHqofUzckvQOXFWW
Na64UaOH/Wk8epIXLhp23flqHJbWRe2gDD2ZGQWhE2FTAK9FOZFB8boSuUBYdWGv
VtFa+smuQWvhr+x7fYbkFZF1Q+cnw13oTMrlq2fgmJiiyLUjnfzd7KEml/k16eaj
zpTLmbMJ/Hf/LGu3xHF6wdjH9mDkyfjfwwHZIoJSj/rI86cH9X4UfGj2Ba2N0GfN
MRelU0JQdURzIS1/G18lt/xfJlJHCv1lNdsOw/kKfByD6cbr4fJC2XwGWZAqbfVA
P86G55icE5r2K4+n4L7PUfQrWprGM2YjfxQln5Q6yZikM1LVloypAtW8f0AyCZBQ
uCInVCXHrZXP/KNKf988nm3efEuqdGahNcCUeIinH90G7cAVeTI1vECdGH6ILuf1
/TOMbteqiu81T6zd98CueGVsjsol/Qk1GpZsMC7XEiQzhhC7RC4hKh9WbV7Y7yXh
HsJ9fquh67MqahbcDEILlf2tO8c1yeA6MU0B51gOhZ1zvj0URIB/2pLjELSOV+OK
wBdv2KBABb53xWCDSzo822KDdZN5JE6irDue00eTAxd8xkeKK2Hzx/2VHuc9LIle
6h/uOXawYgVcGbxdqVVmhWV0E2O0752LYs8w65aEqDY5AVewF+cwHhgVtJqpw3Nm
vrhSxnHqqeLtmZD5jh+Q1PbuDwPErmNFsn/if3DwLGE+y5B0WkBocDHs/B+uD0Yo
ScmX8U3USvuooWjJeELuFf0dVmddNwZhzq2BSxjYMHuImbZJMSJqAA1G395ffeGB
5pzs7izzt4CkGLk4l8yirXefw1J/RJTrHekD7wRhdonGdt2pP1bAVnBkNbWkZEUs
+6EOZXhk4NowpJPv8skwZpfbxtc+4tZCAKYobUU//Qb0tS8jde9+q8i2e/1bG3vh
gCqyVgQMIFyEJgwohY7QrHKrW3m9S/uMIFV8LYK53O3cFjcwkVIH3lBI6d0LhjE+
5uS+/KJ8OHJtaRbFAbOvsMlXzQHB0MLU9Qr1NSYMe9wYyHjtgXWqVmA6VL03UN4V
AMnS4kcEK46UbdblB4qesj/d8ZqT0uW5wN2odQ68Md74RdE9lTuEho9/oyfXweTJ
`protect END_PROTECTED
