`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmJAxpScAsvmjHa5unT82ZYsE6SOhnxoCuVJocFBNywFkeeyMvdZ3/7NTuGYEfFw
qgUerStmmXO/9Qsmdis6xn5OAbmYU0NzgclTq97Ibm6DYVYH5HxOz2XVG5uIm3rl
3jNKhEJUGSUOzxoGxe1N6nIu1K9yXr2L+vwAnvYrcnMeG/qigkK4KvzdHP3nCv4Y
brifZRF8Oc+jT7jHfc+6rtipK3FISJHAVHHJKN+dpwXr3hwmQ8WUf1mEqaZEG3vB
RtjHhi/T0JJHX8IIzqSDhSp/8mOQ1dBVARFwCKit7yFN64FbGGjRGJwf52FOQyzY
5ptUSe0b1AWhk83OIfpeZzr4IAxbN4C4WY5sAkTFg4mRgmG9EI+KZART37IHTnrk
1tVnVINIC7wDlh5xKmx29kubt74R/oA8c4A9THg6RZIBAv2PDQMqAt9KVTzNCWOx
yxtjxFrOq+mG6SXp15V0JlfCjE6WtwlfuM7OwKz+1GYjXULG5h6qO31OwZnOnI58
n+A+i7a6dT/papgbX1OVntRjICrA8dF+qScO/uyJMk1jPdaBfUtczDf343p12LyO
AVVfVnZ+OtjdhmWQtsmAwLH78ZAZNBc7FZS1k0Tv09ZC3zYHm4iRdV+EqDNXqREV
fdeRvECrkBh5Ks3C/bmb4Zq8lFTFN0U9byvYDQrKWsJ2dfXlnRkiGHlWkySmew/1
DqL8GQMRMb+imdW2YJ4aB6DOzpNjioz91l3Wt6URcSxKmxQGoOFZ91YRjaMc67KB
aan04ng5SEQOlBOe3RUX6PntOnqV4BphO5kQyd/3iVKw7ohsRXQiqDx7R2L4IvYh
V0sLXxjtoHpcSQoR39Ea3L3edWjJIVUXCgF19HJOJvbH7Qs91DDjFspn20Xw/J04
9+jCUCeVlcjOPDx9jcmvijsaxhbLD6imhumaVQnPfnkyA7DYWw76zY2s5/pgPRzH
c6643Dbdws/78LdiQSi2tqt9REJhVyhYXkGwBAJqmwn23VIH3OZrVOVCGqa9ZzCs
p5V54F7hiKL07yMasWwsvNzBDgI97S9ZdFIQ1gd30mJoceq7k7cd4CoIXbfywFJI
IfEi8zsiXKgjjYgw5jtbjyecObx3VkWxvKzrSdQZ+vzRxmREXrUEl/Ro86nC82U2
GI/QMaBpMvS1cJGSYSowdlUrXMR0tczENXV6TU3gzcRoHS5Rn+2MObLnXYS42E7G
D2/kVCsR2idHR6NWWjSnkaKdcMIBE1aAX5VskhzmCh+j215kYcApClpBfLNFK2pe
TBNklqREV5EJ+efK7pK0942fPSnVXbPHKu8KUas+iEr1VMAtHuVQ79Q4MArrbI9w
qX12RNedxXJFnOj3VlUXB6i1RadHgoHD2kx6YHeErvHA1mNJSA75JXVMMuCtCBVT
zLsTbgraybv+yls8Lli5JHNkIT/SPtC2joW9oxXJ8saOUdQp6UXgt7LYSvyvcSo9
Xl/8UmY209oR3QuShs1EBpUxwczD4UVMaoQ1T/B+a7r1nhYkakMLRyYD5xcvmn1R
Obl95FZ6KGx956bUo040FsHgmdJkE0WFvsg4PbrwJH3JOgHQN2PXKywii5Dphn68
C5lHeNcalkonfjhSWZutpNGaiw8BlzJMH108zN8LmRN8uQssMtr+RtN0UmWZ/Cdp
11DCcSS+20yQIZIKv4zPbgSPc436ARb/oZDqg/8C7N/aAye5XtLN6Hiw9g5UQnVN
KXEWPckVUzFRPlYrS3YS/CSThIMN9i6WFxaJwXWwKyz96AhTlTG4ziMt7/NGSC64
zoz+AGIrf8RnlSSeBoYo7eCZkkRfoPz2owaI6Tb2IrvGhLq/15mxpNyJWTJt3NvR
tYL3E2ui7YG1Oic1zuDtVi15NRm0Zc05eVqzc3HcTrhVxjEudJxfRMhwX5rWwy+R
HQER4EjC8NAOfMyTcmPj6wcpg8VC9GU6TO/qBtCEYcvdv8y2pWFdE6IUc2rHRPkI
dAS9YYRjLEDMDLa1ND8sRyiYgvftC3DzfxWS8xDdyV6VL3hqp06s1djlD4uofnGB
RPkE+j30brmnnfvfAQ/os98MVq1crRY68drM4UgCNej+8eoL42n3d5Oy/Bq/kImO
NxhMNl+Exj7zhGN091JP5S0OdFg1SkhyAKH11NePDWk2PkdSW71dk0Q3nndWZXda
lhccYemp6RVL/nh/JJjBDq7C3MG8+YdgpdLzpqA6R0opQpIEzJeh4ynJ23wovwuL
A3KJK5650AIIJ88HETyqeI+OCGQtCaVdSmAeNCZ4kD6DPBDU5YVuP3qbAO6ozNmy
kWMCdrqd13TNJF/Q9TPx39uN079hbS50ETcCKi69ZFUik3ZADhJ1M6FcD4mwcvuy
z9bOjW6Zyfqax/mg5xXTUGaf78X5TSZUSAkAIP0hoKKm2bu6fJ18FRtBNFWzIJwe
`protect END_PROTECTED
