`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7dmPqPqiWENDY42/w7QjcRGRPGpgOWSIzrePDZznUgTxOI1MvXVisisc97T95eOX
Qot4Kad10Hf5K6gmMiLLsoLgbsJAchs2wKsOqmaXphj7KevjLBPYi0ACOQC6ImHx
0yv9uTGUE8MALD5QOR2c8kCakQM6YWDfihIDrswz8cBV9JObwuOa4sxS0TALMknz
UdRDOt1z1G12CavU6c3N+WgCA9371NrQgrH7Y8gKnhRO9Mq6jaJNIv/D0qTADI7k
9qbD/MPUYZXED2bEAcEufjePEzU5pjhHNXNS7LZVedd0QARrpEA1f11+pLmExVPp
4+aFew4H4rnSPaQX2Te9D21ze3n4FiCtgi/NJMvrdnj/xEqZxDxQO31w+lZAAMs8
deFfkSXJcayXQhoXBA/IZVtrII/E7Co1+m0xpzzw1i5c67A4LYIl+ARG7CFE48jU
T+TPhHErAISFXVuKHPO8UzQHsJKW9vNclL04ukwVLFxVNvU1I7c+RvE4GLuAGBq9
+uS0Af/h41ndeKgxHHMj7ouqWeC73K71+MI7K/wraNjOIri0LwK1EVEpLS2R7G1L
eLnabJx+IV6N97pvrHVXaO9IGCB+Y5ASIRxoQL9iyKPMlslHTYmHwO0yZ7kpP7bt
LLxilRnxQuJO/gYG4JJEFIO1UEnTHIpsA/rTCiwy5aepJUnaDrPlrdEhvuJTeysC
UPpSDdOGDD+y/QOGYDswzOE4WNvQ33+Q7P5eGj6ppe6ZhO0ZBggXI0t6+7qcBlvw
UYIpX0p1TQ6zyKNeq2WXVaLTQKXW4ir03Sb3vL2YJzkqYkd0xwRENl5L5/OoePpz
S+og80FuFlm7PrYJpjrx72ZvjpT8WG4CoXHuD+TlxiVbCdcrPYUzdwPdDOSJp5BX
aL4VgnGKUXB69KSoHsy/EZFamBqWeIpQVuhOGm74uhxjuJ20eWjcD3ho65uEZJ6i
TeUw35c94YuawAyS4Cvm2tal5b7Q3aY5C8xCoU+IUfJQQ+FHVpqdILaUMTF+P6zd
grrUP7c8HQdSnAz50bnKT7mN1PuW/rm4ZZblTeHsq7Nf4zZO1Ta99H4kreLQc596
8KgTCNmg3sx5PqBIQRRUy7J6ThU2zoFMFmXRaLisg5CuHy5e8l6MOBspjPU/3aFO
TnsU4B/+PsxNnWzuK5lnuY1PIGA8f/6ss5oe3uO66m9PTdrdJ11/GbH1V13ERHRf
RSEnZi/Yr5qnb22srMHbXVsGT0X370vCoHJtJNUwB0A5iTvZ9OMGmglgNYfGvzlV
aTfL5GlubAa8g2/WrMqfQ7qpka/wueDuFqtp3gC0TV591lb5H2rRNCRGKOT/QCG/
3X/Dlz8keddhixgoD6QIRXUE7npNxk/E9DNuCxTw+vLRg9BOdXF735Aa3qxkvJkd
6ERVqVYcxlwu3Xkur5OOAMf01e3k6X+CeamU2U63tJmsdI2XJr1JjZVr/salDXXc
z3g3iUolAbU9Ls3P8TY/++zM9FxFZm5EviI6V85XIcEXNEXQS0+qQm8pVM/M/eT1
M0jc+ERoGHWMk+l9suLNlh6wykBx8zsUg/S9MrlGoqA4GuUKnkab8W1KkpyfvnfD
LIrsMjL/Do99T5u/j/zv+GnYLEsXtg+sCruKt9BzoDYPy8V0jJEOAnCa7Y3cUeQL
YKpFDnYCHZ7uBKi7HjYkIXfZqTUJyUoYbNuYdenUECletMYRFAA5kgBs/i5BvEqE
hJXETeb8+xn2vnXGte6KqnI2dC4Zo2FFLnCNpJWE8hmE/qU4WfHaMoZEXmnrzfwN
Fgv3aiGR/T7Ur+z3NUowRQW3rGb7MnIgnvzTqdpmYaIaCh0uiEx01Wb90DsmYGjx
QR1TymTgD4IoVqEpSQ1ojfSGWXommfbwETuTbvy370KeJAeZ8KRcxdIx2vwucyMC
x1CWDBMwNdoy1UiU05/duhKiP1GsaK9bMrviqf1ZyhrdlI4ieNOh3AfERxVhGlin
4O4JAQQb1aoc9XSTXvh8hgtNuBCkpgK1ze1l0q7mnPswm1i/132cC3ObuQhKkual
ehRWcaFKR4O5mu6YgI6NmcroXNGJfS9UoA62j8wPQDh0HwIblcs3gRj9ZUEgtS7F
6mpZycsapK+lc6J0QmmL5WVfJMA/FGGaDY097xk/iVz0rB+Mc5UcOkpVkXOXv4ge
DeKbATRTZ/G0qBPwylndspOinmbNjGukexH+IX90gL+hHYkdG4T7QYSmM9m6XCtD
BkW+RqOmI9PMuj0VZXpzLMmAElQh5OXue0Rul0C/HnZg6DIZzNxSzR3EVJi2vNQj
3PQSyqyUZie8kOYiVbQLNEMhfiD/Oi+Cb/34yfI0SdLfJenpxw7BELidsy6dK8aE
E3w/S36OkWZsLemEkxFtMfhJPvmpey4qiNlqN2ZoucA0gQMQq9nOEljBCEMyLVwz
xE6Uk2rolbIQSfdzrbBw9+Ekw+Y1ZMJuEAhudjXKARob3HCr0VKsVvFJ4qCi12rL
OtG3YCtFgcS/fhOx9C/pPK+V1Zf6W/7AT+czviLzRrFYHY6ljftumu/SpePzr5XA
wMcgAYEdke/I8hpFx97XPp1dX5fdTISm9a9rwkg+yo4Y6NNYE7euWmosr6o1Qi1I
0GtUCh15WOGgmL6qVXFkE473DKVU7PhDD4F0wSqnKlzJGQwmVRDM8lk2COnIvp+o
fyK+O6EOQSGCN1EtquolZ7RzmniklThftW08PNKzBWLN7nx/QTuIp1gQ+z1W8+Un
PkrkrvRZ9iJcq/3ksZtmtH+rh/rsonoxe2GSqJFsnSO7UiCVU0SdyNoMLUT0Oa3K
IITs5x6RlpPzRH/YcQZB7vmsL/mqy2HvcqZCqJxYzdudIzAlW6KWlYYSnjU+Zy9+
Jk/tS15F+ef/uFfKIF8SLk4PQ+vf8bSnxfBKssgJQPn3hi+mrSSWqGf7EHWHKzgu
J8SuL9aOD37gphJlaC6f/Yrfzdhd7yQkYaMwd2n5crpYBj5ZxLmfFZBaG9sssD36
PeKo3L/m07iXGgxngPcLoGtIfWcawQaNJyl/pRcaBY0qCsfAUpq3UVNXmc/ljk6X
jo6uCN4Ik+wB/fKbR9jtAIzFChm8dmjbdYfKBXwz+i+2G23F5W6FvQutH3+8FC38
VFaMSvTtEqjKYq0je2dPwL1qswlDT6Znv3Sj8tFGowNQY5KtlBHlnodj6z4FvS8T
MMEug6EbS5OxvOKUn62MckUWt6CLnE7gH2BV4hs+CubK2JpTLy7ImD7upATh1iTx
Ahp7jzODsKEPhGP/8En0gUtjYJ0YnoIi2C0VY0kw4Th3vim3t9fGTR+CyeDZ4GtD
zsowJb7zEWnXImekUQ0t0XPmT4XSKuNndElZTiqraCWyOYqzGvulfUxuo0Bcs0eh
3JrMm35a1Rn2Qs9VcVArTrQdJloG//EGmdIEbXa0XcXN9wIR53GPJnU2iP0/R0o3
1LWXHJiuvUInHexVvb3RomILHKex5S3dRfxIx8zw+Bi4VlO+g+GIUjqjuv6V4Rwg
gEFEJYP35k4SZGXXoiZW0rS/meQhE5XR5WWzmoLz46AlGU3nfQ/FTF9FcPgV+7f7
HtYSXS8IE109hTZVW4RQInOVx+Pg0+iSUuet3BAgF0WG8vVSQv8tXNYORk9N+shX
7+rwZNVOWOIzzSuZ54SkUzwdb4LXCoF4RKpwG6dBqSsm4Hr4Xu2ifqrceqg56TWS
gSdqYWfBoqiD9W+px+uCJWZXkn85qS4r0BLDLBISWoN/sV5wLAhk1V0ZSv3qK3g0
zWYSNbn1tNT2blSWZ1yxgnCsbBiEOyQ7aeGBR5Nwh6O7mJZ/V6CyTAyFU8U334/6
cQeQQEuCJGVcKV5tRDvWbJJzhzzNQfj0af3kkLQ+6Vn+IojEPi9OK3Sip/+HiiOf
6Rxf9DCkYR8EDdKlyC1IKr0JQLKMuLZxjNayhBLvRGLfeHQFeQe2z3pTGZJfCDgD
6Uqp9SZRbOyUi4gYvkb5Nf4mIIGViyR+n2TGFZQJAG+oMKDnY5bUdqMD+UO4NTJg
qIJdA3xMWx/SG4neIrXK76bUdLk42col8tztF2F3qo83SgsZ+UHWR5xkahvu+nsK
TI0NB11oXZqgP8xW22FlHmaS3NiQ/V78M5AQ0ndfYMNYS/eTOr6XAOgYqHoezfqq
lWIuu+fl60IOhMwl9z/kFb/z3jWsMGgB0+oe9aNwCN+14AyDJWuhoTnQEFVFqUj/
d0JLNqSM0/4U5/XI7ueMzL+2DY7OLD6wY3ozZgcAK4IEsOrsoU9eRMyZnPh8tlf6
gR4OprLBh0L3jDa0syOhmlOgKVKda0+flgVOajEkiab2k9acn4Bc1M3onOOCaUtJ
gcvMo+Y6w5QLKGowNwRpPo7SiqwnsJIJ/Qcl7W5jIGk=
`protect END_PROTECTED
