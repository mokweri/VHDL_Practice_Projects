`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YepEtSX5UZcvEmZV2j4BVmoGYBkKf2YjEFPg9yHlvjPIqeMSvt9YY9oRY0tPHyF
LbL5F4EmzVMWXaKfPUAy6B6BJPZoRXk2LsIy3JnNoXdikGgmGrlmtd8FGpemAk7b
bc7mqB8Ei4xhSRuQxC6TarFOx20xLItGHj3Y3xmxDBDG+r7ivTKLeV6FM7gaPeZJ
NiwF47wPOpvLJjN0zkO/DAtg36WmHGBBuuAkMGUhM9UJAJvPNQJWmoYD/WV80XrJ
PjQyn5N/Sd0+iVmzhnwN1iAG9iRzjFm/l20AFBPPNw4hWHDxMW/8rd1KxXW+XfrE
3k7trgkBQSY/ozkce8+94utpOBMJ6RUQ0W7ZKLSVSCWTwJiDuLONX6iat78Vuxkz
EggArPLMJJ/s8L8X0zNkeE1pJu3US3/iSvo/gLuVMT9AHjPx7OEBj5F1tFJoYeVX
0Lgu/UO6YjUJ97WgU9/jX5Kc/EbUtMosFQZXzy8gSNhmpgIf0zCn1xSPduiuSuAP
5994mA+OAGUv5Ce/oDOtXLlFBeEONJKPTUHX9/Nnhh28xmWoQqjsOesH4EilJLQg
90iVuHz7UEkMzsc6IZ5dN1pskOffJ3+BosRvEpLUWHmQrUw3VmxKqeiv4XhemAf3
czQuP1X43wQ3olV0klH5lPVUilsaBYzSHXA90UFVb811XNwCkjAINLtpB+lFbJsG
cfoujx5v2FJES8sUBHfNMemoqn7gzToh6XGPwP/YpwcI1w+MhnMvM6pEZ2DnNS/e
VwgmecYg6OHat7y3uIQrbcvWBR2bpSDuuuKmzEneijnq1HRGRcAeaqzP5GI8U+yv
1mjOE7rO//ni4/bMqU0R91X/n0aUx6k7r29zD9es6dH0PJYlEg3eiwpi+/mbfUL/
GgwVaKciJDCTM1n24D0xNr4BgGPZywSSZ9yXZ7BMFLBmRjEwbrJBhgM/5RQ6wBc3
8nRTXvTS5/2T5JmAkoZPmqsMIApNNpP7M2SGjW0PARqNhhXqxFz5pj+Th/0keJeb
LbXqBYW+Nyj5WjCZo3uS3sWVTMWMp2WzhO+jZkohKfngB4o2xRBJaxOUOmp81NBP
JV9xpKbFbsjsSPGGsvMWmLMozqj5QbUQCZnlS3yuVHbWyz4OdNIpUIYC8e2nbALT
qc+U8VZLCsQTJHPON9H1GBBGA0dujYTqgRt5FTnSHngrBtZUxE1AQmDRGgn30Dy/
xtTi3jjUeoet5H5Ov9GKNPrVVQos3hwNKeHuvEezilusVLAhDxv8HnqY3hYUQuUs
wcuG81ATX6xh5K0DYjLM1sVJwp0W1UkiDuVJNkpljIoW5+8Gf36dw7TVdPjK5rHT
Huvizo4uNeBLhynbeo80vGQ24NKtahjy+Df4pzQhHVboFS/tyXrtBYXkrkSqetCz
u0fTtcrh4cqQEq0U/z5oPrqgjBLfkE77qDIH/SEs5gNdUf+4XDLpX0Y5ISNr5SpZ
/cA7rPLnu3IhD8u38c6A1H82INtggGFrNALWNeyemcEqVkdTSwepSrQ2ZXPuPNlK
okWNx7CQbrasK/djqjcXqeKxAZ64wwWmxIMbyVlCU2J6/JuCojXROxzfD0mk2Upl
/9bViYY+tvh6aY6JIElyAOa5OYvuEGnVsDfsZKLRhBYaYUPzZFgS3xVJwaMCHXPP
yoJUumbjW1S+WNDknkbzXg0Pw6VgueyeuoN8PL4ra6CZq8bcdOhseOA4VegQKbci
4y90hhnP1l0cI2ilr43hPcwRws+4uMO9k4gMkQt+7e8k129ymyp+OpyzZk82BqhH
lVbIgw5czUCDWjtrGyGcXBOtFa53NeVyS7P/SnrlrZiJNUi2qjcsRuxgFhk4XbZD
VBKmNmIX6x/QgxFK5kl8NoI3PPSJd0WARt2biH3xS5/+leUT/BHDA01DkH0gqJOk
zQ0vlk6pUagCNYPVCZyuNK8zj4Qi1DCezmwh5LnGTzFvLjciQ543ie7OdHDkj9gM
w6HeXhFSv/Oija7CaeABbwxYfKTxcK1bJc4oI69/Yytp06bUNovZdhpev3UnRunn
TfXT2/6j5sLLiXi6faHuDmijVhmk7liyiGZ7g4nrI/j+fPR374UHv2Mej8gjRa4I
09XwYbOLBfBaKun/l9eSw4oF57dvCLK5jiYXXORxVmvymUnwOXAseSVEA3Elk9ro
goFyWyAL/N5wA/OiEpWigkounT4sdi3DtVxt+mawQ4q+pJHOcHqTqUoFp1bzleb2
8V3BNl7anwlGAkFMWM2+T3Uip9y2uWrOmj4DI6bH9j1rRQz4dCxUoBQxBOUmDf35
bMnoY5Uf+bFaCxp1i9lSRThV9y3Xe/HQ5EKHaBpZqCHAN/wRfDiA+mIq5jI2PDVB
mPf2AeQdarpsEHKiGRvsCI1UdZTvDof2UNZkkaS8zH5d92ynw4BYMqrs6b17FBQg
e5yDI7jX4Ok8DRHi7eK9BdnUZP80UKnA2Fyog4UJ1wOf/01X/aEZ0c3iNl4hR6Ib
H+LQEsH2M7suPVkfG4Rppa8U+Eojs77Oz0bBSuybahP+IKNSn+11VKhXVw1yNBlE
sLTGpfOfHDpetcdy7M5VG4prVu1rRwMqf/gj4STQHBr2Edq/T5YH9kEEDQhmRHIS
3E9JA1g2XuednRqP08hzDz3KKR/5dOyQubu0NL2O+9Gob55dFZe/SLznhZt8nAjV
zdgx844+NBfwidyj7yF+M0EYnGrWNHNC6tKlUY6D12bfn2h9HL336jwneBZReTp8
kXeAcoYTW8mDGTcJAbpyR29b0wDxFWp0PXZB/xMR+iDKFDHgkS0HexzdjIn+8mRT
I1r+asFIMw+tT7CmnjK5ibC6ODwfdS6OLZJfqYNo7TWJBlYHDHVeWGTj1a1qREI2
9YheIzSgeO5A9zkGHjclfGtZGNwm05zLFoypz2hZgGMyazwMJr0PqdBHjNAILPYc
Pt/B5Ht/S2PKJdJtZ7xUxrac1h2Vm657doUt30VbUOR85C1QLcXHjRdgrLVi5zJH
VBrwf/vLqZlKhoVlnomgH3Ub7ytA3+4EtqU5d68xRdOpHwgsbBfRIYgZ26xkW4QZ
pFBYblVfrUcfOU+Fn85cprMQzMAblj6kGoGNC2qUqBG0VPHTs75BPp4JQeQKxrej
FAZzWfFARrekKhsckD1emImQVuAW3O1WI4XI1TepP3DWc1yRmvAUMtyb+C1kNTzm
x9V1t5D0kq1muUVQlbXfxXtZ5ixtaBx1AhyBV0ok9KEwoOYdbmeeLu/7973mwJgP
r3DC5vswdjDeY2q/RlN1voUcPaaJBdWiZg6OTIhKlPfYq6xd92/Xqw6v9NdF9bN2
ZhoIHZv/2t0COkNOn8a4Zgz6zcuq2rdRF0uxgNxlesFv0PAtNojqzzNijo1XYvKl
j3leOmlSpdi53lz0RPx80ny6g6CQzYPUtIv7JZ/kXqtb1hHNbl0M0VE1NNLtw3jb
tmntAKiKUTEjMU6eHaEYxC2SRSHsbF+w+WfdAn4rMdi9e/nMYJt8O3dX6sK1hzOj
hChU2PlwVGYxrKVnc2zye7ndF9WlhD5VYZ98r2OGWMceNiyKuEuqUbq8eTTTu0Ws
aWxnK9vDwKH0h7NEcHNAdlLIHkuW3zXS6hh0ThUVrpjfZT/71CxXFsTuswKebpY2
LkZZswKLD9Jn/ReqS2TtsnFt/u44XQbH/BxVF8Iz8l/fmKvPRSq7CCqOn7PMpszh
IAcrXVOPkeIUJtMR3dyC9308rag+agDfCS1PMgGQUW0Q3i7EgCLFoDmeGF0oeJ9c
UJ9tODYFo4FEQlQOZqJmcszyEFPbFatG9XeqjHsbIIUU2NwIKtPDkXQBY8E8ewiG
5bPUhDgeGflTx2jM3f4bZB31zFFEhjRTgAcCHX8XwTjZI7S14pH7y1yjxFXRRD+P
ccsceF1PY4U8qKhbCQytauQGiWhqwxbZTdj0MdUvDO9Io7qoTSv1VHfrLnp8W8yL
MPLtjIKPrxradJ4ZlJbrWuFGcv3w7GUQPQgpyiInaDVX5pKVfxlGLef5nsLkn1HX
pLYr2cP2NtcBo4dqKgEXclfjlg59NVtli84BgXiRY30/30mwUouum9l/Nx38TB3U
8UeXe0m0QJWIG884E9bfXPxl2U5fNHUn+/AgTsfbNzGj6RsTbA21jx7iPBlfILDO
6YcD0B8CgWwmEoEvxiXw/JyjJECOjogz/6GDVqJBW/Xa/Q6UkrXJcX2Sb44qHDhd
+/fXDVLhx2HZcmQvpo4svu1yjEaEJqlbugdDVGkSZicblsbZtp+RQhKYfFcpq0KP
OS0SbrMKyhZLRi3db3OJPz0QR7i7hb9+qHR1nO+5zPnvtsd4CGnZLnxD5b0oz8xm
XynqlWKGtHjYyQfN6EXCshsFWvllVvljNujY+Y0YcLlpTR5f6/DuttmgYFyScaoW
CS+HXc3P6yzW1k7N6aZWilZqy3bH2jJn6y8YyJUd3Nrs38H2hbTvKLmXTmlq1I6m
mGkbP5eco8Yo7X9VFLLSQ+ya2BNUx4o1yyzweXXXSVe5DFKvW0x0EBPWi1oQZsUJ
rIOAmWjl7M40QKJPUS2vJaZw+5Z6TbEANBYfYa6G5sVF0CwPDw5VPZpFZqWBSTqZ
nvak9jItY3fc3/dIl2K2UUjDiNoODymd6u40vHYvDO9l2Sdwy5fAqmJgW+Kn/gwR
dCwUeEy7cvO+q0RzqWs8UHAYoFb0HUP4+2ofJVKNOTcIBigVV5+3/sQI5uzekZzL
wPMSEoPVxiR9eZQJZq+jT4ZNrsyPsg0w7KLLG+SXDkeuYtaYw5Qj+jEzo1kokVjv
2edgQMNTSWbA99xbL0Sef7eDxBd6+Sac+L0MYqRIAzfd2oDISyJCNtPf9+ulWTlW
92RRMNsZ8SwOUbB7eYEyWZDxJsxkmaJzjPxFm6uJ/JRdc4uE00t51gGvpyofnErR
RXBNxvhtKs+sJw0Ef0Ub6ewTKAr8cxvhyAeaFgHTSlxDrrNQY7cLnoduzrrU6pyM
o2MGx1qbsYGJ7XuTO+Vx804RDSjFZUz1wxT/FdQwmBpd6abfMOAGs6UzYyP/8BPr
pzgbmuRBnLj3i+cX2lze0bqmi0iNNUScMnmAyC4+aYV9DS5RxJpozQY0jbxJM/Ak
3jypIbZYf61RXftD56JpN2eYshfplhwsov/XGKAbpV/rMDM33+ODuJHDk/RpYG5Y
R98tV4YZbrQJi3LdA68cW65aYqLH+dXNXblqjklEJRXFqtlhGnIx/XdG6ikwNbnR
M7WmnihKADmMfRCwYFp4qKwG3zrH7dvY7o2oPO1ameXJ2bABtycfysM1Vhj6ivAG
eZZUgYcaBnxg/3HwQQ7jA2wkcwSJyniprMCdX7tDmm+eiLwbdpjKNeSFR/nNquzg
dtQjZSlQUZmKU3Tu4YVy7wNxzFgAnkYkR8u6Q+MIa3Q7u/YnXn1OB44ELILlBXWi
LC1CXb5SD5eBbXZqrswUA4k2FDBT2bncdd9WhpvqT2lnZ+dxRAA1LlrFl8eSBpt9
KZStwwikyF+ky+Y9CB6MlsaGcXEx8yZLoMg8CTtw7qd6ADcZmV0E/k/VoL+bc8r5
DcvxhfLWpwNhjIwgDT9VSBKe8Zpp0HM9BeF3boT0EwZxAaYjqUGzrLP7+ZxRJUCF
qmDvNMqKdyj4jCe/Bnk8QfM0p2OHjOslTFtAq5+aLISrNkgZokXGfbf6T58mtgC0
0TlnhWoehPx6JfZdNb6UTZuf6RNeO8c/3h9gCeoYEJ9qsEUJK4n7VWvS/930aDHO
I3+/Cpy/S3XPOgyzSaFfo1Hp5j4WFI53fg4oT9bTRhhplG0WGZ9lmmpVVC0VO3SN
FxVmHzQIa1sD4NREMF9lGjsrJSysPnal2Dbuj16lRPTXnRnu2ySz+pAIflnFROP/
GP3sSbs84B53Eh4kJWtbDSdesEu7yJodPwCZwjF9Wj6P0y5hUBoA7t61hyP1Mk8z
xxKa0QbEQuiZZKF27sJP/lbAqWxgW2Jg5+xdCE+W1iMshbJhbNAWhXt9XYZpduzN
Ra+ZxuwdUT30/ks6l9YvnZPx1JXTPiojU93yvoyyiDn+7lAOdzD2ZoTeenGhbjVG
nZO83UklUIaZqc/JIqsy40sTeu+hmHXLe6blWrJRPFeiLEpPQhMlFmpYpLY88jg5
/sBh0OPnhqhVU5zGsMhZB8qZyyWhHds3DeonufeJondONsKKeyw2yOdu8RMpgDrY
NBQkmKSXmJOwflMyX+ehYzIV5SCA4x6cA50LuMLg3+AF9zMpmEIgq1RRSVstEHR5
WVH4YkGGajCy7Z3KyeBfDuIJ9caAnW5lNh/b6I0ixldZTp4cAPCNFD/dmnZ1h/kG
E8aEPbG5nEzgjtGOUR+HgyhmeHgZO8aiSOlt1JO9l+HiOC0ktl5TCPmvOQ4KPkrv
+S6b4PnlYNDbZQe7ev4YFPe/XNLPqaQhGD3k3dwfq1PeBt7CzU6EaFgzZO5vcWwq
fM6NU7Qoq9uMLwhs0U1uyEpuhn2ig6X/y49GRII293rgeBdkPuNEOkC4V1yJGOqL
F1pmeCvuv5yAYCI0Crmu6GlhFVZxyi/oD8qzZhaQc4LVkKEuYFvyWWAtEXoMTxK1
Zv+sDBPLoJ0cbffPnt5iJX5IAqQhrLQF9QnMkJVRvno0RtiVGCNQxmyom9a+lCmJ
PFc5ENw77qw5yYtbaCwxekGf5Yzjs2Setv8cDKRX12IW5UIB8hJHsyWmTMXom+8j
/OW1JJ7kDq2oYisgoYDimwFONYzF/G9MZsGaXR6RJfTA5znZVNJOxFjJvHqTMsDu
Mpt5oUn2EJlOzgXixuAp9a/Qd5sPyWPvrQnO+Ultcd/eTrQQik1/mbj9No04a3hP
vD/BnNrhaWoV31mvgcFzHu8hwcSrz026+n1fPQXJs8NOMXtu+RcvzywZ5Y2+1X5K
l0Zmf9cafI6ndOKo4GxXTtfLvndnTOSleOdEDvat2y5vgaBMEn1MAhPkBjSaQm6J
0/iAVoNZvt/h7AxNlkJGzsnwKwmG+czdKPqmVtYQWiGHY6jeKAdU30o94N7p4ARv
geAYaZ5dYJWvZbsjMahjbFc7awOQZ2XZhBsaBCJLo9mcZrQreqvVxmVe4C5lT4vZ
f6F/N8uJLvn/QWUrvaB/KNgPmK3ycyoYsX14vbwBebOxUyUFT7IOyoGKRKn49F4l
/eYtq4eYjsfYVsdX+QA4pmy+F2UkGbryUisg/RxRsdKSNQdy2LbeI2IW/dXB8H5j
/k5/d66gCfAB6b9PwqOJnsXXI/4kT+nzvLO5RJIzfm10KVBq9wtIrb9FPfyj60wv
0FKEuMzElGA+KW4LHScdfbygTn3T7O16F1mLPRjG4oetKn2NGePMeIlnF5HGOdIR
MZFY8FyZprlHNjDSeezRN5nhC5LS6MxvK/tKz84ZNREo5BzuL3WP3a5TP379/9vN
ZccYIZyu/JsC/EMG7hZsFRrxv374cfWfe0aWAGzBkRwpgIe/rk2uPSBQ0rbjv72y
wvXaVzouYHtKXUDnGecD2RQLOJ7afWYA5RV/TA+5Dpx9WF/A7tI1QIPDp91I7gpU
pxbDAB4Qqr0VUEsJb6c2CR7nBO221ZW5FiTBqdUEco4Iu0rbgTqRCRy16Yg7Teu5
fgzJGnFz6cSFtzEPzItizsrBOUBrUu7j2Jqhd7bVuuVt4OWrAR/Mix17Aq9SGjnD
9PIDYdSFguKXp7dxobn5hAATkUfC+rHQH6uKCW/0B2PpeD8Ax0qRO5wc0dpGRLeU
0hRuRT1ZyPWjoR4G7DZbkF0xzi2Zy4K+87w/1YYKTkAY9bE0nwpRcGDUuPVl74J7
0pm5pxhg2FA8nufsBvAqIAWOSfl97GrDq8LhDfj+El3i459GW4Cu6fKa1jWdENj/
u+L2lsJA9NIsoa2T4pvmM3v2qOFZ7JRDPulXjgB2i4NMCdUBeLJpgUAEXo3aPxh3
gAY3onmZ1AR/sJQ495Pak1l8dfr0l+YUiYxMOvwL8KYMNLyFS7uNC2evKRCkFuAY
IZQax5LsNozEw8xApQCou6eEhXzacWHhAHr/6AUV1h0FyGw9qLstL7RFUDexugpO
IIpyYtMYo2Jw8g6Ic+rOaZuxpVag5W2+/MFmkKRJeQy2ftpA3UIDOCTT+83ctc2V
494I0ggOostR5YPhsVoEvVQhZGXs8mHTQ10PgV+MvdmFlwKkEU5jz4xjUv/zo+7J
3GJGtJ3K0QzgTfTwEMapDgLtG7Ua3/EQJtDPL1cv8yl1Xq+/i9g1TvxKrmMc5Wsp
bb6q5pPxX9Q6gUN7Nku/a461RXHzROyTrC48wyVNqe8rrmBXmL3f+OzbY1za4UdN
KKSIL98soUELrBQhIXbamv+IEdCh6JRqKnYzDuCaaot+q6ZJot+ZwEpEUiLsjiLt
n1+XkitFBDrbBoT36OKxSPKiJnBbiXjePh5JzCzWpXL5SX49VbmhnWZ/yss+3VsN
zbAjqO2fl4l8zk0U774p8RjcttQLtcuUiHq9CwFigcRzeVmWhjJl5U6eB1DwCF62
jhiUQawWucKtJkpIaXZRUwzipdqa8zvO1G653fPoFANCdj2RICG0pui+7sCLMt7v
YAaBIibJgcVOPRTOqeZ+5x2xcSy//ZSd55ujnns7j+G5qtmVrCJrRbR9dCjdfOb+
nfXK3VUo5eElBZDR7PV02dvnFERyr8Y3HcM/W49f4a3YcbXwMZ3LxGA1BBkPU5od
uAR/w2iHh/LRQNRz28Q5luOH/R868sIO7YPhtIn+Ehj4KaAOLzyB1ibNmhGccHDF
NLazl7Pnem9pzgxEj2efK5+jFHLsdONERZta0qr7iGeq7AvR+L+9gAgV7vMVEW7h
Azrnjzd4hgcu8ZZa6KSKVSFTCdPTYsUxSwFxvetGMulRxif31Ki/4Z+I6CEiaYYH
k5/iNXbVNTLXEsNF9VKM2Th9Us/qYvSMo1NPgmSkm0I1oA//kdKDi2IAobgiSBUJ
kVoWfrLAHWLn0WCO0y0YWbnXl2q0BFn/MrB9B2U5eIlb0ynJnwt5i1Zl02FpTu/m
QgF32YQwqninE4F7WoXdA2ii/eneiZLGKUL+OcvBZIXv7wvGsNE5OX3ask22xxnn
XeIah2Tel5aRQqWbc/e8JKJvwWLff8imn8IKqXYiPNDJpxiKvnHAlXmQi7UqHT72
NgB9sXsQuoreSWZL/V3OpcamgDmzuTo6INsb3RqdvYfWBOUuC6x31I5jejKvjE8a
hx1yp4tZP9hOXljVApe8BCgnIiB6phGQ/ST4K72qetTVVoMyUvvcP7RkW+MePctM
kU/lSQQePD89cs+R3jS5+blJeNSu2HcE4ciQvqwjGrdWcsC+Jf6gC903PSyP8dZV
4Qh16B31GRKvKti8TDc8nQMwaEJOT8+/cnRgaA+6eMfg/MkniL7MdKQIo68pDo6s
hPTx2Ikqgg5MPYC5JaOclo6di5C6A7gatg2xlTZ0YqDn/lexj990V7BPW8ZZxKqq
rpSMHm78KLHXygYPSs1/hjbPhQfE6x7hG3POpDEJCeIVC6GuYMWEUfTxqfWVa3om
xX/VLjo4629zpxinXg8BbYfmytiOeIwbpJhqc/AE7dQ2b/tDNOmhmv2bE1deWjau
4mfM19chj3OBGG3nPA98ITyVzdk1o54Ris4dxggdQ6HwyHNOXfohQEed5NjKvn4R
UO64jezl3/oc2fiETYD9BhWtx5RSgfUeleKRf4X/41HPKrPc25uS+8iptgTbws5U
o5pYsj27UhleT1fK0u2fAiOM+GYMsMmaIi5ESyPhT/goGvIw/N5ALHYF5dZd+GRW
t1Dpoj1r6NsJtK0Yh1UvZe4kXIzpkxvT+DQ3SnOt1/w=
`protect END_PROTECTED
