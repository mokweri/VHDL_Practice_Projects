`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4tNK17nhIC3QuZ8ptPainpiaMWl0JFpVwTmLctlEFudYVtQN8edfCrif02oP8o5j
eW4Qgn4m4Ft8987Hwob1J355GdQ1p871IuMfFqyCX3xt24xpf/T+PxgZveyyCLGM
p99ej38Ec8MdrAEScIyOvWUJnAIT9J4m89rVFdrp3U7L962KAWu0zMgH6XKiQY+D
vm4pe78Ns/AGkmdSGWuRUL5v3jC6NIzN/5JyI6sUp0In9e1i3dYM49cUo7oU+2ah
lvOaw0FPGHcIkobQ1yTn12HQoQCDQvfdNJibvL+x7FuIzhgTSwOkMWnGWamxVwgz
2W1rt22wICCgjKjd5FstXBwllCuksyQCOTn/9G2xIynYn6WtQV13oyIvA1EwnX5K
5sL5pRbW+35ejhZjoHPFAEQ6ILO4XlLnTJTd5i5RTP/hyeGdIp7rpJ+GiVoeFzge
cM6xea+aMO5qdcPeBHZcSfQK7lJtabjoEbloCfK5RPK5SW5xgp7aPlmLCSGmgjMc
bcwmMKkpUSHLj8fLXtyKHv8ljFjS7JPjZb36bXS4AWZNU6XAKfKPh1xqFfIEGqLj
fQeCJdwjox8bRJYCe3GJWAw+QOot8cnp9V7jSsUoL0hVqnhbvyzOiI929qDfWCyF
GC/oMBY0enA2y62tSjvtzmsEpE7DjVFX5kU0lQ89uXxS6j4n3UEKbjt7BIkgDGCT
XQdJdZGs0kNgopaadFWDZdOwRvZ+CArIiY57dMDBU4LINoG+LZh2zDgV0b3KHtSc
fcIooszDZLIDQK/E4R04KFUpKG6n9T8BUh8H4XFsCbaTGB7oKC2r22vo04r+nogb
XKUWRy56KG4QOloCFr9Nf8SpIAvF26nGfMA10M+4O2D2n4Y5KLLlfePI7eCo/sko
FRw0AdKFaV+s25yg4TCN6wqcQUm6ZNq7+ICf2c+iv0qyNTtM7sfVxg+cnyIuPKvc
uhr0pTYmN0+Vz93INVuqQxakoqFhenR3s/K/jZx318ZTThztNyBiwZKT1T4AtpdI
ZOYVHlX1oahCRDEISHTPA2iNcgWE+o5BHSMiAGQqHgXaewZUiZFSUEHJ3X8BRShk
ZSGGcmWa8oZZ9xZTChE1NgIqsu9Vhyc98YRZ+McLZxfFL+CaLPWjUJQfUH/ZZbDE
5LbkGCV6H6s8l10NvizlrlNfMgKCXJGi/lBTfdHD6r+AZou2fRd9IuNgqH3gakae
E487IBqtdMb/EmJgjzFCNX2qImnUvJpWFT1GIJS6EQfbKyfVWCqFEUiACpKRYo/P
bNOFZ2P89XySLxmyf7p1NNVjnM6XeYFiJddRLUzkXK49Njua+VrPXgK/V2y9yDvX
lxwBu8ibIrRvmHdTeleoTegv0qtmssrwnQUm9Dhlh90MHDSMXG/+SH+swcPyzbet
eQHyF6JaaiYMz0dZI7CUrBFH6xKNkvd+Mp+NrTrHFBsAe/5bXd50BiR1Ekc/v/Ah
G61xlYpcRDyqm5t6+f+bLQaS1DcKhHNva/PPOo+5T5gL5ierKtHaJRlTQd5u5Jsd
NJcmku4uWT4MJwLkJzZOR55wPRXQlEw45RNTkeYVB5CDUL4U/kpaCiydDyLj72Xm
reu3lmG07KemBqYN98NxnceQG2OOYTEZ8W+bpb6l4PYV+DBHnYxgwsiMWM5JysqV
3cmh1ez7BC+2TkHaSUjELuGMghoxCNj9NYPwkLyfVbARjR7pI5vZEDsEanixLoec
r1z7E52F8N6RTDI09JmRyKNcHdfKA1NBrbkmuHmUGyLmyHsuReRx86VvdgPIJ/mJ
0j//S+QgQmuHnszFwK30V4kd+FeGtMPLudKWf6+8HYTI7E04190WO4DOpChAz0hM
`protect END_PROTECTED
