`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oagfihk8vN/aM9K0muae2RyxT4uGu1+07VA9m7aOHPuOPi7O989qHupUhgAn601s
eJG+OLGK8ZH7vxuRIX/6rbQ8q8U/2sPVgNLwGvxhT4E2ZRwUPT+VrUmvz/VI7Xds
bej+GvHy862565+iwsKYnQBBybORpY+KEouOPZF8Ymi224fN2urJqqXghHO2MYWT
mWF2I0iiG1R3+tNBdRanwoSCf6uVLafJz4R9uKoS2l4F9c3bQIfsHWT+ciVfoA9q
y/bvx8S7JbKZxbbDlFPIOx4ngnznA08dc4uMwxIzF3/X80h+VBAYK/ndahBzZdLc
JwggpC/R5dh6G+4u0Wlt9wR6lQgHOMf+P3ERtbU8yozWaBUB4BxWyKXmJJj7g6Xg
2t4X66YPQZ0eC/EJihZCOsWk9yg/6rIpL4pJnoaQWO9dUaxG+WL0aiOPPiug4B9W
eFfCXNHl/iNjuG2NvzQGuHA7ItwN6xDLkU+uXi3n/v3UY1My/FJdOKnbYgCN3+Km
RtjnQk2ObSZXZ0KNHhUKut+PElANK4Dw9hv4+yuo4ixNCfxzQsaCbEdvuZH/eY2R
tXa0k6mp/0yylHc4YT6Thlw4GvrQHWMS0+/0EFNC9Ko/y32E/wulyVAFtqeSd84M
V7W5vBjIixMO8Z0VVLLvP/P5MNeYHeSzaKCD0tjfrAKb62yjNOxR994IBYlTiJ0A
/4OVFWzgv+KkoarKkkp9JP7iOK6bmaS8GmyLk8I92cI7G4b80d73QCen8FcDs6Lw
1FJIHdlyf0nL01xvuoa2hBS7XztjOavJB0Mkcf0GBtX3JzvmZ8kBeRU2sblH12nT
ewVbEbbj8zvNw+cDd1oW42mhcuHCp35G28zi8aNwK2/feYGjQIYQjVFjVKt44x/h
NlKaetlyoxQVQY7F/TyJzT/nLZ69gR/XQXAoWBpGPAtPsJ/YuxdhD5b77S78P7yA
2Qx8yB2WcGYSWwuI0PtuzutTBks0kGCZhpUvjw1xgvQWrrlUDWHy8ROc5WZoxvv7
zrUkirtkRC9FgfUC5WM9fd3znc2W2QbBVp2TnNSPb9W0+akErrWy+VBsv823PjWt
KfZuOOXnttBSpldxhyvLCQZwPPcok3OGkvgmfF/AsyIKUeS5iiqRAMvjHB7IXVW3
nvJA5QJT4SYEsnvBj9+dFhosqKHxbthVZJi8VM/AFl1+QOODY2WFvxkw+FLo5ESH
bImOuhjbufiRe4NTX1k8hVR+u/mzkaTi7D4hgx2JjH+cbMomMTZrTFzfyFWjIMdk
KDgp6TciK3QOLwe2f4QnfruqnmKeLoalrIO0Z6WyGpTbyxrsLg+EFOqkCxmMvCAe
zoc6gl6shLeTu+IYikqDKNeo6WGmpO3n7KfHHVR0EhR/EHLCXYC27iPxegvxSdAm
Uz2Mb+q7Y60Zp6IYKkT4mehBrJV1EhwD4T6klIZsMuoceNp3bZ1cOveS+Pp2U3SD
Npb5c1c9hZAKkzkjJ61a0opIsq4Jt0pclr0+eWfDnl/TaqjlXPdUm45BqHIOz+qC
pc7yVAWLspBYrJmSnKAgpLpBoM4BJ5kPzR1hbAPgSbrBY/8sK4EHTICGNPI+Bdmx
bi6bLAL+z4oU2HlQvNf/Acg81xVgnuTJvea0bTRt0qAJ9/ODpDH5FJDItWAVsOPb
l+enX1QHhpvGvmujjfMNXw8d+QhTXUo5teGcq8lEQpEqs937Bd4nqra6nwI4Y2uD
734zHihMq+PTZ6g3aU2EaoXEAAzPm8iOmmLKmLfEBFEoa/YkVK5GbH4ORSE/PnYx
/lXjoW2QgEL+OtQlugG7YL2YXknJhgjHPmbarbVVZ76PN4aO37t86u1hvWO620Nj
IbzQs3T3s/aOmfvyHT24dfl4tR5Q/KuVCeTMRElEMhHhiPt3iOEtxdtDYtMZZtU5
+vac+Nt2gSHic9AS+iv2mhhDcP9f3dIeVoIzsyXvkilhZRsxHCG9Bo+QKzE1C4mW
Bo81pkPpTfnpe0UmXCD2+kXBiOgBZUlG5VD3z0KUjn5oG44hklfZ1d6+VrzIGM0J
X8zyJH21gXP2IjjP4fpjYA4cMXrzxiZtCJGDxibByfRHVQ6Ux32wsXtq0YR1i89d
AOt556HQbMe1LCRVGeKQgqATVQVcvOuXCzSuwWuZlKOl8SzOGUKyPx1k4nlBpjNm
zCpj5rIRHgaePRm8IthSwsV6sjXR/FD2hfM3MIfZzpCK60qOok2jM2GGEro0KOoR
hySmeRXjhqIi56tgaY07F8W1WNb//gU1X+KmDoH8OC5U+Xco/LtfPDe4Q2+TNMPS
ykE1ug6UiK00V3f/IJrpC8/cV8/aWqrGrqw39hff9diq81OuooUYipD4r8k2jw2J
ALvAvSex3OoJUKKVQVrBaYysXgpg6xHzMVTTQHeGpX94lNdw2+2kxRfVMMVfiufC
shQ8700NqCngbKkEBcxYag3Lh6LHuNpkmoXY4z8f8PAhdaI12+y9M8UoN/h/5iWp
ZlbFXnnJMDV/3jtBkmxnLbBWZRhJavXrrgrcrZ+9yDKYgo3+jFqFOcmoBC4NZmYR
`protect END_PROTECTED
