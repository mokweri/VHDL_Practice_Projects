`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfxEjEuvcV35/ZFDeh451LetSJ3ABcg63PGuQ6fwj4kUiypp8jrkDFtK8CJWKOXu
Ea7EVxDbLDtC8q/581GqCbEAFQg9FrStjpplJqBOOzivAmRu5XZw+L/cj/jGIFTZ
ZQhnyUYB8UiF0Gb9Zhbfq7Cq99wzdRMuKmnWR87rxGMbOkQhpjmpQSiR7NoAPUSk
JDT3jeNuhZ++WHCIOCoL18Lxl9Cjg1KCUbze6awmwNNJXgfcaKyEGeFNeBFKYA1q
8mQvvYnKi2aaPz+Z/eWMJoso/1dD4F3QdS3gW/uXU7vIdnY05dwM6vyXm04LrTP6
2N07u2f2HUMgfol9/3Lv7+f6LWIZ2ZnlA9dIzjhPnS0Lgs5m0WUFa/catp+AvIuw
k0hfYCZWaNYu0JLerdiTigySCKvpkN0vNx+AEWDw+NEmdI3UdqqBbk7k4Mz+mwKm
qlG2LG6xhLCbQGf7SMlvU4yiu+hKn/Isvls8waW3FpV6FRtwtrR7Pqln1dpOYEI6
Dg/2IUPHYQ/zwMGtCbHNGSk4w6yx+Wmy9uztUyHzdKqAuwl/NLgP2A8Zb81sLyrX
ZnDbzWPsK93rTXP9olqjIuuBK7aW9KUf+Rk7d6aUHSAkXQwMgMX4AlK8LWqrWue9
0IqFYNixVjALwWeUqWwRVv8z21Ia1Q49Ic2aXOoZ2w5dBu3QZ/e4wDhfwjJCu7qa
IUuDVdmYnDHr9tCT/X913/lLn1jWe47guU6DtN6fpvajUcg2+hYW/ba32qvafg9h
MLBXVsm5L45+ArHGgPZ9+B+iGX/11jA4tFLcdtZQOZpslmTi1kpbhArqMhCObW/p
Yu/rCvd8FN5SF+xS0BuVm3Z/C94RqpbKce3V6oBRTWSwy7jASIic5ixHAeEHc5Wa
Ivg+ZGnS5dtFzuBhoolaPqc65OTwn8JxhCUnXVAXUGAXEfzHkxEMc3mlIS+ny/BT
KRdgY02qRV5ZTekJeA6mYesxh4llK32YDLZRFEIY5qd9CcwzY20L5Y58SXsKiUOs
SVBxhk7W31CsNj6CEiu3ozQdx+Zk03eakSaUex/fuNsBnLiYYKCHOhpwcOnnqoNk
PgYpct+bDrh/BEv46dCGTx05lnah/8wQEFc2z9Lhzwk=
`protect END_PROTECTED
