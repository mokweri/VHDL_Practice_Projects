`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSY8S8HgyRfKq4B+6hFeUvqAx9k6o4b2ADXMYpu6Teh+vv48e+ZZWF+plRQ5sxVV
i+4F2cqHwAAcpmo/b6W+ewZq7go1D1pQYP5pXtxj5OgzsonPpOiB8HHmdVoKm4E2
ejkPWooXV04agIYm0KDjHeVk8FXHfTU+aWKNPrgdR382XsNd6zHj2a+cBs28jSyB
561n8jYHC8dOXi9SSesQP0gXJnHvtcKivqZotQFsntUiEPbfHiaJrnNQS3rgjTrt
fvqJGcYgJMiubSjqKh+hl4sqsZd2zMocXnYV2Gd3Iuhj5uPa+hXOtYatSud0V/Oe
NWrwmob8pbWnjBb3Q99RF0c7Kxnk5XkbLQ4kHOOib2Y6jzfXsPPFWZSa60dTM0Ir
ko9avaCuy/9IhCQoenE7iadhG9CJGEDEOQwwvceh4rkJ2RXUgoq1xlpqZqrBYMON
kSk6qsmW9TZCTg5pb+h+JGCK9KrZHLHX1k8o1TbNGdQtUF+MtDkR9IarVA9zS3vz
IYg4mYp7DRIzzsj6rIBl3Q==
`protect END_PROTECTED
