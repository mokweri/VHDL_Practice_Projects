`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7LUZBteH0/6iv69J52OZd7ngRV8XNhO0XsJ4vh9KkTwowdAon7Xzt1GsqIEGEQYA
rtV7LHkSDdORbmzHNc56utbfWqXVOp54d+Eg8Imwz59O+DXbOpBPu3N/+8iEooj0
M8zalrnL9pTEO9WQPIMlf8LtBxOEUja11x2P9gRIqZv2AglUbOZUSlYIb4js5ik6
VDBikY8SkmopRjeUI54DLEvnYck5m8F5hJ2FL5lt3CcSAuLFTp+m3SwpMvExTSTH
9/jvRz3rskk+E9YN0Q21hg==
`protect END_PROTECTED
