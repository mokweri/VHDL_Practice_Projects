`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfiTqWwvAuCgs94kgrOIQRB4U67cpf+DDpSl4HvKl/UWGgGzfhBe+QS481mv470D
iyAU+JKk6FuHUE03y9GEaCL6T/RbXPrTB90rNrTyip2EJDr2No5OF3xraRZ0q2+r
dkpqAXQ6qnMXCLH1n14ycT5PCKbtVhal4eu+eNfktjuNkPO0xjdk4WG2huUVFDyr
rte97im/lT6Mst8Vtrhyd45mdR81nr3BKFFaHcoU0+yoVT7NnNvoNt+IoGrl3eMP
yqNczUzqLYkaRkCZxNyf7VZemUDNnT70edtlZ09KZLX25WOZure4BOAVPxt0OmjR
Ja2jfXNUo3RVX/T4/tyt2KffaOcI1zvk3HreSVUovBVA73slDjaDo7RURG4vkQTp
SQGT5WjBVqh51m1MotyxW2mjPGhPFn/vq1lC4gYIssQQ9at1Dn7UjUaRG4wP4cV2
kt0Rb46l70rBVNEWSyF/1I/FGvVhvyj+fqNZgdDYr/HgOoIOFXQkZX/RjYiqxP9T
ABAN3pHBzVKzm6sRvlMbRFtgM2lOpry6PUQ8LwHJhLyjib9KN8jqJvajUHpV+/5R
nBLfPctzBpvkHRG4vTnm1+N5plV9wZKw3zE/plqsFOV6F0rDPq9qn3CcWU9VTa0u
JP2gJJgkGjHteL1VQL6StGsQYvCFDiZRjBWjAcYeXtO7P9kZ1IlLwtGZi0XGDftW
/X9xI8PgIr0bFdnKXHNX3x7zeb7MUIqOx2JmwDJlkEiJBfWYN+UmUz+0zk65kPgc
jRBuaTSRmJqJoDXlJ1O5wceSDFiPZ40vRZRoXdC+nVm7nUPmvq7xIJLxXssGHcEv
AukNKDfZhM+ys7rdReGQ/aw1eNVRyn616cT1we2lua+/nZRmW/UjuR3ftlm2YXjg
btq9VAMtxBP3J6nmRwxBRIGp+XlzfRHItBK7RDs42dXK0yCROwiL8T/R33hu0SUh
fC+L8aS9FofEQAKyndwhpDsuQ3d6wpEstTZQkYihFNMfylT/7Shn7rNWjy8ODlOs
br0Ue034wZgPxbBvNxk+d/G6Y5eFcO+Xa/ko3fYtajYWdHsOLO4mEJSQXNJgr1xm
VxIW0X6JCIPhtm4MN/U3V7sO++eQ/U1IwC4GU1qVQtOdLfcB4tQouGfNgimpUsbV
a5eKtbUWeFWtPuY+kOpEPpQp4aUFCgeVBeZw65QfSDd4AmVzYv7zPuHw/WXafRd4
cYYiWtT42K5550ufQn+7hRXObO8dDAqMIZZqz84GRcK3z9pQB7Lyhvr5tkNd+uLj
ADThrCCl+KJ4y08tMiV2eDxDPpofl4JiTc5NFeR9I8/d1cM8oS1sR/Rg+8zxm36d
aRH1mO1cT+QDylhA3ugb5cpsptS6jMFbfQ5mkf9TelVkiAifbEPMIizZxK9hLurm
IubY5GEU5jm4LrZv1vu6p748osaOdnGu8FB1zi3Z6E0DIBw+IMKbkRyibxqJ2gyy
CdEcw1Kh5R6qytXEZ5y2GitPrfQsw8cgfQ2hiKZy1eE6XPO73fTMl2kwy5jyBF0B
OG9nz1iPqFK0bYZynX/JXhOHGUDNU1L3zJRbEfb0d8JL3HwY/3lBR86My6IiPCfs
HbOA7zUPTbMRYy1W1jclJMUzlCe4//pdMOlkJdm79449HjqCZKZi4gzyg32KXpCp
MUa3ypiF25ZZ/78Xusj5wuAhODqc277VSKTvr+QtPERrarl9dsb5uWBo/Zp6QaHH
hEvV6RQXGm3S1ADz4UqL7ZOQ1y5QODptshK7zSs+Ca47SFddmvm+9CMNrR8uvQA+
7bScLCLkcrtP/G7wbZ4pmdWjdKj1IvLOD7Rr3iIMmHuYQqXzYE3GmKJx7B/UZsU9
YIN/y3Ltx8dURXyFRX/K/8lqmNeOEAabsqONNuCx0E5fmuU9lVyeMLFBryVAZ9Rj
H40zOZmAWKO6L2Mw6yfudq9fPb681NxxRPKeZEUza7jUc3+AbeJ9ql60VwDRtCtc
+ESrtvdadlU0cUdFSZq3fVB6dD9tf4XbafIOgWq0clRE4RJQlQnbs5I/l5Q37X20
EDUet1i2urAQ3QvPrK/TGtsZYX6nzG7Q1rjEI1SVKYbDmyazHj0EMOx1qOceESQ2
Oc/QNgTyaDj/bzR858lHWtgO2bOg4m7OEoaQSz7s6XOFyZTlv+AVCf86zQYDZASy
1cVUHq1IbvrF9gI3/GY3z1BeSJa6vROWMnPsqcREDPlKaj0S+5oyFODRnUqImzT2
pwSpldKvZGpJAtZWDGxX86M1tr5uxsQJh+FbCX4f1dA1/Zu59srt9kmw0tc8hH7j
gBjC6nKTE8Ph3OXlZqJNAKNS2olmRN7Kf+7hUl+ao/8uL02FgcFaP2vIqZ+/Lrwv
GydjTn/29j2tL7XNm4Q06NbcTce2QjlIYmXGBmOxvERLdKMJi6ebIUBa6pqL68/c
tw9GPZbMPeoqJNJRnx4wFg==
`protect END_PROTECTED
