`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6vxSHh2oH3Thcojrs/sM2sLmqTgdJyJKpmoM2rNyNAoHOhHQzfvZRVLgyfSKnkC
aAUx2s26bsxeuVv5Kbtbp/WDg4QZ5x5i7h8Z00cO7JQRgrkJItkKyolrfCk6/xf6
+7dD/XIASLdOPuiKTjvDTXDRECXs8BQ1/kvNltwnEok8QlO3Dof59M/a+b5/2rcy
mfnBr7LatU2G0uZwcGN2KU7dU0TL2xrB4wFm9eUkxOEvOi9TezMzbkf7dqq/j3Uf
4JJkoRHobEiFOxye5zQep2C0hIsm2EDV8AnvjNuXIF57U7TDAsJSpIYCCQniIgKk
fidZeOq/QaxEGSvXMEnggMj4UiUen6jTqY4KHQNkzLBZ8ByA2lzK65+VO/t5pRoR
jjpZu3jvpsyZ49iSHIT4h8N1Ud72I5LvEl9qAf9Wb2jqxO/n+k2wbmHGanF5f198
1hNsnrcmIoL38lf6BWhOXJ37hN5rTUJRiobZJ69W5BiYX4FyWxsI3ayUCOh7IpCf
/in3tt5Q/1+unqIvPA3e1hbibMSFUU+8WMrFb8ngF7SEHP4ZN+IU+mxnix3O7wDx
ccCjyTO/w6+6Kqwkd85NS+17Fr9o+XHOb4DryRMzRLLKjK28qH9tWHF3WEdTOjBL
ZAjnnLkh9EaM9X3WTwo0N8CMSU4XfTdGpUurqmHAFzP9p1BGJNrau/fiAQXfsa/9
jLQr8FUOgJxoRyUti0i+ASosfgtXySOlP1U74tUnX51cgzrQYtbk+IXsKCkZBIxA
e+IsN6pdVh17JDAkGpKrMIPLeBQ5S/BjG1K+W9Ui6YzfGzE48akuj8oWYVC2RJ1n
rXENXgzKDLsggpHh33K3sB6Qa3ltR84xws85SYqGstgwBfLoG2NSf6gb/OXsQRKs
/8wankErnfxzics0MedpwuHO/KHMwL4WZm6roH7oiVX6AazWT77ox4nAXdGoOiEC
vxPqy6s/bgH3Vr24KC0ZDh3Go1nrLEtg4KjTjxAVLxrqmt++L5ZKYdQoyd9rDFGr
L5bNsjJwAhslfY/GfVIPpcZa6L+17LeSMOMcxKGF8vHFX4OWGPEod35ylYQgEYaa
z+ADWWIglr+QXcx6OfSggeom/at+wO1JTPRbZWPSEGozrn9LnwxkexIiSqt4FMJz
QC8Mo13bvKeXBW2alryQ+TPKHT/ss5PvBSxr0VleHUfKJ3l4llDwU7wvACsNR4WF
FBq8ALSfjUOkMW09OX/Ej4NGbRJEPMCP8EkjM4R80JAsDwp1E14eRJ01snhey/Vb
/z6m/rGyN/cslzDOhxrxaMPz9G8SxVS3sivIcJlKHM21AXKKAC+p4Y8AbQBenfKN
A2vxRMtk3+v8biLRPNRIIDxwVroRLwN+s0jJjbWwscaz0y16vL4SRTckTZxxAFOW
spvG6qq6WGcxGrGvmfkC07cS1VIGO2fVYU1kNXE/AVsjiqLJHWmz1gLntkygdJY0
cQGm4rJGbe60iMyzaz9KxC+AEkfpldMP8PcDhCL0Ig+X+pS3lBABfGCiN2NZeHvD
qI764c0cQFooXfWQvL6Md3/1GxdkdPV+CMkca7Dlybj0RXoYsyji4Z8CT4UilmpR
4RS96o9VIWRWVrRfK9cjfup8fOY82E7fUNzAatRSPtU5AqaMDa66v3s5k+ObV9Gj
PNCROMfzzpzmiBh+MXj6WYoElqnakzyfUHYv1y2R9oVyokXjHcPSLUPJdFboFSXY
JXXRnrKAtl8/jA1zTcKz83Wa/9krn0/9K6XXF0RLcD2Y0+qoXefBetsZ+S2U6I5a
EjQHwr+La1TAKspegzAIStsEGK31Q7roA8CiNoAHXCDaiRJiFHnHIMSb1HVOBHx1
v06OkZVSr2eed5AMw9QzwdD8yKbmTv0y12huwoXnmCfgj7PwtdtjBfGXSrSfKG/T
z081GheT8aEHV3oc5Sf+kh1P8Ffyp+aQHx1bdJefvcxRquRwtBB17NVVxWvDI3s1
2WlPKaSQIq9kEiJxVuHpWSrKh20E/S5nhKSqZpxUCn4nKPzK/al3aqoLXuF1Un6Z
mmBmJhp439mH9TleOVVmGOQrVfhQjocTbfDYqnNCoKcuH/SErH0HGyJoGAmoyfLP
9q/brg92+3cdTWppLU8bbe2kquzN3yM1qEgwkJItH0ti6kpZLtmkXbfBQ3Rg1e5E
a0617cXA7b3mpN1Q6T4ppINn/8K1+whT4st8zIwKqnRKw2egn+4px2RiJ1yOoA3P
3oEGNiWamHOQVOGd6nKZsKoLTKPiMSJ6d39YxomjBFvKAgETZZFmWsoQ5DJvyMHz
RdcNWHpmZL/5XAFT6Muqog+w3tqhRiiocrTH3v2IOor0vta79oRbkPG61bXktsK9
wcW6xYD6ojwMjSLFlAHQoNs93q55hWwjzz1tMcSonabc5xBiCmHrMivHhXr4AH5z
gFELLEbJMNleb1PdbQ0JIDZvYSeL4d/cK0tINRJ927il/+3qicwGb0D1uV6AUPMs
WdfaI6qFitOkeCWqdA9nfvgk6pxDLxSoWAEQhF7KD5c=
`protect END_PROTECTED
