`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
777LbjZgxZ1Izi7HsomnGhVRx8nyUYlO5unvgqQRNkgVIiXsvFlS9PMJGfiyt88F
s//+JJEoaiJ1HACc26f33vlZjtT1RZ1rDpYwy3xxcOHEZmArY18jVvJxiaJajHxF
L6gVXn7VAPVKiZgTktiRcWg1FXfG2A5qjeZqRu0QEq3X+a/0e8a9jffl44PWxApo
89ApYKStmZiGTvYfsvAm0DkgUmTFQRGyEJpvB09lXy9w6L9HSJl7DKt2h3FA+xSK
LgRXPFW63IvEeaN7fU5zoyMqaL0sgOxZEEupGNlwWbhHxHAF39wwiKvSCN5C5D4O
g2z0Xu5a40jGsapji1nMN/bRbvdfoTjIWSYjHnMj6Yr8gXTlXzyQ2ospvzll9Qxs
/vQhScFcBRsuRk3ktCnf7IuybXBUkiAs2pn6QLPvTpKUYhaXhvpIWonpp+l1vVaw
mVDEwxsYlLjmpLrPzlcbJ+PhuCKyGzHPPQlsTlEd5OGzL4oHWecQ0fzZOx8jhbGq
/CJteQzznw5dtHFLTKcZ+9flJRq0gpJQ5lu0CaP6BdEDhlB9hhSL6vypduRufxoR
k2GM4AOnanfk1IigCeQD/esibCEnAhSSvO9mBOZgc2DpmIrvjbFTojZmM96TuA1k
D6q6ZqzMfZNxb8QChVuiqPbTwmZC9Qb10E8D0AV8OSWfLtOuPvdM0g8d0b/kKhGv
pdaZHwujcN+o0zprRHWaySrCjg3Wji5GEwlvBjxjvGiatFtL4h782a/n3trOZh5T
gEVf7HrPP82BrVi0nxpgNGNP58rpjokCghpSOnlFnNCq933duIgEMSgeg3+eFsPZ
r0FfmQGXxvQyWiX9MNs5LnKQ+Tb9+wp7mdnlpnX39u4CWtXzGY3WOtn+cAWDGhpn
1dkuNDK+mr10rYAtkPF45oB6BtvOY3tdISNo6c+LnYEwoyn/vKEWuRyiA7U/Eosa
jeUhg+durHpl+FzoEaLih4O0LQ76DIUPR+ocwuQFNPc+Jgd2I3+/TWHrrfeafucB
C9rOHvjFdqXM3btcSb3GZWipIDmZvx4R7MJbrz09DAIoNt/ESO0NVgoE+jKqjXkI
/5prvy6TKf2KYqjijxXhKzL8CC8sy81tTsa9/PS0LitFnTghZzlRVE8BYFEECVKA
Z2ibkvH0GyEodSWrvV+5ovyj8l+n2HyLskEVIf9Xz3vmhj8ZcPtkSzWHCoOOXvT8
w4AQ5m/XQjDntlzxKZcTz9P6+VQ/dGWmTI4PRQuW67O7XdQI0jtlEL1LETvd11Yl
ZEYRlew/nMWLwZ3Z6XUHTrn+Y/TPYvMFiGrHsvGZGH3L7cykAhKb8iey1EVp5v5W
9h0oYOo6ikYckvr+1kYfNDBaWUksX/dR7vXAHvf3/y2frD28Sdt+eUMJ/BhuJiwt
+aSATjDoNO6dwZI3CUqwx1+HSP8aGixHXEN/Mx+KGV3owkMCflNlxDyuiHsrhz2D
1UkFndKHYDa/60H2RtbQgpgG+eun2EvVrQiVS0bEzwomCmCHHbwnD/tsP5uHsa82
cFruOoOlWsSrOC+KhyyQBxTHJ+ekE8JSUcNMdD7eMwGW+Gy5Vt60uLAjh8R6VxCP
lsYhCFa110zMq/Ue45P6Oml0V90K8SmVQywKADvjbkEGBnpB/0MLxTJjhOhQVyCe
NR3zg26CnAC6Z8mOZoNYf5stL8FwBe2znemTjY1HB7pBc0A0hovMtwXjo0Bmo+7a
Rh39JNyq9L+GBgKBMniIBotvPFw+8CQB09IW4feIs4Iw9hELgk3EAD/t2wBgAUvL
4Y0cnkxNsNHvo6ln1U1BQQLEfvDT/VWHobL6eWHBibQjmKKw6R96p/oD2XK4pWB1
VOzsDkObnG39NA+vgQsw+d58sL9fOHMya2q1Bswf/9pvxx24aQZEKsBmdUPXV4YR
aqGtvLl/zTB2GEOP6yxU1yLxKR2vD9XaGB2SMH9HTqvigB01Yt8RauC2LRAhCE9i
zJPh/FU5Te1zAeSTGenhQnEgEieELDLtfcatiud2TnuUvY+BvX9FKcqYZQag1XRu
3SblVcUKoeYrh84wr4k7OtxA2quIVv+LwZhak3So16MViNcg+dKGlh6Dtqvk0MCS
udaYgiEOPBm8XvTieOQEDBTdPv3050z6LTqOKhpoJAp66QXrZvA8uK3dggDWWM35
s4YWcVYBsGF4D0kRfi4Gwsh2lc6z6J4Tae0QBKeoDhjGoH/uKXpQTCuY+HumvSRa
IVyzPv/X0ghKC4Xm61y03k93Vfs7KlHTSExRO9AyK0o/Yfx0K319sN8o3EnA12Ug
958ziGTGFKnScre6Xn3H4bPuvfKNKdafiYEgGmhWvQh6rKsG2Y1LeEKz5ZHx1V1T
+7Fuidh9aH4MDAx1EJ558ledTV0ywuCcB8UCqvGLTYR8bWYvmyNvhuyO2kvbqnNI
zAPcPMG/df8SHCVBYRe5jlk0E+yKqz3tl+hMk96t9PrXlXrQgRFnRcFOUaxnx+OS
sjJz+32kjLGyXLzxl2MMgZgKIoiOYU/oLANUPy/ib/QkMstdzf5Le63A3/nKibTD
RviY878bnbu2sn29JpESmZnxt9geXzLc8EMJop12YK02K7U5+pQxufMbZgbgJvBS
2++ISqjvbBD1PvwzCdmBnsPI5t7o3o2vsvYO1ZgIvmhd2/J2Sp/YS1pbKTEjZnzt
0RviMrqyVxQL6ALZzA6uJD89C5G0q49pUo0+gzYoGGW/9mjFePlQy5z9ZtcpjwGh
CE0JUjtd1o95KWPpAxjPklekGUlj9YimsidOWMK7dm62mETNmAnjL25s50AiKu0F
8mhF8FwHReP/o0ep8q0npAMWMLah9sD7znRKL3YKWSLzOE2UHGNG9rIdREfw66cD
LmEDADBUBjZ60PmTyeuo3mN1cMoWDvwFWljYRSN+pO42JUlaeuH0MoCv7Cl+AyWm
myCRFSdC9p7cU3E8S78+ffFE90LVzU95MkiBTjvE0B4hAcjhLUc6yVX8T/cT8wza
KR0swJh1FhezbkKsuyYeszjDdUU4W4M/q4mAiGY29yI80+jZO0TChMvYYGfpBlRg
hGpvh/XTCphZB3IpDJAbgXPOEkbOncoTPZ5NuWyeAVNyO6qUWf8UaEEvA5oXGVGn
4GNTp+MOzKWVTz8BRDFlho2Xll94tb+s3aFsRznX6nyiN9C/23XTZb/e2+7bZDW7
3p6RiOPpkqDzqiGYD9n8kxZQ6D0CK3rDjm7u8O3fZkLPHIBydro73L3UwyB9HjGo
LEcMsFMdD3CdsgTi7HQEO7MpVrwjuS+h+pju2qFYWOpHKVzhamCk+/Ja3mg0nKps
mm5rSiOQ5mYUxe+iNr9DBq/Zu3P1NqRkMr7MnVF3o9Lbxee1xJjGT7C3PcJS5zuJ
ooVqXfsT1e0Gl6QkFKN1p39ZU+wXAkaRNn7pttLzDivO9WeNf81svMDCX+YtkKA6
N1btDsXnAIFc6u7euZnelXZCJLZqYlro8nJo0neXWOvWEZQhCexdpZvm6L94E6mH
vQUXquwVlYe2XfLs/YiPtCbP03M2orZpdZEc7on7HiKp5kbBtXNoIbuc32iSHXyf
BWWB8AZQR7YEfrOrFq02FeHnfnIE0wzBVeFCstK7Coa0FBxs6UL1JxVxow34Mc4w
kUxFb6z4vmH7qQjC0Kspkb1i54LTZQXubnys1c+pVZtbTu7m/rsQ0QzJPwO+r6Ak
ZaD7C3UnDCJvdSNryZEdFGSpVY/iffUeSfcob5O/KzQspIEz0phKHClG07xPqxd9
URQL67In1fa7bRNmTvk/Vtjsxu6Abh72anyk/f0gjlSRLkbtiCVMkz7yO+M/nUjT
yAP8/0z5/jLmvkwdgKiMa7GPuaHCnu8E0dBsKaOdU+8s1ITMrVj0ynmvnQMEm9Q8
KJ0l7Ssq+7XcUb+F7eONBENdP/HemEH++tVYSHMRcbiTlmLo2HLUX1fugckn+hCS
rGl7fMyEAulhU89G4QMPRrPBJMVrcmfY6W6yFA92aIQu7uHplR3UGQF2I27xXJYI
z8pKyCz7rI2DJ2KDNqmoF99V7iqhbzv5NsR73hu5S0M8+ew+kJSAdqb7zqp/5veZ
CUrPo06iQ9hW/64Y6oVC797iggXJcn6ZNWPWzPsR02PQ1bkn6UTUzjPvrxqwK+FU
EbJndW5j7UOeszGbDpM3kgi43BodUl0s2OfOX1v4Klgk9L5qgQIhRsFthHSh56GZ
8MXiSPkX4q07/UE+qUH7F9+mgXWn35LSWfSgD6gNc3EVQjCx8Wm360rGVV2hhryN
u2WABwEH7yAywNGunrn6/6JnKm7tVYAiXUsXJKXekfOF4UFpJmqIK3ssp5pZydJl
B1YMSB6trBNYYB4BbqpfEn+upba3i4Q8OtPhYY87mmG4zka8tea1l9L1xQuycgiR
xOyD4h6+W2BeXmh7DXqY71laIYx+fGZdaxnnt10e3Lde5SrNUUuWrZFA36S3qtze
xnn7aTC+zBEM1ejJ0ieGee8BO3PCn/oza/LwF38XotrL/9aWEaeF76rjIsL1P7ai
enttg3OG8ZZMc9svvgh/OlTS/V/AaeTpLMkB11CrVgJ/7wEaD8ecyk1riGqpFNqL
N1UI23pnV5Kl2hMati32Dr/oWLvpOrCNrR4YyayctTX6QQHudW7djSaMIGA+rEdM
foO9TuX55kDwusT46VJDLW8HpJYIs7JOf1iNcHp5bWdZpmYuo+zpVie3g5cEsSk1
tYtZlXRLC8ybnKYro/4FY3xUJDCwqOWUhLHWicYSmKmdCk4FJ1CE2GvRxL0kpmj3
KJqxzpCPvb72j0wsYc023Rg4xKEvMzWNK9smiX8sG113UZWOuYAddHGp0q4lw5OH
S8yfVoMzmLrLUYfymiuIH1/Yf1JxNXvUtVdkizR4SrK2Fbiyp8Vx+QnfTxbkgcm8
MN7VOhKfNXXaaJkSt2ms2UOqE0M/NSBENMsbex7cOzjls79l4FCOBfBZ5O4TvPVB
8edC71p7QAHO7sjs47f8kVgLaBpID1uMuFoDPh3btuA3v7wM5SsGG8pC7CfTpP/B
R01ATGSABQslgWa1S8Gr+FHxpykmYFxmbWcnJ9wwk37Nqhe62wSjYy/hfhwENQfG
pkem0GkiLWGQy6RI98mjGfUUd0z3TcrmqELNiGJWD1CQv+9dlCJuFmEXRvfBJHto
Ee3zJtPA0cfUgvMFJRKuHxAWeHyduYbezXNNDgAEJpNNphTqpmfgtnxce2PwCePE
wcKZN/pMUsIZLsnpITChPYrCuzHZFVriroi4NezEwP3RYEVN5GWXDb8FyT9XYVeV
7iJQ8mCGg6kMtUPagXJ2eax/MyHY444IEFnMPLv4E8OEhW1kY7Kd/RyFTd3rpzzZ
/iot4+ryX6c+280QoeYohH5UHNRtcIyALVceRL2vZ46QwACkjJJ/ApaCc1NtOK/f
enTcz6z/CYlDEr2vE3tAksvcwb5d8RNPexCvyPIWR/Damt+Il/W+B7CghHxBBYxE
TDSpAGt9+YCx1GW+6TbcVGlbmzbETAZcL+HAv85ujCQue8j+nIUqAdbon3Iuk66q
HNqlSGjfF0apBIURk+w8r8m/wMgoI70Lu/Ta6i5N4Id+628bmy80rVaaMRJEvWRn
Y+7N7GAACzoCN+He3LvjC9gqD4eVEMb0RAUYMz6YihKy2g6Au6GIy528aOZ7GD1f
4oDma4MuM7EfvhmUFXmL7HidsOX7qprOva4XXW1z10nUa01O4Dy0iaDmskGacVZb
cHt+bkH80Ha6QaL0mZzt8xvzIpvXJjaaDYFUU8O9Ku4IBp/19oDp1xBNQVHy79m3
f3eIdC+Sj6P+NIjFJRO9NLl67nwVWwOFfMyKgbi5P0IeiKO0W4Mwh3GSHR7miWrm
vOGfBnekKEXRUb+Xwu0pHrh1+bDKOEg8++11ysByfbgoMOul54vK04am/QPs9Dkq
hxjF1iASAhcI/1dYUjslqVUEeTLvu5Qv6tMm7FG7rBu8KllhWRYckGTAPR9uCCaL
K1GhHpYjm/6zR7u7IHF54dp4W4pMqo/uEj7JE2P6+jnUra4YlXyWu6CNlLMguvCG
M2LQlvHhHXrDJzXGaHa/nFg8GbHPQhomiB+l6iN7l/1kDG7Q+YQR/9AZu/8EUPsi
+NWgavIRD8xZ/aelS4dBBJ3TzniZ0ooyfmtMEe814Bwa7UrSTNSFS3/ws9xSVBDN
4YQ8cTcTLao70jIbWIFBOFE3SyzZUlvImFsvi+TOnWc4RT/AlJqq9nPLq/dmSqFI
zlub2N021EUz2drqkPi8zybQusXEx187oXpNMzNX+8pRH33vA6CR+MWbIf/cPmO1
HjNkVeKbC6rF83YRBzyKpL36emMuMYID1iPgUKahUPq4BAKn4uymXKKPyQf8JmS5
reWI+wq8v5obHTwyj0Kc5pPZkh1rp+w5u9NuQ+FPjEZdcWzDgLJaKO/PItSLiKgw
HF2sucwCX2kV7fGPtoRT2KZaI4pme6f6V2f5GSDb3hpZB6LxnOBU02A3HBl4xquG
73ij+K5ub6rYSGiW819h5Bkz3tLkkk80Ay+0RA0ub/QDkT15pht0DOEXO7+PH3RG
wes5gCVf5lAo/YEghGTLFkZLbBoIfuHd3gFnaUShjKAXyYV382y0tdTMZJuRjUg7
L97jZg2xCCcqeQUT28PhaXqv8y/juUKrQs7RgLo7ufh2uDMDN4hzUsFXzc8hVBKk
Rbljc0n124sbRncdkcY7fYIuPSld70K62ANWHUzKX+2bcCeEA/S2Kta3MXFJ+/TF
QPVthYjwVLEm0tgTweHJVvqVIdeyqCr1p81F2+dgzNjKJdGL+JZU27APvdsTOI+Q
o73q7IkLqn3yO61/H630CukyGETFZ3TNaFrznJI4+nwLYbozzZjj+rhZVxNEy89D
xUeto0OjhFoweE1A4kzQJE+Kd49uuFxozIHHnYZ8Lnb/tETS7wQH16wH7EQMm6eX
sjlLoZs90wTzzCZQqJIY9iulTr65bWBIsL6B37dT9okh9ZUiP20kW3SooqYdAPYV
1rtiI/qF/TQLg8GmsjGq3PxFsqyHU3hDk4CcjT1KU03LPrQXrJaG8BZPIs5HLLZB
jj+RMlXWPuGp+YVa/tnlMloVDxq5HblWoas9O1Ildlzq1RXK4dzxA+E7GDt8at+r
pCjJdHASUPgESAGGbpOpXyzRRG/IPHgQOD4qCaOb+okYrAh78q0BCfHe4qbW2xLs
KtLXa7dewOvt/VIIoTXORjIsrwW2MaxDG+xCoTlIlOXalPgJTtzyEZHH+7HPDDQ/
ZqiDt69qqVNMy/IutfthsijDlGSncpFcHx2V78jONOBu3kkmKJ27Q9IDeSSHyBBS
WFdwLiqKmLPLu1JFqWhJqcq7bsuLJKNroB9jwHuAQMZfCILQ4euSNTFlH3mnjNBf
RGuA4kn2gvPdMnI2a+3huCf6HmEGVAHmGmPReZmy0E0iYaMeYDAVh1h+koEAtt0E
ioqlZle40fNnDteWabqLErKN++/NsnmYYhGmbPOsa6zSjQqthTa660IQF7YdgKM9
8YImKu8TIIC6WWsTCdUghc9KvElmhShcZMJCoTabewxVS35WaIXuwFASZ6qkGaWK
Zd1LG/jEaylFXtt7nwWG2speww/NbEGYrU1J3D3oaFy4DLTGuDR5Da3uje1Q01TK
h5AEbvlEspMOF+jssVaOLf6IU8zEqgJlJm5Qmr/RTihZpCOL51pDlbin4fjcx8Ns
mIhizlPgmy9Vky8B7xTX5gLUlufpEGNsl+NKezrqJdhVyZnmY2Hgy7bn3wl2zKJq
qq3gwt+C930pGkkMPkavkSA3TzKxBluQNsM3T6oq1D1EjJagw6YbOT6L4i5mtHAi
FWh+bd/GEAZd9/4SEpPSlLFJ+2BR7sfTvK+vyKibnEr5V+4pf7junZ4dZFKQGHcA
zHoUYmbHTIENnNwVrAx5KB67Kj1H7fL+uXaixygSSODOg7EYSavEHLBAbp51DZBJ
zHmxsG8m4y+RiD8/DKKTDz3IvynRMfjZrviNZXrWDi7IMdkIf6q/StP6AFq1m30N
CiHRAEI+8qbLreeX2VBNdvnnZ7CXMg6ZFBuw/VwuMBDB0B5noSTd/9TjmLbLSsdw
LyQck+YLI09pfrbq1fOvIszrxrPYWCM1nyak0hjPppYFol/cWK936ruO64sye5lG
Pdsn5nei3tEH8Pge+b4KvMEjTQ92XwuGXbpHKMBFoeJ0sWk8Uf/HnuTYXKoIcSdW
KQa6Y17XzllUxro9BL+OJLP0imKhdO/3la1386O7wS7/V0DaEFUc7+iK+/Ux9kqV
F+ql4SMLziBf939rNtRkRZqfwuULUAS7EB8TdT4ZDQvmVvBqh9zqT+lm3YAnlWdI
PuemoFYWM6dd1RW8uI1N6xVlYXrER7yk/QRy+XFXTjeOunSGcm7W4cjLjXmXzrdF
AKeWh/e2xa3cfEbXGcuGHyrDYMOQN29vpsJtWq9aD5o05M/QbmHSFxHU1Ar6dRN2
sHPctaAk+dULJN2f8WVEXLLdMlIhtIb5DwEXpgLYnwsnLgCnfqbD8v3bZqH23aAw
QRJP9BdlzaVk6KPq02CfbsYoMWNmSNMsn0NLqTz3gwppnaJ5wU7ZLNxt9Op/2yds
bxTftsaG1t25jEL+MYLvEEoVdxH3p2VkJu15+R4rGTRGTAo5Ejgn+LEDsw0BlekI
KDdfOlzXqeHjNrxApjK0P8wA1KCv0B5vfIMnESRanIynjzTS2pRADOCpUiyT1Yec
lCpgw2e2x520cBa1pW2Xxla45ToDJr6xkWNzUW3U1/Hh6t8me/FzaWV8lG1d1hiM
g/aIsy1g9fXPrb9udxkvNb2jJBsmdguMCw4s2QaJ+bFVvOVISJEsv2jBzTkKLdXe
qytfSzG5UnYz3YUJO+yERMTAkAWo+ex0SYezkiHIysfK8lNLYADqN8tg32kdaHja
Q9ws0C4627g2zoSfBo3x1IeSngDXjBRJRfZHFZJE+lrQVg3wCYu6j8gMOAHK1JRP
I1icKz9dZf0tE8qxDL0FVzUIpwsm/feSAd/k8+Ie/7FSm4+XzOVJkDN0Yk8j6Axr
6XBym4avgre4zeX5IqjeMB099GcbnZjBlU8uUXpzDDrlGRZRyys1WJ2rm2tDqvjo
5y4PQutRkZefHlRQmzhdhOTmka9q+KjCF2CYHct2A7iYBJpjToajDhMMv8yjl43V
bzuYLYMGugbSc9cn3Twzn+Zjqd+j31QGx8lvE/JK4XZkSYFNcL2sOd9/qzhbUCYG
LxIA5MHzXEtk0jSofaa2cs69ijaPaXeXMQQVEbEyiVa8lf19MVXHSQFNz6F8z+r4
RGXpGHNbOweUxbJoKzqO/8i0Z8wvT6suYSJmOsdB1wkXPHMf1DW0sS29/J581WrE
l/kEUEQfz7WolS21tHF126xtM2Z65jfk6sRVmSuvKIO44jiMGcGCribm1KwiSjNz
sYOiqody5gdrY2FuA1h8bfrNZ2j9K0vcpRZ1xGvNcfUdaMDRfcQ7XY0TaOx4rBfe
JuhmZ4OXIR0vrkqnHHKmomdT2ldyxxwrmORb6+hCGiZmHRwe8sXazkMv1lQGaFtS
JUpjjRsqdeg7C5CyDKLxHq/kaA325J3jDKTRe2oACwUyMIANDviPnAW/6P/Z/Xtn
SU08IdFUCh26mXGtRCo6QBIZ9+7Nh7cpf5bPqLi864t2cP0NVJyb061WZAp9GSbF
pZ4nZqh8wfPmpXUb/0XYekvYkYs3BH7TwXWCrbEPuBS0EVji29y0ah5zw9I/kmm2
/fxMWMccUP1SbOII4XzdJlaLYEcDgFx6fQyhbzF1hHwOLL9Q9hhg5XIXNQE2LBbI
AiKWlrzcXCcpwjfhSFJ9gx/ZMNvFEE+qzOOceOJC6UWPO/evKTnZmEbcM9IBM09v
SzxiA2stWsHTU9sbIEG27ErH4R3VYm0RLABGYLwfuLkWep7+x6lzki3suTQK15hu
TwMQsUmZyGmKMHiUxonNRXVDmH/c/OEs0UthJhIjVi4f4Pw31miBVJFy6Zr1+CGQ
EzfnBOT4LqF+jArl/J+lGUV9g2tA9hVGHztjfnCLN1zt2z2O5ybE79OnzfejzTYY
ETIfTYOLM7iKm30PjfZZRgYQj0vMxEz6D58a6HItbcN4SCEMSCxSaCBYm0XxkGyp
TXWUBqERUDJ6/RI7jVGFMIIPmhtDVueiV3XsgAM0AGAUoMk2vkvN99roT1ecMe8/
Hqa9eO6DRjZkluuQVT8Jpsylaz0roSolOqkYZiej5hLShIjFNJ5wWTduy5YREjI2
hh8BooYmoQ9iPIUcFuIKOGQjPJQf3jk0OOdo7b3sizsuu2JaFTgoPtv8/C40PoGC
dL92CK2yt8i+bnZXzjmCJQJ13v9HOrQXY0nv9BA7O5Hnd4XVPibYXvpwYsX5qsyA
4xmtrMGzmjrEhH0pcUNaCDt8e+hbn8G2WfFVta4HD6Ofa1SzyCCoCUOc2neUh19z
0Ymt4V0iz+AnlZaTRH+wUw9lnsrwJMc42aaBsselKV5quTP6tslooI8C7GBuy6fo
KJJfxFHzT0KqO1nFMva2aLQDwWryX2lRW3SGF1Um5Lu4Zmd45ebEalZKsBXrjZFF
xayde1vt7kYZ5IVfGeUQschVv5DEH0o0+qmUzbxQo/DvYA5hjtlBse81t5FqKYo7
vl8BRZ+sipFZ6WXMKqSh2T0rXSVgD9zlPUioK0d4sO+z8v6QTn8yPrmskgWlHnO8
R1+il3HdZhR6jaM0U1h1S2dAgSzFfib99sJsEUURgByF46FWqmwy81cA7WfHVVN5
3jfGa31UuTvIMs/mm4C/04cRBnj6Jz1oslBM3Tei++mXWQ8rtY6Kiyn+ZZR4e3Xm
pH6YaIYx07C3qCIgcOBqcdCfGHXpAq4FDswEbceplQmSJGeToqs9LNbL5VZmopUl
DxWKfendWvwWO+7hlffyhCZOcKucfv+ERq+EFBBKBVpJsOCd0hi7JZzTfbsHBdOq
Dq5UrXscsE6O8vHQbnrHXIcWNoR+kt6zbUYrF+IPf0s6Kod/9MxhIozg7OsI1333
l/ZracHpmquy6Hqewy4iuQjspuzuAKBUG3U2faW1muLltbkUkDhsbkyVfOd4zUKx
EYIHrnWoXv6RzAuk4pc63ajoehCczbzl5HyMAY64j7IhzdcQe2rafYUC3ptnuEGS
NdmftXWxGJLqbbQYV9ec8j2wU7TWBfJXAHemQsmDNFmXPfWr9j/4jj+U4Gi9Gdxv
26Bc1o/pjsiwUxIl2/cjUaSdQe7Lgh+0bjpgnTK45hfKnwDNbvKci2Q+NH65xR3H
ZTdG5g29TkogiZC+unb5w69yUgNjSU7NRx6vYV4nUZT9fdTsuoD7/oCwCJ7Z+uoh
3/2K3/stsJTt/cPqwu+y+5cs4/kdDk9oTwFnNe8UabhZApDh8C2x67HdJWKG7202
dw/X2nhgwWmmddKrECXaDw40fDPhJICHukNyANr4QnhIA/Cxd/6b7R6Lmgs64YiN
FzLVr3MpzI7ZFATWAWgd2XdlRsjpkVHwhtCdH618k6jhsXL0RTDBrSWLo7xCUm7U
21FitfWSrY2BsEfeAzvQRHPbrJhrIVsOrz106xOKDUm6ywLupq8+b8sv4j75W0Bj
NYKcrSomwyupJsoLrmfx0jjwNJ+hy624pYcrIqRmCLTecy4JlcDYgtPXrbx/etrS
p5txviy/U2pw5SUf75V9bfp598uhpX2rXEYRqy0AGlWE/5nr8HXUfObScMpqAz0B
VbgcP0rwkIfk0zS18629SC/q5XckTF1P2Fai717k5Pl1HyC1qmi3ui4kPwejqb1T
eLwSP4UGBb2lnXEAe8Y0it6KcTCd0zX9B+szAF23OEEQRVdFIDph2ilCcBVVEabl
wlxDr+eyHd+Cd19CnPR1xY6jOj4/n+550VdFhi8AE7Ixv+SOl3Z+74zZRYX6M/xQ
ZvJD3PBJsqE63kZXagyawKEoDnaPITdEGcuJrPSwzmCU2e5Dreoemg/dARZcWC96
XXgTmSzNXZmmWdlVPBAg+vZKMExRUwKwVSdsrGW9Ynznh6yQfI/5UxeKiPaLhRYg
V9W+EbPdIc8aiBZtmWgN3WCv9B1wSeCN1AjCjA3/dWmEnpWAYzLu0sdnwU6zQ8fj
HIXoMkVGOafoCHAErMJc4v+7/HqRfWtzCxAmGVETw7g18rhabgKrV0GcGk4ihQaA
X7OWriRKvmR/aIh0BHIEetZ1YucWQ0c52NQeBTLWDIpbQSuv48HnpSvFwRQZC3IJ
Y3LP/F6vSyU7/V+ZraTfSPcEU4P0WXV36j4wdWcL/AOIY/nIsm7hOwztOe4spQg1
PgG2GKPVj7MECbpZq3r9qxyh6WJ5oA1EhreO3DBHMvl206z7o0KWiAR9ZMmGGzeb
iQfMeaLltwPKCJjKEFOrSaA0RoQkq14AR9w1RSVUBmkKCYxiYf7iTZsPyMgK59UV
/rinYx3fPcA7BTrTRd0Lm9seHOeT39x0dnZNI9Qd77tgerrh1USHskRpbJ38Dw3Q
dSo01KlVZjWeclfqERUPUZlGwKsTBz5hOVq/C0+bfFRmucmodbTd9EhW4COjMCfl
E5KmcIU0Pm8QObd4gVn0t82Qxa3BnllTZLJeMoqiYDKGjEwy/YY7ULjrzaYgFYVt
ZRtQJyoSCdhpdhD+RuXUpXT6JvW5F1jD7Y1yJjb1BuY+Zurk2J2borzgG0XkLuwQ
4p+RQHN2ue9e70Z7ONBBz81vEaRrMnZT3iIYMqp2LDa5iq6mKeIQTJOYbybcj2cb
bqpgPsVSf/TpOptn9lP+ukClNbJtDIolGHZu9vLWuf8U1NEgBW4kdMm/1r7RbYsY
OO/YZjtliADNlq8n/cWSssbrnAh+Ux1+mjy5cqqSeKE9RPkAQeUIF+6zniGrfk5L
zaJriKwVFrXy90UFA/LOshpnXCYjtpt71P/tDvQeGuapz1kDQlSIpp8zhBo9CwEh
PDtraF9iVCA+t0NxExFBCflhbOpPzharTclgf6EgF7Y98ld6TRZBojno4trjD4Kv
3YHsoExjT0wPdb5/WPeAJYe3mGoOh5rdiz7ohbmU2QQTi8amc6AkmSG3JRnM4gF4
jgXo6kj1UXq12R44kW8a1dmeQmNuilycRbFryJXc1CPqK8Wger4WkqTGz/BgRB2J
cuHebu+T46F4Y3lms7XqPpYma4Vxcbw6f+pbRh7vIowU15Ru7XWCCGTyu05Ska+6
mEHP5EZ0HNL7j7SdtlaS8YQTDMs32Z30RdU2hmD620tRUtK3xfO8j9p8fE1jfUYA
BqsKF8MQaR9uQhpxJ1GIs9TQenH2Q43jPXte2V/KNliDgR/NYq3R+wKELDzqfD/q
86Sxyi0kW4L0+41BTUFAcUhxdbU0Ll9mnKeJewXEBMv39KjoEffRNFPOcczG/dVc
mc1frbNKeWqhuBsKA5kieam4qHWx+4CSRJ6PqqPShww06U82K43B/j09lGsNeNlr
c5HznGosaej30LdiamT0vXWSViOS+y62zRYfUe/1wyctZhfkUvUVKuIbBXrQZryV
aBHuVZ4oU2F4cNjj1xtZ9LjsheDOpjIXLRdXWAnQcnkZ8bfVs+CcGkAejYbuJN38
bhIxd670uJITdYIA/TT9OMLCYC4yNTyJOW2wAdxMyuo8NfCE38pfnzKHPlVSSV8U
Sps7uPjgpTD2AsxdHpEEtGAiQJpYk7sAafPVXek5bAaNEBIXEU+DSdMKsajgSCL/
rK8OTgLV1W6qt7vlRJ3Ok6Fd11IwBhZ2cclW0T96OLeKcBXVv6OgdDOmGEYvylcG
bYVXsHM9IAFlMP6p2VTcmXGUBYP6/IyqlPKxUPjRCoCgWb+/sp0IAqboCjzSKR++
7O+S6yst/F9lxd/UavtxzzHDSscHdiDtUz4SiXHKXhe/dl6ubryNos3eZO7bXikU
odntv9nqtBfQrEFX2sS9yNqfbs49tCx+pzEwQPaASs7lE9PFCqSQBRwLWR8gzIy5
73Y1U1+/ex9a24O1iOqga6MtMi5kro6i4/AG3+S+STKFSplFOKvUYxwMlXsMvNjl
Hzxo4R4a5XlZBsTD+q8CL2f8BEYirO6DtJDi1JVTrATFWiS9gn/mbIKIRPFH8fFD
he998GHO6iix92b23oW5vCYVKhOY84CPa0g7rYOBHdHwByDeYkgs+hCNyvdetnve
LiA/IjnV4F2F5xnqvRRlAS3HbgoGWSLoxDn9IlE+uauAzZocD1Wh2oZz7uKwUIF7
Bhc5be9OJIXHS55P9PHN9n7e5vF0mMdmRlqQq1Ty9IHhER6gosLQ6+5Li6+bnWOD
M9NVZFmSufhvq9XAsSlKjx68tL4j5fkdjLyMR14LrjzP7vGFtHDzy6VGma9wTmWC
H9kUNN1SC0dQsiXVVGAXo47/R7W5+W6G8nWnddnneVV7RpWyL7jpqsIbXw588u2X
5vuD8tzsNCK1RRx52srexJVKtNfN+HiOPD7jP00hpl0jYL9KXGg+/t6UWvMODuT1
zzH5/RR/nPisnQXIvLAKA9AgKmF6mIFmWz9XF5r/wnnMkmeV/0KuagNYnByrpsAn
mNpQ82Q41DS/GtCmbJmTN5jaeW0JQWNkGjkv1LMylnfYU2+44S0ahmx8CLnwkvYc
t6NcYctN7IG2ZPHDLiQimA5+p6EHa4z3zR9F4V3nGtp11iBgSqqgLzjpkJpsKbd5
Qe5jxLQ6AQeziDM0CSepSjWQTyg3NCmRp6qeFKI5jdAkiIhtDAdluiaKnVhVOpK7
LDh40VKO19J82VUBM5+adr1IdUd78tCPbtjo74H0nyC/WOmADH3rvoPpLDOexGa/
hMdYriPx+oZJzyUmbqHe7E3UgIBobaY3zhvGQQYE68JzTNKqeSSscBnXPuOLAkjJ
FQftlKuNlY3L/xP7ba5tMoZtSPTppHEEvCbci2RNzs3ZOY2OY6O2Rr2+Adj8cITr
c1J+VC3Q0wdz9gbjYqzUsXOSN17ZonsC/jjKxtm30W+y7bcMNJehHtDhfCxpGstV
q1ndkmy/2io/W0nMGInT1W2xFioSTX6IP5vHXvNqlvZFyJ+OUz1hXZbxfWtg/6m6
gei21g/Mq2f8PITqwGi6xHNgYsPbrM6RDXweeHY2vOVZ3rAhzVDJ3cvGWFBVo9LT
U1mA1fbI1VL8JOP24qhhGti2CcddZLA66MPJXOosA4sEcgWOgoIajkMR6dx2pDur
Uuw3AARViecgGmdtTxYMYfAinLOcSize+NyDXkHFcm4vx7pvNG00szul5HfvQPr6
ul64W3ywNw/I9qe8hG1KpltwgsNO89z91ZsX8Z6uEELDiv507RXfPJfySmdA0Nt7
CNtMt1LWrth2P7ho/LDVnndpg5m8BMh4X+EH0rFJF3CMaLuM7yRtdO3BgUCUxm2B
iVDV0PYYjWq9HkkH2tNHYaOhLLrISqCbwwXOGKzYg0dnBIntF3jizBPfySkmOXhU
fZ/90hvJ61NVBf51ZvuooB1DJdJia6uOrxhJ2TYcRUJ6t+mxuSqgQRhGDQDMkOXS
xkzhOL+6tORUCIrvjrFc7ZeXZZjN/7GTF8G9m5Lcg5k7qWhf0oWHwVl9M9fTtfAd
26lqsjM7qwWQ7TUimquCHw616m5Ebs6hPlEZH10O6hBCMZuzYioqqXhfsx/E09iG
zTqELSD/b7B4WNxUz16rsNhvBK3lddPimPaWdprt4GfCncMhSJvwqeWVtBmWECcj
QV0fQuEfhegw9pJvTJXrkxUc30VcQL8lknDDE26zeagUrB0XZXsYtYRAUBeTwrrC
lG63SF0LC6Fwp2dBQ+nYvMbUXLBuWadK4c6fkZKfjug7kCQ05L6ZzfanGj8MCgJB
534+OxVFW1+jlgV+Vfo8CiBFLb/qQ6Zi+PQzLfrZm44Yd8smbSMS39MlqLj40flh
wruzGZbbd19dHcCayhVuSFgxNUKfcdNnuYqM+wgqoxQq7vFU57DAFnZKaCynsXEV
fzZ9jZCB7jnlf7H3y0jzNOJ6O3Bay1jZjH4ZFkE1CIo9HonKc4e2Pqeayr9jeNBJ
MGM138KkkcKm9CF7SNgHoC3hcxojRCaP7AFbfibMSfTDLEEndG9AJkHqiKRDmV27
T/lR5I/bfR5Vp76Klu8s4fS3SqTxrPboxy1E2DThXmOenHQ0V/NYAZdmSzQ0gMuV
GodE5mJfMSzMkEn9Jn66IM+H7aAePZVlA/wXKBXSA6H50cZaVOgN3oiYQtpr9xQR
oQKaRv+OAFb5rNmRpk2r0M2lgp8XexzjKS8tQQLe8qU9QMkQTMt9uAvMyLBPcmlt
rwfbiEbxoI05JsekhJrvGd376YU7tcqsGuMBklNuehLc57z+aOEpw52rdpcp2DXA
GgG2Il5slKUamd0KwS7YzK3LYdR/k/G1uubeLWz7Di2acp1PpN/On5aEH4gqIeDw
gpYRAMln9iTuT7ytrlbTkptvEz0Oj6LT6fy9bbBPET594HYNU90qusc3Arck/Q8k
J6cYO1ZwOOr+MVj7VFnOYR/jI5Mw+BKHs4QYRs1T8M23dH73vLNcf4sn93DRn1Ay
KIdj5CvYRmmWVs64+Nb1Bm/GA+tZkmCtEGauOPfThQZ8r/30IztRqMQ7HxfNCtUq
T3VPfB1s/jEHR4ZlUKf6F/y090r87vm5y2qopn1Z5tbg+lKL/mVtBtYU0Px38QVi
oNRJpISMayUrfwP3kzbTn1KEy2aYpedaIKy++UEtW+gvG0lI2n/G2401wWGBVDwj
lq8AK112y3r3C9OJ2lHLYYU8cMV6M1G+uzakFzBklVYfN2EiEnabTyR1deMbM6WD
2eRwYFGWdhlQfwCP3bj6i248t/TSgJIosDsnHxmlEBhHdol41WEOcn69098zk5o4
5nOHWOkgQtn140LvzLTIvbBHxOgWyb1laugu1dh/smvLe+RmqdZ5ZmQmmIlRRt49
+Q0gJP89vrDXk8lG8YUdbEpzqImyMDIedNw04xFcostY6N6zWU8ECGr79NoQTt3A
ycHIUvtqNEptdGYN5pxSlKadARM15kNreLNBB41Y8GC5Qdvg8ZpsU1kGGoW+QdZM
lGaH+5gtjwNc9UvwHAAXTxJ3Ap0roLGQYyc3nrH6V/+FmoBStoBZy5aEJT9LjFr4
6jYSgp2kR5MXrtSxBfud4Q9flze9hQDWuKgV+aODbzV1V5Fpf4n5bw4iqOFmw9vP
No8BSTdlqp4i9LgwgGZ32mphjtNKWN01teNQoDOkT5ZKT+s/vJ9k1/2szbEoccO7
RuKT7rxsqUnV5jyU81laGd8xB8Ls32nt99Wfi0g/rLFt1OCgXEpCoMPTKzKD1XPT
axlIaQ4D7ISPXKpGtDmbufyJPJtMVr9HJm6tAMBrts5Z+/Uyq6F7Ha4XbMkM3iK/
CloJM8C6ltRbKjjzRI+rkcMEVedGJFKBuDd+vihqSi6SwwFYb9/XpM2u3qtHBLAd
+ceC5RU8PBVZ7rAGkB/kwCePza1HyZsvM7XObom/+ODM+rBHwEUQyz6RnQMemhqI
bbSWXHKX8AQL4aqguY2cWKJseIAhQ9VwicEPIs82n5aecTvCb4OcATnAD+zyslcY
PqqiI1GdP9AI8z+mj2m4I11WBLHJU6jqACqF7mPnvDT5vu9MwaW3VGjnamiAw9G2
kZHh5KpUAZPFaSmCjwIiIDCSI+mcstQ7Fax95pY/GNG0Dun4XyTvR9+DplMCYJKG
Rk3mwviL1upDdMYL3HpF5wGwVPJDgC9idIhnhXA7iPMBW/eFgHl2lHaD/xkL6nbE
mSWVQ0khD38TzRqlCPim+k7jw+VDJeSviovvbYLLRvVcRKlutjXJ7z8No/43yCX6
GNYLHoVHBJjVq7yh0UV1rNrdDMuwH3FS3yBeA95NyaKLsVANnwZyka+/uhAlvEDI
7pfmipi5LuTxd0FbheOb9NNF2K9qb0GSa3CKLlxs9jgj23jtBQBgUb19XNeyJ8h+
HINYOxvyAsM7vr45a0eU7VZNITlyPWcDiMlz9qG/l5fwW6C2w/2zHCa9UUMUFGKp
jw6aHCcuibjCmjSBHYQfBdpRv1qIwkLr+/q1tyD19jsECkzwZGPiIhFXahS6N+7O
7rqjlaHXvm2b6KXdoLmzhQA9YT8eSW6jwgO1tC0K2D+6rqgCq6usV5TGaMPfjGbF
bS1wVt7VJ+gXlL79GOQ2G5cnoLwLUo83eq7JURHHAkrKadzFtPeU9drZUsrIlK8H
Gkh6rhWwNWQ8qE770UctSlTUWWP3m2JvfvKSCeW+KMNNddEZY2glp/2iKT3Ec632
UT15w/zOLVl+rhNFtdXEwQ2KiIWMsY+/WdbkQAzbhfa88HvmH56+xvizkkY32nei
ePJ+mi6Db9dxrh2rKbIc4mlvvYoyLsIHvBn2qwIv5GybXMQCw+QNzyMoeaFCEqqh
gyLPkKlKEuRZj2IRZBFsnzuXpvVODh5r7LkuS3utKsrWQvc1tbewWScclGSIZWkK
cITJh4f64BVJF95e94om7Ius1U7zqA8TQHSf1wG64HgO51QyBhWoInbch8qtgThC
sqsHLEfEP5ARxE8ee+uDU/Lymar24cn263ENuNUxR+z/GeIjoqiBXqofgIlC/Abs
BkUF0Q3Cs4d51mN+UyxPq1JzhYw5frySC0S9M11nlpIQl3bDKKx95in+ung5av2B
ibEsuXWfJ95xmC/wx7JM+zKMSjI1S/g0RUfdYuhQ+lFzG2ZDXvQv/QzqHVfdjekg
u33M7mSmxSbSIvk+LvE+alvYMEIfk8jEJTlIjiF4PjfzPld4R8HdJMB6uGEWYQYu
iwtlnjktlNmaXV/eehCmWFIZOsk5XvSZtnu2rXCGzZdX7+Ex1sQaXDgzS8NR39oF
J3ZE7jdswhSQfmBkjmZhNSQvH8w7Z3v33zijgzBginzi1DR/abACHgoZ27SHe4bz
7yVsE6C6I+kPGCW+g3FyOwSC8TRsO5SzcIXFGNA7Itz8tcvVJT1cJ4Wmq1l/9rK7
CNldDxoi+7A67IIiGJWBMYX29J42Vh3eAvsrGoDxwNyMUWq4YM/JZqxbb3stQST7
AvHD/w50NCLha3jBGHl2EZdYfAvZm5wGxvstLj7vdg1zO59oknmlhD9I9sGmZ5QG
jf+3td04jqoTh97yEBFj06tDd0kgisAzXITwDll1DubiU41ZWZyvbK0hQQ43aojJ
kFUKp3gJAtOf0giLLwWjLdY+zA+0A4pbDHoPtIH0zfKobPqw2gLwLBmdoXvjEfl7
hZnOYgT3g7nvttIAJ+sylkncgxeYJO8rT4lIyriuwOMsVFr6RyYoSvpWPr7fxM4M
mm+Ma4MOZ3CPigmrKRF4i06FgYWaP5URnfIlFRY5knCPSrSJtVx5nUMGlFd82JxR
BGyzq1temoq20wGlnTx6h0IRVgwYsncMNIM+Sa+MCEkm9Qvii18Y/m+9MCpE+ySb
SvgSliHAYUQiY+kD+ju2UGtvrw9W+MrV9XdDZnVyy4kXqx8wwFetgcyN3G+AKS0n
GMaK6cpfRzd1xvOxtFCDFLbME8DzMBrGcjtlGZhpWkJ4iLYrO0UYczmgwkbtLZSa
fHhkwtjhKLXhcExRCfj7jmyjGc+F2GOM8vKX8pB934O8cCAQNxkqul9dMQuF26Jz
xn5NMyAgF8IBdR0EOJDuTKOaQqIob9OuI15FDT1rjU6t1EbrNIN9/Znqb1jZSMvH
LWawNoEx3XfsPM+juJlKX98MLObAaFFdK+KbiliBGguytf8oR/286XT3IliVTgBl
BhRxTdyoVPU5NOGca7mv7/0SGpsn+5eRgCtlv/mV4IS3x8duU1xjdR79qrekn4+7
ZqjVkntOME4dXRnmu0bwU2+6KRDfbBUAxG8LlVWd+wspDSTERNmFRF6B0/eiE3Bf
l0A3sLYUyc4eXh+9ASvznPbsAklba7FYbk5yE2wJXxWnfB8HlFax5CcvSQ/9T/P2
49MIMy1Gnh69mxX/5APFjYjetaqMHYx6OX3BsVISwwlpkWxTrObg6YuzFFr97rWd
1YeLV0ZnM1pJVEK5yA7wnKfR6P5xz3ASsEVuEznUA9OIGVOc7DwL+bbIffhcdXZw
JMSabMO1FHymT0Vje5L22ox4kZJ90dEBghvGb07TxPlJzOrE7jG+3IUHL8C5svtq
rde+VGCwuKXi+AMOKtDQ0jagOMt5cOlBg5+utM5CIKB7uNFi4nWX3zyOi8hW09/S
hYb7dAXdP6S0HbMxIlcmTFqEhMxSAFUACOHQ7hvX9Bryy6Hx62jZZG2tKOEZCcCc
i8bQ59hLz/9dIv1wIydpD2x1dlOnsRfPqDeJr4tqF1YFyF6JDtXdcCGCq+m+ZN8o
3XA6R7SwdKPhPWt0q6jh+SmihGajCy1MLMvf/Aye2ikShSsniIuKLMernzg5geX1
mTk4exbeOoqyrLxaw9GabNhRQOIymxgXUHYD0z3Z0Ug/YMenOq8LT55DepbKnq/A
CKgpbhPPY7ikJHSKLMmWdcsrEuTliIjeaVehWOkzEttIXTEG6j70NIOh10K0/rsU
py78mD4fh/Q9IGjXQpBOuU5Vpls5rDMf1nafYdV6nxNSl/JPejmgyEjAIBXGLII5
b+9BCXdBzZVlWkBpBSC1Vz4jd1gPwbqCPpfnZ9Rqrxb03w50bKBXnQ4OtO0pI64y
A7lYYWovoVWZ9ziZbWr1Q1DMTOYqZ0AaMg7jZyMLES793C2ik8QsnXK9uaUgegM2
8Xkg8VcAqLWztUEaRf4VG6QAljVCTttymcliiRevgS8mtuiNqGxxtrFOTd6wj1RV
Z4iqDh55wWMzesvXWNC+WYDiGjQihmos5mVnexIeiMTkG1s8NiaFzcPOBhdbuDG/
1uQauJzIjsuM6RgdR9GEXXkJVrhS9Z/FTsLhC2hT6mpaz4FIVvYKd0yr52wkymP+
xAaOs2pII+1i8StLTjftHkQAzMpoVmTQOsZm8b4c9VChPk0G6UTflueSFoj5mzYi
tb2UUhZOHCiCNWtOXebY2fANel4Nij+TnTf//hxz+ZhBjwy3nyUWCLQQsgzQ+hzq
OwgBEmXaBp0K57yncPZm7aEOBCE61iyH+Rm6VRYXRw23kW71pwCJgSMsRZ1mnWTM
M7i0MsOmUOqwh8h9OVWCCpRM8GxtGDQ3ncc0WKzTrFq27qQmg+3HSKMuhiEZ1ElD
V0bTwv9a9dLTMoMIA0gdsv4qaJRzLgIy5lyprhaK7menNSlcWZS50BqMTijUldu9
k6FAlrSzVxo14MBfuA3FYfMipcrrDBU211qbYIv1X6IPSCztRZlG+r+06+lCuSXo
2ED0cZiDNol7oeduLJoTm0oiOKL3EvHzY9KrcR1eSbdVpLnc+zuYkTMz1GGoATG6
1mxFsR6MDXl7+hhw96wW8itsLIXn74sl7Q5DfUEsjqIjWjSQmJawQ6Leq6N0QS1n
Kc3ZjylavfIIp5Rv9aUB+Pk5jQw3SGrXbc7ViABdCGsS8AQ5Mt4k0F4pYky7FHFT
kMlw2bJ8mLbdc6gUgCPtZSthxrLQVNXhw00XNnUdtfN9PEAIm4R+9Yk9qBuQiA4U
6g2K+mm3i7zwJ8dPEhq1fmxkeGAreCZ2D9g44OHIkkR6ERpVnU+YNV240Ejp0IsO
vZgWv+P+tgF60s13mfcXoogq4sC876jS5FDzXdgayfdoNX5hMOcl+vSsC5wwWAta
h6BAB4q5JAhQoVg6M5NSMXYf0/bUC9tbseV4X0br7hKCi+hilL/LFzQ/o8ZCO19t
/NSIO7cy2NtBR6rVJFogZaP23esbS8A9iQedGc53w/UiI53dLF9v7BpZdqG3zeO0
gfpweXRbD5zJnbpoZZXaz6pwBpipnptCMAwTdhMmuP+9+VaqfKr8iBBpaCYqEJo1
4lb45Ao40gZvZMaaW4ZSzBG97EHOWp1zbNH03FabkWYnLH/JmPba+Owc4Y6qhI2m
Zf5AHvuoDS7zNwd3rbqJGXSTDUOVz45zkI7IjGc2zjZqiVZxd9pYJ/RBM8E6jEFS
UabvZ3j3zuabpAflQhLE4cHe+sFQhjGsfGYEGevFOrLOwe6Rdfhd2N3q4Eg5p7EF
yc0X22MTgHGr88nujGYCLWBkOx0KFDiCnvO9KhyeOeX4VF0VqVdwOOSLbeX9QrAz
qH6UHpDzoTbdEC+pA6/LeZQeKNZCD72w2MRZ9ogm8OKQkA4YEqCh9dehuznUnxu4
Zy+XsolXJ4DghuVRcQz1lSZ6TxwKrZRCWUumJbuYNI0p9sX57302RVpZoYrgUq/V
o9fn9xFdN0VGwm+u3xzGbFFGvkX+XNjEmDI+X0G+1Ov8p2IoVs+aZRuinvlI/4wN
pclmr9JlnYpd87qBJuyOj3X4FJoOH+dSc3pqdRH6Qz/XOX9nRxyOohVUQKAcEXf6
PsnxqUk94XrJKb04nl168FvEmY996bWUfmK8fZdSo2dPBfkF02uO54iEEZGXeNMT
1DofxzgSepu6Ls3biefc7Oj7spol0WWq4Ks67jGBMd4Gxt5M1zReOneunYteFe6d
mVKydSy2398XxSm0qmEWqOUOvwlhrc1ga2nd45Y8hVc8SldZ+8Xynqx3ZycIZy5G
a3uCp/0qjgSUQrdTmJTwfa0GNaT9dJK6VK1pFhELxwCGG0Gxa0oOIIYUT7wvxXH4
2iNYwRiLEmbc/iyZqbAWHRlsWPCS5tBSXHl34kC8WNmH9LdOrInDNEopZYN7gUtR
YZYWxe0LNBFvSbI9QZugIYB73bZMbJHBih5oX7KPz6+u3ww6TPxzNcB8szyLLr6Y
TY52IrdxQnpLcE5ljxyCJSXh534pEAN3STZCnLKV2GyYD0I6lPvFA6R0bOiZTro5
tfequ34fx6qwGmtfI6Pr1ZzxcXvHQGk6IXBABlYDdDN9fOcssrdJ8doLYl9L9bKL
B2TPlgAE07Ix30JUHo1ecufC00O+sv+8+peHh0QZXNzvlpo69LfdULvJTl8eWUV+
7qtt57Xcg+MwgL40oOH9vZd5//NU+qtOcGa/sVO0j+57DoUQ8pK2B9igk1xjCM8E
rjcEppwSOfI5Mm6wa3MO8pEop2ZRamIivcjeq/m/8o24BGZ7rfv2pSS9gmadWqI8
Yh2MFWolDFjueWE0IRYhm94QpKsOMHAibF19m3dHi+dHh+Pzg7BTYXFD1bToejR7
XZocZjYOAC03tYFf9i50bcWDtsh9dDvPNH3B1ZV/17txpi2uLfeH5haEJt9yVXct
3DKLyFe6lywB3vKb2Bf2TthWY/DEuqnU6k1Tiy0I2P2jQVnbxFJLRHCDqGHX+ZYn
oifmPo849kAfmx0eTkrfTiFutFD85weGFUF8zCiqkXKC1S28TCquA+rl4T9VQCIk
wDUiWmo8t5lGf3ukxNIFSAtW7LKBCs77LxIxWBVT+k434IJOc+/qWVOPHVmeiTY3
LDyPBnEuJYAkoIOP0IYr8GATorJS9ZqONFCdGF4oBX444NHbdKLyJqdokqUn7HTO
52wg0SqnaVxSVAoBb0eXmgjW3YpqtACQumK5sm0NZr8DII/BtLzJdUl/pIFdylur
MLUpwaOZw2LLZrvQPMCS6nRnhVdKHkqrM5FQSwMWi0UgYTPUdX7M7rOBU6210w/s
F7SD5CwurAO5kxDvfvap00bSlXiF72c664sqKIWEGW35am9D1oyRSV/7TAyJ5wkZ
ron9OtE+dMz0UyLu0odecKUgCpvFUvikjJ9b7ZR8CleDCU/czrrmntBeBBNVDRhz
05UHBUGhusM7ZuxlbcVpF0td+tz+56kMZQKOUn/XfhzeneRDzezqfAALvaxXZaSN
INRQTHpTXQDicLaBJK3+w6M44i3q2N1QUPOafvs2GCT4GMlAgM1/TXsjPHMWVgMa
plH9wxDfoPax08YdPFphTyv8HLkz4jkoOhhbAgBjLN3MvS8/Zt5LTi6jtiBkBlEl
AF1YZyxd9dn+nj+L0MsId/deS1l8QJp+xSzkgd6+q/owIYbLOK58ICjPdiAUlZpJ
92DyYUzo1g/ucnhlbLCCEjigEB3Ga/1pef8jVrWL0BmN52aZps9kpNB1lVUuPneQ
Mvpdg4TyDc7tSJncW8K/EG8t8yfhNIFYM71OoxqV8c6NuJ0MEDgKLJQCQFqbNwi+
PejPMFfO77rTURKGAJe5T/tSELG6QMq0klKwT/XZD0geeJu5yUFNyC+XzqLbVAq7
9Rl3JTHUmzhU1lqhTvw6X0CqGLenTGNKhhPMfigvCnbcce5Z/YzNbAfrZCdrjoGS
6gBfjE/nXE9YAihAntkmlLDoAwMWex0MGPgMltPcGMTtFAEJvAoW0a8tR+Kngj3h
qBFN1V2p1ZfF7NLVN+TFLfq1AFNQgOyFXqZHIBNsswos4t+JQaWPxnMrHfFz8fUa
OtSI0R88BFT6LL8rkOsjz9nqZBvQLyeBAifBhUNeTXXU6sEmdjchNT2wXODLd69J
5sFwYR/DTMqDreLP59RIs9czUyZytgtkoc/c5p6PERK3OQPsWFIqIBTQ9y7jkqw5
zL4nzbkmefxRJO4l3FVBwgpDHpQGNgM+Ry3r5+QDMv3/xDkliZST4WJDMF9/H1Jq
XFey6aF4ZkQwdM66pNk6NXpIDUp53eSKtJ1OnNo5w82nreVGQGI/zRcljd2+FHse
8AN05tHvA447ol/3GwimMqytH6ruPb1wWONn/QOnwyfN2qsLDLobnIduYnUpJ6eI
eiyzUuzDe6+cN1MiHz3RWfs+x7yGt2GGVsptO9pLTtfCwpb/Rp0+pwqWXaV99zWu
VJSPYTa19bEIMdO6kg2d/T21l7Ue1RhQ57RR3gIKC53kwLPKcHFmlZ7RKssDJjdG
cIWOsWYK6A18Hbb2vbuw+tXL4laKF5XtUAqvK20L/fnb6Fqt5fNRErBu3OJQH675
T7dgyU/+Fwe8trdFe1niKNh4pstKF/lOUev3xiRmBNa1adAIt08FEKj5hT1ZjrXM
d9GQ1NCV0rC0bGEbcfnUKcbb6j8XF9ESTHm9qGCzZY5sHS766ttWKXKjyniYs9aJ
M9z6lsEDuFPjwywWo8WIIY8z6Z6ZZNA3bSjUkoKJxIeYaXtRHDIO+G70K0WGUq/0
SvqoMpPXmR+Bi7Jg/WZ5X+tewjDuBFQ8ulmDulIQf5CfnF/X2mPXXGkEC336woEZ
FAHens4H6Yivzt0uKB48R0iy2SSmLDcLop+9zswmiv3CVaPPKWzwPOb6MuqOpT8q
U5XJoR6siygpQgMzxFlFmrVi2P8A78+sx3eBOrTvEtmIu9NrOvsMjMBjqlJP8c9K
pcFh19q5ObawWC+5KXhfQxlsVpJFUhWslG2kPO0815hEiOoBujIZFs2Dh9RfaO1Y
PXLHP1PurXc5TEavrZVM39K0Yr06lgp8zBNQftLGQDc6dRx0mf/jUt+VM0FOSr9A
CQLLsm3WlFe8Aed67QlMX2vJ1mHCd7bW7xQtGAzPS9HD64RxDCUerY4GAECgI3QA
JpjarsJK1ezqgUIOn8afr+83OMWIHljVY5j4sdgXL528tPz13MrD7rKouu2qUzbl
CZkdTmdJSZQ83RiAW6aWhTquzboHuse9kzkpcTHp9r/hTdQyGTYqffe57QZtsy8N
Isyhf3nWqobS9X3f7xqiKw3ASzOW9mZjACKJyQs0qEHt5gum8xzn0oTdOmBFIs4F
iewmy4FBI0EbsEMwI6MenubAOz7jgrWTCv/aix+A8PwECBJGhBr6IyqG2GgJFhfH
shMvs1CNUfpQf9P254vrRBB39S6qQhpE0qKP3Wj2OEUVgIaj/EhtxRysDfE3J5Gx
kLxsXXHnS//zcEw56FFxNPievdxaIeYBShbvsfGb1aFDWeFKV7t/EQ0MOrPWgOnK
+AcIg2aNc+ZfJ5OlgiQ5yYuYkjIQ8lvwEV+8WRSantNV+pP/BYMzsN/SMlm/fLMa
XWgpEuTvQlSUONm8EGw2+agGWcBkJqJ31jgzDXOpzcmeS5bdNGm1YmOQd9+LZXO2
76AzynOIvqXNSY9wMluys92sxILS5eOmrutOChiVpQffDG7wS3XW5bu37hL6WCsf
rrK/Kt04zFAJRzyykc6qs/Qu38ZKE+mXX0hA/0jf2PXe4zFqgzSb6DzzGuj+mUqR
K1QVIJiq3B7GUV2iXrEGJdjqVvrj/7Nea3quW539tcTGt8wYiCoFryycYkma9Z4v
3/NL7ZVCYX4tgaUQEYiLCM/GdE4jWP60IZpODqe5lvTBDhXzbU4wQD3wiXOE4dq2
mwgm0vuzqezOr6XCbC590J64OI5bneOCUQWZwXtgCmIhuL2ox0qMsYQVPP0yTbnk
E5cdE4pfLL/fpYi4qpQXXWvN2gKttSOXSY0PZKTIvWFNHk8xlDNwpAP5gWHUeDNe
wz4XlRGCezI3sKA0x/I/VXXhR9eBNCCjU9pSjF2eBUodLQJDQfM9QdcQA7FYx+m5
wvL3A70Vsa9lBaVnP/m9f6OAV3QVl4PIWxWiuzbGck2LFOILwpoMzeTMq3RmGzgl
rRIl5j+G8bTfEFEuU10t5iXSmouWkPu4TMdUmYfNZVOeyHYcVSeLwZjbtWEMNA3c
WzoA3yLwYU8d7apxk2Pkw3HsZ8oUcEDxC76WHZ9V6C23FuqfJWvYu58oYcYInIhc
KwBEKAFcx8w1W/POMbPDTJr5yYIsZfrbHpFWNZwRgULvYpP96yYK7c2wN1bElXPU
MH7p0W9/ORz1HSNxnNKP3CeRkLbbO8Bs11dcDtQBZxAcL031gb8u6qUntqDFpcTq
jgvxir0ExPHEq+1QOtSbS3g6axVOjzX15ISO79YxMFT/HA4J2u+SuL0N9LwoddRW
Bz71CQEUtnWCzmD0VxZePNs7kOH1aL/SiO5maacvuCnoAd4vT0w5rotzVJAaMvAt
PGBFcDiiD+7IT6U1KQG+YxhPof5dd62/YrCC3f8sFE9FquP9N91DeedQpFxSHg75
QBLLViw7bJhjnouXqzeLOrbp41PEp49pXx8AQfjBf3brKKIela//+j4DNhZUKklt
rUcKj0DV0uZ+SVaHky9xlOhB8BrH7XRAbzJmsj9prmUqFmyA4rmcDuM0aIXs3g2Y
ye+8e3A10LoACqTtqordu+YBR9GCEs/bRfH3ZJsnZemd8+OMyFeIGfMO2MbNo0u3
8Vxjc3IeKKRRp4WvdG58zTxoKoZMTQKadrg040XaIrK8E/lGmVnE2dnHT7ZT8mXi
0Q6TxEzhRB+nyP9W3Ak2gSoYUjhyINJFtr3N/n3/KLS6vAW66BkKhWChFVdJ70zg
kxfvkAIEi64CECG1D7WYFMlj/FoIwrqI9ZP8pY2J7JIT3ziPatCxibL7+byIxehd
MviZvWWMpSNcPrOOxeLkQA4KXLcfox5cvhv+AkL7pnpa/46cYPg1NunqSdwdGCEE
BTd1aC5F2+0SZAEsEZtLgTYAmmYwlVv+Gv3hIUyXzpMM4elxpPhGozUstQErgxym
ood6FxzXUtnMYr7TldTFkWTUSH7snIoArUeMWIOT2uXhrS/5Se1pgNRNoe3MAGm0
xMQui5N49/crb/T55N51dAI39QqQgN5vj2pbu8sJPBMwavMPvbvxR8efDEmQ6/Y/
k0MpJrnL1bCx1yc0YXK8RM6x3uD4at9d1MWmINyZKOwdwcJuvNWeTI4xP1STlP3x
Sx8LctIbDUEKn5o4llmHnjbwKdOm2Y/z1qGmr//VlPj+DGK0IdhBqt5j+yMUUqTW
UIKcKWHiq4Of7Z3sdy0qUqJBFEMfo1V7fHjgEcIs7u+HrL3wjtYrG4mk3cIdk9Sl
0byozRh2pF61mbS0D+Dif1an7Uk+HXX/A3L4rTc+CugPVw02VZsTm41U2JIoBFwO
HhCATbeYRmbVRZutL8mdguoATMT/BZOfaw7KWD/PmxK2RJ330u14TuWZfOl1/QpT
+mMUEHu7zv0aGIu5BEiQT6TvEZ4wDcLQShBFMbH90JQyodYILNmO1G2LY5AOCGiq
m9kNq9HDTt1+bb5f8iuLxFvr0WVMLhof1r6be/uKUuNWewqpzkatzXSenjiycQ7P
B1km8BaVYtrurEE36ugn4paI/hFXGw34scblldMZn/7bumdeLcQfMwOUN5CLMuW0
rDWvXpGa0lfZfUCqsYkCTFesE7/ibHQaV90T652CVuTYcvl1xvuNVueyWP5O7q5X
VA2arO1Hq4mVKSaYeVY1YEPhHKHsRk2anNCvsubg3xxdh9vklW4T+5s3LcFODi3J
vNOOzbhLljfli/bs4nybahbeHHxt34e3VzF65uYezMROYvVY6quSjNPQAIDn6gQ3
mDZBdmcBfPp3amZ9Yis7soCMGJBWKdVuVUu1hM19dYO1zZVAQsPJqvekz682puXB
cLr/r6IwNSjf/si802qlV6DbE23V+KIlx/aqKMyaM+QsSbDrAEmtQj6bwFn1nASH
UTtMFva0ya7QsvWwKTwg9AYq0LKTo31uKZet2IacbHcvFlPZvFBag0s7oSJAlzLk
8W20+Ia+pNakvaOxw/pD1K7yT2wqGOgJjo6+Bzkvl3PpkBpWWj9SklXGJ1b5xNGO
mqmRcwVq9lxtE+OseLzv9f6J8NRcSaz16BxDZQ14qWEULjxKWJIE9JjlQVOx7L3e
orJdf+xGg9NJrxa97BHk6ml80GkXK2yxkFKWKGZ1gTkpDIcBsNUxK6C8boUKRZ2J
apAQmDumUjtQ2JF1RAR/IqLTZ179xebN4uVAdmySHFHN2FIMOtteqKdIYAyjV+0t
wywmiaNNTlU537ewy501PN4dlTpaF0/fEVUsG8jDDZbWlz4am10EB7Z7q7W6qU3H
ZW4F6qwzyeqLMEKGubNqCND3wy23F5wGNg6dYG7LWZJfgDQjAkN2qyptq6Vp0CfV
xxGQwp0cIKxOfvJv+HU2e2M6P0eHNR9OfiyV41n3lYBZXwWFkgwoVrSgGMO2XXTA
jEe81CkWiTzuohAMv99Ahmdrp2I8ibwsQKipjcI9ny4DDph0kYrC8ZNjLeo4qsHo
WO/j5vNss/0xVBhULzZigXovFgxLZBVqvCDW9UqrMfhNY56xYe0ZKvklLkmz4myb
0crB8xBD0EMx5wTaK/Q+4jMGLi5vAtsxju23lIydweWfnCC0kUa5MjBbrwucXH51
oPPzWsyFUzi4Cj17NwOLaatP9b+vHcyINklqMD5KqN4/+t2sOOXX3iv9mZ3qhcT9
f8iL2EXQoukuVMLTsBM/gqyxqs70Umsm7UYRP2fs4HEz6PxqAS7o0tEmBGXLq2nO
XhihYgTikC65WgvG0rHJ3ztH0GYJ0yZItL2azjm/tYSf6orDOQuwpTMXG9r3yo9W
BNBOIeXKwHM6yxfNs8zkLZJiebYAFG8H1VhDlE1CXnk0Pue03tY/DDhrB/yjZvso
6NnjghKlh9pS9cZsiLSXsP9PxuG+39VCX1J1AQUcamZS37OyS8cshedPSmLLy2a0
9FzBFjX0ZML+yYyFX0sOk3T59Bv/openFkXTD4Wkmd9j0gfOUlb5BQsH2/nOw6Ib
mD78B7SlquybiF/DaE3HDgaDLs5M7IXcaZVGYVkQDqESDZJeTzZtY1oDFWhfKwaR
XDzc4lZV4YwCIQJc0e4ucJmOeBylL2sAyro8WbnVGdgtB+Kd3Zvh7j8uq/2/uszy
uI1uB1RTkxjkUaDkTVNwz6BlO1Fv5ZpeI0Cn0VCG0oHsCVKWrSQre0rVGCKz8iBN
oISwcuJ2z7Xigg8H96YWPC6/Lukxp7aQxbE8G6eslQPlfcxYE5nlYSEl1R2SRHrU
I8rFtXLwwHjkvHGazKtFy0gVNh/YNy8D/+X/EeoItw213797qPteSBEgeK22as5M
FVJEmljuoeWvp95EV56/c9EPzZg1NA5uECVHF3YKKg9swXaggRRJq7++kvS50yHi
BWmm8iq72BYxuctTbAnnZgmIsLwmpPgKrPFfOjl5XAbvXBjZ8O2DzwIpW7q3Ie90
ciLwA26PAPRz05Iz3lTV2zrFKVfj9Vxnp0m/3FCoTYSuASCPWK3ZefnFCJR4UupP
GfkexNGeSCUvD5d6ESK9VcjWzs3pnTGpi8XD3Z9kFOJ3pscMn1LyuldEVzpUAeVg
lwG10+JSTZiAsWQdC6TiC2W3g82zvjcj991g0GcQQT9j6jQPkIP2U2TDw9oWhsfM
9KcQUw7HxYls5WGk3qstJcHq/xe+WCdGRJvPzpBe+9ZQuZSLZD3JkX1U2T3OEDXn
xIX2QKJYGthc2/OzjwYFRqlKTFqRE6/bdVyvP7/h0kzLjExIR6zpqq3vTQILftZI
DwAFLxdyJc5xEETcEflFuoxv7DNffjQ0Ynih27Ww90P9+e0posF++TaebciAjYP0
U0XPR8FvSmS4zoLrlMTkVlHeNovSSGydmTmqnWZaKlzb8cu+C3Am0Gb7mUN0oRvb
oKdqxneeecJmKE65wCHFJpn/LmwWCbiZZdMzYXRh+gSfVpZ4hMaWflXpZOGlTlPk
JKXk3ZJWokOgXe44/XPrejWZ6jhMFUF7Vuow4gnLIT64LvW9mq0KjpIwZwn8R6nY
DFeZWfUKCbirwCgKyAccH5Ts9pmSup0TxQEcVLdxzgaE1NH1NYQB1PTe0VQ0eDi4
ZxxIkCT5q6IgbhwsICUT5q4Tg5h3QUtQ6tk07PMXP/kwtjlWDWrCqFQb8610KtKe
YEOscdq1UHqlXlkBMQNeecW42oB0eWHvUbtFgDsmIGbfGbtwLTZHFtYiIlX6O6Qy
vP6yYBeT9b6qScSqRB1Smdkxhp6PosSNRHTxnJe3N9fbsi3xKa7mCoI/Wnt2h1UJ
3nseQlWvFR+xDisemZsO4Ruwf7rPZO+q3DVwzdGVEFQmNEKfCJ28F21WFj4ShdTn
m7Z0Ej1d292qmvl5NQho3Vb3rF3LRaF4HfMxP7zjDzwkdvXuiaunFdDCcJXCD/4O
CDswWnzN5Xukx51dM/AUL+zcMF6RyHDr0gUk6hrOBXSE13xgT/J8jXwLZW+RC7qu
m0vLrpSre6HYccCV5teOun9/YnOPJ+0xPtRLABsWkPIhtOnOr/HHO4EP0h4LjWPH
mSuADbbzOyKBpI2OeneNwwgiBXR4fh0aB5xktVPFDLzinPrlrSCjD1idFcttFkPr
YY0rcwZW3ieF+6IgIDdDw24RRoo4ROoqbX/gJq0Bye2pQBKovllGItny+DjvtRwG
pFi/l5vwujolkoz1dL12TkhYkecZp7Xl6EvEpAZlt2RDwwFc/r6mrd4lMr/YISxF
7VfwqoLHC1Daj1budyyGpbRLiXfjwKC8qpdkp1T9QN5oK/e1eXeQrOXtpOgAx322
UMqOOxpnYCvBcqk4pUsg3tPVq5gCBOyJn+sgcfqPV+JYxqS6c51/+qXuaeZLyjam
uV+jkvfUcomfdXH0lIqrPSGgiuQauChK18F4ORQOQBMFCo1Si2oUZsle1QAwrnTx
A0WII/DoIMpjk/6jDc7OGjTG6NCh8LyIm/FjvG2li8mxvg5KvQmHLiBks4Eqd6tV
VsEMOTSGclMwHbve+7n1Owiy4WHZGD1asQP4JulDyKMGTiz7EFWtYXpHXwSFqiiM
AmBu8QOsFlJLUWdoVIHznk1P59pJzRsngx0AfsnzVR+3iSr8587Gn+AlKfGNASDO
PH+Sh4hOA/fq0B+Qif/ddbyz+kNzkZSqXxGeLxh5eX6CekCRxUiy+KBBq0rIZ35Z
67K2bu3eacZLfqPuVQiN7J7AeUIe4rbbiiNLOtGIP2XOmNoUHio0FLFzyQdlQoI0
yyKccu3anOQmVqLZQmX7U8LP2QVne9jM16Cd6n3bCozoI3CjXvKxgyOn3Zml7y4e
AmilvZ7pNoZ9mpxnOuxbQHN9P0zq3uk1dGNw71GztHdB50rw4sTes1/o0zTTfQG5
PXdsGhJRq07/SESfIUQClZszuV15cT67xgm/Dv1djarw59HyM87A0biuZF1mTVuh
AInftinESxNZZ1TFzDUqZ961c6Qj/HUBaH2308KjsckqFPH54KsE4FqrjRC1zFB7
OJ2qgW3yTEdjnDRnxKACz/X6CCyC8k6app6IptYTDTSgfZsfXgWPKzH5CN9AbEF/
X1tjrlLc7RFCPa/3ENwvMKxWlsFdcgf0cCzvajTy/lFGMPZ+kV5pZsMc34P8uk6s
JagEeClw6/g6von3JIFIEwRklvoasBBpSH7haZwdlV5GL7cZkONBduD0TVP5jKQ+
GmBEwRFOzo6UBIsyafOt5J7xRV1ZO/5l4BOfJPUM97XYu15+cRiqQemedc7d4NIt
kKnchVLQQisj0qDM6l4WQ/9zKEjnQAyJ87n8NjvBrzyVfhniQ8Q3Kgw+nZxB5Zjb
Azwl7BZY/iD1qUa4FfzdYciK8xK0Y0q22NSBq+Z3aehnOmHvv7G5N/83F3FLqL1h
gfzwQXcwbNmj5r/Q2+PIo/hyKiAHxhFkhJNtqc+EJ/ePAcqYjTlsgRWm7jvig1nf
lKWqrYfw65JGBdXvI+g9t6xRjC0ZAbB+ndaHRQsHsaR0qEhMCkRF6i2e9Lf07L2r
1mV2cuOq36a3QOH+PXve2ae+ZRwIn4bxcoB6hGzwr4DQRoOgfPkArkdJpaVK1tSE
V/vA8a2Uwex7Fbv/V4zxIZKx2JwB6S3SkuS0+POWLuK2UIHfsoV975AzXdQkwqlp
mIQhdlFLBMAFxFKrHr1ORGp1dAlFDZNqYKA4SaHi+8EhhZeUAVXQqkN8zuFONMTc
OUIPIh3cGxCAm4Df+2ZB8qSGWF1JaCza/KZLraqpW1wIuwV8PT4XxY01qo8VEFju
PNBCfi20tFKseid0dVlAKKUtu/RES6hzBJ+v4Etw6IgGk2rFEnII74tedxkPOrt5
tJISv/apJc0WUum+IOi01L0o1VwkECH1YTJlchX7WlXRDGSt1DprL05VUy9iEW2g
Z7WVvD9HLkhK1db4Jz8R7NzVIo3xezD5YNzN6sflQzUHTyM5C60AsGbVcPi+rHBR
WlSN8XNcMxWtuZkOPNk1aFfg3JZVzZZl39Gw50ZeBQTn0NBa+lcKUXWY11X7oH9c
2QBVhBgoXSFJyHS+tFAhsI0+fIPiCN1vY5lUMQoESuk2cOtr7ySfiF9pDXIO00A2
cbP+I27ySHwZW9AsFqIHgJX5TbnyApUrpk7Qk7JyOKtVEljrtuvXnVn423H3SOcw
TcMJLNfi1g7v565hqJj/3gNKcevWhXCYnA8WoRQS+rmM61c/x+gxLRTpUCAIfu4h
dVZ+0CQEpMPeN/ivxmX4JetXWGEjasxjpt+n6AslPL6rIeby3zyHDX0EFq3IgGqq
/LDgpLEvyAFdUM/fT6hkhGCAwOBgMZSRyFiShf9mwle/f9VaDmudxDD234jRMmQm
3U4eTt15suJQK08z64z9AxFf6K/ImcrvbwGaqH6YyJlFQgxwxoPJJ8AFZPUK87yx
YcIZ7zzcATu9TwDTKrUJ3DpDix52WxP6FRZiIeNwgWUVLkAloznWHoFb2eA7X6+5
0Suvxvg3uzJ62ja5bGSJwJH7lmyrxrlnr5tjfLMEQqu672tVCFhZP+E2oCV+Qvqi
n0HSrDLyG6/MIC5fd1OJfdBCaaxTW2KyI7ynodvnRw21/d0p5O2exREHQx0FrPiG
lEWm+N8uk3JYquADXwSBdul+NrKr6oS7FZBYrWYink1EsYqAcSQB44kjwSRZLoco
xBNyLbDB0AGqtHrpTnPqa7mMVqIfKGn2mWK0mR0o3DYgQxmnmzfeFM0n3lvd4m7F
xFmoPGL9tZ0nUzQytmFJGFmmH5CApA/m/zGVQhufrKMvvl9cVyKS+ZglZlD5WFqI
/KGIfSY5l/WCXt209dkdDXlufB8xQpPTHvg+lCA3K2nvOpWAdp/vR3DTqvm+EOAA
mO1LWyRcU+THweAkpSPyHDb40SDovkIfTMxhOGrE2wCco4SS63/bzSQvkgmTHQtK
YCR3MDE279jwJQP8mvXTxsbpe7HE+LHT0qSrCF1AcS7px729ArEn7lbgaDTeSfLX
TUAi9P1EeAQhqZn0EkojLjRRRGD18n5OhQUgvBiI/I/SwR+feKMa44BeJcEYYn7A
0fCVC+RXKCPbMwucQD/G8meJgqelxVhDfF88D6b3urAdApGwkoMwe5LwJ6OYNaCu
XKgDVz35scRyb3qbDP3nJoAONU2yF6CLdWg2FJ3vLDh2LxDGBdZRWgocwdh0lDkR
BZGZ7sy/voD/xrBierf6pVph4MIILjtO8i6AY8PhpG4dPc0IIzdIJcdaUk9/C1qr
7aYDn7fAajmwTfMXovnQUW6ChK0vaj35PrBbG+1d4YDK+bpI47FewECG+xq+vaCI
tY3Wh9tRiAueRjicGZND7gPoxRmKXuaxEhWzf7Z0oHfvxD50KCUqvcHwrkq2+PbC
bcPnobp0VxgMU/KEvPq4VK6oTc1uMANRvD/qMzvhr1Nk1Nky3X9Acmou6mfpHSGh
zzjjI5XT4JxrCpaEWx8EHucbjdb3nFI7l8TaOiJuc3KSOPV9aOn8krI722ZK2Y01
Y7HDbs8XCz/0f2s9E0tY8yWh4apkZnRK/NRextWDysfxt28emSTUKYM2qraxOauI
dd7asEKG1KzldicJrReW5DVbCzayToUv3QUSM3imHtTL3FK+9eB77Z5JSsVJQfyH
8GmBIn5THunI2j+orbV+WojAcuSoze0OBnVX+vywdiZTAEcGZj/uPkQ4en11kp0V
b5YfOEfP7eHuRWn00kVdmgqdACIHwOfjM1VTaALZQvrCL2Mqds4ll9wb6PcegVQz
fv5OIQkGFvmY5tHWe4C887TWB3+xikhaDHodTwOWbgHdDNo0fHiriakeDGyin7HU
Kl8F8Ssc+Ckagn+NipULYn/noFzFY7vZc4seSVRC0kb3yX4IVQy6ylBK+gOSMg80
W3h8WgdvTeFT1ifUCz0XuRIlZ5jNlYDGO+wxxPj0RuSle9gmTHyMMXe6ch7sDZbr
xY67aI2w1q2/S2gUPgXzCKIAa5eNPtt2O74aPwn9PFBoB9B2l/cg8wxxh4TFjDqk
qtETpK+XQ9zNt/12EuMTqvVcCfoUMsXohaj5lv8DfGe3hJWg9cj/xnCy3YBEk0PA
km35f3ZaNKkwgiMxZbMG1/dpd6ygiNJscHM4euAuCUDkIMi7U93Q5cjv75zb+6ia
0rlm9PjKAQ4OiJTnMIoNLs37v8e/cb0oLUf1UOrhypuYJ6jQhJul4fqs0X0QFM6B
+N8bmiOKpSKnYSnJ1uWwONT17FkDBi12Kt+vNKtkbe2aaJ+1OY/1FDy2c/XbQ1Ui
/5VK60L7UXqYH9P8INEeU3acfbK+59EKRBFuwOr3z86dh+/w/ZSNOxR7jqVaPlVT
mQx6t9Nyc4YRzBXTfU2xqCA+QJzJMKX7dIYnBUfAf5pWbw42aJT2ZVeniCpxLNuo
XLAf5/doRCkhrFcleK+JS8GTyXK9yohhr16SFUv91lgAVc8jhMl8EN1dR2rhJiX3
WmhkEKZgA2xJBxMtQPKTkcVKOYusbQ1YogPT4Q5mt7J8UNQCTqUZjMiE5FH72u6f
u3fvTIXAhwWg6zrTeK9Yz6jw27j7AJ+41DpzuSuE2J4Y/xAR/Sgaid1TnstyNv3a
Xh+eclvvXp6PzgJ3lOJVaW2FRS9RHSluBAhauFi0FhaXz2WqljKO07JrcA1BNz/q
8cK8FE3BISGMhObo1UiA4s+/TpSuWFIOFDdTyGph3CgxzB2pQSGTWShmh6oO6qcI
YjV7Mxx+3ogVPjreZ09zoqhjzGAUA9G77CNajAHZjWUIv72tbPJmhLZQPJ9MDlwU
K/seDdziz5tx6mCgTZepeGTWeZMWgsBMPTlBpXlPu+7ZdXOiJUIrXxKnyIrMchiV
152WwB7ENT9Ciipgx53r3UMa8VFNpopIbCWfj+ezDOqMsNQ6688+0Ruqy6YrOq6Q
PnqmEs7cDlC8x+EIhC88IYJrweWOg7jiKBNXVZanmRfvLHHOvqGuD1sekzUa9/J+
T/VyWlKfBxd2OwM5FWgiinOImtArfefabA6WAu3aLREkwbhNfO6SXI7T5kS0Gmjh
PRtQo1sU1Q9U5ivpW6RHFuUWN3WMbySjzahSGA/fTfPt2jJBQ/PNf5MaVQ9DQd/z
vr9TTNq5yA6+pnhizqScKwJasuI0/u/QwQZvm6dptl6nBo8be05QwiFXzdvJO9tj
lfY1f7gFtaVfnC7xgtpyvcqEbFeIt8P8Ib4BmWPGxK76Punnr9k2vTwnAsucH73o
OJq4ymDD3PXApYbBa6f/LNWr5JTO7JLsgr8dQt7MAi9fUwv/WIWy1D9MxgBgPEgQ
0yh7OmKEOKyCWJY1PRPpAghxTtk/rTwH7v17xYfj0RbDzhXk4RyFV2GlXy6M2ax/
NjNP842q8ZCySgLHcfaQj6r5+9lb3+e2m3RHbprT+TTMiS+UFNlPzHa+jwj62TeO
i5ZaJ0cdeygspHLWbJ+GrCTiTLS/672t+PYH2qUdSXnsNTUpql9JXvKZYDAokQ5b
iBtmwkQ9wT2caNUr32ayyiyM4heJXet+Cf2VPqkr5S6X1vpKSJBi70EasSVm6TcA
LgPnTFEBH5UltcCjf7IvXVbc8Pi/0Wwienf3z7qSI1FUqZUkhEtJuzfB1hCfO+HX
W6Kg93fL3MCaxxIcXyzTlEoobLnQirj8nDTAQ3bvlAmUfrvMndjzBdK7Fd3zPRN1
IiNBKpX6b5vcHtfcHiiv6CJEwM0IJ9Ni26D6VruQ6dUkGPC954RXKJhCk+mN1onL
25qkVWIgK3PaQ4Fmx+ke/yNNiThoOyyQZgbeVPwaGI+LDtnVtQYqtDN6C0f7H6vg
mbCSHTyv6VDPIa/kLI3dDih8dPnctkGVbQQgw1TIeShQLShzw7OrIoTpJsWLeyxu
K2/WXSjad1s2G8mkdI9I5UG6e+LEuWNm6hWKjNtLtEHnW0YdliCuR2huTA56wmhh
sNRWf87t/R/wKhI8hNSMntoHT22TQ/2OQ/VvkjfO51kLO0x6SeEHJFIjsqR3eHRk
fa4u8xEmm5ZGaJITjBmmI5VRbRe/xgNHKFJeecy/ZYsOjfd6CMNhl/OGiBnxoPWN
xPYW1PcU74tLUU27PSpZh1MaWDuy6qVo6Xr8Z0BO5WOJMFyivnwfB7ejPxElskRJ
SHRMlUZuIR7py14DyLuUBPTbAtchoCkywS8Whp38IJQZYRgU2561TyFmS3r/Bt+7
AwJjMGdCaI8tvMN8vlUTY4gF3zYzodXA/2eHjSQPrpfhMNJ2wbjTa0MKrXFXgBWA
3hk7OYDJDxosk3GCFeQSbLLNJRqpKomOWVsuFFKfnaV1HIAQBwROOI80l5MEwBI0
PeHrUQwiu1X9UC20bqH0BUM+HRqR56fTqzzUcLoBHQSw7OJG3/Kbj8sDUGcNYUrB
QcQ7FwkaVK6UsttN5H/LhBj33Ltv93MaMOel87wDPOAKd50IP9AUr25cq6JS8cm1
LedVb4HG7zcK0UAo12nH5GF+Ahd7Biz9diR5QiLF5im31/2PcvyFrbdVHU/J6+2g
xEAzBXdVYgZ1e4HFgjVP1g3UT7STUAkCDOmygIK1y3w7rRaG0yHPxgQ74q2owQ+W
fnN1Y9V0WrP+sjMrWqHXSKhFvoNui5BrkR0X+sNvUssz59fOwnUVTuFxFr1+XIPD
DE2KfYAWmAVUJ5wK9rKi7jxIpgZV2X5r6EMeE4Z8GbTy/FnOwPWKhk9yT/YrpNi/
lpCjTcBGHCsWjkka4vIbin48zfWT1EgLZ4OimgkEP1wkOkl1Ft1BqSf7NhZoryTu
nuJ0ZYYPxpWZhuCMuyxmxM6i1hxI6xAf8j4G//UqbFnTMrOy9gtmwp5P0wGaZ0dv
TfCsbkwmYSuEojWK96dx6rt7pM9a3fWd652TJ0V/g/Wrcqf1hmeOPQTn9qSfTdzc
fHmK6hjfsPl3MKVSUmsqSu67S+Jeo93LODrN2hVfsBm9biThHVd8tROuGDdRrdH8
y/ZSjQaSbx4rclZas2hdbdS3Gv/wIDg1mcUr7XK97aMbhEhcp0pLIv+zrq260FGm
PpyJRE0nE6+CMTKM+jTrWpxRll2mOFdQdMpsNvQA36OrHj18tAxhD51SQVxMCsvn
XPexRhbET6fVqj0wSW1yww4XP2bEgUW3i4JJQnRZWzHFI4vSVIZOtJZKj/6swWo1
drg143fcpu8vELXHj8pWIcfzh2LPR+aXZpdFsa+GrJqqc/rduKweFVEGrVWJfPGy
5suYbs2AaEfC0AChRnmdwPa9ocLixKPTioi7pFRVhhnp0/PK91ZJhxvddsjakCns
gZe4FLhhKn8LVTudIl0ejcPl22gwmyqauNC/PQwyBPj7ortk78L0x0LemNYheIeN
AuZYs4VII0FlBGHdp1MRuCM4/kTEporKq0YjUAW6VikjcA26elIz2XTKpSGb0s9Z
o/ZLKH3XnjgMXInIFvuIhzKgXH5rFBXCzFmWeGdeHEVHT41zcJStwbxbIAr2Bmuh
R6uV9HjuE8+I+RLTh25/EXecPKt0y2H5VTYWdo4zhP0zMOqgRfMTVSeBwpQltuss
aw2d0OmAzUrRcNxF/HHasVoQNEPTi/insBVZCwc6uB/m0jqLKSFJvF8kWI4dnaQ3
djzxPZ7vGcduQAAhbnrQZM5LU9YXPdBTId+U+RGD0R9zOFUJwZ0g2ohYclzgu1gf
F96AeOuqxIFDu0+tX/IP3U7JdTd9gHv0DlXNrAxL3rVc1h6Q1RySrJbN1z2hWA7s
b3swhhIbcpoSSEG15rn4xsLu+4TkYtn8oyNTttBKFL7JDidOgQW1XFAlmm+yxnGE
P1LjqQgxKtDR7fpxQtwTdyhPbNB+uYIjk793thLoMqQYz+ifzNW9B4QU1MMgK8vn
UydWAHnsijH1t3oxsSUtRA2bBtx7lroUxnVmNsvKtPgNnSistE9ZXhgTyVFZkcje
tKSkpNDnF5v4ufdokeV2VtshSJSsTTwmsDycQ7M7p/bKURTBd8D/enT64FxDhRYl
EIgky00o+EdlutOATuOyLvg03NAWLW/wBGQHpM2yURfjlpOV44EOEqhnoULYDONd
LovreQYtfbNQj3/7mMWbypnV2X4YT7EkT4fsZC2jF8o6NjhTzTUovfJNQjoAwtke
baA0AscLU99acUJE6teLyU30G7o9SEeihcTM+v2bjnGdmFDANmF/V5ZRkL9+BElt
/bq7DFkP03xVMkJcRc+PAl/z3M4bo6FhmYjFIaGoGuX/9g7ys1LmLCOTKbG0h85i
HRRpppizsaR8XC2Xb8J/irMaHjn7YJdJrbqLJz0383kIfuspnddkVTpMVZ5ayZ6e
2aHP/5yrNxkq1yN9czeBumHKREG9BaMGf7cpMx3RVKFHeOyFPA2jZEh48c+6zZ1K
yuJ1RSEsV1TvDW8yCjUcmq4z7tXiewUpXUUY91n3wDjTNlJwysJwEROKk9mwOVpZ
l4gUkXGHxE1Kxn7oTyASnXJPvUT6Mgc3maN+1cauRHHNzeBklR0d1Tk3yeZOBBEv
xdi4moEhYNmHXueWI9ebrhLWA+TaU2tjgQnwMpReGtuxAkTUYjXFqQa8ygg5ruCW
bk7FRaKK/wLimjeO/eN9NFJHz4m4CFapwIVVtHHTsBk2HsE961ix5NGdHmuix2H0
dNnQcWgIxGPkLNhl9166oEt1+y1BOZ3glqCyltHd42kxiock0AA+RTJjqujS+pUe
Ci+mHwo3cOW+Vh7/Y7jhR5NsG4rld+OYz9TkrsargxknKTP/8lW6tyt81IR4UHt/
t39ePTCtVa3Y+wjl3CYq9DRh/siS9+azTOGBJ5HgKQbLkvq9qku2WEGiPSbYqKCe
z5NRO8gm84bBtblgOZnw17IruurVelKYdK3ZA7NtmCGH6HNxqE0o0wUtrRg9mDcn
cYS4mjz/eiiB1VZvg7XRyLtz3dKbnG4YRRMO3EzCa6Ptia8OkViu6mwY0b88lKqq
k1FnRLk2md4ez/7qiHWmcpylZpLb2JVl/62scMMJuf8FWzipi68WUKxAR2XFEkHJ
yRzydbZMYt6PCYZ+bs9hjr3r3b68xTnzK2be9BtHip379ASK5WTilxffm8wu5XNy
kb/JkVv3SXwwdiY4nCmKFRMONozU7ceJpJvEsuy6QHHJKG+9bCfCIjchQzFJFmn3
Avtq3jPpbeoZ1EJhk4waj9z3KeFdOhbgW0/SOQribTGmXsgia6egj6WPrBJJAi2+
rau6gt5HjG155B4uMuzX7WVOIY8bkW0kwhKw/CllJxaQ6EuoIBd/ImEvifCJf7CZ
6AO869C2r1cmiNLyKzQCqrwvb5zypc8y3WnFv7Xf9VDjXEEUa3e5KALzJ7iBRTZL
g1uppwFeK2aHjpqKdVxgz9Ldh5XwSnc9G1rx4Tp8IrfULKLM4RfcGvnh9qXVw8RK
bfkuh/Tc1iw31H1edMWJTUrfRDjnbkd66Np9xZ930hXcneZb5GIbExGxNK6yVSBO
aG4RPrKtWQRVKseXYT2NrLTklORDQm2IjSoQU82xkaNJajLcw2sV2swCFAzsKV4q
U/l/G7prEqA470gkoT9+/2CWRFKfQEBPbt/VSw3m166EgAVax0/etZw/hquJOV7b
Y46Ehr+T6jZsE8uIPE0P0rYNsLT4PPNZ7fiZc7rePAB8eXMdNAd+9D6EQaD4NwGR
qk7+4PmZ2mXescJw0+WGhY9EUeAUmSySOkG0jUebMLrMRDo8e7r9F/42wU2h1syW
IrihGVWn/HnYpOXc5NDjGsahwuUCf0Tjelmq9fV9pzHX8I4V3dzkCygF6OM6kEz9
+snXDuY3dImRE9VpQ8k7yVGrOvgXhcv5zTrtnWflXNJvmC+IdOoAKT+W5EvhAUID
gigauT9UiXDdDKPH68F20KCwYLBNw3kX4vuZ7SDd6XSxB/Jvc2rx4a7Ki2AheQwV
5KnzlNoHUyY+t/3UsR10cMoF25OMj+G3Y8zEu4VyeTWTUUwqOit+7LxxyFd7vZt+
N03u56V8d74WRyF6PtDxeWjWcH/ngEnqDozyrjofhmrLqAVEWKz648pCpzWOjZ2F
gVTrjFXLZCB5DnzMHlDo+/f3tuw3FeU/8wMBTTjSzgdFZ/YIyE8kTbXHLkjLmM3P
cyPVqHOCZBTfrD7IVDwWdGal5QMKmJGOfSdu2s74Njgvf9msWP0yH4kZjBv1JX3G
mQwJQIfKQabimWt+adPWw9M7GzsZezhujmWE+91KnpzwRmvjZWHGcSlalGyuoIi+
OrDnpfSi8zvOe704KNq9uRHwNhFWO5+SnNUkq97n3KbC/dUeHCzWOhx1SYVYGFRG
bYfxKkQUhYbjxVvEIKoelMec5VfMMvoLmzniGCLVMFACuXEhTCKNRwA9IaLP8gIq
MWMZkD05GdEE9DtIU2fxdWjaeSl0UN6bE4cs56B7KEZm1uJ73VjGko4NWP+WvIOo
MMlmcruxbl0d8FsNP9L5BVrrXUmxBqVem2AViguq4Cc0DNITTidVJ4MYERpsbSlO
ucDtDNTAWB4WoUUzmEsoDCxyqet8WOs4rVyadFnGWzjiV7+mQ1nSFEqOFP37oXB5
tYshLwaynscUVlcHc/lhz+iBqCIKPVONVxMAdfxSTug392xtcn9ZjD3ae0n58Ke1
f7APTVbCrxinaXOxQBMWnVpyIokbTMVld3d42ZG86MM2oand6EOe4jVjQ2ecAnME
EvSFhsr8UK6dcdQBXf9BISXremlJeomRwxLyl1tIS0A+QNCYvCo5tSlrwjMjASPh
dXlkjDbsRGnPJ6QyMwDaamqdlHHVFQua4OH/ZqUEkVpOj3wt9vwZWa1aGkA5xF9k
X42+6Z6bWdvp6zb9ZuWi9x6h6KJrc4KavL8rgsuTNLv22p/QgRty2OvJHZay96LR
xZ/H7R6kt2wiRQYuZ3KO4jZEShdvMquxSy9/eUJBFskD2tWb9AY6z0Zicln4gPeg
nZjm7+LNkf4EGY1uFDDOiRPlLbK5Uww2pedabmmAE3KRpphKpmySI0CYExbTRqU+
CQ3nvD3lhmq6eav2GltIAnW6C9nlgPOQrNLFa/qANQCfXCAuZzRTIxeySUyIbus/
94XjlNQpd3gLP5Ni8XJ9vMRDcB6BShjsf/7V2yJgO4HpubTsgll7JONC1bo4A+iz
WQu3eKhW8UlNkuOZHa46geOcpO1rOirl3scwTMESFb1kPLEG2Pia3dOennndzmez
/Rjk5tb+ysXZi6JBJbfwXfM1LkGfhRu2Divsh8eioC96ljd7Tb73ouz+98mGYg4U
Xuhcv0Zw04A9OUPYu/bEjCKXF62kAVNNcvk4FKJcYenkjIsehEBUb3PGsEWhjLoq
ol6A84wDoq8MmLO2UZwLJCK/ZkOhRpmBo1spxRDCHmPA/IZgNeBbg8LYW5xkpXnL
LIpYKXyKs+Wcd0U6blvSFwyC8CZAkJdmaOiKQpu/x4gOySrnHaccuxqadWLnHhAR
H+soV550xgvC/6O66s20+9UOB4wyYTS3lUnj2I3i1DyXsyVqoMvx8SExo18uQPB+
waU5p73tNKeZV0z7wGlI0nfGva9jirR0wdbLt3dgsPehLjb3Qx5UB7aOMgQYhCtd
InWg5xR/K694OOXo620gaQ8KlRJYsKewKtNjA49qvw9TN4yFENIknJk6LPQfADVh
UEPKBxEQCEnV86IPab/UigUH2ZdLuEgvM+u8QHxulo4OaftXGT/AHVAV8pJ7p4x/
FybNhNprnySMtjvcISmYJbhYOZ6sb3D1w/A4PC2G/JAj32g+hFT7w967SSnA0EaK
7KnDO/frcDFqV2iPBR0eS6F6Fm5cEgxwPA7kQDJVaozoNPd4KHPXbsGfIhjsEHz5
iOwQ/3ZKcfRNCHSfVIrEWtsJ3xt284Ycsye4egEktw1bRRcNRzrIfKFGJ8fBT7ov
m4Y4WWLNT3WLpQL8/bDIKm7SmeBWU/FKpT4efudI19JktcYMma6m45qiLC9hxUnz
DP4uhW6sXQ/ZGEveTh+VVbN4SCq4kczQZQFW6kK9ckVF+mZSaEHdLiLSStgjl+MH
H7rctlXTGqsRnMiAgrBCw0owU1siyBBjZOvMyMW4tBjph0wYWMzguTbetyyPg5Fo
VEPNKkbaNAVAvRmDOkMb/SeMqiiU+cBGUuTVVjiZWAAiG5e/X8tA0wVzMhZ1NTrv
3RGKLtV89echicuzek585Dyqxiey7YcN62RbHHTfkS1xDRpSNBmYukOhOXcSldkO
YYULYa5UrQQ4ARqpgplUtFSblca2h0aSsQRhsrB0hw1nWH6zNinCsLjypmf3gchl
aMu4SYwjTowrShijgwrd5eCCXyNvHbs/9QxpyQF+ezqaDIzfQzP6AzqJWm7TbCmS
j/3LPTbVD/tk8xtuCOkplv5yAEWaAJWICkWsYffJqWa9iYU6JviKAyjL+2kHPs6+
pgfC8IDa8uV3iGJd2cl//EdivzCbkLsn+CtoNNsglhWAOz8gQILOtqU/Wfw7LE8X
JS8zq6f5vaPtMVR4SCDCbGMFTHQ5J52c5E/IkckR5LBUvapmz4okojGOEyjlsaRn
GYSmrIFhISoKVHaJ3DsBP8ZPmG7twTEU3EIxdLZhnvScEEk0ClIHFzj/mO3K7WJq
iX9CSrNBVuHYiYTxu7ka43I61ulBonTCw9GgniGdfAcwtaBQGOuzMkMgznufuMeI
tKf/5OhZkeMy7DTN0r4VcVfHfbO1/lVuZqFWr2CVALoBToXkQ04foYkfbfHjqwU/
ytTyWN6Qa+f0iOHxND1yDzDd8SNB1F/FqCS6pwGohfCFI4IX2pcsWh7phStMr2+j
EZ7tNqPPzrJ+bNh7UonFv/9rSbNCs4mWQiGQeFctVizJjMJVTtxgkjcA/PGfeWUs
/y5yhElnT9kFyEXEo4USIg52kIG16GnNfozR8bA+JjXTv9I3buUEYRBRl0+zWDpx
ZvFY9gDdWc9gwvOie12VvCSAB2eMk3yI25q83g3WyJcnFwFnBonYXOvLnPZtufjL
I9kDe48SE3nz0K227hinYLW4KYRKQ7dp3aM4WNFEJSosDXVMF+joYwpJRL48ZLv1
kW1k3yUqZVB2yvX9Emlbkm4ybTagAIYuqrx3K2DCN8WwOJqRAEZTGFnDZC3IK6n1
4gYN1mN8qh7n6s5PARrAo4+oKrJyCKe40N8yGQ8XxYxN0JeQD9R9LPJYRNdgK+FM
I4M3JLkwtQ18Vuq2nStWjPAnS5Uux1Xh//LVEJedQL1nPbiU8caCEDMDCu4Zr8Tc
bJymkpI/LiTLikQGWs66acWwb/MiSkYoFceYXM0T4wuvdeI8Z3/IKPZj3CHDd7Af
itO/3d1S+CRjfFbAZfXAaLSpGq8TkS9EaqrIfoDLS0KSVwgYKj+r6JQvUQN+5Kk1
+Pd4/9bcUNbULpq6vly7fuF6jIsgQbPLyOK15pV6tBSB+tuosljCowRVH0Wmmznj
OUFr3WWP9ucFIcKzV2G5XwLsbkhao03PxBXgnPVXU3QlgmJwadOJx0pUxxb5rMP2
eWzsSp9ItFa2fouFvqfSbJj2+8l3OhKZXRbvAToHbx896n7vd94y9SZ3Fb44oMsX
VxZe6FTkUIGgZR6eQk8sKbR56zXm969ACzNUlBHoQPNRCnwbsVm9b5ffFSReqf0f
P2nYMZAZlUrAul3SQoM1XeeUTFBWP0lSnuZZPH1bdNdBm6cMTHrmMt7WRuAhmkWW
ivDLXGlEhMA0ZY+lWiU8/Qy0jLBHT8A+2Rrn2ql/8AmsHjlivgN9YUIEi2vpFVuD
+W+PSRPSsYxHLy7IDbJA4RWFRDDytGtYwUQSXyoUc/zkQNUIJtZ0w29pUhfg3NBp
mfiBTqYfnn8UqaFlWcHfxQCCFWGVQ9VWNNmuVQXpsJJAjZ4yT37J6u9CuhBqzGq0
OhvQC0sKcvL+96Q5HxYTe9cb9hh6LKTulhCJIdfHL6e6VJ67LhIB0SdZhRnyyF+0
xcWlbdA/vQpqmHRgB0sKBdSQx9Wklg6pAJvJg02pI6ymMEKQuNhewgJBbkxYshE3
r+myC8qE64Up94Kjqxh734BWBa8PNCK1urVa2YDYmsAnichYrVP5gxinShOqxw1q
IbR+Tbfjmt9AMEYEMgLvRZY3pb6VbR3fb7mqjsFJ1LFE9PnvQ03PBrT26R5itV7e
KAtKDRBJaamVkXNKtF3fUjz9dfOA1D28+LQCrCYb/dJ56n7mWph/GbV2DazL+Mex
RtXoB6fmRFpB2ucKxFlMwwDc+Q6d8yaAk3yapsu0Zv2lY0dDHF1oaDoLBbcFVG4T
vTC46bmeGJkS9dDaWVOldOYSHQ93EdpM7rEcvr0AxXdiSSCa5g2UtPaHTheHpgQr
qgBfZGr20fz9Orvc7D0V9rBk+b0fYJTCGSkkzH+gy+qhumjyO18iZ0Ty6wYGKT/P
E6SomlbQvcJWvuH26iedJlPsV5rzoRTmZQnff0eo5OViToYJnOPwLDF8g0USMrPO
FevmrQ9PfIuipYnnu0AphKkPJE5xwwL8j1i6g/Wa7uTl8CxaGK1J3eNtOBfxBM4A
GYShnYY6kZZshdSQLq853L0aRCZjp3IueCdiwHxiWtNsrfmgfKqkTCQAgLvOBUVO
TGta1QQjAHZ6gUw1HJ/n/UXNpPaK2hCVoS/10rAFf6QvnXMGihisvXpCiDg/VZOa
M8VHGCAvQ3kg+SJCbDrSPJ5+NuIyeTDGkKcZJZP84CxvB4a07QRWhPM/JytB/7Ou
grnGsAFAP/3aLrlMP6tzj7m4tdLL+RUJqjr20B+D2LJRtK2LOL1mbzFSON0+me9c
nQllKoAFvrFpOtFedv5v1CVmCOxE5RjzYukTE5XZocy3fYkSfPbm7yubFx/9QDkX
cTwrjUe3xzVTvHE358eMvCAiAKBYS7otBAFnG2by3sCL5NxL3DYMKbG0gzfZ3HJk
+/Mdwg2rguVY6CzJ1bMmMj0imjvMbSgIO7skjOjRVVkOohfzrQ+iYMErK1fi4BSc
C5DhKgmpZb25G9ePpkMCZXBUTczD3GWmzGuJ7xHGdbo3GcUvkIBse1Gok2PGLJyg
ByWDsgmVXVvCS3J36D2POtFZOBZsTqEzjnoljj/j/X02BO+nqWfCqaPBKCgAwsLW
ayLg3XIdBW+o1+4Bus2EADwo4yOo+keXBkjlAamY+JFbe9a7UuVVOHdx/dMYBQh6
vmFczReUEUUs9ktkxMgjNGGtge55QSGNXegfE2fj1cFHRySpONE7Pxnjna2dM7lH
2g9j4jepeytRV+AOJaeO/mGUH9OVFFNnwt2wZRGlSVyfzb8daABg5D2ySGOrbZ8a
DJLnJcMGZMOWFplbGnvH/iikEBV1S7EmYnHrESohmxk4AU609j8sosXMx4HNqVMU
U7y588Sr0WJiwywonuI1prEQN8se+c2jKhMUgnBF7YVQrMwVJ6sKrNr5O76sFyoV
ZC7Sr8VI/sTlIwtaYij0JGwBrPjglaEIaD3yjyby3uNxUZZuHg2bXsN+P22lVza3
S27GSeY1j0Sv7Mz91vTAvC4df21ZE4eFTxYhy1Ix+vnMgvaXlZZoMYzXHTvcEAew
L09xLjMUHdT75FT4HtVBHhk5xQDcJLrDKlS6z/uZDEx/bGn+XCHWNiWklyk5jL41
dFWyhRRZJGFj/22KNHv1QnbkYB2SQF5x1KzgBMRsYhFHp9wEtwoATu2pLKo34P+X
mVYuJ9WL0kn1eZJgKNmSnRtW44AFYEdBaOa/GpHzP35bCmNp9cNctXC6WLXuTfvv
zFXL1fgaH48li5fyQnIHklIUR/pwB2jik9Mu6pqonAqJ36SVwMdW17Xi5plzMA0b
IGN6KkSdHVgOih7evLlYhkYbNxmqIRPRhelF4bvHnvp/HOjYquGrK/4xD/ZJ8jak
Ht1QdUq3F5MXSPA45XFbRicCL+T4hTbzdCRJHIfMbza9gfQx64zwvPqfELejj0gO
PwocrRVbwWFhrkCmKbYF0+6Bh9cP8lTZRJKsnlR9LXaa/FSSeY+bit0cAIY87roy
Du2PJTeaKV0HzLjd/lYs1I9NsB4K6/OgnHmg4wk+2sdngjwjYKU54ifqGBDVgoqH
DL+r6F8s9GDvrTZrXM7WMyVNf6g65z5ugqyMHwBLhqDHQ3F3AZ/4uS/FPiLeaNgq
OejxSjOIUffrwc7GsX1zFkrJapz6K7viD9NVrvE3OqTKl5rO5c/4siXsXQK1lXXn
gCIsrPlDxApQfBTQM2JWvvPFiZMvmyQSDT+MKBH0i0oEunhUQtJQ40tEYr64CBVz
Be0m5XoYUJiEjtbCu5+hQMBCVRkOwZsFJ1CA9vsriylikavtVAvfuvDZjG/nH74S
u0dzwCutTMtQ54ZzOUgKbfhgywHJvWTpGanLI0d98qi5zV1lzh1c/kPl84DE7gd0
pcZ8/GW6kh9DWSqA3o/XWV/DzVVb0DecylEkAWaDKT7Ib91ViGOO2lOAKmGkL0kM
4/W1tpWQ0+/Ziserr83WNdWJH0wQzgxYJ5EWwXKgQn1c/iNANlnEw99tflWefTXG
dYYd0nO/ZpKRkcrHGiJ+WLxruXBeEV3rSsv9dbcpS1gpN3GIjaBwWxLlqtsO+D/A
yuJwN/HoeGckJJQk/Wd5EeleH3ldC0sZvssjcKdDwp3M5cuGnMY0ruxFicjTUF5E
Q5KPAFdFXWu3EregWunWW15AtQpRJgM+CJ0J9tWy1taBxIHyqqP5mIsfvR2ayCkR
fMEGiaOf/7/YyU1ndwSlWNcQ5a6cl7+MkKQEqJk+lY2CtgbW0oPiZ2nLxuPs+dLR
tSllP/E7bDa2epSn09fuy+sPv/UTOJT0uyMue8y/ypRK7qzIT1Q8WmHgUpqrd6EC
OKIBQC6cWK2plJMpPvR+pNH8aVgn+aUZPXV+9QqoB3Ua/0c197JuoptbHRWKwCHr
iWhc0l8mWJNSzs22LQuf3HqFj27WSju8NgeSn1i4vsg2NoLL3xV+TaU2uEBz7E+Y
VOjbzxHyiTj8nO97ztU+rzFNrV9j+ryALvOwni5DJdaaQ/qvYE+LP8Nq0KjYOnQN
/I5b655SsnOHYBomvdDUXWF6QJ//a1wx5gX9U6CerDKBJbH0FrrZtP74GHo4yHHK
VB4DE9AtAuS7cor4fry9Wr4IcoEJDAka8sRNNm4WisndZ40DNngSs9+9ewj+50ys
ehDMP/5BBYZViOzw/qxAvVBNqKaMqMsZmTo9B3FQ5JkP0KsyAoaDShBsv912kCBI
P6Ymnx6sGbs/N2NZfkz4dPQnlOr0t3fSjXARKmedpTcAjiC1bwFwzL/V1fgeDoFi
pzJOW//VSbiqVGxTMmtSnLskaGjPPi034415O9p1eIveRubDsiabzYnHIVJG2891
JvVKPpUGBFR3e/236Z5at7MljhFUkVnXMvz+d/hsMUmiiOp7iKs3Zldj946FRVxX
YJizHQwW6t9LhL3SfYe34T9bPUbPFe+umwXaC4y01tPT7A/vGBqSHErsNIw46nfD
a/bvHVlDsVL4eWt2NANO11V4668T6SLBl+LnLL8nAqxfCTcUn09Yl033cwk+CuMa
BxNzbLRRFvCc6cLwL3dlcdiPIUNnieMk8xeZZvsz1x8J0zn2v6GwouQifHJEprXb
texiXZxxBN7lYPM4svizigM4/uX2ahzPbqN+Bj9Hb8TdOWb9FuEsQQo3EkguinFK
zuH089TNL+EupdUjzLPInDPQGb6LwzBtUBM/nChQP0D0EgqAtT+TJdz7uKjxTNX2
PG4iNhT5/vSzhCBWAiaMRodYti2X/J7UqB+8/TFyXREaeeML1Afq3ofEBr0UxhyT
z1u+SQaUXhBfkafxtssJgjpcnpK97Qv4R1vO1Eotge51k662E/RQoide272Slxm8
cSdzQ6E3EbjhAm/k+Ta7K+bczJsmRohEa/PBYEOMUDlXHLt58wgjyhiWP6R7ovSr
oPujugpmrfrOcyPNn7cGhBCvPb4wHLBcEYIcz/eWsOHhVBEAs2bR/kAqDgLwmBXN
asFWAApmNgtB0fMMkKThdRHLXRoav56IcQCT+HrO42wpdJpk/dgfK285WgCghILz
TxE6w/5t32Ug9CaUUqGeGJE94DzJzqasci1X85jOlwzhNy5B7HBPciCOpjrnizFo
atwZNxaw3dNocYqjmmskCDwGhAtFxCKppLk8pt5woxnNa7TyN44Ji6t3D6SIqg8M
Cp2usmk7IWxixjQICopDm2zLkD38B7TyJedhAyFTEdMZZT7wq2fphAbpRlgwtE9M
uaolY1kp0MgnZnH/9Lyo6HXQXQPSgT1W/v/XFKGhRof01W1UzAu2A3gJyKLZruJr
K7hNLYR9emD2Bd6P6ZaAiLv8tDuSwg6n6q5EDqdaS1R48C7dTBvVuS6nC1Qk6ING
GFpMhQd6ehOlR5+jTs9x8XQeKhbu/FZH8VnbuD0w5oFGGeOZ0EjzrrfQgjR/l72P
4LvVaISTT81FAcenUqIj0bvUV0tpyXC0qzku6w97UYsT49BvkBhbQ3hmdclwZE2p
R8a+CL0keTtETcDqMJa8b+fmIqqHjumRJPuUAZqOgJJeys+ReuryTI/x0CgFzoid
nLhcgNSvr+IzjI6YTBvIIHXWnc7XHwiqkqPjQaI3ga8/a7VtXc1y+wxj8y2LTnAe
2/RQs3HDBH+8+wgyzSQ2WpXiibdegFwRevOZDoBMhuMe5e5HsghGGJOV5/xRf/dw
jxK760FJeGjX0rFc7/XN7LPNCImKRWxm2WUNzWEHsFHimgb0P6ATmSuxec/T6/OJ
ncuSlEAxzhJIAr1lo0oDF9KD7yQgujJo59MRlElrgbZDPxUeiH/03Me0XGYH3Qh/
EK55/mfeJXJSKnsvKmFm5c4cDjKwWMx/atAFXeZX3qURK3XI1HPmSwF0sCmfcDVF
Z5CNLWCCOV+JzZloOpjw6KIcG/4V+lCpNZ8h5X3K1tM9Nvc6va6RkS7tSP6nwmBu
d60seA6zNa4Sh9mA5Zw8L+xmjbGCnYtxPIk9qgAJc06HCH5/gciZeyf8sqTjjXpE
ppmN+MO4OMifRTMVgbxtx0kJt3IdVDTvahDCFXa4GdU766UCb0V51cZg+ya+gE/Z
CoYBXIWEXRW5B5gWL4h8zrCm8dhbpHiSYVsj8sPzgztT0DKq18xFX+T5j9aIWdNA
UF7ECdzEo0c0KeZ3B1ou/ygqx7UDYuL5yTIkzazFtlPZE4mWaoWwvXpHk0/v6B2y
mTXhSAqCiQ+tCA5JaaEHrRV37cBeS7aVhV1CPKJ72WCOdWkmCMOIwYT97/j6PJJ7
k0WHKeuIyCHSWOmfwmrHD/9cxbjzzzdAkYPTgPlIiRfbkDv7bl8KN3qtzMGkiZeg
00sq4bw1gva43TJb29qilTsX9b5dS+fn287zuGISB9vnxd4NAViiWL+YR7L05Rm2
2XyE4HF50hWu3/1+wsNeVrWYFXlFOxE1eRDlEm3SwlE6EefyqHMphHaqs0Emzb9I
nrgcoQIhrEKC6SvrC/cEhbqjeXPPQOMGtd6RfSO/ulfxgM7sR2FqKodMlGPUDCou
AtS6noBZgIg8iO9mYoCIEtLkpoT8sxf5YY3AwTM8FcVqTPCx6KFs1Aq1WXvVEobv
v1VVxLvJ+9mCjX/7S7jZZjV/BY9+fYrP10tZr8Uc5fO3BMTg+15l+89gJi4sO6Ma
0aMvlqKFf5cOz5pEd6ccVKB4C43KiGpBiRKOB+B6IHI03PKBe6pDaTSi6KVBnnRm
jh4A+guZ+FPtjyyyu3bCsjnopugM0Lbwkl5Oandeg8GJUsbZfYxDEekso0m4lfUu
PPLn6Fnv7H8aag0F72I+n4FMzKWtnyeLUMOSGDB45BekxZPAO9i/v5GJI9ayvBB5
K4GIt5lGuMaCu7OVWTRBibbnw/BDAYanvZtG7iHynAGR1l5L9jwdlHElMzBUgase
Ds+/W67IHVA9dz49DT9nO6HmIyJzkksfVORKywp8458OSdwAw1IBwudEcTOq7sy3
kUBLpZ0LMdGBqmPNkCYruu0rCtP5LR6AfyVvUIooNO0DtPZt4q7v6KgPGAE//pgr
uvC60ewajeEAMlYKoriWF/CiZccqysfxfsqZsMYFx1H1NUMmkFL/QNjJm2rmKXpS
CamvKong79sEy0yvFw8bUbB+bD5OQoX3KfyH9GZq1nvmxGzYdmeom7QYkGA/niNB
U2ARV/4oTcalN7g9a6bzY7PV9WZBcZcjKuKHCKB5xoy+D0vUQssa/D5B15YT7zV2
KmBkWNwAxKgDrXqWVoSlAZAaWgTj87sRfYWb9QWkbMnxKwbrSyOgNg/lN4FY0fu1
aCOX4w3+PtBz41wIxXWb64taPb+ZMzG/7yraoulX/GdyJpMn/PscJlZVclT0OQxb
lD5Idi0Ml73A4O+HQnGUEf7cGzX+tOvSUDZ9iVBnkUL7azoABF0/7Jrs52FEZyra
8Q+xXyDSMeJPL9fvmx3+ZsIk5DH/uqaP5mCAYOb1eUJNoo89xwaDWDLkdyTtrLwf
HcNJRr1GFi+ddRe0Z1l+e5ZRVvvXLBaOy4jJbDTSlF3NwmIxXUA0A/qrgbY6ctTS
bVJ/ljA8YDvwVf0doEiVqqgqgiClmQDEdm+glDwna60aq1IfCUEI322VFu5ZW8tg
YCD03w+k2FQFFZ8i6fQy8l1qCS4SupeVAxI+5xCcpWRProzqncCI/fVLBuUNuJTb
39pY5STK4MWP1XhK3gR6OJAp1+UUTt8wy3AX/9z0LtDV8POa/uZYxraVj/gMDbaP
kyY0xI5KvWxhbDKsuqWcCd4BhMM2VQa6cjvritjp7L6dwLf9YGFO1UTpbk5oNj2g
ySYNdbOqFQ9mAlixSnJEvjPDqQevqxBidVbN+CuzrUOSWGWuZ+HRROadPRQTqNQ5
19Y7F4Fkl3ec+/jbjT0Ocu25HgoZfxqLZBM659r8J6dSpMM53iRCZkbIlA0ki7+j
9W/rh6dAd91tLUkO2i2mhBah+fSW0cgTt9skDyxbXm+8O4p94EyenKBpdrTRWzxJ
DJAPfKm1fcLHTIDgJrBnEOZPV6cqaT/d9Sup9qtlw66z2ck8DdArxwl5vKs9EuB5
BmiFQ2Z1qNQaN+fuZwN9xipZ5cQUcPriO0zspy7AWTWBX8GQtHJQ0ve9icM2SaOf
GltsGROmtHRO3X3Ot9m9XvSpCxBx0AShXuF565gAZ0oqzgKwLr3r8o5CI2qn900l
nWqoT7W3QdoK93yzBpckHnBCohhkJdbi6Gvskj5Tha596DZ5ifF4/EZjCoN1fFQE
FkXp4ucumKqIJ+8fumybIigfzTxIaM3boOvhLWBluuNHBabEnIQ7E9J8gtI98RmC
HlOqXMmGzLAlj6IdkWTyWn3biR/rlZFnJXY5+Mb1ovdRSbJv//+JhMyWImnbuOn1
ilFkHuWmV1kepWaz0+exvL+labaoNmvg8MP9wTSnxZ7kGBO2wy5Dr2ZaY98xA797
Ep3XyiObzzl1KW+PQYiKPoSp03kIH0WNtqvCg6i0xp23VdMeawcbAws3LYlS3PcE
Vk9M8ZYsZCKqoLkOzw2oMvLBgWLlcfbgmQL+YVSxyioMI7m1PLWxmNpJ7xNLvyjg
8QyeQ4MA/FsVKr7B+ZJQIB/5PuGZQwKoaGzKEyNFUOPBR+cBluFduRe6t2kAubWn
whM011s5YsioMnUctEeEnrlGMge6rDR4jPpajxobTZXiRU4NM9khtJ+X01gKh3Pq
/CZ++Pb59VqCYQ1PS9nhcA/jact9BBkCmfxZNTh28rFbjkfoukMsQQNztf6/PEOr
V/LopyhBaft/SNv/oGiQ5uVGJzGekTjJ+TkWGNU/w+EbIMx0XVSvxg6PpKvMXbDF
jyAAKVy0/wrYYnNtt2c+DGCPTrXwKa/XI2oJnb2x8NlacwMANMbDkNZGwE851chh
vdmJ4wIW9HArTn3nP6z2E14aeU6/We4OPaH1bnpnHEGyimfZKIC5o/bvSWyhmM75
spBlCt6CJGMJKSWRXuX/C2byt8xwJvqLCqElYe3TBMbGx72uEHehqXLr/RXSL5DX
n0B87UdBq7h64KOhwBzpQQy+nt9sb5G7fKTGuO8mnDRPhCSJReuL67gmlSrh6U81
5OUPLsxXKGUWuJJRAxEuGJpNsQAwPlXQ1/CyY9pQFLBi2gZpSVu7m1co/Os4QqfK
PPaX5hoRr7cqiLO3REJwsqbyAA/bfIdFUaW6JB08nXZhJBSuwI9gfiGJa9TOwsWr
0mzCWF7pQczjWJahl/p+i5wOdVE7i+gmC9a4DQDyjHrIVuaM7eY00od5nBJ12x00
L8J67obLTD79Fkz/7Ki8VWjhOesFMklyxEKXQBiqmfuAaG0cLsz8dmtZfRnA9E4k
Eg8h65O1OkN4Xefow/zpvG69vrqrw2Su6YFM3QWo4KsnJQdUNW3NLayNEheNPsB7
T0Ap/obN6uB0POJCFR1uZ5dBfZ2dKbOyWHT5Lrb80ziK1ZenieVycssjingAtpWy
i5u2vbnL3kExDwvFlHnjzOrlMZ7ZFF4R+TiIIVS/cXJE6oj6yqs4+GV/cDGxUztP
Ukd2dScR34+z8qFnumZ+Sr95rGeYdbhotvalhPbdTSKpS6lJFQY7GmwxpDU+TjZE
yL+386KrqjFrBR8eVHJa3yA9xEmfdSqMVqrNcX2wSdaTkCNoDzcz4QQqK/H4zynI
QvrPiLt0/vSTnaRy1NI9OyzayOk28EfxIXC4L2QdvTtmtZpY4qoIb+jMoXdVfCQU
Ufhx8zPbfdC4NGz9SI25bzGPKoD99/Nu4qfOnwpzdNuggsWyfcG8XiY7VQjWQE7C
ue8LkN2tiRpBGFpk/YF7H6aB785Xc2jxKCLADxEjSRD+oFahpbKUvJCsFssnEmM2
as1548PAzJ8TBO7cq3a3Tash90LTPWbA+5dJh+Hg52J1DRqE7eNA3IWmyAzvNzkp
AmLtMcwjbHDSnsXQhD2SlY3SAcIKyGGze4AxwKNl3TMi7G6ciW4TLXECnqPCVfjc
aRgONpK710dNg2E79J3M4/2/b4MvpCXF9/3v5HQj1iQmPijTHgnPyy83ZcOoV8Qn
4j04MKTze7KHvkqUvfsWo+ne8QInzZqgyrOQVG6WukQDrdTx5K9VdImuVxOZ629a
7bvgtJn0Av7kgLQ1EvM+lczLROk/8GTr82k/c4/ZoXqJm0h6TnXHgJ3+fvp8Ma4F
1O2SkdPT3sP1Y8XxMPUbiKV76ft7jeEvkZJvgdClL4g5mlohykjQSp+aWMjTAFI/
vw7OlxywKlJpNvtHMMerUUOWJFcjN1xtdZZTeLGLhSxHsdBvIZewnsks3pPXAIRS
v2vEmE92wp0QiQDWhF3l2wD/XFxFPXL+j6znHP1Z/VZIONYcpRowmbzIuK55Z8Gr
oh4LX0U28tDVCeJd7z4biFU9sPp4rOe5yP0XN8dT6mOYeyerPoGw2GnyBR//y3dx
WkuTaiI+Imdy51XUOWf4Gsh4Kqir1EQaRWTrQM+KdHyJXhMpAwXAnf8K4RGww4Fm
k0OUtBigkWr6RMkHiOFpvIla1fGF1oPqPXYi7kcWg1aUrciUd8tFRDs9ipQyIo3+
RdfLJAlbJoYJ+myKrfbEUc8nEYylDrfwRYQrZM5UJcM9Hz1bQ6Lb5O1RnO2bZcJP
tOSan3C99Kje0yojAGdbXoYOs9s2rGv0proXU8dE7mfpabamuQPCi/GB6H6Hp8nH
WqLX7IfGKVCvVYWum7z3XK0aBaxvf7uBu+X/iegi+u0yNaNQyVcFuX6pxiDmKoDJ
wdgGgqhLr1MaqAAXg3wyzfyIMmWgd0vclh2vYipoTRqv6y/lYwVCCpempexDxODD
omRftV94fx4zSIBI8J+3vDK7BXrZAt8fZZp9HPQMWljQHxZ7Ioj0nSvr/vXgLbR9
iZVVHAX6iG2NlpqPcOPuiWNy3bwq2PczP2b5tGEVJMxXeYwA3Wb9wgHNRg7hXV8Z
qgHVNJKx2Np4UordyUKj/1uGOuYRqRNq8NO6UpaFc5g1cXQTqC5plYYoJpfXa+4H
tsDmHxVsB9DhpL9NGGcMyNgmMU69xthIaHYrYtpvOQCoT9J9IIsdxFMWpI5DORKE
Cenrbx/8OW9OxSnb237MXH568l2fp393JtLHtRdxpNc/e/GXwgaovspYx5oxdwLb
/ygHDqNK30iXAOt+16V463y2Favex3kO0kL/CZyf12HsnyOrHnXrU+4n+luOZH4D
mLbSAxg+MYyIVx8MhPDqvstnFc3MWItaBpOwl5LXgHgEZEqx/A5kgpIZKbCq2tIe
YJ+DUrDj9YzTzInDVTtxPiomJknVLHrYLCESkHwbXSiLNljdj1Jhb0gjTs0hrhbA
NiZaGly3FEm3EZy2iHoDrMpK64T76eSMNDz4kamKk0klMJ7pdNGwBPaOD5cvfhjh
OqJmTIOinBwa6NP6LGKekFf8avyjUctkZGj7UWkLEQ35LSJJSWtzpN2mz4vBZsvt
ZKixNblMhwy6DNfPiM5lG4BegsLst9GePkfHJIbsDu1zhwxnvFNuD7Jlnw7HaidB
dtFE68goe+BObRt3FKdMfifK+t1qXbBL9yQVgj3OWN/9YLoioR3C69Y0zZZEUgyr
7zkeEJdfXO3DwP1x9bJTfezgQL62sr5vNfENVopOyyP21MGrvJylg8N4XCn/uR/h
diSrJojNEVlXDoScJOu6e4VeQmm7aicUl9hoUl/8KY7Fcy3BxKNAN1xPCV2bLQ47
X1ipd1SDL8agLbe49nqa/3qNrFjMca1tbEZUqvgs9RwxT9PbY3IsDNaPGiWLkoEQ
N6ZmFzgezJXUMzD7/vCWhbCF1cmQL/JYbKloMbcCw01AEgtm6oCHoW7hZSsxAPRZ
sh0+vKSNWwWcNwzeU7npEzOuO6Is37jXrfB0NmD8jeu6qLUVzizMjCB+xzJmfObt
XL99Ejgrj0D0300Sn67Dbl4ozI+0HrPh3IswupZ6/fGIOdkVRiSvsgaQ4OaS7e1j
2SAgqvk7+vwen170VdmcfmuxMOHolCvKTcCAmhoH8xEmJRK7E1amuRp5Y1MLGxSj
/Leb+IxIhdJn/HdMUjCb3gK+b+qaAYzPjDcDc6mbCMbHpGiAbuWcYZ483Mc70q8A
/8wSZJaxHg0BI/kJg9sBtBh5A99kgQgYJROpxz5jP4O7GFCbAMdEtZwwTgJxgkrE
u0zldVQveVCLc0a2bdF3GmbGT42ltBUcWQefEOWIYG+bjqvWKu3+cMAuP8HGBjdY
ojIvDaeJz1k4V/OB/5KnFOCPf/IT+/vMniLvWzORAOII8UsfpFReVp+5xth7SUh1
uCLEmWF/0jRiTro1v3lK9UD90/RW50XkSJ/40s7zV/+nkj0Cl2Vand7nPdxwIGwQ
v56S7iXMaW0bh17hwZc0D8hw7ozG970k5BPsS0MN/C857aKsLhk+WI7eT0Vi7FEB
ze+0RI3F+ws2BHgefjMdQS4egsP5J9dZvKH1quAtorrQ2NHCmDQRlHVD1Nf9fEWU
5CGr0xRXgKZKh9aTI0g5poiHstBqLpR7sm4ttNDsOSIHy7UmMJg3puxd/DTMK/f8
+H3rXbMUcEcvogZA2mw+xINztk6lwiC0TQsd00NZ5vywgiM3JEx17Uf2J+hYgcf3
0RfIq/pqk3PH94AVhkdjIsZuevLaB5fSdbK7hHIBtb6+xGvVJu7PFq0LzjNRxViR
Upx37FzVlMqVE4Fy3ymztzGjkCIuPYZGjbfKCU4w+h4tI6Mi2hd0XSYQ/jf2ApJj
RqhYWwpEFXy46qAQdfS6OVSoOgjWW9lf3ngHihBZdxi9V8N4VL1unjSSXYE7RyWi
XgccKQFDRjhvXH8vHSb7u8n0UZBg90aIotoJByxqET60vT+y5uGHzpPahUuojDS4
S2WljQy3Y7hbHGwKUgv0ho/dWtQqg/jb2gfokNjAvg+/RtWvQxYoc0GlH5Swbqig
sAWqMfHucqTzoVYnU9IitqhHG/7YTn/W7UvQbkuhErSmSvzGMC2WyD+Qreg4qgMa
lB12y4Bv8q5TubiE+LMJ2B33GsPyeQKeiy/bIo0J5o57y/BBw8Bt6iv2VGtgsWOf
7y7N5n48U366lnum3GSgdXp6Fxfqg6rvVQf3mlcGKSoPV+Jliz/gMjA+Ja0c8mnb
mVhHzDExoaxobtHjpIGXIO3eY555gvgFMrEIfC6TlmFrqf3XFQVY5w4drlUDud5Q
m4G2mfx1bqQbbg7uYHY+7MHvVW6qvinQuRyMwNWbJbuWy0YX2sP7LhZEaMrNHZa9
g6HCWBoEh0L5sFkdfTVhR4AfqPeJUwiauVEQ30aAXpIQBT0TgxY93p6eD5d1xOPz
aLuANEzhFvAOFSDEMpzsSg+M7/z685el5b/+oP8PTFA6IHv4zPGahJmV4LYQRBbM
sUeisjAX7cpwHMjkGhVP3N7hyUnuS7T7OYR9xn/Qw1BXadGvMQqGlQezaMuJQsjz
qYz/YYGW9zApK9GFrnxN3nUAhn7MYG9VOASvtM/bqtV0FWFSmg9U0CQqYS7EMmXt
7YFKVZSdPaW51CTdthX8JvYlaC08utsJokrvaJNO6DKP1GzrsF4lcDPSPMDbyWke
0CjlzE73Lzx9a+Q6zBcRYr/gBPAb3QOSyoKtVRDo3aZR7Yw+xaXu/y57Fd2P/pwS
rvoScAxUq/kAghpmY4zlzL+Ao2qn8Q0H4rmGroQozMWMiuUj2HGyhAEAoVKc10Yd
fm6P0KMIyGAX9VM1BvKFf0Fmu1tbetqYjMhIM8c+u1gWG1bHSk1VZkXmeiRVx8OE
8nFYACoEHt/6jODTijkyCt9pfZSPyJQKSK4FcZCHEuLc2iZeKRiKRZk1YVWTUd0w
Pi1lsyFoZlfyn+lvwxlb/yP7aJO1ocijwAJfqkEYzhnT9EQZBPoAZqkSfZAZuJwZ
paTrJVvwlFxjvjYJI0VbWmEBx383Mqh8gCfO5O+q7KmLI3OMzgRtdOwvZfRP6Xb6
P9SFKAMfDUHqFok4T8K6LunjvpSGhllbd+BQ1ZuGkA0YdwFkGj5KpznbZyLy/tOI
rWc5xAcDX6t9Cy3fpeJZWxPpJxmVL3zX7Ho1XGhAyH2MCxkSPBa3pakxcmt9HIqg
ledX2j10GPAayS1Tfwg4fnrTjJkqgYJtI1BHc2pImzpGlDviXkRdD130GT8BR/8K
P76QaGfTNN2lttMej/2vyi4jr4m4alBPGqV9BxFIfpnigA8x2cWUIn7jJvdrY9TN
gzPs9kyKjzE3TrrgXNXIsoZtPSolNJpe4Qci0RNWp4CClTWyx8KSdyZmGe9MQXbR
FgUnLAgATa9CLoXo07Ju0GZsMy3rBAT4aWWSfwKV9PeYTTL7Tgsweuu4tc5clE7Q
5HpElgvwdXvDapzMIDmOfU7Sv3W/L+y9hswbrY4aGVbAocpxXiodJoZTTU1McN5j
XTRUNugyxsOYqY8R9kkmS3XR5YVFD5x58AolQbP9Zl23cxo6K72mqfDGYtg9FqwO
Wp5xZyyTsX8j8+rHWLDUFGdde/ia69+mBcnOAQaf2vAyanhzT9y68pQDcZp9z0cI
C/bQqgY/V0sI7sHCbUH2VvzXpQQv84uJ4Ur2HyEnu8ktXpnzJnICv++IO/FXgIP1
WaYgkr308fjlMF7MclgfE8DHFyXMubjhVbqn6u+lK7cM4rizAt0jy9ZKRYy6sXdd
zRiQ+Y023nLlJLBOrNWPnjdlv/JAGa9f5/kTBzqvFaWabu3s6VakD9agxT8EixW/
D+pGZcRReAsJQRBu5vduNfPSeHZkAe5FGruiHPvKqFQS7S2NiHt0m7WaqrO1w7zr
737CIDfp7XpcFnEwyJRl1NArJo0vBC6o7ORqJ2rNTmhdBNnHeSNLni5Z98Wlfuqc
c+YogcHOs+6l4IDT/Y4iJtXi58kie/mQtCU+W3RSWnDvnltxBAr8RnoZZYk2k+sy
no3p0+8obV18YEyThC5KgN2Czl8AThC0M1EN1h8e2rnvFzl8k/s6ElFHmiABRIzZ
Q27ZS5QL4ln4nFfcBZfqWj8OQaiM3F5mqKxlj8+8Udt0UKYoGKkLp1hPwF+RVZiD
jWir/cISnmDZN+zJIW3Th6o7bq3K10g4IeZJzVnb/OFIiYUShks4FxexNEs7/gTG
QNhicY4TmlvfUHvbF2TNotR6qjcJ1OAyB/lv13hTKAOQV9licWianWMmHVmByzqX
KUrxe7nrUO7I+fA+dwPTZfmmywzgXoH3TxWs4qKrd4JvfAtB19bmISvaIYVFCQzt
qKdHLyIMHKCShwqRS3W5PqegbbUloo0NNhxoeh5jeMVxjUjGz9YkvZaJVyT1LA/N
M5OEzMmH42KMCyGe1j2Qqukx3fPhQzYY8qzaSAiXFzczUbtykyocufrpoChcBIEQ
xAf4Ix0bws+VHsnDNMuNOLkJzlx2qFFRTtuCWyvix3QSUdpcP0OWMPrGQ1Q4CvfH
D1F2RpIq8l/W4wWGnhr2oHI/esFHPCkR1bjGV34CF054DHYxl3DE4yy7I0a4/GYa
Pqdas1+xQFuftGvXpYJrTzxrpvyDSFbYcoRVr1vphbAc1VwL1lhqs5El9bb62i2+
ynOWNBjuWIfzmiaahkdq59sOV9bzOSP+cs7OFCiuJnkDb5Ysgdmcq3K3EGqPxDIR
vXoUbGMwuN6Lb2Kz1QdTWCA0vaqsiGPEzTRp48k10UnOSvXaHQxfvEH6FebfPK0q
naNp5oH0y2HPmRVnAD+SFRN/y2fn56SHFpTadXD3NJrTSOJgAdP+O8wXHS6MWAxr
V7uG4WunJraEZQaxx8UFb8olvkCHFxAr2p8m8vP8D2WMtcg7ZKGNmLxWexLpUy8q
ZXzmFWGfffEQU/4e4JP2vR3tyZziII+92nvhdcC9CNcFaINfsdLdYvjezmgNP6mx
ao2HxIgXKtKPaZhUNVakyQAOWtQluOFMNZsijef1RcuVNTfMCQZSGEX/vKwp9/HW
LG8hXZGBSEY7I3PEeWaJuiBFzBNZvNrUoQTVo+uGGSVOS2imyQIoRFLETn+StrJu
jhxQFmPQTpEOwJe/GCrBRxai2lV4WlRXOX1ergxxVDB3DbCGNbvUZMTfMTTz/Sjx
wqgasp6ZATkb1eee+t2oehkbZH9KUfjDoDT8AHTlCvBuUWQ7LAMLfmTpgNFib2ZP
Dfoodrk7uXGvbbHFoYpLJ+HeWPoUyMMZ2H/6ifKmNrgkkkfUHdt3Qeh4iWmHvNRF
KrFf2ieNGEee8zbVXJOdLDY7ixgERbmWzu9BOzJ/LtVi+hU39Srv3+99dtoDSkqT
zksEwQ97MGtXj+ACW3YALmjxGcZaQQumPS5rDtohPGCjlWFWMfdel1gBSs2dJS2W
jN3jbEjSYsRvCAZNrFfkhQWtXM35ZaHf5OsvvTaAT1Ojnuk4Ecdc4V1NUMopPaOi
PDh69bYgtOqfGi279Xn8UdbMr0ZVF0ONb4tiFa6yl/v0u42yn1puh6QLsbtr590y
mZe/gnHeaa6+aPO6XcBHS0WZS4zu1y26cemD9HjVLZgzwfRNvbhOrfnC5vwpFJQH
oasOkl1jGurTVSwzVTRH3APq7JnenbToRUMqO0eC1KQCTxSzdPgkWWN1qZ0f1lMt
dRrUUJY7EYPoPUWym5cdPOfHrSHueznpHdL3X6emmG6t6JByY2cjrRdejp24MIKm
h0ySvCZF9SoQbwAAfiIz0/tWq4mvwnef9iZ6BfwPjGEQcg4vZneetchQ8rrVTyAy
Ic6/VDVPwpaTkzKGspGRFlKcGFkfgzCxaCQYAhNW78vkbCp83DRw88YzNFJaKeCI
K+ozpdb1w8Y+jCQTEk6TWsoUw5LGe/5AHo7DIJhkeMGoxJRRHoNwrx8SZC+6OhC5
YZ8XAFoIDz+30A16Pz7OHpAcOh+DBjiR87TIzjRXAVg68gFQQSmTXL14FbNPZzT5
N2/R70hPH58VaSvW2GzqBfrMEBfn5y+Su5mjRZlxz1ZDq8cOi/cIXEGljYwnI5GS
O5+59T/s1sbmz0njqhdTRpTwd6Bj9VI43TUbY6FrnS38MkKrqBvz4wWRuMo5Ux01
rxHayDX/ST9hYISsPDeEBOB9tCXEk4xD9Hu/YAjxAGvZWNeEWt6kOYB9G+KHRJY1
6WCipdxICJOZFykLT/AN/ClgH4ghdncO7GbsZWy3/yG9By8gsXt07UMXocDlHmEg
93vGw8YrY1xj+/L0EcsB03ReQDIbDJQlJ2HA2xHH6zjLg9ZGegczCVb8GY4d8KsG
IGA4u/SFI+ic33rqgj2sSlEKUanDEDWYDBgmTFe+ji+Ntd7WCgDJGB88K+c0c7Ye
ZX8ADXGM28z9gXzCClZ8QBD03Ag3Gs9EzqToD1L3QeUvcZ+mVaBo1WGsaSmxURjl
TGSkXvMnUmumoY70CWFokExfgxitpq7XvIO4BzMZednw8sCuAvjd4tjjd6uSLPdj
fgAo9ZM+yW97WfRhoPBIzSvI9s1xqOi5Q+n/NZQBoY59yv7kURNBv8UgmjrkLYtc
2ZKqDZjdBdgA8GhT67t8RF2y2zQp0nTvbgSRtotGKOXrYyF2S+LlLUOIQR8ORAb3
iZlLgKDh4di5meSY/LwT2NT8xJBnW60y+lpxzYiY50jObphlExLaek9s7ZVUyeXN
+ynHoXI6M3H4o7DWmA/JE60kI4Bm73T+X2WDwFoTfSbW/tG2qhsLCyYDbB4dOyMa
teSbJPdhYZhcHgrBppeDxSbTL+8Wm0WS/ne9gRZocGNS2+G8pSFRmCQ0+SHMRiIl
yedH2tr2qlG9dXhwUx3eKfTtdCJX/UXenEEsoxOrEgwmIkjMcynz5t4cCKdRch4v
xWZKmTXTLVvucR7IEhscFJr38YQBazm94Bp9MWoXEyFoqZcxHIbQYpRPsU3SCGa4
JN92d1qo7Bi7x6N7HLLZpQsPzG+9Vy/U1S3eUmnnkfhQ5yX6aeoNqZtLbxRIgLYd
jTbek/Q5Xpi4XqMCAOAGuEpvlwMyApx+makJhqQGekG9RskpYKlBJFt128yEBmu7
p8vUWVa5AZJqcU94juS6zJVGd4iKv4YlH6bA0myvU/nSm6k2EdhKRoC/6hfrJGSs
1uwbED77g4m6mXDixSqpf8XEC0yJjkYFtkPgDDr1fGnSNe6+5zVlnd2SeQzvMWVb
lI+1ItXdwhNTSAZDbv1VZRaoSkrbrlVgA013/ut2hQ630hU/MrhOrnfOJ6QEoD7Y
05zLR3b0GsMsMjAbpH+0oZgA8DGgKesGYzKEKSj1F/vqVqNcOjywXwlyc1/AOuL3
vlJQkO4uhKuT3sLfHvSJASMQgEzh8tIZDSZNQ/aWBbhhu+DVsTo+3pB6QIP3bg21
zJyQ3VXt1nVwudBdjZ23cQoZtQrlV3JLQHONkLV7DX8QnSIKcOXdrV+bsYyqf6Be
Yi83WlwFnGaIF1vs8athOk7ozeMz1LObfdohjgpnmtPQlZ++S/6OR3M3QKPl+lYC
gbtIczOO7peRo/hCYGraOOPv42HzDSkmjY9U/wGQOxR07T3Hf4SoBs0GtpORfo9O
bQTSk1WnXKB3wZRYDqc+ZXE2cZCRTAX/JrobVMJ/D4BQQabATbuEiyQNs8bg3O4j
sQs8Slrf1SW1IQdL11Yoloc1m3hzkfMZTW8nrmRy7UDWNnhAL7nyZrrEDUJLwGmk
usDFVuHn+/VoDpUklu+0NqpedmID0G2qv29VPbVeR8hhQKN6cBvwvvd98A+C7uXj
jkjO9Ooc7jhKIlZBxCzyIrSK7RJ3egS5VxIUOEZOLbZBZJkhc4BydrioMhaLImNh
/vbBhpHJsndyLPg8yCBkPFSefKzRJ1dhsGH5bskD3NVG3O1cvaDtiv+0AMqEc1HQ
LEWyuoZmAymLkug6NbsRq19rRarWq5zVG41mxkICH5w698JvxlKIa+7htWhhs9BU
zj2e6uA9T0ZYfcVWs+mMH0aOz94q7In18JAoqV7A7K6d7a1483zG8IMiuKq90aDU
o14PlgWR7YTER3gSRZwh7w2awDchQGk8bxCv6QMkUaF3tBGZ0D0Fc7WAtH2RBLxB
jZZ0K7xt/Z56jp/cBnHOjoQan3tk3v1BY5ILd+YbJuY/st01zZcxOxGSf/xUyoNd
ySCjaG4vHpndf5uqZZFkr+5mfFJ2Ehd/t+KVdM7AD3sB/BPIXPt/X674wFgpr46p
RFCzxTn7RBcibdG4bXuyp9TFn6hLWHYBjPVhBjaB0w4BNpkxxrDxHf7KOb74TzXN
vPYa0YbWc8wSpsVjPEgve6qLKx+Vpwmo0LRyZjNAkZPxWFDlWsykWOsSB8mN8/BR
xX2H5b3C0PCBgi84CDtg6myHg1CPylYrzcXhs+9RiL7qx3szPx71lAwD6sysB3qQ
otrzwQhhSBr9fW5oJydfhfZjqKgD8TRqvl8CjevAzYtXpMHWJJIciB9hs+w1LEit
EjR+kLr855UvjGaLTjJ9WWDGHCh1IR/F16k9a9lqTZh7M/Hp0WtWQWjlRr+kG8xV
6Jn3cAsQ01X+NxW0dwZj++NdjPo3+08O6XDp4Yf8AQyapUto/FPVmIgFCkdD6ZUu
ULQ38b0ncUQfuoV4i8//h1wuhhdTKKuPCL87UWGL28RrDS5IMpXDDzBNXtOIydWi
U5uJ5P4wC5BePsFzRt5rkrg9F1gMmp/SBA+Tq9bnmsC0c/4BliUCJs64OJcuz4iq
zprRRiyuKO+ONDHYYNF6EsSkKhUFe90CQpN+ILY8vq6WNe6uPSM9zv3CjcCaCtFz
W7P12oV2V8xwsTksHMG5uOezb0NpQuYrdoMN/pV0DMlpYP7inmdAkEuhQplGbQGh
CeO37oPqcfrBqCvxKpoOQGtAJDgN5K+lm3tWJowLyPI99o8aCDeJ5E86BhnYXm81
MAF4z0OXdjK3GWdGpINaGJiac/D/vPPCE1yFnL9e4CukRIHgVjQKKcpTnwT82E0+
amN8v2LnBSZIJyfk7AOaGZrLpey7Me+opdtHzNx4bfjUK8b+Y9kIGN65EXIgwT97
QfpXHTlqETNNZ6WloLGq6CLZDCqJxzozVuYhGzlAlGOKvqRu/SsNmhKPFdgK1i3W
yUACz/Nzd45XIy+4cDqSm2+RjNG7cXs8g3xTIvbrAbuebh4lBlrg/TJ9/X9yXdD+
Mt/2IrjxPPxgYTWOkW/ihiMiPayJwOcIL4Tblr6OJxzwaei0mWHVSDxtTypS3XI1
eWxLR9xuI3sx0XbZBJOIDq5p4rB6apjfjiH3QdKHwE0SsWx48FwwMnERBcBMFgIR
nDZmInjl01S/snARWwCJauJ6py+OTsYcZfQH1zHvClXdIWCiQZdqTfmuaQ+wywYz
QvjUySbPu86+mw+Pf1B/IGDSjVr2zx/mX0o2pObFbjaoDxIKkVzyv3nmWYkpUS10
l2+x0opy/MXSISvOi/7z7AeNkAvkdPyoOyXZNwS27QNOXL0ls5rfvBwfmZGlE35p
ZqrTrpCedx+d0SGyhP5ttQvbG5IcIyhOWnHPVmiF3lSsS5MPoA1JLAWb0HhtEjwI
+WvTAIVYUrCTYHqmiVYlm8C0TuZa9moHjtw6QG2H92TdF/T76kO+yKvOXEhk4W7Q
sA71+3YHQl2dmsETUR1daAUnuaLVyhYhISne28GNOm25xCAWjTaY+GEB+X3TK6oy
8/XGKKiKn2qPX7zABCRpJ6BXcaIlUXM+DVSbwuSiOC5y8RuQui1sCEa8wFaUL+Ok
hSA9E6aJ4XfDnTERbiSwC+wSJte5FV16m5zc1rnUqMWZ/NVA8QiVCwnQO+mMURkc
Cs92T59dd1oeD8af8j3vo0Q6wHT8/+1Mf8YMR7ps7w6QrNQ5ywD+VRDXgNh33bzL
N3JL6W4AS6DZ5YLG07Vj+FH58Aqhi1McdWH6CbAwbwFreMcv4KV5/Xt4aNjm6gWv
y3gVu3gGK6YlOm1K9izn1Jxb5norqQ+dZqso9EgRKRwOviVfa+Ki1ZU8Q49BJP9P
uLmKeh8p33qfsj7HgL2tpykghnrFZl/bLqrA0vMq2B02q3bRXlY8V2d0p8WY3HsQ
0UC12sYC1wU8QcdJgkAI+kJiYceDVZjTC+M7Ucs6+oXSdHPqkOkZ4duLu8ppJjOA
X2wYqGv3UMCf7ohl/w5fK8SiobSBZmboROuXrv0KeTat0tZFQAuYGOmtCQR7aYfk
UQBVCVTE+NdTQIMmieCguDgDESj63PBH3fx9Q8dXnylSuFOtO/s40Frkh+dKNpXs
9f4IA142WC49PsGPECE4Mq3FCUO2fOoJlE4GAfGCm2OlCjMkamYG5wdizOQExeZf
7NDpyPZcFctRoFG/WD1vcjfu7fAXRrT4AjcLxoTkBPZHY/kbVm5PWpTnmzkIX7u9
jhlgWPE34U8ICSIlHiC4mJoe8KavAGNmxPiqfKnr60h3e7ctEhLbVZuNIAlEoPHS
4gMy7ZL3BCZjddGfRW60g9/PJdcqwZieF+YFsdduUeuGVidIYpMKDKKDmNK5XV/q
CwFw41NlhAdNztVYsclikZhMvGZASqykp8u1rxA6Vh+2VpcFN7ujIo35YUlj2rBr
VH8BojM4SWUqcKmUu7S2m/ckoJgs7M2vyITz4qwYaIN18bpmkdRmUtxLWYdtu7gu
lh8ydCxY9Ad5BPRgvKVlJD6dJSC25KKgZYKntB6hOHGfV5kxCIaHi9TAbWCDGOPv
Cs5JFZ+SP4j672x5YnF3S3GH+gXQ1yB6OEr02PF/LMobUPaQiKZQEuRx20gljYjB
lXN6j6nuU/hW0bhkybtOXQDbJim5noLSZic+8ITqcjAHAUHB+lioT8buE3iN180Z
0zugKeH2QtMPG/G0QShOxWqmPJ8oG8mLzyTiudDUgAcjBx2qIWH1e0Yucww5ZamG
5SRkLHvowaGkawN/XUxLkUzQFH9n+9ngoGTQ+ywte/8XHKmvjosq5ypnSJ/s83ub
V3yMvRUfZiGBmpyQMVvtX3RkDdarfLOeDX+me9n5fx2ECzncZrplLl9u0a0aGnOX
JWHCTk8RKZsfiRht/MIIWVw2y0f8OsNIFkgEM2Re/l4/awfdXzeGtRryob8Or0dJ
+BeQ7zlPlyRGDn2Tc0q5rQPg7Lb0jNZwETpu7CylBGM4Luz7caU2h1Vcslic2hgd
u1OWYy4Gpt0h/dvhzqPzSir5qY6z5okZ7TwfSZRWGNp57sBP9XLaKj3N8a+Q6YcO
QsYdWv4sLcEMqA6jRjs5HCEwuKwwjEa6bnh7H0d+9LVZUwmzAxu0pifDNjxFoVu+
8YlsaiXQ8idAC6zHv4eqGUpXmwhR+SqOPWBSWQQ1fmViiLKagZwyfNg3t9TtL+Xb
KhyyMHQVCSEdeW/HEscO/Y2i/qC6fGEj9kmBX+XpKbJevDRx5P5fxFweNsaZIyMB
akIKwazpf71I9m5w/hMzRMaATrEBU2yLGWtx32+BcrnN8ifAEkCXr3s0qBnFsDRX
9JFzoZi2/JsB4to5OZvreWEDX4c4VZ173IxHrGoT+nMxsyKS6zN3yZ/RnQJWw/7L
BfDLV1E9wtAHT26tJOS/jRCHp2qukEKdOFgNQ1hWG8kU/uFPEAQ8Glq/PO5bZx7Z
2ppCMUS5Ng11oJ7MMtTkJbdMEyy7k4AQFG+mnKQn/+rDySlkcrgdj+QCNo/repH3
0O1uo6Udx5QwfdV6N9tIzJhpQHCJNy3BIWlNzZc/tqGx+bifKyr74dZpWYisRGyt
POY2m6Sq23uCSL28L4MIbcYp8yHdh/CJ934M6hNghzzlUemcd1Twn4opHrvj6LAg
jc7aM4/K+fm+grW/JJRdKDlJJ1YrcCVag29NN4r3MS+BQhKZhNW6bgqZ+87tSOwd
K5IiusXrM3oQ6XqL3Gl588v+jw3q4wdZ4Njc/cAqD6Hjrz6gm0DaPWbetmFa/23L
NTCGCOLT6PXOSilT8oFRqRnrN3vc1R3gpBDSOY/Y5rYFxdsTacjbszqsT7fSBmU7
HgHaT7PwS26u1goE2xsN7Y3WI8Rh6z3EVYRWGGQjTvs0Dfz3lgyYTXG38g582URi
clpI4wnKcQCds+X+DOel25aTELSGjJXwSFXQhmOuGKWiuvfRcQoQb3lw9WKtCUk9
5FwI6ptyQA1CDx+0WaJ2TGsWByvw6SenvGR8UE3Kk7VJJbnSOam/XRyJzefKlnl0
e+5M2PlenarMJVcEs0MIGPrB4peQUZcZE2TRMkOBilAzWz/NsEYpm5IwzseMoNuI
VEXIKWgYFRsyWoxFNPcDF/XR39ANFaXOlpgNXz0vN9Nlx6SqDH/qQSoO6b+GoCYp
iL41e+d0Ab12r0fSRjFf9HiimSFL/Q9kk+q4n87s7ZY11xMfuc5YGRsyAvtdPkty
1ABDsbdO43HMIe8KWrAT3ZAYRIj7h6iJeDQyMEoU04abuZCOC7w1AnNIXCteK2Yl
LCdiGt7cUsoT9GFui2dTkpXc930p73iPa2wCzbgwLEEOKocW5UJ3VwsorGgvo3C4
VYoyTucaSvYLCj0uZPWLyuSXFV8HF3Xh3/NJySWBdwH7doSXm801pmWCnlfMse2V
aoam0jbi4AnIRQcAYsK6+f1Nw5yk4MGADuy0PqbsaqPh2Sb122R7dt5uhNJ536Gi
CACwvrfKjqbieVJ1bxHBLiD+y7vs2NNO0vtNTkgjv6c4aKrlnCLpiZ7KmxNYjEHp
A5efLUyRztyQGIbJbsQggoW8DzeOYX7k7dC+XSqHhx/TdXGxoxMRzm/iaIVgQogM
V+RqTsyBdrMq58W6e800/4c6f9QCkeBgyBwYRYw9ZcK0hVWmtKFkHjW/Ets9CKxm
+C7zj2nTnaa0Opq+I5zxtyt9ShsZDUkjLlQrIR9IdBpfrl0qSgiSz44LmgogDDrS
i0gQA71xKbvqrHt/ufr97/50eTIFRLqK1wSY1B+M4RO8VyTDJKUvTnD4KtfHuER6
vAE8BNxnRcern+609t2hTDJiv/ICc8o5tgWhwiOJdbVLvXbBIqTlAfZVdan0KiMq
lEdLFVuEC1VEpEkOmixnkIkUPBs9l/6zQdcFc0FNRVaqTz7lamj7T0Jg3V3zm93z
nBiNpB7xHYSEDTjrkKRyNiSrufLJ4QWYyzY59K01fvDXsJg8YjZ3TkcOGyIxJLQg
cYfCiENqFT56zb8BDNb9JY1S22KwOJ+ta0Lh8j2ZSJrnOYL4cv8bQW2O1aQt5tQN
oam4269r2Wl4qeNlfXK8UdK4BzPGUAYRHyqGpNo7dkKxJbMFf0zQLOhDinHlG6Ga
kQJlSdseXDrjEE4nP+FoNcWnrzkDQYPyvj3um3nLlvTkurMZuyd5nryusU85d4bJ
OcoVEuA8CFMFeajgARt9URT0F7KUBmUf2KbRIhborPiMj/NWoZv/RgFtw2xwCDYG
TlIdDqxEV4LlgZNeYgMla+bN64xhk6XmYB8U04nMT76ZdwsLOefOp55lV7Ve0BCe
StdQNHpyMEbVmDYBKCBBozRV/PsvtYT6dJ6e2fHsQs+dydSXmcpafppbfWCvNgfj
eLfLFUFKH3X160pWp/7QkB6d5xBFCgVa1ugVfLpBWqTNpAAXBxHgm61a8jyA3HT9
6wzhLu7rmFDG4rX+goLLrryBAvtpRYyNHWF8gsrFNG15phedxTxP2MHBsnBRQQja
YYUBI9dY9o2MQNyjCVWSK7W41gngo9fcDzXtJr4iPvXEqeL5wie8dJnOug0MbX2W
K5jbhl/3X5Nt4o3pwSmUF2sErKZiLhOY4Yyzkn5fIWzmpCXsEsTcfjSuHdCu0dpM
B0iIG49CYnuHTpmbnoqtdJ7Prqy8HRAZif9bBGgLusCmkG9d8C7mbhpzTbbPQkUQ
K5NUybpSIsNO1NqGirSAwntIj2a6doTlN/99Pna0xp0sEdyhvJEYw07u7pocumAI
xSo+t7geDyjfv8YHtdTAxON5eWuULwWOBfSa0Q5+5qNKugrGlOTU3OIKWlUuVNbK
wpebmaBaM6Mb6N0DMsUhjGYoEZrEx+92T+rhXuAovaNdr5NRwgM68rAoqbazYdo3
b345tEww6u8G+uMg2C6tJpa/GcClYca0yL7goE7GJqcj2FPfxk+eiOuAUDcmjyc0
AIe9QHEO2rlmYrfyQyY4TJ0iWkxogiRIEjVoeGXGXvjE4GbMDX085NRRihZtIe3Q
LbPMc3TGNEZi7/6Ed3/4iwJD+10WxLl3yjPwHrVujYSIz5c5VYITTgOgeaDxgBr4
eMnrVvn1Ah3ZolZqJmBgiO6D39h01wxfBs51D4kX1RcYTKWFTR7+Fh1A0QTu7zf4
xAy6QjA/uE6oqV0wfYCMUIgHLiTJrwhNWEtoDZ8Fhrlku5HEmyQDAI0qAmTp1RLO
zVf90JsnFUqJXE/PTEwinHMg4bJzhsOyKlNfkv6bfl1c+OcoCyQnyqvbeqiTGQhc
jHu6ykha1XG1r4VrM9yI44PeIYrt/QTIlFMv3Nbw0sw+2pgPWWAWoq2k2gvgE33G
ohFLGKcGLYUWqzQriHL7+zJCppgpqP2RDwr25mrfTM2Tq1QF3Ay/f+5U4cTXxgU9
4psbGypEy2nIRydNfa1aSIbn3zP5YC/lZCEqe+IgZ63TxcMQfvSyrjfqYXhiCGpy
5PaDJxyCb1RmPHiuAfksXPhPnUJ9D1VqzVR41CV7cii/pv7BRIe8ko1fUjYmRYYA
B8XW3h8G79oo5QZ+IEjD4nSGq9Yl2uuuQZuniaIahyfh71y/jEk6zBWf6IuEfXw+
CbbwIejjfamPkuoB3QNYvoTtY4mp0gtWpbGQ716qIdGXN9DclaZwewQ5bsXLM+IA
BcWAcn4LcGwAfU6+A6NQDnTu4U8NRPYQ/NE6+zgCdZIm1LnEwdM4yR+lU4wl3eyP
rQ6aNE3CL+vs2WaQFjmkFv1whpU3AtpAXvyD8/6BSpUuPQBp2HLqm3FbT5YZ3BDa
/APuhbwTuvg9R15PLAN0sxoy7B7re+4wKBIYobqCxeN6tmQO+Cj0huyKI4KwO0vy
I1e3nCeQv+H0CgAH7RrwpKE2blIgsj5ptzvnwLaFnA6gCW9Hww5+kbJcxrddAZJC
W9xB3hwQcvnKi9luwGj1DH35uPYCjuPwgXbY6cHKsvzzSPM7Pvmwoj7nKlsc7fcx
Pt4nkJnfsbNm2pSVk8q81PPGqItZwROpdizrE1c3ydZCQPRpDZIeLkpwbXoV6/on
yoHbGZD2D2yHFlgvAbZ3QjfqeRvCfKXPHp3TUcVjQ7pbpr2aQp+iDd+BXivqgNEd
54OqmaCY9cbzlYd0Aukj4TduHPNFz6mXpL75leitOHjOOcotvLVgM33UbIX4ed1s
I3htdifE2rZBtkZyIyjllm3X7Sn2L2k/+fBReNI6ov7a0ObE6yvht3neVrFHxYWN
l+E2MxAq449AbSwzcX9Tqdw+farlPH5lf+uE/wDpzE1wpbgcfnYn3W4Dftn2KxZG
ncBfNQmKFDZjSS5TAdjqKLJgN9xtRC1VJhPIMBWTOHbsYEOZWZusuOV3fhQV5Fwz
CMzEkDkGoX+cWSfQbaG48q9vVinmhpFxJPSDSNvWWwVjdILMXjlEWCAk5N1halT2
IDY7mUlXJc2Lo8WCYYy7IUmUQcq7SmyKmSYvbX3Pl7N/EZx7YOUIhfOb7Gdmfp7Y
fy56geBffSBDWnKx/BcBaJVSVRu0ejbHjFuIuNmGqp89QPvnvkyny0izi+Q6bskI
Rs8p4wBnnaz9rntaPDDgG48wqBElrzGV8oFH2hbbBNLYgq06za87IIDzOTw1dxNX
8C2FG6EYI94RDynU5xCvc/obyYSdmEzrs/suTDGV+KT3wYWUhN6dzVqBd6LSGBRG
7dX+p9n8Jh21Rdzs92pKGNbl6HtN1h3Qt69x/5O1Bv3me/5cSizROWg5TYiEeJL2
TH/PHIaDiDpwO8NATh3CbWa1SobFfH9J17ZIo3i0e7z31D9eUXx61QIy87VVmROS
OZGmjRlpaEnLsiHUryA3TburWoO+Lcs9syvTpPHM3ub8lSypyZM82Iv6EUcWPjA+
VGjBuTtRemB6yGaSWi7H0fNvsvPS7Jn9m/dWswrMkNsIsPmTeksR42TOaMxRZC/i
wVzKDlRip7cQxzdPFzQRxQ4jYrcNZzkJMeFskeZD4JsKfCuq3gKuGzKRND/v1l8B
3B07J9H0MWEivNZG2SOZ09LmjYX2c5j2gyRk4Z3eGqBuxmTLcR73UfPrLyHFkSls
7N84Iq5rpsT/aU7Q44fLVEGh4W37VAcP2nH5uIN2NWcOY/8pBqlmseLCI7i7rnbc
VumwmSLLnXZBPGPEnIb/iuU1locaLdPWa87Ej8CgsQRHozFtlOCZ/NMnlYJXbHR8
GdEpazluwLh/wsDRuRzbTe1/6+/jR7rSe0phfEA8Js9zvaGBOJlngc4jLLUzEEDo
MByzQPvQjtjdVGpIyKmCCQFY6d9/iTv5jkmj5TMsgmEhO/QG+wfu/M5lGLm+Skuw
3JcFCko4hYTa3zJzbwbKeqY9mSBND/+bcEHlioAZ3EF6+WIVN3M4LubFq/D2JyDt
o/vZEmFlniWEFQ2SYQv3Hu68aIZnv024aU5p9c/moH49cxuIeLKhdtxFK3YjCQNR
FZ3QbA2CxM+I9kH/8GOqxoGqj+vZ6Tya0Ziw1wB9+dQ1xgm+Qs/NV+oJpXFgnBhA
kJ568etMqKSZVckHEj0TinbBi4OK7rUnCj8f11HC1GhYKRkEOHGa+ltQdjidsp8K
DtR4Du9+bVW+MZwZMNw23UUOMkt9U68w9zKKU2AI4ghpwU4VaJJkSq04MIAEaWr5
p3WmzPzo78TQrPudZVxfisLmb4jvR6X/0q6HucrB55/JHHWoPjHcaLYRWzj8O0j8
guo4U83m97H/X5vw0AOsV1SpSbWeQuv/utPR5W/olwHjvup1uC/jWnRVIc9cpscd
4zsr84c7YKh3gOxvh99noeosYJc9Xp9TGfPZ+dpzBQiZnPTjNq9Y79VboXsAZY28
QDa4/+5L3kMSi2i+2LAPj7iSeTeFICYTLY8AJ6xfzi4EGG2hUzM/AQQCktOqpXKg
IlUhTYEn4eCY8HNetNCgCkfRUc0SIqvjhq/82iEttXL3tIq0g9AkTf+YvWHhPvuO
dtJfM+aj5v1mb88NYYlSsurv4mFC07b+mqwvCTsra5sIqWKg0mRvgmfKczbnsfU2
YKIPJc10X2VLCGYoMeueK6wA3+SnrmWbmkDqXqq6vcYmX4GBmYDPweIuSiV15Wx0
LuEbILZH6fYEuT+aB8O2EIojCyc2FGCbJC/hIoJVY2asxibWvHVNY0ydU++paV2t
N5OkAAq0o4uNSTFWCCfBgpngK6/McbDc09dnelOYHfuZulZqqAoktzB/Y+BawI24
5JGLOrCkUDYeRGPUvMjBiWAhSZDCjReqPZajsOUH4bU/wN3Sjnt4JZ/loTQFNuF+
FR6Qwp6Uo3t4AynPVF+qv/k2ovC1fSmo57xI+X1vbVb+5IxjTS1qgogrDwT3v3sw
sYs4xt4T6XJ+AcD3YvcVTxJXzGgZoTreMeZWN11qN9vUvreYC9rp3JHzcqm9iiRt
YXT7nHHLFtiApZnxN5ZMN8gfszLTGpPXbJTE4Javacj90KDkvObalotWS6vUEHGx
As2kHexWpJyxdJKQwmF9pILnUzJrZeBlx5gGaCjOtyP1EbGcCh5JC2memolzQyVt
+lE61VCHLKtaQbA0yon2XIWtFCuZ3xaQq6018Y01g8UK1Ww6ZmHBdSHAh8k+HCWL
WzchS83W5t7LeJSIRnBhUBztM6v3t3rT4H8FjKx0cdWTOatkF208WiQBfX/8g2LN
aifcgVNqkydBFuqvdmO1IhBeQf/xSPWNx/OfZY6tSnwtVPVzTS5rXPF6/HdmQv54
F3mbeKk7TgFQHi6MbbO3ukpdEkJG6XflNySx7OyiwIzhV1cH5JYoBCcyU951DfBs
My5D4cWEH0OvOEp23RlYsavu8Ca3SxyTsMAFEGiA7BoX3xfwAdJX4kP4g4KfKt3A
obouulLOejJhSPzB7qXiYDpQtOmhf8rGPnm3elQTOGHPit1HDxp7hswWkNPP7TNy
EQJScQbxc8+aD13DBvoGEwgpiegpGf06bQLOkUKzafC346T6arNmtKKJ1uynYryA
htLGInIwqr0XZkCOdkt2cMCE1LTtRHCYswung9yzRgSSVqi57KN7JJohybU7Ui7X
THgoCLaVuupyucbxKHmDTdOFkXy+V0GD2Z7sizvBtY8Al8CU+0ZuJmeBEVWhxXi/
BGc0yGQHqGfdCZEQclnk1fUePkqfVe7aOsbYEtarj1UAu3IReWqnjPk+mNiaVStK
723tkuSpYdpEDpiq0IlUffIen6lwqXlAaijdS/L7N2Q3bfHcNyto2hpb4lUP+E5S
NnUyGKuuF1XEK9NqzhDU5rKkuSJqnyKR0pj8H4MnvmaMYFPsZ4i6LbKU/hE2L5up
WruzvrgWC1kEZte8w1o/hpKmUbMcuH56UWK/ntKet+N2z3w7Y7Vz2JJ5kDnD4/e6
btorGr980hbG88ZZREM8XddrSc7FkjZAezvmmN2fiXCejXzOOA+GxKl+eeuwL0Z9
cyOwBas9NFdfpU9/aw8Fdttz+NIiHH1b6X7r+taHFZc=
`protect END_PROTECTED
