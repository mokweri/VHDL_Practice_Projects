`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oCfS/H/NpCItNx+9PNzof51AXDPK+uIhE2ygII/CgFPyyD08xtLfXZxYvyv92VTX
JE7JMKe0o3updSPIeb/+93aqGeOykUqhDy80+2GYKiqWlxlQJ6nbnLoLTObcAcEk
rMWOexoK4w+TPWwAqEjeepoLiyulR4f7a3cGZJtDCHFzHrFbQyMn/7BLu4qyCztc
NAu4pm2UVeiwn9Kf/SIbKImuJ8Qm9NBRdyVBusxonrobW14nsUKNdtIu+YqDieyi
PNOEs0nFgdglt68q/ZNMWofAn6CcYIFB1lWmxYXRaw9zo7FQCsKJGJfjXobMebKn
6f2JszBc73mLpQ9tlL3cNJeY5J2TNPJATH3Aj1TsFeAgzg/Hm3+NulHxUUUdR4tf
8UkBkm0UN3rHejkzcHk27qlSU+sE3WoU8g2Ia+k7aXirQSM1mC/slOn1OpBrfMw4
`protect END_PROTECTED
