`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTE7xtaLoVpgPpv8p/z/u+kVMQ6Z3ssNwx0DIDqpPg6GvXgKCBp9W7+psAZyalyo
r5aeiMxbZT9WgzFTZgkJ8mrN6J9/Ob4xRJn3lan1RubUjQD4JuoL42bFqwjIm/eE
xrzwd20rLpb6hfeFtOg0cU67G1qqx8PQtl5MMKw/yFkDzoJ3JLkPC98vC3WmkBvn
oofUQHhweKuNzTVDJp0z/cGubnmNqno6avpIn3dl8at8IYWyXULfQrtclmwRCDHc
tTYd9TI8++bBsP0CXPo8lsWemT/V6ZFvptK681YoycpwQGTJLJcyps9V7D57RDyX
BdRLb6fPECWt3c9EOWxkguqTIMzZd8dJ5p0b5Gq9ki5eRN4ypVw0/uabtifzm2dl
ZMyvcwif/k35QKgbxckZKTjY+sN1QpbA5atVLiubUQxh0hzf2RdnhsSOnLhaniKR
lp0sn8exGQCiTk5D5HaKkYA7VBIurrOsX2f/2vlzbWHlg17HgRNV0GdklF+SysvP
2H1itJvrtxki6n0opYvuzAJAhgvgfhNDwYd8pVk7a2pxVp/HnnlrS9hnsn9Qi7ku
Ghb0iFUE+zZ9AQmDncEUJyRrDE3klvdsdsCAOX6FcpQDdUjsrXEFLBlUdDN6h6NW
t2yR3Vbgm0o4EJlog9smcSaDoSDEULxjNW3Z5XCU85C45djQAQyHkf0INgFAX/k7
CVjjUGYT4Qh/uwomTbR43RGKKgTmAnFbf4ykdkcRmvDOGSU6cYDx+UM8iXmqPCYG
OFlrjZ3uvQlR1nwWsrMv0imfvcvEVr5w0xUmsTGilKbOUFCz779Hsn2OC7xt7rLu
Maf2gXIWaTcSiK458COyiEabWANwMrRMbji69zmSvHT/Ml7ibz7kxUta+FiDyO+P
6Kf3B6c1TIpdJhVfgB/48ifmM8cCJsPYZUYwx81Q7yUU6H8KXkxustOWzbVvqBcp
i+wnuwhz9BdqVRHHsy414Bs6ipx9CHYMkBR4NudvbX5mlszfxJIX0SjZRZ51hq9l
Af+WTJP9Ii63PLmEoxaY5EPDnCsF8hd01AEz5IbdESjYkeOa4gwZ6rXgMvg/I++X
TNS2GaB9w/S5pvR/jXh1oyiaUKZqfT/an9f8616bgyQShY9N+hTjNlPJIdkegnFI
0p4AJ0R+pzQwEk+2FG9s3eBAYPgp2OaGZWMycAVZk9GDto/TPtJOMKUpWWgAM6mH
hETi7gm3GKykowP3F2tjP4tp6stCbuPrHY6FQ4ZTZjLD68KFdf10LO5ogeZtinwq
xmx+C7tGLSozdrkkedlwEJDMit+Yg0joEb4FrpXL9TRT2xnvgVviImPYqNWCsTWK
0evKodIsMVcpDkxpHt/jlVtRk4k9Resx+zN6Yh5CDOWHpfVK/ywusvwr2hlg+U8X
J7PxSAw21Pbmej8LCIX3Oqsj+SJrxFc2UE5vBy6i7QguDeJGGb+39ljrTePOspOY
M1SLQOOsdS1HGF0mvZ4sonin7pZiiiYi8EuHVR9HVdXTXsHzSl2rKe4RciqXu1hr
eXrrkef1a/PbFdcCDI4J+FLi/Dj8x0lcBxYnwBtAU5FskMe6dzclyspWfK+g1Cej
ehFSaK/anbXvcRBMX2zTiX9mn85HmQGa6FhjWZoGTvSQHr9RTZTdfB6wenIogtUh
aMgXQFG/o2pxiUCaS6JktsUG+CjGociC1Bxyj0A6cu8Kl7xS8cRA2xLal/Iq11W8
mPWEGwegVjVBE7jKeXF4ZAY1eOY0vAu2riZ/g04fYvvh9HaQv9gyqMhBHuxgV4kL
+Se1zo/jzeRI3W15ENL4SL6wmkebztGxhx+CRQV5JQLGcw5tJ8jW0eVG17t8UE8y
WnpcRsg0wPwBAHyEqHPC8mjh12zvgL4hajnOxpDkj7VyL4Sf3n8ToeMW/CX0/h9z
rPMvxaev4g4kHlNosGT1OA39O+d2cN4Yei9xzHQpzMz+LVkvCCl0pC9MEGT2o38K
7WieZvuFKW+acnE7wH7f0IphUY19EBMIcWl2dE+uOI2gV/fWHyMDiN99f+hlYp1p
x8vtb0nprh7GBVwPlSmmo9yrQME99TDIt1nS7Qkg1Xhr9TwT4UTlpZ2s5FbkcUvu
Pu57GxdONTrmbrlXOeQYs9DvV1Bn237K/Du96QZB8Egov6aEI5KUAUujpOgXjavJ
q14qx1x+CLQen6kNSzWlbDcDBtFmfzcythw03j51mVoqwGLgt+CTlbX6rwk4wUUB
W4IdX5C5tAKQt5ek94nHn/fAiLPje9+9u7kWGDl4MshsOZU2dU78C1ZUN0HJoIYK
WSTBtL6VKp9GRGTGbfxxyIx53Rq35kFsx0k+39UGAemMfNYtGwnD4OiQUMPHpLj6
AJQaFaWUJGp/W3y8tmkI4UAR2ENSf8RewNprnaljlMOxiPq9mm8IDMEAVtwepLdm
qor6Kcl2jYh0qPgXPi0g2g41f5BdRb9NrBMJ4/SLNi15iJ00AWH40KArUxe/cnGu
EaHqu+BZ37S78wsQ3vZkwTDvrBEQM25CSA9NZ9r0TzzkF/PfDE2KhzNU9NyPn+bh
V/AoYXrvT7fxDHLfajuRnYxVyr6at92DnpKbHcNc0B/9PBRCXaUPh9qy8EJCXvX5
d0hZyqtSpgnc+A+kvC9xEEMtbUhBngxUjbYBFZAWBsYqqLXSttL4V2mtnxqbguz1
IufktMN5jPvXHhAF75mzsqAdFPWTM/hoXlIMicXPDXwx6JLs+GSQy6wau8dj704Z
SVqDq6k7LJImkBg7dIkyJ8v4T1e+O38hOgOtHXPGsxE2okkegv1PePn45PW7f7Ds
xT9u5aPTs8Kx++wO9ynLacVIttJ4AYOEoBz5zfSBpYqvKUoBNV8wNAYkylI9dAh5
VAuNNBXGkpbhvF0i6OGTiaYN6flsWF+92Tiz91iiJVS45gZePx/f9/OZPOWYcQhe
Gu9brAZP9ugNS8Y9+ToJVg==
`protect END_PROTECTED
