`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aq5UfrwYq93H50U1XmL7raM0KnF+ept8ZoTDUxkoeIEBunO5NaLZngNQRzTjP8eN
HLHoOlz7p4OqZj0S3RPSR77j1GI5oDQb7+BrJEIbBK57KoXjWMvY8nfwbn080RuE
dgMKhmYAXIjBakz9+c6Nmj4oPyKRLmCdmN5GKQK0nfmwyEuYySzPDWMEhhFeoa2e
1fNalcPOQdtRBHs8P9WOO8S7G6gu99mtIIGppBzlv4mr7ISCoqRjlkFEYclkd4fe
yfH93YoeqFseyf4od25vHoGSwxiP1ChrUkUNn0OSdnbC5LTEOLPm+CVk0Vvm9zVR
UoMeQeC+7Si02mYPQOMxrEDPRqbNkQifAnHa9mCXhM7O548RHL2+/Ogf06jNnZer
`protect END_PROTECTED
