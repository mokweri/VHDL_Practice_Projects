`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwiM7oXbY3acuO6KfxJIS1zefZBUaagZHkSnxoy1bDIhzA3U9+wXWOFL9TvvRRA2
UNL087ReZ8dZN5Cp5Pe1xXadNOcGXZigfbI5q6bgB4N6Ff+J6Plw1G4uuXyL4pUm
Y8PGyLVKRJw9tMBEcssbrYehnly3GXUI1oCejwFazqAE9hMctCktbmQYBKYFMBbX
FCpN9283B8vi6nG5CvYidLlbVt4VZ0AMSwnyNpC9GrJ0SpNA4Vh0RXGC5WYrkyr8
BruUoIrvHY+5bxt7HJPFHgkjO58RZqhZiQnG1V5d8ZuTVXptJAahaAyuDajIs7qv
xKHpqiyRDenlZ0QMtNtKh8FZsBH7CtJvLXDvMG2hvxwFaBr160G4AY8Q+4P4j9wK
gmwxHQTxREJm0DVivgUZdiC9qoaYPYAug/0qTk913+QoAX7ZzY8Ptzko3BkVKDct
mo3RcX85Em6bGxFRVnWA+58+dRsuuSDrKCuwOqDHo6ajJOPnqfGPIH9QPIBXXYxd
BQsenX2+QeP+n07JFK+sUUymPV2khIFgFhQip29vFXM=
`protect END_PROTECTED
