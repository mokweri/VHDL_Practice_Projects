`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xjR6N6ZdF+aArBmzToiURIe6s1z9brfpAT/XnTW7zx5k2PMRpWE5GLPnYf04LCfE
BLZfuPqytqo9NtpjQI7HB65FlSqkeFUKCinSTIMeBt0jqD5ZEtt+gII5bQjBsatM
olKbQxrkb64YWE9JxzsHc51RqKbLBHlgBMsA2/ZKTkTdDVWbd04nXYWp1gN6Hvye
TR7mIOx6iGUoBeFoJ3pgArnWgWU8VPsUaXVbKdXvXx4rVrAsje9pxjy1YomIr4Ml
YZOah+jI0N0Px/gQfnVI2zBAc9qvIMKeqewjE0Na/1EXGW02RIWKAzTYmvg447gW
z72nbPl0EOFWaMuZc9qxeu/AiVo2qTieNE92UGUuUSgKT8MI6XB1lYbr7aNIu3I7
AGTnMenbC9v/LiSK72dTIv49BnqCKsoMgaM1VUX+3m2kt9ANGBh5aRKvxS8SgRXn
dq2m9OUFjSKDv0LAciR0UKglqi550o6t7mMSZ64wgMTrs64HJ+D6nlgRzjDWV2sH
lvno9Zd0KuNbJ7dr4ZbWrHtWALIdNJlU8zV5Q3pMPLMYHikU9+sUCJF+TD45bvQ6
`protect END_PROTECTED
