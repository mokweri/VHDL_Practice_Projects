`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ru+Ll5oT/GGQ4R+Z6g1PGeuIJc47PfI0eY/dPmCNfzOSSjyOVgBnYTtSsvbzbG7V
e+/A8jzp7atlZENay0UVpwwqcXLLA2cRmT1LB//XBpTlRr70gjv0lZeobmqXQym2
+Qy0jA2qPVf4H2Es9JA5R7GNydkgfKbr//xqga0/EsTZH67gFTaBxR+mOmOaOl2T
05Z13IbwC/0vNFaemB2IvJ86b48Evdb3me4C9rx8/HU00S9ffB4m+h+YjrPvPT/V
9lwtx1hlDtV0Tm3p/9uwHYF0FRL0JaNM1hyE2I+5Z01FcUoeGFxBSwj2FKOwWMBj
+x7S54GlnGiNxgTXHZQ/g8uzEp/4MVR1+EqyI8lwZJpi1ttvlTX/YRDUvOy+d1av
JAiclNTGrj5SPUOl0/dmCPi4J4uBjXA37c+8G2pc9d3PQ0deQJ7Z3OlMWqJeQEWU
fae1+xUaK42I2ADsOAYgmx9xUswu7luBOsdaOCx9TH8TFtyLnKNMm7Bz2pGnd/De
SWo64GjDeIYLRpWcpN6Uk4ueGZeZ1ar1wdXcoDvUPXknhvXhaLlECeZdyhE1jdet
0OOVKJNEVV7ORHRkWAfGHfeTxo30zFc5HAlPpTqnCXA4Iuq8dkFDxoALlIvc5/s3
MEQ6eVQ5HCDOCVqty+MQC3MpuCQh/zQvkVUqSGx67rMXojZ59jOt4eDT8iumbaO7
ThnXWY5ONeMfQyktTx94WOe/hPg/usEHOxR6oDWkJwQ=
`protect END_PROTECTED
