`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVZOj8ZKNeQ6AYp/QHBRC3Ff6d3/0zRzOaTa2OVLQlar7jfSwK7TI02b7YxRxxtj
yuxnXWHM9GpaeTV25RUEuVHeQdtXSDAfkTysFq/0YTek4Nn5DH4CnjN75oHMndop
7G/3AKgl0ePt+nCat4Ko8E6/tyOU5TkTPn+ivwUfmrdV78vaPO/ljsE/1jbtGVoS
O88SUoEamYexmeION9+xFtWgXLe7DEyzp9kIgLdjBNzKhhBQ+UE2scpql8ShD+Ql
/yTU2CBM+7JBQKv0m+z362qniUnGJi8nh+QcLYgle01eb4AwRUCU2WOK4nrvAZR7
5gKNBVxa2N+aDJqH+4tBbUnDLuKUHuO8m81qP/23xtF+dn79Od6MInN9mAZIbCaW
wHIAX7QUDO1jlHv5jfO9vA==
`protect END_PROTECTED
