`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgR9JXj40j5n4IfH793U22/+e+k1mAKMqWfYfR/9YsUh5/mpO5SSUkhZ5Bzr/pX3
ICSGY7jiwEWPfNxOslSsHAyUJFmjQSPERCQGcC8zWe8jGs9dIhwlL0XLGkYiRo/k
jhFMh+e8g4h5iQTKz817PaS/4f9djWeHmWyeMFc3KuRfah27CsibpZoYc0qOWGDl
+E7ixBR2w0Q9CDsmiLtWlBxxdl2PrHV+7gyjX5ii4/YMu8vsb3FEGPfGCHBC0CxB
LinWUsEijmtyvsEBiOYi3Qi7fQOPz/tExhd4H+cQYKk8engeZhaQEQqsYXUD2NFK
AtgBmgjuW7ONFI6sc4ZqyuPbWVpJN3TJZKkfBHsmCgzqiKAX0724639idZoT7PIa
223e/Ic9qptdogVJ5g2yKB2yN400XYh+Aquq6zYjayJQDcWWPxVTsCTvSwsB58y4
1GpwndHV1gq7VaBi/r5cDolnjjWM/aOiwb/Xglm1dT7seKGa9M/3oGafWDxONM/M
MR1zObmGWQu5deoJgCyn/NRAlpOBPQrdodZ5CFaFbobtxXi0XR0P3B2veScjs0cd
jlQEFdnowVCpbZ1E3sLIvYXc9nvALzuLEba1jUoIrl7QoZfz2iM4mkYMRwhWiLxF
CMwDDVoHd95o7jYfAb1ifjCigK6iSKeMcK3ABiTC/Sv0McOQXWEKIYvLOSe3dDJK
M/SCCgZ4UmyTRPPnkrigBqgR9e2CjxpDKHGGgxn2G2M=
`protect END_PROTECTED
