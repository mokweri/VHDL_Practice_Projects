`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOUooIXNrIkqTxm2AbA9Wu4Gcjjlo+Q1EIl69evyaoLlp7sNfsetKb4Pzd1jX+uX
RvmUnf6nJJtVNtYjV69DHD7wA4SoG4OSlt8xovAmPMyXcnUeS9LyXpatyigoyYnL
NXl2e10JH0AgLLpaUCS1OCj86E6GpO59gy+tvR3gIelBw9QQBL6i5/9+i6pm72od
zvyLIfn+lMNFQnOvqcdnFcIN0WqmWcVT8Oio8Vlyz+7fYAQxL6u6Mpn3uZgWr7eM
WtD4N4djdM7vo4U39UU3PRfM20TO6bPxCoc/kTP1/oQfNk9m58E9ihNysE2hlLjp
IreOyNaul19pz1MVo1n4pE6JqNVWOwjOmQAxA94u17X5PuH1s9nf+nmPo1QHvnIk
a3Xi0hDcPHLgW044ei4Mf4xlgpt2WPtSGLok0DTO8QWrdfQBsQa3AUBjstid4epI
0VqfSpeYBUnA3CNUGm9VHuB4ZGcpIBmjgbp0ZsdGe3ulhIWIC28xhn7JIzce71Vu
llPmKmQVJMJWYrJ7E4hm3C3guo7f0yzizDQBLsglyDqkF1KY3WcQYj94S39i+KjE
1qBurtK9rRM9lhfBZNx0FD2urDdlR8Cw90dLP8v/g3MGuhFtu1az99dxDy3NHL1w
qUBVoIzeQ4g3aKdKHDZk4el1KoKgD8vXPrCO+OKEsvpFA8Yc8/e8uk84kjhW1uUh
yh40afLW6gM9L8OBjXfTCeQYn7kFx3izizr1JaGgKcuWe9njZwvaWcJ2zCfSOTUi
wK6iXntOZe8T3woi4z01R3TLQ232tqxKv29K2cF1fF7Njub8Di5eCm/GtqzBK+68
a0DXxBMDThDbbkabRw+28JxwOutz/HDuRG8LcswME22uyceej6NzGoNJ2Nj52HLn
tfAM9stfoxdXGNxbD4tJP1QDMyLCFg9QA9OkuZbj+4089aQIaIRKOiTcLfn6VWcy
DZrs5M8vpu+wjp385yO3yuBHXdFJGQieLwnv63V7zRtEB4uCUdxlAp9s61E7q1au
PgarFV9IVeD5juaT7mE38QRad0rrtd/mxt6z3UW3U2goA1D1uWkdOne1Eb4VOF+u
UTsfBLkfo+JliBKYB2aoND4cr+n41sUM5ilOR+6wL1TyUgkwz7bKY9qgEBv9hl0c
gLGqTCh+ahvvDavhIotfYn0Z4nBVrwQRNLqXQP9VwpFkAwt+Q3OqJ9SsgABnNiGV
/oAIAx5xdqo/YF5qukmcmxan82OxUponr0bkaj5uAAOgcUD9z6PiCVPqYcWB4G41
FoH9K1NNp4DniLuH2YwclaiFN9CaSabPBGE7ReyGAXSur6dQlHf7hYBE4nLFK+UZ
cn371dJeXbMbHvtRpNY7qrpP1ioQaXQMCFNvluybSTO0mypiDD7P+8XLtSG5Ci6p
iQXglhUgtTxK0TEjoxGhSBoE00ueZk3joXuTobDVrNfljm62IyeIeqpadHQXKkxE
G55NmU1gSMjaiLLUHIlGg/968jbN2PLVvCuHH+plkuPTJO53Q9dOoyxNQ0ksBs+8
jzacj4BsxInnmqLKVDMa1d9X9KuuXe4mz+cUOFlyNU3Jstjfc/qRbjA1pvrNx5T6
yOtLpjdShUh9TAEIn4scGQ9rgPD8c0kI8o4naQW/sWiEczkpOM9K5VE4uR6j5EMA
zfw6l+yoUX66unh8e1/58OB7F4ZzwarUaXVyM9zRLDx++z/zkJyuDf1acavbvi66
/IjxwunWibn4T+r3qQPzaLpokbIlKrkWs+c5JJ8RZRQeKoA3yX62H4Gin+QrU3/t
Nnj/fO7gDqR1oISjoZyArntGUc6XFT6tLUGyi0hbteUfONBuHF6AfpIyL+i6rGxA
YaAtGDWNhJQ+EH/FMPF/tD6akRn+es6CuxIBA4xnnvrOnAifqZCv4ROHsui4ZP9x
3jfdKj1r5LnHXcATAlYtdScV2Sik00B49p6B9K1vZYdb4MRRugvKE0D84zcBrzXB
qaCQ+zbKEzx9hf5lpE2+bBpKiQQWBJpgfTZ7nXsdLLUwayIGxrjIEHmyThOqZGCJ
k/UhFAGNMsuWofQjkmeqii2qN0Pu0jM8FXdQwA0xSDt96pICff5nmStJiiiA22v2
kndZFZZ7reOkpTJA9F+COAKD5dU3ynpQ0NMR6RnblQHDa+pxnAFDyuftgRQS/8d2
2ItgTCUUynjF9dqvJP3vZLD1hweP43/QN72418mN4bRWZ2GPN9sxxHCDz+cg+E5O
Kh3KTLWSVZjWK4S7YLEygwxGBhWWhSQvaehadOsr9bgJXOgUOMIjzFbGkbDynoMD
g1n3Vow5Bsb+7F7PURqtM+urppq0ms/+J4Q9EQUL54Bk2krZ05w9g1W/CyuyARrt
FWEOhCCCj+N4vYJHdYwnX9I13wq13ITAU/1Z5yjY8KxhJ+yb7UeLai56I9sV/WPP
D89ETnRpH4VtUYFPZMfrBD6l2t4fog4wXiIgI2ja9xMCwsgwc4kULboKk0JAeX4S
2huKnaLnth+MHVaWyjEAAMT0ww1yTZd9K9oZv5iu24DAXwVB1275JKCtYVgr83TL
iKJj10CZS0poW+Z7zs2e8Hk7GeiR4NcnOJqlsg1E9MbcdLhzMhQqpaNSvrNxKPkS
x2KnHsOARG5vN1rCEWHth0eXJ7Yb3Hro6EeBAMHkS5CEV/Ud1PvLMV63k2o0KZeS
Hie3rk3tOr35sCwLLyqTiVc/UNr3Hr0GAo6TW/4/bEyDhRC/sOkUJdKrwgTbDTP+
5aR1D6kRUSigCGvJwoatL4RTPAaivBORv5lDCwnxP9s2TynatvgWlc6+TSgQu4cW
+pD+nFoFjCFG9wi7SErYIl2lWHm8rv4XoVaKyTsCbOzLkKQNPWuoye/96DFB8XOV
KxTEV4K3dYhvWRZFE2sofZSLt8Z9ZjW5MuYvPv3JP+qCyLxF64a/9Q+NXDXtrEVH
eVkl0p9OHc96ZD9yy4DmLPh+dkNvCwqfIMFxXSa0E+K5FgPf85Z7adLXsfIc98Vh
j88Nk1mtNvc4zmhHmuCwJQZW3P3OnjicMCn+j2+THu5WMjRw714b0HgoXpRLcPc4
iNuI7dzGQtUu0zFL+xJnaGeJFSmCWRgKhVN/9cgE1cmfTGXmtPP0L37rrVAKsGkB
c5aW55u/iWKh8WI5VEjikFHRYTbjJmH8VtqLsgOcq0vNeNO1kI8w+0apR/iGiS6d
o8Q+AV6dxWlNyqu3FSahLAZw1XMmbkM4/Jl8lW4ndu0iZ3b7X1j3D4zU+361gxUy
XMj3m01PbMhK4sBfasEIRIO6QaiPfcFvIDRC/vfh/V4TGHl5bIu7rJCrWfpBmR2C
f1gwX/MR9Wklh5yaTbhGIb9bwO7KDhZI9W+gQo+9jQ5ouL1kl6hRi545IxhosIPI
/5iBKSH5WR3tEMM76qQBd5mJFL5AfARIrrofoaQrcZFRFHjO44sgJx8uWuw4EX4g
QGLH8V3u8VrQA4YqDgvfW4vvjdODvcy9z9y1mJX7LZLT0vZ5f3bZdsZD+NEylgEk
DCcfcVeHGhOgfnjzMm0QUwLjlQF13ymLwDZApDELLw+zWG8z+8WN/zjZS71oH0N7
WbIaPyGk6014F5yi5PQ0ChYjbyKapNwlykAdj5Ldc66L83X9JvuO4mAaGU+qwyfY
MhFtBHeNisP/07h+YljsA443nLpOJw6gkQl+19oaKez+FakHDtu8aC7qcjoJd5US
NH10TRjrViJCjA/P0EOjKJn3crusJ/LWiyLBkoMuPt/coaiI7aM9Z5i7L3k3ARgj
u0VBsmqb6DcNyig83AnCX+OJTRBCdeFVVDhGcB+m3SdBF2EFg2aDodi2j13Bupiy
mVbU8GTPaialpAOZ9mSyNxQ4mKATXoc035QZ3uiA8lVPB2bAhldB6037hZlEmDGW
gf0P+btbKRb18+Cc07VXuH57ah4D6tp9nqGezZ0IwUIf07WQhu79G1bxipvIRKWX
oS12Kao6AyRyeiFu6DeWeKff/Sq8+FJSmn5Ha2gdCE+ITw0t8wrk3NQXsxhy04IF
o3ce3tX9TpbyTtEuePFWTXTRahiWXru6FBx3WYYklyxrMJ//nMLQOC6Wlki5goWK
QzNLW/a1sM1GRrFOZU2edCbb6rADW+diJYCAOavk/pci3z41Sd1+sIO07wGB8Aq4
MqRbz+WCG5oJQ82kei//A2tjHjH6MIZ+GI/S8UgK/sHOLRRrsNFJ/AVITKdSuUIB
FBm2VIo7g1RWeBT5BV8qRDRu7KjSNfdQXnjpuFzG5+nAKqR9Bvnf809wV13yRHhx
GgIOGZqUIKbC+MKNXDut3NYkSu8quCEqaPQakrrz8noC/sBnc6uWdAe3Iwctvu+R
gbbmSnwVE6qhwLpiAKH7iKBIjJunmXBChpk9YDJP6X0hmuKAcjGsoTpx+1HjhBCc
780KNmkbewuwcvNWp6MsBH5+/pHqaZNvgO96yoUtBNvUCv0Tw67QBHCFiMdRwykg
aMSzjgIM2CiNBGz3oh+Ul/oWsmLMxJt/n2KrT/6cCnFgexLggVqGSJQ7SuzBiTlW
cM6yw+qZLmkIC7smqDYCp2EEATDAnm+wItfGhaMlWmeoYwaOC6zwgrqc1Fx2uvE1
oz5m1NHwF9QHoQSD/7gjXYLZnEVmRthiPNHtQ4BEuJn4ko0I6DqXmQTYw5Tr/787
bDPg7yGnHIliaHnWi9nYNAxbSu0JzXqMBBVtUD58deaJiXN/UtMH7BrE5e4fZfqI
5o7TOxejfXTk7cXkv+qvEm/UlpYX5KUWUuPkc0DeZlOLRTPIFShaHguv7y9nBNdF
LrCmhClF+cSmPeoDw62/e+SGs10lbUyKVgsuFFg8dppmrS+wSOx1H72mbayQLLnW
WLBzbM6723iiXC2EBGaWfdPVD0il5lBvDn4ttaF5SK0QFbov+JoRPd5GCy0PIDrF
d9B28QYaNjGNU9zwE/36A2lPmWAYo555GrOGglsj4R7e1Eel7cKXLcCdN0HKulrX
+oCkdUKqi091rJOX10kbqhpD9XcNHEJHK9AlOqivagzaueniJfFnHN6hPhgNBSA0
mOLXH+3MGDVmjnYFwYqU0QNvQVvSRFSBr66/CFp1qVA0ktDrzcfN42xvWak0Dhce
tk2ykg+BXe0FdeSkoK0MwBD3htYyFfJYkkBJ99bpTGAFeJpKLpSD5zoABkxMYah4
vLgMgYrooYJ2TZR3siUwRL+HAauvxa8mHyL0HLjRKUW126ajT3WYQChgMxltHAGw
bCxDgBlbob+Rxdzl0ksIi/77VQzBa71XCya4pOdqrFzdnbIWpyUPYhXmxD7gCsBg
+nhfRBw3if4R8XKg+IrzvYaX2fDZC8QZMHswQa7UlaM4sbAYgSCSCHScZpV9EA/E
bF+9LUuv61Xjm2oFLgLIy9+isB/i5gn9OBsXZSBsPqoXUL3qFffLzYGalcvOOzX2
C1N/nLRTjeHKxYJNr+iEC8hprLUNWNSKGyZRt16UZyUeE0GsodVyALFfUWTPYvfw
gQgt7PbOIG9yKJpZ2fo8j+NJT9Zc4Or48i1dYpazrHr7mAuERmTvH7H0zzroA4pD
yeN0k9IOyPxfJVbZvX2jU+zKBShEOmq9xFWZPM22e7UQj7oM2P8GXa6W/YxHIz/i
6/bc5Ba5I3iau6+bdZ0uSpW422P0sBTunjfevd6DPyfU/wlNAOPDmWCAmT7qpmpe
bHT5zFmJEgalnYzC6T9ZFVqE3HilNja4FGCzYQNNscHlx/KK18DeC1+US/euU8VH
Z79jdC8whm6uGvjXTX/6iKyfGstTq82UksqlBKbLUGq/jfiJ06qUNFd/PiTSwovi
Zd12ky0fdKx9TYmWFlyNOXJ8cTYiSuXH4w3PqgSPt1kSt3RRkIuVM61wysip0LDQ
Qtvbw+4VwhJIDDZaVhgfkFin5FSgZVWnlzeR64RmaFAv89XO2Xi+rSH5dAj4aQf5
+4xX5K04oNWdjryALs7pVITZiCA5tU2UC1J+0PlzrJlaF4F0EuqHqyqILcRTdkzy
x7MpaxQWNm+t/5bQy/s64K5mAk8fT/ofly7qaL8BWYIzX8ay8gmCTxvcoGBHCwEu
zvYZeq6AMKxLRqVlG3Ukle8djk98qK31ZK9GPgfhZY8rSv0NR94hgFpuD1rJAsmh
HB9gtFzLEHEC/w6n6Rc/cHv04sX1G8O1Viktxv2Q39myiqoBfgtW9o6xeIQ8Zcl1
zNfSrUeZhEgBMPQUxFWa7A5Pdor0llzTz7l9MX4XJNE/L2xIkkXAQ+77Qf4df8g3
uN7oNllW5OE719EC2bzwcmjQmHs/3ObBdngvHV2e8Hbgbxhhsavf5MIuJcBG4CXV
/gdN/uxKF4CMytLrusS4OIkaeAi2+L2Q3HkpkjIgTLt1Y0zJTi+7ENDj4KXWCwyD
jhhkLnnfczq8yQp8yTGtQGnHUeOqZpo5rMoYUozw7Os3kni/bscoJPhHGnpKLWiY
cf2NR/QderGyWuxGtoXi5vCX6tsDbByBj0jygePW/DtOgqlJqvIAIMVpl6VbXNDN
Y6Qzmiw318tTgrijWFSFldYzb2YrnA4LUlmWar5CYL+DRBiNstYA3vpjD0TpCA6U
bTAfmftaZ6t35LHp4kI8luRkkpasyrzZiAE9S5/w7l2UiXvXyTVurY3yQcYdM8+W
DzoYXMrrInzZZLroTu6jSlFc6ryRYe4wUmxv5eue7cNxiWrxecDJnJPkiy63lvvI
7PvBlv4+U9FlZpKWorIBi6u5yKEJr3EjPuuWGVUUT9GoOJHAIi7x3DHGTara3dMn
fUoWQh82xDkbe4OdaZwk8oiUrL5KQAtfqYJGCOgiVAs28Fq4TxgJ3kdiRyePyYAF
0h8jvhMDzsPrEfaLJcPOQt2f64Bzeus+9+yv3EcL7cU86SKqTtj+TTzsgPyAtcoC
BOC3Hgkgx1GtCKEUs3/tEhMRwzeGhsw1cfaXABm73FrHsBSjGnGEqBh6k4eTNAf/
0e57RHbPy8uYLqMz8/j+l98qmtAxzRMnkpGD1bn4cHIct3DrWg68dUWcb/SaBBw5
/50EuaEDpy7FhMdUpoMMTH39S5sn42A3Vzma9mEIrqRgcwMs3rIacsKJyAAXjFj8
+/11Ne3RRx6eC3mVNbmvJAMCLE89TmMhjpQv/4qc72VMqHtZtExpWIaQrI8esG4O
MWFi+gi9jCK/X3yyfaAV4lZ0JVsPJtz7VyNv13J03TeihNJWgMJeuIsXKBc8UCgk
xB5tAL1y3RY4keJQWbtUktv9MSAqit5dVRSdx4v7pUxawP0CNNIR8DmCskGHnHzC
dzWbInPgp4CASDU3sXqrpDS5+rzGUvsEt6ZwwtxDzEtfBzysX6+KEatalUxm5miF
0cQYv43G6ouEBo4l2D5QTfWAl3LjGFM21xvGxRAArgjsZqy5Yxyd2BGIR73pZ86M
RFG56uq8p3qHN1cVSiWwKzDASpbqVGc4HhH4egP/G8faecrlkzu8zrYUpb+RI9OP
mS9sprfDz+2D/R3RmrzAakxPDxdk3DwLbmlZpf4r2hQv06lDz70J0y31mwV5OEMb
TmB7ULe72ctvyRupWp2ekluHrVCEb411awqwI6c6Jl+uy852C8vJINTp4AVYvswF
LBYKklNXr3ipgFOSpMMHcOXTdsNmbQanTwJu6p+jAQm+MCygmf3PiZKFNJCVAPOY
MFbCBSWUQL393kf88jAM6VtM7HmJJt+yOUV/XNQLM0JcihUxwZDr9pGwWajhfWga
0xOi49cKNnEhcbPqC6lsCRR4Lm7Wmhe3V7P05lZZCWY97/D5xM39mXNMHnadM4Vi
S+cB1mYZuX8FPW5lCHu0fQZhzTzwwq0Zo41S0hegYrtaQTe8xMiduao8br6ufsLY
AxPLKGU0P6q8zTJiQ+Ved+4egoEXvLqdSGf0fDqDXcVYXecBLISlLHM98tcPWyQe
InEXOyzp28SXQy/YQ9QKEvDtdroOp3tmqQNny8pso8aFDNcfsaQC1kCLbORn0On8
1N/5JzmutF52sNulIqgNu1rqjpt7qdRU1HrTrnQGWP2UGVfVJZYsVpiPZjZLyMnp
SerjPyIB8Bej+x2u+Dmqe0LUrvjPz3z8gNcJQ/+eZ1IA9ulrVyryLjbu7Pjdq49j
i/EM5zBaza3A9h+ivIAHRhyDKz5lgpyrmsUBDB7nptK98LSG4HlC08wdFR6QMZIQ
2kMYaZyaqOrUmDd7IpM6E+Aelx+Vuwpe/uuMkocY8gcMsvhYaNtsZ1La0CdA7FUZ
KQqV6SQRm5NIRgzjVB14cg/OeooYxnOnhghuqVSungyRsmcP+NIpWBdFERNOXjsQ
0CyANC4YpDzBjj5cMCnSz4rK5bNRnfrJFiQ93r1RzWrVkvM4S4O7RC5Z0ETXv2Ne
PQHp6hX2QBnC5FtEburzMp2JBYg2Wd7d5Pj81DAujT5HOT3TmSuLPd0caYxQe4pd
Im+A/AtqYxvl3U9mrnlipSnA0W/p9JKyRfXfjosRkQaSMrYBrqYlVZ2wPKXSfHwL
xKL4d6RM9PhdiNaHaWp7cZel89u7vMk+et+1cFMoxaWPQm3fzx7wob9bQi+ARmlC
2oPqnDbncEySTTuoi0hBsfgo/ltv+iioeZ5ldQrlrz63yLGPwiEKExZZ721Ih8NH
/mGU5JGTC5i9V4ekBrjzSK7/CiF042A/74eGTr/6XCNn9B9/BGFHvA7smO/OPq7T
8St4lQ9PWN0KiBtgwt/weNPozO54k0Omdn5iG1hNK7w8Yh2QelWtE8y/aI8HnP7W
IqiTSSIbcSjBkbiyaRBhbPcrQP5zIQfk6dQ9MO7JiuMHxb84lEOYt0PyfvXcW0Nf
gZS7fVIe/r3Wi82YMafsdzQKDu2qCYgCie9/Ahn0oEHQnwpEc/DM/Kw1pdsBp7oj
Fa4RPKeM3CSyJDAj9Gr36YSTrOSUZfr/jToYksEUCW3cBLveK9wvfjEAT++BCa51
CU7I7n8CwVIFGxNhKxbl+tf2d6ny6WJOzi/8tVragt4S0y2zLLhkDKhnyKcu9lRi
vhQuXl4RyIbC+Cy+fxW2rPiSkWe8sG9w+tyxV1oFDz+N5ghsNHcDWWS79Ct3W/7M
EsXsanigDVS4HeKngKZiLfUcGRIieIkknIj6RmYJ/a5pBlVDhwRNPLf7gRbTF6sc
hjk6zYhA4ywOV/wp00tjenPriVjkeDiXzIsoA1iX94l25hryxCAsBeye35MKGd+d
ZT42XLBqIzwUkWHI6I/32qwtu5JehJYzVHOKZxm6YwDTCliMcpITd8AIQgIiYgmH
pqszXvtiYfqklIbm8KeSWq1Eg/C7weC7IVdfkJexyjVNCcfb5An5hZzf/L/5uG8l
hO6tsGMW2dDU6oLOL9C1Yw+tWksvyBwbRn99dRbuvIRdYQTevGjkrwKjOR8Ued6E
K0+mC040L3iyLfRA39WpXGK/4/gN4+nYCipjlx3nXoXrGiu009kv0UfKZBWWn9O2
+ASfZfnR9OX+MC/4rdmcPFouCM+Nan7LfWauHmN5iIoZO8c+MwbXb+koOZKmYPlR
BIOOYhJOYZYpZQVr/eNMKTrHzQ14H8KqyrudtYxK+syhtunXbHpKLVkSas687SP6
IC6BPbRxY7aDOXaK8Deak6iGBkRMEUjJkitsHHXKbXxKDdnLxH6jg7JeKmmtlpFc
e+pE4wRvLR6OHaZh9NNzh3AF6QgFEiBaLSpBqVzPEyX8KjaLZQLlkqSYBHOKqJ5a
rwXNYOZm0msgAMnvua10mS/hYQn351MNV03VJj0hc0knkQkgHDg4npBytG6Sa1bz
SclwchVKuU7ovLTZU9V/TVTNW9eyZDkphLOpYNGYpFTMFD6mMEKCLCj0u7DjeQfA
ko3dxNcJzoY+25XFn4ptqUXYx6ie2OPNcWNyIwHCDb9za/HSIkE34RQXub9Yn8me
Xpe40T4YHcQiDLR1kGDo03Pom+pWDFlE6SdezyAPJpNvSRdQp8zrnopXfXwGvhdz
rzFNbHJwq4ZrWk1QIaAJoJ/04GZagZTUAiZZOGKfl8paHGQpbj/E7Urt6By/qhdI
DGW7dnB7fqg7VSpZTXdm+Qed/KMa8ialNkEA8HRcfHxm7xFg7T/XnLBN1oNhHo4H
PdaDBUThIb4tAHx5RjY2bA3nXnTNGB2P67zN+nTq5w/zRwDRe2xZ1JICR0GPBO7u
lFI3hjZpA3UcDi/rIwVuFqpP4WtEoeWrvSdLO1wsTV0ZRokqpnaqEZFVXYX/sB28
+MMXH6mfpC4dzo9moGNJ+6a/2LNXfplMxWorI3ER9pPjrSGN/NOduH9sZ8/4nFBq
q6VLP6qsYhHYJa4JzxcVQyi2Ck7j8qbYTbJA/UU7yHLqF0JFlCFxJRhfkrCvSV2U
EtfdQMnyxrVKdgcmD5UswFH+AaU/oZk6Yq2yld/hlOyRrj+GCpF3bGrjqr6ENfzQ
g34KhqB6FyZHVRhHm0mOGg2i+e5FAUxYkVwNXrKOJQgf8kF2xwmiultKVYWiznd8
eeamUKA/WRRkZZH/+vXOyk1LArAxd0GHxQiy8uWUXvqh5w0yC9frPuV73+Q6UZMW
y9tSP2Q4LwCMvLkA9V+uyst/Ak0pzUd444kXchlkUs4Gv/53bfzB7aVYaXHP/8RH
w/CrignXE+Rks6RQ4xKTbYR3CNLyF9nHbRybUvwzN9CwFutKof74vn0HbeBCp8Es
Gwc3GBCumOxB1ZGbSqRJluFzTcRUdR6J91mfWgvoOCPEAOBE79STNSz1RwUyo+Lw
RP0ypMbypGg4kZGlF/kuE5SZxizwD6OEbgAaBNjW50ewxUv/Ol7Sfrs5GVJPr7q6
uZyYfJ7yHUY01gYJqlANqk2HIbV5PlPtc6tsgstjIr+X7Mv/c9RxB1qszmnwTtig
67j4lus00Foj7M1wKBfCdipheA8aW27tVnn7FSd9WcjJKvxl+ablUB0nE9SsgpSQ
9zB7CGLRJHCuYnjD+SusHSfP0xKlsrMzR6GsjDvNVb79RO/j70ul2dLrJ4JmCuUX
WSpILz01eyijFKlUIe7d18TYN/ytYWHASjuwYg6zCXA7XDPu0g/6s8CJ3uSBOAkZ
SrWnas3AXbL8D9Gc/2BT1pu4No/+XvjUCt2MDhRwlZSIV+mPuYB9wLWREJUNy1U3
aN4JoN3lSUYNZVHq036q5xYxggm+lCr8EVDHhWH1hNHoxK366ZWqj/M6BZmtdgMV
08ynPgC1Eq8vyiSDf1VtL0NcA6XTPJnCj+hS07zGVTIfKgVGGh+d7MYYLbrrT066
3QayJ4i9tbo4FxidpaIvwqh6jKtXpP1u/A+nLjFQtwkdR4lqGNKwV/oeY/dqZXSB
bLihRae6MYIog/9uoBubCh4/k7lylMvudI89CqJ/sHRPxexW8QTyBCihl/awgSvM
0ZTNNBaXqkkWyUvzb1qnhP2mXHWehmaEAv0uWYupDT3BU774mccRIK3vcy7pk5Tk
o8lRcrFatIPN8bX8D3sveONOTbvKt9j8iPJsjc9YjN96GJy0IGbsFSiWcwCWnjor
QVPxvGkUdRc6FYZ5yUOrU/qsRqtVmFhoCFjFQYZ2+Ao1+3d2qt26EduBjcsW4VLS
BYV2ZWlfSxF9h4JnJBcPtQivrWD2yj1sTdQzaMAYGuRZpLoVN6hQjKNIjEd7IdVW
lA6b7pe6lW//HOIGENB0LpIwlqV1+JBrDCjn5R3MyTddBw5iQDKHhoqgXICCvdn+
5Gav6vNkjr7Yxa8y/zrS+fISdP8QsfLFviT93pkHofanpnytvt9QDsH2QZYJCKAs
G1nJtxSFfEu+yTq14vNCc0ooXodf+8lq+Gn3C8fPxpQWwfeoacVrliGl3cLwT8lW
lLiXZjxczg1J3Cbqa1vlq5vhQh4XuKLE8ULiC2SWZ2yVRbGZYu0tTW/vNyeme34R
mlGG09ll6KKB/r0/vNDY2LQlWcxLfdIYIgVkjFOPLXy15Uz05efTsnyBQlw5koUc
a9vg5Duy9eIZApV4CP42v66wgUeF+5k5sOPiHYVrgle25/A2/BvbBPn21DeJJYv+
inTIdcYOfZapgkXN4mCFuSXG+2YgN9xA/rRHdHJ9xlm9eF/JziWXc34QYTgAcvkL
y8zgvtFI4zVr2wYPxQh0WU2YEHe1KCh2sLe1bNoAu8pL2XoKTxSEc3JmjLD7FZhT
zDxNtqXDE+e3i35f6pgtf4cG5pxwFkImDZh9f5BFNRQG1GIh7bWQmWAsqTRPjvg7
0bn9imUng9ft+Wl4TeAOmqaqTGbmQUIyaQvmO4QdDdoDhtrjScJTtYbKYOxiwng5
qjfs8O3zsmMSFE0cXz215gyOOBHIOxrN7kGP2nS98gEgSih+21qhvGnfpBHZ8spj
5EA1ZhfKjy3JrQiwPcBeL8iW7t6UE5tfszM5ILValtmKn9DGOzMxYq4RB2J1KBXu
2EgQRf0EM0vT6V+spX/QjhQ37nc5yU0qVyQvaHAKxhdPhws6i8NK/V5+gxJ+al4J
cAtTdsBkx339D4ziWTt86VhDfjBUcKfpMJNuGF19LonfMI7SHa+/ATa/A/NFO8oL
9/owd3qgpZn9G2EziViYeSiIAx7y5Z1FE0jApMMmzE1nzSD+RBaT5dCAyTi3mkrE
B42mbOx2CqFEkdtw6AhbJtGAEZIPczHUR5oDqp8V7xvlMqlHsYq+bVrpJeczW+in
Md2ng4aWq/rGrBYPuNmxp/jPziV8GzEuGWUBOqM49SD20GCpcqH2iJUU0QFPH2a3
L8ysdKlkm/yGQ8VmTitunSLeEsaqAWE9jTzHkKZ+292/Jtj1bvTz4PUzabZeKNJO
HaT5AssYQiVZJhshLCnNKufXY43FjBntNTCV3t2wp9hy1x9qS3+yzgKW26A6tFHC
oivXroMH7a51BD33cOOUlwA+QbL63SaxAapXYLhhWxhbW3ChSuJ0p2gTNB+z2MeU
JjKIiNeWoC0vV3VwBbIyRaK9k71pSpOHmGnHslbfbJzbcI1zHlnIA3RzNk9j6cgD
QVDICMXLLecfwYzE4W5VFCtESb8c4wOLYrBU5hO7kxfzrPbo/fPkEEdYw8wYiyxi
f3zmR36XoVSxglbxkd2gEclCZlJ+YHy7BF4y5YmOCj1GwChFp0jIbEFqWrxvSN5c
YMoD5zup5N1C4dD4/W3WpA2O5BoNVdgEvDGqlXMFQ5E200Laq9YfNBihdrOc1EgT
PVAGwBmVwc86FLrhYM17ZSNvmgEnkZJmh5cuNK8UTqv3uaBHv1wFvAjoSjE1DrJA
OhUe9ggFDId0udGNTWohO4Ygv6ofqTS9E73zH4fGObhhZkOEg0ioDDwh5NxxCUGg
gjbdcuqbpLNWiR2rQF2xzXtaTyxb+FI+GHdltt0d5bHMwEL8H9Tt8p+wMFEOuec9
Kz8v8dQV6qogzdUU77qLaX3mFcAJfIUeTx32XLmqVl/7QZrVHt+A/6/uQGe89Ynr
I3YnuvxOQfCWnR/iVngnPJ4qweOxVGe9mcLPiJyH1OO/GVPq4TGn3IpB96PoFMJx
YCAJLAASIEr7bOyQXCfRLQ6LXNbdygv8MbYe2H1aGFvcm+eX2lUCJ9r3pGNJCW6L
FWd0aFX/DxNLmcQ82qHfNW7V5076TtkIOa5Cx+qiTTADddOBa2RFtqF9Y1IpTfT0
jKtio/OM3NPwSdsHavlGeywb5ii8rXmK2S/ODyBYUDbm/OrFzsTbR6MhsWf29674
8HaX6GFH5UTbqJIaGZc35XozbJcd7MsYhrunKVldvOn1fzQjQFrvxzdSmJ6jQZIG
UP2+m57GDEKkBNGEkeGlhu6PnbJ0VkQTyNRbJ3VSXxmMuQIti1ufF3M0ZDgIPBmQ
3NPnJubZo7h08+VvhURxI8adRShUs6qkgiPyk6Ta6ZS3EVDRNIENfbhwVYgCX4lJ
eBqglOaa7VNrh6g9Ek/8Yl8OG3+ui975G95Rya0k6Skwl7osSKMFODBNcBKk7hYu
MbJ7HTBTievPANUZFcO4tlF9dvf7eGeZ+PKCQqF/l5HoJwF+c/YyjgGPG1PCCU5A
Bldg9R+N55I4vTPGNzaNZ4ecacSv1XLaMLCFT4nEIOMZOB9IR75DKTFXILya6U2e
39IzAM9FHmtl/fJgcSwcjlfKIAGmCP4jLblogKRzvJ5PPP2xjxvz5AO87Y2sBYXc
hhy5VReTEc3XNr1DHFfNtck0/UuXw2TcgWJBSEfyF4h3vz0HFEJnXQwgTnDa6XBm
W5Tyu2pCUUfA4InJqf95KSvYrPZKVxYdw+V8I1PA/S0/zmYY2J04P3FE6QinIGM+
uOkC6NsipCbbEyPLgtGbnxZVxY2zkIjqXS0Og4cAT/GLPO+gEdtd+7PntuGbZwsI
vsAGGBpyAPFsANTVuLyqggZWMeNO8fmun9JGb9BTduQqf1eCro8RcUaIdZ4QZYbe
FlgZkUeSJosRfLPAFI27jXxdhS9RlrdzqI8MB6py26LFEkf/mtd31rAXzzpGJvpZ
fjL9+q3XEtvBLYTYPInUkOxFThS38RbPXfxIPyu2zOgLrYOJup4f40vJADuNcwVF
QmrKfBxxYUJUJ1oIaHa65H17ArdvJz5qifwmOmxDDApcwqiytqxlXvuqPwccPaYt
tPmgMksEfdygeF4GwAv/RIqsgoAJ5aF9YAJyqWYD55I0gTV7lb6YzRya73H9rncE
A7KjagFANGF8VFSna6Zj76OaFaHet06j0rqppxtXF4K96jmb6KiXGh2nOeFVChJ6
KRkanAfUABzXG3Q0eOo4Irav5mL3vovnoAlvaFd5FAaqWg7n2VUw0QtZEAgYJXBc
qZuc4ouZDGt8Wg+8SaKgNqcDuKND3dIPLjolVdUmOqnTqXvBf0LKHzY+NINDhlBi
FgM3CRIdj35TSkyVfsO/Mnl0TJZCv07TBgmrIFaoKBmxXqwwpNOgRvYoud9N7NpL
WAZHOSjhCU6L5kMBLXzEv4yrfFCjSAFJKa75NzkESawbLKUFO6XSlI++vJuqDByH
NEieGBB6H9PIifxK+S3OBhZ/ZqOc11P06XAfF1mFesrS5DrSuWUVOlzYDvVaRS2H
UQ48TsIH9Wc4lCMqsVwWzB2cvmme7ngYXBAkS2V2HkwGwn8e4N2yAkyEIHwM25VY
wDl7sxKCDhGsNase9aISQHlLcxdSedvTqjb8o/MS+LBfMFKTT1TNBRo9NrZ3613S
MfxMyoThvRgDbP2W1mMxEG6PHDMaW0nHMsQVezsoVzgmJFlDLbc2UwE2vI3JUhUa
hay0A4GEtMzbj2ufTfEie3n9m23T7k7j+GGqFJ1voCZP2qgiOHKlKPEatpY3LLg4
03uTX2v90NapX3xwHIvrbNYZJwoY9bp2CHl5dZvvwEnyl0X54PvI/sRaGZqAgPV9
4uGV1JzOQfHgoRUFlnaQ30oo5i1JBEjuBqmBwzBya/ifDdvjRCGa+pEaAckUh0fL
O/BGJRDF6ZUXNGXGCxBQ3tNOHdwF+EGVfX5dYabTJHNMr8ui381inARotB9K+fa0
k1h6NchuOSvev4K1ySvz18+zj7pHoBWxBtSdjEgw4kM1049NT/hO4enfd4Qj5R1n
4HUV+x+cbP53ZIdBhSKKv4hWChscm2s9gq4Su3cC6ihHH6Nb4qBqvYWQ0XP4x3H+
VNt50BBY08oODgi9jb9dPLySQN7LT7DprBXiLJybBYHSGDeTF5etMXXz/O/S05tB
pjbduttwHSu4t0jzaCEVzqRLhaVDWX8kFR7Q8YBpvEZHNwdVNTd2MAUxzjGAN28V
GWDZT6u37SnBldbjtayd2i4pnEczjRl5t+foicOlRtWHD2mT2n3KdhNvHhydQa2r
PHsmp+gpY3ZqTWYgdjpKJaa8HYrkPKDIRC/BjvC1DhH9LFD5W0sqvPnbVwhGljIL
9adv3u5Cm0NpPmOqECDn1oRSWeFSAHUJs13hFLKOsK69TwEre1vE9YgdHLDFcAHw
3RjNN5xzBzHSUVrQabE67XbLT3yh7l2fYq7zbxE8+qYd/rImoiT5zXuC5psSHn+v
VCiH18t+brRE7qcYVCIofFD+phMLjUWx4TSy8O0kRs2JsfTpYK1aObxEetuamixo
i00CqGn/4nZXIG7zAndreOUAgZLlwkYyHkcunIH6+H1XDzFfLHj7Do3dA4AQfr+e
J1hrDkpRZjvA6OBu7TMhupJfFgBpLmEeEFXvv3Dq5aqEZNWGiWop/lZ/1ohIfxn2
HJ4ip+xFNtgtoRig4kGiDvQ2r6zb0BB9p497yHHKw04aqvqcblWbsOhql9nTx1th
Jn+JB/gIUEwqIEJI5uED1KEo8zE2rkWO4WcyVL0spWMN29Y7osiNezMY14btrv5L
2zUZOISDeHHi8kNJ9SWgvyTioXvvp+6anR2I5g0WVVNsS+rSiLhwaTVrbvcRU9u9
tf0sO+kE5oPB1HsiUxQYRSNngTMsY4H+GR7X69XTLBdFJR1iuVPgL0sbFxz5sVvw
W9o8Sm6nEtREh80tNM700uuN4nnoICUwbU3GlhgklhyixVHE4ox8gDMEydGS+jPk
sZaBaWFwMQ20Usj/IK2EyBqgGM8MiPwONpXr3dh2vOu8XhiKJNkqZ1oFvPCZocv/
Ev4ir9o9coFG3EALemldc7hv6iAPheooKGyerjBcorw1ufKRTqaWdKEKAdS6SNi+
hP4WmwZh2QLFO6M5SjylVfphNvRQYku/QdiQhNywFg9wvIOlr+KURykz6N/VaRtK
rIy4A93rPskrlHfGTCNlvE9GgljfZESN8ktPv7FLY61AFVk42DQI35QiNsNtcHL0
qOFhpBfUtH5eQtWYyQemEjrzqR71k4OE04QJFMfi6RvJ9f0qOQoipPCMot9N93Hi
++Ij5EzkQhOP4USJWve8R2GfAB6RUb+tB7gRgCPZiWis7Eb7Pjz/Ikwu5PgesQTn
XxaaZoHqqW3SiOTL8F6VsytDUxyT5BJhlJqSHIfO5PCOT6QVIUQfE93VrV+1KP9L
qtpcHXy1ap5wvMdRx1egjzhP0EyvLD1SxA5/zkVmscA84RvqZxwZT2Ga+Vf/Gmta
qAsry44HJXwQwuypkBm3DEB8g+oXMz5MPddKcezZ9rE5tYOiOTelXLYqSIBjAAkq
l8jQtLCyXdQMGTv+wYCAxzhQxWfPNDXtkA4yuOYYISz99hbM57vpshL6y7OYVV7e
hdYGTlJ5Ytsxck187UuQ8xICFq8dEfCL/ApRsNRcX5BxOI2NUgyL+4iTHApJ+a2D
senaKsScc0tqpT3yBN8fwrPyaAL/QNY+vE1lm22wBGiOaZtpheCedsHAJcLfx7vZ
E15fJCBnXB41ofkxo7lh8R8lgWi9ngbXfWmEN0W9Q4WDROLBT8FVFY72mMqAUhP9
FGK2RWGxsmkxGDQwcwO2nBO43iBXbPZE+dOvtK3uSP1LOWmAgh5S/sCM6KvPU260
ocSlhq4hgK24tFD882VChweod2Hhmq6GXIXq2iJjOqWrdFIRRtNtWr71ny6F09hq
7jGmfWuiwQLt5H1e32Y26sRqhSL+M79v4hmX594MryyQHsQaZurNnf21CIb0RsIR
eZdYpWYrCo6ULCVOd58b5cydlG52DgCYyq3BasYy8HseZS+i1VnnOHnkiNsHT/9E
o+Ok+42vqzU1e7R6kx4H13yGxiIQYVH/YhOFGIpaDYXG/uOwdFVF/DcKajnJkRIx
Eo+XaB0XCSjfyrQKFh792uIxj0rpSEC8uNvXw90UJ6zd4FQnulfFP6hOhTgZat7p
cK2PLpYK6BMWMxKxYYwkTxwnAFlWr0lRhsQHQBI6oLayvO30iGOSEY3yW1dqggO4
7hdNcwrefVjPNkX+GZaxyEJP8xLPQzyPIyiV3ECbBErjxt09UeX2EdHOBNZUGdw8
sMd14jRykO4u5ONf2ynUOR151zPkHKemExasEiGLc594yaZVQwVogoR1YrGT4aI/
DJYsEOBSDOV7tHgtv5oPWjXENEggNBcuSq7jY4ozJWbc4h3ahUlKarlUlQEdO5eU
k8ACu0dExlKlPUWOHBaSdvBQoJWgFsPTwSlxXnqAjY4CG7GLUfDKIorJpz+azMgk
WJxPZ+ZDWtDXn9ZcEvv8vtPKSH1YiEqFmIDcABOluNraU5FaLr0dfkablnHtBiN2
5Nz2wAc/AVB38FbyGFh8KKwJcsjY/roohw42trcNgO/1HHJATKgT2nZtJb1d70Af
OFj/5h5Lq2KwllIztC133TqVwnTrT3EnfSOdNbAGpUXOuVSSBYR8fEENBTNd5sf6
XWiKrBheSaplmtz+NsaK1Mt9iGeht5eJpvQBfAzxtx1w12K4NvmAGwdi6aDJHztO
kwXbue5lAES74Up5RGWnm7AX7YQB5sEhnv4ZZLDh4qCbTYAFbIK4bBk3n8jyQn/n
LcxdkgTahG3XXhXHRboS4nn3hC+tOKPcG1Jyl282vYWR1qD4FyQM4x+x1RJcz02d
7qVlrZLoadcMNNTJv2xIPo8pDSDuCmkI3Pc1JEpUAwwjrf7TWD76wNHMP3nYKoNb
fjqN6OOXCWJtoMG02Tvq42bf30BTYMXHDEQ51Cp19x2vbj1tHsStTiJ0XbjFiEQg
ZcbYEbHWDSkSAx5aT75upgrdAeFdI8lxCtTP62rjxcJGFSUFjyUk/2mZL2BAdd20
UboFD3KZ/twtr49JRArn6uCXNKZH/8ojLFCcFCtMwv25P4JwdG/yPtgfmjkBslw/
jlaoIBLUFasEuAhIlzIkuqedYBmZsZ9gEZuOizSg9RCI0313udl0l621vQJVpXOq
86qmD4TqyOEtGOPo+q978e/ErPoGd0IZpCphLHldUWI+JKY+WkgW/cr8gvJ8Pu8s
hGer4st7KHbRIT2DH66ATR7sN7EZsnph65CMfK0yesy+RNKtPQzs3qGsmsVJO+56
b+5nfCw7jtyOcY5luWUKAyTQNIcKZ2a0jfNA8RMkM7NW8uOXM8tz04hLERgjaemo
/ixDpRRgbKG/9d0+aDCevgm8D3/HhuOjfTsw7sj9g8UFfnJhIbbzbbh14DeXfQib
FlKZWfPkEtivvXbpFWwumAXKBDohEmhLwlFO5DUSo3Rn14XAa4QfxginHlXgBRtP
isU9kkvjbow80ywMwyz2XCfwJErZR3LNxXoj19e2IRzzyqrVbMFZwpowdQ4AN5oW
qeZTKXNu9xB/HJ6ba/gApmmWgT64I2APvYwCkCl/GsyteMVd2KOuU5AVwSxsYPjU
wW9OiCEYF1d+MnlXsqa/fO57LchmwXyThRD4Dwah5JjN7EV6nOSfQmlhYVt7uYyK
p5oUV3HLbvLFyQw267qCWqK3VtQV810JNTRJKVEEZKqCiIS3UQxUR1xIwL+uBGET
gBXri+GBELZAnLCYe5QBF/nJ0nWpBxE5COioAt6FbXsojeVA6Kcx1KziGGnYy2M3
JOvH3Nobophkaz7j/8OJdI1xhJuNv6+mpjFG8aCUtinS1PdvdDrU4c7oT5fBWGi+
dz8mc26Ee7KGrck8YWGaHdcyqux+UI9HwGsC1JX6i56RHsAZ7KyKnmS7lZmR04fN
yStmk5jFdFzqoI3vORx9hue9qVx1UZWi+EHSwS2edmq4WYeDzYkCMUAgFAkmXrx5
5de5a5bzEKbFbHyCes3ZZmUzCcKmgZ3EofLPUjsWNpL/73AnOpzkzyulDpDmiq1s
fhPKFds3oh/OaL5l/1eUKESX6VTkDPDPnG8dhD88i+oumJO8961Dc774YztQjYGZ
f4hMY/h2cHCS4RAjXMBusPgX6kWXyg/h//9nw6gSR7E05BGXEwJoMgdE0wb/dgfn
ThEBLKMLxDzLcNtxM279aQxquTFFNgfazeEOiFUlnvGGjg/PAJeIua9z+FyJewzm
T6rd7aiF+JjnQXiPL+cKpuWQ7nCY22zZkVNhf0pwNgxJ4EFw4J3HfQfJm2C701L4
13U+Vv7+xFcn8H1Lvbpp1CMoFS6fnmKTjbNF72RCkY0IM2eF1t0auQYxU+iJ/Ugj
wT+LXZbK8RdtCAXa7G75p1AKkJO1tqguE+bE8R/8g315wJh9vtM9qAase4GduHfF
ZMVO9iKCZM2VSJQxBRePbmj3836bx14wmj1Hk30Krfl5PosxGxgbntMdzUHQEvJ/
5GvEYp2S5SmL4NUiF0i29kfBQsZvw0SQED/pvZkV7cX/lnseV72cnc2Ws4wFxRPj
xe4e6vok4zCe8DzsgN3SbZtCdNm42pIwty/nsMZ1yUbWOFrFok5Shg3p8uUmcDs1
XbRtFWV0tp6mtHmy1vkiIzakWH7G7SWly6hPqtN3oo7pdFq2i4Rs+uPlJtBdbHqt
vTkcdESZQpWtpBl8Bi/qGXeTQuLYqHnlHMIGfo+QVw9kNccYtRL5f/UjIgQSYQjk
oqF4QLcAxecjD/jK+ECIsx6WgF5vP0Xi7bGEojw+Gj6S4Exz6ttTjbSlgbc9uLgX
UHmtgWQy8WqbIrrfOvL8rxL7V8/H3rD8tSvDtEKvSIdzbVephOYaJkc66tkGpgBY
CH71nT4i3hkYvRAPsaEz+hUzoj6QwwsU7ixgoIfxBq6ZHKX022amKxacCLWojYM4
tCSd68cB0rd4cVW3nICGmbxqvXTpwkGMUbrFbiD1l4uk++V1QUQpGxw8D0w0fHep
PMt4iB/OPd9LH3cokIf7zwbjk2wW9DAjjOLn6smRGIDfr1DvEvYRDP+gmmnC1Bk5
SpaqKJHTtZTIJdWAQdgJ9CfpPinnR5EtksBTex1+AO84hoNF59uHJOV7Vt+QgdhN
665YFdGnKmTe64iSb4JKMZ9e6PV6Z+djqQrG0ReQ5UuxKuUDrsWyAOmJ8k1TobG7
uGch8F+vTVZf6uKk2pT3tt35lU70Osn2VZf2i5MYqM0Qh/PesXH1qoejnphHFhYV
IvDNrwieu9ns2eQRoDzZ46JJx70JMbV/0PNpBUTGLc19yRFG6gK276d+WnyvS7or
vY43mR4e80Pkus8zZZKdJq9A1F1CpEiR2a3dnUtjsuSxt+YMJIzH1Ir7dpsH8QVZ
HoVOqkSy+qOwbJEt96HBxv+di8SuIic6Qi2+BrImBr+KBiwvRM7GBmsXRsoJqAVO
jfAJRDkU2AqdNL0OMGpf02a4AG0aney4nBtSlgMOS4UTR9K627KmMhJi1eRFXR1G
601l1XPIEGWii8lp39Jel4SdS+kNt8A8GTwAMQRaUYg2sZe0H+xWU0zIo628tSQi
wJoHVmGzw0ZRdRM5ITXZqVhQHnrZmpC5/vfuo1PHFSZRibUDQ8IB6aguZFF8PrRO
eNk8UGqr4jXMjL84pxTBgAl2sohRtAIQEFGuWjnj03SFpocA8AimKSNNo9U3zhfp
SxG/hrhhyxtfAAvJ3abYOwbDpW1WE8r5xAq028nmvKl9qkzKbV/GIkLtR/1w6rLV
6TlZHs/8aVm0SxktR79Ov90+L3+7jx0zthQ4JPCmqsoCRLhi9WNsNp6v6l0kmH66
xzL8D8a0vHU36Sk8rskaeELhKnLpslgPSDSIphwFRhWHDPgLLAOTZGxjLhfGLePW
Ej0PeKjhd+jHZbtcNN4tIfsvfyX2uTwWDunl+hKXhu0nzy9la3UagfIy/SA+RXF8
5aT2L8J/QJB4fS4uwq15rn5IjaHvOAkpNI956DuW6wq32/rlXCXAbdU5kApuVdNr
LGiPmx8EISPRh3aKumTJQaBelNC1ALL/7IzXcrKDsH8NDcVY//tyjJUqzQoYPbpy
hwb0HiIxW/JyEwJ0W8PhXQApZwwxI6TdkSiWHoi03EuajxlBLKSuUN8tyyWmTI23
W1tc5YJMSMIihN8W+XKHHsTmCVUFvEUl2+Y90B3eLUzZS7yJ6eu26u2MJ2Rz1Dto
mzOirE+yOaFEky10adUGRSYRiKcsRxD+h9ihdU7bNgrat6o5CJw5OZUJlDAqwnqo
Ys98AdVrqi6kKt2GFVehG8vyFfaCYsuDlHjYXgEIFm6ZaI2/Wllu+OLHYRfIu+sG
IToYrT0DxCpV68VP8r5vH2CnP3Euwj/UbKAW1JE55YqWQFuwMF2w+vhO6CKmEi5B
18PmB/x187l8MvdIJUDI3LgmxA/O7nwbjpw0oHVf2eUYy1zwgNisjjp9vOH37L/3
p2WhQfNiI2Cr904Qdv7tG7Hx5U8WglfNJL0KUrFLcZdtJCWHf4RaXV2OtT1lYS7h
dKMx/eVawh3o4AHdtIFegUXSyxwylgnklNyvfoWfgRjdRXzxrqTyIo08lGvWjqQ1
7AjyRuoOPwoFnYsE/IZHjfHc1vLbJ4V98XqwV/nMEYYrNzQ4hjyG+wO8xY4wVI+J
O1P22tVsfAb1k3c7YyhABaKIdGQp03wFfJfhcifIRzvVNY49OwIYPdSgpJTDh1RG
0VVKqxXk8GPfqVt2dvzhl7dpnHpSl27b/AWTCaKdFoTh/ifM6RRyNuiE967GbglL
jgCwK37yiP5fFd0dN2M//8npOEEGcPsQ3VHjyp8e+W8EJzNYpW0s4WVQ6fNuwndL
Ul7K5MsBkdFyzn6BvRAIgZMgWBkmEvFFM5srZ/THA3OeP+W5KwzzaH4tFA1XSDmX
e/g09YrPgpP0DHZjJdE09qO2bR4XRRHejyvDUt/srCPSVwFcK13WtcoJgTeJTdGS
qNWC9rwG04FqGudeBvM5KvQMiGquxnsNq6cquRSF7gtYgYBPKiTJ0VqxehPBT/XB
Q5hmRbhKwvp2OOkup4DCCcGhJYFSoPzruaVkylEI3itx6VF32skRi0JW+BWftf6Q
1hcnngXcVsyoIdPyRU08r5fpdPo7tnjpFSE+HGPeQuS7uHZz42Uzg+T6huGQH3Ba
H+0dcE13wZVus1n2iWrSSwzbA72OtsroPUIOrmqgtTZWNSd0n7jaKCsC8YOWhwVi
bCGQXxYPlhkQ7IBYivOIGJduC86ifFsAx44fZJcHh99HWQxUDqS67anqYqONsd2y
RECO88TibX4MtuaUSVZGrdGDnarCFsgqTry8wTcD8Ty18K36IqPhY+BD4x5TBsdt
HqYwF2A7VHd2YTv1L7/tDPSgDiuf+wNaXpPK8EfrJvK0VQOQLDaQxlh1qxQIKMe0
u7eBtFqBVMSoxIoHBF06oUZ1nhXuEeSTunHG7aoYc9DllN9RUAad2ui55VtrA0G2
n4i31L4NWsWcmyE2i9byDsT+a3MnifPP9z9sZSCWdsHxUYsGSdPswWa9pqaEZ8je
/KbycJVEEAmK3wdtacIBhjWodOuJMfXcKRwsx13PzJgMSix+BuqJZLQr1ErDUWOP
ZRcqNahdgSQkCkOxogrZBciddZMI9pPUJ89VZjWvJZFMzioptdQ76hmf5Wjj30YZ
ssQcKXJTAvfQWXlQsPEr0SX0Cwdg3W2lYOG/4NhOUTCjjQU3phib800YIpTUhaPY
iiD2nm0Q/oAWpGsTspdA4Aulaa2O/QqrA8mO07LgOYjfrKQ3W2dhL209vrXlRFIG
LMn3tsiPUz0FvV0wv27yGOuV6XUOtz6mpws68QiEWh/caSnad1x0BwyH3CohWig3
OyRdcsiCfxSokPSoNp8g53iVQ49GAH+ekC35tBozpgJMnKdJbSZWKDeFPlUFsMvS
t6fgvxLgAznW5pAs//c7cCXsUGlkl676bJfC9QvERpF4kH1W49sw6sGfZiT0tbPR
7ljZPzHoxjOJS5BFkCkxWdKRWna1RDjnWDj3KrFVFSyPhKd9aX8WezQE1yk0QDxP
UEe4+VxaGERrRZhrFpb21lFE+DCnS8JacLicalG7KBVqc1BdJW6dVuK7vPNC5jCL
rirJ02NQTggVT0Qb6woGP9BtFIpKEaXEab/AhH/Gp/PGoUm6vm3/19Gm+Vu8PUuf
xxkbQKS88/WT37mo+ygDyHIVr91WpIGb0zLMlRlp/8sIaYzMBt4embmdTYqq9ssC
/S/Wf25wDaq6vAi0eWtLy9LfGHQ0RXMToV+g3phBJC809Cg1GZSDTx+5q49IeP1R
tJRIGdszsI37kfnSwxyxynLwYTE/++3kM6yRMbhURsrJXZGzVsZsJh9MF338VYoy
RWPH7gCYMEf4vEK3cPL5bHsM3q0Au47+AFbowoaGWSYbzXCKl0wSAvSe6BN2mdSm
OM/FesarjbbPv/Vy2sPxeMl9fXjmazEMBMeaBj4rgDbLIbHgTT25wx5C5kFxKYx0
ZlA39dohxzPOaE1xL1D0/zVANdnHmcVis/2orfZWazVCOJWJa02NDTgxtNpvVvLx
6pVtQgZBU/jW9i/FQ7Z57isitXOFC4AHk90DobcCrXTPSVaZkO9bdEopgOFSFOC4
jQ7zANhmvdGukhxnlmEc5fgQOi55sSnuPvqO66kfbzKERAeE+mf/Teg/kIpV2Vs3
vUW3W5djHrCgY9FkVgYxvZSpMVjmf4yMYkgMmZolGqZ+vysdNE7I9gJjk2PUtuKM
QYxDsJCMxcMShusvOZg4qu8p+BKCzVwllB2zyds03+c6Sz2Mr1HO1Nr06tdRNhyH
s/U6t62ZtEnZ1NMuo/i+Q4iAbm6UgV6PFYlGSkfbPMzseSEZCMWbUVRfeFeT69Om
2X4YgnhtBEpRjVZTY7/RQnTU4kwTIRYa6254MrubCBLliCKMjo8RI1iw046VefgB
SdpMhbJBY1p7wYxeWKaVgxAZ/rsQSdXW6RbZFPySiuoW+Uo39Y0sPuRA6ZJYqSDv
bfBb0GPtt0NeiqE0Vix4GuVCz1MJMY7EVT8TwLuJQwK3iP+S7jljr6/XIS7XdlJa
7Tpza/VP+MYqNl9YODs4blGGYrvyr29k50dzKmGqBFNfjk1rMVr0MFSNumxFW8hx
c1m7atClk+bnLN2GFKZWOkRhX2OuPfXcj6FE9Yi0q4n3MuI9xhqD+vcT0RZyr2iN
PjFhfMOWFf640wE77K2t/iH37f7iXUNU1qFuDniscS5ZnZUq666fyk+y2449Aoh+
kQcFFWNRbQlfpRH5tVGZp/fD/8UXx8Ssl9fNZfmJoKyuuYtBTVVrK/u7NCOitsIC
z1PvXuqHykqc4GtaJ1MJbbSBkwVyB3e1kUuiVUtRCynfI+/h9h0tUxlGR6h7odZY
exI67x/MuZv9myn6ap/pjnWuGd2W1v2I8FQEhKB8POGxfJjVl30t5lbxQxWvFH9v
AjSQK6wCG9RNpsvh69O3bjaPmEE9ZIxW11ump7IDFPBdPZI7kxvUe45JdzdI/oKR
UZn4RXRhgieRSd4QHOB+4giJ0GzGZ9tMIM1Kdm420LKYFMTXUdRxesgxfTT4/9pq
cTyLbDM1oLBFCv55WTBdvpcmL76Rm34r35JkD4ya5N8vNZIlqYTGHLLoNiEIfovZ
gx81WGlzTMu5JMccRSt7fxJawt1UBkvVwz6vdYsFt4OQawKSDQNI7u4dck0zjW/M
sdDRhCRT9oT4MLnRrmZ4uIaY62sKH30cGKJErUJPqvvdfOxlYcWmPm2nQ6JuXXra
Q/9Zb0/movhn/xen7NaqlkGsA3twlnU5hU4Oql7DfkvMz+Z19XznOR7ayuEUtAqw
WoJGNjtMEAmErhWewdQsTLu9d4lRQ5vovS9YuKqgdptdO7Zr75h1CDBlpkIVFF40
eFG0qviTJMNxLsZiVbykMOcs6Pf/C8KDTxvJhqRgYQREZM0h6wwpDlR/O79dwsdN
OJU/Z0yZ/El+8+aL/sLdn6jpyvVocnWD2tbf7Cs3BcHDoSsOhAuOCTEbRdDMQPSa
rrvSKkKvfe4zkTy4fdjtN0DGfZAixfRkndPnZtvPbBB06RJg9Jdm3iAhJyy44vIa
dSpUYDjVLvzghpXYDpOySusCn3pJpm3GY6vGyOvZM91JZofd7lQqm5ohX/grWech
wE5dYWO5XztX6AowmQoYngPE+Fhk3eGUiZvSJPIMRb1fxBcQ1CdR58fG/wTQZ4/H
gKAvgFMFSENgNdmLmp8X8G1Fwo1msLMKgcfdEzE9CNUu86xi+lrxUvhJR4qJUtAy
wONI8G7YNBXJL+sRiAjtneqZ+W+rywg9V/0QJEQDEOXGAzzjzxzIxRZyz08MFIMW
6voqOiyajjCfoMHRfm0u5RZr9W1dAXHfbdKJZGP3fHZNctPY2qfkdXJHYdDpYPPN
qPHYfrzTbm5zzgCVl1GS5or3RVolcZdigm4HpqN1ztD3f6clkwTRpd6SwBU4YIP5
cA6ydALXRxqYaEo+xXq0zK2CC8T5GFOw3HzTY4SrRId7PTd4BhrdzeBIms9lvgDw
VhOkJc9MVk/IzyRHuHbqOSGK0y4pNyqEMkvMx+1mA3R/MicLX27UyibGR0s66l5L
9VmR/ntpCwNZ6kbObzBF92P2B9BcmZH6s+BkUChz1vbXVHRWCpODQRyUucWZLX/p
wQyZleNPgzs02duCntdvsvKvRUdt/jnZkKzwr8b3xUvLTdUgmMuum/ZnvB6/c1T7
QDy946DCo1W8Gie1WkjbPNfLlNECW2ByRdmeRWpJ7Kc8qYTBFqGnIF8D3LBoWlwy
5l2RM9JAN/Q0jE/zgKl8/Vd9mYfCU3/kXUkhjM5CFXRcgUJ1RHKw2qtOloptI5zB
/Ld+DIgC5sLBMm9BmcV5MpWrgqVjgJVzHgjyokaKYL9EBqYRS/p+ggDToZtgu2SF
JOpWndwHdPZx9dN6pWqX+4e2sFe2Yg7Erri5IC/M3w8H6dKmVIG1xqpBv9LjCUSx
ig0o3YqBkeH4Y4dpRfFNYttkkQj+mIInhRuRtQbPudQ53wcWsxbwBstto5EXgiGG
aat7CSu25477X49iM68xOh5QUY8n/8/7YFuUg2Aa99qQVAa8VjiN5eyM1WiVqmx4
1Vkv0RGl6lDjp+yC3OjtKpJcXlJZieNcqfStf2o5YmybLK7au+7oZRMhW10jB95n
7HUuC+hB6fr44s64n0bQsfmnBQSiwZnRIrHz31AtUxlTDhKFWU+zg/4sSo45ymsZ
eGdektMSccqvwge3pBazvIXSdrTVByom2Hg5wz89IdKPp3yfYO5E3/wKLTaR41dp
9mzr5qmsKziLuGqKC6KaRygrbm/UJF7sVOP6VGBwiR6EQPxkucfRSfU+wGRiuljJ
U2W4xk3zdF+I8TN0zqnifmqsZLjP05rY4w+MTUiorWaVm+GH78rogFvC8lZbQ2sJ
/iHROx/QNGTqislPxKvc1x2NmGDjull5EQJwcURkxCirV4uWKDVzuYox9iX1hKTc
uFYMCbozS7nCEc4NBJ0lSNA6JLdNWV4GCSWgNmEgMEn/buCe39R2w3IpcduPtPSn
ancN/3CtneiJthkjt3iXWnIgK1fs0uzNmTEGZZWg8jAjAc/095KgwQ3haaVaoVFU
fwqpT6PV4XQEDI1R3Juki+VcSLgvfnKgsVh9FJRjIhSWnvNoDJJ3XSU2SmNy2CZ+
zXLAGklD0K6ss2V1jHs1KRmZkKSetEpTD/kZjV0V18bNDmp7DoiGciDFvl8UXHDO
/n4m1N2Fwxfo1m07+hUOV7ztg+dgp3+sVpcUOvHL7vlFU2o72QJsOqgeq1dITI8t
O27xBdTtxO0yiUPY9bgoc5Sx+4C9gFmckMfEJiS0qQfLLIbqhNX1CeFsyWEhLNv2
7rhc2Roma6wwHtB7ut2L2sKO6KFJOj9u2xYcsyyul437Bj5g/Kact3WfuQiB2ukn
Nq2cS2z2UqGcSXDU+PKzCXny7FMUssAYc2jCuiz2uj75BdxM1JHsBxJsVGNA3Rl8
ERO/nktw0K5d/fC55Hhhs7uhXks+ZrIpZTeiV4QbiA5ck1FBcdUp0ZJdO3sRi4Dm
0jS/4ic5K+xEGBLi9K7bRtHUg6sm9DP56PfLOv4Bxf173XDaTl8EkcMhMqtvdXU1
qFMsttONPE+xx2AgpxbqWkCl92FLvUc0KmbLLck384D4peQIGWkCXwIC8jxIQzUq
PXo8pzmxCHof/cBBZy+JRZGN9VONIqp9pKiqvEdENHq/hJ8ttz6Z7BuJvbuF3Wem
jm7+K2QM2IpFStTYkH03RbSxMa1Zy4/sJ2tmVpmh4lBNobwtCaUir5ykfvob6JtV
CgiC/ttodkn5z5WswoRCArrK2OU+CWrb+tZ+tcny+x5gqY6l10E6l91Nr9a5vNE/
p4WZlTWqY6NElJYFeer3xR7AcpfwaC1j+J/e1j0V6aiSxQt511d6N7ErPtEKbfnY
6Jlj9+mFdU8PEmuMeeH9BjtcT+FE3rL+zIGFFZR/l/fv4ssUucexq21XOurYCgew
8gPxEQAHAm3esOUF++sYPWfE1gEat7E4MYywkDuUBx+4NBUKSlO1IEtpGOAnvRyv
Chqm+TXrhAzP/JsUIT1NBVIxdmnv9HbsbxvmBTDrPW0cVRKjZGYc4s+mKGFF3lig
zEwLQNya8jqppHUgI6Q7l5QbV03/9EZNxSfqZZgMrX6ECp2dBFUGPWRDX3J63XZC
i9VaM/z7W7qsESWdRkNB0yBr4e+ibIJ5QscrnJXYztVPCyqyNfYHWxDegFe1LK2Z
Tp1bmOTAHlBoBTm8DWudN7XUZ6V9U3TPAOpJxdN9ZfZ9D4TxHP7NkqjveP6ulHLG
e/tv3ROlyZ4tyE0rCPqufzI0BzVpjdIxkv4OT8Ey76RNgumpoo9Y5hyiPPOcRUj0
F0Hnhfq242QYNSHLZfMR6fXNaQdcP1AqybMVWrtP7E6uQzzGrs9usXVykwgKvQwS
D6gOLCVZYMxgDg0VwYa3TPwR+Q5tAhsXtEUWsif5v3KDXlOLnk4sB1ATVel2LxlJ
7zzLWt8uMyNm9f4caxjzMl7BrWDSmykN8JuGcSLDt/j64SYw6CC5DJ9ffvX/Xcez
CFHEAuYhr4uuu5j3uxemURHLiSzk5TVaEVv/QjP1M3iuuwZ2zgdKYEX4YWJKwICh
aItnN4mTjPSvOjqJdV79+yeRWjz27Bux87qIP+MLY16azL30MvW9B1d6v7169jsx
ylT/HO6CcLbFxqkuILPFq2WmbCtBIBg3rH9Nh3WihnNGDaGZu4VArFNsLm9fZ7PT
0kDSXjFXqzd2A/TAiO7XnrdCbmYSEA/owXKHmWUSAzN7/uZPmVxtqvYn5WbVVdyt
MkiU1SZr+CU1ncNFPa7J7mVgSdFgCsM0H+HD0b2UtyCIxV5Lg3MHNchL25UnQtn9
MvOdiAEJyLG3ozLk9AAqMZg0aiD/HjilR+XTd3nTLB1rnqX3/yk+nJzLY7HEK1AG
Y6jct16dku49XbtM5wI9fNQHJGI8/q9Ju+tlAnLvvvgsOcqu4rvJdQhRcsn92LQd
uLY1fKrex+PNEkGgoVZp/DchFZRZUGfoEnT4c28pk4d6TPVHKWmL91IXW0emCM6h
yGVg37391r8EEIzpIdjYBVCuNgSxGS57VdsEsqvp5z4eWN6E2rvmcCZZ+xXzh96s
307eAq39wX7SkNwSlNZYdRcKzPRtdSgPPiKARWdnedJGJRqsRVeZxHMoNbStgFCi
eIRFnJbuP70DbJbtgwBmOSRL7bLEm62qe6/seJNPlpiB1Vhe7jpbttTsDrLUQ3Qi
ns07nhxss4WsUrNgsKcFP0E6rPmHQ7B7IrXsb9UWaKPvS2McLLRI4iiKwXJwEsC2
NwP3Te4pNjcS5Kn2ufNbh2BHvFlmTPMUbQzTeoca8krx81DpnNI+yQ9sZPduHQQj
QZ9hd2ufA0liMqgp9qdgsBvm/Q81/wA+xfCAzfmatlZ0SVDdy2I92q38khGB4zSF
gscN+vUwdzOgv2xHmOOQQs5P03ruP3mP5s+5Q0x1HPO4Z4X26X653gTt4QTaZju/
703H5I3Q5m1c/5thPQajPzKoRpjYLDciWF4sIsuinmNXVJoNPJgRWsKV85TGXCPY
s1PrJ2W5FevlOzwcz3Cn7iAeresUtPxzsrW0t7G+me19Gz/E7ZoKmFpJ685cI9vo
JS2fJXssm5hj9QHn9PsFqAEmYi8CmSAiv0Abp6ZSmf0K61welFlzMkc0g7hZr5Mx
k+DzdnW/iDsAHZ/WEroqnWcKS54zDEUFh2dvgkeLQUexUtpT9yl8JvehMFPZ4jk6
x2xDbzGuAfY/nvaJI4TnoEy5kqFgkYupeuYsryv0qXhZt7HUdh09fuHfN7VUsgbH
bYg6FNAp5k4Zhq7m+DZdZcZCGjG95x2UJeAlmv1kOusTzVrD/I8cmXfNnWxdqEIu
Xv5SXwuCTpUgsFcrxbSwNOAs1GHVHZ52JG3WlUxeXgPVYggf8iwBgDRrZM7O6FEy
rkdL5Y3XfaPiUc+JKiO6n4ihGPWzYh9tE4QUORI5yEoq+91FKEzmcjCV65K57Vix
+/NuTknLKNKt3ixQWdaE9n91zK61LtTdEiYUhbSO1OtaR2RgAxh8L2W+UeQ19jZW
IufEYYPbgDwqjIy+CZX40uOykXSjp9xHWmFpXuf+qtucHYIFwm66ZrQWidh7hBlc
k5fKeSrzjQoeb85ztliZwkpSQnRHqtl9L9+z2b6gT2LTCF8MRHGLdmUF6ACykMqN
XDktbAxApSf8YpkFjKKpCVxzEh66gv8ogsmmbNiZvHZQEMbYeXtQkbJ02kMZXqLe
a+DflpP9qhDfKo4WpXz8xtYVfxWQvj7XHnYpA/cBoyJLmePjs6+FuHkV1qcPyml0
lchPYeosUiT7378LoG0cnC6LR4GaZf1YYGeOT2EsDid62cKJ28yXSeHuQzgJgAo1
tibfzuDX8QByEbe3uCoKkzCuHI9MW81t1tlysjA2iIjinswpLQJYzp8Y7Hp0OPZz
mSve5KRRXtlmdtBK/ztGiDogPSaQkjuOm8ev3f7szfMELg2aRCuun/TOCtpfwSR4
Rv5JG0+GrwnK8mXQ1q7HL25NYBvOAlKflzptrjQLjSmHNNPk+46ZTqKjBkW+27l7
VsgHnoIvzMQmqyJOZrFh6FOmQfcn79CUILtlqo5E20YKfSBYca/Be3jMnq8e1wJr
UreagzOpO202K+RKXasktJ22VH1ojVj7fkhBiwkKcBpstfmDDZlUfRRloRz8uh0U
qYk7KtwRroQKNeB7sx4yNvcLo8YAxxJEuMfSRVFVrx82EwLpPzJEx4xlYVAScXEH
CWlRFTYZ7KYgjCzNR4RbKt5vCeR5Kj8yFHqhayJt/LkSvrQzRgYLxwxJ2STN+Do4
IOjmpxxdy3rPOKPCx5SK5kYtZKKYOimeFGaM+mNeT8wYfuS8S6UxeOtYKtfkcZtZ
Ie8Q/BiUfP93zkgd5WlzoEtFSXwFVuI45gI6wTOp2Bhe0BtcTVpVxzEXsqQt+HrV
JqoOBQuq4sTcW6IBl1ngW56wK0Coe6BmGNUmfD4ClmRs5tOK3zDjUdqRAUoX+YtV
QIStIweLurj+ZNCwHDkhmmG6mAdocXVw9KLS7bA9AWWHq+L+Awzj2pFcS5Y9ktfi
Wfnv/KSUuBrxWZ4D5E7Gr1ww5mlMTvqpdvSNeIA9k+jD6u5qelD2i8sV5oYzk7/D
WR2WIZYW2/ifnnYlt5CzkGkVCmsXLuzAwa8+38ThvMiqaxQUzPZg0VwQkwuWo0NG
npuRpCAJXttYWVu5XNU/i463wIfryJfNUt5CTTT0nb6bQS5mvUM0lBt0aPceF0fD
Y4mahYifD1uMzwqV7HgZT6qFgZLCnrns5FFifSI9adJTx3p7MBfLxAgcwnnjEnHJ
KdDTiI6yXwRszdKiiYKiDbmTsZJZs92Xxbofz5C2JT5s/NqaCufrzgDuq9Cq7qoa
TslNrsVZVXU9PcnH5wKK8UP4Fzd4EYYH+OXkZ/D0B36OXVqsGjnyeT45YLbkZYP5
ZoDS/IWpvERmo93f1LeJqwPt3eCE8/DhIPxCEkVLTWQqhPm/HYMadr8X2brGfj07
x8SDW2vP6OHjatWIu6KERpB+EsVzETtg3dPRT84SU3/p80SXu9IYLxK1ldC51aV4
+t541rDm7yBncucgrr+5rMzwR9xI0/yKFBfAkr96BFwOzG6Ii9JR3pVcm0CkujXX
DASO+KTRbhREqGQfrvXoIEUWZJL1IGNlMKaTIRCkh+cQWr42pycdFhYqiAB0HJTM
akWQf0nmC6YnmPJWDDsieIWNVJbazrSB9DqO9XKle2ceiSbNxtC30n24zn1/4Ht/
FesZZ1rfWNRr7lUaPg/6dB29X5MZAZGZk8nzaQhl3rR6X69+5UzGbPfzqkz91SUj
xjVRHNQO74dVkZdW7UiJ+FbI9mutTbtu+VEnvJmv0nW152d+F2wIophoFNP5UoVN
/tiUIa52HLmoQkSWjfaBDkODd7PNBmVmPT63gIvwB5qBg6PtGleNsXGn2H12uzyZ
lq1aJu3U0HnlUqWO566kdgps7Jky8vs4qIOnQ/kLC8CrLpli6TcvqlDam5ORGKUb
Ad7UFj6Cox7UVclzExay+5ZGy2WE6dpORGO4/5N2A+u5il0kS4snZTUf9CcB6AN6
wsvsBWPTJbF8ARJ+2jX3t/poJNG0Gb10FojqODBGMqZzQcSEICPRx9tK6gQmiiBV
6BXHeWzgVgx287kq9SY0lDJURlFPX4ECwjB34Fo5F6ol0+cytrxpxQcqAmiT++D0
OYG5GwiVkHbHDRpRov6dvs0vjDz21W2ppOi+p/D45W3zzl+DfQlGII62+Bm/o6g3
+jFZ/lYl6Kuzxe4Je9D55VxQbQYpdJ4jw/aP+eSRSGbZH2Nk/DEloUQQyTvFfvFu
bhYxIYaaq+jpGEjn9jOm/DKk1YhPE8UE99QuA17NmHdwerBMEisIWT7pQAxWWYgk
EL3aQO1BzVgqo9aNkW/6ZQvoq+DGFLfkiqZjVn6Eju/8rxXz4gIPsUaypZVDHf70
R6NNCjY6Fz548i5q2xXbKeDd6GmkEgEgxKasWL6D34UTywBRozN7+Svq4JKxwgIF
81AqdftRmZxssuLPjx8n99mb70yUTBEDN+eJY9gzsMEKJkD2qZ9CpKdojxaV/rF4
Qhv5mdXBMB4+IxCH8tZta6K3pkfPpSTTDUe4d9vXzk9fAwrKooZCLmI6xupaKbIq
qY8/AWHKUlHKPMoF7B51fWDkWg6qkBga163go+dUmBijX25P/e6R2Vv8pfgwqzPA
X+TlXGRxxFT57HpR7H04Lut+UnJlAzk8IPfiP07doaHXOgtM9ATpnMA+Tc420Y8h
wZ2WfWi5Z/rnt95wJHiGuAmurg9QLbN/IhMjeiIatFy1VKnUJ4qlEl6RXnDvL5ob
t2BFYLsGAGDaPLf6+V9mByqDZdEigvSDNDRzc+aGFW+yBl9W60vGycFSI6vA/3JC
ZOSO4im7vQiWhJCDrVIeGwP0ymhVyF5s3RB6Imh8wIsLA3LIqVA31y7T+fDCkGd0
jBHJD5VmEvbKKyEE/dMtN+fibyH/MHNQ6dHH2hvuOI+fR1Oad8B9lIOKmyyu4dXg
VfOTBpb1QsCwOY2qYFo6je10+9ov0u4vyEeYNsv/bkRRLtLeYG89n+p7+HQcFrI2
ti+Fvlj94o3BKpO0Ry07vcG6xpVyg5NXvL5m6gdpgav3J7SHt7u/OjyLIYTgqwus
GMiaE1b9ZzGxkqg1YE5NuKsFBQzk71jmrmyzk2C3auqbndu0SMUTl3BSp6airvHZ
Rv7okB/roGNNoxfuDavmOPwE4LJVEOEF7qA2kM/bkaPFVABqU0OhaeOeCbsgICG8
0RQijUie1m5aMbyi5K22EuoKnfS67t0O4QcMaRtRSypWQcgqhupZMP7ESOE1Ix48
zcu7jXn4mBwL6BrwBYwR4q/w4t6mpWjgCt2BWiFRIFqBCB2Hfk8QRzkrWYLsKC4+
VopVeaLowQZ/nmtDGyjckGmHasG0EjLQyKFGGRJOrW19GfsTZUTznBUSeBTrDJIm
yAvGrbPwYxNppD7xGBUiNZGT1emCXTa8SAbeXEK/VdIrqRmg/0d1tuu5Q6xpJP2C
ka5yq6J6YxZ+qsNdOlfZsqgywMrUrjUTC7zkfNsa/tt7htzbzaP5uW9SQ9ZzbkwF
h2Cj1KOMWc7PUn8ClDLu/ygFTmrRoavTAo9eeQAb9Ma6avC/vw5JYgrCSOnjeGJP
8ti2wzK2G9yR9iTTeYflItxUgIRsOnPk8PZ28r/fgw0k2KW3I2SOtnSUof5W6Ma8
M8nXeU7Sde046Fe1sm3v6NJHxPqM1JI4PPtd3DZWdYtDdglB+G4PYh8VZ8ZQhKBZ
6eDbHrSgVHy+Bg1Vc4SARwDh0yeZ2h4ZXyb2HQFQoJL2ylB1XmWyGYRvNa0s9pqC
H/8S3oFoXz/yixNZPvR1ap5zzLEHnoBZF7nWLdP/vfOjE+iKy9bb4z5GScOZ9x8+
ba6veY/AW2/j+TCSQYY4LlwteZL9XprI4Y25iUmRzY5G4n6evJgCru6ABx28E10z
+KdkH4fpPfU+rqAwWAcu29g/PIV4a3tBPgxetCzTYj0y7ZJe4T8WNjIxn48pvySv
MEl+Kk1UFtdWwjwVwklaVpx+nSr9b8PuJZXbsKBCw64kIu5CN+E7UaaW150Hfter
k7i5+MCVeIQnVIvwFhLDGBkhtg5+tShW0yZgqcD3L8thNdKuz6dGx8Sgps8Wv2mC
vjoQNE9F/B+ECMzQmgD2TD1KBltPOzNwLel2DpRVDnlZVzPHBacmOht2ochDJ24D
0tTVufaN5V+dHExXwFhHGLwxXvWt5KaXzD8oRGeqLQtFLBtYiMgpn4Rhl7N1H/QM
P059c2vG6kOpv9ydNNDziGF++cN5cR9FPdxPf4tDEUPyR1vNrjNFqxgJWWdVdo1C
Q5ZAp7fLkV4AWOSXNhRUdf2P+CHCf24mxHFPZN3jOwCqmiEygB9c9/GvpLuMJzB1
KCNyB3mufATIfKKXI55CmpBqlBwcNhhFD/zWxJdkgDPgzJLyKy+kwqo+K6uYexmX
uV7Z4ponLMPmBw47JLxt5tGB4xo++faMrytKNCbClIS18V91jaECu/O3GPYm6xpE
kQqE+X967wpjszsNZk9S8CJlfabyhzRXESI6yrIayITj2U+UJkAxBow5kgyyFOrf
bMDIapbV1DjfiTRNjkCuRzW7w6x6PfQ6z2mere1kk7r6MR36qpJmrhQ8lnOWQxOB
NoKPXWFSeAF/sUqYdCtTYG72Qf90/9OuoepqXZQWzWiZAUMlztFZ/ms2cKUq09r/
jR7Ym92dV4l5vcPJLTdibTtTtWy/9hLp5Lbqn2aN31/uZJVpzsufcd4CfqPW6ZCN
sizMwiqEbDoYCav8ps09FSQuEjh5guv8gGX646i9WvgNbkZw6aw7xg/ikGmo2D4G
H+CGUfSPxDF6u5GW3t8bXPjKKw9P2ImYlzpn+hTs6AI5SuCtdTLmHSuT2AmlUV6a
m7KbjMysAdK6pxI92i1RwOpoL1QhI8NHAsFu2W4WbRRIMGyZAualNI7SeTcxxhrk
lmHgQ6PW3pBefxVKKmTKWZCyvxDGi67+7lrqciGA7ar213LnWueokffBJelUOfv6
lf0Q30Oevo0OuZhyv+nDkUxPCXXIlPKwtVxCDyk0QkN3FfDPkQgXGZFvsMOVA/ng
oiBmHTWE7xQHUSCTvuXVSXADHBZ13vPveWTKyhenfTufgDqXliCYTsXPDCXe6ldr
Ria1/VAoJFB0HlhmpHouk7UhGoT1q+SAnQ2VlyYV1VvigFjX1DMepu8cG9ujyc7w
rUYYiHykFP+irRRZVy6qtWb55hXMa5Y3gTQ1YoTNsEdVX6anzO4iM18NvojNN+Yq
8Ro1EaTRh7PvK6K9jlnfjSi5fFmI4XPw4rsesaVKu7K6gIp9D0Oj1O7ImmOCmP2t
5sUZZuFHwLMgoaYikvQQ4XPgOI7thyEq0NDrgA5rKRGpM1I0einxkwxAGkevBkOI
1wX6SRM/qoJGVQpmyH2NdYQmFTvC4LOOlzFatmkT1jGra6Gc+TZ4tDQpilxyzzSr
VZ3ZtZsPj7CVGMh4YyrbcBV4wq6nD0RJrSUI+zZYgHSj4TN7Q//1eTVPzrVGeIdv
WNQb8FGuVT+37XEq1gGDJPCX+g4Eiy8xoQTR2k25ndD79NiCEAqlhgYXPpASoyu9
TPzheubSEPtPGM8YSAPGlZ/4AQRylhqyL/sToCYbYxVhbPFsNWIN8D8yNDtPdqXQ
o2hX+NeGShqIJS48VI9JMWBxACfwRXpoERnUGXIXHyvTWXsoO9orIDRZktfUXuXu
zHImR4C6ijV6gSThTF/JupVtk1YCe19wSGRQKfmR29nT53kXaqXYzELIMY2NDbQh
qr8Ex8zswkAFOCVyjpCwkYpT8PbEB6ZciDVYYpddrDI8xxWmhW3+Tvorz7JU/lqx
kVW8yylQQzl2q695fflpE/uwvhcv6AOfgon4VFrlF5VqK/PtZezbCkhBk5wcH8b9
wgce4U9lVkpqYdB78YNZV7HciGFlISSJ6UHTudTmKmwjpwT6K6SBUjKW4YnwGm+3
Oz6ISY5OJx+3NGADYYkfgpqouM1Bnn404Tv6M0YODyiKvQA/y193Jpvigcq/0Ye7
JE5AyVI/1XAd/LZ3jHxZquVCFYfkXg04ITL3mQxMDwnPiAgIqB6Un4hNaDasKxk4
v/++55HMMRIgA3kK2li41HKLB9OnGBMhnqitKgj/QXB1K/mcfAuq5sYGZXonv5GL
BWEi2jd+nEateHxfliWK7qvr99o87BmZwHyOrgBTuMf9pLIs4/30WWaQyLbe6MWS
LACyzt/1QvRuUOCQKAgIKgThrkJrRbnhAGHRwi6Au8cZlkqMzdWe7/1H8xbo9uY7
u6y5Z73ogDn+YpI04fbeuiQk2VcD9AXLkaM8xZHG1wsAJKCilQkG839Xiwvw2lZP
fBbuc8rVLH3sNcCyZkc8UewoT65W/mzvAcfPVhifj4FfqnbRbVJh7N+pTA4+1qTK
IJ/3ktTaMh2HlXS1M0xyC0LrRm0p5Jd/mbwuNWw1E0x5zm5zqtrZM+XZ8See5rwF
Zu0Y2yiQLqR4yEgOktCvCitTwreKtNTxghVYXIU3fG8O5NJ+vJ22/JrUtpk4kSLl
V6Vn1FR7FztAk4TxNkKdb/EY6DBCtd5j3jP8oidM/eU23HeA1hCpEkWyjNiFcvhH
E1SomwHBC1IPLi+1d8bosOJTR0LPmcCV9u+tIgqGaIqL8A2kqUSQdL9D0MW0wZSF
SImkfFK3rvUwu66Afb2oAOp2bc9pA6bp2m+EKk6M4ND4FVId9jjgj6NrVaRmZEjK
h8garQ/izRfq+e16KqWXl+5JXdUmNLfkqIP6EPJi8hZNtlF4Honumn2tjFklDJ3m
gOeYgUmm+CPM6rfEG4+3qFTpLwj+qEIYrE1EAq5Dm//b7UMPfR1jvzW/K0Tloy46
Wrq+sWNWi8rZXmkNcRnTKDeWe6QSQ5mPhrSzNSEXCTB8HVOn1u8hGS34rGWGhMTU
FDbsnQNNlS0MWM2GdIyHD1ww8v7zhT1p0LsYNNroCHPiAC72kDdxrREv0Gtu9uLK
g0ZrtfJjtWIhUVxke020Mc/t8uCUjZ12m+6/bS4cU09fZOo5Pq7LLj4n7aqueQjA
5BvkE3dIhrUcPdqs5c+DmP58Cdyz04nxyL5c96IAMztheLzvQ6C7c7ph09GEvyUp
vDNeqlwRnsTwBpr/+jbno3/6oRSTKw8Xo6BHa7oBz1Aiz6LPIpQWkv6cz3a/2pZn
VF8pXtkLGauQkO5z4IjksbKuxBfMIBaIfPIAVmc1V24Mx+BOqGnWdxeJ0fQTo/gp
7Lb6J+63Wgy6bDIz2GgvdVMcOtEfFceXUGg6gx6mr23NaZ7QzfhKR4WdS5i65ous
Ifk01J/9WwdHsZniu0+GsTX28LSAMWXyOoRL28KK+ZFJMbQFhP6Ca4NDvY/S4EDO
2ntsk5LoxAcEsgL6/wlH9iSO/n1tJXLM7KHpVtyyZkz+8I54DeDnaF/G2noUPNwk
fQA1qsmHmI8KbEegFjBSY3uJU/WpxPXvS6Sgt8xDVKJC60MSFNlTVnYaOL4uHJgW
lmX0nUMPjfbF2n3U02xCrueeMu/efxU2Vd8CcSV8ZHMPy7ppCBg/FHtwecdhZf09
2P3HYLalY7bsO9+OEoRjrLIj+xMdcIYtDmKeGyd3tJX44Tt7F6C/5d8QdeWzhQ8d
8sYCY9UxJQACn9LO7qe3HDfkUXj1hge7RyPmT2f8n+wUGSn+KJCddf+3nZcOVcLU
aCdiACRJIu9pYOhO47Bu4p8bBxMfjypyhOwYKqsvwVal2BnUf0OIAUCDfM0zrCgd
aNWNDGStMxupAxW6GiUKOpn+2eRmjUah1UymiQ3yOEw8JRCWKGEplgR4hDK5D5uj
MdBdb1cmCDgHCyGLevptvQ4AYgB2uMo3aEK+vqGrMo5OaVHaAZyVOBbQWSJe6Akh
ADPHKCiK0n808iwMSSwxzqupt6fWxSULBDTBDmGB4ybgBxXuF7zF9d5M5mUZzNTx
0F25c3iv115vyj4hCWf6LI8esBbfh5ugQU0UN8HP+cBzu9bvl8HilbcPtIbkUkP8
aNIXIlkR9o7VmwM9vdYoct55qB87dEt3aSUk5WTE9jAbLPv8ElOHhINM7sQxSYTx
JBEUyGKrTDV9lGyGS7V8yZhCTcNWe3BZA1IRFbZIapx7Lm12wXWNQ4VsIC2QRnZB
3jMrp9Gz9xPkpwPK/kkAILFn9lhEsjehIpJLVBR1YDLWqJtSKnivbtJ5dVeJBLq9
8PfxRdrJN/EMqZ6LirSbfLe1gQdmhel+u6BY8+LupKaDBxkLdTfcXt44VvEUogp8
3R9XNyFKS/OG2gOYEId7H6BkzoGnyTz0zeMQvoocw5qx7+Iq10+Z3GdY/53VcP+o
olpBb57Ox/rTC1kh7uyuzGJM9TvI7frfIO8Nwfa85DtPT1LmVj6+9B9A1M9CAIi2
j7MCjHPwI+4uTNey2KotamJQiCNX0A3mJnpKBwrXs9Om/NVBq1DX0AekY+tV8Dzu
8ccv+TWB1xLAvnIhbO9vzWD+pfnBHKKtJa+bMH+ILqN+56+g9N77ta/o/Fgw1yfm
XKzKZhTtVd81+YhtY+oo3uzL/rjsOMXk7zVhyKmbyHLiTp0/M1e71ir5kZtspJKY
sYLea2rpCcquUXoCqFxzVdUgp//nhmmSJYa1xD4pFjkbTLh51uUtVWkpRyvN+8wv
YM/aJ70IpaXX7Mj9Ll6zHHY3jru7V0huBIe4TRuy61nAwLC/Ql90tz9VTs3f6fY8
ZKaYxu4o6H30QRrJyybi+YQR1eQbvp8teI52Vz5pjFR1U9p+TKyqaxs7bI5iG2TT
IEDr8cqjlJZ79ybIdLlcBSldbplefVptCAci4xbta/WNu2VyWuyqqJOYjCfGu3BP
UPUkyeqZdSMxBAoGkwdhzr70fMmIr8s5CLOI0I0kNg+N4dJ42shKsUxxrlxqWjHi
gACtbly0FZ2Y7+aU57jMi88qNkhSxtCo+NM0La4ioVo7ZzIp7YPcXGoWNKjNiLxn
L0s9Sz8kHlHWRYFOfqzjaUzIUoJ0QSNGF53QuvAZA50Ypyr1OV26UfjCGBLW0zZa
IdgnIL5duMQJxcg60/qFbGcR98j7GebLdk9wrurORKvvqh70T8DEtuRS1pxcL+Tf
cWT7Znz0i6sg07R4lsIiS2KvgGEdptef9UZWI+77TwrINdPxBbnfq7Mu9hhrIPCW
9B3IxK4ZpF1vuozJPelErO6hjrmvSgOEZgo3TFD45pSAkyFqNSPijgpmUYfyBng6
yannmufNrwM5+q/BTLWLMP9IZS/S9GVzE1+btmM/VRYhqlnGSR19vhJpwr13zZhC
rOQwersnW5HC5VUL9HhWryW3OEuwWr4+HZOXLOerW1A8830tifRIqrTbfLYwEt3G
lUA6iYGcrxjndvgzpw1vW54QEwfuUbj+qWWsPyoQWOIhdWhLDIJV6RutpZCKM9D3
Cc1p6ljCBpO3vbYL+e6p5EDKDT+Ddk2QdhR/WLDMgpvC3qmi3DZvc/kpWpSpFkAa
6XtSXryc9ZLvuAiycNWAI3ubAItA/nyc2kokWJ1VOLbQo6RgXvMGWlrdzFomyOIo
XQKfz4GTc5MZqCUIk8vEuOlb/MZ1MtpCjC1OKx9bcsWyunV+G9s7jevjVuSVkrLk
RUpKhOu9X0UQ0eLyYxkEqvBu1JyRG/OXZ8AOMR8N4VRzgtorIvnrSCq8UntR9gTg
lRsthWXlkkVBehwAWC+wh7r55vnLes8BUSWYR3y9BbVQYHP8sj30E/Y1MIL75Wvz
K1vHxWpca04nYe4/gO4UlwcAUBbQqJwNvoRUm0Bxj8jF2xRWFxOm6TgF/uUuZFmb
0/HtlG35Gkbx/jfWxMeEIbvEXn+pQqpW1HDBHMGoWbKWYuH9MKWPAndm0fC/BT3E
q/vjEPNfo/teCnezbCMHSiCESf+kxU7QEtxHw7UpicqLIU4JbyNgl/oyEb7fasJC
UWeNm1XuNjNpRIg9iTWMO0bztnmik3djNxc9+1H5eTn6MWAFgQLeeJjjbwu8jXts
53lmxMCc2Cxde5Yl7FbIyciS3vPKTkCA+S+Ox03K1VEfWRx8vK1Z//GUdsut6c+7
aKfsURKcNDNNTaelOElHrHmCCTI76OMo8halIny4bNglrru/kIsi0MPrRQrS0nuv
ebikFPeATn8tfMgazFEgNUv0g3+AwU7l66+SfJj0WuRSisJ1uVLF8RRSpl0cYVh8
AArmCcjpqRISv+hSQwKQdZpZlc7aaMZjDdjnNG/BehDgjhTlu9Mjx4W01VEhLbse
hlBsyILgTCq+YtBITQQhnYWKpC9AmumXclInc1hMvUKYsfNPZhjRpkH5jT1RZ0cG
Ep4Xi9p5EvZip7HK/2U5NB/oyEyaz9cUd5w0YpykP2wy8woSUQPvUgC94VKGN6Wt
szRrJjxD+1gVp5GJVpUkuJhZHbA3lukBPygvVAtS/xU6mbem8so7bR2LY4eWawpH
uJCNdWkDHnl5V/3yxkdZeg/aBgKXGhNEzpeVaZZ0vwR6Atpu3kcufC4rBpm3G5Ki
LhSpxkuEcf+fek4TKzKM/12wyuZZeqybLkag5MVfu2Z/4ZCS75FDuGYzGyAiU2lR
2v0RbYJcX0ncacMUBYahTtE5LAj0yIMQITrZiWERcz0mtWOx10YDRmVBLanQc4vo
C8vO/B+FAj3xVABeTVqG/ph6fs0TI5RbkGZBFRNDKoD/6wEz1NAg3UCPapAn0hSv
cqjFZqa6Cqcl5WsGc0qXhoy8gXMvlKMBHj/7KyOUbnrt65aQHKqlFvYBuoesYU6t
XOYyRf9fvGuABKDN3/NTM69Yn0+//B45C/wLGbsgdnuIdTO+T1Xzo6NrGIGB6cPz
WoOxMDqUTs4rjWUh2SJ3AL0c7q4MWnAjg4xeMI6s9VZaGxgfSqXUYQOKOQ84ZIPc
6qwlZha7MmNKntVPATVUa7ZFl5JGVvzghVTMm+Y1FvkfpDb/CISBK4tjntuoCsoU
71NW39Ex9ceISBPDPdD7g+6wUCN02nIsvDtHq4rklJ3EdFGX1jY0t04zK4+htVk4
HQoHwv7giPykKcj4DsY6Gi3wT19UOElWXeO0EfIxthJQAu4i10H3SHU9kGvSt/TL
SpLZE4Dkn+Qa3guu14oYuJjA+cGSwTMP2RyhS3PC+8u140f2P2nnK9NNjB5n4rHE
OHteIpDDsT+sdlHHZrrCT8F1N/pt+0h7sBt+D84sVFwwRaSnQrJjo4eo9oah/IZY
XMt3Mgkjwz6bHKwUXOJ51FKd7F5vw91vLCGoYZwtK8LiNuCS+Fwxr6UMoOLrLiLf
gcX81gb888WpgfNEetlK2UhrfDsTzNWN6NynFtB4nxD6skCL/mZDw9DyJ4v5oBSw
Eb06do1gWuaxaInkpGPWZT9wwA9xoUq/TsvI9USath6HdTlwWVw8PVNPt1PJl0uM
9byIfy3lO968vPBAJZpDR9cDB9fEirCnKU9LpowyXwLQHEgFEbghKVm9jBEyg4bL
D0nqM537cLZCSwOBm2umSAl+x6ULtvutzeZEGGxs6pJ+cUQNEjjZ3A/7xmdAwWut
vxGyXahtx4iqYJBej4ezttqzDUHs7jwdgRVG8o0wU2rNAVjplkHvSf1Za4NfymCb
7lNgf22EM1ylfR9o033bks23EiYLpx74xv9sS83f2YVlXg5oPfD2XwpLzAt/Gpqg
Lk0snvsz9p+029dIavif2Krc5IDuX5qnY/MRhZykW6LRKRKV1KQRxwpnyqc/xr2g
r/sIPVsyq8EPIHuddDZb4lRglby98xZ9Bwiybd1wSw3HJeed+QNwrNz+Ga5vne09
YWNBo9VaLIKxFCTTR11R/Q6pLj8CsneI/LVj2duvDTOL0t43T8SUlurpJQCQUDBL
KPlbQDWXeSbB34gcIBW0qp1fSdkQ7DB1e10/KK+VXY59MPtaHBJM9NK9AdT7EwdG
TwAdfhdxNxZdX0dz6M4t8zYsngtliClp26R2WTTlnU0VZzpPILjI39rXqgXTsx8P
JpH+qb9fo+8gXhH9epSxPBGzcXtlXnd7we7pNkEZhEN4T0hJUjYbll//7uiQQEnA
TjVteYj4oHSphYAzyhJRFRtOz7GSJMSGWmdU+UAKoY3U7+/y5mqbg7XeKYYk+lJl
SZ1hLimyaygWTcrF/nHovYKCm2gsiki8zgoPZku6TqEzoXzhEArvKlBd1Xv02ygT
eIWoryh/qfHORmwyEARGaRl9DhCyNJ9gaIZ+cqpMiP96LLy2Ev9++4Q3hELq8Df0
wcZ+NqZaB0GyhME41uw2PYnj/GAR1NtTTUwYXx0YBA0Cn7H5+9zVgOwnklaA9AB5
8h15ouYxwoH6ntm06igJTu2AR4pu+d6ByyY4sFfMWq5LOquSWXd46yMTEJaP8LGt
TBUWkDGd9bX3mBHhSjjvGB0e59tJfQ2tGK36bggTmFbyy1L/3RqLPhOcxfUao0am
ymXtHdQsBioytOOzwp6vee+uPfj7a9oAyaLxqJgpyOg1nB5xELC/MwJXLnhTI7vL
HYaw8Ts7Zaime1xEhx2urofz/4MkwryOQFGPhw1gPVgXelF0F3WIStocH+5PhRuE
75CVv8LDg62LzFtDMorif7ceSlVRcNHPdALg1myPKx4pSGMZAyRjFLHSblE+aoxK
XqsUvMMmV/eFvUzMcxmYfMpyQy0GjDVqdBpSRpj2yb9rPIazcVce4JK7bdW43yg3
qf6bHBKn2zRtn2fTKyiaiP7gJ+mh9pkGFCYce0yAfjbNwv7ydxMFbtMOkFTc5r1/
eYg1LT1TZjAUtdPjlD/5R9ilCMjRMt0XzIUGmCUermPYAMESiDfeSa4POq1pA7SM
CdHLw8zbPTaU9odcFZFfhBKlmqaRKN6xnAm7iwiTNf/qDAaaf4dFdBUv1RI1ZWeT
stmTJvQA4Hc82S5N8mI/LC1/EsYvlEfyxzPd/Wx3SRW6Mh61Iq5mclmTKQg4wE4K
8GPNaqmagPsJnJ9LLen/knviMlrG3zk5L0XWGr5ktJ1q7atukt4m+EuOmNNxBv3S
C0sQ5dPU6Q4xZ4Eoeu8BWbMJMH6kXGrlxCBxNBTz3VyHIy5OFQ01eNM56y6RfxCE
WJom3k7V78La5Z27P8FPEBA2LYyh8MfeQGp81OjocAc7R2DdgQDJe3g+kDNgEcSj
AkwiqK30qX076ksV4HNU1qMGgjZ45djNDkeW0h4fe2tdc1CfHgwBQUEA1SCYcqwL
G7sOw8e72PZPX9upJ9g04P7sE5q+soB50d5dqqGURbSFaR5albwkB6kRA9/8Usu3
RgwSxdoOK+LPyLfTCihz+OOoanhYwD7EqB95gZyBGCh/j5WHFiT9HlO1rIJgysU5
8VfXEaODHGeT+LrHmElA8ffDZJ+aUzn/LV74DEKy65cM69mkelPKR5NdbYZyhoTf
lF+sB57pa9Db80waURaNm1L8NgGzh243BEgk2TIomf0N/eKB2NzBTbHrPaIL5ASj
O9gELCKjQYqFVlfn4r4BisZx5I7CVGsexrbhX5AAb9KCo0Po068qTYcG9KNd/bkd
MqHjbDPtzqwRowTgdyK9hKvF6KfZuckCirSl1bYloAjeJ+4x/rHIwmog87NGjAHb
DLhzFoB/RS05pvfbIRhCNQzhy+edfyo9fSup3dTD2cTyirtXWK6X2LfCCSRHzxrC
8qvtApSGKwFSIbN8gvvpmpsI3YHeJzr+N1l50xzOws1hkWikLlkNtTzvfxHQDI5o
GYVx188Sa0QZW68k0/j+eeFkz8xjykeKb9/8sEr4K9sMcHoebED9VNcmGmsqY1p+
F7q2n/O14yOJkX5MmEvtGrsgWvO0uWUX+QjyTX7Dj3k80rwtNuPZlmi2icClSe5W
GSGpbJr8AfbtIaiSuam3lZ1DsZ1qhpSfUjWSVt71GYpU0WBWwDl3yDLB54uLsTYf
4k9nRPgVJNkvFsBet8rZD+rHHyoOyjMzkwESVlv4p27RlTdE4rqMh61GVFDB83Er
+catWVQYpinUqZVavGUd5HuoMZ2qmeOUBWJ3GXREJ2w+bEofmXjHQ9DPhceWkif+
PNv0a9nom7WtbBTErbQUOhT1J/QK8bLJYaFhBdBj8EOMSvJjW2vq9+o4AepCqx43
XZ7saN4sM87m9aJ19fzih3CSS2BFMPej8MdG/vixNIF5m6lS9Gpuw0f6MRBilnQy
xQ/cThI/RefvDzofN9dBu62tqI+oU5owmhumRF65cEAeAwgo+UFVVaK9+kMFPG4S
k1skbGRewQajdy16Thm4lBYM1qhBNrQ/BgtHpuURXcE5ZEADSa32PoES4Fo/+HeH
ZmhTfVdx6NNClUT7DWVR5yN3rLhCKBmbXvWfOrcrVha9hThxGB7CbUpKDnBO0ndA
wH0Z9E6KTuJ5Zi+04gzwiqwUol07PW6fptY6Jm21Iie6f2ce7U1uwKUTnBeeBeF3
+TOAvCCowwi08SBOPzxlQP6YvG7NN4c0h5KXS7aEzN6Fk30TqRE2SCIsA+Gqs4qJ
iaaC8ucRt+p7+yP4+2nLrcbQGNGhFi06O2yKEVMRA/A1BfavwrF8WzP5aEULhrhp
lJuV6BTDUR+EMqeVq1DTFNtgk5Xbzz8BtSOw14AeM5uCjh+KIrXsw02lp0XA/8CV
N2uYEfoXfj9R8mc82m+tLkCD7ZOXSPAp2ZN+D+Sm6YWVsXVaLeGpnr8ppn4fTY09
g/On30W+6MrwWz7BbCsxq/MJRzcI5eWgqHFBajHSPvnFJd+9UpFPNblxlsEwRVGm
EY9oMs03nNnq1dBp8+YzPeul6koLPmOHeM596eO1DB2ggijt6z1DgzrNYC+aPIbN
rSdiG3FJ/ZFrD4khKh8vxhjRg1TlXmgIy0hOTKXEgEwTc9cfhN4z43RLmC3kwBt4
qPBBfi5OrbFeJfboN1HbiU0YHkpp8HEb/YbSHh2sri9/DvNOckjZ6nbR8AKoLsBg
ni4nsWVxo5XFhKQbW79FYHziEJD1WTkvzpDWE67qkkqIch4m/NQL4DRcFa7gBfJ5
arqg8Rtw3rwfMg/A8Uk6VKyRheZOEfKJU71q/6UPjhHaq7pOC8p6Y8gwjYO/5NO2
wIzfn/9JlBMVUMBo2BwTr7Fs7yS+ZhtL6+QIo+U0fDzow7wp9YJXoPvQr44bixGH
4718g7KzaW8DaHK4NZe++rbrjFAu/39ABlsjbqAnxgN2zH5XiuYJBEMqpcPgkWq2
ZJGovBlz85oIadktzDzrU5r5UX+XsuH9heTyd3As1ddhfyG/JaLJc6/yTyJsoNJd
e6w9/bYxaF/1cXTtplJPAMeZMY7UhC7ybiISOKLnI9wg8CSajydCjqelRWO63vx+
sJUx64fQQUsW6pXLTacV2qeF0xbAsS8JoOubs9FPo4OLwuft7yCm4JnAYhKdteG/
E7gc3oc26P3ifp8b/RkTFqN0DKA94Qs6C/13jMfG3QXMAQaqr+EjWMfq8XWSNsuj
/YhHdbGCK4e4Ynd9DJ7lVw7m+liTblyLQ0Ip1/fVRZfj+mFQFliQ/UpUj40dvn5t
TMPEM8YXGGwf6QobVWqYHzqzbx3ea54p0Tw5OWPwPlyXlD7LeR1xPlHNdYAQnh3S
C5C52eqzKSO9+9R/XdFfNbiw7VRkMUjrWSmNgmWHXZCdty6unwhxN6wu8alezfGW
6haS8k8yc2z8O1UfxJpxkEQCVMRZU3XVfcsMjcGXFcj2xYjcZ2kz3Yx2e6yKLG3j
eBRSwX10isiYKG2hyn6urtigFFBgnV1DgTnNOXSBafu1CU6JS14U8Em7WUKzIb5B
QepMA8zOyNMCJjPQnknMls/WZGpB/NFTPvhBzZTwsvqBeeFr0b66jJ2bpOX4gC1y
68gF0Ue/stdNXgtRTVzDbSywbJAdUYc5v7za59jgEXPbb72eVsHTJqr59jSZihp/
WpeQIp+MTyMJIF8NO7p0mCf1S3Fy4HfqMNCBiBP1M/Pm6Ei5ntJZjroGEvHeveMk
4llITCJLHtulz8sy+hOOc1wIOimLZ7NopV/AFsZeO+az+5ri6RP1Ue1ka19044uj
iM7vUBkYcOKhDxsdkZj3dL9UftiDXXOqPzdME88zOoVf9s6HhzjnLLzib32wC9D4
wYs33RLq0UJ2zc/kl/5qluIKoHLloYLQYnhKQA5efsfj8Iv+UvMyygxrOtEppCEa
tcOhSj8CGWFP90pHM7qZnAk3xAvsLktcWw6k49CDc7XaGnrKyUcRDNmq5djsGx9x
XcZuUgY5t044rHhWZSWBo05634xRBenTWN4D4V12nK5BvCArEHzQh/mg5Jm+pC5I
4r/Ble9rukLmPmCuWD7+8Hyz0j3JaY/qbgWu46l8xxQDJFWXoSmTSUCirr2WDOXa
KzK/5M/V5fpQCygSMW5/IPpoqin1hCB8Tbl8KrlzkhD8ZdJtOGuUfreo9UQ12HKh
FWr3o2W/IZuNh43kfa88AEBmYFP/En+vYsqrUyvrCJrkRxS5NE/8XitNQdGgjR30
oW0s4hd9+6WnGLdMTsIS3HU4Cx7hKPBX4qnidgt6+RPh8sKaLhVzs7emI291F36l
541QiIDQ9MmAtcMd+Q34ZJUNIuVEFkVKPlno4Y00FVBKLfkICRHTo7IMGP0zohpN
nMwmMff+3mevYXhoqBZho7T2hWkZeqjr1kuhFHl4slqhPCthLb24DYqolMltTQpG
v/D1n0JpDakvHIJVxAluB6R44H4cqBPn6I81c8EYCdIdkNjcwcfRzVeG0ZRV0r3k
Hv2tFxbASeqT3NrhoJtey5wzag21AUdL5YfdIgJChysOxCP96sHKCWlhLtwFpnjf
TUzeevtbvWZ1Z5pnngY/uWqWDM77O3/BfwBn57Qdc96ON2uHtoCH0Gbh/L7BWPwp
+zRZ8/Cn9n8EzRzLJK7uZThY6njZ/NKKouQlf8B4+7qyxr4pkdKpvybtS29TTHoD
amYyIMAySb32bssECf0YJOpeWFVoqK09BFbP3tkagJzt7AKbycYRVDtKYS4JSGma
7I5kuiVy1PU53H4IDoDkGp7gc7Y3bzMg+Kxhw0U+o7wDQ9CrIQSacXphGAG2vg4j
R1mOCSmh2tZTzP90d4PQHMRYeVAX/Iri8O8a8Y6iW4mFZSmEITpLV4OCj4mobeCw
0RIwFB/GrzREZuvjQGoAhJ73Pdj/bsi0+Egi5flcWBpPpeFo9Zt9wDzOuX3+aArO
04OFJEAINQoRyClPbcICS3FHmYFc0IOQHWk1ieliHO7QyknEsmkUEcpkI5djRd1n
2RZPXQjlyiIfKFyaQA6PFXr9tkQX/Y+t2wMIPbDqhXyOKrz8CDoLeCtx+BTKXXaY
75SVIK9WB0l2qV1eidjE+eZunbDvA7JsowIcqMpgHV1IgzOmAuB9xPhw0Ru4vF1R
AhbVKltBfmVPppB2XwQF2uf3WegQtpbJCRCLLjmMHJEqQ2bWkwbt2waso3h8tk+K
uFauWRK84iOjhFkN8YzoarmeYzn922fw/Nj/l8p243REyvgh+gQDIkUcJFPb+Luq
LbSN5TLSKe61EfHWwQn04NnLy47fnFcmMqd3tsYI6QZQO8o+oozsATSvLPbqR16b
L3Nmyi/cYcaDFPO26jLdv0PQOF21aExRgEjdg1igz3t2rEUESOnjFrM4Vze35lhF
UeIWAtpkAiEvpEMiOOb4zH1CYHA6rpv1XxVpS7vuYiBJfODDpLhpfkcR+sZc8b+v
x58KMe+GZ4kcRpGaIfHvaDPipePfa7bxmyNk1yFrw3DP2+Za9onkrd00kAMlFYya
fZCjBlat0MAKZb6m+jR8pLBdrHspMDocWhUxM6j66Sau1Pv+2AZmJqHWc/tZeVlV
lxXkYUpnRjC3S4H0B4mMWM90DJ8a0W3it8sMHCHLgp1X4FrK3rBCD1g1nOZmlqK1
bMI+Ctji7Tnc6umAyvZOndzyBf7LcdT3uKyAtlbfHhEA/CHG4EnG1xLhmgsJ9UOT
eVQEOVybhR2bUMtJqpjwra2lz9SlBP0s+X7zMgh3WfvXy0Glc9WEpvaZeldlbpoz
lk6YnqrV3xr/CzcgkbX/yVNBqWiVn6B7AEc1PBalbDDcMSPbBFjVkwQanC2W1F0z
MARcRLmgULDh1doBy0BtEM7KOwHNLrcoP7Z9j6wZnui97EgdV14VpJpEBbGpx3c6
ZPLUHg0uvub6429p3F+cJJf8ze1fVZrDRqfIw8Al7Y+sDP8QKKHoA4vh+Na0IHr7
UDrx6kfIAhHs3AoYMihJs2uQWcEf9a4C4prXyQS7TDX8vU7Ig+gQZWKFG72sjRRv
AicHmcaC/zpvdDueykYY0i84VoTYEHv2BQT2p+cgks1NjhkZP2vYpAvkS7LlrTdn
PyDdEYDi8xSn8S388Hxd5TanZEPZ2WEdNoQzEOv3d1MjbLH2VtbDhhihSBux+o8B
nWkHCsS89aVDhC/7eOy+ch88LbIOAfmasaduKOukFltYrQCeovJogo7bo9Bl7uuT
N43vrN61Bm43W3o175EOdsmQuTUn8V+VFaJk8ZO2Dg3OdbeRb2w0gARrOTbCaOmF
PF2bN6mAnyb5eHWQIB+N0D/G+bmCd+ksFwF32BhyKuyxkwVW2eybAldjYoOP1pFB
6OZydu3cKVAF3nJqdvKXONgZLT5OeHvixjqrzMEy6T1bRwGU3EdzFeXbNhk9qcZY
N1wmfASxk7aeKj4fepLbg6SFyvjvsNl1dVL0MdeDY1jTnmB/wgWD/kFpUUjFkmfm
9eh/Rzt/lJOuxIYBjSU74UvKrqhJM72gMSlsHlBYNoN1yheJcp1Kksgq4rUlnRG5
VpJNB5t+XgZzy5VmS9E+8akb9N1L+Z+nBp3XmisEK/RNu45egDMi/EXX56JVZ3/S
LlvrSaYxIiwDelXDYWLcteUp6UH/yDL9L6tR4jCRyQ8631tb9w0+yALWB1zgUl5a
DQRF4ZP3l7T/U3g0R1gVPK86U+yiUsQdy7eG68JsTt8aLUZZp+iCPv8F8wV5TR6C
RCiRF8v09+SSpfoFqo83t4kh4dFt1QVt/XQG9KlqbwcVJbtIjmclAJJV1wpChElT
/s+PoETzxhBLj1PH0uv768gMDLuPO1C6gMJ5UiUZJmJrMtIuIVQfUddIrlRoVyax
+fMESoOA0NiIFoG7AWNlba5oU51pJKwJhqZimPYImOMxqRCIbtdbDVOLm5Sdj44d
WWv4risoEgb5Kysel2zDCcXAk0bJYXUD6ig8EFzBVW8nSg28RQk34Gj4VqMD2afG
nxk4gs9tDWwyXDTz5rEv3cm6n0J6kSXs+OhKCXh3J+4qEEQrURzXCP0JlnBZhjnF
ZyYr3FmbtXFJkB2HX01B7UxYoJrEGOmY5L7Xy8JvzisaY5G3BTLx4NibYHP7zE6i
geRKfeKSCa74IpZZAYW17SjA9NYrqHgP9E1DKgO2pdZu/9JJxO5WJJfJh2BrqGdy
OsHnGPPeoYHOldlSBwyII3rttJOAZ/RnkNSHQjaoVCP7TaOhXY8wzDokCs90/1c1
XIXlaEg2C1L58jHOSgrp52uexU0vAt9KZuDuq3drplgHUGX5FKl16yiHOS6hij53
gf6b3rf5/rAq6TEZjNudnAOp79/dYX1Ay+L13lFDk3Ww9lCAajn91FYuqmYS8NxF
3Q9qC+6FHIepI/KvSJfY7YtH/4HTmByzg9Bc+oDbTx2IDFboxN4SxbK3H62GI5jb
gfJ03v/RMiwG0DnrZe2SWri6e2K8bV4S3wW3WF2MBuyEhGWnpDnDfdW+jtKp3B5G
ATF2DCItswwOg/wkr2ERrAIadQkXgIDGlQEGfbj7zZfWudQVMFm5p6QVwy357gXj
EBpBfQGSsDj227lPF6wFNzs99S1QKokzAxwK6S0qBvkaGB1EZdYVCPG7hOpprP1O
sx7ghq+uZUclPt8d0lAgmSGb0H5sBxpzuF1S4Jva3uFtmyzdyACebFu9VSfRemhk
9ZK7q+AqQySwCHvB/JkVE2N2OkhyorjAEV07PWg7Xb4rdMF/619M4E/1YsbRemSx
kR7SAkP5WJd6VcNenn7BuDk5PVbi2bdTGwyQzUXIHPy4KDDifi5HlVw9xIsenHm0
qDhVf+0Gp3Fg2q8ls4C36C1kOajAZQg+/AScchDNOHipSzldEwv43NV6szjHKKbN
+TIanUNwk5A/pGVepEYUR2oTiF7zBhHPnu+H8mCp/8t6dCUOp0lXFTHI9n4QBL6v
p0vkdXUVXD6L91NHRbD5tCiu1Xmm7aCQwWOmK06hxd8nyb88OGMAGUf3FiSv+HZI
7oQHdnSNCZYIk9kdcXfykQYRIxzo/foaHDhDQwyp5X3Mtyve1O74S9RQh17YOvfi
8McBlBDozsO3OsMTwBBekZqOShb9jShLZeoizHaa6jG1EYmM6ML8zED20qbm0Xy+
YQT6gTA7mdRn81zhLJeyKCcZsu1gOzOlUysNnNNVoV4aM+84+RH3BBgiqLmLGGZx
MFF7zhUZSNX7jSZWRhVcfuEo+wb15Zqw2TAohbEYr/aTzmD+pmvpqip3OuQY50Ac
L8tdKnfRgNltVjXEcd7aVj2pdnHqsCgbb0CAVibp31wOeBecxdZChWWq1XIcCo32
bB8H22yd4k2jso/UAgX8lFr9iMTLi7BR93OI+DQPI8X5AfH6w4Sjkl/tqW7HgD3y
RKk2a1qBY6W9LsmHZM+oTUJRIVxQ0Z9iZ9Bj9eCyV/soe7Id7K2oNS+Vd8DVIuXU
lCcOFctFovxBjbR8DPPc4pC6WalUrJD2WphCiwnmSCWIrfGjJXCncYbbizDzV3Cd
ht+xmP/bmSS0GTZFG389XBipi6LWzN9/xYgsByHjPtp4QkfIBgVRhadWHM5qq8IC
9aGpGP7tvrIBpvQlTpBX7tX1r4QXCXnvvs9yJ2wm3mJRopT2HzDJsM+G4SGZnpmT
4RibcRu0xpPwIJ9vRYwrNzsK7gUgZkWuXyCbonNTs6F4GGaGS4O9ssZtsu/z0RIP
jBupw7pQvO49DMzFzqApXya6wnr0hnekYyAMTtzcmjKjrzNW6k+t1UpLlQKlxlrf
sVW5W8ltGcgf/kREWC4DvlC/YgBYwAk8M9hPPZUtzmZyiM487nwn3O/Zyu4KJtK7
a2t1PGpXtrUSh8DFO3FtleSB1kHCxp3//hJvLab6G4eokLxUeU8c3F+3XlnxO8ux
rdLbU/8Sv9DxOKU6P8DdsPNtqtgxDi+kVzn9rEaEZX38Tcw0cw85SB5NnPaXIkt/
HC6q5UC8xKc5rknfEKtGnbnaLeVtvhlgatUvhrglFSjkuiFGxFNmvPmCGKeJLTNg
62tlISOaLOyTJYdQ+dtj2UBNlObZk27wBRg7xWehLEjXBc58TogDR6pszsR3YoDg
dBJPcaR2bLTPoQc3ciCVVtQT9jkHLsEQfT26cHM7VvGR6wgh6cr8b6W1VlpBS8GV
LkBCCUyloWFxzbQSLzyYuF4nrgJzjCnUbk7q1Gr4OFCbJvbHYKNVrkNHdIkKhfBH
e3W1H+k7fxRtJAU5El3Vy91cNJZ1r6uuzjTYIInHo59DPfbUdt6wkl1PIxMTw3Gj
trVJH591LHpg6Soef+bmTUnymW2ipQRsSauophG3orKndOT0AC9eiAAWt25dtoYA
Cy21Dt9VMV0KKSZNPcEaayRJxikTeg6dnRq5SwgK38v97L7raL6D+ywyPkbRlrq4
6jPC2UginWk5zGdCOYS32HhZTkhGRqWNvpGnSGJKf1FxJdnFUCJEwA//ek3SQhIl
H7kWUtgLly5maoYypl9JdGMRX6k1LIuuR5rRlDFC8bSn/LFtXYFpQ90eMGPxcUiM
Z+gxVgTXJkc8r4BBzaV7TZLo4GWPysSr4Pw72RXMg1TiS+H6SXsitkn8rMkVzDr1
/loT9vDcLzyPeody56+mCkg7XSIIzApj9NXPVlXyfrVIaPVuP6496a3U76omTs9P
0a7Psphu+wHdipUO/mbflrl5CdTG5VUtAdoPm55rllrzk4KbhYOe4TCF51BZ76gP
0u7VQxOb0Vy4XuIfiF1rBRuDIUyFTB89jUzGxFmSQclXB1NuCG3pZPfynV32XtAD
wZuP+EoibogYzqHVPEXXRMXx/iDHPAhKquFQo6XF2tbTTJkGprUzX2jfei79fxV1
8OVwexC/xEyEwZb+RIqTMQ2P9mv3u2fk8Zcy8pS+ebZhHDwK3YJ7ZBQdqbvolT47
XbNqnS0PWUFNopN1t6Y+YJhqfFIlQae6G76klKlrGvRSxWepilT96SyoyswnPugi
NsWd84wGt+PspJYMY8lJCXYJHuzZzLm6WlezIoq1gLGwnWE835ZxE1s1Ha/aAPQQ
MIpeimSWiWG3oOqb2wueUbnKZBN9D6Uq5CSX5s6xv7ymKGuzAHFSL+c0M+bvqjQv
k4RREQu+6tNRl43lUt01ZKf+B6JTl6rKEiYmYA51GnCz5IodWnaRBysLJNYbcRza
jpNkpAXCVQCiOaXDOCsgoCRs9S1cOeiqXCxOvJzsQ3MVWx2rp8uAsWhUvPBJLWCN
xAOD3DxP4a39j5VxCf9/0/U5Iqb7s+MYIyqhTXX64fSmfuZZl3OhyEnlJbmbx9yN
Fb7X4dX6z0ZT0P/l/+1VlRs8/vshU+blOaHeXpAAPfVRo3WuWfxr0ZtDGA+7ozv0
wfvnQtFvVfMDAnFNIQ11QbhI8s+FQE/T2L1zSs2RlPe0vg6Q68bjQd4PFZgxUzNd
IfM5c5ke0tAD82V2vo4eRfN1sPPMmr1/rTYxfKos65eiU24W91XJzmBTptnaXLQI
yKZfvwaQ/fx13mVzM/18d6TfprukV4S6EKgmnCQv6Lxy4cdteVaE0n9oMECqOIiV
VNFwCKPVXWOLMPDlT2bsSufMN2XBnjQ4HLNDFxZ+1A+wgqJpBzSQ6SOyZ1K6j8Ma
pX5QcUxbwJoHD+F5DgkQil44OnubmGYXe7OYaYtaFf3tR1BF0hAs44z041JVYToh
bo5ckAsiEs9lPRTnx/smeUQZdmDJwHAImCSAUUygGy0ho5FSEzr+k63UlQwDITQr
/RUsLEKmQx6XN0TlHLfl8sAbNRLyTYx+A8oYuyWjAegndr2wjI86rnhkZt7sGRmt
js2UoAE0EhiqX4su7h440ePU8pubR0RHqYtqXYRLpbQiRAeb6BmvzxcFpvfVRl/x
5cr+3qCuifDY+9SjSUE79qPM9xXxVAHfZ9X7Qbeua+R57Phqkt3JMXP5Q3aiSuC6
qfO1ec4TR+i90TECaRK3L9XUF5R2S93gVjsX1Y4wXfVPBpd+qp+7NyCii8uEx6IS
Ce3JHGTJfPcz9f1b9PMpgE8LJhR6A3j2qzF0ri8pdacN/NqYerUOhVcCLVCixQhZ
/bzN59PGUMeV/DtGjW1CMN77WbLf13FNGJdz8XREJ2B7k+2pzooL9aMw55koQKgh
JZ9ZwxJD51jNzqBqscMS+vV/wK9FTKxGgGdnICZuP4+VSu53GMxggrjyZg87ACj5
VcH6Doaz6ncC5OwWu/qNh7HZ7vBrYJ8m823eAM84z1WoeYNhtPnVX5KSpHNznnD9
dUHyylnmUINLdKYGpvAcIsKaOl8qRxnOR74M9PhMUqR7fOcZLiupUNt0ISR+aToh
syxwN9GjCpPHvBh1eTovlurnnzL0PO2Uuonp1OkHrAC7KXETPw/l0G4xJTakzB1o
jXQUOBkOxdW5adhE9fl8JYa8pNd753msByPxWY/UACB7TAEd6VZUgEp0D8Ibianh
/qeBSLmkt6NT3wxT9HYvjwWQ4zXnuta7cdC4F7ePcU5nmYOqB+St16PVC+KLICGy
4ClPhKjsfvciLxsJl1UTpDbe/ZbVQp6W/10+Tzu6A/AiF+bz/FxbXCCg9RxTjo5m
UHqe45wmD7QEhim7Lz5dQ9h5dMtO08bQQQd7Hqghci4FkOi+eIyLm19Tj3lLrALl
5M1NfUaE4/nzB2osXwy9P/kUwPecIiPa1/aB+pC+QFI6zj8n4UllldhnK1TQpItW
qCiAujkXxd5hfhdM2gjzQ7Neicpu14qtuTZ4hBLx9/po2YKZHnAXpBUv6n5QbFB/
ZPw44vQhvgtYmKz6CIwbHn1qNqbHLH3sQIWjmGmgflDIimmg0GJlYdr9Cj6EHi+6
TPtR4JMtQ2qt+FI17T5DncFvVfktFKDSo3Tc7Wh+raDHH+dvwrX7PL1QT72axwf5
uWy4xO5HyRc/QzkGcE+Sd6Bb4rgK+HdVQSXyHCxKSEH1Fmcc0erb8mnxHViQfSpW
r3MLsSGSmh5wTSEtdEeBWPvpW6sviLLVZkHl2WRMSl6I/RUPLAY1B7qbjV2v4cyD
9hrM8aJAMG6cghle0hN9ZWKue23Dzot4k0+Q4wVOhJrkeTwpd8QgT/EicQFzeccC
aPGgB5HxzRyelW9hZHDmBSWNdaP1/LWnG5LLh4K+RXcuzil8CmpdSe/L3Z/iwJtG
D6WoiP318HsCdkBxdza3XvkuzbJwXsl+K4EcEaAduxIfQK/GXpcagt435B32lwsQ
p/gT3xjslu0Wl5jb4PzOKEY9LBhWeE74iypPBlQq6S+zkJvfpASFlOCR0GZzf52g
NKKhxPDQglf2mZY+AByVf4p9mZeokD8SGrxtDL/IsLc7jstRgMQHEMG5wNsGVOyL
6JYhtrZrgALVirnDHnZx40xXWMn7295LpuBPSgvMlUCzMAG74zBbCrcqYbns2tbM
EqQcZNxAIvQIv5T1BKM7nXj7YjCIMFwmZ0n1tUtq/vFebhg6l25OgbpiTklyhC8Q
DUKpOKKYojlOcoIqIbgcJrI/XE90CFdwwACHBw3FtKktLCefyh9Xe3rKonWOcNrK
hLxd1LTF6m2hSyhudObZHyxASYXu8owOKb/Y5DhIFbQuo9U4eb96Y74dCtSKrU+G
7/fvAr/xD6/PyPKptDmdpKSPBlqrJOxQJJpxiyqbR+La9l3m2t76SMWsbHTeb3kK
tZ06WPuLTUmoZ7p9KWTzYzUXZ50ppA5SilXnk4L+B0buXFPH/uEmkxlYCtR9wV0e
p2jXZg67ETEB5Yc86aDcDRVBHniCAr2R8q6sL2Y2KWCKtDzXj5LyiTc5zFB7A44L
gyDtFT3c+gKbxIq1+4AwqHMvQ5mEwI57up8HYZJ7NDawMS4RAGrZLcXi/SImoHFF
3yTLm/034+sx9amABepbnw79XolzaeLnSo+eLEpxiwGtIb+GmqVq2HFjfw+Bh+1t
S2tqrsEKXw9EbLS4Ao/QiRqgiEj4RsrCUBvSBoG/KBliiAAKPArbPLsz2OKzfYqa
C5Ou8u53nXbZoNU6xmyYnfwneFyXRBTddxqExyEbOQv4Vkd7AwkJwJHdHcG31oGp
cO6xUbXgAZwUA6yI4pDSkXAw7MoCUaLmuPHoB7s2kfQz+CES1DfOgjYanq+h1z3V
2q5SjFLXU1uAUA2UNcMzQk13e3cef+F98Nak5+ACZ6KmugvL4HTO0UpRQGbYFZTV
11UitC9Pxf840S5w7WzonAxloWBcPTwWPooVXo+WsTNohlvf5dyp3mJgyB5KUg8g
srgRH8RsmwRS52S/6pR7z3wRL8dPrpDFIqpsS5iJxMiv4pz0fisCXh+Qvk7w+At7
fyb23YztZw45AynlFQHQHv9v4PpHmDuhTBHy+HXjF2Lzjjt+Oft8MqBmhNHbphcn
2XuU9iKYMM+3A3apDA/eytwdDUM26yVysmtP6mVrO8Kkicq1Tc4mz0xc4Dvzfn0o
Joljmq99Wv8Lang3asgAdiptpwLykHjf1Z3/2AfuctgbW/I6Z6nPXSfSBccDL/RW
Lq9YWCjcoKkTTInq0DXQia6riKwW1CEYo8jUjKtkaCFsBObpnhZQ8gStYtGED1aV
pZ6t5QmOACyWDw2G/+aXbhfd07uAHSpYeUtIBkvgBoXkx4ldM3nRymbUGp3+0an5
MFn1+oayKDUMgRXhk9MESTh/uS/p2RzQnaIMO3AGWMyDtKYrq1zEDBj506hfUgoB
kMRzRIyle/xjsphsmZUTLYgA1FTXhTu19vV+pRD0SMTrlzERJ76n8869dULdNpqG
G+WlgG1q3hlJvSI/caBayz2tzkEx0evrNENDetRxT4vOk5C6aC/jqyHZymBCSZJv
ZGK53zbNioLz+3zkLPWraYhtoJx1knrx917KedHSneISgsL5WhDqQ/YP9N4W9wNX
8XtbdZpaWVD+v2VdlXgz7bU5QDSmPa5+55gOMmV4NI71t0MvwUkIDgHuLjXd1xcb
GK9iDXMo0tj3408bhop0k1IyDLpmcAKs28/27QmHNqEj2hlD2XFOKo7i2Z1m2fiW
eG0zb3Vi5FunmfEZWC6oQm4+2w7HVLozm84EM+gHgELgTU+jpwBWxEVYBmptSGah
fcPCLCIfYrWXaXbXUkzBjjinmy/HBNGlU39BtsuOjw1ELOs/zU3BOaApOCcYrm+B
1vhzb7muSjtlI74zHkgNa2eS+iyHA/SPjTVuSUAvKum90DZ1yXZNGXTy2KY21REj
q1NivYnA4mBqv5hGcKlViYTTcU3qDROjD/DXy/Nrw05T99Yta1Ei+l0BVqZyFfS0
+6iAhEl/1gNbTdyPOiDwN7YhmAXMS2b+Qdxg7FsYMl9TrVOJ3HTkn5xEhXFZeVEP
JaHoJjxNk9MWZRZR6eXk7VCj8JLaP2TCqPx2RPFbnMQI9yruzRFrY5B41i8aE4KD
gI20dsRQpoMQl5OPUe+5zvHdxDHgtKPZDoY/Yr/BARd48E5/CsaKXyP0QSkb6oDB
tAHAr1eJNoqLmENQmdtkzWdEboI6ZNtfy6Q9TlTPD7BjIW3U9F8yFWAUl61lY6QA
c8zPfKH5rakLPSEG+bB2CFDl0684HCg5XxOz8fTJUfLZIkdCZ9RfHq5Y9INP4Oyw
CU3h90Ty5qr15lM4WEQaERm29gaup6VqrsfZruzx4CaS3F0yyNOr9uXL2gFeaHLr
ErQoOB3x/s8Z3bUwWS0XrHHAtdOwPZRTlXbdQR91qy8tU8C1Ss68oV/1mPJrKTC2
W0VnRMHPPLbpDdQdrh3xoCVr1V006QzSQLT/ya2jR1JORfkQOcLghO8fddKOVRrk
9hUIX30hFe+Nd1M5gvYPVX7iLDBZ6dTWZ7H5PMtNFcF4LSMiPvbsevQtnSvyBLRB
5dCwCPu7I9CRsSZg68KmjBAh8jEu8A/wNOuRwn7MceSGYuh/9cQgTlsTt/8OjuWd
Qd2B5U2MLD/sz3bzl5Z2TByjFEEziPgmiWdm97YhiuF6iyeh6vhBUklhW4ifg7OX
/zrO0Sx77RWTejPP5G1zkKqK+2r6KXC1P3VPA/TU5x0KQFiLmE/faQ5Y5sNLS6Yt
8XbjQhKrrvlaH874MRenI5EeK5cSmUmSSrziZbbsMFbePUWKhyJkZ3ME9My7ml1A
a77H2q/3SUIL+hLuwTfui5Xj/Q+CkzeiH7GeaORUk2/JPq/a7/+QNrIRpE2uq4qO
CkdzGYnhp5zx14r0gM7rZjq9EV7PpUEQ9kk7TBgGoGe2BGyAIhr0Uf+9cf3NZqd4
21J2ddBhxGlCpCbxLFj+qLrOZuNEdqpJigz7mlLFX9pivDm2RFsolD7JTmoa3pCn
7+4tmQL6+6Tg8MsA3nzFQDByeaD+T0EaDJduAytfhNh3JKbvlfnNEEMwx5uMbELC
JEu9ZbdJu0iU7aSc5oV7LeGRPzxfY2EjKGEx33ehWpQVXh7ZUZ1hkeUPI5RnTfpj
8vQEa24m36LQKKr8CWrMLGBnvC16ETUPb3jNJFPFjFBfCoC0imfeaIKgk5kijJl3
2Id+H4mDbg5f8EKG6AJ7vXLDp0p88YIjN0mif9N0+1tK3GnXY8RL2qJKWi7jlGNn
avrlnEOO/xeJ4+J7XRZ88Loxb9gGk8ox2FmIQQ10pvSNDvs1i3bkUJ7oZ2YM2fJC
bCteOusC9GZ1f2QY/HGcaMomSlOCUBXhTAYatQaIB0iTM187vrF/mfr0lQ9sQ1AD
gAHzDfeD3kaEXyVblIYvREJShdR6E1yPDSz+ja8EbzcHLW+B8AqMty5bgyjurVi3
iLWVNtUgBObKfr4Wd7a+CcqRcF5YyI9Rni6W2sBaaMDRl5ttVYy6nJGMTpZ9AK1Y
im/RKQt5+rzVvMfiuLuOTkhr83OEPlnzn+ZDMaHU6zWEjIBzlIvvexYjx9A8LtwZ
04bPOA2XL9PzQ7g0hjm5Pg3Mkb7coCrWR2+qdLdOMfBxh5wh/WMCw8AuYa1hfMFb
l4Z2r9pFuFqnqIKWlmXDDRHUuyPy4TOQvwJtQfFJ+lSVniDYeUaZxTPSxYkf5Au+
zrwalIucbI4RCzA7spoy/ZMTI+pqx+o5ysNeGd17KIwUb5Kqy6wQ/pAmNfGwu8Jw
ysJgvyiV7yb3ydNCzXkuzJCC/ftEUsi8P+2qpZmqFe8u4nxWJAIXYCt/UN9fxD9T
kuXZlK5+1rT34AgM4hR/qB2VLnYDOJrw6uq2DTew7JyKRpebPflAJe9yk09L23ym
9E5x61/rvTGJecyeG/yImydW+UcaikBLeen9CxU2ANPsySTlvW6enqKIHquQ9Wc3
vrVzVrV01ywuE/SfKRuGPUSHgN/u0Sz5J7oyDmdkk32mJCxIDGBR87Yv7/rHwlNI
+W0kqahgsnZWRfYMlThpmlTxNvd6nSzrZ6b8an/bBCB1UMvrVb7bjW4ofpEiqP4Z
UHxjETDwwjrb0D+j+fe4y1Dt+E6CCSZY29mzKEz/D3Cbb1pOZQTBeJV5VIJmrEy8
5aCWA3Wrc8I3fMExrqjQ9ksnuTctTbOCNiH4jFUhzrQdhiRbwXsvJb9b7p8SFyTw
BRvxutfkQPswfgVs7g+zEWHvsIlkkeZpCwDNAMU8ZqRpBh80T5HR/7rIQ3Eq1a8F
dTG/GXYJjvw0EugVBTqzACNLvcHtItgw643MesazJSucaJfjrFVP/l3N1fk2H8ig
OJETz4FJcdp9Ti6qFdeTht1jA989cqZtqxM+vxuHDP18penbJUpoOIDqPkzOFrqm
BgIN306hY4BJf1c5YSCiwo0XM+3OEikKSuq2Qcsj7VIiN9QNNVNaWy2x6JkES98j
SJrVS/DVMdMwpqUj0EgLFQpWrYwvt5itXScr0K3E9j9j4y+HAFU+tcffJhMBnndt
xM2x5Vug1JkGfoCWklNlveocbH9GW2C7saAXEPo6+O5uWVIKaA8gxLZ98fLO3Np7
64gCqKQ1J73mwkYs9glBrFuCiIwl3lF6YLIxlyrFcd38T7wvM7PS/FeVg43+voce
tFxUGqkWmevQs2/ZHAq8q0dwiGfUTNCLa7ttAqvpITdmFMD+11szl2KYSjnyv94f
3TkIBB50PbOiwZ4doZ/sJHt5pFCls7k5ta4wl+kvZ77c4/L5UWySmMZpE+RgKGUV
JS2Sbqzhd0/wvM8+0+xd9NmPyacD8RHIxowbYb5XJCXoIJ2dnUhSP6M/5MlCODLN
xaaKqRXc8Gn/eSymf4beeyYFcAk6SQ5RWpiz5H/4b5a3q5DnuUwTXdn1b+JbxmOZ
kok2EJyewY1sRb6C6X4pP0aUmzZAbk1mi5r7vkzlg5D8KljhbANrqw+zIJTe3CwE
5mPpymZy3qladKqPvoTytnXtwlopPGzhtporj2ZWI3S6C3EsNfL5HF8KeaZHI7hb
ZSuDt3z+f53H07FuDWCTvpWnn5R13TVb6+NtFTJlyveBdkBiCnK7gjpfmgIeX9yb
ulD8aftTzNRS+IQOvRU/LFJ9DtLG0R/St0n5X279xp6z9tl5X52OoubVknxD7XCf
RJpmjU60hJV9FMFXcvJLDljlO7LUeliB0/uErvECRYH7wnwz9oNuUXTlo+Bsb8a7
hKj7o11BhZWTbUjLFMee4RjscggQ+16WAK2aFI0mKmeonnXRx6G5FT1uptd05OEN
l9GKQtlb7aMOF6fTmTEYxInn47jhGAySyGiyTu4DVreXxiwBM9VNqDKLJ7w/Ud+J
LUvF5odUUFE0LZZOhc2/0h5ZW/hW7dPv/eYGWApe9PnKXdN2/4blkJ4PMHwY9buY
voZ6AE5ceXNU3g+nwy/0ZjDqcG67LYuklpL4ADjE+qcmHJVtjxEzSs8saxKjyQAC
RtRIGChtoz2NPp0rWP4iECj2+hGTvA8cal37x2w56OM00fG3Xl/HmIiybUCKv4cF
MxGLQcMQ1EWX2pFZLv/HKdl4cFanA1MN5B4ohRMZgT5l5TIr/HF6moCLNa6eOCFB
T9RoTdK3+y7/XRFg94kK1okcvKv6ftnV9nxMuR8BxQmWje/xNO4u1sXdvWAh+y61
1732GgT3JMKMy+FG2ZKqU+R6+ehtHXsfmJpIIEbwVVBOrBWEwK3A5kgoi/r7+fEv
/D3G2W0rvmTb6uF9u9TyxFp6kOZ2cmBFNENmm7aGl17vdbuT+pYrJ7aBGFiK+uOX
cTxkmHgPJn74A3j8LKDcpLQsQiRviPs2um1j1RSXY+/albRbl+yul12IfzNwLruf
CPhqXqQ++nULJkKmOIeBG7qE5nVJn8U6xoCuSfKoR4ghq5U2/ucLUvgvnVTj7zqv
YaZJiVnHAS5OUNSU31zwiFiUtiIDD/BwO3Io/h3Fm4T5URKfccWIPr5U5H6fEma/
59UXBwIv7LN+QyA89oNflkVFZQYhI3miyGzibD/Y5kGczJ5ndoan+gnwgnF0zlg0
XYDpNXxw6icSPNW5ce7AXTGuatzYe5h1ztyi/v8p7ZQ/7ZFxULsTjZzPkq6uT9bm
FkJbdvjBlL2RbB25Gdhl5pMShGjT7XjbUB8cz18unMAFUCbgu2pugAmzI4Wry9MK
ZQExVW9b8Pg5cSuOUbl1Ct65SGczN39y/tBqYBFxmnUZCF2GNnsJMQY12BFn9C4R
PYw4pKvMFGTWQsiFFLRd7Ij3P//giM1WBHAy+Wvffnu67cGcv1EfviMloLthgIkI
O6S685kfYD2X0mFqn0tDMLQgx1KePXpILA0Q+5T3LLdZLHIGPyG+hIu9A4ntNM05
TJLfACoxQQ89AwOdR3ikisJVXcyz/TQ7X0E/fLfarWAv3p942dsovG+R+QRW85C5
Xeni+EEi5sZNV3yFaqYn8M0nGi8HOJHphZjL7Gp6i6c11kQrmkgWgrmdGa7lxzvQ
cauIh2ejBYSYLoUBZGXrJsy3UVzDUMfbF7Bhp4U3tpeNcxEbM8C8HaH1b4bywoGc
Asf6CxyRXFRsE0sftatdHgKYRwGBUBr2U2ueXZEz7eNhLUrWHpFD8sKfREBNqnhF
c8KlHpXhsJCSCuOGLbdZJr49WyYZq31uYm6A8jPRTAnCkw9coGmQzzWt1UscpXFm
oknd9P1X4JwP4Iejzhkoh6VrXEr3a8PUEzu14gK7uS3USNmOZSVHChplJg6h7p8d
TWl9LlsZwoza/NCXIXcYZl03VR+2TOzGOs2qlGRp04yEQLP8TopLvhG+W9eh2SGH
Z46+OPJ+TACt4qVyMpdHMUYdhrN7EFpM2O/onCIfV0M6JW9Mn9Zlj40X4iBqOywZ
JWCs3wbzhSHyp5alLB4Hg4/n56vHedze2jCXUilXC5MPUCbLb52bpqXY/rVzuVyZ
mcpADF+ziXUAigzqvY1i1/9+2GsvBTvdiv0sLqYNMY0jNDqAlVQduPeK1jD4WFzb
yxpUYg/EygKrMLl+X/YYLtHsjc1oNkDmjQPZxrpKvrCkQd+ZfJ3g+eJ3ndjwBz2Z
4kPU6KcKgk3RkX8XN4MSl/yZE/h5cCdV7RLyDY9jrb5qK0FFKDmOKFHvRSb7oyTI
NVK7bC+xXJEBgSDNIg1HrjhKCWSKExbWHADppUX5WBeesKxRX0RgMGjcSGIigdSs
qU4dPEzeRALYKis3q1x/tA6S3NEO9sr0Yc4A0zk8LA6Tlg+E61FPJFEiNvzeVprD
Vp5MS0tVKUoNeZa4hIrdz60h/FAT2Y279To/RKHTY0VDPFHNuvDczVXpScMy41G2
3ssuE1KDwwiHOmaB7zSQxTbV26VrIekH8eY1BNwsRH2jrH9WciBHGBGb5BUkJOM6
w23ryVm2vQxWiupa9qD16dfdCamqf59uOFq3Pq7cPNTt9OSi8C/sghrJ6/KqWaYW
11eZnDhAlG1/XU4QNRrQV4mRY+50eYxh2rpEtjn6/HWRjKM08fTOP0kTNXxeZtpf
pWLDUZXp/0QK92ik2OyMjcfxYAYf+xQNQEZaERJvvDmNZ/4kESLaaVIQHKhmRq2t
INZRcL2HsUMSoxvKWq6QPDt7M6PEakt4geH8eFiKeBgqE+L5/hsJ/YMzjBGmz6QX
aziIn3SMcY14xMkBNOP08ajCK31b+i8O5OkA+psRYRN79srXcdA4ewqjIPiBmxnF
Z/jVINXwkPC/CYFbXxhJacuCOitUgcGswpXG6EFuZZ1L4IPNavRsXr7qQ1xkW6Jh
l6qXjbgIIpdo/aOXe+4PDR6NrgjmkGGjY7GUq+1b/sc3NO9KO8hJ6oaq2vTHEkFE
i3IqOxCEOrB+l4VlIex55RWxfUhLH/S7iHWJimIv0Vx4ct9Xod8dXs3kbsGg8JsK
wlcnr+1wRuGYkPnuPszv/vtA2WYeyU4OyHfU5okOzkKmiBpR4JL65LyuctMa3nb3
7nwNEuGi825ahdakBpe2n3lZgXnwgv9pY0bpnSw2wBYL/2zTyZGIIMYQOoi0W2LY
UWPh2zqW1jWNFOARWZbvjjE9q1WHIG22cLgZSdRZlv0k3587bB6z+5AHZlU2J6vk
urHC1RCyajaOcA3Z2ZDYdJ2UVf0MVr/VrlUmt92IzLx3dz2zLi09RhxM16Jrp0Se
sQh5oSZnbID5oSYd3AI6IoreVSMmxMy8xdhkpckdeT69+jqbEkYrHEXPvILZbJuQ
Sb4KfqrZrjXrzAqpVWROvYCngYBMIno2E4wq9yOB1a1O5TzeEwVt3LqM2Arcjpip
7Xvtqf3I/vzVG/ZO/1n35IBCYBo2/qVX1sUzMPBulScpuH5yE48pU5hLsVSeaXVd
tVTq+rN8mC0YeTCguzFw4DlKFHl3u20r5nE8UkONgWlwFO69svjqz7CYtMhF2CcM
97nylG2cBTlX6loRD066/W1hDcfOKrwoDk4UdRl8sEOJuU2X6kexb7uVwX2rGy3Z
4Te8/VmT5+htVK6U0ygTuJ/jaUBY1bkCizlQVnqy5CSi6MGOPE3xL1VX+Jc8mM4k
AFeLyFOLABvCICoTOh3+ODYmRYxvDGYDusbQhw4VjBltXhWYkcKvr6bffHkxReeG
492Ia6Q97skvz+xYveIa9xjUc4A/fFTmJUZwwGkVEMMP/RFhnyoBIBnQDZWHD/1G
jO32QOqMvYIO6nLxMu4GOoKcs1PbwrPBU3UaFLOfMSIfGrVWmH8o2PKLth220OK0
0bPKK5edUpm+yPIxVlgHf1xSRkKYfwVTY8xMqUDKBz2tGrkaP72dQqC3SuFJg4hT
V5r99tgslXQpzXjE7+aDY3Oj6LlbDyfFy4vhGUI0qXpj48g8aCv9d8+Tt8PV9l+N
qJRS2JNPbiwKNMYwvKslVEbZTCfneT6OnuWFJu0950Ib/39xyqCYokpCMgO74Ggq
yiHMfO4gxCqoGtJk2ghj9eVJW9tMxL+vFTeagS2NggQEbmXOk8ibwOmV1x+SygL0
gLSDSLxS541hYPdm8YdRBCotdHBp1sddOp6tMYIh1PeguVZayM6UOQ/yPNNmEIkF
W9Vib5+vbS8QqYiv23ppuVf9Yb6RA5oeEoOOjBNn7odbng2F7bUfUICzbPoR8VWK
qVFx4puUBXyO7UARJANY4U4fWcGhfI2sDm0e3fXsYBFZ4LXFMzSJ4QkiwEIo8aCv
ul+zBdfAKrEeMuyifFIEpjXSXFhybiFqGhlkivTU29QbPl+B7wbHTIY7GjduYyae
PGB9CVDGfIuTszvbZamSTVpsge8uIFDw7PhAzL37NQCW0UieoNe7fK1CyWDqpuNs
whr5p8zyDzyrxKzZQ7HxrvBP/zw9Bf3gq7MdS5p5PrhPIYku8RuY/WAyxQMXPI+X
+COk9kHFrkK/TNEg8lmj43xmrrwiS4UTe62NvrBe6wsCNfTVAd77byI/rbvBbKP8
F1Aod1lFXBjh0/YW/C4Bj3h6JEvAN+TjxfkN0YlYCpmaiJ+rjocUnYoUl9rsxVEZ
6XIkmy/8YV4f1JqjE1cICVur748DeEidnyAzeN2YoFcEVT5aEX2KbEKQAjoPmWkO
TP6R3raCCoapxdkm0Hd7Mg3QZj3B70qKPVFZqjiTP+FtJ4yDv3ZaAyfwlDOetH2x
PRw73wSfWnuiylTpR8StmhIT75K6Xnj6xdl8bU22mkEnGrFim7GLIVeU72S6N0/N
T2aEIkbTPnE4pChZiysm0Mk61BkJ0VasNK0tYTi4VG8/vZnpNN/nfXZ0qRNkRZ69
3dbfZkBOOXtu/CB8Bj1u+m1rq4erOqSSQH81CXdmcd38RCQihdLiX+Yej2JY/C2O
t2GOZEKoxShOODv5zjVodX/xZEn3PK+DTU+f5yopuUHyyniFWLOGRkTiK89K1d3p
uijp6hCK3zJ2yBVkO4UbFNABsVhnEeV/CHFM8MlBQDG2vyy4WR9yfsutxkIZx7Kn
PPNqbQBw69s1fKBF+93uNueIKIP9mSXdTXmQzVOQgUbUd69C8MytToq+GZ6GMJA1
HCAFT6hVlOWW3mdLc4PrMjdHimxPrjPy0QfIyxai+Lhp7reus6QC1u9hjrISzLsm
nY7tiaw9hmBjxyIJvrUDYpbP+lW8IJoY4QCMrdrnFVhGroXW4fC3SGoM8tsVszUA
kLNJ6ex4BvgBvxu57g8F8N0Xmd/0awbynDSpS0Lcfh60FvM22149XMlVj4euJS0+
aSuYQTizQyCjD2jq0s8QVt8Z1LzqRiTtQmMWjUb8ATgCb0rgJ0nQee+ybxfBmGiW
fXuQiPuCgS2xhT/0zPsqcyemdvUMJoBXWuCiNmZ/bOThlRJr0CGp3td0VJ4+XZKD
2vXTR8KhI2gUMfjMlS9LOrqY8OkqsdvL/orXgO881wvCOh8shub3b2AcxzSy/zaE
9HDjruW4LU6LLIJfdOazkAbiSznbcHv80bQIns4i2ZOH/0VWzJQAMfMSMbv0JoPx
XruJ2MRSp0DWYE8bOYHYt2WaqhT/BLt0f2+yjvY0fThNQYZ5qSh5Cn7yV8f7EzkV
BjOdJpuLlCePkM1M6OP5d6kG6GPVAIE9XbHY3y1nImXJ/FG8u9h/M5iS65QJGqRL
ZvkGNsGzXQHlvmEsqVYPyVgFx7UArx8DWbOE9f0FpiTFn2FFyksULrOAD2vsCCqw
CmyPK1qIX1qeSoHf8RqB4++ux7m5JYwUK+QHhdh6XUBmzbuw6n5/tDl7kQQhYDXr
EnwzzVdKrl0fvaCkUK44OV7xv+nAJPcPjsEVDVLpBcMOpPLfofRJRXD3Ftv+mofV
jJjtAzA/g/ZxyDgIbzU2bllNnL2trJ6RQAGJ60AL1QZVottpAcVfGvTLhJ+enrAT
HYrh/cIpjPbp9OXT89cFdcMxLmPcqLQQGfxfM1+9RgQnLk302wOloJIPEW5rpUPW
iaaKH3y+EtLkuC0Z1ZpOZOWDvKWvGT+/YlqpUnMLMT/E6IWHTpo7ZTdJe8ZupGEm
kunZdsfuPagPmvaTXRiop0a0J5Mhit48bjVhMM+mVnX4+8wGv+Fcfaumf/etxVu6
0emHs61gh+yUEZuextAesi6b1MvpvBdEpSgyqEciVQj4k+HrzvY/6eij1DC9Cz69
p9WFO3MBriek09TqStyR1Iv8+/dRkoYph2P3AolOgkC7oWm4gsULM/FZvS5GHPjP
SVo/msJggTNgVqFnR0p0wILBzjXlcq+LMIUtg3u34T8qw0xZFDQ27Kkt1xeZBrFT
AAd5COram5ZnZ//cTSJxEsg+dpCD4zJMw/GEgKeXVWX6OoEhSizRizLV4eQEv0VP
kZkcT4LsFpZC0r2rjf7/czfkNJ8w/G/cZNe/tI6LSq2PS3CgXyyapJiBMNWJ2Mr4
6o9Ka0zpOhZwuGGWW2TCECnE35vFvGibnNoRe1sNatkbaaayr9DYeGPz688HjH/s
DBYyOzpen7hwdH5tEe+XS5YpbEkkviyI70QpKLPRMnAlBKkoYTUhHCdLOzO/3Onn
7OQAEf9WovT1/xF7vD1EpIMU9FkBhfdLAcxFTgwa2T1EVVltDxfRn5YMQxBKlird
4zaP5+xXv8muYkCqYCJYTcZ5rT1Y2wqFPdugVE9mYykP3jP10EkVYbEWqKHvhO4f
155/T7N74HtJzswrjr4D+3twzgDtWO+9j0Vx+m+tH+Ys93v33tJqK9tpizPIk6lo
eG9rejyZq8nMYCuqlAbD6pdGMUH5HbJoGtRs2XSXwZAkLiu+VaEWY0u1OzU6YWfh
qQ6CUy+zXRMl1jxV95o5XZ1rgGimYvfqqhTWi7UHOZS0QLh9UGyD41stAbrUOapA
iukWf01R7rRBsV94ylKynuD3BzafTZFMGzgx2ysoFWKdxXTRCsoTJslPFx7E3QvH
Dlf1cT2lgHZCOK74l0wtM1nmelFowP5XmB8eq877zstropgARVwhB2yKOqKspmVT
FJE1wHRcwtq9FSEe88vPRnJVb6gDMXmWfHa75dk7mI7Nyk1CakXDaj/0ot/zoji4
Zi7sK2718GSe0SxZhZsvvqZ6FkNoEA8R+4jgJUKpKCDaHwEpm8T3RVZcaWenqbxj
EQDWRQZwsqbAOyAj+zioNj5rZeW2D3EuosEXzr7NwaLRKEobdApjmuk4JkQpcDZd
a753aRGi3eKGk2L1CnjFd8fC9T4yQieUHtLvjTuYypye1wLVBYxg3MzGQY+U/Sm/
IUgWJaT8fDQr4ywCiUIqvhi3wWxD4SfUhUqG4OZMlA8k3GXhFP6zTLM8nGT4XNUt
w6Ll8vd99BnXxhzH3A3QUBMQ4viFP1IN60YLbsSA3Px0JvY099SrbYc6usCRcy56
q8D6/zsXl5dzuYClR1ywBGnwziq2uhxPEFMmG0tgnnFQT1Dcsk/8mVEH0Feh7g/k
HlBYcGHV7rzKuX3M2JbtcxAIKjCVZ5kTWN7HNwdIPY3yEo2jgWUVylG+4thVu5ec
OzqYpDPGAU+qRREFPoReXpHfDWwwuvgZ3bp43LaK7FXQnud8oOqh0R428DN8F+Ef
W3FXc0TF9tw00BVrPFWyYq8zq58g4tmTmm1E8Zpb5b0hzQwajx77vftZ6Xzwk6GY
+1twyri2Awm+4FE0bKpQYQA1T/G2cD2LRqQ7ME/HavtANdzyoA+2Fa3h7olveESM
HniYq3DGOpkj6o04CMYdCok3cDZmDVgFqXsuXtWn8uBLFu13UR06V3QehxLUqlX8
Yvn9LM+xvEtCyFsouVSo+CXtRta1mqHYywZns9s1bEqE/yHeHI5Wux74KiwKVvfr
pKI3Pf4LwqkoFfcuhsNclzYoxyC00jqqeYOBSJOZiva9H947C+578QiUnfzWr1hy
U14Vl++LC/M2xDDRKQ93R39v6LZDTVZF7VCKtnxfMLF0g97ja6xrdEqSySIctXWx
8y7l1IrSBdMFfoUM6AEdHELn9QXpAWtQrUeZEHPtvf3KjbJ1pe8XQt61LAk24oOy
0LH7YS1w6sn+PiRNdDDTf8lVw3yOQbFQI6+lcXzBxJJqtJ+wpa7QsTgIzBBuSB+u
3d90ivZTX+ZqkwEHnv3L7CDrScjnEERDJGtgJ8AlP6eCbWFSn6hzsyNE9aJnI/Ne
7+m63m5FgvzveJYPe5odjpPyTmOoIjdwj6ygRWKU0eXcSczlAF06HtRRyXx/Yokc
CEW+w+vJVJ2E5+KOyV1zoBvrt59l1OpWlWCSR+6Z2ThJaWvyGzFOyY4QDNbHvRBH
nFgiPQw8ksCJ03nRrHhCUuTdZt5NfTgpgZdqTHDur566LjN5wHbfDBe8m/Ngr/4m
t2LJtpNJapxQIHiF0OM6XWLvwYDxKoUhoqM9d73gt9aLhv3XrbDQCxVwJK5a9WNA
udpcj/X/tMOnllHdwulCPhS0LU2GhSBSR9RUwrUxJJKBDYyYORFJ1D7gxki2wZdl
1bHPBDErR/GufiwDc9uGoCFF5SFqA+e+gB4GJf8FXZeXw4ofIH/RVw4G5oQ6nRIF
+ndVAimYuQhbhRTl2/xFpfxZB//tZ70ZKIAflekkuvJBep1K4E+AveUVFpRg1Ub8
i5NazoItYF/YdHQMj6xxotIoB0db6GLT1kk1bIfSs2B9vHj1dN5nG/bUFvX6fQwd
0Mg0vYuHJGIrWtCd1Wna6qfM1bUm1U+ydyNnS3SAwdDSK6gEGEdQO0O8ncbZwva+
p4zF5AW8bMs177t6RLjs36b8jrRqqwvqyP0+cWzGHKeRJ6ZGj6Xq2aKRv5JG0bEp
VsIR34AxaO0FtvnGFOqQNXuyM9GxFQLnPPmWdi7gw/xfiME3/7rnvckq1M66k39c
OGmRbH2/GBClueTWTOm/wBm6F2mYt+TjZY+G9MdRPoPAlhxUPSeQIJnJ6ahFa4Sc
bNUYOAB4iHrE4qhdlpkAsP5qSW+UKRuVGsbArnBKiYBdlFoPtP9gB5KMzEh51Hij
ZmaKxRWCBeNSkdjOtC6CmyvIEpHg3Cpf1hFB5LkrGFX6f+8jU39n/Mxq/AeW0J+0
HMFvrvGriQNCUbmJ6Ci28AEa7vg4UWUF+LRSIzSf6GbOv1KmHLeSaiYnCQZnrt87
etUcy3nvo36RVSpWdqEzxi1uatMIaZIpYtQtudL+snyCZslMO3ukJ78OHVD+zleA
NYh8qyupKf00DvmJgsBGOl5fuveAq3gmaqbbGNTdvBCtdVpvTDWZm1KMMEZFmTcp
AqM8Fz9f7M3aKck9yB2vW42nFo/VV1VWnoNPYHTrAs5d/5OwmpbyT70wty5aHfFx
W2OtwudGbrg+x7CpM+32DQMRl9AY99rcgdWEn1VJh6EjjcLZMuJiavzGGtJ7VZ/O
YM4gh/W0wJWHl4kYgqDcxiP18BXPlkSOomgPVDRhmGIHdumPrNswkswMa7PC7vPi
PkYP3+NJSTtQbv03bDGSMLbNbqEyJi1IMWW0til4ycUb20tYOylivtmkBYHcPb5Q
W0wS9NSRfbBqqeFPJK3YSTBrYHMYABU9MTJGOT4SS+EYOcJxrkQt45lWhHMu0RV7
aVS9w7+qAuxFCzrmgkudZ/FcdvG12UM9QnW7WjEJe639ad1rX2NwCojKeo3ybpJD
H9WlFYcS332BF4t3Mv5rCcogB1I2IX3j6AzzMKgwx5VSpBRkPmXzDZliz8PObHmv
uVbF1sPWbnPJnthPnncP1b7UWGo7NFBJ6fsjNx1RFLjHCqCSkN88Vrek/lhChmt+
M+iVHPdJDuspsNW8eEPXhLJB5Vr3JHA/2cBunbxEnmqGB8Rd6A1M+o7uDJ09FZm0
X9DPpxeIfCaPjUXxdyfIEwmC/6x1vTpM9tRfYCsRXbugNGNWNsuTFEqIGkddSrmo
LdghLo0mrqX8BSwTI/jX0onDVhrjTyBV7QdGg+Y/lUO1ImdSfx+C+9cNkA+wLsHJ
59BmUspM2SXW4DEjIt6H9egZ7RPX6bL2bdFkUlD1tmK1rlE2d0SDBxRYz/hn3iZY
WrC5NDHe7T5FMgru02uU+EMRYwjJQ8D6l1Zfvi0C+EpiM2gHB9JvKeJsia71JuXc
vcUjvSUgKeBVKtQnwSYbzW9opbKpwoIoMh2hfAL2wKxZaxuV762J1qAJwMUYaQoa
eN/zf6ECH1GaSN9iTO6GI5NaUSy0CNhz0LqGPpGLLfKjSTjFdY02grwf4ahEwa+6
lrYKulRKBvd/MXBR8lh6MazEQMIfMlS/Q46MQ78kx41sV9OSPRcSpBjMpEuGWWdT
qROZX79Nok/JZayL/oAGcTS08YgvPdmVniD7CO0Z0k0R1SswWzDKVo/1sK1dyxS2
ex03DOAdDKiPsQ+DyQiHuY3x1hVzHr7c8S7/zakT1VQmU4v/L99Hj3VUzha/xST6
E6/YZAHaMKmR6/jwSuQKPlrEBiRIvKHuENvr1XNDMsGZNt8Eu1XVjxB24bxt6Gl2
NzvTxnq4DDbe7tHyQJbm0cjA8Py4l/crTpiMATyO0/nWTU3youcHnynusdzsorP2
k/CTzp91weH5ccH95xgITS+bMAtJL9cB5tFKK66+cUyHxOytmnXneLXcl8XZMi+W
jhxoXPLwtcOuR/IIINTeI1QR6+t3qeSOuglL3AF6ZdGpdadHDM20Yg4Ou9n5xRIJ
d6Bvwsf/0sPX7USfN27BNQcj13F0s8EgOdBVQbNPJ+RQPeEgyKXIWLsSZ4QOaeNu
8Ltg0mjqJaennUv764TCgdOOFHfM151fxoXKY2gI1rTFT5Jx+5v/zJ3twsI36KOS
oQVOk+AIvvK8U/5pkjBnqimF8BP05lyj081ptCrRe96eFJ3OiPONE471j5gLk4Ir
3X8BkApwYRVr/U8+i685tzhACE4FtIKMM+riM2ydEedwtUjnLdCstZtx5cd58IqD
z5hD7Ebjlf4H5uzXLtUnjUlgFnBqkR+6EQkWAOEW+oHvaBGPMwiAt+4i4h9NNKR+
GHyyDRiP9utKVzQ2iIMqzBylfnQ8H8lbOQvOYn68jYsLM6NvL9sfEuu/YQBX7szM
SzuJRTOvXC2AugjIG81SpidA+SIob18Y4tpRlChFQ6AuGKVrGQP4uPUeAQxWBz+s
14x1TK3Iwf3Hl+TsjLOilUpPdmaO92ALUIb4QhTfbh55408gFt83a6YYWpI0ZS3b
mAXeyw4Os9viOeLA0OXD4q3EvdGzDimrSNjoLkuLER/X6yWLoCReTl8e3b44Fh0h
+2AZr8lNpl9CKGya1wH2moOqhI+xnElSycKaHkpTuqQy/nNQhhdjnvCBto4t8J5/
jypJreI/n+95NY8yLMLf2J2JWcWvoS+43JUFnbAgNQkEHgf2o10+5XXh0az8hhEy
R3m8oESxqQXwFCmhaFoozQIe0w9tOGlOb/F7HjX0IXFbrLqC4i5t/um09541s1Th
UW7LXqlL39Q4TnGUkZd+kPmuTL1+aOZUBhww6vHl/R+dYrfr5SFGigsXv4CJzgJp
lu/taDnDjQgL8UK9/y5Aed3QLEPj7PKseFdURqjYE9K9wI3fsr5WqDDHIND6uKIq
Wg3NeB9cszQKZHzsEREwCDtv5VQUZYN53AykRAYL0KlMbEtuHHeXPbixqVdxlHBG
KsU5CYqMkPey6qsoeN+JKv5NWu08KtT6fpfdprZUHeEI7tSbouYT8fOkOQyPzMnz
0/jw+SP5aIACHY024eA5UdeQLSfkQHsfakHakFi8MzqDLgCxDk2cGXlDXQCUty72
7RtzwjDVRRCtirBcCnt5shIcl1NkGAwki0SHbQ9GNPAwJ2PIBlNFd1G00KosMGxd
6alaXKRKepuAjmCZ2dxYgfSPF+GkWkK7IZK+3jWdjlw+tciSLifikZJZLMbJGnTI
Puwbe1qzl+eJzv+OyDwz49WjNQDaDTCLBhro3NbTwA5Bf3YDBPy4zRmBsJCu9woz
hkyrCXLnvDpsCGUriu45rpSsi/78/iEd5/FYfaL4foYMSz2kgvkxKklLOnWb1zMZ
a6gnpRbRP1nIsaQLrs4+VVnSAYUEfnXK5lDZe9JshQRDmVYQVMEmQieHeV4h783m
onS+fip4jDIk0bWeyxUBI0ZzTvJ1bOBFAh0rGz82eX7EVvhOa8B6pI9cvCKUwXXS
dZiSa914qF+Ah9ygHlErrDjEB9N8uJEXn7VbiJg91ZOmaB8TQghewqpQEAbl2che
0HVoUxyEiXGp9I2Em3JdyR8TeZzBQ9SiI2KYlFiSPokvCpJp65wppkSrI6dBzega
b+U3lvfwQedfY+NBTzJ/+MGKVxLpJ64FaySlHXNxoXcZOD7mXMnjq9kN/YC3+uRF
rCrldKzz9m6tyl2vZyDewxdf8NNCNiC8e9is0hBPzon5WGAlyjFCJwBfpoj/76Ae
l+X0Pn9SYboJ1HHylMATV6bU34LqFZssulNf0C7skPpOWRYaXwrsWrsIeoleq98P
ZR8ds3JXgP7RY8R1lmY/nbqS1peeUpXn2esO9V5EsSC6baVWzUUisLNSSCvVox6f
yViW1V8GPlCTAed53hchGypMxvej/EQqSbUPKZmZvaV0idqyTc5HmVQMbOOWRw/r
KicdyEztXeIe5rFF0Ny/lDe5DiwWSuu+K1t3Y29QBnxBsYXXp1NtaQUXxK9qylJS
rZX7PLhsz4/iGcatzSDjEf+IMN0F+sXaGMqBK54q7AmN/3RiUzNaypho6Ci2k2IQ
qpUAKhmv2HxTFqdrFPJ9eSK3SFZuoDcSxN4TAi0UrIDirP6VUUT0AT8huRCoUdm5
+WbTaix9kmIEbBtgobqr5eMW7lZBYxOasqO/4gZeL4ZiJxJM8xM0UeaY7xQi1TqO
e2mVfEuG1ZVMt5veTFs6JVuOquqeK/m5BENQxTU3kjbAvBqFrseBWYAch9Vlrd4L
vkLBgjsdbQA7Fz9iE0Kw/BLUdb24Xo40QKg0UzWccY59sA/RjuPW0ENgaZA/pf+i
gGuz+cUNGx/nQYioDJVFClT7ATBxI6Ur2YlvANl7CsLiF7KIOPNy0tz6j9DlF+p3
QOMhBqbMI6qITHC/B6eX4KKYYDZYN0MOdTTMLmWTjxrcT3DQymZdCDg/LXRqfa7a
QppAT1cAMoo/KL7lFAU9qGtB0YL9F5Qa0DX51KIlOuNGYyWO/WudAH+XE6ajxyCn
fvwVppiQWhyXLE3oOW/M8l5epFdo37VAugHbeC/y3jJIVbSSp0RDGdYl+OPZKCri
UPwj+sDCuUExDetRnf8+WpoAklPeNC7PODvv1WCb/7bGGfDDLs07J4RAeHDtJzkj
B/u2GpozKF08Sye+P3kul2yUqg87dmPO9OKfri9eIjft9Bvv2hU++APFTVnYcJl0
PdxDC1NYwPnNcGojlU6K/fFBklUQCZe9bKyRcwmeK7RyqSMWX85la+hTTMydEfED
b6RPCKsD87pKQwVcfzdiJZVrLoof3kOIKRD1iiQBrQCO3n06tzSv/nrV4Vks7IgE
sflenYfgZ9ZP6Pi0Tg0y4narie8IbMOJuJJd3TfEkUZQoZThgII77EwBwaUcDeTw
KJivyZqgN6FjZzpoad08+SzFq+5NBY9Pp6g9o39rf8iXGoqnQ97y/etnXl+bVexp
fex8AWWNz0oO2REQmqWB+WKzp188Iz5uq++3s6chLbw8Aj9tENpWSxqtql1GlZsc
++5+DzTZDG0UJ8gOv8Qa7g8/HFwI41K3giBmxK/tgOnttpyo8sg2TUhWsS2z/Jyc
LIMlFQ37eHyPceLq1B/PT+xmaDXTBF59dIXG0YEPBj0zYuKpc9RshAMha3qdPQMj
zKwNZortgrDeiS6looSB6Lv7tTo/nKfAzBAZ3Xvj46s/CmLrCT4NQXoFeKGfCgrO
koR+ligfPTRJzD0eepOEHDOD1sJAACDspk6TYHBbyDWaXmdTj99Ei80EPd3W3pI3
doYbfsPJo9Fb9CIBl7wx4lVxdfJi3CcjwxzJqFdPPjYu9CvQYh53QMjBbqbnziLM
NlP4HXziZUOJR14gsSDuCNJ81gjCuvl53Z8uM/bDRM6gokLdrM1U7DQSElxXZHlo
zMxIqa1H8uecgo3YgEFEiL15kf2PFvzdKGNqpt5ucZ0NywlyeksgBuxlSH08eFWl
vN8G6d+xcCW/BZwQx9ufVbXl4NJJwoVEPMI+0G5hSVqrEi1CeQq4wgTaWzMY6Agv
esUecjwCBDYMHZFZnDNAxF+p8QWN++1OWCALToyCIBwBFAvvwZTfNdxj+qG48AD9
jyxoLg72vcYAfPTPK1ScEMlO0oJmDlI208Y0+iAYQjUfQBUZjtm/FsZ71aUKyWMu
cjcg/zhr9cgTEVw9iAhp/yIOuy0ydaAuLe3s4Q5yfnCLLbrbgBwBtBCBeEylpaBI
3X/GmI+oA/oTKT0IMGil3HvnXNCYsFVrUadWQ+AVj5dzvNP8SSWnh3o4qjoodt44
61nnBFw+KZPfiusAKu5ggW99JFr2Ig38xYTI/GRbdeUMwryMA2E9L19NSDaQIkCS
W98NWEAG2q4s6RFg4JYTtoSdFvZ1LMQjSCB0bB+AGhRDMHwj7+vNCqIu50C/8Nod
Ry0OcarM1mMl61AdxpYdidsilr708i2Pfk9xi8e7I1HCo8Ml1liTEA1aJlCr2KUM
9yg0FmIN4+kCU0ypKcX70yzNlLuFZIb/KTwq7au9xeYg9RciYjvxMV+ievzEl55n
ctrMT8qIsA3lXYg5Y6t0YXi0OC0uvOEC59iMtxfU6BU0j57JkGee8770nioLeqYY
u6hyq6MxRIn8uHIuVVy85bqnOYlJE+toauyS3TdL8klNwIlG0HNwCa6COqyd4nxG
wjxgbl66zEXVa2KVfpXM3BMgjegP/3r5PtCKt48labRrdxmQhhoY3uQv6iFBfohQ
eL811SfFdgJuqoLigV1NYCoYUgmQjDAx2hCQo2FCWrE0c0wHwqv5dbgtGBebXq4Z
TV+PH/Jg7j66O5vjQYoWEvsjc0mnk3V0sfTZLApEwp4w/nNK1a1aa6uuSs5kesPW
NtnF5kmpDVJ5+EgouLe/Dt+O5Eq42azU0nn6vo2Ern9Zbqos/kTMCM04s/2efzh/
G2QRg1vs7/eVmJnRK8t2Sj4/EZR96F80jxkyD817K87V7Uv1JaY+0zMVl9Lif/d3
8mYGVXktG7IUst+UJLSvmwQjca1tJq9cLKVRfXNvX8TdJxdPHzrZuDkIIzvEBA+6
1ZVJ2ZQx9DrSciVC22g0uCr9n5z6gixSv3Lc+hIdqYUGka3WZlRhkRipWvmLHTSC
VGZYtxH/uug0yExadMmQVpi1tU30CwiaAULu7D3rWCuDtdsdaxi3ZVRZA+dgx9KY
d98jopn+V5F6IWXzKWtifcz1MeOTrUFzgSdQvNTd4zd/KWzNlBzsQtg6ItwuNGRl
2vusdQTYW8vU5O7MuJbMe6UPvoMZrt1mVjLzLQwnmEeLVeGlgLZTnyItPeNZQsO9
ihZrF33EqFIhoncXoNsNDoe/rW9EI9h+GizbCxyM+4X6D19fOWJK7xe6cJj03R71
KzMV8qRjpC582xEHXb1XRcFX9pzp5I3GsJJ5EmjLoqsYuhHOfafFlGFRuuYW3jsI
gug6Q72rfQIKl6zq2jlKzk359XWz1/D/LzAbopdC//iQO0M1RMSU15BT3CdjsAeZ
OiRwkGlOxb6U/PTrOy2SKNsuG1WqHh8HWyPMGzdi+o4CWLSlx+fpJY3EF4WkjdQh
c8FhYLhJc7h1OPP1YhA4zOnrb6ItGDIerYHbGL38Y5x5fQURIgdNx6lymxeRD00C
PuHUaLwHJYNkg5oNiE2KNO9J6pL9+GVpZQC0h2xPO8zhyMY+RVo2Yh9oFBL6AcId
qxu8OiChsB49RoxWWARxAKGD7aVEgmswkk4EDXa2p2SwLUBEufDjQ02d4qq8u+3O
qUfp79kHDY9zIM0kpBI1F2tiu3dA/6BnhTA5qZbRTVjyuGsW+2MfFoKrssFpFvSG
WL3lzCXI7QxVoVCQWDiM51AVhRT1yPp28LSZ2hFak1ZfOGZ022UOeBsWngGRzukH
PZhPRjt4w/wpb7As18eLGS92oIcr11lq5Ll/w4XqB5uUrj41hyZG3zjmaQ3kpgew
i5A6634LObtbM3a6hY5rYj2xcf2AQDe7BIKgQk4zXI5W6htEItg5TTvdtizHzpsh
hhF7CESHBDnkrEi7ngDQ6MR9SvOFekexUk2zWzWvJsEcJB6ulNAJrUNnEAupffma
Y1yXNOeHdlpIMjNg8RETbtPaSedwfo1L8Xzvs48wA/QG9omvkWR3byaf8VkswN2P
HDJszZd3Dn3jQ41/lO5RYo9MkI+yvKuOfqSvmz+fyDXU57LutrtUMpMa0asQGEFO
V/ynGYWvpF+wB5NHIQlaQsx/4xWcYpnljkmh+gwoXgnuc57mqpibBA37k/LwjR5/
WW+WjR6zLo2wOqcq4r8NQQNXjbuFLaXlDb2SISmq8QRBI9tANCYwokBNwt6TTF0j
eRxy7WKFg3bXxFx47h74rXMZLpgoOmyESWgw3Th/94jJJsWK49bsHtpfi6PINq69
TwiRFXbUrZrBQqnf6eB4rjRxv/TWbxD9c97BmAnwL2sNS2bxsywBtQGYJkGNXRr2
4xrscnxnITLELvyG/Qv+2HOlrgIVGQrnCb9o16n/HWqaUGq7SiNxgVX2O0WDtk20
3t6i3QA5WiNItkjvRRvLCFjNrtS26ItYGWo2QQFStPnl0kMuYIFikAHMYVjDyDyP
1sSB6H/M1XXjXd+VG/0lbqsbGQ1nv3zSnSMbQH8zBePX7yu6DWxdQsNnmC6+0bvO
difFWvdI+Xeb/bMSmlHEvOMgqs3cd08k9tyU0ZqMr9CKkHxgWEHTrsAbyRI3mxS/
BcyxQpGzROaoUxnkmIuayY0pXdvXhNhg02hzULQoo4xibEUXjBuwo1EQMnVlpyfH
FUVFNm4XCgR7d7EoFnhWkOo3uKEtdqu4tdMXSgo7I1clTjXSLt0tUuiDRTeqS9eG
7CDLmH5fiZDDbpY2bB0PB0f65SXrCrsRyAqFblgjeJ75iCRscsScixNjxy4L9yNy
qjfY396VYEr317OUx/p8uxr5KtsveIKotch06j4mfNO3WpYMnBovaHfk45fCnk/w
ZFQRgBGMUP8qcrcsm9takK/1BHcAu6psbwec/+iCB2cUt9iNr5h5IwQoZxWFDJ5O
7QTgeJ8wcITUkdgwnxYHvvxFsYgIkvnezPa1KpPLVUIai1Zlr6m5CP188TrUNryl
asafNJRJzJt1wkL1WsD7BH+FCW5o+QpkPYbEympuimXe3FUJ02oDan9NkkkzIsVZ
IBRkt+Dc7zXnTKxf+vH2iO3f+r1ts0qxxVXoF/bQeO6t1c7p+VQXof9pFbCS8iic
9Jc14CG5V3BXHQLDt32mPIQxxKrnP4RB9mNH3WogNZGTUdtl63NdZLtjAXFq18XW
OKjbkLe+teorEK2JfaocJe/KFqxGR4bBenxLnRJOqb3ElBVJBlTuq1pfowJ1sI3U
HrRymtgBx75RLnkIGa8QzBgvjH2sK1fV4FeqYXNTFhwa1E9H+crQt55Y0IbdXjI7
R8UPWxzlzRTJ+ycJfyboMNF8ymyyCVgD8Z1sVRL6QyKCZTXvf1tJ6DszXjOY+WES
cnDINNNCKR9hvt7IWLfBFqotq4goh/tYNnGskVR8tH2hN9piI7kRwoyi8+ecrvqi
fNpv1zraJQDbNvpJp3Gde8Rys+GU4tdQFc7Qgf1HhEkfWf0yYNgnNR4NBDRUF7tH
3tsQYsr8eHVnjP/GEHEtZcMfLmhNtWAQ/sw7RldGbMR71aiXdO9icBZq+T+Bdebd
D8vsgSr7OMIp+b6nnnDNO8I1ZVRRiJULSUzseCFPhxHo2YRLESZ3fNmL/OQN99P3
XA1JIbaUtNT3Sow138ppMKeag51mxK1rj0yq18RAVDEZGbtSuXJ9pI7e/fpVMpbI
bNdqB0Tz5+jdbj5CQlFJeV2FhNYvpx2hHlaholtiAIw+1X4M9rJ4sfk39B0JlKYe
TL2ItRTXPgU91ExCtbupVfUAJQglPVIGEQpxzBMLn4MXLrinbK8WVAXLgbE08gpi
nzM17qg7kPfUwlpStGT0vhT9McYP2J3YIzwRoalyq6GiY5tH+o34j0Djg+NNgiUb
wl8oVPEP9PHY6tJ0wet+5zCgv/OeHoFXRPGf3lvLmr80/SQhZgStfcpTvPwdJTB1
TsJsN4JJBmh2xegeFxbvjYjYzcOpUVz2nrKPb5EU+dPNcWoXEqaprfLTN8g+sV+f
LY0oQkRSsg5XUqeHuCwfRpbiw//57tXIO/15GU2zOPs9dJJmGL8bOJK/YaAJ4ic5
hthB9Ed453xM65pMDFK80ofNGmKVbzQ5zRsuqDaiH0L/BJYUojDWPK7PJTxJBoVk
Pq5eyidhZU0bNVx9yPZNwJfRDk/QTWoyUs7CS4LybTCwhQd7uIMBjgcYZa0AEGY6
J07R84wAyACg88sH6H71uSwgxbRR5aqveYiDqp4lQ+VMZBOfW0n4NxJCjixj3KYb
P+y/Je6OfQIflgAReIAqB/o2BuyAYvZy0aBuFNCDif0NtroRU/UkGCMbMiNTN3Q7
ovlRv+ylKk3eRLqFnR7Ajw6Qo57V0I2ZAnhP/qZbPPIc4lRMD6uf//iBDHNHElO0
c1lxCYQPenkEu0jmZ0iS7eOpBQzEJ6rjRQ+bWVj4yF7ZgzN+bcP7Tnvm94JbO5uP
vNRqceC3oSKJT4+QVes1Cyun7+LcIC+KmAJKGd135M8CLUDFw845jJLPX7MqiUDK
NP+OXdS83XP7WzfDOZJYurCaRUc5hCqKg+4b3bNMjHyIIz9XYF0ldZQvUeATe0fG
h1yBq6k7YSaTNiadLVhl19Azy0jU1zvFRQeYOPaiIA+CH2oxnK3ORpR0VX88W+x6
HHtpK6fkl8fZz3GsInEnIZbSmwi7Nk8BxmhlwT4ywke8hA2RDhsDUiMpsdYaNB6J
rhLCtkH7rBBO8MNNgSGMNxy1scjxd+z7uYAiPKqUd08xgXNMEzgSs+Sw/K95i2+B
dmVeIr0+xQQC2rdKmaqSNkmCzZj38kdfCQdBc4p2ID0UTPhMBytsDT0fsb8GgOtE
GhHMRE9C4H+q8NPCrPXzlANcsfMmFeARnKmgzSaNP1pxr494HpVVIfZQ1Rh49s9J
iXy/EhQ+5hmp13iOmh6aBP8gdIH7m3TlQ/NY+tAu3m+eEl3TpAycSoGvt1DBSNGU
9D9jwnhv9YnYl79C43Vrckm5PNelEchSL4QZ9AE6bSNFV52IP3+Sk6Nwg2Vfr2P9
01MrzTM6GA+s16+ics5pLGS0ji4g2rL4tuSwsMu+3boc6xadMwgoOAw0USzbtJS3
Xp3nrWa9IhwQapy1rPXr+tprUL7NZsei33FoFwq/kOiKriTgXKS+Kux5fFmDjGpy
DxNPbzS80qP9sr2W9F/sPAHjBJTjmWOhAOlrEo8hoxM+l9Bu3dGqoz5b4RTr+Ohg
qGp9cxR0ITXilYfOiGcpfGr0MpmPpOir2tIoTHvJJCaL9dObUwBDrjUDXJzCHrU3
uZOHBhRQy2IyRZbWy7TVqPBimK4QTRN1ubI0dfvoFgInarfC88Qatg17HC8KErvY
Oy6gRHptiwcJ+MUWVGf9L/oFQ8NdhSqhuoVL5BtrNUbVZ7sWYA+7U5zrjwuxwzNc
9vPW9euFRJhaSRUrcJdNYR2vptrrkBgIRvsbV2itw7xu91L4wbpDc547wBsHdwtd
/VNY1CdkT/pIg4V3X4g0StAlSghaSgEVjXEHTqGSiyCapACW0qoM10jRgFea3uv7
Y6OQQQ0jy57a+Inr5fo27RdmcjLW4NbL2nZRcvQC6xaF1LQY+7Jy+YtUQ8tb+JNv
zMECDc5KdP5g80UitCXAfpArdNwiZm5fGV2EZKbkDjztCVHYKK1p34NDOiMHwGY/
nBAga0CzUx+0zasz6/fEiE3guBm68BotNOz6wMzNXNDSSXJR2oh/QqaZ5ZxsiKsj
p8xxGuc7DRCsu1wHpX7T7F7jm/xzqjIflOBkY+OnDc47LAkFcs4aQYkDVZYwiTd+
i0BD/AvPf+Kve39I61/zNNuAO5qHx8PYq8exAL2PdN2GqhR0s0OGLqhSYCxtoQVj
EFTubMlXA6EbY8FhFZ8elKbn12y540QNzcZzWjwOQxLdkfp5vwlaO+lf7Sb7ZvzH
5kN8XwWSZS0F2Oc0arv3U4BSd3oqrVBr+u9U/IjKwXPNEDoaSObkemNgQOCT0vBR
/s/I4GBv6O5017OuUW8YODh3YuLRcLNjjdu59OIBM9VUdCT6USUSGlvees8AE6v3
BSSQ17QPF3d3x+03Ve0ZFjjW2/MI3Ar97lV9wh/ytD0ao52C6HDzVyz3bncwXLgu
GTvphYR2b8bW3yURdOnvp7t8GJiUCVX7Z8DVif47ZLhbpmlxImD6s7poXJr3GLA+
tC534rMcnXLbnhD/OvJlxzPkRQX4f7+fUhh3da1TvejL3DLNhqEdyeouRao7EGJj
1yeN9+T4GFKSW3G+IwC5dOQHQK1HHUfmuFddJge/fglPOALKmabu42kH3/rpO6dc
JwbneKLU4FB+PUqlC7bNmsRzoJoQx5TGnvPowkTOYw0BrBFKre5h1QtkbNBS0sap
GsrABcB81iPvg88Fny6L0CNDp0OvNc489HvLsCEwFP3X1V4Cjqt9Ok2y8QPVtTQr
HfoCxgHDkFj/0ScjuhZztyPO16wVEXOlfgTfETqASUDUEqb/RPtiticYBed/TDIC
2m92+sajmDze0YKamaHigL/vaP6Ow4rxytQNDmgo8xX8Pw7UvDLUmJejx9hwgOu3
KNK4qLi6KvLUUjwwUnfnhcyiCJ/sOR/AUYihi8pq5O6NKp9whs88PeElCV/caVFS
P9xX5wglld7z1gtJFh8y57+2Jhd6KMbacwRpRxUbU75TT5wz3GLDBy16B8FA2X/L
Wm8ZYR29JdxfY4CQxunoUKkcImmtfSSOT23lfMv9zcvamkv5QRIitWI+48j/qoR3
uyfZ3Dadf1+wiCKPHVgN+A9MU20EoSm++gkWUPSjRaGQ8IKOTIIoWx0G/+DG0CAN
nXTaxi6KdwJk3ihYQPuXG+91ik/gkRD07Sr+RhkNnOuUbNSjb+WkDOPmJUphczT+
klo+JtOou62TX50cfLX3J9ns3Jny2f2oqtWv1lXy+MFy/Zf0khRR4hs4HSw/8hje
uXmHSBh02hPft91NqTkn5QvCYAMKWqZ9HFvbDLf4eAsNdRyICq+9WuTGVSAzb9Wr
qWNL6GCrmu8+0eQk970cQjBPRXO9Ad9VdzsSw+AOb+KJuBeLrFHZrk36cl/6X4uZ
8wiRx9FUGJykRZltLwpm4c+S+Iqd6lU51q1FPAUBtV46+UZGnZA0Um2TKdEKLmL3
Bm2m8/9IWbn0iiEyp8iKYMnCFbxtJPtcL1w9aI2XI2LLHBJszroj5Xtc3bUntJK0
s576y8OX5mpRBHO5J4hmnDFG6E964TNpr7QFNphY8KMFr4kSis0KHB1rSsSIY1RC
grl7ukKmnYb0Cpdk4uehGUbvia2I6xfswuTmm69RbT6WVVchRHKKD5eTedoTOkWR
DpSuPGDJP/LQGoN4wYhrIDNQoetXAJeneV5VZiWlEhiKyorlu+H1oXpa+0MOhnSu
9n+yKCCR+i2Tj/GFY+K0pLOnPEfweXMydD/a1ARY+9j/xxrYUCWxLuBjBkd39kJN
geZGdmv/ZhPy79XtCOYpwUUexVRNTIAeO2JUftncIWggkpFEsMLenf7KgWZsywJ4
jFRH+sjndsmAXqG6OFJKgYQKrEQcX2YdHIn7FlJ4fNyZYGbxMmjVn9KqQVXQaB2c
l7ExTzT731uhwb1kGCSc30b0L2wTWmsrhHvdi1VssAf8x0klaW1cfOA+fSl0tbTV
aoUlBP/vy9whHOWtbHFuys5azXJAmCct1y90snBJgDdv8xMOPpZFpVRJHbv2dciD
lQ6N3etUdEO9MmKQriWEIUbtdgihafPqADShl+kc6tUZdkuCHXiWVHApMd5HLJIR
7IVNRnwXiZIEOKq1v3uHa9JDi92bKHMv1krMsNGy7tcTLERKiBjVWf6SV25d64uM
bNr3MqvmJ1XtR6/ZhyoEoP1mk0i6v0OdyympXKIfTgMn+Sm3qosY5s2cpeVLA3by
ARsbUdtm0S/ELOmCNV2zYgNafOvgeFLs9z571cI4jucTszMi8/tOI1w3VVHsnZYX
xZMQqfnft6l9008rWy/ZK4kG8ROisR1hpgBPV5ZJ2q9ZaZPX8AbBrXSovVgHR44u
8vMxHLExJvR/tNzRjyyZ6e4HpUnB15Pn3+XXDQOrGlNN8KtV7LD+On1hxyp4isMq
IoUhwF9e2ytLAVYo8Uk8xlkWyRBXRNgB0COxWlfWEIYpht96Vk0kgjflefMVf8yo
q/rFNpnc9qbctYcaHzzKR9WH+EABov2Nh6mbDP5k9XWEqGV0gqx6NcB1gzNyPFjD
mAs9/pXC0g1+88mdpiImLHKc5aCnGFdOQkiHFKNePrAm8FkpgyKoDn8+2cYN6mUZ
xyznmFkT2XuhknHWEAQz+7MeCpgx4TSRMWUbS+Zx/CMK4hmuNyjBsduQYxwKLLJz
qLLQuc914q8NcYfp3Ai4oRXO7j5het7RvvvoGUpkjQXOU8LvBzD1+XSK2ToTcs5V
mdxbKH02MmXe1yqnjS7Rm/iLyOxRoPEWwr1IOCs8rmZ/1WgpgJdasuY8CsdTvTql
pskRhUOdP/S8lBb76rgeZub2bJNmGrb52ASaotGoRykVevzeNj4Gioqoc6FNQiG5
lKUhMggrB2H5a2bCGkVSDyjoPMSKtaOhsMA5bRCHDpgf+98R9z7bvVsOeVVAk5zV
k32H2osWAendoNxoRmtzqQ6diVi6Z8NTq3BGbv5EUDsL2UxMFDYtuHcoo0/WeN6B
CJtf8hrk0n0AKvRkoHI3H2bzjyfmlxCxP9i3TL71WOCp3/+9VtVuBaT0/i+7q6W9
5RbotIwQhrIytQ2ZD4/dB5xPlMt9RS9r4NlqW4TY1IXB114S8m0mdgM2Rw/hIpAx
8GzovHJgzL/tA/RWyqx+rgIVRPbEO8Q+Q2EHE8zLdmWsAHOTbfxaJBKc4xBbDV0J
01lGCRoXXUvmGYH5FQCA3phf87QrEfaWcv8zzKXrDPng4ullY7q50SsAsP5hD0Kb
CYGHzGpeexCG4I0NlNXXL8LyGlyk9doGxaidzjoKXGnN0L1TIZKasG1gxKxX4wuS
dGjxBl3nfAPYZdfTJw3bKE4bdjKk6SuPlyV4a4yPU7/lqWavOW2FdavIoE1oq8qb
myjEreZIRG11OEKUL77vY2VbUr613atyzKssL3mHqY5uP69ulo7Ao2HcKG6+wEOM
5LPMPuq4ckoAamMss31f49Wd3eIr8gvmYwYHnUfpkapObYChyBKh6RsOTxBf05Eu
5B91EzoKwMruQLHa1oKtbjqoJnT0lnGhfWY2YAEA2Ze7IZ3cBVH3khKKQbZjSh8w
rxyCYS1DAAsikfFxMlhyt3Mk/21gZ9R+S56SNO1Ev72EgiYNjimt5rU5i+KrX1YJ
KfIoUiskRXJzrQI9QMwg/swg+I0tQDZB1gnXO2EUKlI4Y/0YUzidkOvbatS1V0x6
vrihZYymoL0VfjqtmxSET71tlkJ43cxqpM1G9pBDSr/5w594Ly5iB9NYiBfFfzeQ
0oBDUVfXIeybj21MurdDVI8rnOIVL9sFNZpu/99SdCbm8/qnWAzWX4JNVcVq55qT
S78ApvAGgQfQvkFlXPt9a7aT/1m1rFKvRZk4wsFo5aHZnYj/qGcz/QlZ/DdAiIJj
YJrT0nTkBE/AZNJmMfw6/Ge/SqwWliVYEoxvj6klQvyIK2UE/pfpb2D7wAsVjt/w
Q8TiubwxA9vqnIDMwoY0mnwDFGdmPUgOe3TXvuvyvtIJsb2G3EeWw0AdtXGH6QWB
xR7AfiQARFSlqN8KZxrGkcVKr00qbLSaP3jM3AF1UcLKRP7BsZO8wMABYzPwbVyz
lZHW1jriyO4Y67cLS9iuFPX8v28NzvDegeWtJ+FqsLWsnuaje+kguj4bWqAkS2Oi
jwUp6c2+ym6Ov//TIMeBUlWsvcoPWGrTR9QJDzCjr68v+vgGGw1M5JHUtcnlyHvy
v39rtbAebHyDfpF67dK1F+GLG2FdZ/sUr6tXXYXZK1tQwyuUJp1RmHFhGjXWlG2+
uQORwi8u66DxuNnOUbs+d0Ejj4Vps07lveGokO38R1ctLgg7B88vlrT06HNli/xJ
qn7CiISeao4UJ25YwiMhzJ3CHp4cwvQZdSF0aldPsaZmLi4VDwrv0IDfYqln+mZo
lrq36VkuQYeUtaXXAwmgrFicc/eW2b0nDd+LqC0Z8EUbeh/6mRYT7zya5fTDgDqY
XnczSVsM8cDS1/8TIxmiB7TJK2T/QQFRHUIykoiiuetTUnmaWqNy6KaQS4vrsAlK
Zu7zHgvvCb+oif963zVDhuCgHKigNWmRRcWMlwPnz2lfWeVSoxXsukozBTQKUYIy
liiSwUzxLusP5lVD7ty1LMSkofA6/eCKVw2pOnIh0PsnG+AcaOkynchRXZMCOBVX
cgrFvvQalotxl3M+Lnz3RBT2sKraGoj7hrhs/PDvW713SXWwBAB+UuO27FpMtvS7
qLDyJHWNBQVSbZ+6z0NMIzYYMcCx7EB4Dgptmup8Eddb/qOIGievfUCKCbvt0J1N
xD0AJ3eOClV5xcOZGhkif6iiOelNBEGmaWDC+kLwddRaHD+86jV9unkz4y2kDAH8
de1t3NRQo81C1j5HGZPdghFWovsjS9W7Fusi7JE+5xIYugHwtLpTAdpksoLU2C4T
o6TvGiyIMOSv8+z7T0JSAmlrLckYdSFLDrL5s24mZ8GQYq+PeOgtb0SANbFOgGIA
VI2GB/2PQKnWll60PKiBITROtKK0DkwlR7L9MkU1zIsvYvkE3slN2axHDVbcp0TY
ulWMKagFL800eLua+1oMVpKUk46JkW71i76gqhCYCle0iYqUDa41bsYLH7CLsLrQ
WP3Zic5O9PuRkcxfTRdgYtGpNoewC7KfJ4ALZRq3ElVb3QPTG8kWmsvqUsnNji/g
lbiU9ow/ZVgqILHXIjCmJFTmGQdbSc7DB6m6fBIHLjlI7RyS96u6IykYorynOaxn
8F5WQjwchJLxhOJrmGd625+RpPd/WcXFhIoDgFUvb4tQSvJiEeKee9mo4rGStiZQ
38JG6ccz/ujxk183wILVSchCI5DfCy/WXC/LKpUYQOwm4Zlf485fpv4W8huxhqsA
fkGS0JUo6BWa2513m2CHMbLCTmLq5rHLTKVYd1s8kPR0OGXrnM17IOz/TNb0JOve
RkvvkQAUvIGLBOiwEy25CMPLfpRDIzBYeXHFzT84ZfCxI4EZh4SKl1Hgs8KZ5iI6
fvac7ZAtlpgydmsmKktFZKaRnASuZ5cMMbMEePlEdQpFpGTUX58MS2Ta9PyLR3Og
Yijp8+HPjDxT2mw8/9XfnbS7dwFE3ZcTyUDPvx4bl0O8xVZ0t1IJQ4oUH9qqQxrM
5GUlxtVNal10BMZEtdmT1GXf00tTjW/Ndr3gN0xzs+9h+oYn0NrVwMM2XXj/xQ1j
J3+SZY0xHQZAStXOZez4kZlj6HEgDdm1jP5xso8OVvWsT7+dzBv2LA1cojbkUSF1
AG5N8F6NJItcaJEKfuBYT2D6I96+jgH52TgEUMDDb54wlw3GjgDu8P6sla12Htvb
A3St/nShiyNSu/tg62lcHDYuIOVU17WkHoKP5qKryt9NeeEd22eQGaTaPQPSyYg0
t6MwdyZhC5FPa0vgDxv5WXVcr1/N7xJYTe+JmXk6gQuKgFMwi+Df72T3QTdl8RCQ
xdanO+Ku7miTcf4F9VAtj8yrRiwKi6X5sy1WovuxEzY6yXk4RNW30t1srEBgQu9q
3GcxB+WhcdvOwFfUf8EhraoqqA8vqkZYuMmkJCS6G3MQe+GIFRw4u5KMMy9lj4Kn
CrFpgBXADEQVh6xa+fxhTFlUYqyYLdUIiUal/uEmadrTpqnI0irC8YnQ6knXwiF1
UrvFCUaqEktXpCtW3pL+EnWd8QjOfBMPry2M57k6iJzQ8DOh3MmF6DXAQFliX4Io
p6v4gaSdiJP+v0IY2RG4S4euGHN1w207ZtZqwAVCV4bx9uejzfBAe5E5n/8YF9Es
cm9jVRgHbnXr0wOBUOjcVp6nkymVOvVLvu5z9GaETmuQezrSh8Kt8+Jd18kURJgN
BevMP7+blAqtvtwdc8fLc8oNysNM2NiC7eUAJD5lfnmU7NcfNgNuIPkd1l9U9aHv
+KOLKyiAnU7Qc4Fq2ucW7p5vgHuM74cbnjcJzi1j+FEA8UkrvjeVArIur1cAVuQk
PuPA3sFBV2g3iFWs7Fdb4Y33GYEe3oWvyaHlXFy/PhIOfUXkWFKHv0S2sZBP1WGZ
pYYdAJOA8wSCiKeQNScmUvCIp830+sacWX8xS5h94Qs/rokOGn2gfvKSiwsdizL4
J2tTlXwDj3bd3Fg7eJMYKDkGWghZe4Y5exKMqqxp0EoEi71O0vi2Uokbgd2g8yy+
qrIZVAUE+yMQCT3IYMW6G55VG6trs9i5rO0oJoY7zFq/C2rHBreo35z38RfU25ml
1KG9qa8IG2/w3V/yH2DjIajr9TCrkF9OjQnZJ78KwqKWt6S3jyrzMdtHcPWvM3yV
IwSNNoNd+ZxqaxN4xVpK5skN+XCFF4LhxFlmYTHTijYZKd2KDV+31gtG8EGq1mS3
cyUJALa4+vhHc+DaEFcveP74xr5wtwPnMyx0G5oqosO7cqt1OdtyNf9zxBjoekdZ
gu8QtBK2IGtNGGqwQheAoefokOhSSjlxnQP4vJkrBaK6rx/i77gwekS6cq2a4Fep
Wsl6zTiXxte4Mv9dfySYzULCYTePY+nmve6QidMtuNQ56sW8iGonbbo60i86ZJ/f
MrudCTxn2cNG1/3z42au+3jVMK18FyLHwnFRSkETJtHub1tFf1s55ghbynRfezZu
/5yXwvj76ntWyKIsyAWqQfJ1rqPNKNmmgWxvFUnXhfTkZ4mRaxCneusJgpeMZjmY
YSW+hSVI9z4l0JU+le+7mOTIm37q8uep9pVz3Z5uKbsXWFneGJe1G+BJSa/wVvgO
P1H4bYVRjostyrEk8toX3XNYABnhbz3YwhUHE2Wv4wJ13vRIhMYKGyOZp8ShuVzL
yDN/gTsynHHuWCPBleBAm8mL91ig4KQjjEeBDIQDrn/IgIA6+fZC2BBLx+58X5Rn
Zi90qrEQKFzlBqtU20hdLXP86OGupFRERAYPooPOiBhtLH7ZXqvZ/OtYtB5H86vc
nekZxTlauBrI0y3zSslYsLfhF0DZoGsAJJvsdvTxc+e+rbQPbs6AlcnuHmxjRk7Q
FaQoM68TVy9Ph+LDBladNf9V5Ed+gXEY/V1Xn/OnMvT92WsQl5cnvpNdENWqSdb0
wZN2jr0GJ2NxfGwjbDkNdujQN3Fr1LnmaKja+Zo5/943oG5jIxRthz7h6VO51pfu
JNw1AEFN37yyILL2UvhZ8cujEhQZvHAI/x+0CbMcevFxvTmvW4JgOJIESCVTnq0K
KvtpGI6fC+dsUp/G1zCpyGzc+8vf1MsfdsXdGfwlCNloJ5sxGMdz9F4l2j1wtBx4
Mnh0/WYY7UWpbNYod2LqgKjVozd40rbI/ZTZaU6YJn+x/GoYYl5FUTSLJsOCNYmC
GbdoBoojn5r6OgAdrEkTHz+ke8YxJcnTQvAFvLrnNFfstw6imvh4EplEuu0UPpLJ
5CFXqxqSXlFUVWYrRMFAAIYjLi3HBIy6e0nxwRda644zeQKZ8hOJPQi6UgCSqD/v
jDSwtkcWYuBLJDA0z4FU7j/A6NHvgK0OQbZTbGBuTwfL+2rLmm1t3rayKvAJ4WHn
iVp4o5PTBtH0KoHBc//8N9il+eG6fhSViI3/JLQV+CmnGywy91lYkj0jaMJuLRrN
z9rnoEXtHMcwxfZbpYK8b+hGFU78ApEe5QUTbOoFz/MivnDk0jP/LfI1EuzIeVzI
UICm6JXIM+TnVN2IJpYWkZcjMh9GEp1r5AKYY2o2ZTAjmDS6OKCWUWVJStxWNaNY
VSEyVDm2YJ8Tmnr6lF2NyJPEVV4IYGZivdAPJcIf9eQWuTgqeZHKMOVkksECIXh9
Y4MClKkj/gLclPv790EPVUuE6gN8ogzP6do/6J1xvdBBjXKct+2lJLcwth86vhp2
DgxQwQA621b2MlhRTElH4OuNxF7vPNexMxYoyPdH/tvjurwwHRX7lKyGQRGXYp6l
uSanYQDrl5z1Ugn4bykGcL6Y1cofQhSnMReWxVhHnQD0v7rYGIDjgn0GJI8anDf8
uVNZrDg8j47mgH09YGzbIAtZSdfyv3liK7HorgQ1yrqYvP4rxJi4gdH9TnRql+kt
dQOVstNVUoc6BGr18fsBpJsxdqGNCBo9Q9mRiZIn955kolcmNpemRYTTwL/nWtJ9
aWlDylU4M6LSYS5bWARf6iPaZcldC5jbOlmx02UzQz35ST5TDm6vi7GoQLfQ+0kF
BggXeQB6OvSLpviPI7tdyasOEp6QxHSEkbib9SSCp/9Mw3/qKLD7eY9WWXzC60S4
FbP36Ioo0bTX9kvW15U02tmN9tl42znJ0Pa+6ZsTfbl8V9wKACOEF2pGI2lSHyRa
mFga4HRs04kkhjtoGXQFceEh2FO7gfCsuUfemEbuRladp2wSwi/ISPOZiws/ejwZ
isnOPePScNXGl810/JXIPUvXYQSPZW6xB7nqLrYIvlLAb2ddy7VKDm31JMeMhKUJ
Brhz2rcVwi/bdfCtmWInUb/gNpA+NBgpP300+pbOYmqqi2YBMgqbX/gGZBFnrjb+
t3HwmmJUhFPmiTvZNE0FSd9Jqaw6uVyRhCAo8GyfK5h+NnmT/qyvsNDjTZjNIcbq
GevNKY09yq2P9tyAF2zXH/Xc4xaAaXAFeVyJgaIBWYRwe8v/Lk4Uch+BfQWtT+eV
cGwFWzhEOBTDfe/ZGFd8+Ek1wQslRDGQZjsxckAwyi3orLPYbO8yJ7uQxzcAYCVl
rqezHaTdVxzqidAiBK+K638/7VWkVXIvZh9TdNwnIiNMAbWvJHylZq3YzE5IkwbI
5VKoOAaSTg859SXqBCHdcrtWIzxAp5SjNzXsWuXFuuibqzjm8+2Qyduppdn+MZmE
vuXpJsZ7Xj3CUE7GdDnVZ3hLYqmXJxSI0cQ3e38zN079PuGN0DuagzstlPKaAV/K
NOBH+CdX+F3j15cX5avPYRIYX8ieSu5HjP2l5Zk8g+1xyBd83nbMPk4QW61jt8z5
/PadpM7u4BK8q/2tYAHRJjZ7dk+gT+VK8sa5xM98FbchIUb+48gwOF41ZtQiZ7RY
Ktc9+kfBVXNUY3iVLoAO/+/oHs7seoLKlXsPvHox6FJgio6Riy4SaysDExtICES2
lRjomT6+h97CR4O2cWlnnMr19peG8I8pr7IO3+WEWSBbMszMTgJRqjPQ38QaTZLh
58Vumx9qcVhCZRyEeYoo37qWcJUGItpZLWMbv9PRtceqo1MvYlzLGvU6/jFoL0Qi
EG4jpaLMvH3ytLTl9gLlMtMu754ek3cFK6MGOG1XXMxi5wK8wc1ciOFbUkQjV3X+
O+a45WykExCDu5xzpkpiGOVZDciVz/XeW3ynmgUsQoYxUlvYDRNnSZwcCQ6vGX/s
IXPG1hiLwXJuN4s1J6dZAtQyk6pOTqMfh28YCpRE6EuDCnveFe6O8PQyxDK1w+d5
9toQ9bkKtAf81KpDN2ixxqUjBXSVZ7xbUaVtiShJmzhdkG2Ome/b0UTZSGnFv97Y
rT08NCdtGmzBLtC5IeXXwogXVitAY36BwDY35aDkVvh1V9AKcIy4FfmaLy7z8+nY
PNJ8zNxv21zPh4ASmhthuuuzHxpWQoJRllPkw6gL7ITMES4EolDQQAiGzo5zNSRk
VjEKK0ksHdBD9OupjPRI1S9kwUZLSD8iqMfg4cxWgFc2+XgxzOJqBDnqV4E/67Me
t1rFj4JcZW+y4I2/YBMAeStHwCLNs9MtxVJDtvccAXmtfmesmFaOCNEGnEh7xwEk
WFOLBrEEQiKjd5C7uey/vZ43jPEQp9FIVFDkNvAAp0xlbKnBs7wxDlFtSdDnPnAY
T+tYOhQql1VNozT3XCS4mNa2Yj4kAl46kM/XYa45r/Ef7AKjhMMgULZw6IJvHmv6
XENjKxW3ycyTZi3vp8vI4PAQaWc4JpQ273dPtMwEOlRfGo7GUoYQeq5zIMIrX2AR
10aYUL6HUt+lNgC3KQPhGzquz2zeWm3j+RfzpjAFk7vqEgvdAPjiSUfPhgyTQU/e
wUAk2cVd2Fvwqj+NDSOAwI3xSHWOWHw7JM96Creeqa2rLWoE/CalcRT8Iyo+/zik
2pTS4ieEKSR1JV3P2BcKJDBbpri7Z7bXGlVIbIQx1zws7pczkHBN38d1+48cyG+S
QFUBgcIB4SrET8qcQZot5JLPe4Jq7vtckQN+efw3edB8fh8do4JIql4HyvsTY/MJ
bgb+gtTFIzTqgKiwEVa0MszOoM/AL5ZhunWOdvPeXn6DtJ1rEF11MSPiQSQssujB
oW7KM0Bl5Oi93xMNc9OW/8wjfKIsSR7NcnTGedy9eRePBMdcqqxtieoVJCpnLJpW
TVELBxDorJDJqqkDKGhjNxNnxgCH0JcYz48SggtGbC2GJFxcMcnOoKKChSjuGKss
mFU4Bk20ex+sG/K7L375V3cL7bARzs8MwExXlfWmZB7hq4Z9OCK81TSelveVwVTT
Q6dA73gbbx53U4oFQAFDI+8Url9j8HihOZ4XeJRrNV1kCQyxx6D08F8b0xzr8ZUE
RVOlALxCnTrXBnSSUgb+PaRshf5FRKJGoRkD+nQObUlI+404gqfDpGMtsFX0j7RB
1OFp+hXRuZKf0QcWI2FoYYWu39Oiwa/rLnQVpq7po8dO19llZuvFr2k46xkO4TVV
YogxkQozOnkzf6oyBn/RW0QNSkALljmBFyLWhH7tE0G+LgfG66rVy8g6AhqK12B1
25cPnZRmujypdmT/rqG/Y/UDYFdP7QQfwmRlf3a3hwsiRyi8dRr4MeHfI7nYfmBy
WDeDYAFLvegd7SKop2hwT0GFoV29+dYW/gh+xUHc3Ga/lIplENAnSJaraFXkVUaM
FX8WAaLrb5CezWrvEmaeKV3nbrQOu9fnNGCrTYHbYWodn1y0pxF+1EixRn78JsW0
CeZc8vanCw3XVX0nZiBoQmREgplaVEeBHIfX5eW241mXk+9eM1LbRcUzb7kObsfj
AjcCsb3Pdl4V1+E6XfFGxianIl54iIBQruuwEmxI9z6RXGooH/fNIWKL00H+1bhC
f4Yt9FqYibccX4K2RNHTnJ1p20bhGT/D9SGFu3EvWkNIWKx0zsb7xOtOnlDuqrcd
4bWIaqeBx3fhTEmvMH/HZ3KPzsecVJiYpEUH6Ua7EVHNNkukguHdOLj5sIJHsIP7
v0dCBYlWvx4BKjE84xyqZGpk8hHGuW8J4PoVdaqCLp+z143mJwgsnCjaQy9Epjvh
B3pcDhNCa0G8DFyzjvPwAcKP7ntU8YMPCBCbk6b3dEDJ0Vq18l6SBhuAqRi/NhG0
dSXCMacqrzoDR0CMKTIpj5vHB2v1O2MRVWFxvpyCA9bHzkenzeOCsPyQRy0uIltH
iVbDPs9VSXYB33tywKjwaXHYU1Uqutel/IT4q3zRX2yctonVDXgofHwR7eHxE8os
+6kdg8ZT6ragof4eCV/TZZKBPlr/7ejA3oKGz7WZEupR/HQ+fu+M5Ya0bs63wdqy
TFHDehGq+DXVz2uRqnJJ11qUqfit/jh4zAWOf0eD+jIlloMTRItKPC4wnTJoObsD
V9Pa7vL1ZghkGtX9bxF7wptvDdpIlLVa6Jpd9cGllpBW7WUjKosB29PybJp5YuCJ
wsTmwzoAf/CcSFvMLbGLcSHg57EFRxfECsd9olvNeeqR0XLaQm0qCSIzcaz2BUkH
CglC1FdPk944c70magrMvEt77ZRUh5AKo2uf2/yTdPaGkLrqkA8bcTCQ1c8tafuZ
9BwsjNxcrcMpBPLQwAzWEBwPQsX6SNE7ocP3Tg+ogcfjVAatBGN2Xppa12d7z4EX
sWiXb5jcd+9PLiU1juYdk65wZexf6Y9WSBzsedCu3cMNRVZEU2hENur0FQ2nArbn
QeTQELkhZrdjfhtE6f8aE3R5wmrf7B0n8HnyC/bOLZ/Ud1NUUfxShNQidN/KI3Zy
bGgVl/jag6lae/JD9XY5xM3cLF+UaBtc2Wo+zWL7FcNdqM4ozfg+oMPF02dU9OHF
8Y2A/MCOTGvmA2GETAMSA9931a/DOHQFM/Q8LEk6xAPW+VIB54/+pKT43Z/80Bga
ra9/UNXuss+vfaUyO49dykRnD9QB4IAaOi/BW+tpwwQOp4R5zAYeoVSDAeH9zVXN
LviDZswUWGsYB0424K6LLFQ7Ob+mHuKLz0zoeFaNWke+LpJ/MVjRxSGcnK3wLlLY
GforlJe3k1n/F+bulHtla6iC6kwOEM7oKOySWvZAhO8kSUMzarJN8nXLiZMej4f7
T6Mg0X2/icZEK3HoXjaeJQvz5QwSLzbRfr1/C/ctnu2T9UPjk8bwRaI0VynpY9v5
rwAsQrkpdIjbcv3MpxUO4lfRJOch7/BwVmlBeoMrfxesDXvBv6F/sY46eut8t4Xn
QC6xT7oNuuC4aD6osYb9iMj1eFEkf0cABNEGCSxNC0Bit8CeAiMMTHkLusAexq1T
53n5vwutW6RxV3oDUzVbZZxh0+42us3Vtho4SlQQlWAONWA0S2t4eKA3EmcGnqRz
GpTU2jhUH/T4/BlgYgWph+1IWQAmhSUUiYCatwqZUXFhHfFLDG3rXNwkiKeVr2II
zww7JeV9H5+xmRUm5EKu6NQwXo40rXqFPdbvIFb3u6i6vLpNg5BHwIcTKxFe9ySR
tJld+iDcKkPRPpWOdMx3Gdd5DETZPn0kQijvUcKxW4/LGY5XlKOCTF61myZ4nSu6
P65ifC3krCjT9H8vTYlmuOclY8WCK75nhRt9+SGAAS8PExJ0TT7Z0/iilaI0cy6a
NhueNYQ0/2rqNl/7e9PAhnv9UX2BJzqxZE751VDErk7oa9YvRQ7ZZTHbqolAVV40
RIGapCi7uBDko+bQgEshq+mQj5Gz8aNG5sEbsbbv7UlVUrcMJ5WWSHYZNzE1dUf6
DIeOai8sYIoQORtJptVyhOL9cwZkhk22GFhKQiFUybUPqBck0kkkubF7osPbYQCl
LcoH0i7Q4s2e0YtNFFJc9PgkvdrbcfUdxveuxDvzL5XtSHrTMMds1xl1iCYct8Pn
y113d2e+xw44qKijfBhyRHkZOOsfmj6Lw71bE6fQGJdXGK1spXebJa8pS0gmOL+p
nuEkqNtJe2ImkcyoaaiD2PiToi+PqtCRj4sWYQai8J0n4vSlzU9El+UsqskaNXH0
1t5qQoBHwq1EcL9DLsSHDsv2ZZPXljXnkgiNWJGC6QURYWgLo6q8Nx5p4btRSreT
7q1KERcLAA4rJluqvymc/4h6XwYfXa6mYldepBtfHq+RYr8HvopVLyqzcCDf7bug
Tn5KfypdnSRlIe/MwiNpgsNCmLQMmGMRt4n7THD2Lo25/MdwtOAlTB7Wqv4wfANj
wupfExffVq61a5Jl4/XeyWmfBrvyoAovM7MLfpr79M2Epa/62pnRPl2GmZlYgr9c
jSJcEvagxZEAipms0OXhGVHxSs5Licrkj2NXvLG3K/DniHSaB7x1RfxTTTFVUH5z
qsIXyJO1DyfEBXtUcjPbq5FzNunXV9clmpHh4eyUn4JkkOhHfpBnY3IhlReSB2Uf
KqVqs2NA2YDYQ1BB/Spua3rCkt6Cuum57DoIL2Yht2/ff+Ffo85oGKPUFymqfcDg
k9OCMBnfaJ/6UWMR7nPr0RyhmLsEmRYsmOjW4wV9UQSQzEf4L0y7YMehdVCoN83/
K6d2Scb1hsf1WsZ3FAtsXy0ef1N4uYqLZZlbIEolKK7B09ncrMxYlolJ6IqIZWLF
kSHGMkLiiwFBQnrL4gALIP2S7JPxyP7ojYjQScyaf00jqTAk+N5GDIUN3bPlByBF
k6OwYYMjqQu+afvkSLaLfuw8CEzhCZCT67cow1hqiL1vdG2MdkLMf8RBzzEAyugQ
l0PkOLxMXftmWFIhiJCt6AyoD8r0yS2RyUThk2AOJBOoBGNHzE3D6zRdpNN7B5FQ
HtUdKF4IUny6xMFe6NKBFhCJF2LEaS+MkVfGGZP4ahYdlzhx1/ELhNsOiFz1nyy9
tTgGSqV/EOIYaVFlzelPGbvO4Fz7qQGnJcNEhF4/xDwJGgT0MgLJB5kqt1rbf6ys
56pYM9HRgmJY+KsPisr7BmpTucMGIcm2MBauGWiNElSfENCxCAfwPaaq0hGMr25U
QdHagm2QgL9/qZoK+fRWa1JZbCxKmyXWLTiXLUU3WLqL9ZF3Jjr1EjgfeD8zfGh9
vTHN0KFeBPeDDFn2qUOJhEAhgV0nHxTrYoOoekg+tizmXWC7gLep2PackSX/4m6A
81sQZ19d4lsb4DsfExjZaB1O4ImWedrJeb9IoC9Y0Y0smQ2mQNUx2LtwDDtrHX/j
VUXvVRJPApkUjgEmo4p4/cPKsX2spJDhYizlh1IFUvJRu0Sr4d/U59rn3htakeO2
rsdpwATx4Qu+8gOhO35SfG5M29A2bvdvD4v/g1twAatVgZzemABBKrjQ3xTLQtDT
OHBJCOotNl3y5dzQ8CtkLEWKznym+E0mHBaLRnp6FOzwagi2ut+RGm/VOfioj/ge
8wdIfBO6ou8lCIyoSE50H7+TvZEyKM3c1m5yzPi1gKQpiQZ/uqGWB1thdyVBnHLB
pa70FgWWce+pwuGAg4Z9lkzQfP4Cdyk3bJ9KZB9iJ65ojpAndPQ7DsmCVdG30G1t
E9wmELOrbzt1wNCCHwA1ui17J/WUi4OkmLFAe8+if/nhTFC23+xerMUAv4QCsynj
v6Jhmfb9MM0pivyCkEVzVBHlvisXOR/rcopJVdQK5XQmXRozBb1/aJLV4kcwVa7M
ZZheSZih9R2finZupLvaAonJVFIR8NqXAJAFu5OdrNxF3UzscTEaa3rpcAsF5xFh
7UxR8j5XGCGcvSxU8bfUo3S7KuUqRdb3oaveYFPzWrqjs2jEh/liM68dTUR+Z+mL
+aLxMgKvdOmpnYBPeuEVfliXWk3FQoI3WnBJ3NBXG+6tLyzTzvKJoSWSkW1oAPnX
e5bzdaXbAmOgPSPdigtH805BdAT/wXFkZo1egoR4wlWVjk0S0JxBYejUhOROJT4f
uHYOwJ9VGQdvf3arU0e2Yw56kMUt15tVeGEEfd55nCeluHaIIftYwq9pDcsEocZP
0zSmkdOde4LfIr1VlODuyltsNTMUxGj+Z0vIxN3HGFRGGFZgfJieLxwTMYkZ/HT/
VELuUTXegnYc8//BI0c3TreBNEB35Q5cNwMhaVC1XIZsxcl5b9t3HIFH+2mUfMTS
PEN96NCLpHB/oiWjhU2IE/cCtHUnXMpua+zNsQsX68kSbUri8mS8frBTr0MVS497
iZzGqM9c5n/5B5Aex3tFfJdfS4f0yqqKWJAqRVSCrqHicwb87JaRYP8nY1hUWjNv
JDO0eFO9Upx45N8EeYRCcbf/1qH27UBajj6EjGAdF5Ohz2kDJRaj+bbDHm79MXg5
Ygp+myj2jkTHCQA69kDV/jO4cd+S7D/GrSNutQm0AUaJMOolNDyVgtz3X51QR3t7
VzB97eSLveJ+YnUKkMpZM2TLV5+ijWkcEtGmzrp++ny3ZcgOkhxlugaqBHIbmgzJ
nC+WWgUTN5hHu0DGsujT3g2ihzZKg11gaGkabsOXYa4ojXHndJEShyEtSYnEtvnc
b1IIv2uwFMGSp6t0Ub5/5atANkUqiS5dtdxW2MmGLaUolVnrdcFS5NkrKow51pW9
iG3DZy9QQMOX7wfRGJdgBJ3T3YPhWceTe9X4GXsVAEvAgq5xPRy45jUyfljBsG3+
yBDUnztRmc7QSOLS5HBV/KAdp8beTpxhDM/vtHhbQxYl9g0d2dVKPyH8Mpp/N2iq
1uxULzta3ExD2CHjT2LCDpV+UGXjkAtGXVfvZoTBDAj6wUpS2TGkrq3Z8CklUibw
D/41J2feV4rg8tpnENFtJ3lODry9LojnuQWAI8/oOhioBrIljOSeHmamBrocIaYu
namcoqlUrHpdpIH/Vns5N1Pj8vRnCr63UBuYaPLlprUlp35/DBQL5uzoTCIMNbmX
CnbgEI/O8LuG4MZqJmO6Vo/+aLYQQkGtzlzpX3u3/cLQ3oOBX4Z1cDUzVGvGvZiI
r9TLJP005MW+MZ/9QLquStbEhICBGuYLHoxkPtgaaj8fD0K3vDvxwhjCfugQTySb
6yIqPg2z9kRjqRwqFukfWijzqBrFv9Fi12aYOe0/8+gDlp9EHq4eO8TA3PVgV2m2
BfiupK+MuOogu7qdYVAXoaCcj2pyP+jP3JWNWq+Zs5f6EBTbWnv8BDPvtRlUVP0R
ekwyn3aV02ppLx8VuyrVjlCurSeHidGdzOq08LNMuuYioVc8xcs4X9EgV7j91zc5
u530sP7ALnxnwa27f8Rfd1Ja7sph6n3KBAO0MpkGuGBH1UG0nO8pDngU6lU1Q8uy
kv5+cvKzOe7qn60BZXw/NLPqQd75fzkoUvQ26fayuB4ciqw8JzKj7A8nuPE1Gmxz
fVM1vM2xthw9Y8TwUVrqRdfjAJRtT2IbC3sMYA9OEaEgwEkAtlgVAvo/hPfKbR+d
RmjbUehejNqObIcJFZBw08JJZ2epdN8WR5UCoRm6dZtmzYdySQIrXZ5qGQB07SRW
ivAtJEB/wxa91WfeTSZ89Tpy/aLdXL8Q26/5sgqsjDdFbTja4WIBWHqQY8gFwsH8
duc6NhYJwUiuqliUzv6TwMbj8a35xEX9oZ6CRlsDGX7epE/6vcQTPIQ4UbKYDzRi
tbKmjU4WM7HQqmdMm4EtWYQQ8IRIT9i/+pt9h6A0bcx9U83ZkL5kgLDHNgI52n5s
cbwQXRLxVbTbM6mTXQN+jFP+UgiqMVki20aIL/kGtrSRNP5UFSMZppZu0TK1Jg3u
gkFG4EllpXLe3UPev4P2UAaQBlsWmwjpEkj/LrQZPSy2U7rPM0nig8s8WMFhy8eG
5mtlvkXj3A7dyMB0RkvxkYJV4yKE62H19QwnFjGiKjRGOyYGAItjq6by0MMAZ+oH
iQsRD3tRo5vHB2el4chK5qOse6ALA0yayC7PuqlbNhWXeGMmVo/8PE1RReS5cL3r
+lzV9yA0r+vLLCjhVBFM2lFUtNGHTWwmsyEclNT4ejZ26+PoQSfgn+hTzh5HYCgf
z9N2WqCVlxl2B+ZNUmRAnqDd3BpsBqxDkuzEMq0FzhTDvq+LfbQoJZrDWPio2ir/
9kNMqq9c+uwueflHnifCOfAOW55wg0c95jNK80SdraTACaoxqPd7JjFSPVzuxUGH
CQnlYazdpDauDcPjLCtUykF0+KjXmOckq3f1Tn94qNj+02BExB6DLomIZMXn0uY8
AqzzBXXUO4hnAK3M5ejEnOgZgDD4iNQUEcVowcXqx2Q6oeq90TN4e9/eirOLkrsr
NeCRDbhW7NgFC+N1Gitc4zAV9eWus1FRagHtB7Axaz4L1qt0PiGXzILSsIUgJ6Tv
EA7JA6RpBgnMKzNCTEybtgeLmTtBbPB1gy2ZsCDjn9o+jx2tB3vSkhW16NRaIwvQ
eoP9UeGojjXByw/wcKi+GCBhGYPWG5SZeMW9Dwe6czp4ddpm82v4NYZWXU34lO11
LtvB/8mnxzg2OBWAJIA2mWkQeRnjFue5y63SByiCVFbSXUKd9NRtWS8k2Rmc++Kr
GlCCPmuRZliZAtkW/uJbXiAqH4/csE4a15i60P02Q4wQRJ4T9HpbIT13sELniIOv
du+C9rA6OsHzq3+A2z6a70U7kdQTq4aa4SP88IouBKgM3OjzsCCxFqnzCvlRXNep
Ra4DROTpSfzT9Vba8ESPK7aJ7+ZDSAqQPR8KPP16t4k+1yWuwCSyCv/BO0/U4iF4
nIipY8B5X0WDQgWJ2nH09aGC//pjyp7ZTHLCD2zVsHHMjgh+S2ryApdhKoWUePr2
nAwYN+/GgUn+dA/XXszKw6VRAaIMLA00sqAnZkRLlGZAxqezUCm3BzuX4qMTbEw/
SNt7gcLoRt/XWLPYmyGII3N1bfXkFjHvHFuxnDF5U3bL5pKfgCBUMfIyHErOiRHx
wyIhFERnUPzoHkVcp3C2C6dBD3jBeZeiWeJ9hPR9cCLC3UqlmZj8bd7PAedcnkDW
i5PY+2es3y74rw5JoW7zqhqMUIjapcbM5IQ4P4LoGfhbkQ7cWK17Qxo4ZOyXQr6s
sEMejBafCUM92FNz0EY2QgJBOTrj4TeuvcBz1ROn7pzLgGxH6CuS4JIlcnpMko7B
sEIxJ0bJGTUZIYQ/ZDU+ptAxW97rHOGHElGvT+bXUOzXl2yH3m2aBoB9/VVlddMQ
OaO8X5yaBvVKmYFJnth0PZg/8nladp0oqkcGWOX9LonWwHy71mjYo8PvV3D1Mulv
mvtouV5vOZdJoUQ0zy3i6ZXWvigge+zjUXvzc0h8FnvnyIPrJDUrrP0EHECQ0oDQ
MY93xdalKG+hgxC0D0re256z4Zo84XewvImIn5sH+7d4Nu4IVsYy9iub8pjwVwXC
h5Y9QihSVFUc8vALajQPxeAEFmmAg163sKwVDwrz4QEFvU5OxVYCAQBH8R55+vZz
ENHHLSfktCEzq/ZPqnsyC5poclQPs8o4X5X4kRXy4VCcG7XNs6vR685NZ4mSwpQx
gan7Mh4xasfJdKaSqHsG7MFtj87a4CTBLbDAEqNvnQfE+n1I2DctxA49pfR/SGlr
t2gCGvFaGSxygeisD5wXkAZA4tNIamP1BS5pHvMOPdD5m8bSMn6znFP3Kv4+om2+
lkNegHNwxd28MpY9Qlh3tVsfTTLdpxS+bd5Qvyb/roo7KVT48SMF7aAbVhafRLMq
Zox5L8yAVkQMbjzhhrnma1yQK7bQSaaiCgmW0MtKge0WktjtFnDl+p5lbjLJ5Qq7
NG8ro/RG2fQruYY1cuQzmdWlf5lJn9mbxEiHbYELFI6f5pYJc24cQWu70I6rFR6W
kkUfJDREBXfNRE7ldknaLVuIefiA/inR61/CiFlamkZW3qgrJFtUunCFmAvTtO0E
57gAyTXJFY3um+gxFup+ESEtByYFiX00vF9O5jowBmaeW0NEnhpXoSrzXm9Pz0dV
BSGdXUy443FRU1eAi8ZMcgKO8f7aTfdzKGSKQ0+ydVzs09/qZ19yfX+sCqJV9xYO
KOM/EvJW9gvOudbtfA48NSaB89xGBkrH6KNoSgjsUSts+Q/wFrysTiUVr4Wc6mez
XMVR5wGudmQW6ulAoY274GAKjNvMuJ72iIdw8uWgxT+IzE3P+0Q8s2gyqLiVayX1
W2QD52cG1DvD1lrAx1Tu2KOfaEqQ6Ra94GYE/CTUJuyFGxYoAIaMfr1EpmyToELQ
R1yCY7dfP9niW7drimgjoBgdn0vvQiRInT6GDacvuTUvur0sWAQb9qizNIg0f0mU
bX11RwAkf7z/mIIWOvsEd1V0xfWi740ht+FlyVKcyz5JYqsOHfCie92XPBWfSsUH
umcN9eNbOUfIyFsA9SxI8hDfqUHMpXp0M5DBlyKirpsxKTcSYaLzp3K31qo3JCY/
98S8ibBSPxQwQ73PrQnzig3h99iWa9E/wBFQPcJYa7/R4dV1FqCSY1IBExTvOTC0
39SgBZinw7rUrqE0fRZg7iX7EAcZe1mfrt2sUXpLbw45qFTGrPPEojgVSrjFg68F
te6K52z4XfG28d+I5HzdgaPgvv275HHmXl6QR45PiuAIsNw5G9Qw2S30MH/1Q0Uc
qFf4N5pPtT8TrgvARkqDOQnsEQuZbtKZdbMzPrUtMCulBQRPimnTWa4cucx5e8e6
bziMDUBoxc6dF3RqVR9lbo5V8YnV5ACGFyp4pMdOcRa1Qjxj1z+ONtKlefMW9hPa
E+tKO4EG8Kotv5r9N87PzeMHQ13hBYF5ufyPn0HeVF8PeWScu+vCpFZlMGGexOzM
/qhcufJtW1+GFtA5Sh/HWbkSNrgLR/rju8Nc9G0xMSQOh7mJJKpaFccnTB2iHx4J
17TQD5T7cLIXHlE5Df+Ia0QdzR9DJA/oJhpRha55NskFkJfz7Xe4grlMAye8KlOY
ItoqWnti9U5VTZWLdt8kBBqY/W5HxbKFLE4Qo+Ko4a0rwIM5EtXtcI+OaiBRVgYl
0aTb3FMQn3aZIdDmgw+xnQ+jbm/NOBXJEzM0+VNzc1NFSiXSOvt5MLiJ3DpUcvCR
Mk2x6vVCqW4yc9fdWr+Hud3RMu5PcONlDM0IEZQ8WN/u5RtnJsMfzdSUGr+8IZpZ
xPU07Xf/sAPwSFsEHwjE8sV2sLlBwuut1kckOrqrGHlzmfHLP2ntt2IUhe3KHOe1
a+OBT1isbUGo7SkBGVAxjglyB6F0eMBJoASe/V2xk2A8sSyobKauC2w9+iqXBmJL
OI+ja4jXOnP6RN38bEMQ2J76+Vpy/NcPvx+38ecbRTq3cKu6xPs3mUHIKV3GArEa
Jeb21DX2oQRe0QJj56JlaZZKqdVcdSqUEpUagcjNspqzAFHsmEVaOiL0Jo56jwbj
p/d1gNy/VWRpMYO4MiqaqkUX2fgnxcodQceYPimlONl/lpscdYIX7sLIAcXlfce3
RqJIPLIpij63JEaoQKQcuUFf7h6iWldFUewvzcK7QGzmU1c8ct6ZWKGBdSyeom8D
g5GXPGbjTH8QbbTIdPxI9uC5/deBPZsQWnwW83oQXubpGik8m71pSPkflFN7lOpB
KFkZ2Fm1pYvRQaaNdBHBsLglmrcgXIiWKims9nekfjwrc3jBeRqBJUwlZZ230hAd
DlkpEDv30srt9IDCY4xukFFn9vdWAgWU2fzemYIGnlccyUToM1hdq12AGJ6DKIR/
ioC5+KO+1ADWZMVFyvZHnAjuAl6OJdhaPLu42NRVpZeK7HpBGNmWsolu7PeX16QU
U9bdrIjZ+NlCfkuRMfTdKBRLR5V7yYk1lt3b7RSophAgv4pV/vUodFQRJZbHki7Y
iR+7McEIvCmhpG42Tbp6ukigp7w3UtAZ/VPvCI8EznkjN/+NtJfYp8efO7TqVoqv
R80O0kpBe+kOaPk7yEZw76tbQ7L9N+oB04NQVE92FA3Rffhe7e7XDkl6LrP48GOy
y7ksfM2PHLp9y5fgQUTTkFXJdgZLZq4EIFheJ/m9q1sAmUmnHtYtAl39PzDTHE1w
ZfwpOYWfLQ1NshrNRdJ3WpH9MLJeV82Z6g7HMncTwwBK4fQxdODcKrB5HAYyp1yQ
xTwXCLQOYE//Lgm+NTAEnW3vg965eGe27C1HIlYRYCpFmv8n/Fhgw3Zd1sKNrDGK
aKykt1JKWRTkMKiWn0NAlj+XdJeGSVt2jhwrzGqEQ5ViuPEQ2/VzCaAeyFeXFPHJ
w3lR5HdnhdQEfAHndiloemicNIL2cADvib9ds0iXpFn6L2XPT2iAbVly6ks5UaHg
awbgufJBwwBCG2tu1WuKC9qwnirSau3HHWEYdKclEtz16f4gea2zoAbOpY3IUDFf
BmvZy8bKjiooVXNoraFRpMJT6DJXnUGisClmo1iLBMJmja3ugFJS45VvEmKw0Cdc
kG/0azXRDqlUA2kNVHTe2wLSEi4O75CaIM+d8K/dXY1tcvkJP057lw5N5ndECRP+
zSqTl6VT5vVXgkSbbzCk8zTyJrvX7ZrrOvpl9Hi6K5FZpBRSG1w8GS5h1EcnAT2E
cAfUC3dip6y2F+l0B7eLnYPtWBT8VhTPt5paMo37ySRHjUBGK8k1QWQG013Wj58T
lFxbwBDn4K3Nors1TMc6z3ELUy/NE/W7mB6S2b3SL1eadOTu2RoPo+7RKyMJvLvl
PMeTI3RjI4r9lJKTfN7NNbXE2weQFIEo3znDaFfNHKvr+WLF5opvKs0tYIEWh3mx
WjKCV02JcUPpIMn0oQUZoK9dkj3D/LHA0/GWJ2C2jmgPqT8WEbYmLqV1gGPmXwPY
VEFMS1pp/IyuUW92ULspmam6in0mm+6AnJSdjghz4zQSmbHM5WW6XaW2bqPWpmMn
ZMOssMeGsToSzN/+3pti0hX0juQgMdE5GFc3GvmvSuOSIDEk3e6w38JbEeLUTAxQ
0qbc6FtRWUAM6ort03CvfmWXwfvA3jwGGY1c0fkvA3I8GCKdR1HcgxzwMRLG3zlU
gj/uCFrBhQ1spC16yorcMjI2obZXOwWYqWLhPG3nFzxGvBNykKtU112f7F1HX6Kq
O1PO92GF1JblPeDe2FUtgsFrBmKOI833B4YWA1ogleWRlF1fWzzgzI+EFZB60c5j
rlVTyFB+bPOVq3SFKgYQ5k34dKEVuVZ7mfDitu2/VaOzX+wnxDx9eU/YgfNXrjVH
b04zyV1DdgJ7DhN5RhuVgFXRGaHjtLgSNqewJFrN8EqtfzSgwzbgu0WWuuzaYScR
iF20ug5i8UtmZH+aqFP3/X9uozAueHqIUkTBorUkVfthd9arO7m26oZIl3p3xZW5
2O00bVsXFYHJG+SMHUtlheU9v8T+I4gm+ce2jm4mmBTOdZvGegyP+FCFTYccE8NR
kJKRHWVIGmuiBfIJZ8BxHK7Yrpp68lLosdyOV7uMCXyWg+EN8GJ/MYhenyYCTcF2
lJ7cyKC5oEdGZrTCvrrB69g0ehIQhXpp6cBxEfPpb7VWCWqrEbWK4LGiHqcmP9NS
j7CR0fbLcY/rj39GHATDllsKjk564ZGrwzvHlAmbYNKftJHsTXYaO6TtbjJ/mMVM
+ZP9d+q+Zp5B+aHKVmIlv00ZA5xtyyPvqNBakBEoU2PgI6x4DS2O3r+ddzz1eNiU
JeU1FaaTW110sxBNoDN41Nls9i2327z4SbMF4oTR0xP1dNkCCWR8gu4iciPk571+
yZoBwoWqqPzvebe65+K8LVMR2tXcyMIUf/Ndi5eWJuVFSyMooKEdzltmO/Wmsuv/
6zOcxJBBk1P523e/a4LJI29Ng3fAVxnE/h2Nb69kkpqcsmL5fRWnRoc5kA1hCKOj
k2P8wepLaLGccJUWW4BTKt9jMw/QvllTrl1WDqMCrMWtLQryIRuOLJbqK6HVuOZY
3qdZOhoclq4FOWnxXZfjrwo+qWepJj8bvzyAVunnGvAQ9fn8Ngk7VXY4a/lVodCB
4QxOrrRIZvu27odRPFijOtKSWy2LVk3vnL9nL6EpOwahF9gKpn5EAFO5a8lsbWgu
lL8h7jZb+5+G+6n4satx9/BCSmPzifE+0w4puq1wZkyN/72CrLlgZYGR+Uf8TPuu
0wVWMjCKTYJ88NcBAhZfJlku86YYFZkpkspzfm7k4n0dKADYZ9t0GUhfLryM1Eex
/Xl2QJV4G/hdyl0gWAiN/3dW9j3EhNSbND+AtB8ve+Ws4BtNdgmLkW5RTpdZWxP4
rj9Nk6GfpQ2X4YhptxD00HK+U4NgNohnoY1kLMRlJYzS6Aky0W9VnudObFVvw1eH
ZrsQvTd6ZAM+AKGne6XABtGTxEBBnZjmN1wkpzTCAQ+YwWE/f/OLw7KL0JHbpSq5
wmTYXvJMLo8I5ocja8k+6FHZ3OkwpHNVVmYzdybEAV77aCJXb+MZGoW8xcBn6WWN
31VlIFzBrJ5vWk/L6orRoPcMMmg41RoGAXS6iDNEltHa/2lX8QXNWVs5HnjWTVXZ
25vncnLTabXwDW+sr1YAV9uyYeCVhbKJRntCC/GX29xSSpoFyAsYpclNLDgs2JM6
WY9mFvCX6T6HGaxv8wsurKi7HZzGw2q0qlbO5sX2UzWKNk4+kd3O0R/gzcgWs0Ya
uiw/+Of5opUtZPosyIG01tSUfKFF3St7xdFpIUspex/LO4WLa5NLCF9majcuidQO
DXsOUKoo98JElWHJ0QT7mS3w2Y0VLrLNYC8EsRX7W9xErEo495AI9GjNDLo2GtdS
/BdDE8u5+IKIzQV+4KKeRA2u4HocNJtx1REwVZFFt4VJ0bvvNNnBmQVDkOHyyVEX
28zxiF60ROVPjBYX0xW/cpGIXdA81Ez2hCPnCKZUHH9Xs+EeUw9zNsYzCFI3I2Nu
bTjhPknXRdcPe3sVZ9aBcAN09OvRBr8hfFYHqHmWCL8gFpsRtWx7RJNHPefeaTBn
+5MrRMXyABHXy8JyPzTa/cDANt1Wv1uhV8CNacygjlon4l/UqO1DU+bYId/F7pBN
mJW6cuetGzCoGLf8E/YpcMOWd/g0HRQUq4fqNlDaQx/3GrzcuKYAYXTFAYDY+fbp
7jFxqXHIju10/pn4iXtBKILBJ0hr5wkoFn+dMK/GJi1xf49jQw2ePeOKo9bC24jd
5IV9vUu5X3zgZfThWooqusxwrfvsU9Sskcn/fvxlLbkRZD9jt07sgOcXNexXLM97
14P6Lt3xuyFPwVTJYg173IhB70/zS4YkpnhsSOt6tCdS49CkzgJd1gmkWtx3Q0DA
uyvt6KqmIaEHy8l6hk+x3LRM7zybmUIbMIJTh8uwNE2lPXIzGln7imo+QlxgbqcN
yqptJIMLqcMIXjwR9fQQvG7xtX/9IgqzncnE8ORbcYam6MVn4Mqf04DYLXMOb1kz
IlUH5WqMAUrI6YlHl0ra1zc2jBaOmCV/3klwGX8vcRrZvLh2nLKgBco9ltR4dUd1
3yHMbKaWovLUkLfyhSrUXM+nqYJExRhqBSWxYFwwxaiMK6LlYXUvertv5lsJXDkg
gt211knYheTaDD+0YIVSYpBgZ+EurzAwlLaJyEw86gL/ZWrVkFQ8qrEx7pf0bXG2
oHyUcpwokFYIxopoZuevlt4p1Z/qO1gJqhyvxe8O+XvT4SqriSu0kJIBMG3fRe5d
V9uov/IvUoowytJ84yubZ5ecMcRjKcWbtQp8UGldxEJwGYP9Cnepb4tUdvPZXoJT
FGtNSzWJeAQEPNzMa2xVrCFIssLHcrSyOPEdEdSnVVPoAwTDBXsPZZg24bRkBE06
A+hmweggImg089A8TFbLq9g/3WQ3gl4whmPfuaXpQFf9wQPgIV6Ax6etrOLAuQui
qvr7hOWVes1reaWNLw5Tl/DiO91FjgcsswMGDMvgjRIpZAK2QmrchM1zjcrTzHio
rFxapQS17y0olHoC3/EVK1wTyKr6xtZz7fuV4X7f5WrXc2CdcLsynAs1Rp3X1Nf0
cwEkxUZlzX3MBuktdvp2+zzI/VhO3HsXyB96mOm2TKctH681XtGi5yIb8hagyHFd
B9X8so8ysyf52ddCPj3/09a7KdAJpblXQyGiI6CPCrLL0cpkbHcPm9MvOVNP/7cH
CaoDyJBKHGhwt4ojroQbT9M7TIRKyYUOAobdnNdGcahHle0B9/2QF1usaNa1ka4U
bHJIQogGzXOGReoI0iGf8Q5ZvJ4nHYlNqbgTafUplJaM2E0Vbw/iXyiR8gVqi+xB
0i2FUdGBrpuh4HlEfPa3zlRgDww4Szhb1Qv9QXZD4wAFRlLeh8lNevLAubln1CZm
I4on5tQiRzL/b1tFVhkhQNtktX52Z4btZHnnw1jWkfnsvJRrB6lwx1kDFufG52My
gqA0Ty3cMU6hJfRkGR7nESV8hzzDMLU/W23ipqd9R+x/BBnNYsWv6FgakjT140qw
+V5zXomOztf7r5FoK4LwHfqkMo6k7zGguOqlwOOiV/2zEmuiMTFPCsbvGvK+M3Ll
LK2jmb1QHF0OgqPatarWL95rmaB/YBwYszIIOemBgNX6aoffme7NaNs7JhhruWW/
U5pMQAp84cxYYmk1N90svMXyU3T5p4bU+EVhCOQPx3dBaeg24ioYocS0SQheGoWe
OCDbMNdrNcvJAsMFQGRphgwgaP2rZ9YaZ3S8GbOBN3lttWDTERDmgyxoZLP6xwdW
Ob8eWKOB22iHBWm7zkTVLScqCqjvinR10cDy1Be873h21UDFuyXNyGDBBNhTiOIo
ZvzlPu6hkDMFA9L6i0iOH5voyPAOChmppX8jMMfyBJQJoZK5fiPT8UW9OcByEJ/j
RzAkDSwogIMlSa9drBCnm/XgYOiTy/2TshmoJX8WaNMEp4J2Vxq1/iOrhZKUYN6w
TUM13djXT4qvyLyLu0FRL8yldWEjLycxhqCs3ZANB0xOQRH+957yva/p2Om8Euda
2muRP61VWh6T5+j4EgXhr5UPTnnqSlmF5xQBzaT2EVIPtTvvP6HV8/q0/GpfCEQd
KLR3Lwg+q71nk3p3ruIehogRm7KyLZ0FHfR2YEkOqQ9w0WFIOf6ttW66rrITplK/
MyLSl8NcYezUDfjBCmebb7XHULC1ApxZJmde2/D1pFB9G17nzspxe/78sgs9cHYz
FqD1DBx9AooVwCXUkIa4gl1yyrZiKL8JG/L7GEsWk9N701oiZH/JvIQ6Ncq9Nnvn
oIwNb/d/f3TvRuZ9D7YFeJeppuDGgmLD2hiYxjtbGNjxxngsA9VN8X983KVDRSXE
3sipA7a8UjRoG7JpksnDGpoL/cSCaShLw9S2iXvU9ELBKdaczHF4gsZzujRaw7oj
iewTrkH6ANbjNzL8AFpPZ5YI/GPvFE/Y3AylKiCGnUqGnRTsfcVlME/bdTcogges
NK1uYV/MIpwmBjZZONOTWP5uH96mfqoX0QcxISn8aqnUkBDFkypeWQpkiYh/hyOH
TYhrW1xXnTb/W3U7wfR3xv1rWldshUsmiqs4WfGUew9dCdW2jdSt0/AS84nh8/3c
04mTDRXhRhjm7AIXDavDSkS/Qi++liyBA0HACQpKIHL3UxVGjAQssw/PNE4bfjPZ
gCiFHlLQ2vw9AfcpXD7/Wco5BVjDYvggd4opa91UqqfkRIzEFBaI5v4yGGnaSTLY
RPbY5uRCijGxM8d8WtCmASP3uVmcWAzTpyxfp/GFfDNiL6yHduyDEB39mPqQrDLt
mmlmG9qJ7BdBWREev4eQTxW5gBTBsuliA8iPWZto1v8WLitx45ttqsNFpuhpK0RE
cHKF8PYOr8JLFG4i9C5dwc/NlkVRBRLiI3gUsLOpQQqp7p1CrdL7CPdP6gzvKZBF
cs4b+idcmE8Gys0kxIC2jH/oBccZHsv6b7dbJ9wT+A0+KRAktBHiZ7Dsk+5pNM/l
dIHf0BIZ1SylQ9osEZERYEC8h8HZBgR2IVvwN+a8/FkvwEc7KdtIAgTpWj36oacL
8LoZF1WGfX1V9DVWCQyVRjuZJcPtD3WtmLJNZLUMowoq1nCYCtfFTRKFfrcmjFvk
Eu0qiiiUnOLtDm9C8XKWh4eveMFZzVlFne7Q/Qc1ydDgQmX5xWbzkShqM1iar4i5
fLLt1xrN/FJ+DrUKM49Lc6mnbWpuxO5uFEBTm3V3lFAyYlERoEscj3tTKcgwFCe4
koR4dEVj+pXTkV1zgCLy3vhnewp8abm1VyT7YCc39P5O8m/7NMdpld9u5CsGmGY8
RWZ65IL99yFiSscnE4tei7yGXaf63vZncN9E/ViLxVtJdOE4LVx+RsFxQsTyw3aY
0NlkUYpyvAbnuRRnrfXB/kGMdinf+Egt1r2k/s6GWxqFSrEWfiQASYQlOd7gMckw
DP7G4K31BNKMTrG8osJLyeeqHsFsWFctH1cwKHhmFolIcNzf+1pyBfSqgHeOtvO6
q/jq9t5h+fK0Qm1v+WMlMApfUhVoL4nZLVQAwyJiFxTz3zqv/0WAjvxo7g9hmsKq
o0fmGepV3DPq2sybGy0WI8dzj+iv4o1XOQNnUU2x9ryRf767W1ITesFDpuPo00J4
hKx8aotNlNzZyUBop7xiM0083uDyLkGNel1KdKR73vOefrLRbW0HA/lySANZUGfQ
VVIh3q6JMAM1vJ0ie0tEfELHIS9h7JXmijTRV+0omwkYqhE3z6Mb51hposmSvt9D
B9UqMKSWydCcQDy87tlTK/nCEhB3kFUDKjnjT+HfPptVKiWQShx0IyyPP2+hwYrq
vyHYzq40A4kUEJBL9dQHnOBB4hjGXHRP3xb+vDXNjiklj69JUhyjXcG3BSygbDjG
iN8RY1JaVt3aAqF6zm6w2Q85Zk+lPhNIYETyqLvQyTcv4+b/GDql+6XibukF8BrX
7vTZK/UUYXONEdiIzXfmt7uNecIFhOFcwWRKlMkjICEpvamiZKq9NCRQ6sAU4BGw
Lbz3Y8sxVwemhem/6P5QjiQNM+mS5riIk/zgg+9K8NLkGO3ry7HUnYjrjb86SE0x
Kn+MECED1zdJ8BHLdcZNfstOjvsE1Lv/69rMMJ0IBbbVTyVcSDvRP5slehhtFA1z
QCRUUEyBx85Y9cJqU4O4MLttJoAQX+1kFz50W13+TvXM6o8M8lgqhwmfIecE+Q4Q
PfaWvwzeoqbeFFvkgpFGgN+6rnOV10hqoA7Dszt7agI8AS02k6EpQ+p4SuJXODO2
gf/mOmWH1xc39yr3HgNzgpg2F/5hSKg69bNxzzi3RlUL2FKE7fK+RlxkrHCKSEVW
LD3IzEuMDaYb5mlfK82rfFNk+4yTYqehhucPso2D1kRTgZi9ujyMUOJkgWdzPMA7
kLcXOZT4DxHXc6bixEYrDdlaV+zzdIpzuTHweeHXcfbatnVYoZPX1Uqjn1MGxVBV
cTuS1xWHJNAVzvd3SoJfj0GKP68OJbcpFXOFsWAK4fmrQDo/VNA9Ad37hcgyyY1b
rNWg/f7dTCydwQzZYrFErEDoMsuVDs2fQzPJuqWbBp6AvjxczZfo6idNBHsE9pFh
bQ6Wcta+3yz0DfmN9f1j7zBauDpartBLyb/4Vzk9Usi1YibQoI+xeH0ow7Sp0m1p
VI23ObwbOjLEQ6r7VG4Gouu1B8duJl7UbfPAh6q5QA0drF+7CIhWK8VawG10nBEq
L2HT5AGDi4mPcJ4PQTofCuSSdGRSpAG6u++5wINIwy6zcp2uhN9vHw1w64C1XElu
VTPIwybRS68vn09aiRfQZAUOfNMJhN91qH8vRd1y5mGBSYk6AEHAg0RW+a7NBg9c
NehUPGigoLTz43ix2+Pv7Gn0b6rVWCNkjc6T2XnYLsQ+T4eo4kF6oUtwgAvg4iw+
+C2ACH1gZu+u/U9Y2PiysNVV+hUGdBLB/oQ/yS/PKwNIgw7WeuIaURPgqnpAF/Mj
FBHn/BBbc02PFjUtpNJxpMunt7KdwHJN5Gs274Zmk/7IVOQyv8huc8nO34TmlJwN
sr+3ZhfL+SOAMLK5Ao3jkkvfDDoir1TvJjVbc25TrVaOv+9eTFRxFSYzrY7Ix0zb
gNhPrvinWrNp4LLA1FhE+HHB9mmykUqPeBMzjubquHR5kbBX37VwKgsEyVxS0AJX
BzuG6it08KsLzBivu1cqoK3TuQDhaiwYbxipV+pXhPBV60nt7oBlxKb0T2kMjbUZ
/P/R3WbEnFFcLpIM/jMi+tlC5KmAcwWryvXM6YBOO+UyRwyBwwf+m84wwP/KHg3M
UlgRtBuvSjJJNIaqW35wqxFtxrmbjZPcc1t/wjthx+8QegfyeLjtIXkHlh6YFrWG
Jmfjt5QcrkjyywykX7Kt6WEODYiPzqrwvAflLLEOokeYZPwtEpS/K+R4xuLQcp4y
CLr/C8O1riw1XOwcSP4xE2Bh3phrP4HZUNf1Q9pnp3/yy4fK4aHRsmZJlbiAmZgX
YzrmjbyA+JZCy5FpmTDMx7MdUYM6hBXDSjESx+fJ4QVkadulgYU8bNQvkixLog3J
5ZSTiCKGROeo5gfDSuECSnWJ+4fHRccrJIbnlPLvKXteTeEKlR02/1TZiIfASaa+
xjHbH+n3YRtUOShr4wuDb+L+zJ52+pKnMTlJWnN3SX4535AXhmKRdrvR/pc/S0HR
9TZxXJNIi9WmTYLBmy274USnttKQ31w2HkXBb2bFpOuRPp5TeV+QDJJc4RDMsLGu
G3GOgXiHjrvM2Q3gh5E25P7gM0g5ZyLArwHmy4sEIK7CZHGOYbMCU6520JL68DCL
M/cmEmHZ0G+uGoXAG7tg8zwBZIBtR9BAPWKOSsV6ZsJUuFKEqnZGjLCjN7R86BbW
iaSWhZDIASxXpBlha5Eih8po+0ddYFUuNfSTu595bXwP0oDL0XqaxrH+uHaCdHbJ
URyH+hwHaMgselwWA8Jv9Me7gCyS87WPMCpo8gFSlHH6RAiYmdKqXxyTOQjPfnRG
tv8fUXm4gekCJDerl/N0XAfOeHVr1XEwZXXepVY4ew6HEeRi+VrhWeljPIlQkjee
DfS/nf3PQe4O6gnf34jyA1GoZ8AU/Y4mdb6ikMrqIDDA4D3u4eQsb+KbF7Fxs58F
VU7Y1UF1NtjwiYO9p7Y2Rl5IaGr9/IXeYTQTQGTKd61Bt9QtgBHYfG6GXhrza2My
PjpIWhcuKEbOetVjbpIA9Ze6jMUncCquFndAvxrXOrEnXB7Mvt9x+PLESuThQ2vr
oWdkP+0a3nmJdDv1lCJMYC0dm4C5KWfoAQ09sHjZQo/TUs0IH9HTkZTz7hA0SHAf
CZInoVXrP+Q86/DIdgBk/NTNLvJGwPgYd+0GQUfw6rEV4ERFosrPx+sTwIpLqeB5
RBytfsebJYqdbP/1dg9YfYR/4cdacu76vkQViof5aw8/v+VJfhxrPP0yr3hSoeUd
3zL9qsxcMsSiBZ3rNAqoM40io637C248AsYD7i1TeKQR9y0+wYfwFQwNXfTfNJjE
uKOqZ62Zc4g9vEoPwhrC0gdpnl7V0AclgdnTZf+DBJV1oK0ymuqjv2C/qfRmbIdj
SBlH37k9v051plD9mr9qNZm3+98isZlMW2s8+rUZ6pHJ0sF6EhpaTBfCqGoGEcVE
S8+g/ZiLeCWL/Au9lrVtC1pGZuCOKTAuKbT8Gxi46HOhkU9wRPhDkr+jhAo08lDD
ZP1fspj4ln3v8gJIAiyXZ9Ib7wUT9w0UZgg/CS5MkVOIZYhVPQIgG/kug43ZcHm/
W37aAS6VWoVpCQkNp/3xtn7CmfGbR7SZoFlDO1yVZ9eEnYpzIUk2SNmz6pkksXoG
E1APTFA2UmDT9vgB+owovSdVuezPZvNAaCvDVv1wLW1GSCmVaEIO0ub4sXc2j7aE
F3+hJIhOk0t5Tr904nUU5AsPl7vUCrPdHAi68rw7lY7Or+f51EM/rDxSth8FNxka
I3hGt3g/ptC5Yk3PhXTcmJQWlOP1xkMpF0+mILoSd9AJydo+HQmiryhG4i/xIbgo
uB8q4nv+V9LJynKnsUoJH3yI6gfCwnBC9SRVvgRIRd5l7B9rk0D+3Bmb26Nssp39
9rSS7xm8G++B/+3v76ZBWEMJMusr3DIWR+4RWOgxbEMWOY5KRE4beBCxqK42yohD
CCyOgm5tDdBRmipeQnGz9lGuY2t5xsIJnHH5trdDI1zPAuSHXRBOr5BGfNULUc1T
g7dPq1HekkSv0cBjhvdVKjZMpZYx1vt+M47Cyvs+jWYlAU7x1ufvbes8hxwgWR+6
ARi0J6XEJwjYsmJVE3VMt4+OWC1kcqpFpCHoZstBzMSQjuGmVHOtpqwdGG6WgxOI
2C7oAyFOYOkLv4FkHfnV4s4fOElkQ8xI/jpvFHq66UdqcG160g5UTv/aA70TtNQo
PP6DVCamXyDxfLOj8LK/Y44QaLCwtZvdFC/IJUx4Qer+M5ZYl05ukOvKYxjQvPnM
IBH2kE8Q4g42WOXTG59INrjkr/T/BehklVE603emYJIP7RwOCHjCLJphCwY4dtY5
RQ9UanvmBW1y83z8zt7xJYWb9Cz17V6OcSZrPusB5yTuGKKHoql12n/c3RsKlgL8
tzb8wDMkVSAMoe8be09UX9tCrGlythr3uu6Oke/WngNsYQm1nBdxdHN3rVk0Wofy
9XBuC+33yuFjRx6fcP0gIgX56nidtAlW8jXfiXM0rBEKNlUfFSfx7mfH6lOTX6JI
4/LDmLIKqwj+2xp+irf7kOJpVdycUiLSmm9Tqbv68RBcAkuDbgq/KyBID+d5i1bu
D2k/H8Bn8ZzxYtRCkE0TaSef23sIRnA2f83yTGHCRlHtwx1knBYGsycZ5sWq7MqR
1cJ1vPJ9JiJ6wD6c4rP+aJdatO5lR+RNfsbu3UkLVslPP2RYquoiel72UcM4slsX
fD5GfxcH9fCq/tXOj7JMko9+hgRJbmueev4X5K/R6DeIUJZ7wHrLvt+BPxjyZgU5
nfRqFHl6iKdUaSgzhDKirmwMYgdUaXRxX1dmHq4mgwHu1jbzSns8ah5y6cmlQooc
cEeydR+VAWM9330x5LBKyHLkWyudvalN4hoc15E9Lab+cNGddN4Ha4FFkWEfLFhu
Dup2VOeqJW2eNQ5HCfxCL8fmhA6oRZMeN/zL4xdi1gY5aaNd21sRB1kCTULyAXyz
6bT3zRUE7pq9JNmDVsrDNyU9cs/Sc8cx3fMjeim7w20jewwiUpxElE/2KrO2Uoex
ZHTt2H+tMj936t4q1+jR3rCQQ6RGGZjG5KoBXiUKJHWxbuQxQxNabA1LFYSGIOwS
PJGC7a/t5KdBNnKKXrSwKkIurcANzh+mwRdK+FGHynGO0tdunQqJUBVpB8kEJ6cC
WbyT5EcoyaN/lvwZZSvsLE6NcDtJIhOFWiIHhzpqksX6DjtZVAQDKK/TB9yYUpws
UzvNB8g4EdGyaoRglHey7cx/DN//JMAGRl4sJoKtquafljbVDOxhZm1WbE9r2y/J
nYBL6fpqJPiboi5DXG3woLkmMCiTkHfAvewvc8gl4ULII7om96xrz1pcrjo0HfRk
jRtMVNjvLdjRypTJ27XioepwVqidQ8qzzNwCwsQz6Fe2QVvsdb7bx08KYqrdjQs6
EpcUVXe1c4jOAtrHnwDNzoKdb1chjQ0jODecvPCJvgjkrgz4VE6wIxzAJkJxZxkw
/pd5uSp/oaE86JR27GgfA8lsGeQGun1AvDcjJXdEVgv4hnzHcdH6mm3E+bxt38Kg
a/9d4wgKHw5CK1o+0LkWAcEKx8QeN+Q95ULrFwqx3walR01DNTtzromTD6igizPt
fGtcm+veMNoGGR/XpItkFGayt8mm+Msh/hTbHnV8HYjGR6sf3ZCQ25uFkoXzu248
frrztzrM9ET4P3CuiBX+VmbboBw28TgssVmxC/kTeB+QuZKxt9hvyPn+ZMWvSBr3
9aupJA4Mjh8oz9DlfgnT3xGXxhYUpJXyLyeiT3ADZmtLiECBpxSwTNDHF7dVmp68
so0XIR8FISTsfyq8vXR3i8A9MfD491/aTntnS6X43tDKBbG2PE0FebIfFJBR9bB/
DF/r2LTiEkYISOF1kc4K0qRyGHvOSuQiO0li/uaszh/MvmqQDLS83ZMl9ewVegBb
vlZJACLvwERVc7L5ezXS/Rzw46BbfA79qF2x4RFEnNk35fumB9ov8+DT+YxUkZL3
GXXxqSyO2JUQ4arxfKy5YP8QVSBWVVBeUE0CYyUIVp1HpFCF+sjC/pK+xFMDz6/O
QoC5mh9YFcs4AzS2ic9eKywGvo6kZ1yrYZlCYglOtBxlKaqnIkmZ3A43wqf6lDgt
EHeZ+11scTT5QHmFJkzTXEBYhBUCxv93DI1rx5a/PcW2PBhUzfYnKyC1eGCu1plP
ojxLi6M05Cx925bOjy5EGnXujWgT8B/+D245Kiog96O6uIOF18lh21b23qpCA4oZ
2vzeN7bfrjM58RWxmQR+KTjfjWLFGoSDaO93vCmHRin4+YmOosoX3MoMU5AFVXKc
eeQ8/LYseW3eJlgXskQF5HmaqDl/I0XKClYp6rkWvyr2vNb5GMUrZwpyHgRC5pSn
EdtitMjyCXgmxBbSpC9hUrYfxq1IJ3YmF//XjuSuInszsyTG1pItQQckBYpBK8ql
d0FIIazlOWEJWsKrHU545UYIEDgXJyKLySu6OgNnzzJYAGvJ973QvRYn2zjkT0r0
HMVZvUM4ye3UkzcgMOEZaFy6mjFEp4nm50DvFqbuRSB8fw0dQuLJQaQzQYZYNmwA
7ZGS1Pj/c9Np1L4MxzvOIyCCwUQSLCUBLYlPa7V7ht2UnVdfXKIIfDnr5ISjfK66
sCmX4rZBHY1SuKC8IYOG7ykd1AS+lyRMYoO1yq3kx7vs1U43+E7IbCyBnh25JsKP
bmqDYKXFun/JgOEVuni2sNfOt5lQEb3mPw7do/jo3DOYKi2Oscu4kzw6lwmwLYk9
9QIphLEBCjF6+UvGrEYtoyZ/p/hsga+MYBxNUFC291uWA6rOls749+5c7ppWOMqJ
QfPZBAtrMcjCUlDVyjZSPGIlAqzAPgVO9F6v3lvG4TM+H8zd84AHM3HJLI4OJpLP
oTglUBp83C0nNmNoxrIPqRj2Zdid0qL4xH7Uh1Mtn07s5Irzjuxkz9it70ofpC7O
fEmIiNbyApKyIHs87qnro27aG0ALHTCSa754MkfzG/9v7eTUyOFjEjzy+VfpezQ9
TH4NtJy4vJcVy5XDVfICTQDi3yMteHCQ3rkG5sUz3X5VQytP9C1MVWl5NkqLHXuk
KcFyrLyMCnkJPy9xEE2PcEGU+pIdrJA4lsUNTc63Nbc92u3putFFiQW/LC1vpFr5
+V8Vwuxd+df366UGE/y+v3OlCEB/IZccjdyzh4DVsn4BDDozVNn8dspINSbOENMW
6LS3VG9CoqOwfM+xnjv51zgnEL8/fVNZdKMJPLu0alILh7JDDqwSYeASjiWUWAiJ
83rZUjpone2HkMQXBfkjafRYwZc5uBdMXD59SYc5hQJN8uWjpbokj2BxKouNiRVq
sCZ7Ju3eONosyV7qlZohnxLdNYTbWdjGwKzRJ8QwklKPWd+BmqucQ0nXmOTgO4IS
xYOdMqWgqzg/yqYr/b2VNx5hA/nN45bd/j1g1BgazQBsDrZ8Qm2ZWj7Bej/OHn77
+r91jbwO7djM4isD4vLzfX89B1iNRlJydDwwG2khalKE34iMWtzC8NfrUysU6qlu
MpLdSiH+0ACWtfvkg2ki9rxq4TYS+kFeBb8h/TuSFFyRetAAaFU+A/tRacYsFn4T
LD2PqPbBN6lD4XP5zCCLnHAap79IH6DqN7Ih1mofirD/KF8deOJdkBefPlvD5j3w
o+r+L6XtJ1nAj5J65BrN+snMs0bpgOWEAw3EJF8mXRKkST5EMBf1qA7gmCuAqail
1j+YalAcF+DAcnJSwCjbGIReEqZqCkUUHqeyj+iaS+ZgRWDzcAOU/mGSoF4kQUHq
xyPkHYzYg9w6YWu2kCIEN3mIITreTJ47EfxdTOWWWeBpH35a24EWQ9UZQbPizRvc
UdKH7EnrD0ApmnOPFtUCwi0aO5UsnzaAM6JnPS6BixOaK+Kox7rIZvHyUGUjkyYj
r0s83Wl64PkRGZWM3nyq6b4zBe53y09Mk/MZNKJvaEI38budqI9MWLpCQYVxwdVn
ixYhg8xI21lvsHZtGfsfIEPLZqAgI0yUMAMwz9v1qTcYcNCJH2k8zVO4iLe2hA1u
Eel3zk7tp9LsM+JaOPljovGJmAW1aBJLaSsT2m/pEz1tbmTG3XAELHgvZWByJigY
JWZ8X0AUJX2wEcryhzHp+cpSAjPm2I0RW2KO8keECWVeK1Ll73kUdU7AK23akIpp
r3mzAFvOhmUDW/FsebwzObE45gaiiEyswrg3OKsi72ZY9Qmw6dundr0qtz9+iwgM
A76i5t1iwAeyGNGElnT6CMpH5RuBteKLFRUfsYQx3oIu5HoAEqnvzHdug1JYMaoS
jKyThBb/LSRq1YwewN/bccolP7qS2A+FZDNr37K9Uk/X/lvo9YKQM8TsIeR02T/w
ldcmU6IGIO2YvsBjr+5WyGScWhwSXYqDu2tCQmvnDiwBd5jdXtzXK7BikAurkGTY
tkqMImQ1y6DFRB4PGmhQDMc9Uxi1Ow31EthWSZyXzmTyBnXoAtTzqmq6Fb8q6X8J
1pC1MS7QZZjZPR+eiOUGJ2KGimsjfxBdhMc5f4selyN9lDzktNPlDEZFNPb0oI3q
tc8tVZ0L+Om6O+KfZZNGqEC2CorfSZw/3/2ALH+60VPaABD4EMBYmC9rh10eriPF
aT9zjcDovAUtnZ4L3MgnzAP3g+Msbv/AzmiJQKBuX8p78/uZB4k1XKIHVArVRjyt
MCg7Husr0HDSSAm0th6a+y5+kS+i+FwaRn+o6NFPKGe3WuRP2zesCto22CEqFcwN
dNlPs1XznThHvhRySx5VEQCeuUdYGVmgwlXoou8uomqHltE5R2hseaffnrVdqBHD
IPoQjufwUj01yLQDVWnpmDLd2xGB4HNaZP1PU/UHsLgUfh0nA5BLPY7Zm+nCPBsJ
i1jt3fMd2EaKI+TYKDuuqw5lly4E/kO49CFBkbKi3b+1ozujSinSrX4RkWLneYlY
PHElmQGd5W+QYlGvdu/BdFMXDuTlCJ1SNQWy4KiMVy192FtBKMHoKTKLnc2ZeOMH
4cM8XYeE5RhiPhskYgzTlf9AXLRKpPCfpPV7n6OLMboF4YYd62mIQXRSCFSBmVWD
VZLORLDHLCkxLeNwbP3uZb0Hu7uVFHwxltrljmhm1qBwcMY6+rlFZj4isNoHfssZ
IzxZQpDGxpNjQeGsgKhQkb3wpArn0tgG5QRjp5VUBXA/k+rrsyjj2HhFqRlyaDlL
KvNOU02VMeAUfm/aF2tW2Y9q3CAr807b0iXXcZREPT2enIjuq+yEJRKz3qvwwHA1
kObtFJXr/0rAqbSFfoOiXi3Qnz29MWWi7FaPZCOWUuhx5yZtxlx1MUBQ35po5Jtt
o0t+yxrFQmmDiFLYeRaNBZ+2qLhlYj+WoOjtm8ENXbvtBuXVMFF339YOE20+2WHl
zU+88mb1MuBN6tsVoNstpS9XI0aeEzh1cDuhwyWllzSNjfFQH9wGs2rF4POOSo7R
GMCWnuUztYce8Frb791DwCP1bO9zcm0t8i+1jt2btthOEC4Kh0F5HKo+i2FsR7EP
5nS+ZX78cV3pNUDL4+Tb8PTKCWC81pVCNlZQAvUMIGL8jVxs1/ObxKj9iLEdLymK
qw3Bhpw+T56gOo6b524fylV7iIkx0rxAYYUqo/MP1AZdKjx2SDmK5FdCcPmyYYqt
nUKcB8zw1ppTaYyvr3s/Ma7dpvToWw3taaUu8o4TvjdgOFtJq+bRyUekaaoqQqRL
GecN6v8jtS5T/4G/vEIII2bVKfNtKnNrG//sh4hoFd4NT0ILzhbSyXz54amlUzK9
KdYahpVFU3pQR+2OaFhZrlENS6iyYDrYyMyTdRMKPdOBGmGmvVl6poHJ9rXB1csG
MEe41ZGZyGhnffFIMIPhIdO4LJaAk5gNizioRFHJ/nXXGiDFcb3JVnxGWQ1D+cza
s0aNWQyLXHjtldBkNJ0WR2U+Yc7Nm5xUBR+JlVotUC8nG0IgJyQxO0uj3pIXHbPA
4m4zYdkq2aD00wyga26cyMd+b3KMNbI2LRJE9AmNJOgTjeWK3kcy+fXBQ3uObtQG
1sJ2nV+9KmuEJdb41QIaSbivLJbTxs9tu14/nHiLlBznzyCFlKNV0iPFcrVC4WLJ
uvyhzH5gyo1Ekpm5qk1/DmaWtHvRAvLxOn3+WnSGhDkZqi9G088vqYKoMzeDQJyL
HcNaIT+onQAnP3VTJuR8rIcueAr+9Y1xgasf6H8KPtCUxt7pfOfJRqsP1HZWGEJZ
cnhhaz7CHF9YF5z3NTe5Co+NFKbVvi7dl6lGTw0m9zmxf1E+L9IMVZj1ZQqjtOSj
TeClhwsfZqGLph8pFxDSUgqK1TdytNKDbzMEN/YDKg7ELZ7TJcMFKdJtkPkm537B
2/xXlALda2h6gDvbT7bavBRCAaPzF21neD0z2CsHXw29i2UgslUbmuA6qCV0aa3L
C8ak9Oz0a3CeC67zZ/W5fzelrhFoPrITpeSPl0N/9GBALeWp7s5QDpJEV9ICUwXV
/juQQnyqx56lOGGvJ+oipmd3lOC7U1IQgbRS7j5WhqZPvHhjSQ/cgYe5anMbVU1w
Kc67ffJYxheIeeMape2ysC3lvDnNHdmSTwvJghfBu9FawjGDiqb46IUi7WVvBAVL
CxbMyjocslx7O/vI82U1Dz/Rn2re5tLHUOg6a8VVgum1gtXJtFVnySW4kbDXANID
BKYoTMC77lhz9rPE2rRcXsPz5Ph4Uuz4UNhp8j7PVZczuVLlAvUJob9SamKMJEq9
DTp9p8pR3z16zlkErODaJUI/JoVmNnPx7fZvo+13ZYT5qoCC4af/hDv7BpMBTonC
HVRIquXTPbN1vMGVHY99F53IBYuUKHD7ZtUlFgvhEwTMANF9odGyMVoqTJFvqqbW
qdWHlrVzesLBrAPj6EfksCrRNePMYpZJotVcmT9WxODE5SdUSQcMM4lB+xs5X/1n
fLsbgTB2w0bUTYEmWjFPoqg6sIy1zIMqYoC458r68fkesDy+aBAnr4+QuRn72DeB
EMUA3duWqivbWDE5QmYNzc8S8gj3HZw+4DGhbCtY3imxNUniM1AkLK/0+0v945tb
RStuAudSob1FkHICf49KRj2SAyprYAKbWxe8hWMUD7XU9vuA/Q3th8/xnxDFzDUp
hO9MGLBhWwqQ8BkRfWZMP+GIcRQCaelwwVuaJk2wcr8PuR/lpNGNOfvZS2Ss5893
iHOJ1mW94LiocvuwCCOVBGEtl/timMCvqwVVYBOZYCD9pX5Vw03apwgP8c79i6GC
cvpr+Ht8gxj1vuHhlE1BapAwwuvvZCjI7cVXi6lf4RnFo6fYdbxtGWCKSuWnWPQK
QpjDUSXT3NoaFeDsQNBkIsNB9rvZhRKazb/BdrvVZ7pdk/w+2o0qGCJZahz7xpvv
PzEAUl2fcUpa/BT2zSMFCFyrogh/BXzApJRRsOhZvwSkVz7dQg86C0ScZI7GpjIh
VEuCQjuYngczsXx3iPGL9wSf0o/2iHwlScQKWua9mdMUy6YMVQEz1+BKCSpM4+C7
7PNge2p3a3ipwT33xClYRfdkBo9KebfMvHP2WPXHgSRhQ/g5pU1ATdMI1XGCK0Fm
xtbQGPyETQuwCLjr5x80oYtpW613+3e/i6sm3h3g5zdHTixKiKyfRy0Miypuy6Mo
zzyV71fl8/QIKvLwIUHyzjVCz9JVVb6//ckquaOBg8arWofkO5itGdQFYhmo1rFS
H2h39uKtc7VAeGyfIGDajRfx3D0sdD2DdxagpQAVtD6enDc1NAm4phcw9TUdK4+p
gDfg/ofCbfPP52BHePzCNRct4LfAG1Rd/DGkOAmKnAGXAys719m5yq1buJbQ6/Zi
0ox+UAOkblrhqrFVyuMaks68bWMhelgJXXvltRq7iUA7xCTNiIKZmaj52o73bq+M
BLd3cW+QTfezhi57TcJosHABvdbb2MjU52Gvg1aSZ3cgfgU9OKNgz47g5cjFL57h
77cm5e8z/OyzEq2xoe9xUvf1vJ4zIBgx+mSMnSXwwt01wr/J4S2zAt3LlQiBEaVH
pckaUu7j+i5xhwbr0TuY2Kyn2bHuaUdhdhK0dZKqV8Av9QHxEh2CW7upXjAybvps
kOmPHw7hzpWTyqB239O0OTyQZsPchxN+xqo7WaeztAoLGqXwS8Nwcb8Au2+Y6tPr
t8TQ3Sfz3EvsfBQDJMj1sVdPriFC/QuvLNKLMlkw95ewhnhzlIQbznBa/A1mEd9Q
xX+R2zVu7uPRbEZUe2KLH7Ppnh+9z+4xKj+wOEGJDAvT/qLuBWxQC4yeRBHM5jjc
hi7+ylv/irWFHwqnJLh2DSLV9F4PZgPQXt0KuP9/j0NsGPb/5gUwr9gw0Snis5pz
40vWXZ2z6RkOjE/zdZacnQPIwkqSYesRelFzWEmVFzjfqNO3/AufhwyLwvjvtVLR
5K2Tep3yaoVRRWTlRT6hx65uIUxBkpE4T9oj4k3viDOaLwxbZ1SLpzrEMPel0Aoi
RFnY+EElXI3WsODXyH/qH+/IUoy+1Ewe0yTENibjOb7F3ihN2I4BWkwqT4UxKrEE
gEQvad2p51w/YHjlUXjoP5IfUk7UrBty+USe8zZDpgHErTgStc1CCGlcuviXj1aS
+305k12TzouNNSmy0jpVU7/JyYUMZWU0+2rcFtE5Jbkm16h3gAhUwm8EWY0ftUWO
E6vBFEUmHLnegAV7AJV5YF0q7DTlo9fCaw+fa2V54Atr+YINt71vhXaKxPXUBNZN
98iFRjEXYkBJ/TNO6XLXPqz10Eg5n0qpiKR9uTwZFR01AMYiId9RV+yE6YygOBKE
6Cf46i4+kp0DR4pe51j75pk1e6/johyLqOKNdyCIaCRQb+OcMonhUC70QYuRGIHT
etsFcDzG0LbOUSDjtZCv1yxiGuCXxObmjoyClbxd3iQT72B9Tz9LLv8Wk+3nBA5x
xeP+mYNG9PXa9XrN1Rniwdt9gEwP1rx/ADsLxgprQyLIGFiLUxqpfa7cv8UNLlw5
AU7aFdbgwN6Q1B4DnmJb0tyZgCTIWMCZp4iPJFrlLyXM36VqWjoZgEFtU7OMORoz
T/TAE0eq4iNzOzJJwbjLyAxkJpM0nwF0j2tqtq8aPj5RavZZqoqURBsaON9oE7eP
HGdDQBwq1PlEr1chc52vH6pPDxgiLn/fELRhJQxLeDGwnlxXtIKr3spYXpSLaDT9
2YGHS3VG8fxNgQm6g4hCde0+Coe0Ib6+oAa3FG1yXPdhO1gXVes8twKtTzRJvYnz
iyHzlDRGHr2CqMx+/COKXChjXRVqt/AWA3xokLQ/G8H8j6JJN7oIt8PVemAzB47/
92YpON08FTp8fyqOvcarux+VYFqnlmMCYXuGb9iuzRwi3uOYUL8G/dUfyXeuQ472
xODpW+PfWhXTw5RAC6ai5LeaQS7NjxPDMw6QF4ZCp32utjapqsidkr6zk5tj4iNH
uBJ6AnYvxDMpBF/binkpH5NEUbEV8La2klM08G1LMQN/EbykumBPRaxpOt/qmEjT
NNLm4lBiond3+De+we+RgBf0jYsgmEvg8gqmQAZDdPcOaOi/by/3IhXvz85KemTt
PLI6O9mBwvv6DkDkT3hngdekcf8foF3ky6n4cqXWOlbSFBlemr0xVad+PouEH4BF
y6bnQDciitsHeux+aGesRxt3ldpxRiHULeUmXCrz8N5Ds6ecC6QyOL7biGNmXOFk
0bIO15xTX6fY+u/0U8C0L9Y6xdimOxFl8ViE/2SSEFwCcl2asT+rizNBAFVM+C0l
Zz1DaA3Tg+0UJ/q2UStR8vFRBy7of+8YNcJLS0C36JN5wQlmgul8R7uAhgLVjSyR
uRfTDjaMy5ikcNn1cdm+3LJgu4DOIlNabSdRDSB/DRrMuMB7UjNpL7cUE3+KfNlx
Z4aNexynI2XXvGVVr7jojziz3LboXaP7AyA9gOhxSrA2xQP/FTH8oCQrcab7WtN6
rvgXzm8DflAN5WS7UH7/ImdN14UTDpV6xeet1j4odfZf6LMYN3s3FDEHfi4yEP5z
NDPTlJD8KJIY4YI+X0JDv9H+2dOQBoXpMQqD0Sn+N4sZlLacJIFh+UfpDyg0Xkca
Dy6DUHQ6erszmzxj0xruGZT51t4tufHky936WfP/+8esP5K0vSRr4woBJ4NNq2F3
Aj/9tyYBR8xZ8XT20PrdCeWhK0JUApcInW53mnrDYFlofpLaysd+7RfB41FoAa8w
UmTWa5bvTOgslIXY9M2eIbJ4R/g62o7lxDOpgstHO4vwondDm9d6RurDDUvnKgNU
Vhv7J3UFmaNbOobfLbigP+RsVBXMMK5xzYtujqzG4hmkrK6DUZhuWT7RAJrsRb3e
9fYb2mfAd4Z5nZH2JT/hdc8qGEFYvyjm9l19EWLTQBRd1cpTet0yz8wgibK0OIfq
MV1uRmGXUvxZbQtDgDxMbIg6i/n9mmXukXyHEDoaK+isia1TBQk5PEq+sFjbmO5s
GC0nI2XGX7eNnNaCDv8B+HQ2KLYRTpjAsisy6saW0hHjNypap5zh7MVqhwonKDZo
2he6gymrW4ZOYjGAaOqtcbtGqrhgyGfnci4m/VZgCe6EBiCoW/FWNa3fpwJ6raYZ
+9oNpbyDGOrEV1Zq1lVGZhY3cR6UJ0Fw2KOm+I5kabA9QGjVp1FcjKK84bx8ox0k
yJ40aQ8N0fzqgi7zOTQQUbIF0jT/3L1O31TNp6RQ4PJYAA2fied/pIFSwV80Maaq
H6IdKoXYc1QrNuHr8jW6DkVt7GxSfigfIbHkVk1IYGD+suFNbW8ub+6/pdPMc+Ek
5xpmnRC0Wx9ijkcP0dCnkDrLE7L4VKA7a+/1qno2QtzrhgJuL2HsX4qcyNZm2eij
U0tF12jNMeLCrDXlZG8L07fxwwIyg4jzKjJXKurCw+5MQOcM8UyyCBW/EdEGoRfE
1q+eqmBk/VCjcdM0oCxUnJuXU8ib3Ak66/Q/ovMw7sa3Cmp+/ZOdEqRQIhtju/K/
3eViNpnNjxNR+ojJNaDvz5c1aMHlG7IVRp1hNWiez/BDr140FxfbY8wIJm7OL1gY
VVcpHh5W6Ei4vMq1HT8Id2VZzN14fmrEHVTTZVNjhkYyEO1Szzy/d6ARbVZfNXne
ckYMzuHn57aMuChBXVZnhqx9Xy3k8qBDweWdWNSnykpL/F2u2GMb0AZfu3p+naYY
Dk6OfsDYqSulLbrXdu9YJGp+SO51F/LE1zY+DgheRsUk2jSasC+B9lkMJXV60Cer
6lBjXq789ylCOjDaGf7TmzxuJc3D8aWuCkGI4ltBwR3L207j/ONSiLeb4IPsZXTa
jyv3ZXn2SbTGOIUuVZYvrUDaT4CNB2rpPYS7cSWKg8pepTM/7yxfHuhJ9clWpFU3
So84JpVRxCMnQuOU+23ks9vidUxXsix/s+OchKA19uFhoghl4gImFDdj2LrkmILY
iaW6J7cchzYRJALD9HY/RslMzznZ4Jv8R4pzMBkaZCnMrEvhcWyfCafJ+E0L9DSW
daSw0VGxzQ3S8BzYBgG4U3+7JWbA7wxaonvasMAl7zywwx+iIG5OjQitCe0WksR1
k2gVs4/NR7E2+yB9zl/7iWhu6JTluNpmwb2goDbW2c79T79RSrV9rePB1EJGEjx2
PIOdihXAUDqiYx63lE67hvrNyQkVUqjBv6XUmd9jAx712RptRb+85XfBcLRQt74e
LS8oK7vh+zFt9U7cV+DV4DqrqVJSFP0Pjqi5IOgXNK0wu/fTdqmU84AY9XlzF/Zx
5zI8zgi45orgasWg1Dy+S4zp/0p6cTz9suPG/XLg90ZAUrKn7U8eq03uIw4Ih5x4
oUaDRYMvfLHkkh2AlYeVaIbL+GoV8UgWkjUnny/ZSE4BAqFcyGDMXg8r4nk6u02S
meGJtRwwtba/l+MHPJP/cvFvyhf6pqFZSdOAGlbK81cBUbdjif3sZnbbnksLDlEp
Y8TNtB/AjKqvzO4KwnmjcIr2SkSDf7Bj511R/E7KqRQ7AR8uh16SxbM0SDgYSi6+
mA4NoEizx8A6UKd9cmOrR2wUxwfUNGxZKKu5KXIBbo9a1Js/h4cu5hvVYNDxrWik
zlfanM2RHhGkICyL89ecEe56Ok0Aw1xibNufrQFtCCC4gOh8zU+S+xx8XEcE9fsn
6GJAJdTg+JXsK9JgJ7rkMDOLdQKcrpT86+vhHTtSUIDbRF56jJcHbYn8oBNKm8pt
j6wJU48McdDQHJqVIAf6Luhp0U5oLXp6q83Nl7yujPUhh9prLLm6r8UWi80PDVyX
FzH6JgzfMGpHJaKVR1Jp2m0+O8W91m1+yHwHIKo2gG60L1QR8GhsRgvl1Ch5Ftan
3GHEmCvSK2Ma6sqoPqCEVono38QOaW41Kh1RcKwf8Ko3b/g3J+yz6O7GKNrxY77z
EKV8EJOUeSyPVy7HGpnCZ0wcbfNVBjkffAXA86eAPNhHr4LORU/jzNK5+6nTPkHz
HLa5r/Z5utI8GepMKH/xX/+gssvpMT9g92+tVYoz8XweS1duuH6ME7AIepQsgSpU
1b84qygcgo3zx/ETMCeAWptlKgG8Nj6xHloQEE5xd17fZZyU3yMVJUsBTuNO5ifM
GcH1dP9pBhHOY+snOqGpXXiLP8x6G7+EP24nCpMlMfiGYYSQ699jBDj7yGmWQoyJ
cdEFZkSH8YTPFw0OOIivMb7tbWQXNCazLkhheRGlWv+PNRfIW74Ljc0iUnaRets5
5E7mj4HWBS2P78Oc/LFC9ypnvYgqGI3nI7O5aSMov9cgLC7xXvyTd9hX48LKzzjr
9kXVSB0uqA5m5gyoUmo9tT5LyxrFDWBkJ6n0gbEvuDIPXmNy5FcdrNa75WTFnIP6
tKcKV5rogxpp5SGfOrP/H4xtPyeCFmToVZu25DVz2ozhnm/5DqtLZEBtdUwStEJY
OaUDVC4h5pu0oYxH327rd35wr22E2/yF5n1JfoHJ3wEmPQZA3iBcu8gHb3T0VWxV
MEdsH6lEyUaixPAsP5FOPqIVHkwNMqAhHKMUU633BbLZGpwZbEcj1ki0c19BrwDu
1B2adxB0JR0JtqKgD2vVbkcsm7RfbIVSKKFDE9t23idibzE+1xRFOTTkQ9bM//uS
WgKlPVsCtK3DYWWdooJhd7fk49dNpBSNo3+8p/yLPiOBuLyZ22NcdC61uY0bR8XV
6Un/fqaeTSEkBmY+/D4TEH6R5wXIbJqEweY6d09f26a+8LyEf0hURqn6dIwGSI1y
W0XwSZW+txZTtDcXBq3qV9sIwa8g4ZQ6oKqSN48i/WWX9ztW8+EagGdMr0LRmux7
Vq6TPKVYMOf17HREUe81vx/ia2vfKVb/OLprFJbI4dasNNPlOQhdr/OmESauruaN
c4bPmTjR4MFNU7RRwnU+ECO2UB11NfsHzGPpVEc8PZJogD8RUuop7EtBwYm2YC7D
PrfiPIorcoXIerAzYic8nCmt9NimIoNvZf6sJICEY78LQAaaU7yTnXZKZmLSlHth
yqBHYEiHQtNlGKIbXQnr2pNMUMNs7RUXJ7t5Bhd0Xz40HRBfUY2QBhMIA3CFTjSw
J6Nole72ewE2r3mVtK+aHaKZwN7YquQVwABfVqfmZD+fI2nSEUJCNTR0qZcKuaOF
1YnDppKXpjzVO7BvMlKUWsIS3S7T1Ro6KvMA1+mUQbIDcUC/Ncwy3MBof93AjhSO
3cv+J+SWR+VJzTV3Nbuaz0qJhYXwymaEfrwLllkKXayfTpnfI8Sk5/C/2BmM1Frg
GzzOn8ToCJbYr4kf7xs4B6B+ilQikV/6L90WmnRZxsr3I0R7FrnhneKXqo6M0hEW
SAqUXHgpGivntKd3BuLqZFVFR7yTl1FTm/WI3MJtbbWiHIRkH8rj4JjPgsSvr/++
l1zbxMZ9UdWXNLpxpOVmZ9/K29thCgRhWkakvOEdupZuFDBg/NP7OsnXSJOQufg6
75ogjkmHotQA7IC9LtZqLkRWD0tL9pVeaiXaAa6mID7tZMXkg/NcRN5dLiWbqS5m
awINh3hpfInbndZGF+BB2yNNNouSzYS537vN4OSmco15JcooZoQraN0k1EDVL4UF
Rqdfr/s+g1fVfsHLtXDYprg7E6uo+aDMlpV8p4p/0RGmyp9FGgHUMTqAgBL16Nlt
kKPixJ5olBoICT5FysiWiu4zPlL0KWrJnAxD45ArL35b0wZlxHx7vRgoZGX7Kv6F
7iuzepgxd8dvY+vXPYyIyUQOMA6AQvMVxYt7nQ5DbmAHi6QKtYHNQzskI4caeFPW
54H1KfnT4lEx6Aw9hpckBM5fipI8jqylY9BduGvc854v00LjmQ3WdARHjMd4gGcc
lpnQmpKQsQbj8l6DGO8Av97GXl/Gd2sRvwgnlLmWHHIE700gDpG3UPiq7U9WIyXd
TjoEkjz24poxwAyyQ/IxP4Jj2byRKYs+5Wj7XEdgWQVQ9LxCuYrCpCN4r/K+XRt5
gNnI9XJITf5bbttjM5nL/F1a8cH8P18X+v3Wva8k+OW40p8YXnOL76sH3FC6KIA+
w/M8037q8ZWF3bG2ttBFE3LsVKcEp9Vjr8xofeSmJNfutlwEK2+1NwRFR18uISuH
WskTbxk2ERU1OMwp3ZSUizxZWV/QBhToq4Lx8ogN8+FiBRMCoKVUD2OS7PphaATm
UTHOqeXusRmWw/qDlV3XXb4TrMDxYI+anIRoMKXMI9IblME5oXTPV3zkYAxGG3ac
RClImSue0GRJ3+++C3Vj+JEC8wjso4yrCt9WqzORmGATq0P9ffQz+rlVm/rkc79z
2YvZ35LMimKZHCgeGEMShTtiydFEfDXCn9Oq5gZ1uJWK86hrh0e2MmSu5D8wcPBO
rR+WClxK+2pAkHMcGHdzqNOWHywnNQ8BjTjV7Z8MCwK2pOwBKhCMnm44l8GkCRef
XQoXFJUA0o6Tg51jP3aT+rgH+E1ZeWaqGPqivujRQvZQKr5AdbmEKIBogG8lRkfj
AxjhHpUCYeprbNNmzeNKHF4ssjUk8z2TLngX+izUL5JYtFBdyePWsG+aZy/BYR2f
CPTNowEKLZYYoGHCCqMgB7XQghtYkWUMVunBsH7RqFgX5c4BqkP3RUt0sdMtDvtd
cNIrIaSA5fK7jpHKJWhtU5s1kBrz0pAFcvFVdrXUFUzUrj1nInlS1og6lokhICt0
jjQGrobJ5SoQL3ZsIcWYUO7R2vXzahu5CVz8A6mIH/ovI877+0/1GI8OI2PE5d3V
I39Vw6dvowxoxexc6rLvDZxhtslRkGXISmbndekst1Y6oH2Eb3osIqEWPLIqF0vc
fMk3OLs+ImXWol2mPsdMFywse/Gpcm00U7P7nLoWhqF2IL+2t5jiis1lwaM/kYyK
yNdASsVsDp9de7JOGZibczTKrtd+YE4MMpYIoh/PB1uZRsiZ+T/Ix/LgstBqx7EK
MGiEERLqT0bQX3B4x9fkdWYdvDjyfnrMzG7FTQhY+vZ4GO89yrtKWhDD/76oi9IW
wsc8HAFjcJ2/CRnmO0IUl9X1Jrv54Pz/pipqljF7F6lq/z182W19JaLs9nVHWpJf
D26Yr3xdR26yPZzonaZ4MSM+M3LrL61NDmXAWdQvQ1oJziB0ujg1RKGL6CF+9sNG
C6SbyR27zl9WD1jbIdgDAVhOg2O7IaggI4DqgLIKFo+mL+MeX/vTYk+Li+P2lrZ6
2B8OaRjyr8gHAB9gs3dAjNJCMb/RW1uayEg0UpSMuAgaa8BPn+l4vOhfC/gU7EmB
y87x2OSizno1CunUq+MAbZtAvreHZ0gyemxrw/sT3FlGgFJ1zzT4iBvHa75EWgtx
6h6Z0eA42G0e+r8V6cw4bcQb2aqsgwaK6ej2qdUYBUEPG+5FQ2l3k880lyflxo/7
a64flLHpncyznjxfxtv96BbQJQwgE1CEwsoTA97aV/mi74DpK+8YB07eyHD5yKGg
N6bOzaQV/nbAbxNXRUPIRUjxE4xsKilaAM1DKPOWVDn8+aVYY8ICNVPMvxTK6wm1
qVOI00VkOJd0rqACFlH29IqghrA1qc3ejXeM0/7wmATfjpAuzaSVtfpGVvcwDF0o
42B7keNMxFt8fXfOiiqKr2D20IGcFaOThgMhOs2PJs5w9KoaV7d31NO7UmW+RjJj
BemIEUWL4cQLy9MnVwBLikcYXIYI55CQFd3mGJI67dmqqm5sRNh7Tm/9J5CN0v7q
8h1Bd6BdtDfjAC7tazLuoW7sVac5V2iWEYi021kF+oQfTj480LE3y/W6Y48yS0u3
fBd8rkDp6WO4kA+UepWI5wYMfW+io6ugXqkgLykROD/ZJXKnuJBZEQ49A32p2MO6
6f6+bPgt5JAYugk6Q/o5gFXdF5hLbGOd+mjQViO+fR7tC2T5l9u/lFUtfq/Yy21D
8y0iAaL+qmKAtX+4FhdYqZ2iNHo3JxcqiPQYrJ4CF5u90nDWuMi4+BuL27R7TGDd
062106sBkr2dBVjjD5KjjiIHTWVQFSq4vkeQO4wab6GoJLZBFYR6dWQyNC6EXVZt
BmbeGB+SbmFytgrNsDJ/mKQAWOy6lWm3R00Fi/abzK5uTFReRuOlRpUqmWxe7liL
Nr8Rtx2pgxLErhn3ciOhER1t+Etbj+9Jd1LoXCQlgPVHicFT/9WRCq+nhJOd0Cpn
XZNck8SMoz5lmeHOuQuvLzTsgajXJDBvw6sguhrcgE8ess16dyXLr3d/yILpmxWO
s2ATs2z3YSmGZF6tyb7f5rV6VVTvrf2OqlXccw3/li4uOWu0rzVHbx6SlYV8Ywa2
8S4k25kN1GzIT+hT4Qheg3vI1TbmedrMy+h77EqblFo2BegrWVLWdFvWDyDcKwSk
vU+FkQBiCzVfmzDI4Qal6sCN2bz/DIWXQjO4EbQkkeJW4GoH9z3Z0tMRyiUwr+1S
jgi8pisJrd3jf3CCwp7FinNynQWivsd8rv+Ibi0tn6Db5+kZMz0jF4yz9AlHxkTN
WBgfL93fQHHiv4qWcR3uqmuiLSAZAva+QqIUjD3mEwSc2JwP7+2W86Vc+GxJ3udT
2Z8+/K/ZEnf3II9M2bMdOLDGdv8JfP5APV5/FeqBsc/k6bI0YBj4i5dEh3yZHjBN
KbnrmRukS1Sv7jM8WC2RIgMCVW8Nd9FkPd9Iy6OJ+cVUMT2vddachtH7kky4Riiq
M5y2rkHjIBGQBYyiXzgjJ1Rrpn9VUGFUjOK8boDdwSTDApXsW7nVdFwvnVIA2edv
O83FJ5kWSGIhwqyPK0/oGMLHQT/P9VAw9tKeBzCnFviE2w9I8bGLX6tS7XIgpLkw
mwsx0l5RqMiAzGZBzN0+gQWScO8nP11JopIKfJq2Kl/oYa+Ogydc0+pqIKsOOBpD
MdyItUS8XFtGeUjS8TA4P//JI3cdFDXRr9Bt/uMJoZ/qgUizNY/sAHN45NyZu5CQ
n1lYej3o/J//PBk30RmJs0CvakhY7JEA1sabxYQg49fDzuEkQIe926i2SVKI+u8+
y1xqkR+FyM8kNvsdANNfY5TEKSIA1bAR+lIE9hghDoQ+yWpPSciQbAPbdkDwp7zs
+F6Vc31C98twn3OAddDvGKUY7/ik6Ksc/z3Aia50WTxgJwb/2iUgxn+9KgNRMN32
+Rd9htYw8++3KjVqro6vv489ljIak7gHgGAPqCySTl+twc3dI+6dETmHtJpo+UWU
Y2vz4NQQtOAvwaiwYv8cFvfHRNRb8nfUa71f1a/2pS+p/GOFIvquZ+3iiVmsyTu6
YEcSaMBWDWnVhuAixc1Fd9+Eqk+frKUwPcx5nGXOqbibSnYNR1XGcaH2wcJ9mMuq
1exCx9CxtqVYQRuUIM+d10p5LzaON7rutMiliPJVAYTUKfooSsbe80czZmPmk6Ci
9n1/uVtRFBXjska9wW2rtI6zcD7d/VE5phmxmnjiDtngZN9Sz7eoXhNDu+GOGFiD
i3W1X6LtnsknkCEm1gljP0s2N2r5TOSrn8s4q7oYwogj4TljR0+1IT1Q6PNv4AdY
N3v/5fJAojtRV5LtSOYFyp/xNOKhAt6GpmY8/gXjquYL9cfkXf2pN9VloRl6Ip2p
WUeQGCgDD1N4TB/9McSxEQkD9KtcNVkNhPZOBZpzTXKq0EjDBJhp+4iB5E9Hml79
KGkB2xnh+79YyMw41XI6KYcxnt/4PLu/3k7uN8fA8PgrIGQ1KgAHQtTpXxSeXmU5
IGtVuA6qcP3YfUMN5K+xGko04ZSYDxChsN1qpScQMWGv7C2zrZVIMpTtwuu+VA7z
cNJOZ1Rx/nQx4V57UxauiOvpROpI34XaXD3bZ+nrv9+zdu43BRFOcR1p2ohbDU8E
XtEmbirBmr7ERrh7yJ9k5YE+7veT3n9sppHXF7wlyFCAJ8CHqrk9RHuuERz6YB5t
N3FGU8CcclFdryhcNb773U4vTD8xROTklEza6UmLJvpPXZaLAdIrgDVgGerrrBk6
RI7EfUGu7poiJxa/+keJF4eusF2olnaEyzG+dPT6lhMBcmzO+vQvSVVQha642498
/RsWMVOXthSRG4NbGDxd2fPulh968UfIC2ZX18G50hukwcQk0bi1FN195AxwkrPZ
z820wZ9aKsKl3A5eN8LoyJXKmjuj8lOCKDvTrfhBcZQ7eGgj8R1494IMOgqXwrWR
U1H1i0UNo2/gA6QGjDJ0yNEhVfdPKgHeajMOad/q1oRVId2Y6e/b2grfYhY3wYa8
oesN2ds/TbWv82GTXxTjTmCW+3Zizu1tOfmTrFDAEbbG4egWYx27oZoG+F1gxDkN
Jzr/PPEOAfUKp2LgkLz3+SwrLz/kmpMzEZd5SxMd5wJgv/g44A1fkbWCMulO3NQ6
onZjy3KQnkvAGatzPmAoTnmT3nDVT5ed/JjoS3j26wb0z63GElExnSobsPE7bkoa
pYnZm/9Tia5vd0IJe0SjWmuxIXwEJunN+7UZkid3QCTCVlorm04MnFL6ZHnnvHOU
mVIaBKgl+YHpUs5e4Z6wQKNxEUGhJGPTRJtOHckhnEB4GWzvme7WUjav8h+jApUE
7o0vBK3Li1ExXpND/N3QvdupswQuiXa1FGKG9vPmLSViEpMY5djAEJy649M5pQ+3
Jo3s0qKz4e6BcyWMZ2CNSyoam7Hg2rKP/LDFnAgVEQpKB77QgktQbaHXlE4xJ91s
Cj2uARkTyBx414krfrX6JER+vkuViBp20FsLQTPG2Ac7VEWOhrLhRtxTZGkQ91I5
ZmxPAp7Sb3FpGnU0M5wkpYlNJ7RO08d6Jjbmze4vOQcwWsyPt8ANE8kSrnktRjKV
YIWfnzBFY52p29bi4eBzmPqzGWauVyk2x9+YD1BoOS6m+mifO4FkLpjO4uNKQ30W
y0KdGD9ZS26J12+KOamyL3Dwlji0ry1TngCnfnRifbf6EufW/CKwipkgIhyTwAhV
4i281o+g8oZbR8EWhtwOCb+knvwBArf8nr0ygoIDlie1UeVQMfSnVF6BLFRg+/xN
JVRd5aidy+tGa/qdSUmkPq9lwCPWx1RSYDxVaIe7A6X+ZGK1RC97HKXeKWhX4O0T
PRDsiby5N3Wwtv6iF0eBYMh57AbxC86FNZOkhFNYdZ6MJUcfoeI1KTjJbX0sjsZ9
c16XPItiYSUXrV/UfgAxGTgm2MBo7wUeQU2MMljT/G0DxJYUaGpS5V+BZhbAOZfj
x32e+LA0Eas3vT+/zvoJ6zmIjXvCBd5hCPrExFdYUoqJJFBJwUQ54ZzRXALB54yA
/bcAeIVZyaRjFk080EXq0jaSSYMCOR4wtpEHR8VnTGNCDlrrnIliYdoJrbZrOaas
INYs8CRO67LCSHsqn8kpMtt9+CkinbHECDGRS2SBsPnSP/mKJUfXbajDxNcQzE6V
nemdgI8UY/FuTdeKIlMEu6dV/NxPXXaLABClhMGOE/KSkerfrqO/ku6Do3gpCuFS
xlCKeOT/qJxHJmiziihA78VChlvSXMM714UCJgF16znaoHvpVQjYtNSGsVw5OD3e
dWmI2rWCI0SvMYa/o717AcHVlW9WKgM4B+B2OomYNugoyr7EIfLx/xLl9qu7nXZZ
VVtCotVFH8QSeL4PdtI9QfNeSk7vv5srppBG0ueGEUTJcvY8WPWxXNRZvocOan5e
9eoPhZD55PF8Dm3+O0BAvMpCMkjaqjsGPiK+dUi5Joumg9HgeqoFQNDPCqxLuUlc
+E15c1WURo0waUOb6KT7QpWgrF1r7kNmFWmBa+V1Hy8Sxpgi7cn3QAFTwV9l6eWs
Wbg01JIvCjWsXPAP3V4ASq7hRrkzsM9X0XoHIKKmLEZGHA58a0wjops2XLd2uaAR
vQTbH6OwJc9yX79EBkFvMTwQt0rr2hMwb3TqDXcZYU4yvaPQxTRNzIFYR1935h9m
CkO9GH24aaFTNygy6qPb7aKhXuhcWGi/5dnunWDtuz1gf2BZWNfch/H1fegt2pgt
YP/c2u0pK1Af+eWhw4dHsnFSjTYQzrBbE+E6Xy8l8PNCXdRrzauMFQpHVCtwibAr
ePOygGlCYJ6k4K55dWOTUV5GR8dp+y/5Ik00VXIdzXkTEIVO+UdYibc9uw0MB5en
MgoUs8+bPWW1FGuuaSMarJKWUJDacISGmzGww+4sCGFqNBSSiT7Xk26ZgII6EsT8
X+zyYmddib0vTDCcWpj+xGlG+JI6n2j/STHNsoqH6zQRKuLHYdsOLW1ZhkynVhKw
LPk8r9uV21+p10J4ANAKNyZyO+Ewi0d1Vs7Kn6xsNYISUYqPzglaePnDFjW6k4qI
uoiqIPjY91h/qRqsAXvhxwWGy1Z71Oy8cps5hZr2GKUkx0hzJ/2S5moHZ5FlXcrK
8cKBuuNieOLPrZrTgurZVYS01/GufAw2zbGETwLgFm9yXTb9ERVuyQZaqr3ZrhN6
lkJfyQAJ7DenRXbRsWyNpQ8zoiIScpDbu+0dybCRz+nXi93Wt8MjQM2oWMIj2N/s
y4AIwrQfefDQDKiGjLl80dF5IxtIvuavklehiZAQmsNGG/s01N/p4IP27w1x6l0U
FE0DWQNk8XnnepOCOyH1L9plFVBqPhMbM1pGGw+FoDVs2pPcZpOjf0a8yA1zCrx2
KzQS9ZUIyX9jiU87IxKxvPg622bWctZRNXOOoxVdAHBKFHSYLp/jCUIkSQmjIbZu
aXwMS+qhgIFHkcERt9Z8ZLcaIJyuGi+przOlhChAfPsPiefTSiFKO9eaIrsXowbY
HCBbJrSHMKH7XNeiXxM96qu5v+Udg9yVktMKKAXFyUcwK8YPFVPvn/ncXl2aIgqs
5rrhb1C3DoZw+4cJeplurfqU6v1v24X3EaxyC3RyxhTD5lOY8aZMcu5/e170nBqz
Rqh6So5MpGV6b3QdJRko+EFwOc8Q8jGgIL4mptzyP0PJ82oLMfpskkVKU9jOgluT
k9FmwJBdl9g9KG4IIZ44+NKuoEkPBO//bZ+gS/RGzNLh8cjmGsSKRkUasc8OGqaw
r7nxybotIy6HybvFYLwti4PX/KXg2+mr+zYFvlMC7+rnsRtiltbE+Cf8KIhYlH8D
2tt9/O5vvpqfuDXMwx1eV7Ybp1IzHEL2Zgfosq989YbHUhdXmBdDBTY8qK6jHvWD
gBRHRhsQ8dSZqmKaGml82AFihKAOCj+5GmVKId+O1nroO1VINaykwpH09xif94jk
Ln3kmJ7QkMUCXw62Gl7wJj3FhNmJYD7ZoUGECEW81AwjnEebUi/UgZUd7PIZe2/L
+HmE0kk4O7mHeHU1WjAZoeLNpSxNRl+XxQStw+TO90b0Q5/Xd2GVwPq9r9aSCA0z
j6O8bM4VJPFyW1RRFKBhDsRO1bv0e22z1Muazv7+Ur8IetVzX2Bpy193kSKAgLyp
aw+W82NBDEp1UWJYaJvjzoCDrHsvlCPmJ32elioumP841qSKyQRU2cgob5CCFDWa
UR3PdhvIV3w7e8P+lx/OBZay/Qm4ardtfA3mvLxu5V7Ky/tc7xQGdESLhOiZRiPJ
y6Yp8qJLiprBCpUesUcL9dGhFy0/ml9jO/aA+GUdNpSDn2ou9LBWYuQjKfrmD07r
cMTBLFW1kCGyuIHpWOF2Hv4X8SB/WUlfra0zLQNVDc5H/K9nEStzsmpFmG03UBwZ
BrFMIjeyqeqw9m/CSSz0Zl+FK1QpQd1So6e7oHT4HBYE5QlGkeG1GwBimm/QkmdS
DX+GJig1rZeWUPhZ4gg4NH/T8FLxN0NWdw9EHlE2R+EeH6WLHotwNU/+2HBEBhjr
LAOUZ6TRixI9nHFhVs/N7iTCpcVe7Uts7b10A4Xbyt8p0cpm8v2qVFkZEl76ZSFL
LXqlRIFamall7PKyWAQ0hnijtUxdW3DUxeX70fTe84BiLm2/vyn/FP182VzZ+FRV
Ji2icCg5mAJpT1Id3d/Wb4N4Ls1ofpv1cFPqlSnSkoBgSye838DfAmf9/DrxCq5+
RpS7qHS2LyPzwq1PyQWJy7e8rGWa9r92KmI9UgB2yexTDhIHL+SMSi5Dw28Bxqs1
fLCLp+CFdru4fUEfTQ+bUEkRLBJQW69ei0v3caEwNpv4rpIgNfF0Sdr5yWWsNJoR
5XllpSnc2g0JmEi8NTDHXhmSqNMkkFClK1qb1SH7+SbUd9ir9etmre169jq/rIpR
A/Tgv1WOpFzOd9JmAZp1cMQD2bQm1Tqia58cmJgCTQl9WCr+0gCD8jPJA0KE1zNP
Tf+OWoZ6OilT04YeSKs8hhedYHcu9EHPSevByKXGVDS8lCxvp7+mhygK8wusP7HI
FzQEVmFaNmqfq7O4a/BaVLnkiRvsWDDupGU2ExZ2upqToQ8ARmi1zs5ZW8ejD+Uh
QR6mni8uIY+kvcd+4uFkab7ATGJsDPW8IauPjzzwMdibnqLYV6WCVUM/EClO9PHB
Fq/oQJXC0C9k+lfPHUffCmWYkee7nsQyzfRpnrfZmRjKq1saiF9YLyGik1tfbtDQ
sTZXTZbxk8KKAQ4I/t3m077L7JIFx6mqvcyMpVLk87q0z318xv5an0S3+MZMvE2d
CiNioN9LNXGc5XMgONS5ktnodqutsUuwM4SWrErW+/Wpxud204rwmhUBWAMhbpLQ
JBHfcsY6HbRb7/LKDC0CCBrFrGbr8pxDQF2OvBDOtU8gy0JCNYydVjdcrQ320LRz
mVodzDwEfzBiJ+ctDwKVxCek58N4F3zgEkQZjjsO7axLLyzNN0+gneBuzvZUXZdb
jWBsivfRDBg5um2dM7nF6w6rjb8oyWlxLXULrw5+UL6uCMUMAb/Qn/x9WMstdr6q
IOZd/b/fX7D+anHvIl0O5je8+8H5rm3vy7aBG3KEvNSjcyecstC/ZPG/BfCDCRIv
6Phl3i4pHnGf4bZrYCZSa8EMy+8si7TSAYversFwCOsP2t4XaC2uB5c+HePaqmH0
JaMt+En5Zn8s2IDGVmFfwMvFeSeI+36n4PEiTdozJesEQdFEuER0U73cTT9MpjZl
fSh1E+6atrCUX6X1STnac7zFsRN8TRj8wJ2fJsg97v2OZgOfgMbeitROyaTZ3GcP
9rngH+3s8C4k3TgrxcJ/us4WSspy3pWOMDqEax6VcRsjW4QMOk3lybimSVwGHww9
Su4mlL3XeczWVXWpL7v4C6OdCGs+Hcl5dWrde0HY30hV0M7LEzxJTg5cCGWiJUmB
Y0QIyAgH9kioSA+doo7pcCLY0jzPCou3BC48ZKmo9QuH8KDdyfwv1XJtK9YLORsg
QTI7sSWXyfWl6ax4lESZtTNNbHJBMyyIOZKYl7rZh+awdY8HhDqKmsmjRf9XaGiF
VykZFjYnIJTjrfiQcHDlfBncbrWJXEiyB9v0iZc3MR8OHicyMncEivNpKNn2T6nm
qJQfknNOvSSlBWDCnFSHR4CrgenVNx+Bjo32kJfgWx8KAQ9TdSqhLt2CJ2ZiYY0T
LNe6rBeOnug8lcAAGwvSDyg8WutQM7Dx5H6d0e4DKaBeE8qiKe7qnwo5Qlfzn/hs
bgmBbzjQjq4O/mVC8rJrDIhi0K0fKl5seFip0TaG8u1NUE6CVlKUXrFeXPEf4qnE
W7xQSf9fKsIedet3Lo/TJVbrX0Vp4KW73ag0m0n85xfJwElKwypCZz+5K/+x5e5+
LJ4kHtNFas2JK00vdmEpMz6MDqG1B3QBbYiZJ6k+1P80ZjdnSZfFSXDQWCcOcol/
SCvF21e6r6I5Rks+oAhHBOhjvDyayY8E0MEiFhvcHD6Eiv1ffkzAQzV7dnYJgzW7
3UIgHGKszOhJkuJtUNhpe97llYkDDQWE64nxIKT2xdzR3NY5bwBAuZPmR0VptRrA
JJ/CgOTnk+ryaZyoWKm/QCfKPM7hbMDskXk6R7Ahbjri4qgjDmy6LIz5tUbAeFkT
SA2aKrtcCTUnDvkPGgE2cA/PvAX+1iSgSSFkP+w7nr6hGt3yE15q6skREdj6Zw0N
JzptySh2MXX6tySDHIFhq/EzxxzV/TqkWoQMWv8Ilrb2w/NNGVLBfacaDw4KgRWg
xwHAuxcQPVW/QpsCchJHLR8j5f+nuMrAQYH48BhNIkGXEURnoQBiFpCcN/Bs+4CI
INlWxNI5JRsqpgeYW21fe3oGnPxRzLEQutX+nL4Cyp8cXwjA0YSqq/6OT0FG/Qks
UMdfZCQEMjBo06lTXhDEN2OC+b6Ub8PeQ0/dyh49uOMubtI6T89DJvAuCN46MVSH
UeJn+Ml7OGEjnRnGCuMiHnZ0PW7D+jFzi/u4U+jHTrKayIsC5spHzxAWso2g5vv7
fX3MYNol9fn/3ePwIJVkzbIuHHBRFzIWANgFchT3lKHeycLFmyZJ9FTOM6O12sn+
ITqmfCr2Ot3YE0D0RuF3gLphMj6YLItdhK4sxZ3Gy6y060IVnElTrdX2xfdasyfM
TtE4I3OIXokDx9WVrCmg960qdTF3chGyaSofQys0Lm0LPVdKtozVhLH2la9xGwE3
8QmKu1laWFojHeqz2jIsBrrxby1noWI98DYuSnDNhTHZWjrqH6u3sXTd4H8sjF2L
qjD8b5w1Uo3UbEicypaT74L0YP3YZEFxWn3KMIzXmbfBtN6WCgRWeXHGl792EVMl
lVct8apqpSxPFiHQxCiU+TWYyD2g7jD7+KsJN8gE2TCLXsdSrWAyOaT5Vd6bY61g
uBgviZ8NaIYaVSfLPulromYVAdcgd6bZdHQxe/uwLUQGIWCfcHbDUljFqdqwbT0/
iviEkTsz5BlfSJWk+37p0QeThU0RZLBjMQSTHGT4hwFjHqAN4+m4kUjFOEYe17Tl
nJ+UUmVLsBbzJ2HulZnsVb9QHdaaOMeH5Hz9jso1NCFcez7TtHHn4vTVIlVwefiU
u6MqvzIzzFCKIUsaH6QkxY+pcDFOBW84HQVVZnEKkSKKPywPAApdMozkd6HPNwod
q+f3l1RyB63G8eLTfhpH85v0aSlRyzzQtyzuwAKaCxzqUIbeCtP7jJ4SCG1QJjIY
R4ICOUYCCaa14RE3uR1wQRxD5VOrGNRpx+ZTZKIfo6IDsYWYgzR52ZCvWgwp2HV2
rHPiDPo25VW1E84K4Eu2aJgDuoBwg0iWEWJgOs+bXfbNT9bNMvCaFVh9tAeAvr5Y
BSkNaXNqa8sTQ+co1IAnwRGtdaa4jEufOqcTwPesm1HTmL1w0RCa6QfkgMaM7VPB
KM2BoJXR9XwNRmACHoAs2KJzyXWUtwjdhkdSzDdqqyDrZNFLfWBnIGVB9ZLrFVxm
zMpoVSXmsDhnU/Vscd5YWNoB5pUH83ukYL8Pyos+dVR1h0OWod0eLQ2uKlfOUfAL
PoSH7dWu6f7KJk4VRBHOMLZOM5Sx66Ft+YSM+hB8BFDNuaOXnyZA2df0RiTDrryy
D8CotJR76ZGmWO/xcIqFEYRK1H6YtkuZBry/eeDr4rZ+dVCnEG+AMQPP8BOLUtsD
LvREiYjupr8RtfQBcxD52TnwOhzDy9FGpB/gdDhQwdKq0axByXqxhRCfOQWNYnv7
ZLMzk/U2/ylGoLUGuG8ehLrJYvq+I+xuBE5aMqUds6F1j3QJxqQnJVaQ6ZyZAv51
vblTxGRBEZXct3C/uJ62ExPxeoIzE70P57Iskzd8RGSE2w0KDnEDP07ofDI/TLKG
x8YbpYaXxKdSEZxX2qcClDkjS3UIxp6d4AhS92xMJWZxti/5T0alfpcvI9nvcwJ0
iT4Kf4+sKBhnHnaBCarvp4q3Fp98MbQlPkgoRltRIqQQJXJlIMgvLZJS1lNXosBd
Nkkk6izPmnhsH02qqf4lsbnL2TwA83uK7L5y7DJudGTbn7oUc7wArsU8zmgMRw1V
j5Bsh78DI+6KE2eL5jCoadCktCHkBY0yUhDGZARJQeCfDXe6Gb9JxlLz1OFK06b7
adMqzzm90dChPqubM1b3F1LFoOXiFdGsW0pYnhugy0Q5lQCzT0UlhYBLABhJRg0I
l4uVWD15i1XhW2mCWYiC9LH+mls1LdmwAk5KZTKlgRMTVv/ZVWzdq/hBXrSmS4Kv
YydSdxDuyLWwCM648g7Q09vkKQ0dp7+zOc4KNYnLs3PnjklyR5zhmN/nloNFXdyd
PMDM5mG6i2UXKsZB+ZU4R4hbVT0O84oPVjf12XTmXk+Y2KysAK+kx+E0w0+MswRf
/eubbKU6l7ELg8VsM7VbQ5+rYaQVL06+6IcOCVz3qrZwpGs7PDnojCdlLQKCPDGw
PIgoaF3Za4ZPnc1v7YFBKa6toik/7zWhoc+RdokctHDZTw8eCesOm7j36a7x8Tvd
JCBoxFV8/4ouB4T8mcBHSduYAHf4SL3e1rl1iWCzEN/1wxg/xacFUUgHI0RtG70j
iYdxxd/4bIvtVBqVNZ3n+x0kH3nDT39SDaFwJaXdbcdELrOxdjWILJGzDC2kn/Em
YHnyLqgAQA4kESmMx4+LL2/jnTUapjPKu1qvxQzA7edkshgARBSLv0AENKF0kZlw
qScdPLUz2wdyNdS8lftKNYlkW7j28kTBa3zfT3lSYsAsCNlJmPpW5EaPALD4I371
knABNq4Brj59bbpmV+muAcbFVnTHfZ1m24zXzqWENLrX2Ng/wseqejKmvn1nWpal
V+FF2eVGwz1wlb7aA/FAWYPjo/sspNeaeschd30OgIXlVn7ptVETPhmAdDK93njN
SGsEYq37WtTNxp6mD6rKVLF7DMLZHNdT+SeQpjD0h0zMomu9zOdFwmFTo87633Hs
1NVzoQmXpbQMQr3RXetC6Z/uBuiGcD0vDWCp5pXRvUHFVPrfrO5EeLzGjztmNQ1/
YsQx5uWwAUN8uR6B76B/+JHVGhR7FX4Tad6/ADIGD/M3F+nMYriZ1xm6guR39be+
vBcgQEH554MOUn/3rWyL6xJwmzQ9UQh+vX+i3kkKBkaj/sfKvSvQ3WNaYyPm2ztJ
73vLBVjPJbM+rm1SRSqpeeIvW0wOke4Oeub0eKApa36FNWVqDz3yeqIAqCupc5T0
+VqqLibfuOw8uE6bL8dcm2PIiRtCq+5egDYpUeFqlowTx7ZrNTSwpehD0mdhgR7N
ot75nGDjW7DQ0sDdAqSn2dZNw/YniLrz/iPsAIvQiGMaSQ5xpD4CFaqcTK2/fbBW
9cxphdlyAVicRPMQ28B8BAXhRlMMnYeyIp3RIHyVHIXHIC2y9Km3PQKUU/SqiSW1
QdkvCJuJj5HLXo8CTA+jLudyZuoYRS7w8HEAn3IFl34MTomeWdurQJIN7haab5kI
3Jqb1q6P39T2EtZspHp4+rJkdq1qzjY8FVFlpxVelTcl4lNrAhmlAmza4rn9SyWl
QITKrsOuHTbJuU3j0nX3GRwdO820acwQfeLfXPML5RFUdYo+Dv6kFDcpBqE45dnp
7eKUBFp7mxWuJjHpJjvSmvNXvDsbFHPKFkpq+2c92vqM6ZdN+6HiKBqzY8ICu9D8
FTTKDLknexZTtcx1w6SvJ/127BDB/yjqFUoMZhGb+z8DCAW+oMWKXQs2FNUfpx7V
vD0dRZ3E2MzZuioMLMd0ffadBYEruzDJZqJxJgbnZvsADVbNdiLhVJKuGw5XIKnn
gX7Fd0wMy+U/5O5xDwyMBuHayPehPut+EZyeMaylZN0F6h6F3tpjGCcqnUkOeC+M
DP1L0ITYhmRz5mxvV10gQc2+rDqgNLaEeayclx9qt9MBjb36euFd6Q6wn73iukuP
2e6kctGVTuLc4J1KgO6zSjjQTvxAL8JaOtM7/NSq+y90bDfTxq8oh+wKT9HMk60b
OOxhGXAeQZalSAPVoFYlGTD3pAfw6X8wkOz/TLmQd+m//rVtgvb4rPPz0AywCgJd
1YofowfEmxogdqmRg0/FLYQ1dLv0qNKICeLa9d9iaMQN5xcjhzt6rmKMc0up3DJI
Gp8bqwAktnAwBq0Kh4n2bGr05TGAEHl9QbAIER/W5zBDmcATJK34pCNuOUjOO2qG
Yv6ArBmW+vvuROwRYLqF7x74kur9uBnUqZQIP87Lm4QsQMq/bj/6jRr6ar4GNumW
h+wjcxbvT8cEwcxkJ3zbwSniaz+gsk6TjMPxKdPrDevtuNpzJKQVWjKlpYZo5RqW
tbI26ZnKlkOeTnNHzG3iJTCEonTAmZeLPv7NZtRDM9Vw2HMkB1ahNScQftGcDqiW
QOrcLaBITCDkoeF8eOPZ5kOpRlfSK/ykbQqqDNorNuA2NBpW2iI0LYN7P9MOkz5x
UlYm8KGvRIaFs5cIuh00JTDQtSqC6rsQDyg95HNYKmuem90vGniwECINSGns4rEm
fusZDowxPFw3V2XR9VTJ/jtzYJwMuoXNWFuI5oPJw5bB0eJJTIGOEIuZG3ZSg5rN
v6Z9yA2mCWml/Jw2ARkr0pXonUFJiVAliDPolTYiCIPTmpXILmOxotSZyhWMcZKA
blFXaEjmKxb6s6R3zDNZ2wXog/xXtO90sziaB+zB+d+Cc4WoydRTCwE25beJBhce
RQNYcNSbhROfUC+0y7p5wPL1k0PxrrDejXZJbsSjbSNN2cSscDZgH0YJujtp1t2L
ynVwSYfzvG1EOIA3AN+QHc7I1t4ydHKDqTqJWkVFK2XZ2ZJURScilJcG2OkcvYLH
T4BKQUQQc5bByhDcu9KHk7kB4koOtFnXnhGzM9NCWdphJ3zgCPoV8HGQg5hjQQoK
GapEQUOvCrUKoOIZTMWE6ErOUVeNBbNzSSAjxi8/cDvFNXBwF40+ih5rY0xhwkdb
OvMzuJFEet2IwcsI/nS5tiFgILP+qVSeUpfySxqtHcNd3njSu7f94xSU6QPCWddC
iPM/bc5bGW4V0TnNgiYPKXdDv2NV97sE7K+1/qmbaJk+LnyScFDkkApfFlfzuGoH
U/Lkgyg/clpv/tG7epdruqBEnPm0qCEXWIQpb8O0BTjYN54qWfV0QPaGdqBPfScL
JHS5n6dRHOy980qYeOZl1KTDUHsBcSbBoEr0Ds+bPeYMukWJzKoKUAvqIJUc6Wof
p1RUsjyaNkmPc7nk7eO2dhCFwMEhqNLuJYo/spWhcGJhUBms6TGuWaHyQRViGFhZ
CcRWfhUvXlbQGSwX0wM/IBaRSkSS4RHdviVBdqlNyfZikTKbGKUlxVlcHnoaXyjV
CRxV9N9SpeYWo5SUkxe/W/4qLjUT2OWB/0mA6+9MWoBdR4MozUvY57pSLD2yRJKD
wP4DbaRGBI7pIY0GO7XnoiQXxwJhqQhXvy8abNH382yTT4DR7O6i67eOi63fV9be
n9/xqoMzJDxhyhbIKe2hw2SJ083jF4rj6//QQsqehH+LWaxdXZBGsZKuZzpvSRmE
xzo2h/SO7mcnDj34i3ug0lQDIQd29h0A1sGLExyT3SGrUgfvMyHGcWvKWXwLOfl9
Jer1pkFAOU0IqirlQO3UHgnqHzEuveuT4W4pENBL7Xh/O643X+iMGPliNyJnOhQ2
ra6HSAfU1LqjLU4wpoFjGWQmyVil3SWL9dGCrYZq2HCX1S1BqdbwTwBe8qRZe8tR
jHCm+PBDY16ZuD/WnGeSjicwG0OscrydCN6sv1jp1EejcWrYJnqHcDbqCBOUN2C+
/BcQM0i2sEtcjod796108TIMqqyQmua1JY1JE0cbrTMFGYJ149v+rT6qw2E/ry+g
u2HfVWOqf53Qd7zMEFuBQqQu6kltk/sPh4m558Y/G8ZEaXsrO+efVMZa0t8iDoyp
jsImpO5FZYYYNmIPaeNFSJVeEGE6PYZJJ/ucfRlm9jmUFTlb2fkqVP0LrBSpfm8l
K9MuVBRlNCgc9pZ+LqiQn58TquWJPl9zeoBv30gq0qohbq/9G0faD9Ti4b2RT2OY
fN/1zfeVhvuVRVhT+RNTRcfaoAS8c7pNxorGLOHI8+M3I46gftCSYsL9hmdY06G3
1hQohcjxkpBxjJfuuhLQ7R5ZvXIK4/ca8CfUAtzhusV44REOjPxTwqiMXAFsbScp
ZLGc2bL6RP1tXnEYup5Vjs/ipnt7zQIlUUsTQ5lchp1cFKSStg7bG6UXKk7j5yjX
yb6aNa8pq8MnmJOpt5ZAIJM49cDZs5YF4Oj3kZEMubIsExXSNwm3FcVRrYOoK0fQ
fNM3VxDWPsiP/Nrf5qxM6vhTQin6mokmcbqLijYeK8ecmE+nXmi9CzsXn1qZIfcp
7ltjE/npsdrVrp5UZvmuoFFTgOU2R5Bc6IWbxFaPDulC5kqE0V9dy2G/oMpit9Wq
6Ed+bX2R64fvzR+yKFJbHsxKlaKBwKI0wtLLi61VezTIoKasdQp8HQg1QVHIHaK1
aNSCYGfbF8qTcmth+D1d7Wp3dQpDAhMigz5u9AWYfqSvAIOggnWG9o8e9L5Ymfqs
DZf90DDP+/XQoDDAZ9AmxAeO/aBJ9Ayb9nfZvjJeSFhrQH1bNNEYSoc29U45HS0x
wm7CRBZS0sfXuLm4jVFDDR97pJoLR590l40nn2CcZglJz9LOeT9ECxbbLDi3O4ri
rHT84uwcGMdKi/+vMiFIKHY1IHUfN6VlvO3tOhKJ+kHvB0ofznQ8dR9N/R1Oh1fF
62VYrMgEKO8seUr6bvvyjXkYWb0vpxAyarvbwRne7qW61ayI/CoI7AYLrWcSkwuu
iVAaU/YzhFpoF4UBOXAwVpAAbsTLg+VeC7INQquSS6asuOLGhmTi0V85ITW05p1y
DpuqBtUeI6WtSsU7fZ+q+GNYcQpQVurlOMh7KxKH4NJAYuipIsYtMqyinOkTMAWi
/SCSKGyEleHvK9RVW+Fq2rYMinSmJBipNlpHnAD10YV8ELX7gua7FFG9ap+gWq27
BEJcqJE+rLy+KcjYcNZzx4ktGy/ZdnAo0HuTcO1j1kxmx7egwaP0vayUMzTzoxMK
lhOQHlP5lCV+iA1y/EpsDKP5ZZkV1st64WM+zECp27xih4yVWvPKJ3L4wcuNoiFb
g/z17MCicfsiq8fudznSXLtpiOIz7Ct5f+tbN4Tslfx0SbDvys1oueXAqW5bWw96
gTJlYnfVQojwniPoL50FEx0bufA32k3seJ36m4TfPhqEcI7PamYhnO3jtfTZxvtC
M9mp4J43KBQbFXhEya3T9YEPpc5+2r3TAlVrHmsEraRGQGmfTCAWZx+ms3UrM80A
0iZ7HQ8zQ0jJk1FXouG5mucA3BgksBuuLnzI9Wnur9iHlUaw6Ci5NUc9wZTZA+Zq
mgedNR+7Wz9Vxa5oNJxAeMMABXfX8T2KaGdhYFprxyJFVfHrrcGtAtvLYoDmb2/g
vMEl8lOj49M/vFfXnyFYk4AfQaQmJf7eGSVchn+sqptP1zTAcPpduMRhGJzX6+Nu
qwLJGOtodXImx3pvangMs8ByHL+qSz47+cGS+CnzlAvGs0BoIWfudUstUwFrMKiw
Ohcc+/42CvxG6RdGe6NMlOoXp5NQN8jBOH589I+A/hebhBTj0kDUJz8WbRYrP9/U
Mv20Ksg3gcR/U3f6OnQv64IRC14zT2l7OD8f/Cspkk8sZVPvcokltg2GNagJ4N6n
atbOQsvJTK4xHGyuHAY1n8tVVB9WCJsQ9aXspCjdfF/UQE3VVPGsCH3g/ZYUM+3F
8cqb0QS0IxpzyZcAemCFR0/X0PL5VhmLNK2iYn5KrvVm5/3xwFacD5ATUyw2g0tF
DvZCby2JUukNeEYhgFz7MOMNg7jTrZCPfEbkBVBBiy4SEpRMIHPQD7Gx1kFVYry+
ba2g2tBQ65Bq+4+7Kiwd5kPXktLGSNnyaFW7MfZHseisrOqs/rqfqPcW9XB+95dZ
PlavVQEl7A3LES162Y1OcjJOE6tzO4ytECt6hIVuvclOXyqJEAx5U+eHgCXu271V
RBjMKMfmGDzL0U+Y00BzW97b8i3g4JhObtd9IPttCP9rLoHqaAoHAE71uTpVOiK8
Ug8zPFCUuDKQF1KzUGPPX1JFeqtXzNWfGDckDDp3PrRlsLo/3usVoNu9E8v5c3jm
gzvQao0sbHoJiGfakLzbjVU7WurOtF4lEcT0V/x3qJMqCGEwQGVgIreHzJ+VOMyW
R9i7Wc7OlHkjg8gwEBL8+lLeFQyLWO8czQqZgrJEbOIR1rOLOyfiD5LwgjxlDADp
Rcf0rrYzkNr888RCkr0F/cG7dVXP1ZpQhWBu7tA6qoU18xl5cEvBp5YeHFHP434p
Z8a9aOTDMjGY9n2Svt8FsNdN0r70sJ4N0EFeZCfMlSAXbNGfkK/AA9AAtcwZatYl
QQQ9hu5dSPXTQyd+DaM8PC+h3vviu5ykCWN7Z5+ERt5tuSBvTKXBqQ48OX9Rp9zz
h6gv2jE3LQb+c3KuxLLKkp+IXzxAtA4+z96p4AZVvwti8UEpLqrZNVhkbe5ckuSL
oevjiqBhlRGz97gaH3mnDAkgKd7b6BLXCaFefA+cnn6f+tXZZdL8gWOCgBCbf3SM
XnF2YGB9ZA67iRJwAXl2K82ENpkMJXB/AG57FNaUnmSUTR9kE8SfwFH7mYD8KTX3
NFTQERhLy5dJPgaj1MTL/mkuxcoaTrX2TDYaSsS7OHQf+2N66xqUxRT4Ws+FyEUb
+gUDy3Pii8SsCwclpdJE8c6RLgesOBHBYkhGVkvj/N2IllAakFem5/kG0ySvMCjA
2pdLwjj2mM6OwP19eQ/ahlGNEhvrYaJBFYLNHB4nEPIXqTSMTk0r/HDGeufr7b6Z
1snuE+qK0K3IH8R3fdJvVPXDKk5eRn0B/14v+Z0JnQAWSc/0hgnJUUVd8MvSxSM1
AReBMIakG2cYaokTTYIuJjhaFKTlqknT1qyXA2x1V5no8kz+PjpY8gOt2DVlYdZ4
2H1ewVLAyaj2dwip6hVGE5YLbAhP6kXp8iwl0Lr4GCFDavL9w/TNFBwntcoeTHjc
FnKkMmVnK5ApwWQruLsVLn4HZktU3j9wcivTJ7e3wCQQrJcO3P4EhvdWOGC8tWEF
Pb0OyPZNaElMaVzXFl4f6go6Y+1hR7q581ZQRIerA/Gxat+iGx/JtR86wa+3y8/V
oKwSTyf/2bTdHjD5wJW6NG7DpMdYjyxaGMpR1TOGFc39qOLw4gMgKVfHuxHuSrie
pUEUtATN2VPSPFFxkEyPPLnhJvy19B6BS/KQjs+EXTdbbiLjSVzmxl9PJvzyMDao
Zu3sxig4wFYZcHxLe/Ce4rzExxuLk6JNdkHD+0fmbwx0shrv5OkI4nGI04x5hr/9
+b13lc2FtgReWHV/NaHOkTtJgKD2fYd2dchqag1tl/9om8Z/KM8RcVTZtOpv8J9m
kFNbhFhjkSigjy8VeWRADdZiErRAEyi22RoQXJUfUWYgMPAi+Yp11sdY6e6uUn+9
7IzUQsRY9O+4lHn5XDZPtvMJlcANnA//XqvVWbffBdc5KqVDPrDRttXqTDCRFqzR
5/ThUzLLvxQto2vxsUC7JXtAP6enIAxL/l547k7BZPAB6+7TzzxdFwvfKgN6/SbU
UpM810k0k1/+Tr4aa8lh7aNhPYsSECeZIX6/5hEQBdTv2LcgbbDo1LeklsG2Eu8P
hOGuLvjCJh2Va+Npy61JS6XqZJ6fWXAJmIUxht5HPSYXgQqHoPRzz02x0/3r0HfD
w4JJoZ0S6ELPBiTSNNTlUDi3rOR415fC0cwbZhiCNQkMX0dKQnWlKyrOSnoOsh1S
sobFI6mppE0Dg+B+aSaYAKzlackvQESO8jSbG0IdyIG//qiaRcTjj1JKM9dGGXjw
70ARouDsIKqcX+wzqyia1DlABeK6wKLUyFPaIyX8Jy82t+mSeC6Xn9IL3jogHsaS
0tuJYy0LF0SCKcJhwGWw0SD2pLX1/G57K21jtSXHNyEb0oyofsWKz4m5EF30u67d
F+6BIUKnpsX2n3DchHkBc84Xd2FNII08wSpCi7UHapiFHTiAWjh1x/Y78p4t+nNJ
kpIE68buDkEMXHC1/DsgHUowZfW1gty2r33yPU32NFMPew9CVBnXkOneHPly7H/s
wD0F4ZinNboigj73OJgLULf4aq6qu0IJXKE4J/2kXCmKLv87BrYklpryFymyByUJ
Wky+bfgG5CUnPg2lNFQF9J+RNJA06qaIhiXzGYrmzKaSY2OcOjtYpNs9ZKSGaC37
5QHJx/J7bxnMiGxCoTzqAwIFEAi5FmvXsjg6MJKkdXYi9GHksqUxW8MdlyFGbkvV
ce82YQRpnIMxEMY4NLQQD4b/po2jwxPKKfUjNgSSYHGN3u0cTD5I7XsA4Qbp4qol
isDwGo3cyL8PDYaJ7LG9BPbb/GPm+zzyiTFeJKX/PLWIOwV899MJ3Mwa5pX/amgM
DyrfP98MGCBgFWpV9Jn2vBhu3QjrQBzesMotuLeDDAkkqMpJ1wPsjpyVKPgkrBya
RWulEQ4IPeNQtDu8zIkaGlNAtFz0rIEx+i4d7LfpYveF1AXSOqmpUgEOAGsLAqFR
DRBj7TWwRiZnKqFn+SQqdyMAEjGstHKITlWrYJTuQy66cIkzYgNb6aKTDnNFHG7e
I+MRFWIILELodJx8ib4daaw6LfLOu+SVQkYjIG/manZovv+hmfffj3J5GtIKLFla
uSjLvGaKfWTE+0dxxWrLQcOw/OeYvRJXT882bBa+0AtyD1ROdon/dJJ2p4Qb6Cdg
qdklgm/co1yA6prYhenCibXzEND21q5e37lcWujes1yRQECYPOhh/29NzVLNiq2t
30QU5w2Ohuk30EO4q193EfjT1IZ5Zpk/GmSfop4K8yojm8hRFfWRpK98UC/GZ4Po
DB4gEoTg8rVa1Ca+xKFB3Z65hpJPLPkC27a9dLVim4wTc/+bD1x1vDE09TXWj/iY
taSkesvfnjgNOx1kZ8C5uJPjU9yjSu88xYLbO/8+ZlHKNWu5GizGwntIZqss8TK+
q+HlEVYZTjd2HyNg/+MZ8oiKdFw3/jNtZszjsi/3gnLnfoADyv6fzSUGywaxHwW2
wVdlXuNy/ECRHgIUjex58x0eAsiNVkCM3dVRtL8v6mUtTRL6+hompPF9oiwuWQW0
FuiZ5e9zr0UwomB1YPKk/AXRVvaaXzYdSRA7tGi0mBP9zPv3cqq8GN5U8pBl/Sae
xehsqJndNXAsBcXh6DhLKPDbLb+iZVpYjXvf7X4srINoKfycFolXi+cLhLfzU/iD
B3PARLIHmifV4A77TxxWiV6F8E5N39viUYWlYcTECken9WhMoAbIA7nkmC9gOKdb
FP1soBxxgZQuiW5oXZdjjTj7s0Oh0fh+LHpieLSki0eWgJI5aveDCl1CM4Vcydry
z6mfigNQ4CfMX3EZ8P++W6fZ1ZmCKzAuzUax1YAu/O/wTqPT5UxsMlJ9M7Ip0qhr
ywv+MScJ7bjE2bA80VLgS6EO0eO7qOwgc35147lvkQ54CUEoSkpi/9MOH2yzEU7p
QJL76pTioLtfg9MK9YRRs+Cm4mW11DkKckt2O7VlKoailRbZr/hx8SHE5M+5GaVI
WMISRDkODhaUdgie5q22kAS1NORgi3TxveM/LQIjKIsHICzwVD/xw0UIMM68JfGX
ks87Akm+MuWAOnH2e9UIHqn2w7dDHcnDfnOKon8UaXeafcl/kq+vSAwHFMpE+Y2f
p2BrovzH1MURMhP6s1qbwkkuSfJ/T9iljKDSSuoa5Kcd7Agct+NgmWMKCYKAQ2sT
TGa6u3Svai4VwjWh1YizDbXfvOzlD4gtwgqV88oDPbUs1bNNQK86WGasL/ijOMcr
AQM0R8mY3jOpIt8b15yVufl6nrl2hS/gU2MDzjtHQzWYVVzMa+o5O3Q/5u8Ag3Qs
DGtUqmOk0VYE6DUwAphzrTZZ0veiN429uk+E6F3ivYXDAHyIi4HK4htfOAmIRrFP
zhUx3DkrVz9A4kvANmgls0JiCCAcuy3ji+cZE4dXZC0jUq2z1KXNvOQXOwDkONhk
HQtehXsDQuOTJ810exZP4n92CeBomt1L2otU22qLSqjkKmTq2egPssv5dUPj6uBF
jqmQV4GyftX2ZLd0r4/i/YKYZfqYBhADZBpgAEQaa9mrL7PIkOnZPWGy+1J5IF1A
NvV2gqQ6wMKZk3O7H3rdrOTva4NpAQ/A/tKxsusfUIQJJBSh4LDE8lZ8ogdD6w3+
bzv8e+tlUU3v/BtE9Hj2smcPbAtUSnP3SUawCT/bhwCQO504hUK9lvEddNV1Gzbn
X5ZbrmpXfzWKAFT0fIRdCw+/jp+QtyFliGS3JErPxHD336YSlJi2mBzVWqD3Jz+r
bgK2cZPmG/A0KXyib5XQ0Q/A0V3qVB7F9i+foRzR0fwkEnBbnt2ehEGOjmygs2Qk
ckZ8Ixz4oBH/8FuB95Cb27yFTHiP7cD5iTe+BIlegys+abdNGS63bXb+uED5PGEj
N2ga8XxQ4NxBakmC+skGquFz/dxMARlQSGgaIQdwliDfQOaaSMalz9b6bxWJV7Am
SKA1OZq0PBZeOksqsuVHljGDAaFlq+agMEgOc3khFL2jWYNP4JG87zSYyXU/m2t9
kJptkxlEG9/KYFK+KajbIL7yKYQeN+v4Z3vyC3x6LD4b7Qrgj088dz35bMrZJd/+
ClCDSyfj1N4GeAkXgSSdFqtX9pHA6YMQJsdWZ/D6awVPqTg9KtfntP4jg7y1aR1p
Ko6vtw8oPmNK4jR3GkeDihM2BniwRt6M09/whjYdgP+2dXhiF44Nx1Vpv26r09tY
XHjFBaCJGmuaV+Iyt4DfOL23zuAd6awRkcbsqcDgNgGDicaYxCc9Gx61IBONV/t8
izoM5mOx6jQWD0uQN29a5hw7P9J6E3+yWC3YGjTASx7qlg8KrrId1ezMWChDvN2x
wFB/Ep/a/tCSzoJ5RdSzf3VdGjO5sKCGnjysURl4Ef45K/OCTeXHYDIChZUdt3qO
6z5QYeLKXiJk1lybIlFaXPzkYNnpj0wHkR2eX8KCrnr8NDrGyGM9uwsWQoqJuSEL
G5IJ5/wo+0XvlutD1LMajVz+h8ZHJHyKpJ2xXUyRttzCKfcB/t/qd89nT+2AzSAq
p/s/8ZK9crENr7sUnw6Z2x0KaCkLyUuEnoTXNDpjqotYPDZgkrnISYiJxQcJ8LCv
IcacP2WrW7tng8rVVkQ27BhBsMzVA0YYazjnbtV/zVnjD5I/nV5P+rCCI4PDI3kO
G9/DNj2HEY8IPYD2GfxNtDFGrpDeExN4GLaSk3iBwQkaKX2TQ1qTz+h+Vgg7ZjTf
tpkLydmNmUw5MlViR9pAdjpaFyYomIw5kXK9+RLpi8YHLAQs8Q6bS8D+2DIJ0Gvq
kilrfSfYxvRQZ6qokfbJWZK8RsURfsu0WP8fdEhvfzAXkQlQyy4sWMF3uqp/02pg
SUecl860z8T6TxjqoZBHCrN0Zw4TzNVPNP748Iv3Z0GrBNhmeMTdmgAH9zdDCwrn
xGawmS1WmapF47sqC8ouBLaYo83dUDrCsei0fqTt79yG0GQ/IhpoPX/GFtCIx/5u
5GCfBue4aeS4XrmUFhKbfWJwu5LYM8iU5IWLRdYsGBHnEJEehbR4w6z8h8/AkWK3
cEXSPzCReIrNkhTQ0GDUzUI/m7WBTHhevL0IUhOmY3f22T1ZTdeWN5XJI6CeDxNK
BVD01CKOcGyF3Oww2Nk6monDD/Oc/VC0jmHMHzJDJCupoYWcUvxiNzlo9hQJuJNw
A0CqSYMbByVhN4dY6yTfwmznJ77TatlzBxpXdqafPwh2gkFbq6Yd58TJFqh0t3ka
epCxtoZdvOFpacPNa8gqVwqjCCDlceKCbu1evtwOo2HioeKGlV/V/DvMwarTt/vR
RP66uyEP9arBpPIIuDs7KxPWEvvWBUBX/kzJNMTYPzFHJ+GriMzLPJwqn3PtgIjx
VOKfSFElYYk/M/+fQnMRaYDClD6e9Sbfu1p1EpZ9LRWByvIvSIc/sdywNPIJ+Nl6
rEpyMVMot7jQKTvcIUfsTI2NJRAw3I4vEd5A3TLwXh1zbCco91o9KnCkNUZhDcOA
zsCwXdVk1PHJUffI3Uae4Qiq6uU5OkwSirqPi4h4OREnFxA7h/IzFN0rd7625+hR
OjFi8KX84nx+xFCA1YVfEoXXccev8iF6E7skkZ1NaWS83z4MbrsS+X5AUIoln+FJ
YSRSXOTTyS5a8TYSZxlVNnb1hGP8xPhLn5DDzJWF77TEn/326J+kNbyxrHyEudCp
eSkP/pgd8mXpHG3/EFyPb38twrVwgQjHdm4jQmaS79sKeO66c0niAHvXakf6J+VB
ahLoWJ1X0f9f6XIMnQWj4j+Fo9Irq2QOHTD6ddpIeV/0Hw9B6TwEt2b/OcZHk6yJ
REnBac564z/RG3UevcEuSI9FBGL1l5XwE8ibxXzZ5amL8fgrtMvNPe0VGke78TFK
pEgWEJJMl5B7thIYC0/dSoGfb/hYuO8sLTzP53XJ+nuuPRFVVsNpRhQ+T5tuQne2
j3dX6+4/1mPJSZtIzdTWnxcgYuvirq2x4zo6j8b6VKyEAiD5IWsg6tNsu1zwDN8P
cVML3LT1qTADW/fx8kBrURUX+cRXagzlwqOjPEHUzeFZ+qG+DBOn+3X1VR8o2qTM
fg2fg55gt1USDKqEkAFmZJdXq/DjrOijiU+9Ui5ZD4mMUyUmFVwF0EWATYq78ki2
W+sVW1gX5QQvDF5p5H5xlx9XLCe6yzmN+EuU/7baG6NLpx8wE7eiCxcblWcHAAA1
AwzwWP5K/8EK7KxEitKfjH+llNXMmQgY2BtkgxXrbuj8/agdsZEXJYUVkmBNU3ym
L4SCJJ5IcT4kAkelxCv51b2LD9xF71Yqr/yOf9BlcCNvdom8iM0XFbYIgY2LoVFW
vH2QIH7SI2jfPjtvaE5wr10ed9p15J1xV9UtuJw6A9J2/S+GTDFxO34FWQTAigMI
+gz5EgOP/6zyzIIPk1OcuOwOfpwkzuY8z01jANsO/cNqLb2aNv6a25jnpavLe8zZ
Lgz4wkfIepX6UzYBJuGfrt49tn6+tU5wnoJi1Cr7fuQkrTDzbiD55o6O7BctoHrr
C+etixuqB3wfad/dg8EDCh6QHz+QJAhQEA4qDFCTInOW1Bt7b+wAmOrgiwiNe+kH
CfdQN7hz3ubZOZzjmHyRo0nUo2R4S5yu5RTmNGPH8oCa/u7IzcAuNLDeKjndDFCE
bOm/jnoVqzGGGSiwKBObWEh7gL5MGlBzSiuKag8KMFcvNX35A1V1b9e/KmkkPWuv
rS0prxBEpx20IC91CGtBZdylBGFiDMMA4m+hbH/EGes0HasMlGe1Te/DjBlp9tkz
aFC6gk5j8BPcOhYk+AsZhudlQTuQiddAYf1Axp9hQUCmH/1BSkA2JhGeT3qnuFU9
x/nZnIln7y6dP4ZDmtm3dh357kPtAkYgONtgtsE/1yenvONQAKKlu3I+/ThSfWi/
EWXum1HPy7s8wUFH8ZfRnBO9a8PEWtL0nDL/43mMRIbUq9u7bV8gutqsQRewdwab
+dxmblb2oARb6hPmab5ZTnR4t+PxNpYbA8peKv29IMwsrE0VaN17lmW2DKJXTDqN
15AObu6kF5AN0tTIOGn9f90wC1ZYNtuKoTSNQSaa0e1WZeyVeiPLIw6bUt9GaH/G
u4gBeONA4hnzuO2atEDwdyn5tObwTbNCdRlE6o9yCGP2LAsNF8fgkd3f1RT2ZfGk
bRldX/pH8emBON67RyV7rYIMkzgClVEjuMMjNfJ6KfHFlh2MUVUeLjmgJNkm+8hW
YqU6zuSHQaSYn/TIY8KX7rUbpBNkF8LjDo4BGcTJxbN6pmFQQG+OXqluQ8A6GBbA
6tKqc7XN0UpBeuvUnpYCkAU5cxypDwYd47HWNqtusqe6+zS9dUx6VPst+3jWlT3z
xD9P9DUvW+FjRnw0PABXYxlHPc3GrD79kHuQRg5tbBm8fqf6OM1OjgNcj8K8vQH6
vTdTYDrYK1Y6wlm8/dMGb+krMrD8htwYCnR5Foq9a9iEAnk3IyJYA2e9I9Q5n28j
0TY0lokhPpobcWczJuporHQFUx5pAcbhKESUxVdZDzVfETIMjtRJeVGjJECPAl4s
YLaVRa1Abhe9GKBzB1pX09grOJYgfEyYykgXNaAKOfFZIBszryXAm61NisNsZok4
aPMo6QWJ70nEvreQ6Q9ia1c3DMmRfK3zqVuK5wddaYkLy4NXy/DNCKRXQBUoEJdJ
O0Ug6zSZIhyUaOJTl7YY4PLDTwPC5bM6DwaNB6ifEAge769c572SKrwt88oVDzid
Ha/2bW0/42npdKS4PSSVx1JkCrN9//Wax9qJ/RX0aPPX1leB40NTkr/S8yJB5k9Z
49VJITa8WYr8gEZShzpmiIn3wKzfXSx30C6kjOGnNNu2RygZC/Y3efvJGrlcqquj
YQ1WaaIYqdLMCiEABQ9ATC6KuEHNOV4uY5Kv2ZoAKl6QPN8A5Z9+fMKuHqvvv4vp
gto1hXsVMyki4hjWIBDkPKJGAzcor22uOs4E85YlSCrJ/BE5HNAG7Gs2MxPIpk8X
rWM/X2Pk5VHUkJWYKtkCdxizT+ctH2ondY/QDyyc32KJoI1zv+jYXPELgaZdQ5MY
PcgORHWyDWmUIK+UoDGomSajcxa3Lv0LlAhWOSBBGycp0YtTvgfjF8eL7J75t9S2
41L505X4vzH6BaE2kOQebsjTCNTIOjlXCMb5jP8Y473CgXCXWcRoahpwKXE6ddYX
S96hX0YSOY6lkEy4yTd7UkxIc736NCWWbqomCtU/hzEF0slmxo0ArgcfYku8SLd3
IsFRNRgYcWxxzKZgZKBai1VEms7c4H+3rD49rCIJUWoAbItZ4KmpsZVHwV+fiLlF
DZqS4c0ctC77Ffn3/Y0d8d45JgZd+ZZ20UoYycNC39VI62f8ul27lpQEy7lRhzLS
dYvvVdukef6TiTHjugSaA8KCTIphKDEORUZHWv7R3ybDx2dGHJpPkZyHJXHypwpR
NETXrMWvcVKur0cQozyhmgFv+PAbs51z+bOHbJU4xWZsSO0/eLYwzjGoiMdUyKwJ
GoUmaf/xRqQvlkN7WDK6TijHLhiwQAqpDzLP49CjR/kqzBL5Iu8Prw6vKdbAYNix
bHjDRdGhPjrE7vUKO/plMOMGLRcZvQ5k+zjgC/KH0iXhA44vbj9ie2sUUfPFl7OQ
8w4zQLKxLPvb2NbvjqA+oIglHKbRBrDZ+y6wnsVbWr12AVpRykyfQQbDPu+elPuB
qQhagSdIDGLwBxujG9cKTinx+tzhmiujj3qtFo8WdCcaFofXYrP5dd70Xq6uBD9T
ssSba6LNdhQyBlkm3aGPZz0WSJlyq89FeVszjnnLNx9U0sErBKNrYKrPFW2Q3VSY
k/u7Bv5/tHn9RqtsAvSFo7RtODpz3U2aoemRkrLA7p59HodfhF/kL9GR4NB+7pQQ
r+rTDi2rZFrsn/OzEKFBf4okrcjkCEyq8qJ9/XMcJcfrOuSZIUB7sBVAZjY3yIeJ
J964mEA8xIiqiaJBIBTD7P0KJ3+sYkqXjQZ8rzEOEXBxjVUbqytZVP+jFJbsbVSb
uPCvql1bYneOVwAlUGkUEQCdOh/s4mJG3Xhnjv/MIyaXzH3XQEoBHs97wpaXOI1b
MGfCYx9nSSQmAMRk43jJakp4spbWTDkzhvo0UM5nBrmBGLTE3JZOR0jwY++4WaQy
CZ7G8nf48Xw1H9MBhhRJPm7eNjQKBt2DnpOlNVngZnDrzLIzo7Ydt/ygDssCPZjU
cWOjzlBIILb9LgOAMg1GZqJc8SK64uC72dP/2Cx+VyI6EbXF0cwO/gb+k/3eqkxi
15SQfjPXrUGwmtyCHCz0OcUKXrbDLfNmH9EfdAxfwobViJFI41khk0VViumAi+Fn
TFmt84fece4wnB6y3bUdzhVhNr0FbaaaMc8IMKCs+YW/d1B81w1aduZWuNZwhXzy
2eXxXnv8MFCpztrelE2weqL+VMKQS5PilzrxYWu/Mqqw2Oc6qPbLk5BxrZUwNDl4
rlaOTF3r8b/1yfKS+5phuLwKXLPOX3LhDBnj/k0uFiM2HaTZQ4gfMi7zgp57VZ7b
O/v2D5m/Yxff31ir14mVOdVRa+T6FQU4+pWIrdw0IEylz4aw0M96QRvXs+XIxFLn
h6YJ0bHDDfDd7ffYPQcZ6Sxu80+lQ2KSm7doGCz5dKXlVa7hrk3NfGeChJlAUOu8
mPE5pRQGKwHCI0JPvuEuMruZF3v36cGunZlwhXLm5FoQ4aAb5bQhREI/F+ZEs8Fh
duNPt0jw3WPBb0L9urxi1CaSOrxv4ppEwsn45hFTPRg0rjpoBF/9P0C5DYD77JEQ
khmernYhVlTI6VHUiv6vTbBsn6kDCYZanZxU85KFKJGG0W/txAWuwN75MLjvT8pB
0PogrUeb7Z8p3T6eJCYklhjCCBPSC9/9zyI5SmcLfo/lOU5pJcE9Whoxeyr6hAjP
UXtbZXse6e3+w3k5XuUrcjuOcR/JSPBl4Q/eyDQ4gInp5FHf6tLsL5ZZt2NtH0bo
EcmU4r5JB1Jg4wz8JKswYem5oVf8k+2ziSfLkuUBX5Xy/l69JCkYXk7gBs3hFReU
3kpkPTb1xj8E24d9eghgGFLDpTIRn8Qefm5O7iiuKr7ADXfgQs/LnMWY+gyJquT2
4y034KxdAovhsoBzWuAyAb4wNlcr3b8moIoVwynOUehacMTG4ET89WMyYGAAjSzm
IF81wS0reXd14p+7Yo9p1kKd2cNveEb7JDZhEf/JXJ9xj64rEjF0bSgZVdhHfCfc
TtGjHXCvUymKbkQEJCZ5rRaX9lA/iUpqf2NSY2V8FEIbbbH0+/zhBm/ml3dasr0h
+izfwCDAPjDjuS4iBZU/B/DxvxR1KOKTFiZoeLGKzngyMFwBHqPhyL8sDe40K2Zk
LAz6DpkaLT+3V/Ls4cdxCuMP9wDQqLBo84LPkIjPdDsmrGYxxg8w9u4mjiXF13SI
vPg0cZMXc0WjghsxPoonf4zjrFW7UBooYWbr1m72yFFJuigLrBa5jWlch92doma9
jmUh8mljr9Ta+LKyBZu2hrCzLWoxcMAB5D6WerWyY9GeHgY6JQ4iGxcdOll+XfhQ
rR3WnHOr7GuGax6KGBOKIxl/AXgvvm/NU+wKAJVwV/FxF9Aze9KN/GZhV3GkMFDa
+ZGCQZGm12suYftpiHwLoEpSINEx+qu7YL7TsUFNwIAaywchWhsznF4ALbKl/a5S
LQt1Yy8T/JBI1XsBf3s4TEANj6W7ASNdac+MVsM0eMwkYvzWDkJzhfXI6FUi429/
v5NWjwo9gPn5Xq1uX5ssb2LbL3Cda18oPwkXzoiiFltsOcji7QdcqhxlyeRGf4sj
q2smUnGdGIEk2KfMFa6YJJDtE/SrmBVXfVaqqYvL57jHCBzgQIap5LsngiakkCRI
ce9a2WtQ9so3G59nPem2b7rBBuyVYtnUtXl//sb9HTAMLVCmn9MG7JYC6leEHckw
z0++Q1i3dIG81KNGW+MkwevUkUVuQvy2CBGjpAXiFEdtj6KwBVT+Fazwtq5EsoGZ
bMJSCQ/eGNmTfAGh0gVioTkYw8WIb6rbt0gbex/NJdAsDNE+QI10twCUvdVvKc26
Ei4Pcj9Cn6mQo0umzbpAgAHDIlIBhu9NVSiFFzPjm/+U2RL5rldIWQa7YVhNZWA+
J/fkuwpMSxOjIfXY9tLWi5uyNtbPQbRFnW0P55hsyupy3qKJOONdldBRC1xZk4Qc
hfnuM5pGV32HJcH+snz1KviEMHlPJKl297/VFe4J+9HYnaDH+nKRxP3hB9UZTZA0
DL6/cnE7BZxZhUXFhUUQRX/bIHyA/8ZRKwpOOzPfh4Py5+kFN7HIJzlnEJxWRMtk
b5UvhxEp1Wb+IAQwrJCIlPGvCDFLk1j9lv3RBiysRAfeQX4+z4MoaJXTDFoC8lqo
qXdop8kuDCdzpxd8Z3wg+vcjYso08ZMAc7CtcKdvvor99VpVoBG4bF9sooH+bM8N
FmBNTI14u1ImxsZNkF//vz0kuZzUydLmHF1YOyrgPQ7J8HauSXENLNPtQoXnh7Vx
PivwC9ld47sqJoMnPqOGb/jxiZ/a0v9lEjCqPzlrzd8xsi1VeM8zwpL5QzGItvCF
jRldDPN0HrB7pe4m0yPV/X5wQIk5eFrRl3/H4HmRVS731jQj3MLG76Ljtv8vg1vB
S4E34ibxcXuR9heRtr0pLzbDWtIYK6uhp5WS5qTL9KCASKSPYCSrXb20157mFHBk
vaL78cA9LAq8h7cVhfXkkCLYu8wj9KSA0IvyShgYgtdaZ380hMcVnAOHuKQH7u8f
oU0u96iBpcP4ufAbJKz9qBml2X4l66gyN221Xevf81QWsISWlkUMMpqJ+Jg32kev
4Ivojmd6JeOZbvXygcaxLA++IVww48VxDTdvkWWVsDNfPw2VywHmZzlJmZfK9pbL
fZStTyeiXUGRAyuGcQ+9oX8xn+MzxInrpo+aa3WDUc49/vqVyhkiJiU/9wjxhIuV
PjiK/Z6lwVvNpfMxnU3QZd/xY9X2gdJdvddIv9i6Gu11tiND3pk/a/pWznOwIZh1
dL3J6a8Mgbwpg/frn9gd0uxybFYTEBY129GtjPNQ2zSJGZQKF90td5DKOenyJfWR
GD9s0O9vP5VMALH4JkDlre1mYeAjILoKxkoFaoNEyNv98rOSjTVMi27Co1lmMdPl
gJnakCgaJpm2HbUJ4t8HOc7y5hsHK8bTLmq3SP390T2BQY/WfXjZu+04YUs/m2Dc
1OUc1NUKHuPC03n1/3lH6bpX0xmRvVpwLgQIZnowoJklw6K8vc5uUi8LQy7WhWrj
mmmc8a+aXOAINsausVz02R37F7fGag0WIvfpI4yHj3bSGKQ68/Pd5vzA+AqmeK6M
A6pjndNi8TUwgCwE4B8q0IhPCOJVzkHr5etof4rx02yDhUx43Qtc/rgVXPdwZVYW
bcy58WZ9wrRQmVgkfF0XO1o6MyuLiq9MHVrDeuxDL9PxYWBKbl/KyqOhOzsf7MGm
OPGOFhZ7ythEHXgllagctIKnkeGffpcAw6xQ58yFkMPWD+5MuAhcIivAFG+blO2q
n9PQ1C02HbUySsOTHL2/0n0+yPPBjqI/iyzx6DDH5vYk8jEOrscd8YgGKp3R/7yA
5NulnJ5b1gaTF6XV5sBfUaLFMXVrKB/bH9PAyEhHJIdm8ZZlm7EB1ADqjyrknqKb
XlZ3D2fx7AUrOaW4flZLZwP7qQGKbhrz5XM99bYwt/FqdKQno72LyBrIW6bkD4QU
9WfkhIdToFuhSXzE0rx2vWMtpV0L5kmfi0NkeCLiSPWo7yT6GP+dMowV4SS98icL
OvrxwgWyYVFBdMW+U8TGeNBZNrOsD8gkovePauofnjXWmgQ70bBM+ykxCWJM3M+N
f3/msw2Xcfo+hr61VL1BA93hAwa23LR/OGYfyu5voBKiAw2nNttAHUrBoHg9ljCa
2B39cgY35FhQp6KtwTIeA+WhlQPPilrqSxB9WJZn0S9WhNb7MEUZmSs6kQv1p77t
l4zzKiIJCZ/33MkLujSRnNkdvjFlLJaPZtryDxtOHvegfQ1gi7J8u0RjGA+dOQSm
NoDHnKroq4VQSIFxbjlHKLm7ZrxAmpY0L03quvpQ5/hClJ/ULMWGSnpf/IkzHx/7
o4JMst/IOgEXDlto72Tk4xE4iUjMtNCHlaARZwXa3CXXQPzK6L8HJj4qWTH7Tkjt
Nj9WENNS8/L38y+6xUqcCs8IHoSKQxY/Cd2Py5oh1oG/qTJ3eCqHIYdsoyrhv7/h
Ae1lVixKADYgaKcTHuQ83upP1wX5EaUDB8vorGVdKo4FliCSUyB4023bp/tMU5+A
GkQZVCAZwZPBBdT8F7VGasmQGH0+vNh8Y0drC8s/LXtzomef/OgMz+p9mKaR/6hn
brWcSttOkl/horFvDy2B0ZLg5z1M7/M6EjXqF9Jyls4+IyD/amr9I+BRLywCyM9c
l0zBcJFp5RvCwKZMlkS27yEZ+jI0UuED3RD8D1irqsyQaNAPAVnkL9tJ1P3OyMik
81zWCyadDBruDa/Yw7hYzGgGwCEOH9lB/7bo8wSlOWDJNcWxiHwt2O0mosknwulh
NePJSnVmV/+wTz4xIFaZ//BSSEOM/3JKEd3NyDpOoT0lQp2Whp3DueEEyAYrNrU9
wOIPikNPy21qXQk1X9x6KVyykVRxNYkhal4MvQmQO+S4YpaO0dX/tkyHYHVfzMeb
wwhiWGV90EVKcHxp3a295bXCpFlf03dfUwDqfFpODh0i+VvMEYY0ORdUKfg44fun
XEnw9UbghUF8+Y5j9H+3VnspNMFmbgt4YeCXTz3h+a/aDIZMTIjwxtQIrxyms+Vv
LOhKrns0bBYVbt34HQFCS0WOYYgdQt7IwPRgrua/O7N3PFg27eynvSuJDxI+BUsK
Woa/qM0uO3o6kEDDm3yGaA/jLh3LWt3Np4E+rsG2kA+bEQifo+BXUxf1ZdhjRNUT
f15aNxCZXL01JU13CVS7jq4ueoIFmAq5FejhQbvxhOalmS2SoXOrFXyYTc+Z6Krx
TWuTOGa0ou1wCibsgY9c5IydKfyUDQNKRz3yHlYKIOA68Kv9/LCjqsvgEqo5Rsgf
r4dkAhx+6xbTaCT90kUlOdloRV3kPfOR0BtcXUXGtZSh0luh9MKM9NkJDPSG87kn
Cn3kVSm+tWb5ksGzoRBKWYoM/x5v9K/9yiN+eTkGY0MEctwmkSDhTuE854hurCAj
EoQjlLGeR1QD4MBrwg9wFmep6er2tN+Xwmrxr6F8GHbYOJCI1kHxYF7/dmYbWTuX
9cOOk4NA67bj/G+sgIhQoSN9RZzJEo2kbhCzeMYQQ5/3oSGAgRqLz6RbLJ1fFpRo
aRBsm7U0DuHz+XgC3+Tu9vlK1Fk6dGszZFb7g1UETvhe+Q7XfmJUCoHPFI7+5dOC
+kmVIwSSSiT8RQ2PSaB2OafcG2vzSSgBT2T3eztcu/ySdWWp14Gik2IxDClhKIFN
iJSKS5E7sfq7GeJEWADlRAezS+OihBVGu91Pv1oTBXTqWRNYMPMS7//wf7M6e2KB
t0RvrTILwpGwXLLsxSrDMiVJpjv8eZJJOeX/IEgTLfD33RRM8IVOakV+mKb1vBlN
51vrpPhlEl9QOkpgEGWMtQqNofAxYiX+smxt4hE9WeSPhVJcwHDR1m/Nn2zOHhXP
oeZ9tihtsYKiCtbA9+Wnkt0zwIN250AUepYUGD60DDbJ13lDWL+e8d1+7eu96ejR
C+Trz/ra9y2uw0lDSu6DZychNZ/rszM13g02DYTtjQRwIuRKTCzBgVoKrdmHVeUH
zpEvrSfL71WM/O/qbEHkdaWbRnZpTeGMNi5RanH2U5TPlrU3pWh1qzx+b3YnUQ0K
ejzwZGy+Ujy6FZ/AgM2de4AL1dwUrumpuWS6li5CXKeSV/Hhejsp0tw03GxQGZhB
WS0NlN3gbjinBZMwC+mfAcWoo0WIABf7gF/FeiepQectzdMKOQ0bh9req+spIcue
6aL0Xsm9ERJ09Q+A3qKpvO/7fFrTLQu+1o9RQjnEa/nxxH5X4pGtXS3xqnIeR7bF
p4ssalaHpOim6cIKMgK+AMd6SXf+WLdUg31xr5mK/8nqrTSK0uj3nXBFnC41ZZUj
QVbiv/TpUGKv0bg6KrRgLktZCLb0kfvwdYtuxGXpNlXIZA1AZ79eJkv1HPU0Vofd
KLHpMzgNjevbWLLXiOSTF1XuEBGLp3oMASmRQ2mAoexJUM85k0STBREYZk8gtG27
SUlZKgRhR8ykPRlwKNJhD5jbmN/biXiKHH2ipinjIwUpg5Kf9z3N7PFWiVwihWG/
cGBz1FuodXVlXgNcDSKDuyfJ7QBQGlKJgeWkUNekocggC8M24IGbIoVGTte3oL0v
rfQQTjkhTptbOAZSPFfg7K5PLCrdWFVSVnrOM0qF72iU73xgUkbGzVcVDcvER2tT
16BSCTIgsbzszffffJsGcKgD5E4eHUq9VhhZzBTLUvmXH88bFg+9BFhxG0BxKu5z
w5CCZeDMdov6oppRypK60st4MEan1jxy1pzP6oIokrYwb0Ol0H9XmEudwx/hYs+N
s0SUGURYwR4Igo/NsjDowv3r0Qgb0YAGAj50YKjqWd01+I7D11ioc96ffZvwjvl+
gpW5ik1NySNsvVugfyg38tLymJZmqJn/ProiV7JsZ2+TfaIvDhzsVl4eHHxFkw2w
t0RcOK553l3LmtGlU8+/Za3sn4NSEC+dPxiQLb3CFR99tBI/canRsoeiyJibO4uc
IuSHulagbY0MJtwqU3p9k3jxf/a5Y6juwT6qcGVJvFGU77r3vW40dr1hB494QET9
+gU5vDbNVrT27BwzJmszAyIfLn7yVLl3xFbJ7Ax+g930Rz2PtNt05ndoLjj5PQFF
oFdnQNF0qbxHQRSELk3BYOBZHbF0bHwLlV5YpYLD8qJBZTeT9A6vCX9ju5HJ5w/6
KD14UpLz8+DiUH2olyfzuqHqY0LyuO0/XaCThcbu3AJ+BY9roXtM05sM2mlRNST7
pv+i0en1JP25KfKiAP1gacHojeHyqRViFNOVWZ5BYKnspwdCRXoiMy2n5IQGUIW4
CHSLow6t7fNsnr3c7oH1PnL4doCjglmR2f608oBM/JfPGsqTjK/S5qUZLMqZFqvF
31ujwNDSFwTFn8RFFEK5MlE4hlsl6eF6VwKu0N8hVxdisixFAbBt9XMjn1tP81wt
xVAa1vugl1h0M5UdU/alJ4XgeVseL52w/5oNClU/dn4Ucgpn9vatP+qiL9/Memmw
5EaRC9KUqfxhSn1hA54Q5371Ma6zzxdrskVNJ3AEROthqA1NyliBWVxqJHKF1I7V
720UUPzCsZ8KXYKWZt1nD8OVjiYg8Hej9mxC3qMF8LxRNi2nT5D64k6le5Yaq0wd
E177/5iECejDzThk/0v5GKFrZb8RLIkn8m7d2QBh3ER9ZzC0aXMMJoyow/7wlmZI
6QvrxhYTJbHemLV/XrgT4xbGjotsvgPbbkvriB6eDzfu67P2MwZpUDuRSBt062C9
bZ8Qqw57ajgqpntfM9/zXlDKiiIPCJoWzXvwNLuXV8yLn46bgAOJDi3bxgPNvjRw
u0sa/uqyARnuJfISB1da+oTyGabDB+46FoUrTc8ae4qwD9Jf8AX5xlFbUHRLmpFR
33itnsEqaVBR/yHB41Faz/eAA2/nBlg0lV2+XKCQTVdyHD3QLehwDeHNqwHTM82o
FNomvCXjbrAUoT3myKRFBke8Y7U1HdYlsOY66Rv0m4/oonTNQ7bCEZ8Btz6Bd657
AJb8CTDZWTiS7qWjPKk49Sik/O3YhAQKbQmxFp0T93+PBuEvzjMG+OBmyXKePlU3
4r3cBwinY5O9OhDcCILUDIM8OzQj5J94IjTPo5GNBJoDdDkHN9eFlVZOOtV0mL+6
ksnEfxzqI9lF8HJUC/R7giN4DRr3qZpp5R1ewdzsq7Ge0UM8NdeeaN0Zuzqsb09T
F6nlgyuD5WQVH8mluk4KmCjWqZNmc9Rdgy2tLzzbRQw8hl9LCp/k2ctId5vsHKyH
vbrM2paoXZkYiczKQpazMqDFCTdJfA6WhA1v5lQtWRzr6awo0aMUkc37TjYcasrS
2K/gsMM31hEsb7KzruxvRgHzfxia6Ps3ygXj7xsviz4jjdJeV9KKFZ5ADpkIn5Lt
PbRkhTteTAXfZpl3YVrWYCu5rHMgueTqYeZLGgd2DyG9ONRwNJnP+EawUygdUDqi
rlDRpcNuno1EfTiB+Sp1PmuZ4hbpynyPOAs3BHfTw3LUOsZOI2HPPM2vE6H36oTN
Va3iVKcgFU2j6NhiIKws1r9IFWl2BR41GGfj7yXJ9HBGnGM/mwGGvyLBDq71MuMx
qWpGJD+FtGWImFZRwuI2V0wOMuXBEZUQjvWspOc6x0rYVSAhij8m3T29PyxmUpyM
pjMVYoK9BFhVdl1kfKIQ0fibp4XQoaDDn4Y45Nn7O4+BRzMBU91uWQyTmdNFIvoQ
rOCYX4/rgFhEuE2jg87Tk4IXWiQnkhJJ1kxj7NcCjF7KGp3Pyf5/ZQvyrPRm3WER
gvdvPddC0YtQHi+hCPZ+InO6fF0e4q1xfSO9Shhj5HtowbrdB+i2dpy0y+f4+z/1
RxBCFUksBLwkVtMnBDlh805PJAu1qLYFuvA73/Iu/DB8sl1KhQ9tufubDrlkR94a
tYcpL70XPgDVNQc3j1CpfvZxyy2wH+SbvGbLdL0f9aepqpL6uan9SV713InBlhrE
7GInzfykWeYgT7+0FUTWMWeAAH2mfuxyw2T0zZwApA1JrO8VR7jsnrTrFOopx1Ld
ni7sNl4yD0bviM4I4akxJNgRHaFxFDBttY+rkuT97y4pDPFwt6vrwpoylpSWHqbK
jKeNzDBtRzXh/8QGOuq7i6o0tZjT/GOdB71HnqL+1iy2Ht+lM4G51iBaJb/1487N
0GrUQGz7CprxugxA2la3NM7GHOLZ33Ai5pc6usKNW30GBX4K5TTcM0LMxKSycOZz
whWG21jDEmcjCfFNE93wOeK3MUBUqFCzbTrLHBWSeqDoft3O1V15D+9dgvfLVHwU
OCQxeWQj1fUH/wRWO+14wVKeYVhF21wpLOHWGnthie/L5rZYDkzsDPSQrKSb8lcX
s+bHFKEscagh5UY3PM48nIf+kcOBB2Lbubq8aPdAbVoRfk510nwDKg9lz57nMWcQ
qb4J82/OPK5Rb+wskT8i0FnsWfEfl1vhiE9ZPOSaS9QexYTn6SXi1+U/+7pCYbUx
jyvFdt8Le4kkvNoXGopnjbfX/v+t22+4wb4uMj/Y0ugxjMT1IKcBrDiDADVwisu+
+K0vPisopm7Iyh/vPeqRN26lmvkoDL4KAPZDed8eOisX/rLaz0s+FSmgN5ykCvqu
4/TUP/jBgk9ZWnasUN+8GJYJ5812ZQH0+vx9iqBbdTcLcN6IFlpoFlGa5vCCtvhr
dxb4XBWydIsTU4gITV9SbZoZizVxY+SBgWQM0t0kIiaHxWKKWBEz/iGDYiU2w5iL
dIQz0iACJKHIZv1vhF6+tjGgK67lofdskjwz9h+djUJlNU0QxLS0Y11GJA9B2HqM
M+jhBcLDsHK1MXOiNo2DcRFqU92GqL3aRXh1xC3h0n3OL9MeTywe0Yqbk+z0GSZv
+llHrUELVhhtcORZskBZQPPXM8X3qz9pjU/AM61ykvlQ3iESt+4vATd9F9VfjcQi
IC+S38B5XJ7dym9F+sw6T3K9B3BW2FBcXxSFd+0TqIoh1wUeYIWG6eaFLiipOnVW
F8d6/2HV71XNZFpeaUOXJZUF/qegvfnZX+OybR3BB495FX5TAaK0Z2jpPhBCHZzc
SP2J2k2Iot2ksWEyFkkcUdyy2LmEYnPWTNRmpzHlaIBIpbCxBDobh7p6EmqtOcfF
RCRZVNZUP3UdB9KipvjUjhwgoDjQHTupbOfY6KfHhspdQNZ5YK3B56BRSEBZR7ff
M2w2pJon66nvMKKRk4jPL6aCSUqJKV3HlHn9xwXcnKXM6adIFFKRMHV3MhaCHTlb
CSlYLPYS/WbGRgocNLIjZ5rF0w5fA05PMBVfUThnIsJ5R0lxcTAoXtmnJxq/zq0C
GMqBan0DeqVdjNP2j28Htkj52wVye9eEbRCFiz3ULh1cfrFunGqd6E1AkUvuuCc9
tZbTOLYUYpkh2hhKWmR6p4GG0Vg3vjWdwIf+FySoiDXMGNN3yCplV9gF9ZUFBvis
ZoGNyuboaoTqaiBdaqThz1rR4k1g/BaiBJUbqFr68HAPEt2iY6c9QtN0ZJMHfBTw
ZLZQAbgX0mzx8cKDWT7yfcYHNJqYc199ku5agqE9DIB5Y2c7KhPLEXCTWKA/Lxs1
vDGL5BXoudQ6lSvUm8ekZQujjudsX2aWn5sbW3WBDCKK6NdPkKaIb90RRJZexcFR
T369+ybpRTzwqa3sJUrJ9P8RzPFxWQFKP8L7YVDQKIklSSFes3ThGWiFX7NfUxp3
7sjbTsbJSoPPUvaUm1SUOBArpOwjRU+ieeQCwar14f5MRMRfogFKLphVU34o4p1O
UdDgwYIjWcuhBFaA2yKFcs7EeQ661Eyfz4FtKNG3uahR5B7HxiamQMQ1twtFjaJh
+Vab7+dof1TuUMd9q8mEWLR31NcuWnLV8HPn/RxMw9Ez49bO/4VhNcGLTRcTxqaD
j+cYOIWFTVDr26a2jEBZKZm+piwjFGkYQgLwSZoyu9h54Hgw/tYXYHCsTQpfZ+cE
LWoYAgwD3WTCpNl3wE33GRZaXBrtowxLApoRknYeTtthgtVBiqd2vhDBkY5DKyaF
8nxREtG4HBTHbGaeU6Pxywd0Q22Ytkx91ad1dHSVRxQCwuIwFFAeCV5n6iGL+YQr
N3HmxpIzLODxnd/wKGpf0DoK1nAPGmKJDacE0du2m8J9g4+fTxR6SXAsK3OtHjHR
H1XZjIz5zlA7d2wGgiuO8D8wzW0vPr9ljQl8WpFPw9isUmwMP1VAxlifM7WvDjVB
Ur4F5rUGv6O0EY1kO34OyfdV5cXyK0AC2+HABGbXbirXA1fEEH2qJ9XASYFw4SHD
LfyieICOP2bAZzyDLPV4CokQOm+tu0Dy+gnTqhnP6nGoIu0uNvXvYa+PiI7LWWsl
te6uuLLOTJ3XdSNpRnOaadYwKt+ETsfQGkpDnU3hiZqJbuz6jrLjKPoXZzuilb0F
gLutRVp9W09EETSUIO/kE34wDDF+ycjUUJcIhZjKnlzhZEsLIvoNYsyVe+lPBo9K
2BhH+pWwYseooQB0hQLrYRwpa+6FiC+eFEG4NcHIBCPZFVPw25foJmTGaL2ZcDzF
Ha8BMW3r2U8SC4VYkBlV8Bk4VSVlsaRY31F3D5bLjYtSe0BM6UNmBQW3sPBO2E+v
B3BkzR0P9ZWpPrM9JlLU1nQd2KSdP/SEjpXfFH0fIAvJMbj3eH3eaCAU9t7FxPHv
ix1/NXmTwcRF++kFOXgWfWY2ltDBhZwmeitDwT3FX9IutGXIb1U9aI6gn5kqDdHF
Kff0p7l4+zQwzdBDVuglTqPDyF3vdNlRlZA3TcHVmSc57l68lw8myy91bUQ1DWmx
DIHVc3sTalTH90tRSYokGYqB8PiP1lk6l0CzgPxCtO5iWW60ccsv4FNr55+G4yKD
MIX6b7ulEtOjWxPx2QjNJsuFt4NbYWEthHZd9KzigFQ9/iU/PBJc7pHo+AyPOhoK
FaqojtazMGePsg+h/BPvorEpc3/b6m17bUwz/ywwYvLG/+G0kc0P4lGBqMWLHUsW
wg6pjdVI97SChqDVy3EE92DcC8u9qOzcjJf1Ho8zRFTlckR5uQ+8LRVRDbdoAzQ9
iZ8f4PhRBrilp1qUTHil1PUbryv1XiRJelA5xMXsirdbA3CG9bzUQ9xoHiBixNLi
FZNqCe+50R4RWyDPYz27EXXDdYCb9s0mCZoyhl4cH2K6Hd3eY0YWVF6LnWQjft/0
F1tKLlRKWrjOG7ugc+Btw7bAQg+lL0pGmfLAYkJHMZ6Ghd1Npbvu9UPSnoai070M
JhVt7VSCCZDq26elCmbnQU2oR7l3L48fZQc0VHvhVcwkWLf3rqENBYfFp/Jxa7ap
hUJmKxo5JgkNmYAkxdib53Yo9PHlDjhSJIVi0ZcupRHOsAv0TY7+5gbYIz+HN7p0
Q3q1b84VKqaEPDEPZGpEx+50/0DftzV/kFWlZ97OOV6+AnzVEknat8smOG23L29C
ivMatztJhZncYf+yrIrLCVe7FZZBVKogwcushZNw/MA67PM0AqOuNqGg1bQjQK2c
hn0MZHjhbxqG91hA2MqjAwmelV6k7/3I/6MAQ3anXVLnLD5NJ0l4qeKiTCDVrW2Y
YM+G2Jm6QqJkz7QxTB0Azj/pT8PUCX67YOvmfpiZsBuRgnaFNqAQBr7bA9mbyVrI
7mQy7GlpxoQvxF+qHWCzHZneJLqVLdCnsv15e5RmCqfOY3Vqho4fyItsx/HxfzpF
7aaP/RMGf0LqxG8bAjUjuW3pjPcKVwbhAhAWikuiWbWQ8U790xdMe8UvISJtBntW
DhzilHW0Ym+EQ+Bke3fRXje5CH4yodGle+0Ld8MLblSxvrTwBgiVL/664yGCeywq
wc8NZYbLDZfwT/o/J7axhbzTzrL7r7chnTrmEJ7AJmRlPcNg9bOhbITQ2CvWN36H
7z6Q3e4IYwBbnRUDlgRvItj7CLqq8x6T/RloWxNVnA2EopA4cVQeMPP6/PeNVyPG
LJzJOFAq00fwUYk+Xii5l+mDloBLpjTvYYJo892YKPVtubTPGO9uRwfWow6hIO/X
/15zUXgJS9+hHIgNjl+TBrfIdmDYWjPyo1kYQE7q+zAbfOfZt2oVpSxY6e+knV4G
IXt5Acivixd592ppf/4+9KmixNXpafwImSZzodSiMcWTZ+MplrweuIPtrBeuhbVd
xUQPU0TdzppEHd0xrSUlAIVafKhAMtqEB3amcKtvqbrsSr6zXsIj5q9zN2fRsvIQ
uB+V+o/qu2+Y8HpeTLy42GmYaqZbYBL1W1dVQC/hKJLfO47rQ8e4zG0Mw0oakdRK
1M5M0ljeC7BXju9vXxQ90XO5T86GvPzp2SSamvGR495WaAih9rKuK/9BuqDvsHS1
jxqjNKUzvOxWGyuJI1XoXjXsCoILAoWWIIFpXMr9tjwYsOQv1+Ka7Qo07tCYh8qO
gA5Q/zNS77wUuUbcerCJX+G/0QRR35xdsZ1TEl348iDUMmKXZdAvK1DgfHMF9MtT
llEhcAwmm7jfAaiqElzQJSfpFy8AHZz0yZK8/uJSSewtnDC36GCHIIi/Lw/3fJOI
/e0SUHvo+nfKb8XXV/MDn79TLYWmfSQqB1xGOWCyptqAshoj+HurZ5rUTOeCTr5a
Wz8s4nqkgLZxPgK6+QyYHdF0wZr0y8go7Vqz8eQQMrGDQuSW4l5WPSvQ8D7RKbuN
t75vi1LfZ7l3/VCQHmWFv2DUeksRgKITbjl/NmGBNMNd3OZyOC5Xx+p8mGQn8U/u
YOcVYfNAITBof1FtGy9Zd6QMkpCV+ESh6mutdyKZJhzX7+w/oX5HfXJ/H7lm1v4e
za5GLYXk8/qAo/WYCq9utQQ9g8UBzlNsT29h97sXcKQRFxtR6GWOIxlKgbOfrVlf
uupFtYsNKgS0ZCZRQVuY9/ppIEMusI1OECRYd1a/pm0Q8CU84jrMiSnU1slAV9yv
qqquS4GBO7BRXpWfpV6miA87BLSXzbc2tGdS+36AsOumS5tB52JzZYSINAuICdXa
XvEMbeAHADiqP/3LphQ0RauH8A8BcdvDNaYLNNwaTdJO4QrGrW/noOCYQ/Rj+IL7
LmumiHqvxU0bPRo1/OZc5inEmPNveKaDGtNBkJ8WhaNpcZXdlrAtBBps/xvRdPEn
jWC8cH62HiJbPsiMl6kxkGJmNH91/vJntDPpiyv/WXRlMf7Xb6VWagFSVBkxHu6A
lzGhrLSTHpuwVYC2kIM4n38W1965TqxHBq6C6dQ9hFo6YBcm88bzpRUPVUIvJTlp
xrrA74MISAYzPpG8f+QPLu1mFtwww9KUF7TYZMCcDiAvkTzvfWyxvVuz7t0fr0JU
/ISPXoNtSPOWpPxLKQNhyaQvWeLu5fSSft/FREgsrxrHDxE84dskvxFBVz4Cbb/U
iuN8/ijCrDS8TmfZQCOyMePLzVT+hYT6FVmBzG51+Hx9FVy2ONpzE9cGBR3aPgon
eqJqZwM1jsvNQ29PCKG/Pgm7c5N+GyBpUrd7tuOQSljiPuRVeFNC9Roiw1qQQUDO
9KvhkMnSwNFCH2j8bTgLsyzqRG9mdMSz5dypY0XxWfScBJMd4r+IMGIlTsjtimJ4
UJdibFA50TZcb5cbQ77sTgM8MU2ghKobvCGTKn4fmpOU+QJGJDH4WCv/stBDRbX+
tKFYmLtPRtO3xuQtKTTVj6M+NIwS1olaMh4LZspBdDcZ1aiUgdW3cznkLSAW813t
P8gdoC3Uni9yO4XwmhbQZF8H8jkJ7exXkVETafR4RC8EQ5zkrN5YO8d8VnA22EXk
de1oJpcDpuGEuWGCtU7Y0859ZAjA4Chk+TxcMAqJ9i1/PI37b6Rp4PXrYHux9uL6
g/JD5wpWict/Fg56Mn/Rnj1AAydlEVD0bgdtCTd1hGa1ZKA+KrPbUs+eVQrpNqZ3
X4ygYZBRV9GqdzJEgE3T8ChpztjBLI+Is9MC5YMfO1DG9kgBhJjJlKTT7OIoPASZ
muGyX+SRt9RSqlK2cC51hP+5WgzCHD5dQsRMrZ1yN9Ti+HsEfblifxRUV3nper3a
dqpE4NlONfzU+ayCU5m0sxFqkKaFXVa4FvyZK0A5Yjl2udHjxrpDFtuaT1P2iALy
aKpCG8OfNW7SFJy4pajc5Q6fROJHvxdmv0AocQxaPZG7it2UXhNXQkkPDR2r7UBg
/OnkrBNogY5akHJysxBxjGTuej9y4Yim0vfh5OakC7joiEXj1/WsDlPCnpHumyql
55y9JjcDmzt8qzZeFptct1mD6hGbKZBeVpOZ4aXgYmesBe8OvUMjQTFK+xXCn+Tc
Ysowa5k2t3bWTOEi3kCJOaScl4OCwBsSVS9U+b8KcEzkAqHgj2gbqjNFO7HPitI4
caewUc3Dis+hFrxQCMez7bwyLZrTPe0gYla+QC+BcLfC6e2zw3/uOOkv83zbJJxs
bDp/zfxquK1JY6VjKSYM0LQ/5eS0MWhQ/MStrQmluwmk0YZShGm4feQeZUKC/Y3V
iqlJW5JAHWtajX/mRqeF3kq/UEuKLRlAJG6+QldVEdOD/miXtwZq+b1LfbOGTWsD
eAKvlqewWHsohNYDKfOFYAgcTz1xVizm1qvX0ZfPbzNPMxDUhEJF+IGUxxscWl+u
cUjwVETFNKC1Z1kiEYyrSOLSD7KF9avJSZuY0WGGAN/G9kootu8exSjixK4Wxly8
hmomoggqG/7CkMmmBoVUGYRWPt9pii4iGxdT4FP3vXjwr9WaPUtI3K2tOF95UNj0
SvOj9oeMl60be1865PVRA2PrmAwTDh1x+0wAlk9j6xD3CQ0uXrNvYlZy/Pbr0xo+
cw5rhgnOxKeepV/Jr/ThGLNtVc/0q9+G+YeE9utn81jfY9vwmE1i8lttKtRJJdND
LDwpgP96olRCWU5fA3I0R6HpGSkS1SZB1kfMsK+7EkjoiukWDp2lA5AACLsAuWlD
w0bavxJmiPPWP5FGx/2n6NE0yqvDu7kkAt2C9QFPaRqIdKi5ztliqyXz7qWV8Ytz
1D+kJmYRPbw8rvb2RllMoUDZsYZIuxJyXyBUoBGbn6HWXdLznxhYXk4m+ZLqe2QK
iZmYx/V/n2gpc1KxvX4RYNJO19/rq2nbf4yrfJOqVL7LyKyFL3q4WZPm9rrJjqWO
ytChk00EtvHPmpB2URujvErUQDM3aEaHZn0EZLDePd+z6g49ai6EiBSly0odKXWv
kOGKrMV4EqrNK4d0QzRfCdudg7tAu/LZY2mTyCgacf7rBkQ6fhnjXFfz8cLc7orV
tyw7FK3ZrKGhWfjPPse6BjZ/BxwF6yGOh8hP1xg2IQgMn6jm9SZIhciI9ImVqiRm
o/mj9Kf+JwJtLLel1ywb/Ipf7oym1YXhqSwVmSxLK+Jj1rsO+LxWBnTKfktIboxr
AGA9qTprJiejL1yAt+zzFR7fn3SyUtsLOj4iAOr2usA/ZQb3hoHXx1udAbO2FGwb
HO6MhOY/+F5MhHeWHvXK4ytq3dI2m/x0oT011IH48AI1kkloQqUX/IOfe7Htc9JJ
d+WPsviWx313LBrukp6QTl8Vapc8INkVrDnZnAiUkYX4mmfLitWIUD+iJZEVtC7t
nHx8+toxm7YZozB5Sm044RPWIQOegJvM2K8SSsJ/FfkVsq7gQ3DbltdY+dr1O/TE
kC7Ze3eBUwmtsUYN3ihgAa+zWY9xvFlcVfYnmVz7uy45TqfCZxoCzZ5GMfWLENJc
QNxZQYEXUv+KsogradUWhV45iUgDvromcIDckwlM05Qm41A7WOFice7q6pRRObZH
qiMbQgd1DuYb1eShueShY2rwA6YbIcMI5DP7s0pYZxbgR/zSJzGKC9s98+KUh9ur
X4k7KwGcS/HD3E2kzIgT9ytLYwVo7DXRfepCm+8O8mRZag7UzdtxoDgc2sVQJHcA
34RmpL91QIcZjQkjOTOzzcZW+TE7/nRg8/iyh9MHxqtQ9SHSLko1c4crAPSfKJxK
XlavnUFCz2B9Ll1g42IOs+k3D+BHGukd+M7IIXISTiXaa6qh+1ujQkT50aqxMJa6
BTO+2vpmibAgX35b61E2RLXFwh6VBT8NX+nM8RXuixsgKnwk0cq7B/6iQXsf/ype
2zm5ANsV/scDrNBoOpypzsm3IDqvw937wHS4IEZr5QMtwKj0Sh1vbHhQ6v/8yRi7
wahy6CIIjsctSyyzCnkmt/gaq+1jh5eYyBDtansP6p4UtXtEq9Z6bu630Eyg0aPb
4B3tmyG1DTUku11ewRuPsatLFmXWgp4bQ30ub+yhb7/MzDFhZUdTj7oAIm/6+juO
1x12xatelJqqcnuvebUtu3vcs5m8ImoLqBSxZNO1hFdyVj3OuBN6QccQEy5QAFxG
HDAuc2o1+yTzDafXuOJefCcILWuzmrceqvj69pjqEfSUoGUUevbno0JRzt9h99Ww
Zd9JZRYKNWr1ufk7kUPYbyaJgB1CFKmmR1GILN/Qm3UuZ95Ltwcvk3MZXA3IgXb2
klZrVOmojFHxN26/uYEIjBy/EctISQOnPprGV0qiIoJJoMBT1wB5UEkd3OWHwVC5
pokWiHS43YwjRGS3nF9GJgud88DvB+wk3Tpc7ShzGVJOrbGk+V4CczC4HM0bk4iI
NXy3kWvd2ilPfQk1JROsiSvR8r8zzzv1Wsl2WPL4FdGK5G71mT0Omxl70yz4NrMv
zp9SJBN232eXLRLIp1zbE1ps66SniL6evp2RsX+uBnPQ7/WD0CJGBICd0it3zvRB
7wE/Nup9LKkCPWmjK3A2p/NG+JY6M++wMOo5lPsjIXsARkNAq0P+1TPqhfmqYCJ6
y0fHNa5Y/39+vM0NYkzqnLyPyLICiFPA+MXi2nFMdK2lccyzDIovBHaw+m3Hd8IJ
CFfc6ugJIvd5ps6ZLUTj/55gkZnu+qvHoRNMMuSEMV+H0A993OvjszEGe+l9IAsV
/wXlM9NDrq4Qg/+x7uItX4ut9L07WfS3fexg/GaJ6z/E/U8bezzeAUj4OTfaP26w
TziXeEJvDPrLenvGvk+wEJU4I+C1coG2if+qCiArpq08CI8oADK4ZsKlBpzShoBz
76klnf8oZM4UaUC/b0ujH7jG/3HCgyx9jHYSGx1PGdZaX6/GdWwLMgQp4pCi3px/
wmDJVC8Hgz3H2txA0x+uOi4eXjIZHLuexOIJmjVrCbFXQz+aLIfHEt4/3T0e2Awh
lkmFWDes1Mib8+pG/dmwNACvG57EP9GVekHlCLsWnsRgMLFWzojzYchJMf+6pRGq
qIagWoofJFVLeIzeMf2ozskzJUEf+3DcIXcyYmx7u/3kyZqLuTa5nCSxBZZo3csj
QeGEUs7jq53f+hpBXLwVNWeQSG6j2JGP6AwmYl6MchYN1/FKJ2zZVkAXw9lUt3BI
DApmWs8tIaWyy0vsSnD1rwasq0Iau0mruM8VgWBpfaycroywsjuTQ9Q4xR/FWWk/
iA5HIAjuB8TaKvZ0C0BNboKu270sqjRP2A28ToJuTaAIlP4GjX3mTYozOxD3viVE
uSrArxNAJ+zhSvmzhZPrgLjzejOEkFgHIOtRKcO9H07OEHpPFUx8LKh/DX3SRvWG
7Qm6fJ5lPf0ix4DEkJrVH6IRUVZbPc3PI1hM5CLxQCs7wR4nQJ90S2qUu9LlVUaf
lv5hPLIxtpc33yCq9QKqHtgq4/onl6EGZ4jydPwsNvYaVGJQVV0K8DNgGQD7exoh
t6ouFOM3b1kzS6ZmvR71NvICGkdvEDP9HaQza+XO5GbkUyxq5Jgt+nxNKG2o0hdo
clSiTRWNLECBNLJvHtN/VwLH9VAu30DoCKZ7nugzujIBpopjRCuUEH3lApWSOBAQ
UHNYX79vIJzARUydpzAV4aWi1/2H1YM7z6vGOyu8Kye6xqkxwV6eFuc8sS8L+Tr1
egv8NjtGMdBu1zCf/wDkvZbOqBxxagAx94/ltz7zWhC8jEbHGRagHJn4F6cZsRpY
wi9CRH8yru+ekNvoRQU51VCHLb4wcQ3jlsw57AcL/J26K1hOC9NHmKEzqFhOgXyf
rvjc4qZCr9EpPUcBmtZ90hcYRVprYOeS9cq+HxPJPrBC6mJBbX5A3CsYKnNy2f6r
rBdfkVGe10V3V4jnEBLOayT+ABZ3K8urTIzH2vNR/1Fk81KRFxR7tZdtJ8xmjABE
54jXj4PjZjVEc0U43Wk97ICwoxyP8Ahm+2hyyp1jNw30aLcmp+FCyVoOoPdvAcWf
a5aRUWFSYsRUgi4ztfnrLn6yEODAnsiwuRJ8KhcqGpHJhPRE3qX9YccG3IB1OfSE
NyTooGThaxKNHPSAuRj0G1MybQJtqXXnDlTyk/47cBmI8BhaOYcjIh97GDBxjkCC
laqmIZGo0bG5zbyh66wiHefb4VPO65YnULYyWHvM2CD3FGW+BClJbKk8NrdIILO2
mb+G3Q4i9jI6Ciebr/JdTklwSjgX7gy0Ssm3zkyaVi7vbbc+8Nzk43fZdS6ZSoPT
0+noAxLWyWT1tl/RnpuXcuH5MYK8AckEGPL/Q5o3OpOthRSrUbQy617CWp0IktN+
leaVrd08+gQg7jdRcO/X70/0rb2y8H7RRs4vHa5qeWCuh4f62ZqX3k9bMBgByE7p
D+m6D6qVkcjEtqQBCVzGN6VvYJL83mjUM/AWTSoJRUj9ahwSLhuts9lgI6PpHIJX
+V1ftiDcjksCFM51iLuL171pJbDLjrBSuPrkiXvi8Cuh2OrF/Hc0iVq9h5n8LJ6O
U7jpZGozNq1mbxEU/63l1pwHl8VKPW4Vdqjjc9N0ei8qeMnAadDjMtgJsxY/WGhn
O0O0Z7DqVQkReGa9Bsob4DZvjLhU/ieHk12uShIMZRznSKZ6wsHtO4BMdSa2KRm1
mNNDkz1G+TMLXnY9Q6T0yDy7NGX9sd9PLlf+pzBVxBziM6reAFbSlmfRLZ1fR9sV
0FqStKw1FmGpUqeMoHt2pV+NA2mfTvvENBxaEU8eikgocAHsqB3qVoANYvj4FI4z
t7PAY27vqR5Yk/Mqa396QodieCPSbO2nyXoJ5Q+ipYi1UAhgdjkWtuQQ348FKe4V
WdjJgqVikIlCrZ8ATj2I57/eMbHlAKZkWY20Omsl134dqxSCsrSBWwYh4fFpM6ij
X2xzZ304zgvihY5G/oeKM4xRJKQju9BR3RBAvMsOFF/LiEz2/YGOMtb4C9TZrl8y
VdY0jWnnIl5QUfrEXJMXRXC7aoDKx3Pxj6f701evI6YAPkFxLk5/b1Za6P3dnCEk
oNvwYKQIL1twZZbno3u/WtLf5N+znopT/5k0oZE22gGnDlytqXNu0PVo5Lw/d2DP
jMHMLjvpSErxXAPZ+blRefuNJwiooKc5qqNJjzKC7xLUYT6UHlESzg2IFU3QMi6b
RgPZ3+5W57ITpOHY/MBl8kJGvMngn694RQ/cLlOVmKuH0Mx74r6+G4Pk3d5hFdcW
L+LeVL29NiEBH9EnQb8fo6HrSJjAESICB16CA4z01CrV8obgn9kbp6WYJDGPfwGo
NFraPrEfPxsAieBr2Ap0K3sJVKAqctlUL5REBQv/QggiZ+GpW1XQgVND3viaoOvJ
YhqO7byEMORaGJdJvG2VpHaz0eSmnfLwUvN4T4KXgPdoINWLDeVkLLTlr/NBUbnr
37pf4fszCaw4+Ui/osT9dG2WyrzBStr93c642KST3m8kk/fwrRa4WBsVzEtjXIKa
c7U/1YLkhbRfebJm6Zy661ueAlmVubbAygHj60Ba6Cnm/hCpXuF/1DywaKEocTAP
veN2fQ0TjNzt7cu7dUy67p/edM01wBcEZJUE0muHHKP4Ri0nRjASHGtekU2ir1mR
ky9BwLRQZd0PbxgbWGQdnR7TSRftt20JbBvzcqWcm/mdL3AGJhfd1q2A/LSFuTEF
2yCGeP61vdnWLpiQJOpqD69M5Lx+FIFuI6HuYfFS31oBHx9v5kPkHWJsOW/mkhRJ
o2mXRZh2ZTkQte9tpz8Wx8GjQcyt4JuYc6cHgX76C/PzYwSHHyml3DUTLhgKlCPY
8KHAb35YU4fv2Cp6EDDf174cIcysySrX6SD95cxnxBQbojQ/N0caKtf2YVDxyf1L
TNoRYsK1xWGEEMPbjEAHRSh+3wNHA6ovfbXhdZoVNsGHvj4fPxrYkEfA+aNhCpNc
snNWDKyptAGak8xmQmfyeoNYS2PubxFYXNeDSmQL0LNHVuaogenETD1CmN6RqjPj
BF1EoAa1A9MQGCcpnH3hzLGdZapNVVRPMOfS3+w8D+NLYobc4pEWEGlVD95q5day
S0np2m6UfAFAtfJCG1kbdeMY6Z90NYbVpqHul9YavffQxKuVWa6Tlee1p4cvZxjD
RDC04VGVgsQNr88WpVkoNlSmcSdaU/hRq/ClsLfD0qDNdf8Tx5hTtRYoCXk4iOY5
XbmwqS40arsyKGmpSd3zc2IgUFlZQPEokA8CK61m1TCp77zgHZ3K/SrM3XmVJxfI
8arCxDchJwUq3jngazZ1dNvO4GiTDjLeOIG9Q8aMTYr1/4aKvLyB2AMwvcZ65zHk
xYZO76qAzVYBuw066vMVcoyPd0J69e7TSBqscFDH5R+tMpGAvcQYckhoe2YK7i85
VAQciZ0S2sPDFNdqQ21dC6yvS8nPhllW8qm6d8RI1F6WRIb3X/RpyiTora+J49Lw
/PHPhTByu6QCZwPlDm1TNI1Wef+dV++K7Dr7KYqprY5P23pMd00C/RC1UnyKjTJy
/vrcNf0XYk63FgLwfyhr+7p+HZGDthV9AAy8CiKmdR2yiBck5qJ3jb2z0X47jxj3
/4O1yEYNdE2U7NoW6/NzuGUZpn2WxbMuO1wAto7DCKQOfqxiMwShNe4WVIuhjliK
XLhxaa20aAAwrAgEslXHDUGLV1JJvVO8P13Pc7TKZlPv9u/hwoFj2P2eNCuwqQZf
dZEde76ZHG3Ej7yd4WrVdEUhAlvPSHyRJvxWXMzTzk0T8juV+/ab/v4ya/0KcWk+
xAMPH1+Up6hVxbzeLUf68x5jPtouIc5+kdBE333fJvlc7Fzney5W/Ip9t+CoEkfJ
FEkeyATcAmhbV9bPIrHZ6N0w8n4Au4iXreTWzX2/JO9lorEpcPapSeWrohAuuojf
4f6PMjuyjVyxFuLpgC78SFY9HGix82Nnqz7x4M06PogHtW4XhhpnyvgoJBrZs7Bu
xbaFprIvksVhwYOoPkfim1dFI78rKXNrwi9PEVMpLsQAeIrN7YZua9YOvrT0tQWH
qDIFn6dj4ci2YMs7bMyvNJa3Z4v3zmVMuALY5jrmAd3sHAlD0UA9RZS+up/V+2Fa
jdnPjdCYiG57ubPeWORoqDjT7BxVy6nv3WhIP5IzrZgX33hRrYgWfdnmLm3t2fSJ
IFzmz8xTbifI8pfC21Vx+YzQETaVtW+23i1uM4dNXH4jVd1CzbELXi41u38qEhQb
maLgyhpjnleUngcJe+YERYut52MxosDIM0IRverivesYOzQUAN8jGNCK1vRtkRxE
CuWNTtcAczXvEpv/EPI4uB5ZCwep3QkN/V9rpC/A3IZTkxiRFx0Mz8sFQBSvk6aO
iTPa2F2LaLuZx25nWFN1GQ/JK7+PU9trSxdYlMv5fJHqrxghFUoWygd9H8yOmRRb
2sMnLH0aoIenm7sQzOMl8lUJ/kGjqagn2UBB4RNgyEfaIURLo/4SSYbHnVdt9RvE
DhxCqtt7pq/5ICEmxromce0w+WnCPyb+RwIvpUFH4aMGEpOPckqaZuHKXotl2pxY
CZhDBmp7nWdIg3GJeN2TLhIkN4FW3X0f9dwlNHkchWybN8c5xwOOfcvsD7XMnpb4
cPJInh0Hw+Aznc6TGcp89TPeu6xW+nz1OINhnZtZpQepQFyffAdkrd8sDsc+F4gn
LbDA6MGwq1qgpenz2lpeltMEsONt1IH6TOkRsjtB/E7tbsgXTRL/DtGEXExCN344
pxz3ZkP1dQkwBlg/A3DCwXbBIYNq/EkOuJyCPmzOEDLuc1w4pMNNFhTaYljy2eLp
TaWBlJI9Ybf4AxI0NWNbFskR86EFefMRGqUvSpjcLhcwjfDHwTsOAelm6kh01bIm
oFRP97uqEA/phAAhkWY2Nfl6O6TfD4LNnoPjNcRUARAgb+ky9JzN6fB7IN1r00G8
iZeJdMF145Nn7Cu/RqK2vi5G49cmi+zUOt4bvLFRdAyrNZZw4R7dDOJuERE4bRp1
VOuufx7es7wmo3AOCUhqfVo/wR8UVTL/8RZkCvmHK7MLFJqBD1fadUSTGz++cWX5
fVb2PfN84TiItHgFr35StcsBauIMoJMk5qY4nE3SZ+ciF2lxJ2jzJWxeC7HBGV2N
hi/F4lVeRcOTP941ueSQQMCh2rVA/58o3nUQKfKY/eAEuI4AKbdbygSQNtK9nRcI
/de+zPv1aA7yeqssVcUhJMm46Thee4nUOaTc9BWNBANucx/E0OzbFOctSEsttPYZ
DXX02qw2Vq6evvUBWsvJKhU5zKDtzEbyTM46ci/NUDxU6Me6ZpbcI3F9V3fu9+8p
TQV3YKkcY4RZTqKqVYjT+EwzFCLBvWcyLd3SI1Rv3yHqK6efUjTk/41poPIlAlWV
j9OmNkVBCpqersZbRo5Rt0i5n+dt592UjPle9SHzgdJNGS9tAgqi2yC5Q3ue4Ioj
lzUTgrd1T1QK/tqJPAerAO7kimaCC4g3WEz1zkTNo6XRb9bbMu5dOnTG68h8YJsU
fK38oGrhAPw5OaVphA314c2q2rKCoG2bPFWtcYmBo/FYAYLmNkYMnEbgMtEn0RYJ
NjGYoQdqbbXBdJ32wrC/xvNB3ro2QE3FnnPyghEE7jqzXMO0Vc0E4VMbsPCAMQwQ
4El0fvKmmLAhV/NBtTkvotdALruJy60G4CaYQEzWKcN3jLMaRDYjgWqLIt7+aF64
z95hyLX+u9tZh6l+4iLs5lQTOM6h3WTX1xL3Oy2ECOSzmUGb4QmlsNAqAFtghkxa
N7iV8khc7nN61CCmUWN9zaeRqvPZGD83EIwNqXPwpX+7zDQ4iVL5lnj1URdBwEEo
6lil8R067jY8tkE1aO5z0NrRs19ORnhZhXVeG26/AazM2xAoVC8HhLuHcIc/y08F
mxIZP3CvLPnUi1gOx8BQfQKndIe+wuzpz9kIUXlbb6UuW7hDMri9GYyDzK2N3pAa
NdjA907bXa7IaWYIdQ9JOlKjnRFxUwPQoynO/acZ05y8P6tZ5u0xgH0s282o1uT9
idTHpG2hfC01ZJ7KP2YnBTQql9EkUk7iv5xifngmDNkDW6zfzuOpkMtSETOlv1Um
6qgMXp+v8DdKgUv39D0rt0uHEDKweTfRbPjXBTS5ddnSBpsTbOPS/2cIgV22A8pX
Ki1OXEQGcBwSOKYZtKORXswJQYHdCFif3Z68/0+iXvBB7EaD+5WKFAb2CmUCcdJm
TuaGQAya92KxkMZ6fRlY886zsi66iFFIRqr/Ea3iZ/2YVOXKKnf1FbEdbGPiVjOO
fUaR0yWCQ5VAa97ZfId2kM88HWIVNAuX+u7gZ+ldhb+9oED9pe+qINgRMGaVXUqG
/Sar+kkShVN+PA5ZJozA2A5ym0F02+v3E2cuiUFgXOG+8G94WsoG81xNpCjVDkwA
OU6GrY9QmzccerqMTgwiV2ayVAompoKUwDP2p/mZtiKsydoYoNckt7zTnTQ65Ape
LaCjhZajbBA4tKlZ/fVwFMxxvXi6FV894jAWLLLn+vXyBf5ELZoTY0ofDQqTYa/h
ZgC7+N2KX2Qtw87zsk2NmmRtA8ObLO/sDqpky3iJE8jeelHOoihF0RmHWioEWA7g
C2hrRXPgD8UDFZggmVC6Qs7IBq3Oc18aZ9I/7FzcEOFfk+xGic4h/7OXmTJIh7qF
IXqBe6QbhIPJXu/40n2Fk9u6jkACyM3QJzTSj/k5q5liJ9Mu4dnj/lIIzNKPNpRw
0rZ+74khQ98Jp+3mnslexlh3+jlE3OMOWxwioFmdo9cIMJ267bTJLsFC3BQraODj
AN/wsaGNF+MZVVHRXaU+9yiqY/XDeKipWWH3UbKEMOzuhiRsRYD/qmjVSq1TtfIS
mGdCIyt1027m7D5Xe/knzeGEwvkNTDSGOAgKhkxTX5NvlcKVFlK1v/huvdCcx8dw
Bxb2qqHctGBBbn0sOdWqOOuS00rto5cnFuLU16+1CRrTL168z8wr8QsHIU3uli1V
GOeVPOczpZRPmyhnhQhHT569wujx+8O0fuRX/xa4qQ9iQyqeAvYRPGpYzb5yBCq4
a0/fqjRwIqbSQAwGxPP5qFsS93lqMe/5cZrjGwgxJ+ZYkolcbK25orw3X2rghuvr
ruXcnKalq031I5rBpirMza+7laTHRrIe/AvMxsgp87Bb4miGoYXUADPYzI6rOSvi
pLuJIwqKUw6UO4klAslgCZ84Wgek3OuLgYG0rtHJWzfeGzAls/40hMwd9VEm4Wg1
OmqrjYYlOqVNK3qnWeYedx1tmbloLKl6l9prBACj7WyqoQ0qYjyVTULkRanmN0Da
IH2bgMpoadcgi0sUtNWkEo+n4jsIhpAYZ5Qr8yTbFjq19ylTtr0e9s+QTPSx0J0i
ZTgEVPazmIEaMwSbWjvHidulRT7pBjJrZ07ANUsjcQR4cmEbRfwKJgOxUcrV/5nr
FxDAK7dUbIBt6dHRZCiD8IOwFJEXiNrggjUktuilX3exhCcmVBOWQmr59tZ+ksp0
raECHV2IMP08sIpku194aPPA3ExVGYnGRypF7RSmftyqHEmKuwWdn+n5V2yANqGb
RkLIwboaVIo3EIUMsVUxhz7KW1H+zxvM4Yc/6krOkAO4PAN/DCzS+7w58s4dAt8v
KWu6F0kun9DmWKvujWrugeB4fJAZQ9lKxN32T2Wx/jiCETvrr7urNDaaKytB4ALK
orsD0clDYNSaVCwR9MXW4N2ThditH4S5Ct6mra3Fh++nsM5FxVzyB5HETcYn0xn2
i/LfDihsE2xAT5RXBYX4GJKe/cBoKhq/E5Nf+Rug2gGjR7n8LU37H/N/DfR7QJ4i
KA0HtC39Xw2GQbE0ihbP/ZjdxzJzXX6DUsKMKVg+y2TonME6Sbatr+qjCE7pBhrM
RfGKr386keigxCrh8AvXNdlWJ9SJ6nlwzeuSmYh6DJmxU/qTapP2QEN0xRfZngLl
iw5AolkurW5yItwWZhvGTfep0IXCJKGFW1fbofHAoaO7O2NxsACJCgQZjTRO3I+n
TU8rtgHYSTR0+wg0jpi8P1iE0EiXD0VdF2gV1+K1YrXbLmkcl+eNEbCq7QP9+phv
4XzCSfHrasTMowW4gCke1qXuXCn5OnyhfxmH4wKH4L7GIp/ten5Hnr8kx8x1DH5G
4rY2VbTwxlMdsVbCdg1ng8PxL0ToD4KDMoKpVGfi1Mb8+iVPJBTRLvTh8U2bwo80
0JzAed+U0CFZV/g2sgti9bBbfrWe2Op5wlWdk2uZjiKM1n424NJWX8RrmioLLM37
5BtP03gkmOjfjdS2Bc8oyU4tCk3Mf1GazPg16wi+z+CEqG4jYl/R2L6Je8K3Dml4
K0OXzppvwTHGQMoyuKmYDjUnBK4kUZes6qppugjIoq1RRtkjOp+Q9AzduoObCawx
30P/t2MEY0RBq6wZUwo7vGqxDH6H2FpzMvmSkDttBgPXA38PMge1Q9lrYuAx9hty
jVBpZODSM0+1J+MfsY2ue/IWYKNRhSqCVtFeMhoLwKC1dZC6vfkDddgJL326gQJu
rx24UlVspPdEFzopSQnLB6rX+7EVcPuZdBNmbiCzq11DkpyHEON2dQOF032Q9aum
s3RltHXTqnXTE9Gm3sXUQSCmhwanycAxRu8Q413LCsUWWkBS7lZo3PjzCKUEO5Y2
hGlUd/aPWyPPitTRXCDby4QsuXdeACe7S9awTJRZ74F1Gl2o2TdrLQXgvcls3qm0
v3vPHwhfUjR1W7jBufPEChFhSqBjKgzM+dTz3khDVFNv1gu8CMTB5iVZVZ7ep8nr
vC3+zONBcg8xQVKDV3bqo0oEtd6Z5wVP5tmdsltgI+dk8WGmHCPdXe3k4UkV/9Sm
vFWRzwt/I+HPIGFJg1fRRWW0b7Vk1f9WuBbf+eSjqfiiZK/Dz6j6P1jYVmXWzJeo
fVZHDqD0P8AvYlUxBbqWhn99Y4UKfRlVDv65GRhNvV1m3DtPlKJzt4T9p7tEY0LC
oy/tLVXsAqzFxoGk495FNpfYGx1uODhWy7XJXH00LimUFPpaUOQNX+rfifj4Vr0u
Lt0uDDJFZAt2i/+IeXKINJlXioldeXcC5ANkgUftwmcym16ivAL26VzM+C/TR0Hn
T8w+cp1EBeip6TWbbZ5kg2MTVWTl9EPBSAxnN++93WYOqNw5FccqIdM+H/ANJMVn
L5hIUmTwiborQoNYzEfyWcf9rPj66cMoBmCrrnASwF1kNkh2ikM76bGjRZiYrj43
F4OdBgXYQcG5RwzW3M4K6AjDrGHrT/yWeWgtCK/o803dVa8iUYFXQI4ImUPGnz1j
In6B/OzBsBQikXaejsyjmDGvD8vRRUSorkBypjNnbbppWx3r7LZPlNGmX3Vs0aQh
/7gcsildgGiblGj8M9I+PH0eC0/ROgpn7XUyOaIPO6G9Kf5Bw/NPwwrVE0Lsn4W6
JnV70kKJUoaEqVC0QWKsJ3GHiXDNT/ZlVfigOsvNA7xix1RFXYF3zk1IAFrzHhik
KkrN/Vk94H8qCWTovQo6U6Qi4vH/5UHIH+UyHWHSfQW3o94+DknYA/8X6id+vE/U
GELf9Ksj3gHpVDjdEYgdAx3VB8tue1ugDhjU1s0vZg0YVJXlg1pmXfXG8l5FPpVl
pIucfS6VBQjhaDmcMEQtwjxIzYiKT3zMOnWeyYvdiuSb8pEs/0MnA/5anCfX1Tq2
IQ2UfPzj0rsKJK60DJFGAz9lhqLcOzuJejCZTslUduJOVMMtSoEBKAYDYCvPWdL+
0q+oTgEmMp79IZ8Y5A9OHzSYddmeu3FIP7PJY2Sksas6ZJQ/1uIjgbcCdFOh27Bf
fT2R1z8rDntCkSbiqzb/O1ITg7Hct4JxlrHWAUuGDapCUT75uYs61hC8vBrdwmzG
ON++OeyOKJED6XJ34axj2+CYlN3/GsEuOhyhCfB9JOwD9mMVqOaW3oHo2nVBdqF1
A/GZw1qSc2SpOB1S2tn1PNSuYDllnEa2xVQr7v0u/XKaeRGy5xFtsw2wF1dUMcYh
IRJF+0z/OsYYyfv86B28f9crt/+HJ6PgyhQZHUYEd6X6M8xGLJXK5EjY3A+rdLfv
fb8WiIW3gIoUWLhcs4hO2pMON6B05hC36B4wwuGp67J/BxLRPXPMRsGXrApbArLA
oolI8mK0luFNujOHCP3V6+CwqIYwy0GERWm19tnsDzfHEPOIJxHlTSC/BDug7bDQ
LHmE5w59ejLQwSJilVgx4NhQ1UbKZQqxuTdt4FYjLRT3vPOd3xhvKkcs7jUk3Xix
gci3MvHkpnxti1HHxMWPVcSTafgRLH8284xNYfRGJh4clJ2aNZ/xQHfvidbbDi+4
r1X/cp4dPc9JaklG7DqpxlJC8xdoY7wrByQlMBvu08A0QHrZ9YQ7upydcHtYY5Sg
vIJ1XAPZ4Gndkv1OHyOpJPqOdvrq6DqVVW2nMxjUCM1+ai9uioi72pfPRA2zWzxw
0q5wMSIpjmlo2sBvSWTXtKD8qVb9BOVEJpT0js+6ii3J7RtYH8g5ZQgHjAYGR/LR
BS9F02yU3x//sD3aVHpVHHnVNOU1zftLhi907Hb7DkZ6KA5nzfbKliwPsEKQySkP
gSOt8JkK0yDERo+VDllcMkItf+ByUSCUmEiVQ5NjSj2Xh3Dw3v69WIUXOuXCHe2G
poOUw93KcY/Qp9PNTc6zKdJ/vf3ZGaAGK1Hd0WROiiuycrsXiDR2z93Qt9f7/51/
5yp0TBPK220WF5V0zk2mKj6UW72znb9q58EkiMM9sM6kANEBCjVx+bSS8gOPhw+y
WABu6FRkGFp9LltEOqNC3KxfCZEJ8ZYO1cn3Cm/AwPtrt0eE+xeS6Ig/W7pkuQvg
dqfiQy3rs0DdyHj6iAt+4JAqm3bdqimZiTZ7vwbyIfUVF3iIs+BWKNQpsNVIajlh
6MhbQgMhbaTSxsRuw5LTKJ8tIJx3PzbnTVHhHfVilyYxJDUAB3cGHynObkgCIBai
9DudTezuqcLvuf4tPezK4UC1RSnPrJoA3nCvDnJnsWSVxfTAs4agX22lsO0bsNfo
QY8arFnB7c0hIv23akSWSCrm5P9u+HnwpqMM5C6zNdTrHXAwcl7NBMbj8YrK9Umk
BVcits5hnUV9YQiJoD1vY4xsrS1isfF8b8YunWrevKW0C0lwjO1OPNHStBoUeAP2
qYOY6U7GaWTXQDm3s83ojoilN3BLgesTvlCSiDqqH2mwm93RT92p2sjqwVRYx1tr
gHvXVyn1Ys+nIns5jjmPuQLW4POtRfEIpmgHakALkfw8+Pytv69onkgCf8ZWt0+T
ehOXr6dLCjNTZzLL7c9Vk4ajha3dfyR8e+PdU1tajgwELiQpwNOEu+S//a34oY8o
f2fdzHzsUbNzfGpc+sjxakxFQlt87VF19vDQF2zymf3KGNyza6as5N75F8ImMfn5
E2LT03mfepe3wcOVK9ir3LDyddIdRQXFkYeZTr5Oj3zxbYL3FC6mC1ovQb9dIC47
BHQ4kwKxK4GaP2+xGZ0MnMO3V5ZZej8Q7gZE+fLy03068STm3CxY5wxRYsXhcNFR
w5UB4y2iYVJ91/DwtlPyzO81bY9dp3dqJ2dwa7N5bZfrFu7c5pInIEhJsa8y9iKv
qyWRldwtmrSIQ/J+GTVbLnb/MOTiHmhQWt4tV2ptTRByc/IsK0PXTjM0xdWoFSpI
uDpRf6tQEuBAdTbHsox2LzJHtlq8U5QJrJD6mmkSrjKeP4JIJjj1oFtGN1HTII41
LTxtSZaP7yAGd0hAVilOV3cXwwo+w24WzO+QtQKOa1OmbMnpke2JkAkUGahlm3y1
8KFHLg6t/AF6QeyNAG5daRfyjxUtSXvuXJA76ME+j3KsPz80VFn+UMICTZGQ9cA3
u3/UuyhvweM8qvwo7YHpDlcGAco07hQTgQIUhvbkDh/8buJqCtS3Ya6CIbaRhrmB
KWS6axz7dH61126/TZ/0Y47G4ipzgT7CJBnWTeGKc3nkRqV2pAPxwNrHEz9fU6p4
1W6PxnuNFv2zmtaDiRRlntBuoEhXUkynGH2gShsXJJmKA21ZitKA/PWUa1IbPX+Q
ex6QWw5WyMP2lr5rSNZVMm4r+hF8AuSx3eIVw4M2Ybl/oZ2PzunkZvIBasgPHERs
OfAOAaSGx+Pqmyg/YBWQ2gSLRzCIa9Csr9FYmXgMOhJNRn0GT6e1fdlGdElSqfZy
i2Tq+tTZtA45NL7a48aOdaFAVczZJfATIAefFqX6xdsg8QrBAt+xEpX/4pyvhoFx
L9TfADNg+G6E8tu6/Q0naVZrYSJ2juP02iUUbeEtgg1nFNBpdBM/hYnemgL0OJBd
ljy2iJ1Tf+ZiEkCyJZjBXmlQ5vGF513YAR4i5LO77fBEeanX9pHstel7RPlwUhzQ
A6/2ZnaSZ4S6BuhQSFwnngqmuOt4/PFsUiU30Z7e7DaWE/GvYiGKsEFhCCoJtz9a
HaZ2U3431kciLlUOF63i+kbq6BPE2hO688lXsfLptyv1kFCe50rDEoD0dFmYknlw
Wowtoyhe64eV+flj+tjJ/hs9eRlmdRWiZk76mLEwvnIQLns3SUgL4AQgQwKxaL90
V1X8/DjH8pWhWG0ah7Hvk9kq5nEZitkSdxQ5QSDyYqpLvtvnRf2A3SCthd3x6nGs
f0+JqOr8HzW6dXPf5FWGMfQnYrJ6mdbKPHGcY70OvTcEPrXe2ev+Y/minxIKceok
Fu43xRmr0M2eiisNA+VXkwKAqoIhq9xEffnnkHBMeJffK7LQsAD/vHPovG1h/DbL
wEPEmuvhBNeAWBwkP4Fbk/JFdH2pNOZ+EynsqSg9ZGa/5e3x3p7iuvF7RrTVrvr+
ZZVofp/AHvat+2fvVX7HgV/38T55PRyUNludbV0vxfKz64Lko9fBj+pxKduqSs0M
xjQ7kkA8x2SulWE/mo45eiQT4nud4Znn1Dhbbn9nny6dj5GvzIDZeZiRxoyKxQum
K4EM4vrRQ9TGE8q5z1ruESgNt0UCVJnM2aBLEGM4jTbFHhYlbMK2oLmFDJ0FHQv9
xmk3GU8v10XHoyEId5DBHiXo/WFm9E9/ihkP0xea0aTtIHaqTCqK+A36VrIUuLkR
S/NmCMyA5mbIu0Voiv2CQV0WSkf/+F1bYFfY0ayRcJ+ufPqnVMR5zL7thyMc4NT5
LxKZTikscwUyqqC4Gk9yyhcD50c+hn0r1X713vlZArzAH8s+8YI46EUqg5oN+y9f
ckLSXV7ksYllFXWDFZLLn+h2Ps9hqaLS80mAHUN5jUvYfaSyuNLNllS2JhI3trhG
sS3R0fB/al6ERwHffdjFPrVB4zWY3D6KjEgwalf+SrGqNAWmZdi1/ulalvKJtpSx
BQFxFJXU2yJXOyG96xrN7YnuY3vS+UEAI24ATddAcdJmTPc7nqC+910165C+kU2V
am823zLwLmYgcI0lG4Tv8rdUm5ilBBdDMAkLa2xSBSHlgBX4UNBarYmB52rw51F6
En+zl7GRyBBC97LC4Gr6FrzkTAtkZXwwiLBms4tt90eH6S5J2g8LLZR2S2Wr7ybv
XsPzoc7ZWmsb1VDlEGe+Q/isOBQwoscxqYrHbELeok+Q6a4zWpE+aBZS/AFAV3XS
jkX+9Lvte/J+zxQM/Ujc7CZ8oSWMlVVPKbSinBLCyqnZh9jW9yts7zh9plaCbWIf
IgoSgJKP9kR7dBOCmctkCBefNsIeAaKuok5U/7OsGiE/5u+cPpl9H0tlqAX7Amhu
MYp82q6Arr/7UsvdTjUs+OsnNX/cUZ57ERwGaGPwxL4b2JNECEginQKkNWa2L0HR
ysehRKnr0vR3fGC+uPsmR/cmTha3yg0NEWno1iVjhbhQkt6ap/3qcX3iid30PIJf
os7ZhLFDuclCFO2WfgJAa2me0zL4/1LzBMOKChybwiMA/LfdBN3GNhji6yOT7zjn
wdPUV1pfZpFKVqYhyfb+T2actPnX2rejeQfBIsZ5mLJrvMGkGLRcArrpHwqJ0F1u
MPrRAncwNsPTLy9Gz1lw9z6jHPzKYQ3ScDtfLcBoU9CGG/wvsNGrWFehda0dJbEJ
xixnf7VfslgSwyonRd02lvkRBdWbdnzbezz6qwznHPVh+4XJB1JOuED/URNMOXER
V6M8Iq69Vq4FCFOIBMr4rJNoEiMXTxNHdiQ645Ie1DgUabElQGIQ/EfMbgsKeINS
PzH1mMNNmD52jrzHrbbIFrEf/uKA0ww0S5gQ9o2U08l/8Iq0WTznh9txouzmOBHV
ZOpLy1XBG7eqcnzWv0jwnJtSAjA4mev26rl7gPdvP/Nscyj/jdjRVzWXPsA5rHhY
qOmTECgRSjULlf0ejrhTefDb7PVBJsjQ2qOYI4xecLidJ8QSC7vtkJm2f/7F0Uu8
RKQ2YeCbEXGCZM3FSmkMonPzJWitFKXuEmTNNDY6iXR7JH5RDs/5F+cTycLjOocA
fIahTxVIcT76+zKYnLWEtLkzVNTO63GDDP1jk4kwsCLXOWz2pw2TNU/fEJke9GHn
rTCxiobceiV9ZHt/1zpit5Evofhd7hUpmAxm0XrRJ7/OStMQAUwIiLXmrGe3gK9v
FfeMN2pVPkHSBUUzSD1h1kSo4kQS7QrAGDKn3B8eFwXPVvxTg9RKohzwxZ5D2Y2z
hzTa5XNXgb8cHOJ36lYXsc5TxvX9EOcykUriGTGLnSDI7h7bqAz8ai/K5C9Bdm9J
oU/cQJZKobgibvIvpsmvcqIlNw5wKWJVMTVIoWqwTqr997HiUaGl0oOKlDbcTwza
GfkTHiO2vdlBqeqygQmZPqeCNSuOKr+/MYoUuI+H5ttxyde+H2c4BPccTylHZBfu
b0mCnJa9Cp38V4KOItR3tQp04NI3ZDeftzfSAdga+UlD5oRdPgw/wl8ldedbu5NY
WTEMUT88CSxWn/Aj2EnVz6CmbcqCq5lh8Y7xV4lTiPXDvPPTRUv5VG0ZPAC3epPv
dKwhyeKAaQQwQothqbOi0YmOAgkMo1+Zv5qnLIPBYb4pu9CYrFhR6HHrTHXfNzJ6
bK9OzNSVJPNLgBHymvzKhY5KBPGcjWa8IuhTPbv9qVFyzf3+dMTNaoz8+IznPd4t
171WEPhd+WCcm83wir1QpKy0+omv3pyf8jr5U3qnxDnsPFlKWA9k6r+/x2hngu6I
13bTeJckYtE2MUhoNYOvKC9J13zIZaijXVZDd5jkVX90fZ6ce4/XYxgIZX+dKM86
iUh72d1ELXeLuRDyZHXMzjlC64AoCX/7ZxCKRfekiTTs73KyGwWw/61VpPxhZVEL
H/vn7loKEU6dVnQSDDJR2yd9fMxUg17/arN1zsZl0wzZnmsPOAiT25fsszXpeR2k
4ahn2t7N2uCKiWnuCkic/7WLwuv4GQTwhv6rlzdkM4luJJbdLy+gmFD6ntNz0h0w
NILqRnr6r5HNzM+8ZzKPq+cpEcZMPwjqcirmZxjuymIT1Si375EiND7ArhJ+Li1l
9Q/NPHd9nV8O2iUXG0JkjWRs6LIHd0RcRX1QJEYFmJ+sxqa7MbgJioiJQMTovwYm
8Ej7G7HGK0XYkHzl6sLDRxTd66Z7Jf458CTtlO5WT+Y=
`protect END_PROTECTED
