`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Xk2CD3gvbpJVWL5StPjjtwQv1pz494q9A1wObg+P95o25yhyrpKFG1d4tRHfz6h
whidd7ww8yWcauqla0/2TaZxZ42ukQItQFSp/EVGi7PV61piL1FDN89Yrwi2BJKB
PJYILtOzIBTviVzz5eR7iAGYqRO3Vvwd/wIovJ+7nTbRzRoMXjYHU9P6p5SpF/dh
TXkVZHPHXY63CZlVmRgx6v6mpncEZGZkKNEevpuf9ox1GrIJPFFUFU1HcY9eYbMV
zZJOor1JBvgijLFyZc2X0VaSpEkQqz9SwPk8EP8x+66eOfKAhTZ2gwkeMgPsZ4uO
a91sntluEvthLWCtElHtfSEswCjYi2G7sHRDlz8w5z0dwIGbWWFQxLxRUKHzlD2b
04TmDY+TbTJsjHWGN0YI8bt9Vmx1x2Zn7LX6tRhDIFF0c4p7+KlPDPlE3+bZvkw+
x5Ge8bTYPRzl0J+SZ1EmuDTpwEwx349TzF7Zrj4SH8xCsJcfF0MDn+P6JBEu3ra9
MDsN2PrSFSvKd6CLtbHmqBAbidG2vmqx3IgBxw5esiJrG+pYPsHv3PJtQwk8xD+B
jQJYYO0p775+kqE9uv7G/Q6z6QlAgmeIzZcLqrLM8Ehy1Gaqq+6fgsUIpS9ESF8q
EQ5SVJk5kTY2pSCrBgQAtpCJ6GV6m6faRyi7X63Es+QzazRva2gEg4vT88FWcmwz
L/nAigTGcNcQ8GxgEfgX6qfN/eZ2GXU8DoAozHHnb+9ShIJUOepl+ZxuS6Op07+z
Kggc9lHhCWqaE8AuzQ1WTCkaLq247CJ2Cl6C4ct/iOAVaO6NX2fJkWIj4WCllviE
/YUD3fR0eCszghq6dz3l0QMCvN4x9l0x+LJPriJbvweygK9Nr1sKaWh8O+0m/DA7
YowfBacQnZIya5Lbo0QdnoHkQLMZevszsNurYrhOTtDmULGtcLLpoyUg6JB8Z+t6
kH7YCUB/kLxOKmh7Gypeue9LrtUOiIQYZXfqI58lbzdCyc1mQ8SSpmXJ21PyKMWJ
ou0wQz38L3vWrJKI59IIennY8W97zlcBxpj1Ef60GCOrh0zW2YbmWYowkT0Z36zM
GFHnmqsoAVgdnAXzszExVUD+Sccvn42jkdb85OROQSUqKCuyxRJAJ4tNXvrrrqkm
PmE+efcP3zKs9vmmsgPCvnmNNQv1qJIcZhbI+BkZWo9Ixiy2FmTiTieP7hRUOMjE
F9H8cGRZnX8Lys40QW/lG6K27wD4B2shePoAbJ34yoD6k4I8LQ4L5GZGA+czzfAe
yI0XbVMNsNu6Ko7BqbwiA7RcrTKPR6wsXTrn7tZwcu3mYkigrAxaDlFqO/3ASdL3
8sGt2jPlsX2KJaK0yIkKA9TjA0FfSTKQjtiQ5XmXUm6Z/lMx96ZKUxcc33i4VRkt
3rkvwoyL7u5FUbinxfdRHL00yWvM0zZ+5GVIJjpd9tnEeoRrYhUfRG5slzPS3368
mwokBxadeZwIH3QJ/NpdMH4YsDTcZ5ABz/WnOSrOAsPUpTtKilbFz43XoCYufRbO
lJ+AlEwlVMG4WiHK2uE7fXwvhsrvw+fNCAqz99ovvyd/91ERWL/gLzOa+d1vrRG9
dnAmjPPhgKB8cVB2zF01eOY/YPNjN/IrpGZp74VYsFoXk7VBYhHGWIQir9kBh8p0
6eaN4L3DRp7kCvH/8dyxhOKWzB6cBd06Gj0iTA9JzEWM+sCvECGYw8EDwZpW5x/W
35RuGfdKA6TDLS2xMJjufiyZjWYywo/ncseNiWFd9NcmZ43+4NTycS/roHBB/f10
+H/XmS5zfDIcrRrwDPG9YbbNOUtRjv/Eaw2o6cgqZH0i/BRm7RY0eQ0vbpqTXOlF
+HxSyqqRQ4Vnio3Ae0QONI6jYyG2tFjS9SQmtxcGoxsJaX0zuQEliaV8UNmfFI72
teN3yPRzmmiNDDO1c7UhN40Ok5fd+MMwbQvDY8z0cmb4DtFsMtMHiFBfWyacXo0C
nCxP98OTx2GXvUfSHjBSNSMq4DID3KRMYAjOGnszErnqhzk1nEB6ahYJzAumP3By
vmUIavDpjRGIrpd7GoKOT2LdcGrfWgvxLvwGX1FOeGVxW+zkwIW2BtE5AVhXw90H
GbU4Hy3pIJqiE/rLKJHh1NrtdFkEvq5KjfdGihg2HmNmAm30tbaKq8WNR1DRu0VW
6ea9+7MD7Ui0gEpQiQDEhhc3CFMh6AYbpppqoElvowm7g/15kMM3DKQDfGuKDpFP
xdzvQoz1ceykx2g3MKsq9pIWn3PDX00WO5Mx8QTpa57dMR/2EklxXyY/BxGe8Xus
50kznmST3+QeyfJhc1Z3hb3Iq5zqbUC19gs3OySSeFtOnBE/lfdFuPK+A1tn7oBy
uWbl8bF7qY/eeNyj4sXzeR8rMSMBRpcLKV2TO0McJIuR8zkuuHgYROLqgyJZEemF
uqB42vHbDSZ/2vQDDwgNHy2VkuDjEK4dJMT51lzBZNVSfeAtsYJ9zfsxQLq2CIEv
jAqC6Y34gP2lOa3Js5PBQZqO+5i6n1wxrSv+5jXdy1p+Wygg6KjofQng0wXyvzWs
pa7vWhSPxrKoR7my0D+Ynkl8h8jvmzYdoK4bW+0uQ40d6la9edETboGWuc+fgX+M
q5SEXy82moCRrrTrTbQPJ9LugXr7rV+BZEkpaGkhcmyLpmyx3RjM0WYqKFUvXLdA
MIeAWkdv5DmgXHRjN7pf/h9I2qOLrL70tBW0r8Oku/aqG5YoPd8Ac49StpnqJ5eh
In9dJQIO8N6mXnhUtj40ewiwH1Oy5fdtzztnF1cyGFAWu+x8dSYwvxYsUXUwnsO2
6x/C8gJ/g2LjlR3nCGfY1RpOr0ABhWtJ+NZFV1MGVjN0YQ3cQZJ/6TPqYBschSio
5cbw1o160wZzqHC1QlwBqtxjyAO2OFQAs9tQa6oPN/ibMxZZpR2ayM96cq8l8xFu
9p4hMTe196Fnguk/JsHSyjbQt6h4FrmrkgvwR5CFFP/bhfLikTLvXiVTy9lp7Jlj
FEjUbAYl1pEpRlBOTuZoZ4yzMbUF/LceZPc+KeZu9aSX5E/nAalWKeIqFCZ50MJb
JCCEwiWC5x9OXXEG3FWDUWZR4vZ4vG/xX1GoUqb4iFWLiKR/QVY2Y6C81V5NzmnT
PvlWsgWE8m1yalA5o4M4Yu8OP8XWHuSaGzvGs4CPWWAyvao77YYmf3+ZGhRajC/z
wSdAPDDther3PNSQ3aUf1eHpTXgI1oZMMKPAw1MLKXyAHdnlQQL15XEclc62AStA
BaK6rNNhmDNe2Y/5TrQJEA7pV/JGtmk2k62xK2LuGZ8PaghRRPpbOEZT0yRZqdHh
UylL+2KCF4d/9Pf5M23uUOr8CR8BJmtP2kwtiTG2+BH0j1X8yZ8iKz9BsbXN8KNl
jEUyaSn0Jhr66M8KQBeT+a91/9wVfsARYh5j8yPE8v0+Kx9Z0FQAEqLQIHY9VQWC
4GPlbQqcwVWMhSocMN2UZmtBD/j7UM9c1O3kIwFOZFfTqOy4DharBHge15PL4iu6
/iD+wU2flO3VDV/54vDVfw16u7Rq8nO09G+Iekk09MyHT+pUKwgIJA13dIenNZdw
rUMeZ44xILTorsKTGHKifWunBF0trQvqQzC4Ut7zY6MgQ33Q+7Pm8y8ntn1fTk+Z
1vuSqNKLWiaqTmR/kKaXR9V09h1Yij8wNEN4NqjbQG5uAGGkWi4LG1SSZvjm6ZKO
FBcqb/j9FTjHHcf8zh0fy73424oizz1tREQ4aybUHMbzYrHTrqK2jAqSXSrSYUx4
y0P1a6iBFbhvE5ODZvEhDnE7cdw5/7hK2qUtu4A2AzSgEQdnyt7aWxzByShRjx5c
DvosQ9JoekDZuqepf1F1QMs53U0lpmt4Xl2liI7eJQSvODPxecWJB9Kym69+FMuM
gAxthY+pP8rVu6k0SwgHsMEEFKS+LpRn8YBVHHr/1Pl8eITAgOUnsHtH84OVl+bi
d6XtV/8ESLGNXmJAFTmaf/Wd9yLCGIG1ElwJ99Nk22J9iD3Cxz2zGjABhgYJ0474
sUnNn4q7oaAyR7jezaoLJyc7GxyFTbDW0DtuNs97uuw2EPbE/Y2muQ6Ifsp+5V9d
7+cpyVmHH7NnMkFkU0RPktZGpeEmHGO4vuXV80TmJOC+WVaHhE63lONy6FK7xWZM
y8jmiG+qt6Eh38aXkji54neqjnkg6j70o3Q8pEt1wWnKkoSUo4NGv1IANUJlAaHq
37XvUtivBVW9wifFnefc/zoMh+vB4xCNPoe3aSR3yX0/farMSA3jdHbIBis9Ewpi
lBxNxGvoKjPSbVHz3CUszk3NRtqeEColXilz/siF+gh8nnhZjHGtzbJ0rSlg2vHk
j6wHtSQzsj6fF/CIJBBiF4HIJRaOo81MbsP5JFHAw4E7WS/mkfKTCXzGq0n/meXI
krKtcSzMAXTEXxsWtvjom1KEBSLf/+zvcKG1nlDBFT7drvjjpVOCPH0+U9uPNn9H
jXW/F5/SmNvxaDd8f3CkX7WURl5rgt7pojUE0BcErjZf3PZkJ6HyCywqbgEsxs4+
I+avvo9bYsalD16A6raFUYYhHvZ5wGMV5lWcqBrwupP/1wkb1zqfXykeR+rrtYPw
ImFNFB/9saWGxfEj1eo1OmlcSDXIW13ZYpyAlcnvT70YhBddrYlHydX4UEs60Imq
5+nL7eY7LSqqvCEM+hAaZiR3uJPRhv3cHlWFNUa7ccCm0ywYrQlyBmX3mKXbU1tc
mt5MFcKhWPfKTl8FLZp7L+WL8PapxtSTRvs4b5gBpRYxPYx9kojDitzs6sgan8H8
Trt65fHuakZ2+yuOyWSfeuS13I68FwkV0qYz6FnH9B9T86iz1UrTEKPGGV3bvav4
vqFb/Y58Le35sJGMKjn3FnRJqcadJNznnA1+KzMzqKxGkrsAQE5Rk2gP1rfRv6sj
Q/MPprU0CjwRMQpd1AV1YhetwAdqGEYtOA0d+ZERRWp/a1AV++06w3uV4YFnH3Xh
djrRu/jNl2onnZRZYz7JbEnCQzhQPgXMus2NzpiPiKUKvqroSjj/3uwV25JjQcEa
76Vycr5vLXeu5vP1WL20/37Axy4BPd0SjxjCo2qnboqMTh1Ds9/jQE4SBVCrhzXH
UOfmELDytNGzJvNQ4ssiUxAGEnQ7qYqbQ1g9GyiPkIB883Lk/X9sBDqV6i5nlbl6
81nEeTzGG/XLoyoZV+UVR1vf/HxNQSa0wPp3+1GQkqANoaEMSkxL/tEvudhL2iEy
0ILGkpakglCuaO7u10mpAWiVaoMLKKhBdz7YYn3AJJSxrRF5UyQgjcEVsRoju7Kw
MfBm44DgYZAw9fCRyjP3fA6PzO5WTudmlPg7m775lb4f6UBOckbVDjD6vR6JXAXd
c/rpJVOwws+RMVlmNK4wUkqwYntJtDf8ZpKj/Rlx8yrlw8gTSJSv630Fy5wBNLEh
XoLouYWcqbyqPOHZvSZV7zaBjVa+g5ExyDZdcgUSZtFAaWDyezfWfcnP4lO0nmJv
eXiv36i+faI1xUJeTP2M0KhwA2uEYYANYjghKcwnEgf3c+MIrjD97ZFPUgP6Egoi
Xo0NXFRz+hbxCGkotZzcNwTX928gyESi7uytYZUunqCvz8I4AlQfNsxdWL5JYo68
jGuNR4oqdXIflWgTSrhApnhIZ/igToyzyQdcwJ6QCJtR74V2XP+E5TZQmomTG4ix
1eu9964Hc37znpQVxTuX6XNuIJvcW14z0TaypOVax2FLxAfDFJ0UGdwnx9QWPCYJ
Uf4TY+8KHYCoVj/Bhw4eICqCWdFuX63jC5JmC1S3wEtCkngpS18X7B9ds4Wp0ySY
pdGyhvLzRhQuz7XYyl6cN1SiymLskgUTcn8ZIqfHDhPooFx/Us9ygoMZk5kf1jmr
I6VUYlveiB8V0AXCA+GDZxbmhNEqpUjNSiad3rpzbmHm4uKNC+6vCwgPRGcoW8/n
4YEc1hYpWfsInHgN0qqSMy7zqqjOwrIR+kFLbpG1XFU0M4Ut962eKbF65aPJe2XB
M+p/8ny748+Wk2Ca4fWiC490F+ho93frPrtV0TqDYd2rWyX2PD8OZ0feUZvbDNHn
RMsFxsB8QH/e57s2j5WZm23Ke0EIgD3/XzHowsAafe18pVQJEHB396gtNrA8hU+K
cjGZ/Dois9SNGq3wPwwJNrROLMupAYYyUp6bW9enGq5IHVLpSuDKpoPg61JIqQ+H
25mWGmyUPmGvLoyWTnkDpsZpiM/XlWTtwzaAqIrIyC3mPzrFA1Q6CLo15FfVEvBO
t11YehVrsrBOjGvSvvEtkqrsIe7pkzuedd5MCSXcV06U7uQdntTY3RI4O305uUxf
p4sCeBkwhXeF28E0/24L55FB42u8prIKv8+jWhf1F2uJGtbYtLTVEM54TIVZMB3z
YgmXpAv4hucv9fH4jtX3QXUIbZ31JN7S7JwciMiFikm2kIDUL8CPgyJ4ximp+eql
oHJhRU3ACKynRan/cEXxfe41nATRDLgV240dSW8qMXhZxsh19u7DodeJ19bzxEh8
RBqptBjI2Xym+O8iVSbgskJw3+omYJ6ERWu3xm4H22amLvlHVLTDacjd6VzpodtF
NJriEVV3cNF3h3+8GCeBwC8RnZYhiwhPpOAeySD8t2wWG8tjzL2YTiOUUHcRfRjo
tfMyp97U7QT6lKgGcCoX5XTpRLd5ES7W7FxrTo35APsGmgfw9mKJ/o7VY5rLlaY0
vtA44RszxbUl7Yy5xfgkaF7y/yrSjHFXPq4AAmreJzKJ1I8T1PYNlSRXFNXKpjm6
l50K15et4pagJdsboJxuaxitCH7iwEDOxQs743OGZ2vTNM5YFTfC5/27nIjJEQBP
KmeIWSYc7fvnek3UrL/UV4fBIh02oosNlPAta2/qiTpRq7ffSFvhcOPcvo/eskFD
4PI8T5/ZsC8yl+eW4yfogtyt/v/YzjL53jr0zhpHkzfTbdC00KdNl6CNM/ajwLHf
yTgp/RoMk+6xZ06bwMd8ybZt6bxKxaaz0WyyZi0frPswwcb8CTF7xQPn4KmIMVyU
jB8QZelf/dvg0ZXfPaCsZAz6v0HXBY0rIe/7VP0hrhoJQKAWEmxCX4Gmzl89aSdb
zyJ+OClZ7+qioZ1HvqUOCSV5cpSs575b1ugFHkrapp77HQinRnBCFnxunyG7xeAs
yOLUPo/onRFn9F7/sjRlV2Z7C2KyOZxunMXuPtMTl/fS7TjFNJw8OGUHG22v007q
x4Aw3JiNzUxmfZnEK2z7+feYmPq+Dcg9eWO2ZEbtLHotGrqh0Sfq1pXdDIO9yyS7
uW4tYOMaxGFol1zQNs2aK4p4Lvflwm8QpVW1znorwxNZLaSPOo80u0wdi9d2j73F
kTLCZDaecokLA8jwzvPmV2DvmX5JXr8LhtPYCeVPpt3wQEpk0Ze3+Q+Mp4RcmBBN
zacFT70HRum6ee9SMpSMyUI5SXmDSiuzXfGOj9sw/Rj64aY7AsBEsnytFmo3/c/u
4azlXpgy1KnI/+V98UbrqyS/UQNZ/34ncL8OBQvv4bo8PKERzdGmYa2ftajCJIn4
pF587CcK90+spCN4DwHT/My/8IXbv8xCFwY/giNlq2tA74DnN0z3/K56uJmjcLq5
5SUxtTsbQPtFsMX5n9lcJrGVhEOAzVwfRt7uxt/9Z02Th1SGiphoL40mFg0ulbBD
CD4Omol3O55WM3fpGOLRJ1cYA9PgjdBtB71nHuEctReuwcFwxW8ayiDs+WH579OH
90hbJfiCX3aWuRWrpuq/k2Pl3IROkWrzVKv8uTQi1908MQGiNb6PWu2W/tT72DHM
Lmjm5Xg+pi02fiLrVdM+zMmsi4zCEcVeOAbWOU0Imoe75zAtbqrHKMwpXpmD5X/X
517nMO8tP+QQAIXzPmMSqXh3oYBYEN1XWqil037Y5EkGWsS7cXoOxpz050Y1RLx0
lTzlbjpcwj8cSl0LY1ZshcJZXOGoglL/kPuuRf/Ruowj/aFXjHKuDfp4zlOtyxwe
LTub9r8K3UooC4FCUAVkexIyJ573ZuCWiDXkxLHwy2+OGzuKm/c5qW1hz3NNEeiS
O+yN4s8gVv7Ab6JOYYLMqdD0o8Lg7z49ip6CHtcdmgsN6eCYiGccTTK6QzruouPE
oVY7i8aJydswpgROXJwCWJqfGmij2co/1/CDPKwUJ0iQq8RrHLp1gt/zGWHNtNwv
y0UG3SK6RTun9eQp3+HbVjdnL/HLuEmjCSpcMvaVh/xyFYWzy7/4xHC73fUfGO4X
OdX3niL34YW4Nmw/ZZlL6sEJaECCAFeiIBx5eq8FP4FQP+HMwiofyyhSQvuryP71
eIHmaf0/e6QgPvoEPeUxHzctbiO5VfZqyqie0OnYl1hjAlKTAmeCjog7xFfVnLNl
bhJT4gT76Ob5nF0/KpX1VVsYqyUkw//1q2WDgyHQeXdVA3PwMBOeZrdKCDoSS6JY
9lKrtTeciAFAbTz9SY2q4mF0lh7x1+s+8n/FhzqQafGvSqi30S1wZm5/vi4jf/+L
rggw1hGOwxysspV6Oiy1ePSYej+IBylh1l8MmnVmFoLL9ChUi1TD00yGfG3TIC9s
brRpHgDne4jHIs4F8v0slC+EYNapjfmcuaDPh88DhkmCWsCMBHUmSzd0gQFgbEW+
LXVsilk3KlqKOcGqR8jpEKCBOGpRGmE3gafzeIOdiMMDadmR3b4k4KlMsR1ma73N
JQFNXl8pL+Kj9XGs7BJIpYI5nH6ddHyDvwGvAqXazbcR7g2aiJMrqCSHAmd3VuKT
6ExbpMq2Og027v6sJeSfb5yH7VlG2fMfDi7583EbG64fsL/aqixn8EpMEafThj9i
1psDOjl5ebfv23Hwmzr+xoRPD3vRHCeY5/JzMNHtwwivYaNld8jCpgJnCaI5mp3a
lGPO+/eCMuJdb5+aE+73NSQ9g9kkIzSaGFoquL2LeuFiZ4vqyB70a6IV54Jbg361
KJWRl9XClDP8Up+I+z97vWjjXucMGaeANemgCwkNRdJvfRHQHYSBzkxF9peQm0+K
geH8fd07wwc97sElZbpo6kZSsK16pmpTZGpnDP4b8Z53awze5mVOZf5EOnea1cTZ
Oe2vsj3xidyJDzddhIHynSqpizK1mEwLVAcwGVEFjQ/yQJcT79tkyb9bnYQcbCA/
y/lRP+hzHiofUcliJg+OwfUK5pKJDB0xs3M7pHmXaBjaZlzFkFuCECeU3+t0eDFQ
II3sm3emmuhpPOH6624U+3WYCQiQMkCDwAH8LGKTlF2Xs2kPbp3aKGJ+5WD/bSRo
fZUj3R33IT3Pqdf/NnriGhnT1Sl4EqwAKXpgr8Fkl3DxiWt1up4Umvpg3/F0a6f/
08x6D0IgD0Hvn+Ng9Y8rxeqYmrOAj0n7JMml45hRu8KGF35or2JwN2YTbvRvQneb
yy7rPjdQ6UOvvP/i5keaUovzb6ewqYmr3ccs/jll03we74LQna5bwVeBJnLF1a8U
ETYw1ZfLl3zBurV5QGNKxBgcTuPaLXC/4b9z6XuBsCSCyZmtbg7xXeQLhxbOjjXp
ibiB8A5wyC+mvhDmTmTAKCDP/az5Lw6M2mhXm0eFq/+mmVF18Xvs8WfKxZmPW8YU
x4LjWuTgo9vIHkRSpGkUyQCe4xEsfI7bJ3xTf6oAkyxZdk02jYJ5oxOCAm6CI1lh
fqmOULNPAB+QzQquI5/W4p3tqRzfF14OtpKb1Ic9eLQnGtc2XY++IVsvAgLL4wu2
XZ+J7ulrFfHCC7wmPH3n4xboUIIqOu1xqVJremXHvp94ttHrzHgGQohGn4msSOb5
H/jkOYJi6ZNwPPj9853g79zv3w7gSfRH6LDL95yoNREA6PctOkNQC8jg/Dj2B6hl
fKywsRP6Dp/yDlbNlFlCBZxJBZculOngWf38t/Z0yOvrfFlgxPSWHhktgcObgr3X
sUAAc+Z5ikwxddFxgh3xDQ82sfkBa8rSTABtK+W8SLKOXSIXqCbRoumEpa/16pgS
2Js72cvLPfZV+auUSQj+bQkH9fYiujKHiVMQsWFh/30051jGjZn6NKMNW6lhf1xk
87awzwFYHtNGCs9cEeaLo/Bc8nZo1dkpcAzCHArieuIMyRXOIffEzjexcK31nPaj
wTGFWAJpFl60UqFcnFenMyZpF+6QjFZ41k7qAN8xckjDTOyM9mQq3rNTTV/qjYSs
vzsNi1tmx7FgQNYaMyGAakV3zwbpWVbC95y6+nFz88/hYloaA8PBNli7tPSymHXy
SBua9zqoAGDYtY6Lki8aBWMVg4qdrkicS0pzKuOYvV/bGDYOhUezPYufnzRMeOx8
gYHmE/sziUtmrCbm6YkM1+wQkUaB1+7aOUcdFTvAWNQ7gpyMb3j/rpAwqCygaUxc
Aib+vsumh4GtHXyoMoVEQyb4GWjgmUMVNEBtFzvU2+GeTs3y7kYDHCjagyyLxH4L
AR9gG9OhwAWCVlIE7tNVF/kX9qN48uMvedZTqtnEP/Cj1wncJlMpNOA0v9asnCcp
l+5mfdLWYBLM3zIPmCbt6sWPuq9FYUPozc1io9gRAM0g5eDTDJqQrBz5/KMNz7Vc
2E6+7sT1ah+0kNeSUXngunwkFnq4FTuM4g07HSNUijbTXiCMnQ6R9PJENJOJfu8i
3KVMkVM337sWgRgvbH4CmrDeeIWwuJkIndleE6zFIxpN4JFD6TYtYtXZz4VHkalQ
92isoucxTGfhSk7eBAD4TK8UPAThnMuqC0MIvWM4EcTWmTxOOaBV6e2jG/pb7UnY
uphGughfKO5lTGZMUbHP/uvwg7S1WREaljTXCxyCKFXlN9mArtzWHb/cAmlFXzTr
bX+vACklrtH9wSq5VLVGQmCmwYhTxp/2UVXGhTWrcZl+IZDE79Jyt0LJyBUIrLJP
j2zrZncvY5TmtQkLmBTn9XSBAWvA8YYUeGau417C8qDelvdQXCyI+B1uULHoi4Qo
nmNc/VsLc8AOcxreizp4EEA5uIqO6aw6erS3BWzHgjC/f8DoPbRr0ZkzIwmqH/en
5K20UxOgvBEhjx/ow5n9QG1Oc/EMMea6OdzKdeRAiOrqzsyLRRxUeBWuQ6M7DuA9
cHLI41bGzlHqNWEhP1AA37n44Ie431ZnBS1m52xVxas8N+9KnDywWLc5RiNK+SEN
b+QGN8cID14DGJe4o16voYY+RAlM+Qy7lQFHcwzPejkOyVNGpLGqXd3pPue1uv5N
2Djd49QNedzUT/1MFqgLKFYAsf189CyvetW819pD1xr62dYw15WrWHlIXnZG7ZsH
V/pdJznCUaSPE2+BuuHclW+tTh1OaU2zfA7YPWYTb1LAwZdejJbnbfuM8fiKB2zI
fgy8pnDXOYO3Bu7XT+RXjjuz4cWg/QAAUPONxzuLYP9r3MsoXRqL6Zpzczp679lv
D88T96ngg57ndAC6Ib4h/WRh1fvRD64kn+3PXeC45Phq6VJauClbbgtq5qyVDwXR
pN7L3yjL13etSf6Zw3fE3flZJKWTfTbQVcDCMAcCay+s3DjLkBRwNT1d/M3M5DKE
aqiueWRhJVgxgKWftC876toNKFTjjHFpx2ISxA/UufTtKOk3ecehFTAenapuz8DP
04jA1K0ArOyx8RIm2x9CPdf4EGMQYMvmTTFtiHTsJ41cDZiHQu1PYOvQhg8rV0mj
1cx220gV5fhzTYqYuUq0DcZg+DVGUqTPPiWMj7e8Tur2DxSHwJxD8IU9ykBQPTM9
sm/FYqZNswyp77D+meNpgVuGZnX+0ag5w6TSWVkUJo7hDeY7ixXeuVvgWEauhTpj
agniQgonv8WQb4C0ycXf76F8r3pZdRCtlWhEGjxYMUf53wJhkUnhL+LtIIqXDIhL
nBhBJWwcqZEQsoH9lTM/9uO9gNSN6kYkCb+q34Vo0hiSJOxo1k5UwJzjmj/J9xpU
TKmHw5/kVlDMSQwhnsKsA44YFGkAwj3KM2Qo9i7mVenZ1XIdmRhi4rLuilIDYq+w
Xi5M5Cq12kskqUbPGM7jyardMtfUUXsfiakhnfVw0OfQcysjd8vZ8BoOSCUNOB46
ssHGodBfcryypGqWEL5PzQxJXLcyoIaZyvjJ43vQvTTc1RgirpiuohUx/wkPr7EM
QaNjDtk/JJbi2RL2vqeyLT0tYGlJdaADtxU6FJ25JZUObzN2mbQJ16rjyK3B0Y2i
AjfkHv7ltg2J4n09l2iS+f5uS/xFTSeqzEIiVOUEsjUInI/AZb1fJ9uC+mkqT4VC
vMbEsqdUZqxG0duYLqJ3JEaRWo0Vcq9pxeOJ8Ba5nsDdzwjPmIOpUar6x1h0l5cY
6BIw7SPdKYU7H7JwZadWYiq4RS7hxDyHyyQcQpALEDEfHO9IvZIsyhFvjO2nJicT
SyVa0i2XQ+PuMZEOVo1hjClJKcTUeaLKnEsyouPlUGlb2RjTpj3i4z51Kt52rSyt
Evnwc0eMwmaD4SL6ES/IhVLB/qF8Bk3sum8Wzq2g2XCbtSxslcdhlBD6QJ3I4ysP
omoriUYEGKNwqP4Kfoe5Emgqm2i+Ihnk920ignc7r0svO/+12eaJp5qkrR1RSAFX
lEAA2KZ9dIX9HMjRdNuLZ2G4k+WMMlGLlxYXY1QcaOPSkIa2fFVfS5zSa8BzAjii
ky4rtIGDlfOTPVON1lRXZlPA2rKTwZ7gZWT+A5j15cEvI6hG8cdk7O7p2AGS74hv
5fcw+nq/+HMM27akj9c5SEQ0/tQk06O+4vqPgRe8nkv+vLC7srRBKtWNIbIaVHtX
vBTShA+NNCVbR5iyy0P9ERPyP134ighchMDRRSb7LaC5iOq60QkPsmb3v4EMofj/
HpciYIGFIlihdN/PihSXY2zA7o/0QGx0FkzzGNnymzGii9tYiTkA0SyzEOEf+axm
v1FXNdyfQU8A5QCZ6An24xtMBhfqWVZSDrw8nZ7Ek6eRdWiDWDqJ1HMN19z5q5Jm
5b8I/aJ7zkvDbnrcWT112vRsyGEBJpJ2DkCp2BwerFLqejT35b6VYHWbe52E6FAP
aeby79eCzRdTbIAg01sSKoKQSaKmjWSf32u19dRBec5fAXfuOvs5kJNjRniCSn+O
j5hnik7kULCfJLVUcv23wcoC4MqMd5SSQ+iYkgcj9+qvAtYWCelEUEaISW2PHkQm
KNvBy9SKb3mFuzCWWFaVfGkBrMxbr+PVP/0HpAE9GY0chRlnFrsqKH21JVUwJcrW
2GzgBv2Og5AixFgu6OVdhTNjKMShGpWBtOSvbciGMuVjh6qvNQAWiBO34urflIsg
Oz7UDXCEIKdG1BDkCsdtj3xQ+JImCtx33vZwVbOzSK7iasSxL3HKHBV5D6x1kwd+
`protect END_PROTECTED
