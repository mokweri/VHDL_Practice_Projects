`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkStxjC5e1T3ek5nBa3SE2wiE7sMYsjthTbc4t5NHWwHnCvZrQ6ZZGkx6S5aYlqc
/Pxblzsvx3Ee4IyxSwz62G4Fdrq7vM4CdWJy9+2J5PHRgI7eFnKzXgHW3lQ9+g2a
sb5u2RNLtzfT5Oq3qJrompdiCII8KzWzyIoGZgOyHxd+4w+Ewy+Yp+GkzEixh+PR
6velPA9nivxfrVCvMUznpBHrxFKdj/jgCrDLXb2uOCsoRyEHYUICtnRe552R6uoV
JzE0X/QmSJCqkrTxSdcM+f54Wk9XEoQ30g5GVyOWPMo8VuLyUWysPiSME3IniiK3
gpFivOtWMUld9Q+i2ATPIYfWAKcHMxuWCV6n+dBT9uWuNL01WxIj4mkbUCKPlO08
mlGdIdxoN2oEW3hvQRdF8fvywqbFWnNxPR6yR2O5QjYBXwrbWnyRMTl0Gu2tvIgb
cdKby553QFBe8VNx6tzFyfF3pQltq5GDVTyQ7uAnzdeeGFS73ySez/rP+x7Xy149
+Cc+NhjaFOVW4+j3s4Xz+NdjsgpeBwTqpqtwwhDoLvEkEwGg8mb0fqmI4FuLuzZN
zvdZEt+uLEGj1Aj4jgwoZze2nTowFOu3Eqy+T3tJUwXav6+4gqJ0Qo//x0FRw+E/
M3tBkZyKxzEmIbjKU55y4KkVNcGxeNn4HRXY4fwQpxqHv0zBZ55c1kF+p3ukSwtP
HPDnHqECy0nETWl/iWN0YnigCoeFp7kUfnSS/rh4bXSz7fpU9taNyASS1yU/8cMm
5jsM4q9dKY6hcCzMKMal6KwDayCzi7XYdMxOEpBjnw4uj3DEZz32T5yNOd7udRXh
SuvpwtC/mKS/bdLegUiisEjMXg6oI5r22Pot4o7aX6asrvdzldiYlrUePQpr1oAR
iPeb8STPI4DB2vMh3mnZah/y94gqwEJbh/VkBCYc0T/9hsODyw/6/4zOCk7P9oMr
kJH9KpeQxXrm1rWxDCUBUdFAIFH/17cDIrg58e9a4prweKz+j52wlZInyKKAVOYV
UfPthgIh63hcfltV11Uqw2sJJxLr+SVRFGoLqVBc2mqQaqoZKvwFZiPK3n7Sz8hs
fRTo7UWrE/hlRoD/gOrIHMUPCw4rwiSryu/kLgtrYzw=
`protect END_PROTECTED
