`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8veMZA8xfb0Pmdse+QO9b4gpSkPjgg7ht/V3jYlZxnUElUfo27nxn4tWyBG105P
0WA3Dp+nrJeW63qph2qohMLxdj28eQ1wNReDTFt5w3n/tnHJE101K3cYf2foqQXL
ZD5W45pREznDZpHQybbhd+pnRaV+xofyANpwkPu9uxWfz2i2H/BfJsnyTDj1hMv4
RXcH2teLD8fRu7+sz9UNFZ2K9vuauujskKydDtc5OkbWrxrNqcUNpQkUo0QoeJCr
5cNHCkqQqiVSFpFCVoyZJHzbOgBDgDEje/jWdsmM6pgRNgF4VYTHYmj2fuUa8iWr
gmlSWvoUBh3hRxdABxeilWmPkHcQXYeN/6P//X5Drh+pAGHWn8jOGUK27bnj8X2A
kN1cNSbkwmNBNCU3paGbyupZfOBSbxm/0OHeGa+YFz0HtlJUJ/kg14NxebMklQMD
9tttK0Ki1NDr6Fk8keRj388QFPdRiA1ootOn6MqXAOkFkSnVjbIsT+OYFq3d6k3Z
sVVVfMoDIUJIpmZF7Rj6Iv2DOoNoxtAzA35ZTIIGuzwVvmbcb2aVDHzKRF/h47U7
bRrvDRmk6FLUhIBGy3En//n+QRYioYEXA4Hzsq8EqUqtRlwiUxYuMgdDAsIW2q8P
0eafCtGMjzbJ9achoxIEft3teTjeKtsxE0DJB1rkuJb6HDPAKH0URH8vime2fKYK
JfOdrA3bK+tJhsovoCHIL6WjvvSU21Yoh53Ut0QW9Q4=
`protect END_PROTECTED
