`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LhhbhUBIT2wo+wHFuPdtJG6S7H3IfA/CMGh0Lpm7+cOoe3CJON66yZDFl0IyNSEq
0vIc1carkIYPUuxxjzndXaPFGhABCtlXJVV0HWDQtpnEZFyRKZxJvF15FWLEQjNX
6FeC9YDqPvpt4tqGwWtty1FsKsuqoMt/oK0B0etIZAZPcZsMYpQW7+iNz6dO0Ml2
10RDkwz31dSZBn6O7i0gx0l5WGdSNAEgNNTiO2qYXHD2HrdsvL2yRGd5SaHUkim/
r4JLOUPflY5piMgqvFHTA26W94nQZ+nfNboJKCfxyA6u5g1SLrOujWCX+gCLnENY
w3pGcWZ97QdN8+OhflQZnsPMyFMREGX15qNopSiY1tQ+nYpFq9fxoE6p798uAbB2
fgzKZrYd2TEiKXh2VnNULU8yFVcd95NY11lSUFrMr0W+4B6BlvDsLbuQMVbqLf8d
`protect END_PROTECTED
