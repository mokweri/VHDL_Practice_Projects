`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kt/clL3WHedjAbjIaDxd+TcdDxqJl7fCMpiLzhogxS7y9R5NgKyunwNzp/8dSkeE
xgbn2BMKgZ14a8JR+hRy/EU6LKdNf2K7gkP8LG2HE1d9O2GoYFJzpyR+XLjBKsUt
KW0t9uSXcuUr8a7fFHIohHOicm/oVd/ywN4lX8ANB1YfweqSt0QvuHURfFXNxgYY
K/LaknsiFslvBC5EuKHdWJoNkfWvpSl9DCu+vBmslbkiBlf6HdeZf+VhqvrERdvs
dy1olNdCaVfo4Kuck6FmRlrKzeUnSt7cPRoU+6jUvzf1DOPBVaWbQIbTIBWqhjq0
qgfiU8BrqJgEN2wbkvddr/im5S2IdOFx7tCM6NVSyTtffIi+tLFDmRCSknrdFgUh
MINls8L5c3sHBLZA29DhsBdEt5GFYbK2CtQ2xgZkdJA6MPqLKQtQKxfH5YL3Vphu
vQmWN/a+Zf0OOIa3AQJ28SwhLYBkwaA6qWMI6S8N/litCorLZwwJycsIJP5KbAX+
VmYV4K/MEnylRLFcemakXNsrkHG1kTFwq4l7zk0fZRmbGWf99Z6+paKMQIQ3JAgO
bJQBX7fKMx2J3827X/3uvHHaikdmsp2nIIx1VAu5hea6QVUZIgPUqlpaON2qRPWp
ZPJzRQsVo4W4WdlX8jq301vjbd3y2+Jt8s4nOmM/S+Zts/RBwFmvlnCeLYa9qNYU
x7D8/JL+Csj6dZ9wwOlTWnwH4UaQYCXeZehi3B3uxYSlSHamc7+bl2v1kNAQ/J3g
RkiSyz6R1IchsOTktg4oNpdkmTHCwPKu/8UNFdinvEOy3Lk+V28H7SajtFfTTcj6
UefgD7PKaSGWJGfo6rsjqb09y1+J+msgRAqXeFmk4lZws/X6zKcj4wWTCdkajb1/
+jEdaPZRnK8VdTW6n6NW3vo9G6EQjAK0KgyLhVLbz1NGyBywtrqJrTw7EAdRl9vf
9eCH/xToFcH2RJ+00zbapcrJrYhGtXT6O09jGnrxWjiOFWw3PA/m9zR1nyjgkPzn
EbO7wkYUx7Q0B0yhXj+BUBmUhfZhHUWSNUy56OMvAjqYoabhQk6erRUb0B+O9EFi
eGryjpvbRc71vW5gOhtWiqfWS+qIIgAQGJAPA+ZbjYe94q0JZyyQ7IA2nc8ALKSe
ZFuFHFJxTJ87hkxbNWtFJKTcqvWpD8B7Fta0aSMKG3LTaAW+zRSMpAFF/7o2jJiK
YGBU/z7qYEkB9KCD0dWRUGf1hsPd8S4zG5rGqGWfa12wKxFdO6ihtCbL/APfVui4
fMnwa9oHZNvly/+eTBnJvYpffFMuyRJZ5VGZH497WoRsl5VninKx8ydQgEGqpRKm
ASYrHe4CwaVNQ8t7VM+e61SdZzc9XdsxyaI7GkZA4QrBGp+FyKsoWgWCzCd9vcvx
gDP9WrR/nhJ2Cn9NX3BzVWlaZsdd29EdSJwUuTQ/Wcj1fvC+Ady/F82OWj61ld+A
PJ+GE0uO0/G9Xon+B11L1+s0hiTfsedBQh6bR4xBUNr3Xr1Uwp7id1wx/4E/iBw8
EYZh4ioph2+fZHyvibBMABkYorIqb1PzjZh9LII3JqZQg4KANIlN70wVYGaKYTXg
nC7OLVF2HaqKmBLMxY2CG3A+PwgDlDmysuQ7z5MUAsGUYq/kTAPHpmtpYDz1SNHF
A8/bK8soytQ+TkcPF9jujit+KkWgmPop5OfE+QtlkrMywY4WxXiNLvnEG5O0hrnV
jCQSHk40dJsNMpL9OW4uGpqVYWDkhYNux5PQyhj7wHpAuQaIWr9PlHX1/mAZZsKJ
ggmm6aBUC6nBUliUf+RXWBAqBRFyClr/aM3GtRkRnMzDv7gu45lBvjwXcHGgMvuN
GZj7RKchbf7nuFgq6iOyHk76BlCvVbF2ksokIQbTgBbS6JSW70QfvzHicDLkMtjR
HPI4HbrT1D5BARqf71wyPCc8b1YCWndwhbnWkPhBKl77wrAfQqWU7XmO19PExTKW
bEv3plqE6g4mcVjKD+5i3P7XEWQFUjfz3DyrW+Fr17crlfQVmzVE3bjuJ6wG0Esx
fVcQymiqT2rFkDoYGRb70kkDu8ASB7gLtdu+lWjQL4YzJM4gUCVdTv1s3nW0wsGY
aARiDPm29SMxT+itkYDcl6r4ONiKjUluRHP2nPzS2IJ4ICZVTzmN8u016X4jZ8Px
ehsI5Pl/hi5rLRuC25JctUV/5xT+qM4CxkxdJ/nadVtiWEka0Ut5zeBYGX2i6pFg
HjqiOPLZtdb1SRRVryq5Vw6KcMG55n+Y354WFOmqDFQgbeFCzZdMINRqsNVhC5Wf
pufysEV9cHrPY3TqcDqSUw==
`protect END_PROTECTED
