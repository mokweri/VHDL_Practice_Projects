`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wC+nVcRj4Qji5DU4OCdH2z6lttYjVwv0xPjSrwszaw01mXqi5SOAAh1sCQxGv9Mu
TNklwL17w92B2iupfVtrYht+ky9VeK8zDaabnC7/gX6rlzBRpUnahibOjtCvTgYU
k1UlwpTP4TKVLz7IDH7brUZnwckoMLyk90iawTSr69CtLOFiB3XIw3l/uS/xeTPH
2Np7OrtA56OLxMnxRmYCLC8PNUH1T4ivYbCRscwNXJv91LJ4/bGq/sdKJKw83nVt
WQbXckttes+uv9D7Tt4Y/xF++AwBH9pNxOAQZPQCsafnlwMkfJGFzSMWZ/dJwJvi
VXsB3ro5zga6Wr3N6QKCUdkb2Lo36MbbVE698B3SNrfkvgKW9NLk2NG9SSL3lP/r
lYOesRJ9ezwi/Z4JqVfMaYox0XIPDOxHckuboEC4273dCho88wvLHnATQFaHCbBw
2br/rliqd3L3G3978rs5QDtBpOu/069mlfvHY2lkRWVrwp0jaFQHM7GAuj6rOMNC
mVu0q/RkW5Y4PDZFWHlEHdUUfzZEBypIpQm6lw4F3il0eITjMUmNoLnNqWvPRYi2
iuzPhOyJejT+kQFYUjVXi3eQb/4CvBSXvTN4E2sKuAiGqSgRjNmlRtPR13loVN6d
R3h0QpqGftpyr1Vgi06VpF5QtTt0vpi6LrvtF5dmO/N3yJtwYbUKVCMycWGdbuOr
jjoHcBRNK7pJA6oKioTNk3qR6Egh5ZXn/WWM69XYkRrTMFIai/ud2OtGAgNN5Yfr
YGSOJW8dNYw6IIud7NKZP+GOxNcF2vaxqIZ5ygQ7YHA8rLA8eTk8nXXQdoSHiSSA
4/NMgxVjRvLq1xW1VhIpRFnGEkolh5pYfJ15liThd3Cl/afMKZ1r6CZl7fyQg/sl
iGT0pZmj9jawOoHbSQ99odiuAt6o0RWsutGdK2iL29iUJlAmSJ72OzFxKPuTursU
wTufWopTKi1Ag6YOZq7o31D5M3eI1bXxCGn5H+GZ/THCSkEdCsAd2lXwcy3qGdKK
fDc+kfxp38vcijC0ji+ZFGABwhUjREgoKQGVCcVL9ti8IYZ/yJfeL8ujlcIbGUqz
aPnwp76DoXH937xk0ColPvngWyuanKzOLDUZ2EeIE1415pN9p3nN5Hlj0XQWw0nZ
KLJ4XknAQQVvEdvj/VWLDszBWMLn8VrirKrfuPSw6RHLPLoM7jhimf3feK9HfxCY
bOPGuf2Y/rX70THoEEOo2gHfd5Ld8Bge2NdQXK0owC0nSaBE+jLlR/T4Nn1PcTGQ
U6AKSbg7PoXXwiQ8jXTVDGhuuHuiyj5pQhKrQGCRXZpC13b8ZCtP5uvLAGSzHIe+
1vCgFCSjeDVcx5M/w2Nryw==
`protect END_PROTECTED
