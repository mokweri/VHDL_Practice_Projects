`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3H5hlRAJSHbdO91a6XaLO5xbbMu+djupUfVlAPag5+gxkQewzDqr+TfsmU8CJjNO
/X4A9OvdWb92vwfY/1365EQf0av1Aj13pBlrRNvQh6v4RKOzE033bxVHE7NwikYc
WFqxQWhxR8Vgf9P0cdN1WyKnFpcZn8+pqtcJ1mELUuxz3dpzRgcZrpV80LN/3COJ
jMXb2d8MV1HDRNSdVIBtrri+q+GGVbyRft/3ykv6Eh1+NwW00/yN0Oo06eTOZXnf
2bTD4WPDqFcKW+fk/8NNMbPdUShlEqB1keeEDNizbjS0gL5VhcZnACVxRe9EeyIl
nV/okdLZ2eSJTnbZiID6rOX2R/GKtueTlDLLzpQ2Jr1bvbFUJtDlW/No7mhMfqPY
7PmfYe0D+IR5pLU+wFwkrQWV82X2Vn08CSsgDnz/a7c7JO5YddI3feptWxChkgmh
Rrku04xWtqHgySfoEPm4EwGgmsUQHSE9koQaex/ONGv889cAv7kGDeqKJAx9n0wN
RhpG0O4wPsvPhDnjLPL0H17rduWHkBKKek6lLkn5AQnoIrd1fER31AjBLzrlAXeD
diY+HHq+LtTE9sZEIEf6sec6nKQuBIYRG69XvKXvKtc8O3KToxKIPDkd4DVzbv15
vz3/Z8pnqgrI6gHq8028ua2QOamloHJ3Gc4aIh6Aa5gSjevlxwyaLSb4mV/KixTj
bA4hx70p6X/A5kAJprmHWFNtZTn4RUBp4CzCrvItdxy+cTpuRL4mV5vSkIXcwly8
Vqt4mCLGt47oB9YfmD7IPasygQ0lZQhys1Pc3DCkQNHJgZHdwyj4FJQp8r9MRiSo
hRTg6PWjBNYv2C8hhqnJki97aii5WDKthoOEeJiNerCZ9H1YULxOUO95vcFqRknz
VO99y1cHr5AgxBIzTRtSi6k6UGkrK2Q7BMZ0glLD2dJF9vdB3j2inJEa4owGtjzd
/DT95r3S9o8yvn3K/LMJ4y5Cdb/ANzGolWjAAaG+KGZlP8tMf+fTpKqiBIxg0sQ+
0AQ87rwudlZ8h3WkcHaOo7sTD+fHfmzewucTB21qLo39GdulJJGwq4YWHQpox7Hg
rnad+ra9E9qlu8sw++pTuhXntl2JxJYpvxl6CvXNeDEgXZmxq8AqcgV2rL1uRyfv
yGI7qPciZqx0yrDXqxY35ZRLLVBqfTB0as9Nbnt/9sUBMVLUqW5zQprjjwnqtVV9
3N8/mz21Cu0FzPyir0ndkp2bYcnEYEvgYZVwv4mYqvrjwCSL6XM3x+oXDsoHGjr2
`protect END_PROTECTED
