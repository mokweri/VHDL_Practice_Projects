`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XgYIniXz+Su/SzjRQqCsMpH16Lz8pZ3qlkojZMf73AOxgzNfW/NnpFD3xzY6oE1E
SfM+nmx6aKwoA7nQUNDiwfHj2VyGhpknJ2NXqf44bfxnOGq9b2WlZVaGVLQxjeJW
nT3DzSH8AouVyovBlGBbdOjqwTKB/Vw0GwSGJcpEOZ2BDb9WDeUQo6/FMsQ3cku9
rQ5IV1kP6Amsv6DsA+V75CRy5Eag8flOQoKaoB7Kq15Qzx6KOqXYEwU4TmhyZaYG
3ErQtLmaj/FOsEaxFavI0nNvn5u/YIisI7w7Ztb5bOHhwCp5WcJmGHkv3DR9LCvZ
4WCN/DwkIYJf+ciPJRqZgrFBuaArhRAmdMq0lib79Z4T9p5k4LaM70w/GTUWIaGU
iHS37KkhDTDk+fCkV7SPNcax7oFGrCPlXdn00rvrLuoZE2nVc63h74BG8SsJH0Nf
TJXTMgdMv1FV/TEIPQzXrdyKhQtaontxxL/LIChJg8OtjqfCqnNFuGyqOqP+onfJ
0trU+zGBW/XIhoPuRn16qzEbcGD5SkHlwOtJQYkuNWu6lyJ5UKnal3LAmQsMyHis
i+ohaSy9cNqAE35JXdpGRrMlcUyJppRqXej03qHQC5Y=
`protect END_PROTECTED
