`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nswcfn/UwQaLSqUknSTgCTvktLDJJg5WbHNWvhElK8z4XI04X2ovWW0XlLEsm6at
sFEVoFNTNubzIlr5o2fQyLlVE69H1J2+I/h7zmuqJKFy1mMkPcDLPXDslUbsZaL2
eDAmmdbmkFkpStEc/3UPARuNCboCxGwFn0aMw5PWM70EjTOFhZ0idFmgYSHcjr+J
15lXa6vT1oZ+AFqtDiLN8/D0/Y/cAB+xeLgLBgQgk47GQ6KdkMMdvi7hD4isfzpk
019U84YJ2qZSHImn3xP6j+2tvS68ngARtKIzlTK3vRMW3y5J3D8ZJt2Qv5tgqEtV
Avw3JH6VvnxbSg+9ShasegF7TUVX8ow07Y92DGANJYOFKby7IQB0CXbq9oxp1ev6
nDOgKpHOI1lJy0CNYUkEfTVKBqUoNzTzh5KhGTZiPdI0r3Z7jHGJB21yfOyN/fsB
ppjjZfn2L0h+JPEdYkQIn7S0t5ysZ0O724fNiL0rauTWHsE3udbOowwJjQCsTHnK
2ryg55FJjm1xoLCXOaLLFmakSPpY3fegCxG3mDocV0bxpb+P6pxGPJd+YIAZVneZ
yugPUpHQ/f5hQK0V8I3KgOJB7PPR6CuQMDKP4it+32yvjB8UHQl8MNSiexs12RNF
r+OeToMhaqQN45AV7APxEMmGWqzyiO7OvZkSldvmndPlTKsVh9Mp8jhfSgNdZ0+o
fQjoryinVjcA0KedkGIk29Xp3BejeWcIB/gjXAPbxsv4+yongRY3XdPj5raZOoCl
wo+ZPOIKUd0o2oYIc8gxtDIcPMBoyljroRomjGSoFbflMPr0zsubg5mC00K9pujc
gpdTuceQha7z74TMtnVXgRwbNPikiWscuHtMZgupIwZHFPUr/h+39hp7s6VUoO9n
4eVoQ+aocMdNm/W+MkOaS+AYaORyp3oNG9SgER1pIruHQazLviTCANrPNjIHI+3o
gFsZKeJcZo0II05RFKeRLC92tpHbKeVJ3m1nw9QN9mRP6S/88ZR+kZDK5Pdhd4Tx
UvSnrne8ENHwjIV35SwKaO4I01MJTRbv74mtSp9uqxWkk56jXfhnAOQjUR8OHqJj
LQSDc8f6GkJMRlEsvh462swOaPBaonuqTX+k+VuA12ssjAQ9huu98bIn5yizUiuO
iXV0qsY1Z7v45EChy5a2wRN0IBzOy/DwyeMmBGZZiIWzDScx3sIW5FTqC9Jtul+F
t8MDM/lyUfIsXmz1U8ebUpVzJsDCtnjfNTYtcour97ejAD+8eIMUGYb2HrN+CYjT
m7puViVhVMP83tZel6P6Dvv0/NaO1TA92ZbqjVkVfcY5aQD+o1oJfmnhmZOK46HG
DyqPeSMbHiHunnU9cIk2BtKEB9NeoQU//beolWATFPOL+8acJv8DiGBvF0mFhk2X
uN2Et2fe76kO2cOxnVv3G8+FSV2fL58RX8Okzqor6ToVNgtxiSVV+A2SfW8vbTNg
D5CvVABG8YfWuJ5f91QQQ2swfWhClhZBPfJ70TqkQSIgUH6SINhzkF5o67WB/bwf
V8PpL5jZRBGEMHDgXDpxtuESK56ry6BSoPRw+P0lksrmnjyTy+w2YObfv8AIXNZw
iFvuCwerAY8LcQkG34eLI7bnErPvKCSNy2Ny39h46g1cICXiz05dBior4XKc+Vfu
oLMgk66lqYDYH7Dw5M+5Ks+BdN3YjIDTkglGURRQWwkifxNbChBV3huR/8jFv+X1
mobcYRWCEXi3PQyDg8NGRrF1BctgdolUBDJyew4g4RWNeO/6EKfpJDpW62mdlDGd
X3n5uCq1l5tj9Wuxtj32LIM+/6sL/9xd4PtxT8xRfoIPLW/skIzZlcC2t2BESJQ2
IyRTpci1cwXrfglWKQfiTBYdoO8AduGr1qIMnVJUvZmcOeNNAJfyNMV9WxQrQBRz
EkeZW2UdINImnoPyDfc85o4vXV1wFcPpWDym7+JhXqP4fXAvwqD6xO6pTtE2y9G2
RZv54NRWd5Cs1P2ZyCoiz+5wsFZv1e+5PVGRQMNdKRwHa8OPeoNAwuoINC2ZZ7//
ZomVB63M8Uhr+3wlMvx4w/sfn1emNvc0Lw+XDO5wTieJnrOUhmFqDjcR496GxmyQ
DJ9E7YTtpg2l2bWcMdHud6oN5SLjkehCs0NxA5LfV/TBYEuAqbos0jz0g1NBbsi7
rWtHDcejC8xg2Y9GWiMmMuENh6KiuRUGl3hGPlTKHnAM0AQPrDTvsuunEfWAQYxq
wBgQ0+fBttFORZlNOIRSo2xejiWSOl3FmF5NhFRPrpY8qPPCgJb3bNZvgwu/Ais7
N+4fLx3cwQChPDW85IvPwpGBXMItukBE+2oFTOW5a6UCRYW+Gt+qu9/xTh2yjUmE
0BabXFOdrAjkmLXxMoxgR9nk4LqIzHq3fGrzK8VgnNql35Wu+STI1ROO5WHeqDvQ
JohBCXEGjH7ivc61gWPSXYD7VBkoKlZv2FudsNqWLt1EkpEMjgmaoj95HxVCKnbP
2UaQMssEi66xRBH5JiF/Aa//k2flKrK7kG6VKVd2gAQJ+oQOcPf2VaR47+Uz3ttp
Zkfr3jrevBwN3v6RmZiHmbzNxgye4SP1aP2tXoL/AFWINmE7+2OMFmyeAWn9q76X
xyVOT6oPGYQM0IjOW9Lc0y6CLWbGdz/yBP7FbKjLSuaARlyYNEOsrsmkEGqCqv8D
oScjQncW43lLmd3KaBnckwPOMAQufmIet0Ol1RJbY16JAoHpHe/BnocwIpBoDeHs
58INC1S09YSN9365KsVFPWLjU1MkzgekyHsqmwu74GCFnJPcciSw0HNjMg0C/bUQ
Z+a7B4ymOvKt4JsJeCEE3bA2YEbFrX6SlQa1P22xaeXJL5f1WcVgFWxcmgKlftmV
Fx6ghlh9YsobIX2YWniaST3aaiG2eMU8uaRgJ7ygVfSEheGkeEVzCQ53PgCxSBgC
gxlEPjGCsd/5gXJ6QT2HfDzPVO+NIisi+bDy08tsGsZuj8Dd2QJ+g6WWE3whLjBP
JJyUFOqcCx4HB2WBuJ23Gbxdo3XHUI7N7KSB2Svxmd1VTxgGl2h0SnxWXjTMmZhi
DUIc683kZOpclqEDV+Cj56sJr3Iwp8HlmVcBDxX08k76gCimWDL2i4eHgbgO8V7C
hC8vSv1G3vCru2NDe/K554jHObdQF1RlBPQ1OxckSY2e0H2m2/qPJHxpE+QyF9+3
SvBZeSbZSXu7tjW+CtzwiKGzeHYY78ETVCgBU+9kGSdNTb6yrhOeMopthDrCixM2
OVceTSweAAowwlbT2EUnt+ShDIqVu0zycbL0TbK3ovBypHFBkvrS/i6c4K/WW5mJ
/EIEnTjafWKegIewmYdZVnwQqMBy9CyUBMeAKeZEDf7edCSt3JE73BG8H1w/6qZZ
fOzSDVxdlJZX5fC6bLVdV4baxrbgyhIdThaYWicTRxBmfYghpcpPa4CoWhw7Yvxx
bW3Tc3J147/YP39znMyfk697e1jMaN3u+tn75bJY36bhl6Xq3yjXY2gL2EVbq9om
xuuWKEdfVxHyQ5vRcPFZSurE3foUEYEpBQmVO51+Q8vC+HhnpZcQpj2Wzbm+UTrf
/H470lRQVxjX4S8J3neg2BJUlT4jdfB72JNz3vDSl/HJWB4kiQ6EMQGjMKsnkT1G
4DZtj0+rOn/cAnYd6hdV+D1X0DFlBxD/iZvSYavntajBPMrZwvEEWzBQcfdz2ohG
UmE1pwZZreDDwZ+ahoxjT2bXs7f6SvPSCngnxYURDFZrd1/Y/TNTBYCzrXz2YnHP
iwHOLnnUyrpxWpjTWSfTtp9XbF7c1MpBpJIIZUkilRKyx2/cPIkIoaO8ckmJX1SU
MV6b2lGsH4SK2WtON2iQ7ugYjR6saOMcRq+X5tCaAwn9CR/G5jyHgnpzhjBOSWTk
ZgYrA3yIPue/tmrCCgFWsJLSp8BM5OOXUcmwdpvhPgKp0iOCXvq6XxX7uJWsXT5G
`protect END_PROTECTED
