`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K4AHPFacEYCRPmtRhD63lBXpLvF5mBZbEfa0TgoAAjxFaf1+JvJC3GASZkQ+jyEq
zg0jtNBzNyJmStfDUizdBXRC1bIwF06rXBN7fQ6FOsFcVBOthGbRmFqMk5HcxG/j
E8Pcfwr4RwmCcAFHcQVM4rGilLlO9+DuayuGL5gdZoJEbvwervHNMKdGxEF9zSov
YNTWoOgyxjEIjlCXc8O9AaYJstHe98cIS/PLvR6UmnAB0BxpufHnh1pFwsvO+PEn
8koCHmXrVwu3hmQNT80Gj3P/vttXTxYj7nHx2TTJdLPE8UBq242Als/uctVzq6h2
3PZPp/qlAxBNvHcIPoAdx7al1I47TXuyxOtgel1C8IrnKZrYNAgktBGkcdEP3gvy
LKiucW9lk6dgW9ly5K1j6jNCVcdCHd7rbei5EON6u9kiwOAyT068nZGbRPet9T43
2qcyUVoTuSfOwUbRQDVineGP6izAikeBQIp91S4/YzvmS04KlKU0Ir4cZoNFLZDv
XLzFVKG8Gj3ArK7aQsiwIOMOp4+fpo6+nKnD26LrTZixFwtXcMeRHM3vIAaMYOxh
ZcGBPE0ka6sucS5+VCiynRgDD8GCf9afm0EgKXIhQHzrR0cYhGJFZTkgzsorYsxU
i3S0JzG5xNGj/QgqKbR/0mYjWU+C4n6loCJf80stOi8alNV55eTjYnDa6whtRc2v
ioi3CRgdvHtyg4f65NSUcHRCswvNL6hcVIlTqquWcvXEAu2wBmmt3kEbCiwA41ia
etfaDYDZGdjOXuEHU2i8XnuxkIIQCXsMhvZmkr6dVb8wrarw7T63aR4PRAizRYjz
CC20G9H3Huv9E/OFrVMKlVr2CRKE3VtFk2f3l63cDWGQO3+fbemG2Hvgdb9BE6gt
ahOBBqu0EYEjUsM7Ozodaux0uMLpAdzrs7I+8MpCWAgVTxC7ZQLFwZ45esTAb9ox
/sbR1kjJRlLWT4u1IL31CoZBMzIbaXZczh3uqD203TwrRP05CSDts8FKd5IYumfk
225K+KbNLdqV8zF+WvwB2B+POg3EgYjzKbkDJ4wbUgb+7PTCHEau6LD8kXzkHdph
UL7wZbyA3TsTeOHUwUL3l7Wuby5PTg2JseSHEX610i8YbgEKpq6oKzqTb9CSSd7L
SO4j5LAvnrPyugw5i8ffwowB087VWrWLTg9bFGulAsUJvcDGrctMH2+1YV0Qqd5m
9Qwcu34PNaLycDjbqzBjoupoIkgs22wF7i2EAimxO+5l0pYA1PTQGgYScBBieB67
fOrp7LlpAOuyKLS0NrT9atmptlhubINHT6OsmlMFX13Bhk3H2we0/Y4597CupHeA
mE5IA94plVY2ekv7zvJpxNohp/bXbw1ev7eqZHLFgzT18wJeUxam9NfxkUtuLNNZ
TgQihF69XY5fmn/6HCDv6txcsM2o2q9AIi8F1ntZY4frLmWTtyfZr5hIMMTwi0Xp
LD3Voc7tBRe5x+QCb0kFwXF/CMn+iIapwUz7GWTBmAa6oDb4q0UuisXbIFyCUD2e
pigjB5pVK3wwalfAejl282vKpaA762Cb32saOgLnH9kWBMWHRcYRfR30Lt73A/O7
NVFENkq9SzpznKy7/WAwruvh9FYwOC0kYJ84sXeEvQG7tX8IZ3cwvrw5rvTpYwbr
i5zLAtGc4CjVaTXielJlADP6fcsaMxkZI5Q0TVL6NqirO/A8UAqxTTYvJOSVX87z
2K1PD/rCMcNMvhsiwIg2iQ==
`protect END_PROTECTED
